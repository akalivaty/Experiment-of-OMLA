//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 1 1 1 0 0 1 0 0 0 1 1 0 1 1 0 0 1 0 0 0 1 0 1 1 0 0 1 1 0 1 0 0 1 0 1 1 0 0 0 0 0 0 0 1 1 0 1 1 0 1 0 1 1 0 0 1 0 0 0 1 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:34:31 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n517, new_n518,
    new_n519, new_n520, new_n521, new_n522, new_n523, new_n524, new_n525,
    new_n526, new_n527, new_n528, new_n529, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n536, new_n539, new_n540, new_n541, new_n542,
    new_n543, new_n544, new_n547, new_n548, new_n550, new_n551, new_n552,
    new_n553, new_n554, new_n555, new_n556, new_n557, new_n560, new_n562,
    new_n563, new_n564, new_n566, new_n567, new_n568, new_n569, new_n570,
    new_n571, new_n572, new_n573, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n599, new_n600, new_n603, new_n605,
    new_n606, new_n607, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1152, new_n1153, new_n1154,
    new_n1155, new_n1156, new_n1157, new_n1158, new_n1159, new_n1160,
    new_n1161, new_n1162, new_n1163, new_n1164, new_n1165;
  XOR2_X1   g000(.A(KEYINPUT64), .B(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  XNOR2_X1  g015(.A(KEYINPUT65), .B(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n450), .B(KEYINPUT2), .ZN(new_n451));
  NOR4_X1   g026(.A1(G238), .A2(G237), .A3(G235), .A4(G236), .ZN(new_n452));
  NAND2_X1  g027(.A1(new_n451), .A2(new_n452), .ZN(G261));
  INV_X1    g028(.A(G261), .ZN(G325));
  INV_X1    g029(.A(G567), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n452), .A2(new_n455), .ZN(new_n456));
  NOR2_X1   g031(.A1(new_n456), .A2(KEYINPUT66), .ZN(new_n457));
  AND2_X1   g032(.A1(new_n456), .A2(KEYINPUT66), .ZN(new_n458));
  INV_X1    g033(.A(new_n451), .ZN(new_n459));
  AOI211_X1 g034(.A(new_n457), .B(new_n458), .C1(new_n459), .C2(G2106), .ZN(G319));
  XNOR2_X1  g035(.A(KEYINPUT3), .B(G2104), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n461), .A2(G125), .ZN(new_n462));
  NAND2_X1  g037(.A1(G113), .A2(G2104), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n464), .A2(G2105), .ZN(new_n465));
  NOR2_X1   g040(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n466));
  INV_X1    g041(.A(new_n466), .ZN(new_n467));
  NAND2_X1  g042(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n468));
  AOI21_X1  g043(.A(G2105), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  INV_X1    g044(.A(G2104), .ZN(new_n470));
  NOR2_X1   g045(.A1(new_n470), .A2(G2105), .ZN(new_n471));
  AOI22_X1  g046(.A1(new_n469), .A2(G137), .B1(G101), .B2(new_n471), .ZN(new_n472));
  AND2_X1   g047(.A1(new_n465), .A2(new_n472), .ZN(G160));
  OR2_X1    g048(.A1(G100), .A2(G2105), .ZN(new_n474));
  INV_X1    g049(.A(G2105), .ZN(new_n475));
  OAI211_X1 g050(.A(new_n474), .B(G2104), .C1(G112), .C2(new_n475), .ZN(new_n476));
  XNOR2_X1  g051(.A(new_n476), .B(KEYINPUT69), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n461), .A2(new_n475), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n478), .A2(KEYINPUT67), .ZN(new_n479));
  INV_X1    g054(.A(KEYINPUT67), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n469), .A2(new_n480), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n479), .A2(new_n481), .ZN(new_n482));
  INV_X1    g057(.A(new_n482), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n483), .A2(G136), .ZN(new_n484));
  XOR2_X1   g059(.A(new_n484), .B(KEYINPUT68), .Z(new_n485));
  AOI21_X1  g060(.A(new_n475), .B1(new_n467), .B2(new_n468), .ZN(new_n486));
  AOI211_X1 g061(.A(new_n477), .B(new_n485), .C1(G124), .C2(new_n486), .ZN(G162));
  AND2_X1   g062(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n488));
  OAI211_X1 g063(.A(G138), .B(new_n475), .C1(new_n488), .C2(new_n466), .ZN(new_n489));
  XNOR2_X1  g064(.A(new_n489), .B(KEYINPUT4), .ZN(new_n490));
  INV_X1    g065(.A(KEYINPUT70), .ZN(new_n491));
  NOR2_X1   g066(.A1(new_n475), .A2(G114), .ZN(new_n492));
  OAI21_X1  g067(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n493));
  OAI21_X1  g068(.A(new_n491), .B1(new_n492), .B2(new_n493), .ZN(new_n494));
  OR2_X1    g069(.A1(G102), .A2(G2105), .ZN(new_n495));
  INV_X1    g070(.A(G114), .ZN(new_n496));
  NAND2_X1  g071(.A1(new_n496), .A2(G2105), .ZN(new_n497));
  NAND4_X1  g072(.A1(new_n495), .A2(new_n497), .A3(KEYINPUT70), .A4(G2104), .ZN(new_n498));
  NAND2_X1  g073(.A1(new_n494), .A2(new_n498), .ZN(new_n499));
  NAND3_X1  g074(.A1(new_n461), .A2(G126), .A3(G2105), .ZN(new_n500));
  AND3_X1   g075(.A1(new_n499), .A2(KEYINPUT71), .A3(new_n500), .ZN(new_n501));
  AOI21_X1  g076(.A(KEYINPUT71), .B1(new_n499), .B2(new_n500), .ZN(new_n502));
  OAI21_X1  g077(.A(new_n490), .B1(new_n501), .B2(new_n502), .ZN(new_n503));
  INV_X1    g078(.A(new_n503), .ZN(G164));
  XNOR2_X1  g079(.A(KEYINPUT5), .B(G543), .ZN(new_n505));
  XNOR2_X1  g080(.A(KEYINPUT6), .B(G651), .ZN(new_n506));
  NAND3_X1  g081(.A1(new_n505), .A2(new_n506), .A3(G88), .ZN(new_n507));
  NAND3_X1  g082(.A1(new_n506), .A2(G50), .A3(G543), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  INV_X1    g084(.A(G651), .ZN(new_n510));
  AND2_X1   g085(.A1(KEYINPUT5), .A2(G543), .ZN(new_n511));
  NOR2_X1   g086(.A1(KEYINPUT5), .A2(G543), .ZN(new_n512));
  OAI21_X1  g087(.A(G62), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  NAND2_X1  g088(.A1(G75), .A2(G543), .ZN(new_n514));
  AOI21_X1  g089(.A(new_n510), .B1(new_n513), .B2(new_n514), .ZN(new_n515));
  NOR2_X1   g090(.A1(new_n509), .A2(new_n515), .ZN(G166));
  NAND3_X1  g091(.A1(new_n505), .A2(G63), .A3(G651), .ZN(new_n517));
  AND2_X1   g092(.A1(new_n506), .A2(G543), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n518), .A2(G51), .ZN(new_n519));
  NAND3_X1  g094(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n520));
  XNOR2_X1  g095(.A(new_n520), .B(KEYINPUT7), .ZN(new_n521));
  INV_X1    g096(.A(G89), .ZN(new_n522));
  AND2_X1   g097(.A1(KEYINPUT6), .A2(G651), .ZN(new_n523));
  NOR2_X1   g098(.A1(KEYINPUT6), .A2(G651), .ZN(new_n524));
  OAI22_X1  g099(.A1(new_n512), .A2(new_n511), .B1(new_n523), .B2(new_n524), .ZN(new_n525));
  OAI21_X1  g100(.A(new_n521), .B1(new_n522), .B2(new_n525), .ZN(new_n526));
  INV_X1    g101(.A(KEYINPUT72), .ZN(new_n527));
  OAI211_X1 g102(.A(new_n517), .B(new_n519), .C1(new_n526), .C2(new_n527), .ZN(new_n528));
  AND2_X1   g103(.A1(new_n526), .A2(new_n527), .ZN(new_n529));
  NOR2_X1   g104(.A1(new_n528), .A2(new_n529), .ZN(G168));
  NAND2_X1  g105(.A1(new_n506), .A2(G543), .ZN(new_n531));
  INV_X1    g106(.A(G52), .ZN(new_n532));
  INV_X1    g107(.A(G90), .ZN(new_n533));
  OAI22_X1  g108(.A1(new_n531), .A2(new_n532), .B1(new_n525), .B2(new_n533), .ZN(new_n534));
  XNOR2_X1  g109(.A(new_n534), .B(KEYINPUT73), .ZN(new_n535));
  AOI22_X1  g110(.A1(new_n505), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n536));
  OAI21_X1  g111(.A(new_n535), .B1(new_n510), .B2(new_n536), .ZN(G301));
  INV_X1    g112(.A(G301), .ZN(G171));
  AOI22_X1  g113(.A1(new_n505), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n539));
  NOR2_X1   g114(.A1(new_n539), .A2(new_n510), .ZN(new_n540));
  INV_X1    g115(.A(G43), .ZN(new_n541));
  INV_X1    g116(.A(G81), .ZN(new_n542));
  OAI22_X1  g117(.A1(new_n531), .A2(new_n541), .B1(new_n525), .B2(new_n542), .ZN(new_n543));
  NOR2_X1   g118(.A1(new_n540), .A2(new_n543), .ZN(new_n544));
  NAND2_X1  g119(.A1(new_n544), .A2(G860), .ZN(G153));
  NAND4_X1  g120(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g121(.A1(G1), .A2(G3), .ZN(new_n547));
  XNOR2_X1  g122(.A(new_n547), .B(KEYINPUT8), .ZN(new_n548));
  NAND4_X1  g123(.A1(G319), .A2(G483), .A3(G661), .A4(new_n548), .ZN(G188));
  INV_X1    g124(.A(new_n525), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n550), .A2(G91), .ZN(new_n551));
  AOI22_X1  g126(.A1(new_n505), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n518), .A2(G53), .ZN(new_n553));
  AND2_X1   g128(.A1(new_n553), .A2(KEYINPUT9), .ZN(new_n554));
  NOR2_X1   g129(.A1(new_n553), .A2(KEYINPUT9), .ZN(new_n555));
  OAI221_X1 g130(.A(new_n551), .B1(new_n510), .B2(new_n552), .C1(new_n554), .C2(new_n555), .ZN(new_n556));
  INV_X1    g131(.A(KEYINPUT74), .ZN(new_n557));
  XNOR2_X1  g132(.A(new_n556), .B(new_n557), .ZN(G299));
  INV_X1    g133(.A(G168), .ZN(G286));
  AOI22_X1  g134(.A1(new_n505), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n560));
  OAI211_X1 g135(.A(new_n507), .B(new_n508), .C1(new_n560), .C2(new_n510), .ZN(G303));
  NAND2_X1  g136(.A1(new_n518), .A2(G49), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n550), .A2(G87), .ZN(new_n563));
  OAI21_X1  g138(.A(G651), .B1(new_n505), .B2(G74), .ZN(new_n564));
  NAND3_X1  g139(.A1(new_n562), .A2(new_n563), .A3(new_n564), .ZN(G288));
  INV_X1    g140(.A(G48), .ZN(new_n566));
  INV_X1    g141(.A(G86), .ZN(new_n567));
  OAI22_X1  g142(.A1(new_n531), .A2(new_n566), .B1(new_n525), .B2(new_n567), .ZN(new_n568));
  NAND2_X1  g143(.A1(new_n505), .A2(G61), .ZN(new_n569));
  NAND2_X1  g144(.A1(G73), .A2(G543), .ZN(new_n570));
  XNOR2_X1  g145(.A(new_n570), .B(KEYINPUT75), .ZN(new_n571));
  AOI21_X1  g146(.A(new_n510), .B1(new_n569), .B2(new_n571), .ZN(new_n572));
  NOR2_X1   g147(.A1(new_n568), .A2(new_n572), .ZN(new_n573));
  INV_X1    g148(.A(new_n573), .ZN(G305));
  AND2_X1   g149(.A1(new_n505), .A2(G60), .ZN(new_n575));
  AND2_X1   g150(.A1(G72), .A2(G543), .ZN(new_n576));
  OAI21_X1  g151(.A(G651), .B1(new_n575), .B2(new_n576), .ZN(new_n577));
  INV_X1    g152(.A(KEYINPUT76), .ZN(new_n578));
  NAND2_X1  g153(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  AOI22_X1  g154(.A1(G47), .A2(new_n518), .B1(new_n550), .B2(G85), .ZN(new_n580));
  AND2_X1   g155(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  OR2_X1    g156(.A1(new_n577), .A2(new_n578), .ZN(new_n582));
  NAND2_X1  g157(.A1(new_n581), .A2(new_n582), .ZN(G290));
  NAND2_X1  g158(.A1(G301), .A2(G868), .ZN(new_n584));
  NAND2_X1  g159(.A1(new_n505), .A2(G66), .ZN(new_n585));
  NAND2_X1  g160(.A1(G79), .A2(G543), .ZN(new_n586));
  AOI21_X1  g161(.A(new_n510), .B1(new_n585), .B2(new_n586), .ZN(new_n587));
  NAND2_X1  g162(.A1(new_n518), .A2(G54), .ZN(new_n588));
  INV_X1    g163(.A(new_n588), .ZN(new_n589));
  NAND2_X1  g164(.A1(new_n550), .A2(G92), .ZN(new_n590));
  XNOR2_X1  g165(.A(new_n590), .B(KEYINPUT77), .ZN(new_n591));
  INV_X1    g166(.A(KEYINPUT10), .ZN(new_n592));
  AOI211_X1 g167(.A(new_n587), .B(new_n589), .C1(new_n591), .C2(new_n592), .ZN(new_n593));
  OR2_X1    g168(.A1(new_n591), .A2(new_n592), .ZN(new_n594));
  NAND2_X1  g169(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  INV_X1    g170(.A(new_n595), .ZN(new_n596));
  OAI21_X1  g171(.A(new_n584), .B1(new_n596), .B2(G868), .ZN(G284));
  OAI21_X1  g172(.A(new_n584), .B1(new_n596), .B2(G868), .ZN(G321));
  NAND2_X1  g173(.A1(G286), .A2(G868), .ZN(new_n599));
  XNOR2_X1  g174(.A(new_n556), .B(KEYINPUT74), .ZN(new_n600));
  OAI21_X1  g175(.A(new_n599), .B1(new_n600), .B2(G868), .ZN(G297));
  OAI21_X1  g176(.A(new_n599), .B1(new_n600), .B2(G868), .ZN(G280));
  INV_X1    g177(.A(G559), .ZN(new_n603));
  OAI21_X1  g178(.A(new_n596), .B1(new_n603), .B2(G860), .ZN(G148));
  NOR2_X1   g179(.A1(new_n544), .A2(G868), .ZN(new_n605));
  NAND2_X1  g180(.A1(new_n596), .A2(new_n603), .ZN(new_n606));
  AOI21_X1  g181(.A(new_n605), .B1(new_n606), .B2(G868), .ZN(new_n607));
  XOR2_X1   g182(.A(new_n607), .B(KEYINPUT78), .Z(G323));
  XNOR2_X1  g183(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g184(.A1(new_n461), .A2(new_n471), .ZN(new_n610));
  XNOR2_X1  g185(.A(new_n610), .B(KEYINPUT12), .ZN(new_n611));
  XNOR2_X1  g186(.A(KEYINPUT79), .B(KEYINPUT13), .ZN(new_n612));
  XNOR2_X1  g187(.A(new_n611), .B(new_n612), .ZN(new_n613));
  INV_X1    g188(.A(G2100), .ZN(new_n614));
  OR2_X1    g189(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  NAND2_X1  g190(.A1(new_n483), .A2(G135), .ZN(new_n616));
  INV_X1    g191(.A(G2096), .ZN(new_n617));
  OR2_X1    g192(.A1(new_n475), .A2(G111), .ZN(new_n618));
  OR2_X1    g193(.A1(new_n618), .A2(KEYINPUT80), .ZN(new_n619));
  OAI21_X1  g194(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n620));
  AOI21_X1  g195(.A(new_n620), .B1(new_n618), .B2(KEYINPUT80), .ZN(new_n621));
  AOI22_X1  g196(.A1(new_n619), .A2(new_n621), .B1(new_n486), .B2(G123), .ZN(new_n622));
  NAND3_X1  g197(.A1(new_n616), .A2(new_n617), .A3(new_n622), .ZN(new_n623));
  NAND2_X1  g198(.A1(new_n613), .A2(new_n614), .ZN(new_n624));
  NAND2_X1  g199(.A1(new_n616), .A2(new_n622), .ZN(new_n625));
  NAND2_X1  g200(.A1(new_n625), .A2(G2096), .ZN(new_n626));
  NAND4_X1  g201(.A1(new_n615), .A2(new_n623), .A3(new_n624), .A4(new_n626), .ZN(G156));
  INV_X1    g202(.A(G14), .ZN(new_n628));
  XNOR2_X1  g203(.A(G2427), .B(G2438), .ZN(new_n629));
  XNOR2_X1  g204(.A(new_n629), .B(G2430), .ZN(new_n630));
  XNOR2_X1  g205(.A(KEYINPUT15), .B(G2435), .ZN(new_n631));
  OR2_X1    g206(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  NAND2_X1  g207(.A1(new_n630), .A2(new_n631), .ZN(new_n633));
  NAND3_X1  g208(.A1(new_n632), .A2(KEYINPUT14), .A3(new_n633), .ZN(new_n634));
  XNOR2_X1  g209(.A(new_n634), .B(KEYINPUT82), .ZN(new_n635));
  INV_X1    g210(.A(G1341), .ZN(new_n636));
  XNOR2_X1  g211(.A(new_n635), .B(new_n636), .ZN(new_n637));
  XNOR2_X1  g212(.A(new_n637), .B(G1348), .ZN(new_n638));
  XOR2_X1   g213(.A(G2451), .B(G2454), .Z(new_n639));
  XNOR2_X1  g214(.A(G2443), .B(G2446), .ZN(new_n640));
  XNOR2_X1  g215(.A(new_n639), .B(new_n640), .ZN(new_n641));
  XNOR2_X1  g216(.A(KEYINPUT81), .B(KEYINPUT16), .ZN(new_n642));
  XOR2_X1   g217(.A(new_n641), .B(new_n642), .Z(new_n643));
  AOI21_X1  g218(.A(new_n628), .B1(new_n638), .B2(new_n643), .ZN(new_n644));
  OAI211_X1 g219(.A(new_n644), .B(KEYINPUT83), .C1(new_n643), .C2(new_n638), .ZN(new_n645));
  INV_X1    g220(.A(KEYINPUT83), .ZN(new_n646));
  INV_X1    g221(.A(G1348), .ZN(new_n647));
  XNOR2_X1  g222(.A(new_n637), .B(new_n647), .ZN(new_n648));
  INV_X1    g223(.A(new_n643), .ZN(new_n649));
  OAI21_X1  g224(.A(G14), .B1(new_n648), .B2(new_n649), .ZN(new_n650));
  NOR2_X1   g225(.A1(new_n638), .A2(new_n643), .ZN(new_n651));
  OAI21_X1  g226(.A(new_n646), .B1(new_n650), .B2(new_n651), .ZN(new_n652));
  NAND2_X1  g227(.A1(new_n645), .A2(new_n652), .ZN(new_n653));
  INV_X1    g228(.A(new_n653), .ZN(G401));
  INV_X1    g229(.A(KEYINPUT18), .ZN(new_n655));
  XOR2_X1   g230(.A(G2084), .B(G2090), .Z(new_n656));
  XNOR2_X1  g231(.A(G2067), .B(G2678), .ZN(new_n657));
  NAND2_X1  g232(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  NAND2_X1  g233(.A1(new_n658), .A2(KEYINPUT17), .ZN(new_n659));
  NOR2_X1   g234(.A1(new_n656), .A2(new_n657), .ZN(new_n660));
  OAI21_X1  g235(.A(new_n655), .B1(new_n659), .B2(new_n660), .ZN(new_n661));
  XNOR2_X1  g236(.A(new_n661), .B(new_n614), .ZN(new_n662));
  XOR2_X1   g237(.A(G2072), .B(G2078), .Z(new_n663));
  AOI21_X1  g238(.A(new_n663), .B1(new_n658), .B2(KEYINPUT18), .ZN(new_n664));
  XNOR2_X1  g239(.A(new_n664), .B(new_n617), .ZN(new_n665));
  XNOR2_X1  g240(.A(new_n662), .B(new_n665), .ZN(G227));
  XOR2_X1   g241(.A(G1971), .B(G1976), .Z(new_n667));
  XNOR2_X1  g242(.A(new_n667), .B(KEYINPUT19), .ZN(new_n668));
  XNOR2_X1  g243(.A(G1956), .B(G2474), .ZN(new_n669));
  XNOR2_X1  g244(.A(G1961), .B(G1966), .ZN(new_n670));
  NOR2_X1   g245(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  AND2_X1   g246(.A1(new_n669), .A2(new_n670), .ZN(new_n672));
  NOR3_X1   g247(.A1(new_n668), .A2(new_n671), .A3(new_n672), .ZN(new_n673));
  NAND2_X1  g248(.A1(new_n668), .A2(new_n671), .ZN(new_n674));
  XNOR2_X1  g249(.A(KEYINPUT84), .B(KEYINPUT20), .ZN(new_n675));
  XNOR2_X1  g250(.A(new_n674), .B(new_n675), .ZN(new_n676));
  AOI211_X1 g251(.A(new_n673), .B(new_n676), .C1(new_n668), .C2(new_n672), .ZN(new_n677));
  XNOR2_X1  g252(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n678));
  XNOR2_X1  g253(.A(new_n677), .B(new_n678), .ZN(new_n679));
  XOR2_X1   g254(.A(G1991), .B(G1996), .Z(new_n680));
  XNOR2_X1  g255(.A(new_n679), .B(new_n680), .ZN(new_n681));
  XNOR2_X1  g256(.A(G1981), .B(G1986), .ZN(new_n682));
  XNOR2_X1  g257(.A(new_n681), .B(new_n682), .ZN(G229));
  NOR2_X1   g258(.A1(G25), .A2(G29), .ZN(new_n684));
  NAND2_X1  g259(.A1(new_n483), .A2(G131), .ZN(new_n685));
  NOR2_X1   g260(.A1(G95), .A2(G2105), .ZN(new_n686));
  XNOR2_X1  g261(.A(new_n686), .B(KEYINPUT85), .ZN(new_n687));
  INV_X1    g262(.A(G107), .ZN(new_n688));
  AOI21_X1  g263(.A(new_n470), .B1(new_n688), .B2(G2105), .ZN(new_n689));
  AOI22_X1  g264(.A1(new_n687), .A2(new_n689), .B1(new_n486), .B2(G119), .ZN(new_n690));
  AND2_X1   g265(.A1(new_n685), .A2(new_n690), .ZN(new_n691));
  AOI21_X1  g266(.A(new_n684), .B1(new_n691), .B2(G29), .ZN(new_n692));
  XNOR2_X1  g267(.A(new_n692), .B(KEYINPUT86), .ZN(new_n693));
  XOR2_X1   g268(.A(KEYINPUT35), .B(G1991), .Z(new_n694));
  XOR2_X1   g269(.A(new_n693), .B(new_n694), .Z(new_n695));
  INV_X1    g270(.A(G1986), .ZN(new_n696));
  INV_X1    g271(.A(G16), .ZN(new_n697));
  NAND2_X1  g272(.A1(new_n697), .A2(G24), .ZN(new_n698));
  INV_X1    g273(.A(G290), .ZN(new_n699));
  OAI21_X1  g274(.A(new_n698), .B1(new_n699), .B2(new_n697), .ZN(new_n700));
  XNOR2_X1  g275(.A(new_n700), .B(KEYINPUT87), .ZN(new_n701));
  AOI21_X1  g276(.A(new_n695), .B1(new_n696), .B2(new_n701), .ZN(new_n702));
  NOR2_X1   g277(.A1(G6), .A2(G16), .ZN(new_n703));
  AOI21_X1  g278(.A(new_n703), .B1(new_n573), .B2(G16), .ZN(new_n704));
  XNOR2_X1  g279(.A(new_n704), .B(KEYINPUT32), .ZN(new_n705));
  INV_X1    g280(.A(G1981), .ZN(new_n706));
  XNOR2_X1  g281(.A(new_n705), .B(new_n706), .ZN(new_n707));
  OR2_X1    g282(.A1(G16), .A2(G23), .ZN(new_n708));
  INV_X1    g283(.A(new_n563), .ZN(new_n709));
  INV_X1    g284(.A(G49), .ZN(new_n710));
  OAI21_X1  g285(.A(new_n564), .B1(new_n710), .B2(new_n531), .ZN(new_n711));
  OAI21_X1  g286(.A(KEYINPUT88), .B1(new_n709), .B2(new_n711), .ZN(new_n712));
  INV_X1    g287(.A(KEYINPUT88), .ZN(new_n713));
  NAND4_X1  g288(.A1(new_n562), .A2(new_n563), .A3(new_n713), .A4(new_n564), .ZN(new_n714));
  NAND2_X1  g289(.A1(new_n712), .A2(new_n714), .ZN(new_n715));
  OAI21_X1  g290(.A(new_n708), .B1(new_n715), .B2(new_n697), .ZN(new_n716));
  XNOR2_X1  g291(.A(KEYINPUT33), .B(G1976), .ZN(new_n717));
  XNOR2_X1  g292(.A(new_n717), .B(KEYINPUT89), .ZN(new_n718));
  NAND2_X1  g293(.A1(new_n716), .A2(new_n718), .ZN(new_n719));
  OR2_X1    g294(.A1(new_n716), .A2(new_n718), .ZN(new_n720));
  NAND2_X1  g295(.A1(new_n697), .A2(G22), .ZN(new_n721));
  XOR2_X1   g296(.A(new_n721), .B(KEYINPUT90), .Z(new_n722));
  OAI21_X1  g297(.A(new_n722), .B1(G166), .B2(new_n697), .ZN(new_n723));
  INV_X1    g298(.A(G1971), .ZN(new_n724));
  XNOR2_X1  g299(.A(new_n723), .B(new_n724), .ZN(new_n725));
  NAND4_X1  g300(.A1(new_n707), .A2(new_n719), .A3(new_n720), .A4(new_n725), .ZN(new_n726));
  NAND2_X1  g301(.A1(new_n726), .A2(KEYINPUT34), .ZN(new_n727));
  OR2_X1    g302(.A1(new_n726), .A2(KEYINPUT34), .ZN(new_n728));
  OR2_X1    g303(.A1(new_n701), .A2(new_n696), .ZN(new_n729));
  NAND4_X1  g304(.A1(new_n702), .A2(new_n727), .A3(new_n728), .A4(new_n729), .ZN(new_n730));
  XNOR2_X1  g305(.A(new_n730), .B(KEYINPUT36), .ZN(new_n731));
  AND2_X1   g306(.A1(new_n483), .A2(G139), .ZN(new_n732));
  NAND3_X1  g307(.A1(new_n475), .A2(G103), .A3(G2104), .ZN(new_n733));
  XOR2_X1   g308(.A(new_n733), .B(KEYINPUT25), .Z(new_n734));
  AOI22_X1  g309(.A1(new_n461), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n735));
  OAI21_X1  g310(.A(new_n734), .B1(new_n735), .B2(new_n475), .ZN(new_n736));
  NOR2_X1   g311(.A1(new_n732), .A2(new_n736), .ZN(new_n737));
  INV_X1    g312(.A(G29), .ZN(new_n738));
  NOR2_X1   g313(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  AOI21_X1  g314(.A(new_n739), .B1(new_n738), .B2(G33), .ZN(new_n740));
  INV_X1    g315(.A(G2072), .ZN(new_n741));
  NAND2_X1  g316(.A1(new_n483), .A2(G141), .ZN(new_n742));
  AND2_X1   g317(.A1(new_n471), .A2(G105), .ZN(new_n743));
  NAND3_X1  g318(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n744));
  XNOR2_X1  g319(.A(new_n744), .B(KEYINPUT26), .ZN(new_n745));
  AOI211_X1 g320(.A(new_n743), .B(new_n745), .C1(G129), .C2(new_n486), .ZN(new_n746));
  NAND2_X1  g321(.A1(new_n742), .A2(new_n746), .ZN(new_n747));
  INV_X1    g322(.A(new_n747), .ZN(new_n748));
  NOR2_X1   g323(.A1(new_n748), .A2(new_n738), .ZN(new_n749));
  AOI21_X1  g324(.A(new_n749), .B1(new_n738), .B2(G32), .ZN(new_n750));
  XNOR2_X1  g325(.A(KEYINPUT27), .B(G1996), .ZN(new_n751));
  AOI22_X1  g326(.A1(new_n740), .A2(new_n741), .B1(new_n750), .B2(new_n751), .ZN(new_n752));
  OAI21_X1  g327(.A(new_n752), .B1(new_n741), .B2(new_n740), .ZN(new_n753));
  NAND2_X1  g328(.A1(new_n697), .A2(G19), .ZN(new_n754));
  OAI21_X1  g329(.A(new_n754), .B1(new_n544), .B2(new_n697), .ZN(new_n755));
  XNOR2_X1  g330(.A(new_n755), .B(new_n636), .ZN(new_n756));
  XOR2_X1   g331(.A(KEYINPUT93), .B(KEYINPUT24), .Z(new_n757));
  NOR2_X1   g332(.A1(new_n757), .A2(G34), .ZN(new_n758));
  NOR2_X1   g333(.A1(new_n758), .A2(G29), .ZN(new_n759));
  OR2_X1    g334(.A1(new_n759), .A2(KEYINPUT94), .ZN(new_n760));
  AOI22_X1  g335(.A1(new_n759), .A2(KEYINPUT94), .B1(G34), .B2(new_n757), .ZN(new_n761));
  AOI22_X1  g336(.A1(new_n760), .A2(new_n761), .B1(G160), .B2(G29), .ZN(new_n762));
  OAI21_X1  g337(.A(new_n756), .B1(G2084), .B2(new_n762), .ZN(new_n763));
  NOR2_X1   g338(.A1(new_n750), .A2(new_n751), .ZN(new_n764));
  NAND2_X1  g339(.A1(new_n762), .A2(G2084), .ZN(new_n765));
  XOR2_X1   g340(.A(KEYINPUT31), .B(G11), .Z(new_n766));
  INV_X1    g341(.A(G28), .ZN(new_n767));
  OR2_X1    g342(.A1(new_n767), .A2(KEYINPUT30), .ZN(new_n768));
  AOI21_X1  g343(.A(G29), .B1(new_n767), .B2(KEYINPUT30), .ZN(new_n769));
  AOI21_X1  g344(.A(new_n766), .B1(new_n768), .B2(new_n769), .ZN(new_n770));
  OAI211_X1 g345(.A(new_n765), .B(new_n770), .C1(new_n738), .C2(new_n625), .ZN(new_n771));
  NOR4_X1   g346(.A1(new_n753), .A2(new_n763), .A3(new_n764), .A4(new_n771), .ZN(new_n772));
  NOR2_X1   g347(.A1(G29), .A2(G35), .ZN(new_n773));
  AOI21_X1  g348(.A(new_n773), .B1(G162), .B2(G29), .ZN(new_n774));
  XOR2_X1   g349(.A(KEYINPUT29), .B(G2090), .Z(new_n775));
  XNOR2_X1  g350(.A(new_n774), .B(new_n775), .ZN(new_n776));
  NAND2_X1  g351(.A1(new_n697), .A2(G4), .ZN(new_n777));
  OAI21_X1  g352(.A(new_n777), .B1(new_n596), .B2(new_n697), .ZN(new_n778));
  XNOR2_X1  g353(.A(new_n778), .B(new_n647), .ZN(new_n779));
  NAND2_X1  g354(.A1(new_n697), .A2(G5), .ZN(new_n780));
  OAI21_X1  g355(.A(new_n780), .B1(G171), .B2(new_n697), .ZN(new_n781));
  NOR2_X1   g356(.A1(new_n781), .A2(G1961), .ZN(new_n782));
  AND2_X1   g357(.A1(new_n781), .A2(G1961), .ZN(new_n783));
  NAND2_X1  g358(.A1(new_n697), .A2(G21), .ZN(new_n784));
  OAI21_X1  g359(.A(new_n784), .B1(G168), .B2(new_n697), .ZN(new_n785));
  AOI211_X1 g360(.A(new_n782), .B(new_n783), .C1(G1966), .C2(new_n785), .ZN(new_n786));
  NAND4_X1  g361(.A1(new_n772), .A2(new_n776), .A3(new_n779), .A4(new_n786), .ZN(new_n787));
  NAND2_X1  g362(.A1(new_n697), .A2(G20), .ZN(new_n788));
  XNOR2_X1  g363(.A(new_n788), .B(KEYINPUT23), .ZN(new_n789));
  OAI21_X1  g364(.A(new_n789), .B1(new_n600), .B2(new_n697), .ZN(new_n790));
  XOR2_X1   g365(.A(new_n790), .B(G1956), .Z(new_n791));
  NAND2_X1  g366(.A1(new_n738), .A2(G27), .ZN(new_n792));
  XOR2_X1   g367(.A(new_n792), .B(KEYINPUT96), .Z(new_n793));
  OAI21_X1  g368(.A(new_n793), .B1(G164), .B2(new_n738), .ZN(new_n794));
  INV_X1    g369(.A(G2078), .ZN(new_n795));
  XNOR2_X1  g370(.A(new_n794), .B(new_n795), .ZN(new_n796));
  NOR2_X1   g371(.A1(new_n785), .A2(G1966), .ZN(new_n797));
  XOR2_X1   g372(.A(new_n797), .B(KEYINPUT95), .Z(new_n798));
  NAND2_X1  g373(.A1(new_n738), .A2(G26), .ZN(new_n799));
  XOR2_X1   g374(.A(new_n799), .B(KEYINPUT92), .Z(new_n800));
  XNOR2_X1  g375(.A(new_n800), .B(KEYINPUT28), .ZN(new_n801));
  OAI21_X1  g376(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n802));
  INV_X1    g377(.A(G116), .ZN(new_n803));
  AOI21_X1  g378(.A(new_n802), .B1(new_n803), .B2(G2105), .ZN(new_n804));
  AOI21_X1  g379(.A(new_n804), .B1(new_n486), .B2(G128), .ZN(new_n805));
  INV_X1    g380(.A(G140), .ZN(new_n806));
  OAI21_X1  g381(.A(new_n805), .B1(new_n482), .B2(new_n806), .ZN(new_n807));
  XNOR2_X1  g382(.A(new_n807), .B(KEYINPUT91), .ZN(new_n808));
  INV_X1    g383(.A(new_n808), .ZN(new_n809));
  AOI21_X1  g384(.A(new_n801), .B1(new_n809), .B2(G29), .ZN(new_n810));
  XNOR2_X1  g385(.A(new_n810), .B(G2067), .ZN(new_n811));
  NAND4_X1  g386(.A1(new_n791), .A2(new_n796), .A3(new_n798), .A4(new_n811), .ZN(new_n812));
  NOR2_X1   g387(.A1(new_n787), .A2(new_n812), .ZN(new_n813));
  NAND2_X1  g388(.A1(new_n731), .A2(new_n813), .ZN(G150));
  XNOR2_X1  g389(.A(G150), .B(KEYINPUT97), .ZN(G311));
  NAND2_X1  g390(.A1(new_n596), .A2(G559), .ZN(new_n816));
  XNOR2_X1  g391(.A(new_n816), .B(KEYINPUT38), .ZN(new_n817));
  AOI22_X1  g392(.A1(G55), .A2(new_n518), .B1(new_n550), .B2(G93), .ZN(new_n818));
  AOI22_X1  g393(.A1(new_n505), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n819));
  OAI21_X1  g394(.A(new_n818), .B1(new_n510), .B2(new_n819), .ZN(new_n820));
  INV_X1    g395(.A(new_n544), .ZN(new_n821));
  XNOR2_X1  g396(.A(new_n820), .B(new_n821), .ZN(new_n822));
  XOR2_X1   g397(.A(new_n817), .B(new_n822), .Z(new_n823));
  AND2_X1   g398(.A1(new_n823), .A2(KEYINPUT39), .ZN(new_n824));
  NOR2_X1   g399(.A1(new_n823), .A2(KEYINPUT39), .ZN(new_n825));
  NOR3_X1   g400(.A1(new_n824), .A2(new_n825), .A3(G860), .ZN(new_n826));
  NAND2_X1  g401(.A1(new_n820), .A2(G860), .ZN(new_n827));
  XNOR2_X1  g402(.A(new_n827), .B(KEYINPUT37), .ZN(new_n828));
  OR2_X1    g403(.A1(new_n826), .A2(new_n828), .ZN(G145));
  NAND2_X1  g404(.A1(new_n486), .A2(G130), .ZN(new_n830));
  NOR2_X1   g405(.A1(new_n475), .A2(G118), .ZN(new_n831));
  OAI21_X1  g406(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n832));
  OAI21_X1  g407(.A(new_n830), .B1(new_n831), .B2(new_n832), .ZN(new_n833));
  AOI21_X1  g408(.A(new_n833), .B1(new_n483), .B2(G142), .ZN(new_n834));
  XOR2_X1   g409(.A(new_n834), .B(new_n611), .Z(new_n835));
  XNOR2_X1  g410(.A(new_n835), .B(new_n691), .ZN(new_n836));
  INV_X1    g411(.A(new_n836), .ZN(new_n837));
  XNOR2_X1  g412(.A(new_n808), .B(KEYINPUT98), .ZN(new_n838));
  XNOR2_X1  g413(.A(new_n838), .B(new_n748), .ZN(new_n839));
  AOI22_X1  g414(.A1(G126), .A2(new_n486), .B1(new_n494), .B2(new_n498), .ZN(new_n840));
  NAND2_X1  g415(.A1(new_n490), .A2(new_n840), .ZN(new_n841));
  OR2_X1    g416(.A1(new_n839), .A2(new_n841), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n839), .A2(new_n841), .ZN(new_n843));
  INV_X1    g418(.A(new_n737), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n844), .A2(KEYINPUT99), .ZN(new_n845));
  NAND3_X1  g420(.A1(new_n842), .A2(new_n843), .A3(new_n845), .ZN(new_n846));
  NOR2_X1   g421(.A1(new_n844), .A2(KEYINPUT99), .ZN(new_n847));
  NAND2_X1  g422(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  INV_X1    g423(.A(new_n848), .ZN(new_n849));
  NOR2_X1   g424(.A1(new_n846), .A2(new_n847), .ZN(new_n850));
  OAI21_X1  g425(.A(new_n837), .B1(new_n849), .B2(new_n850), .ZN(new_n851));
  OR2_X1    g426(.A1(new_n846), .A2(new_n847), .ZN(new_n852));
  NAND3_X1  g427(.A1(new_n852), .A2(new_n848), .A3(new_n836), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n851), .A2(new_n853), .ZN(new_n854));
  XNOR2_X1  g429(.A(new_n625), .B(G160), .ZN(new_n855));
  XNOR2_X1  g430(.A(G162), .B(new_n855), .ZN(new_n856));
  INV_X1    g431(.A(new_n856), .ZN(new_n857));
  NAND2_X1  g432(.A1(new_n854), .A2(new_n857), .ZN(new_n858));
  INV_X1    g433(.A(G37), .ZN(new_n859));
  NAND3_X1  g434(.A1(new_n851), .A2(new_n856), .A3(new_n853), .ZN(new_n860));
  NAND3_X1  g435(.A1(new_n858), .A2(new_n859), .A3(new_n860), .ZN(new_n861));
  XNOR2_X1  g436(.A(new_n861), .B(KEYINPUT40), .ZN(G395));
  XNOR2_X1  g437(.A(new_n573), .B(G303), .ZN(new_n863));
  XOR2_X1   g438(.A(G290), .B(new_n715), .Z(new_n864));
  OAI21_X1  g439(.A(new_n863), .B1(new_n864), .B2(KEYINPUT101), .ZN(new_n865));
  NAND2_X1  g440(.A1(new_n864), .A2(KEYINPUT101), .ZN(new_n866));
  XNOR2_X1  g441(.A(new_n865), .B(new_n866), .ZN(new_n867));
  XNOR2_X1  g442(.A(new_n867), .B(KEYINPUT42), .ZN(new_n868));
  XOR2_X1   g443(.A(new_n606), .B(new_n822), .Z(new_n869));
  NAND2_X1  g444(.A1(new_n596), .A2(G299), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n600), .A2(new_n595), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  NOR2_X1   g447(.A1(new_n869), .A2(new_n872), .ZN(new_n873));
  INV_X1    g448(.A(KEYINPUT41), .ZN(new_n874));
  NAND2_X1  g449(.A1(new_n872), .A2(new_n874), .ZN(new_n875));
  NAND3_X1  g450(.A1(new_n870), .A2(new_n871), .A3(KEYINPUT41), .ZN(new_n876));
  NAND3_X1  g451(.A1(new_n875), .A2(KEYINPUT100), .A3(new_n876), .ZN(new_n877));
  OR3_X1    g452(.A1(new_n872), .A2(KEYINPUT100), .A3(new_n874), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n877), .A2(new_n878), .ZN(new_n879));
  AOI21_X1  g454(.A(new_n873), .B1(new_n869), .B2(new_n879), .ZN(new_n880));
  OR2_X1    g455(.A1(new_n868), .A2(new_n880), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n868), .A2(new_n880), .ZN(new_n882));
  NAND3_X1  g457(.A1(new_n881), .A2(G868), .A3(new_n882), .ZN(new_n883));
  INV_X1    g458(.A(KEYINPUT102), .ZN(new_n884));
  NOR2_X1   g459(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  INV_X1    g460(.A(G868), .ZN(new_n886));
  AOI21_X1  g461(.A(KEYINPUT102), .B1(new_n820), .B2(new_n886), .ZN(new_n887));
  AOI21_X1  g462(.A(new_n885), .B1(new_n883), .B2(new_n887), .ZN(G295));
  AOI21_X1  g463(.A(new_n885), .B1(new_n883), .B2(new_n887), .ZN(G331));
  XNOR2_X1  g464(.A(new_n822), .B(G171), .ZN(new_n890));
  XNOR2_X1  g465(.A(new_n890), .B(G168), .ZN(new_n891));
  NAND3_X1  g466(.A1(new_n877), .A2(new_n878), .A3(new_n891), .ZN(new_n892));
  INV_X1    g467(.A(new_n872), .ZN(new_n893));
  OR2_X1    g468(.A1(new_n891), .A2(new_n893), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n892), .A2(new_n894), .ZN(new_n895));
  INV_X1    g470(.A(new_n867), .ZN(new_n896));
  OAI21_X1  g471(.A(new_n859), .B1(new_n895), .B2(new_n896), .ZN(new_n897));
  INV_X1    g472(.A(KEYINPUT103), .ZN(new_n898));
  NAND3_X1  g473(.A1(new_n892), .A2(new_n898), .A3(new_n894), .ZN(new_n899));
  AOI21_X1  g474(.A(new_n867), .B1(new_n895), .B2(KEYINPUT103), .ZN(new_n900));
  AOI21_X1  g475(.A(new_n897), .B1(new_n899), .B2(new_n900), .ZN(new_n901));
  INV_X1    g476(.A(KEYINPUT43), .ZN(new_n902));
  OAI21_X1  g477(.A(KEYINPUT104), .B1(new_n901), .B2(new_n902), .ZN(new_n903));
  INV_X1    g478(.A(KEYINPUT104), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n895), .A2(KEYINPUT103), .ZN(new_n905));
  AND3_X1   g480(.A1(new_n905), .A2(new_n896), .A3(new_n899), .ZN(new_n906));
  OAI211_X1 g481(.A(new_n904), .B(KEYINPUT43), .C1(new_n906), .C2(new_n897), .ZN(new_n907));
  INV_X1    g482(.A(new_n897), .ZN(new_n908));
  INV_X1    g483(.A(KEYINPUT105), .ZN(new_n909));
  AND3_X1   g484(.A1(new_n875), .A2(new_n909), .A3(new_n876), .ZN(new_n910));
  OAI21_X1  g485(.A(new_n891), .B1(new_n875), .B2(new_n909), .ZN(new_n911));
  OAI21_X1  g486(.A(new_n894), .B1(new_n910), .B2(new_n911), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n912), .A2(new_n896), .ZN(new_n913));
  NAND3_X1  g488(.A1(new_n908), .A2(new_n902), .A3(new_n913), .ZN(new_n914));
  NAND3_X1  g489(.A1(new_n903), .A2(new_n907), .A3(new_n914), .ZN(new_n915));
  NOR2_X1   g490(.A1(new_n915), .A2(KEYINPUT44), .ZN(new_n916));
  INV_X1    g491(.A(KEYINPUT44), .ZN(new_n917));
  AOI21_X1  g492(.A(new_n902), .B1(new_n908), .B2(new_n913), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n900), .A2(new_n899), .ZN(new_n919));
  NAND3_X1  g494(.A1(new_n919), .A2(new_n902), .A3(new_n908), .ZN(new_n920));
  AOI21_X1  g495(.A(new_n918), .B1(new_n920), .B2(KEYINPUT106), .ZN(new_n921));
  OR2_X1    g496(.A1(new_n920), .A2(KEYINPUT106), .ZN(new_n922));
  AOI21_X1  g497(.A(new_n917), .B1(new_n921), .B2(new_n922), .ZN(new_n923));
  NOR2_X1   g498(.A1(new_n916), .A2(new_n923), .ZN(G397));
  XNOR2_X1  g499(.A(new_n808), .B(G2067), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n925), .A2(new_n748), .ZN(new_n926));
  AND3_X1   g501(.A1(new_n465), .A2(G40), .A3(new_n472), .ZN(new_n927));
  INV_X1    g502(.A(G1384), .ZN(new_n928));
  INV_X1    g503(.A(KEYINPUT4), .ZN(new_n929));
  XNOR2_X1  g504(.A(new_n489), .B(new_n929), .ZN(new_n930));
  INV_X1    g505(.A(new_n493), .ZN(new_n931));
  AOI21_X1  g506(.A(KEYINPUT70), .B1(new_n931), .B2(new_n497), .ZN(new_n932));
  NOR3_X1   g507(.A1(new_n492), .A2(new_n493), .A3(new_n491), .ZN(new_n933));
  OAI21_X1  g508(.A(new_n500), .B1(new_n932), .B2(new_n933), .ZN(new_n934));
  OAI21_X1  g509(.A(new_n928), .B1(new_n930), .B2(new_n934), .ZN(new_n935));
  INV_X1    g510(.A(KEYINPUT45), .ZN(new_n936));
  NAND3_X1  g511(.A1(new_n927), .A2(new_n935), .A3(new_n936), .ZN(new_n937));
  XNOR2_X1  g512(.A(new_n937), .B(KEYINPUT107), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n926), .A2(new_n938), .ZN(new_n939));
  XOR2_X1   g514(.A(new_n939), .B(KEYINPUT123), .Z(new_n940));
  INV_X1    g515(.A(G1996), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n938), .A2(new_n941), .ZN(new_n942));
  XNOR2_X1  g517(.A(new_n942), .B(KEYINPUT46), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n940), .A2(new_n943), .ZN(new_n944));
  XNOR2_X1  g519(.A(new_n944), .B(KEYINPUT47), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n699), .A2(new_n696), .ZN(new_n946));
  XNOR2_X1  g521(.A(new_n946), .B(KEYINPUT108), .ZN(new_n947));
  AND2_X1   g522(.A1(new_n947), .A2(new_n938), .ZN(new_n948));
  OR2_X1    g523(.A1(new_n948), .A2(KEYINPUT48), .ZN(new_n949));
  XNOR2_X1  g524(.A(new_n747), .B(new_n941), .ZN(new_n950));
  AND2_X1   g525(.A1(new_n925), .A2(new_n950), .ZN(new_n951));
  INV_X1    g526(.A(new_n951), .ZN(new_n952));
  XNOR2_X1  g527(.A(new_n691), .B(new_n694), .ZN(new_n953));
  OAI21_X1  g528(.A(new_n938), .B1(new_n952), .B2(new_n953), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n948), .A2(KEYINPUT48), .ZN(new_n955));
  NAND3_X1  g530(.A1(new_n949), .A2(new_n954), .A3(new_n955), .ZN(new_n956));
  NAND3_X1  g531(.A1(new_n951), .A2(new_n694), .A3(new_n691), .ZN(new_n957));
  OAI21_X1  g532(.A(new_n957), .B1(G2067), .B2(new_n809), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n958), .A2(new_n938), .ZN(new_n959));
  AND3_X1   g534(.A1(new_n945), .A2(new_n956), .A3(new_n959), .ZN(new_n960));
  INV_X1    g535(.A(KEYINPUT54), .ZN(new_n961));
  INV_X1    g536(.A(KEYINPUT50), .ZN(new_n962));
  AOI21_X1  g537(.A(new_n962), .B1(new_n503), .B2(new_n928), .ZN(new_n963));
  OAI211_X1 g538(.A(new_n962), .B(new_n928), .C1(new_n930), .C2(new_n934), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n964), .A2(new_n927), .ZN(new_n965));
  OAI21_X1  g540(.A(KEYINPUT116), .B1(new_n963), .B2(new_n965), .ZN(new_n966));
  INV_X1    g541(.A(KEYINPUT116), .ZN(new_n967));
  NAND3_X1  g542(.A1(new_n465), .A2(G40), .A3(new_n472), .ZN(new_n968));
  AOI21_X1  g543(.A(G1384), .B1(new_n490), .B2(new_n840), .ZN(new_n969));
  AOI21_X1  g544(.A(new_n968), .B1(new_n969), .B2(new_n962), .ZN(new_n970));
  INV_X1    g545(.A(KEYINPUT71), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n934), .A2(new_n971), .ZN(new_n972));
  NAND3_X1  g547(.A1(new_n499), .A2(KEYINPUT71), .A3(new_n500), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n972), .A2(new_n973), .ZN(new_n974));
  AOI21_X1  g549(.A(G1384), .B1(new_n974), .B2(new_n490), .ZN(new_n975));
  OAI211_X1 g550(.A(new_n967), .B(new_n970), .C1(new_n975), .C2(new_n962), .ZN(new_n976));
  INV_X1    g551(.A(G1961), .ZN(new_n977));
  NAND3_X1  g552(.A1(new_n966), .A2(new_n976), .A3(new_n977), .ZN(new_n978));
  AOI21_X1  g553(.A(new_n968), .B1(new_n935), .B2(new_n936), .ZN(new_n979));
  INV_X1    g554(.A(KEYINPUT53), .ZN(new_n980));
  AOI21_X1  g555(.A(new_n980), .B1(KEYINPUT120), .B2(new_n795), .ZN(new_n981));
  OAI21_X1  g556(.A(new_n981), .B1(KEYINPUT120), .B2(new_n795), .ZN(new_n982));
  AOI21_X1  g557(.A(new_n982), .B1(new_n969), .B2(KEYINPUT45), .ZN(new_n983));
  NAND2_X1  g558(.A1(new_n979), .A2(new_n983), .ZN(new_n984));
  INV_X1    g559(.A(KEYINPUT110), .ZN(new_n985));
  AOI21_X1  g560(.A(KEYINPUT45), .B1(new_n503), .B2(new_n928), .ZN(new_n986));
  OAI21_X1  g561(.A(new_n927), .B1(new_n935), .B2(new_n936), .ZN(new_n987));
  OAI21_X1  g562(.A(new_n985), .B1(new_n986), .B2(new_n987), .ZN(new_n988));
  AOI21_X1  g563(.A(new_n968), .B1(new_n969), .B2(KEYINPUT45), .ZN(new_n989));
  OAI211_X1 g564(.A(KEYINPUT110), .B(new_n989), .C1(new_n975), .C2(KEYINPUT45), .ZN(new_n990));
  AOI21_X1  g565(.A(G2078), .B1(new_n988), .B2(new_n990), .ZN(new_n991));
  OAI211_X1 g566(.A(new_n978), .B(new_n984), .C1(new_n991), .C2(KEYINPUT53), .ZN(new_n992));
  AOI21_X1  g567(.A(new_n961), .B1(new_n992), .B2(G171), .ZN(new_n993));
  OR2_X1    g568(.A1(new_n991), .A2(KEYINPUT53), .ZN(new_n994));
  INV_X1    g569(.A(KEYINPUT119), .ZN(new_n995));
  NAND3_X1  g570(.A1(new_n503), .A2(KEYINPUT45), .A3(new_n928), .ZN(new_n996));
  NAND4_X1  g571(.A1(new_n996), .A2(new_n979), .A3(KEYINPUT53), .A4(new_n795), .ZN(new_n997));
  AND3_X1   g572(.A1(new_n978), .A2(new_n995), .A3(new_n997), .ZN(new_n998));
  AOI21_X1  g573(.A(new_n995), .B1(new_n978), .B2(new_n997), .ZN(new_n999));
  OAI21_X1  g574(.A(new_n994), .B1(new_n998), .B2(new_n999), .ZN(new_n1000));
  OAI21_X1  g575(.A(new_n993), .B1(new_n1000), .B2(G171), .ZN(new_n1001));
  NOR3_X1   g576(.A1(new_n963), .A2(G2084), .A3(new_n965), .ZN(new_n1002));
  AOI21_X1  g577(.A(G1966), .B1(new_n996), .B2(new_n979), .ZN(new_n1003));
  OAI21_X1  g578(.A(G286), .B1(new_n1002), .B2(new_n1003), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n996), .A2(new_n979), .ZN(new_n1005));
  INV_X1    g580(.A(G1966), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n1005), .A2(new_n1006), .ZN(new_n1007));
  INV_X1    g582(.A(G2084), .ZN(new_n1008));
  OAI211_X1 g583(.A(new_n1008), .B(new_n970), .C1(new_n975), .C2(new_n962), .ZN(new_n1009));
  NAND3_X1  g584(.A1(new_n1007), .A2(G168), .A3(new_n1009), .ZN(new_n1010));
  NAND3_X1  g585(.A1(new_n1004), .A2(new_n1010), .A3(G8), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n1011), .A2(KEYINPUT51), .ZN(new_n1012));
  INV_X1    g587(.A(G8), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n503), .A2(new_n928), .ZN(new_n1014));
  AOI21_X1  g589(.A(new_n965), .B1(KEYINPUT50), .B2(new_n1014), .ZN(new_n1015));
  AOI22_X1  g590(.A1(new_n1015), .A2(new_n1008), .B1(new_n1005), .B2(new_n1006), .ZN(new_n1016));
  AOI21_X1  g591(.A(new_n1013), .B1(new_n1016), .B2(G168), .ZN(new_n1017));
  INV_X1    g592(.A(KEYINPUT51), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n1017), .A2(new_n1018), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n1012), .A2(new_n1019), .ZN(new_n1020));
  OAI211_X1 g595(.A(KEYINPUT55), .B(G8), .C1(new_n509), .C2(new_n515), .ZN(new_n1021));
  INV_X1    g596(.A(KEYINPUT111), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n1021), .A2(new_n1022), .ZN(new_n1023));
  NAND4_X1  g598(.A1(G303), .A2(KEYINPUT111), .A3(KEYINPUT55), .A4(G8), .ZN(new_n1024));
  AND3_X1   g599(.A1(new_n1023), .A2(new_n1024), .A3(KEYINPUT112), .ZN(new_n1025));
  AOI21_X1  g600(.A(KEYINPUT112), .B1(new_n1023), .B2(new_n1024), .ZN(new_n1026));
  AOI21_X1  g601(.A(KEYINPUT55), .B1(G303), .B2(G8), .ZN(new_n1027));
  NOR3_X1   g602(.A1(new_n1025), .A2(new_n1026), .A3(new_n1027), .ZN(new_n1028));
  INV_X1    g603(.A(new_n1028), .ZN(new_n1029));
  NAND3_X1  g604(.A1(new_n988), .A2(new_n990), .A3(new_n724), .ZN(new_n1030));
  NAND2_X1  g605(.A1(new_n975), .A2(new_n962), .ZN(new_n1031));
  INV_X1    g606(.A(G2090), .ZN(new_n1032));
  AOI21_X1  g607(.A(new_n968), .B1(new_n935), .B2(KEYINPUT50), .ZN(new_n1033));
  NAND3_X1  g608(.A1(new_n1031), .A2(new_n1032), .A3(new_n1033), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n1030), .A2(new_n1034), .ZN(new_n1035));
  AOI21_X1  g610(.A(new_n1029), .B1(new_n1035), .B2(G8), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n1015), .A2(new_n1032), .ZN(new_n1037));
  AOI211_X1 g612(.A(new_n1013), .B(new_n1028), .C1(new_n1030), .C2(new_n1037), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n573), .A2(new_n706), .ZN(new_n1039));
  OAI21_X1  g614(.A(G1981), .B1(new_n568), .B2(new_n572), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n1039), .A2(new_n1040), .ZN(new_n1041));
  INV_X1    g616(.A(KEYINPUT49), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n1041), .A2(new_n1042), .ZN(new_n1043));
  NAND2_X1  g618(.A1(new_n927), .A2(new_n969), .ZN(new_n1044));
  NAND3_X1  g619(.A1(new_n1039), .A2(new_n1040), .A3(KEYINPUT49), .ZN(new_n1045));
  NAND4_X1  g620(.A1(new_n1043), .A2(G8), .A3(new_n1044), .A4(new_n1045), .ZN(new_n1046));
  NAND3_X1  g621(.A1(new_n712), .A2(G1976), .A3(new_n714), .ZN(new_n1047));
  NAND3_X1  g622(.A1(new_n1047), .A2(new_n1044), .A3(G8), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n1048), .A2(KEYINPUT52), .ZN(new_n1049));
  INV_X1    g624(.A(G1976), .ZN(new_n1050));
  AOI21_X1  g625(.A(KEYINPUT52), .B1(G288), .B2(new_n1050), .ZN(new_n1051));
  NAND4_X1  g626(.A1(new_n1047), .A2(new_n1044), .A3(G8), .A4(new_n1051), .ZN(new_n1052));
  NAND3_X1  g627(.A1(new_n1046), .A2(new_n1049), .A3(new_n1052), .ZN(new_n1053));
  NOR3_X1   g628(.A1(new_n1036), .A2(new_n1038), .A3(new_n1053), .ZN(new_n1054));
  NAND3_X1  g629(.A1(new_n1001), .A2(new_n1020), .A3(new_n1054), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n1000), .A2(G171), .ZN(new_n1056));
  NOR2_X1   g631(.A1(new_n992), .A2(G171), .ZN(new_n1057));
  INV_X1    g632(.A(new_n1057), .ZN(new_n1058));
  AOI21_X1  g633(.A(KEYINPUT54), .B1(new_n1056), .B2(new_n1058), .ZN(new_n1059));
  OAI21_X1  g634(.A(KEYINPUT121), .B1(new_n1055), .B2(new_n1059), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n978), .A2(new_n997), .ZN(new_n1061));
  NAND2_X1  g636(.A1(new_n1061), .A2(KEYINPUT119), .ZN(new_n1062));
  NAND3_X1  g637(.A1(new_n978), .A2(new_n995), .A3(new_n997), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n1062), .A2(new_n1063), .ZN(new_n1064));
  AOI21_X1  g639(.A(G301), .B1(new_n1064), .B2(new_n994), .ZN(new_n1065));
  OAI21_X1  g640(.A(new_n961), .B1(new_n1065), .B2(new_n1057), .ZN(new_n1066));
  INV_X1    g641(.A(KEYINPUT121), .ZN(new_n1067));
  INV_X1    g642(.A(new_n1036), .ZN(new_n1068));
  AOI21_X1  g643(.A(new_n1013), .B1(new_n1030), .B2(new_n1037), .ZN(new_n1069));
  AOI21_X1  g644(.A(new_n1053), .B1(new_n1069), .B2(new_n1029), .ZN(new_n1070));
  AND3_X1   g645(.A1(new_n1020), .A2(new_n1068), .A3(new_n1070), .ZN(new_n1071));
  NAND4_X1  g646(.A1(new_n1066), .A2(new_n1067), .A3(new_n1001), .A4(new_n1071), .ZN(new_n1072));
  XNOR2_X1  g647(.A(new_n556), .B(KEYINPUT57), .ZN(new_n1073));
  XOR2_X1   g648(.A(KEYINPUT115), .B(G1956), .Z(new_n1074));
  INV_X1    g649(.A(new_n1074), .ZN(new_n1075));
  AOI21_X1  g650(.A(new_n1075), .B1(new_n1031), .B2(new_n1033), .ZN(new_n1076));
  XOR2_X1   g651(.A(KEYINPUT56), .B(G2072), .Z(new_n1077));
  NOR3_X1   g652(.A1(new_n986), .A2(new_n987), .A3(new_n1077), .ZN(new_n1078));
  OAI21_X1  g653(.A(new_n1073), .B1(new_n1076), .B2(new_n1078), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n966), .A2(new_n976), .ZN(new_n1080));
  OAI22_X1  g655(.A1(new_n1080), .A2(G1348), .B1(G2067), .B2(new_n1044), .ZN(new_n1081));
  INV_X1    g656(.A(new_n1081), .ZN(new_n1082));
  OAI21_X1  g657(.A(new_n1079), .B1(new_n1082), .B2(new_n595), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n1031), .A2(new_n1033), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n1084), .A2(new_n1074), .ZN(new_n1085));
  INV_X1    g660(.A(KEYINPUT57), .ZN(new_n1086));
  XNOR2_X1  g661(.A(new_n556), .B(new_n1086), .ZN(new_n1087));
  INV_X1    g662(.A(new_n1078), .ZN(new_n1088));
  NAND3_X1  g663(.A1(new_n1085), .A2(new_n1087), .A3(new_n1088), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n1083), .A2(new_n1089), .ZN(new_n1090));
  INV_X1    g665(.A(KEYINPUT60), .ZN(new_n1091));
  AOI21_X1  g666(.A(new_n595), .B1(new_n1081), .B2(new_n1091), .ZN(new_n1092));
  OAI21_X1  g667(.A(new_n1092), .B1(new_n1091), .B2(new_n1081), .ZN(new_n1093));
  NAND3_X1  g668(.A1(new_n1082), .A2(KEYINPUT60), .A3(new_n595), .ZN(new_n1094));
  NAND3_X1  g669(.A1(new_n1089), .A2(new_n1079), .A3(KEYINPUT61), .ZN(new_n1095));
  AND2_X1   g670(.A1(new_n1095), .A2(KEYINPUT118), .ZN(new_n1096));
  NOR2_X1   g671(.A1(new_n1095), .A2(KEYINPUT118), .ZN(new_n1097));
  OAI211_X1 g672(.A(new_n1093), .B(new_n1094), .C1(new_n1096), .C2(new_n1097), .ZN(new_n1098));
  AOI21_X1  g673(.A(KEYINPUT61), .B1(new_n1089), .B2(new_n1079), .ZN(new_n1099));
  OR2_X1    g674(.A1(new_n1099), .A2(KEYINPUT117), .ZN(new_n1100));
  NAND2_X1  g675(.A1(new_n1099), .A2(KEYINPUT117), .ZN(new_n1101));
  OAI211_X1 g676(.A(new_n941), .B(new_n989), .C1(new_n975), .C2(KEYINPUT45), .ZN(new_n1102));
  XOR2_X1   g677(.A(KEYINPUT58), .B(G1341), .Z(new_n1103));
  NAND2_X1  g678(.A1(new_n1044), .A2(new_n1103), .ZN(new_n1104));
  AOI21_X1  g679(.A(new_n821), .B1(new_n1102), .B2(new_n1104), .ZN(new_n1105));
  XOR2_X1   g680(.A(new_n1105), .B(KEYINPUT59), .Z(new_n1106));
  NAND3_X1  g681(.A1(new_n1100), .A2(new_n1101), .A3(new_n1106), .ZN(new_n1107));
  OAI21_X1  g682(.A(new_n1090), .B1(new_n1098), .B2(new_n1107), .ZN(new_n1108));
  NAND3_X1  g683(.A1(new_n1060), .A2(new_n1072), .A3(new_n1108), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n1044), .A2(G8), .ZN(new_n1110));
  INV_X1    g685(.A(G288), .ZN(new_n1111));
  NAND3_X1  g686(.A1(new_n1046), .A2(new_n1050), .A3(new_n1111), .ZN(new_n1112));
  AOI21_X1  g687(.A(new_n1110), .B1(new_n1112), .B2(new_n1039), .ZN(new_n1113));
  INV_X1    g688(.A(KEYINPUT113), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n1053), .A2(new_n1114), .ZN(new_n1115));
  NAND4_X1  g690(.A1(new_n1046), .A2(new_n1049), .A3(KEYINPUT113), .A4(new_n1052), .ZN(new_n1116));
  NAND2_X1  g691(.A1(new_n1115), .A2(new_n1116), .ZN(new_n1117));
  AOI21_X1  g692(.A(new_n1113), .B1(new_n1117), .B2(new_n1038), .ZN(new_n1118));
  AOI21_X1  g693(.A(new_n1018), .B1(new_n1017), .B2(new_n1004), .ZN(new_n1119));
  AND3_X1   g694(.A1(new_n1010), .A2(new_n1018), .A3(G8), .ZN(new_n1120));
  OAI21_X1  g695(.A(KEYINPUT62), .B1(new_n1119), .B2(new_n1120), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n1121), .A2(new_n1054), .ZN(new_n1122));
  INV_X1    g697(.A(KEYINPUT62), .ZN(new_n1123));
  NAND3_X1  g698(.A1(new_n1012), .A2(new_n1019), .A3(new_n1123), .ZN(new_n1124));
  NAND3_X1  g699(.A1(new_n1124), .A2(G171), .A3(new_n1000), .ZN(new_n1125));
  OAI21_X1  g700(.A(new_n1118), .B1(new_n1122), .B2(new_n1125), .ZN(new_n1126));
  NOR3_X1   g701(.A1(new_n1016), .A2(new_n1013), .A3(G286), .ZN(new_n1127));
  NAND3_X1  g702(.A1(new_n1068), .A2(new_n1070), .A3(new_n1127), .ZN(new_n1128));
  INV_X1    g703(.A(KEYINPUT63), .ZN(new_n1129));
  NAND2_X1  g704(.A1(new_n1128), .A2(new_n1129), .ZN(new_n1130));
  OR2_X1    g705(.A1(new_n1130), .A2(KEYINPUT114), .ZN(new_n1131));
  NAND3_X1  g706(.A1(new_n1117), .A2(KEYINPUT63), .A3(new_n1127), .ZN(new_n1132));
  NOR2_X1   g707(.A1(new_n1069), .A2(new_n1029), .ZN(new_n1133));
  NOR3_X1   g708(.A1(new_n1132), .A2(new_n1133), .A3(new_n1038), .ZN(new_n1134));
  AOI21_X1  g709(.A(new_n1134), .B1(new_n1130), .B2(KEYINPUT114), .ZN(new_n1135));
  AOI21_X1  g710(.A(new_n1126), .B1(new_n1131), .B2(new_n1135), .ZN(new_n1136));
  NAND2_X1  g711(.A1(new_n1109), .A2(new_n1136), .ZN(new_n1137));
  NOR2_X1   g712(.A1(new_n699), .A2(new_n696), .ZN(new_n1138));
  OAI21_X1  g713(.A(new_n938), .B1(new_n947), .B2(new_n1138), .ZN(new_n1139));
  NAND2_X1  g714(.A1(new_n954), .A2(new_n1139), .ZN(new_n1140));
  XNOR2_X1  g715(.A(new_n1140), .B(KEYINPUT109), .ZN(new_n1141));
  INV_X1    g716(.A(new_n1141), .ZN(new_n1142));
  AOI21_X1  g717(.A(KEYINPUT122), .B1(new_n1137), .B2(new_n1142), .ZN(new_n1143));
  INV_X1    g718(.A(KEYINPUT122), .ZN(new_n1144));
  AOI211_X1 g719(.A(new_n1144), .B(new_n1141), .C1(new_n1109), .C2(new_n1136), .ZN(new_n1145));
  OAI21_X1  g720(.A(new_n960), .B1(new_n1143), .B2(new_n1145), .ZN(new_n1146));
  INV_X1    g721(.A(KEYINPUT124), .ZN(new_n1147));
  NAND2_X1  g722(.A1(new_n1146), .A2(new_n1147), .ZN(new_n1148));
  OAI211_X1 g723(.A(KEYINPUT124), .B(new_n960), .C1(new_n1143), .C2(new_n1145), .ZN(new_n1149));
  NAND2_X1  g724(.A1(new_n1148), .A2(new_n1149), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g725(.A(KEYINPUT127), .ZN(new_n1152));
  INV_X1    g726(.A(G227), .ZN(new_n1153));
  NAND2_X1  g727(.A1(new_n1153), .A2(G319), .ZN(new_n1154));
  XNOR2_X1  g728(.A(new_n1154), .B(KEYINPUT125), .ZN(new_n1155));
  AOI21_X1  g729(.A(new_n1155), .B1(new_n645), .B2(new_n652), .ZN(new_n1156));
  INV_X1    g730(.A(KEYINPUT126), .ZN(new_n1157));
  NAND2_X1  g731(.A1(new_n1156), .A2(new_n1157), .ZN(new_n1158));
  INV_X1    g732(.A(G229), .ZN(new_n1159));
  NAND2_X1  g733(.A1(new_n1158), .A2(new_n1159), .ZN(new_n1160));
  NOR2_X1   g734(.A1(new_n1156), .A2(new_n1157), .ZN(new_n1161));
  OAI21_X1  g735(.A(new_n1152), .B1(new_n1160), .B2(new_n1161), .ZN(new_n1162));
  INV_X1    g736(.A(new_n1161), .ZN(new_n1163));
  NAND4_X1  g737(.A1(new_n1163), .A2(KEYINPUT127), .A3(new_n1159), .A4(new_n1158), .ZN(new_n1164));
  NAND2_X1  g738(.A1(new_n1162), .A2(new_n1164), .ZN(new_n1165));
  AND3_X1   g739(.A1(new_n1165), .A2(new_n861), .A3(new_n915), .ZN(G308));
  NAND3_X1  g740(.A1(new_n1165), .A2(new_n861), .A3(new_n915), .ZN(G225));
endmodule


