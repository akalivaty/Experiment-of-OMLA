//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 0 0 0 0 1 0 0 1 0 0 1 1 0 1 1 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 0 0 1 0 1 1 1 0 0 0 0 1 0 1 1 1 1 0 1 1 0 0 0 0 0 0 0 1 1 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:22:42 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n636, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n649, new_n650, new_n651, new_n652,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n682,
    new_n683, new_n684, new_n685, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n701, new_n703, new_n704, new_n705, new_n707,
    new_n708, new_n709, new_n710, new_n711, new_n712, new_n713, new_n714,
    new_n715, new_n716, new_n717, new_n718, new_n719, new_n720, new_n721,
    new_n722, new_n723, new_n725, new_n726, new_n727, new_n728, new_n729,
    new_n730, new_n731, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n756, new_n757, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n779, new_n780, new_n781, new_n782,
    new_n783, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n908, new_n909, new_n910, new_n911, new_n912, new_n913,
    new_n914, new_n915, new_n916, new_n917, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n968, new_n969, new_n970, new_n971, new_n972, new_n973,
    new_n974, new_n975, new_n976, new_n977, new_n978, new_n979, new_n980,
    new_n981, new_n982, new_n983, new_n984;
  OAI21_X1  g000(.A(G214), .B1(G237), .B2(G902), .ZN(new_n187));
  INV_X1    g001(.A(KEYINPUT69), .ZN(new_n188));
  INV_X1    g002(.A(KEYINPUT2), .ZN(new_n189));
  INV_X1    g003(.A(G113), .ZN(new_n190));
  OAI21_X1  g004(.A(new_n188), .B1(new_n189), .B2(new_n190), .ZN(new_n191));
  NAND3_X1  g005(.A1(KEYINPUT69), .A2(KEYINPUT2), .A3(G113), .ZN(new_n192));
  AOI22_X1  g006(.A1(new_n191), .A2(new_n192), .B1(new_n189), .B2(new_n190), .ZN(new_n193));
  XNOR2_X1  g007(.A(G116), .B(G119), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n194), .A2(KEYINPUT5), .ZN(new_n195));
  INV_X1    g009(.A(G116), .ZN(new_n196));
  NOR3_X1   g010(.A1(new_n196), .A2(KEYINPUT5), .A3(G119), .ZN(new_n197));
  NOR2_X1   g011(.A1(new_n197), .A2(new_n190), .ZN(new_n198));
  AOI22_X1  g012(.A1(new_n193), .A2(new_n194), .B1(new_n195), .B2(new_n198), .ZN(new_n199));
  INV_X1    g013(.A(G101), .ZN(new_n200));
  INV_X1    g014(.A(KEYINPUT79), .ZN(new_n201));
  INV_X1    g015(.A(G104), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NAND2_X1  g017(.A1(KEYINPUT79), .A2(G104), .ZN(new_n204));
  NAND3_X1  g018(.A1(new_n203), .A2(G107), .A3(new_n204), .ZN(new_n205));
  INV_X1    g019(.A(KEYINPUT3), .ZN(new_n206));
  INV_X1    g020(.A(G107), .ZN(new_n207));
  NAND3_X1  g021(.A1(new_n206), .A2(new_n207), .A3(G104), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n205), .A2(new_n208), .ZN(new_n209));
  INV_X1    g023(.A(new_n209), .ZN(new_n210));
  AND2_X1   g024(.A1(KEYINPUT79), .A2(G104), .ZN(new_n211));
  NOR2_X1   g025(.A1(KEYINPUT79), .A2(G104), .ZN(new_n212));
  OAI21_X1  g026(.A(new_n207), .B1(new_n211), .B2(new_n212), .ZN(new_n213));
  INV_X1    g027(.A(KEYINPUT80), .ZN(new_n214));
  AND3_X1   g028(.A1(new_n213), .A2(new_n214), .A3(KEYINPUT3), .ZN(new_n215));
  AOI21_X1  g029(.A(new_n214), .B1(new_n213), .B2(KEYINPUT3), .ZN(new_n216));
  OAI211_X1 g030(.A(new_n200), .B(new_n210), .C1(new_n215), .C2(new_n216), .ZN(new_n217));
  INV_X1    g031(.A(KEYINPUT82), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n202), .A2(G107), .ZN(new_n219));
  AOI21_X1  g033(.A(new_n200), .B1(new_n213), .B2(new_n219), .ZN(new_n220));
  INV_X1    g034(.A(new_n220), .ZN(new_n221));
  AND3_X1   g035(.A1(new_n217), .A2(new_n218), .A3(new_n221), .ZN(new_n222));
  AOI21_X1  g036(.A(new_n218), .B1(new_n217), .B2(new_n221), .ZN(new_n223));
  OAI21_X1  g037(.A(new_n199), .B1(new_n222), .B2(new_n223), .ZN(new_n224));
  XOR2_X1   g038(.A(new_n193), .B(new_n194), .Z(new_n225));
  INV_X1    g039(.A(new_n225), .ZN(new_n226));
  OAI21_X1  g040(.A(new_n210), .B1(new_n215), .B2(new_n216), .ZN(new_n227));
  INV_X1    g041(.A(KEYINPUT4), .ZN(new_n228));
  NAND3_X1  g042(.A1(new_n227), .A2(new_n228), .A3(G101), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n217), .A2(KEYINPUT4), .ZN(new_n230));
  AOI21_X1  g044(.A(G107), .B1(new_n203), .B2(new_n204), .ZN(new_n231));
  OAI21_X1  g045(.A(KEYINPUT80), .B1(new_n231), .B2(new_n206), .ZN(new_n232));
  NAND3_X1  g046(.A1(new_n213), .A2(new_n214), .A3(KEYINPUT3), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n232), .A2(new_n233), .ZN(new_n234));
  AOI21_X1  g048(.A(new_n200), .B1(new_n234), .B2(new_n210), .ZN(new_n235));
  OAI211_X1 g049(.A(new_n226), .B(new_n229), .C1(new_n230), .C2(new_n235), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n224), .A2(new_n236), .ZN(new_n237));
  INV_X1    g051(.A(KEYINPUT6), .ZN(new_n238));
  XNOR2_X1  g052(.A(G110), .B(G122), .ZN(new_n239));
  INV_X1    g053(.A(new_n239), .ZN(new_n240));
  AND4_X1   g054(.A1(KEYINPUT86), .A2(new_n237), .A3(new_n238), .A4(new_n240), .ZN(new_n241));
  AOI21_X1  g055(.A(new_n239), .B1(new_n224), .B2(new_n236), .ZN(new_n242));
  AOI21_X1  g056(.A(KEYINPUT86), .B1(new_n242), .B2(new_n238), .ZN(new_n243));
  NOR2_X1   g057(.A1(new_n241), .A2(new_n243), .ZN(new_n244));
  NAND3_X1  g058(.A1(new_n224), .A2(new_n239), .A3(new_n236), .ZN(new_n245));
  INV_X1    g059(.A(KEYINPUT85), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n245), .A2(new_n246), .ZN(new_n247));
  NAND4_X1  g061(.A1(new_n224), .A2(KEYINPUT85), .A3(new_n236), .A4(new_n239), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n247), .A2(new_n248), .ZN(new_n249));
  NOR2_X1   g063(.A1(new_n242), .A2(new_n238), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  INV_X1    g065(.A(KEYINPUT0), .ZN(new_n252));
  INV_X1    g066(.A(G128), .ZN(new_n253));
  NOR2_X1   g067(.A1(new_n252), .A2(new_n253), .ZN(new_n254));
  INV_X1    g068(.A(G143), .ZN(new_n255));
  NOR2_X1   g069(.A1(new_n255), .A2(G146), .ZN(new_n256));
  INV_X1    g070(.A(new_n256), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n255), .A2(KEYINPUT65), .ZN(new_n258));
  INV_X1    g072(.A(KEYINPUT65), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n259), .A2(G143), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n258), .A2(new_n260), .ZN(new_n261));
  INV_X1    g075(.A(G146), .ZN(new_n262));
  OAI211_X1 g076(.A(new_n254), .B(new_n257), .C1(new_n261), .C2(new_n262), .ZN(new_n263));
  NOR2_X1   g077(.A1(new_n262), .A2(G143), .ZN(new_n264));
  AOI21_X1  g078(.A(new_n264), .B1(new_n261), .B2(new_n262), .ZN(new_n265));
  OAI21_X1  g079(.A(KEYINPUT64), .B1(new_n252), .B2(new_n253), .ZN(new_n266));
  INV_X1    g080(.A(KEYINPUT64), .ZN(new_n267));
  NAND3_X1  g081(.A1(new_n267), .A2(KEYINPUT0), .A3(G128), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n252), .A2(new_n253), .ZN(new_n269));
  NAND3_X1  g083(.A1(new_n266), .A2(new_n268), .A3(new_n269), .ZN(new_n270));
  OAI21_X1  g084(.A(new_n263), .B1(new_n265), .B2(new_n270), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n271), .A2(G125), .ZN(new_n272));
  NOR2_X1   g086(.A1(new_n253), .A2(KEYINPUT1), .ZN(new_n273));
  OAI211_X1 g087(.A(new_n257), .B(new_n273), .C1(new_n261), .C2(new_n262), .ZN(new_n274));
  INV_X1    g088(.A(KEYINPUT1), .ZN(new_n275));
  OAI21_X1  g089(.A(G128), .B1(new_n256), .B2(new_n275), .ZN(new_n276));
  INV_X1    g090(.A(new_n276), .ZN(new_n277));
  OAI21_X1  g091(.A(new_n274), .B1(new_n265), .B2(new_n277), .ZN(new_n278));
  OAI21_X1  g092(.A(new_n272), .B1(G125), .B2(new_n278), .ZN(new_n279));
  INV_X1    g093(.A(G953), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n280), .A2(G224), .ZN(new_n281));
  XNOR2_X1  g095(.A(new_n279), .B(new_n281), .ZN(new_n282));
  INV_X1    g096(.A(new_n282), .ZN(new_n283));
  NAND3_X1  g097(.A1(new_n244), .A2(new_n251), .A3(new_n283), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n281), .A2(KEYINPUT7), .ZN(new_n285));
  XNOR2_X1  g099(.A(new_n279), .B(new_n285), .ZN(new_n286));
  AOI21_X1  g100(.A(new_n209), .B1(new_n232), .B2(new_n233), .ZN(new_n287));
  AOI21_X1  g101(.A(new_n220), .B1(new_n287), .B2(new_n200), .ZN(new_n288));
  XNOR2_X1  g102(.A(new_n288), .B(new_n199), .ZN(new_n289));
  XNOR2_X1  g103(.A(new_n239), .B(KEYINPUT8), .ZN(new_n290));
  AOI21_X1  g104(.A(new_n286), .B1(new_n289), .B2(new_n290), .ZN(new_n291));
  AOI21_X1  g105(.A(G902), .B1(new_n249), .B2(new_n291), .ZN(new_n292));
  OAI21_X1  g106(.A(G210), .B1(G237), .B2(G902), .ZN(new_n293));
  AND3_X1   g107(.A1(new_n284), .A2(new_n292), .A3(new_n293), .ZN(new_n294));
  AOI21_X1  g108(.A(new_n293), .B1(new_n284), .B2(new_n292), .ZN(new_n295));
  OAI21_X1  g109(.A(new_n187), .B1(new_n294), .B2(new_n295), .ZN(new_n296));
  XNOR2_X1  g110(.A(KEYINPUT9), .B(G234), .ZN(new_n297));
  XNOR2_X1  g111(.A(new_n297), .B(KEYINPUT77), .ZN(new_n298));
  OAI21_X1  g112(.A(G221), .B1(new_n298), .B2(G902), .ZN(new_n299));
  XNOR2_X1  g113(.A(new_n299), .B(KEYINPUT78), .ZN(new_n300));
  INV_X1    g114(.A(new_n300), .ZN(new_n301));
  XNOR2_X1  g115(.A(KEYINPUT71), .B(G953), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n302), .A2(G227), .ZN(new_n303));
  XOR2_X1   g117(.A(G110), .B(G140), .Z(new_n304));
  XNOR2_X1  g118(.A(new_n303), .B(new_n304), .ZN(new_n305));
  AOI21_X1  g119(.A(new_n271), .B1(new_n235), .B2(new_n228), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n227), .A2(G101), .ZN(new_n307));
  NAND3_X1  g121(.A1(new_n307), .A2(KEYINPUT4), .A3(new_n217), .ZN(new_n308));
  AND3_X1   g122(.A1(new_n306), .A2(new_n308), .A3(KEYINPUT81), .ZN(new_n309));
  AOI21_X1  g123(.A(KEYINPUT81), .B1(new_n306), .B2(new_n308), .ZN(new_n310));
  NOR2_X1   g124(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  NOR2_X1   g125(.A1(new_n259), .A2(G143), .ZN(new_n312));
  NOR2_X1   g126(.A1(new_n255), .A2(KEYINPUT65), .ZN(new_n313));
  OAI21_X1  g127(.A(new_n262), .B1(new_n312), .B2(new_n313), .ZN(new_n314));
  AOI21_X1  g128(.A(new_n253), .B1(new_n314), .B2(KEYINPUT1), .ZN(new_n315));
  XNOR2_X1  g129(.A(KEYINPUT65), .B(G143), .ZN(new_n316));
  AOI21_X1  g130(.A(new_n256), .B1(new_n316), .B2(G146), .ZN(new_n317));
  OAI21_X1  g131(.A(new_n274), .B1(new_n315), .B2(new_n317), .ZN(new_n318));
  NAND3_X1  g132(.A1(new_n217), .A2(new_n318), .A3(new_n221), .ZN(new_n319));
  NOR2_X1   g133(.A1(new_n319), .A2(KEYINPUT10), .ZN(new_n320));
  OAI21_X1  g134(.A(new_n278), .B1(new_n222), .B2(new_n223), .ZN(new_n321));
  AOI21_X1  g135(.A(new_n320), .B1(new_n321), .B2(KEYINPUT10), .ZN(new_n322));
  INV_X1    g136(.A(G137), .ZN(new_n323));
  NAND3_X1  g137(.A1(new_n323), .A2(KEYINPUT11), .A3(G134), .ZN(new_n324));
  INV_X1    g138(.A(G134), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n325), .A2(G137), .ZN(new_n326));
  AND2_X1   g140(.A1(new_n324), .A2(new_n326), .ZN(new_n327));
  INV_X1    g141(.A(G131), .ZN(new_n328));
  INV_X1    g142(.A(KEYINPUT11), .ZN(new_n329));
  OAI21_X1  g143(.A(new_n329), .B1(new_n325), .B2(G137), .ZN(new_n330));
  NAND4_X1  g144(.A1(new_n327), .A2(KEYINPUT66), .A3(new_n328), .A4(new_n330), .ZN(new_n331));
  NAND4_X1  g145(.A1(new_n330), .A2(new_n324), .A3(new_n328), .A4(new_n326), .ZN(new_n332));
  INV_X1    g146(.A(KEYINPUT66), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n331), .A2(new_n334), .ZN(new_n335));
  NAND3_X1  g149(.A1(new_n330), .A2(new_n324), .A3(new_n326), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n336), .A2(KEYINPUT67), .ZN(new_n337));
  INV_X1    g151(.A(KEYINPUT67), .ZN(new_n338));
  NAND4_X1  g152(.A1(new_n330), .A2(new_n324), .A3(new_n338), .A4(new_n326), .ZN(new_n339));
  NAND3_X1  g153(.A1(new_n337), .A2(G131), .A3(new_n339), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n335), .A2(new_n340), .ZN(new_n341));
  NOR3_X1   g155(.A1(new_n311), .A2(new_n322), .A3(new_n341), .ZN(new_n342));
  AND2_X1   g156(.A1(new_n339), .A2(G131), .ZN(new_n343));
  AOI22_X1  g157(.A1(new_n337), .A2(new_n343), .B1(new_n331), .B2(new_n334), .ZN(new_n344));
  INV_X1    g158(.A(new_n320), .ZN(new_n345));
  INV_X1    g159(.A(new_n278), .ZN(new_n346));
  AOI211_X1 g160(.A(G101), .B(new_n209), .C1(new_n232), .C2(new_n233), .ZN(new_n347));
  OAI21_X1  g161(.A(KEYINPUT82), .B1(new_n347), .B2(new_n220), .ZN(new_n348));
  NAND3_X1  g162(.A1(new_n217), .A2(new_n218), .A3(new_n221), .ZN(new_n349));
  AOI21_X1  g163(.A(new_n346), .B1(new_n348), .B2(new_n349), .ZN(new_n350));
  INV_X1    g164(.A(KEYINPUT10), .ZN(new_n351));
  OAI21_X1  g165(.A(new_n345), .B1(new_n350), .B2(new_n351), .ZN(new_n352));
  INV_X1    g166(.A(KEYINPUT81), .ZN(new_n353));
  NOR2_X1   g167(.A1(new_n230), .A2(new_n235), .ZN(new_n354));
  INV_X1    g168(.A(new_n271), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n229), .A2(new_n355), .ZN(new_n356));
  OAI21_X1  g170(.A(new_n353), .B1(new_n354), .B2(new_n356), .ZN(new_n357));
  NAND3_X1  g171(.A1(new_n306), .A2(new_n308), .A3(KEYINPUT81), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n357), .A2(new_n358), .ZN(new_n359));
  AOI21_X1  g173(.A(new_n344), .B1(new_n352), .B2(new_n359), .ZN(new_n360));
  OAI21_X1  g174(.A(new_n305), .B1(new_n342), .B2(new_n360), .ZN(new_n361));
  NAND3_X1  g175(.A1(new_n352), .A2(new_n344), .A3(new_n359), .ZN(new_n362));
  INV_X1    g176(.A(KEYINPUT83), .ZN(new_n363));
  NOR3_X1   g177(.A1(new_n363), .A2(KEYINPUT84), .A3(KEYINPUT12), .ZN(new_n364));
  AND3_X1   g178(.A1(new_n217), .A2(new_n318), .A3(new_n221), .ZN(new_n365));
  AOI21_X1  g179(.A(new_n278), .B1(new_n217), .B2(new_n221), .ZN(new_n366));
  OAI21_X1  g180(.A(new_n364), .B1(new_n365), .B2(new_n366), .ZN(new_n367));
  OAI211_X1 g181(.A(new_n319), .B(KEYINPUT84), .C1(new_n288), .C2(new_n278), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  OAI211_X1 g183(.A(KEYINPUT83), .B(new_n341), .C1(new_n365), .C2(new_n366), .ZN(new_n370));
  AOI22_X1  g184(.A1(new_n369), .A2(new_n341), .B1(KEYINPUT12), .B2(new_n370), .ZN(new_n371));
  INV_X1    g185(.A(new_n305), .ZN(new_n372));
  NAND3_X1  g186(.A1(new_n362), .A2(new_n371), .A3(new_n372), .ZN(new_n373));
  AOI211_X1 g187(.A(G469), .B(G902), .C1(new_n361), .C2(new_n373), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n362), .A2(new_n371), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n375), .A2(new_n305), .ZN(new_n376));
  OAI21_X1  g190(.A(new_n341), .B1(new_n311), .B2(new_n322), .ZN(new_n377));
  NAND3_X1  g191(.A1(new_n377), .A2(new_n362), .A3(new_n372), .ZN(new_n378));
  NAND3_X1  g192(.A1(new_n376), .A2(G469), .A3(new_n378), .ZN(new_n379));
  NAND2_X1  g193(.A1(G469), .A2(G902), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n379), .A2(new_n380), .ZN(new_n381));
  OAI21_X1  g195(.A(new_n301), .B1(new_n374), .B2(new_n381), .ZN(new_n382));
  XNOR2_X1  g196(.A(G125), .B(G140), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n383), .A2(KEYINPUT16), .ZN(new_n384));
  INV_X1    g198(.A(G140), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n385), .A2(G125), .ZN(new_n386));
  OAI21_X1  g200(.A(new_n384), .B1(KEYINPUT16), .B2(new_n386), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n387), .A2(new_n262), .ZN(new_n388));
  OAI211_X1 g202(.A(new_n384), .B(G146), .C1(KEYINPUT16), .C2(new_n386), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n388), .A2(new_n389), .ZN(new_n390));
  INV_X1    g204(.A(new_n390), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n280), .A2(KEYINPUT71), .ZN(new_n392));
  INV_X1    g206(.A(KEYINPUT71), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n393), .A2(G953), .ZN(new_n394));
  INV_X1    g208(.A(G237), .ZN(new_n395));
  NAND4_X1  g209(.A1(new_n392), .A2(new_n394), .A3(G214), .A4(new_n395), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n396), .A2(new_n316), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n397), .A2(KEYINPUT87), .ZN(new_n398));
  NAND4_X1  g212(.A1(new_n302), .A2(G143), .A3(G214), .A4(new_n395), .ZN(new_n399));
  INV_X1    g213(.A(KEYINPUT87), .ZN(new_n400));
  NAND3_X1  g214(.A1(new_n396), .A2(new_n400), .A3(new_n316), .ZN(new_n401));
  NAND3_X1  g215(.A1(new_n398), .A2(new_n399), .A3(new_n401), .ZN(new_n402));
  NAND3_X1  g216(.A1(new_n402), .A2(KEYINPUT17), .A3(G131), .ZN(new_n403));
  NAND4_X1  g217(.A1(new_n398), .A2(new_n328), .A3(new_n399), .A4(new_n401), .ZN(new_n404));
  INV_X1    g218(.A(KEYINPUT90), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n404), .A2(new_n405), .ZN(new_n406));
  AND2_X1   g220(.A1(new_n401), .A2(new_n399), .ZN(new_n407));
  NAND4_X1  g221(.A1(new_n407), .A2(KEYINPUT90), .A3(new_n328), .A4(new_n398), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n402), .A2(G131), .ZN(new_n409));
  NAND3_X1  g223(.A1(new_n406), .A2(new_n408), .A3(new_n409), .ZN(new_n410));
  OAI211_X1 g224(.A(new_n391), .B(new_n403), .C1(new_n410), .C2(KEYINPUT17), .ZN(new_n411));
  XOR2_X1   g225(.A(G113), .B(G122), .Z(new_n412));
  XNOR2_X1  g226(.A(KEYINPUT91), .B(G104), .ZN(new_n413));
  XNOR2_X1  g227(.A(new_n412), .B(new_n413), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n401), .A2(new_n399), .ZN(new_n415));
  AOI21_X1  g229(.A(new_n400), .B1(new_n396), .B2(new_n316), .ZN(new_n416));
  OAI211_X1 g230(.A(KEYINPUT18), .B(G131), .C1(new_n415), .C2(new_n416), .ZN(new_n417));
  XNOR2_X1  g231(.A(new_n383), .B(new_n262), .ZN(new_n418));
  AND2_X1   g232(.A1(new_n417), .A2(new_n418), .ZN(new_n419));
  NAND2_X1  g233(.A1(KEYINPUT18), .A2(G131), .ZN(new_n420));
  NAND4_X1  g234(.A1(new_n398), .A2(new_n399), .A3(new_n401), .A4(new_n420), .ZN(new_n421));
  INV_X1    g235(.A(KEYINPUT88), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n421), .A2(new_n422), .ZN(new_n423));
  NAND4_X1  g237(.A1(new_n407), .A2(KEYINPUT88), .A3(new_n398), .A4(new_n420), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n423), .A2(new_n424), .ZN(new_n425));
  INV_X1    g239(.A(KEYINPUT89), .ZN(new_n426));
  AND3_X1   g240(.A1(new_n419), .A2(new_n425), .A3(new_n426), .ZN(new_n427));
  AOI21_X1  g241(.A(new_n426), .B1(new_n419), .B2(new_n425), .ZN(new_n428));
  OAI211_X1 g242(.A(new_n411), .B(new_n414), .C1(new_n427), .C2(new_n428), .ZN(new_n429));
  XNOR2_X1  g243(.A(new_n383), .B(KEYINPUT19), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n430), .A2(new_n262), .ZN(new_n431));
  AND2_X1   g245(.A1(new_n431), .A2(new_n389), .ZN(new_n432));
  AND2_X1   g246(.A1(new_n410), .A2(new_n432), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n419), .A2(new_n425), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n434), .A2(KEYINPUT89), .ZN(new_n435));
  NAND3_X1  g249(.A1(new_n419), .A2(new_n425), .A3(new_n426), .ZN(new_n436));
  AOI21_X1  g250(.A(new_n433), .B1(new_n435), .B2(new_n436), .ZN(new_n437));
  OAI21_X1  g251(.A(new_n429), .B1(new_n437), .B2(new_n414), .ZN(new_n438));
  NOR2_X1   g252(.A1(G475), .A2(G902), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n438), .A2(new_n439), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n440), .A2(KEYINPUT92), .ZN(new_n441));
  INV_X1    g255(.A(KEYINPUT92), .ZN(new_n442));
  NAND3_X1  g256(.A1(new_n438), .A2(new_n442), .A3(new_n439), .ZN(new_n443));
  NAND3_X1  g257(.A1(new_n441), .A2(KEYINPUT20), .A3(new_n443), .ZN(new_n444));
  AOI21_X1  g258(.A(new_n442), .B1(new_n438), .B2(new_n439), .ZN(new_n445));
  INV_X1    g259(.A(KEYINPUT20), .ZN(new_n446));
  INV_X1    g260(.A(G902), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n435), .A2(new_n436), .ZN(new_n448));
  AOI21_X1  g262(.A(new_n414), .B1(new_n448), .B2(new_n411), .ZN(new_n449));
  INV_X1    g263(.A(new_n429), .ZN(new_n450));
  OAI21_X1  g264(.A(new_n447), .B1(new_n449), .B2(new_n450), .ZN(new_n451));
  XOR2_X1   g265(.A(KEYINPUT93), .B(G475), .Z(new_n452));
  AOI22_X1  g266(.A1(new_n445), .A2(new_n446), .B1(new_n451), .B2(new_n452), .ZN(new_n453));
  NOR2_X1   g267(.A1(new_n255), .A2(G128), .ZN(new_n454));
  AOI21_X1  g268(.A(new_n454), .B1(new_n316), .B2(G128), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n455), .A2(new_n325), .ZN(new_n456));
  XNOR2_X1  g270(.A(G116), .B(G122), .ZN(new_n457));
  XNOR2_X1  g271(.A(new_n457), .B(new_n207), .ZN(new_n458));
  AND2_X1   g272(.A1(new_n455), .A2(KEYINPUT13), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n316), .A2(G128), .ZN(new_n460));
  OAI21_X1  g274(.A(G134), .B1(new_n460), .B2(KEYINPUT13), .ZN(new_n461));
  OAI211_X1 g275(.A(new_n456), .B(new_n458), .C1(new_n459), .C2(new_n461), .ZN(new_n462));
  XNOR2_X1  g276(.A(new_n455), .B(new_n325), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n457), .A2(new_n207), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  INV_X1    g279(.A(KEYINPUT14), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n457), .A2(new_n466), .ZN(new_n467));
  NAND3_X1  g281(.A1(new_n196), .A2(KEYINPUT14), .A3(G122), .ZN(new_n468));
  NAND3_X1  g282(.A1(new_n467), .A2(G107), .A3(new_n468), .ZN(new_n469));
  XNOR2_X1  g283(.A(new_n469), .B(KEYINPUT94), .ZN(new_n470));
  OAI21_X1  g284(.A(new_n462), .B1(new_n465), .B2(new_n470), .ZN(new_n471));
  INV_X1    g285(.A(G217), .ZN(new_n472));
  NOR3_X1   g286(.A1(new_n298), .A2(new_n472), .A3(G953), .ZN(new_n473));
  XNOR2_X1  g287(.A(new_n471), .B(new_n473), .ZN(new_n474));
  NOR2_X1   g288(.A1(new_n474), .A2(G902), .ZN(new_n475));
  INV_X1    g289(.A(G478), .ZN(new_n476));
  NOR2_X1   g290(.A1(new_n476), .A2(KEYINPUT15), .ZN(new_n477));
  XNOR2_X1  g291(.A(new_n475), .B(new_n477), .ZN(new_n478));
  INV_X1    g292(.A(new_n302), .ZN(new_n479));
  NAND2_X1  g293(.A1(G234), .A2(G237), .ZN(new_n480));
  NAND3_X1  g294(.A1(new_n479), .A2(G902), .A3(new_n480), .ZN(new_n481));
  INV_X1    g295(.A(new_n481), .ZN(new_n482));
  XNOR2_X1  g296(.A(KEYINPUT21), .B(G898), .ZN(new_n483));
  AND2_X1   g297(.A1(new_n280), .A2(G952), .ZN(new_n484));
  AOI22_X1  g298(.A1(new_n482), .A2(new_n483), .B1(new_n480), .B2(new_n484), .ZN(new_n485));
  INV_X1    g299(.A(new_n485), .ZN(new_n486));
  NAND4_X1  g300(.A1(new_n444), .A2(new_n453), .A3(new_n478), .A4(new_n486), .ZN(new_n487));
  NOR3_X1   g301(.A1(new_n296), .A2(new_n382), .A3(new_n487), .ZN(new_n488));
  AOI21_X1  g302(.A(new_n472), .B1(G234), .B2(new_n447), .ZN(new_n489));
  INV_X1    g303(.A(new_n489), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n383), .A2(new_n262), .ZN(new_n491));
  AND2_X1   g305(.A1(new_n389), .A2(new_n491), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n253), .A2(G119), .ZN(new_n493));
  INV_X1    g307(.A(G119), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n494), .A2(G128), .ZN(new_n495));
  AOI22_X1  g309(.A1(KEYINPUT74), .A2(new_n493), .B1(new_n495), .B2(KEYINPUT23), .ZN(new_n496));
  OR2_X1    g310(.A1(new_n493), .A2(KEYINPUT74), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  NAND3_X1  g312(.A1(new_n253), .A2(KEYINPUT23), .A3(G119), .ZN(new_n499));
  XNOR2_X1  g313(.A(new_n499), .B(KEYINPUT73), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n498), .A2(new_n500), .ZN(new_n501));
  NOR2_X1   g315(.A1(new_n501), .A2(G110), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n493), .A2(new_n495), .ZN(new_n503));
  XNOR2_X1  g317(.A(KEYINPUT24), .B(G110), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  XNOR2_X1  g319(.A(new_n505), .B(KEYINPUT75), .ZN(new_n506));
  OAI21_X1  g320(.A(new_n492), .B1(new_n502), .B2(new_n506), .ZN(new_n507));
  NOR2_X1   g321(.A1(new_n503), .A2(new_n504), .ZN(new_n508));
  AOI21_X1  g322(.A(new_n508), .B1(new_n501), .B2(G110), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n509), .A2(new_n390), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n507), .A2(new_n510), .ZN(new_n511));
  NAND3_X1  g325(.A1(new_n302), .A2(G221), .A3(G234), .ZN(new_n512));
  XNOR2_X1  g326(.A(KEYINPUT22), .B(G137), .ZN(new_n513));
  XNOR2_X1  g327(.A(new_n512), .B(new_n513), .ZN(new_n514));
  INV_X1    g328(.A(new_n514), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n511), .A2(new_n515), .ZN(new_n516));
  NAND3_X1  g330(.A1(new_n507), .A2(new_n510), .A3(new_n514), .ZN(new_n517));
  NAND3_X1  g331(.A1(new_n516), .A2(new_n447), .A3(new_n517), .ZN(new_n518));
  INV_X1    g332(.A(KEYINPUT25), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  NAND4_X1  g334(.A1(new_n516), .A2(KEYINPUT25), .A3(new_n447), .A4(new_n517), .ZN(new_n521));
  AOI21_X1  g335(.A(new_n490), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n516), .A2(new_n517), .ZN(new_n523));
  NOR2_X1   g337(.A1(new_n489), .A2(G902), .ZN(new_n524));
  INV_X1    g338(.A(new_n524), .ZN(new_n525));
  NOR2_X1   g339(.A1(new_n523), .A2(new_n525), .ZN(new_n526));
  NOR2_X1   g340(.A1(new_n522), .A2(new_n526), .ZN(new_n527));
  INV_X1    g341(.A(KEYINPUT76), .ZN(new_n528));
  NOR2_X1   g342(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  NOR3_X1   g343(.A1(new_n522), .A2(KEYINPUT76), .A3(new_n526), .ZN(new_n530));
  OR2_X1    g344(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n341), .A2(new_n355), .ZN(new_n532));
  INV_X1    g346(.A(KEYINPUT68), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n323), .A2(G134), .ZN(new_n534));
  AND2_X1   g348(.A1(new_n534), .A2(new_n326), .ZN(new_n535));
  OAI21_X1  g349(.A(new_n533), .B1(new_n535), .B2(new_n328), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n534), .A2(new_n326), .ZN(new_n537));
  NAND3_X1  g351(.A1(new_n537), .A2(KEYINPUT68), .A3(G131), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n536), .A2(new_n538), .ZN(new_n539));
  NAND3_X1  g353(.A1(new_n335), .A2(new_n278), .A3(new_n539), .ZN(new_n540));
  NAND3_X1  g354(.A1(new_n532), .A2(new_n225), .A3(new_n540), .ZN(new_n541));
  INV_X1    g355(.A(KEYINPUT70), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  INV_X1    g357(.A(new_n264), .ZN(new_n544));
  OAI21_X1  g358(.A(new_n544), .B1(new_n316), .B2(G146), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n545), .A2(new_n276), .ZN(new_n546));
  AOI22_X1  g360(.A1(new_n546), .A2(new_n274), .B1(new_n536), .B2(new_n538), .ZN(new_n547));
  AOI22_X1  g361(.A1(new_n355), .A2(new_n341), .B1(new_n547), .B2(new_n335), .ZN(new_n548));
  NAND3_X1  g362(.A1(new_n548), .A2(KEYINPUT70), .A3(new_n225), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n543), .A2(new_n549), .ZN(new_n550));
  INV_X1    g364(.A(new_n540), .ZN(new_n551));
  AOI21_X1  g365(.A(new_n271), .B1(new_n335), .B2(new_n340), .ZN(new_n552));
  OAI21_X1  g366(.A(KEYINPUT30), .B1(new_n551), .B2(new_n552), .ZN(new_n553));
  INV_X1    g367(.A(KEYINPUT30), .ZN(new_n554));
  NAND3_X1  g368(.A1(new_n532), .A2(new_n554), .A3(new_n540), .ZN(new_n555));
  AOI21_X1  g369(.A(new_n225), .B1(new_n553), .B2(new_n555), .ZN(new_n556));
  NOR2_X1   g370(.A1(new_n550), .A2(new_n556), .ZN(new_n557));
  INV_X1    g371(.A(KEYINPUT31), .ZN(new_n558));
  NAND3_X1  g372(.A1(new_n302), .A2(G210), .A3(new_n395), .ZN(new_n559));
  XNOR2_X1  g373(.A(new_n559), .B(KEYINPUT27), .ZN(new_n560));
  XNOR2_X1  g374(.A(KEYINPUT26), .B(G101), .ZN(new_n561));
  XNOR2_X1  g375(.A(new_n560), .B(new_n561), .ZN(new_n562));
  NAND3_X1  g376(.A1(new_n557), .A2(new_n558), .A3(new_n562), .ZN(new_n563));
  NOR3_X1   g377(.A1(new_n551), .A2(new_n552), .A3(KEYINPUT30), .ZN(new_n564));
  AOI21_X1  g378(.A(new_n554), .B1(new_n532), .B2(new_n540), .ZN(new_n565));
  OAI21_X1  g379(.A(new_n226), .B1(new_n564), .B2(new_n565), .ZN(new_n566));
  NAND4_X1  g380(.A1(new_n566), .A2(new_n562), .A3(new_n543), .A4(new_n549), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n567), .A2(KEYINPUT31), .ZN(new_n568));
  AOI21_X1  g382(.A(KEYINPUT28), .B1(new_n548), .B2(new_n225), .ZN(new_n569));
  OAI21_X1  g383(.A(KEYINPUT72), .B1(new_n548), .B2(new_n225), .ZN(new_n570));
  INV_X1    g384(.A(KEYINPUT72), .ZN(new_n571));
  OAI211_X1 g385(.A(new_n571), .B(new_n226), .C1(new_n551), .C2(new_n552), .ZN(new_n572));
  NAND4_X1  g386(.A1(new_n570), .A2(new_n543), .A3(new_n549), .A4(new_n572), .ZN(new_n573));
  AOI21_X1  g387(.A(new_n569), .B1(new_n573), .B2(KEYINPUT28), .ZN(new_n574));
  OAI211_X1 g388(.A(new_n563), .B(new_n568), .C1(new_n562), .C2(new_n574), .ZN(new_n575));
  NOR2_X1   g389(.A1(G472), .A2(G902), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n577), .A2(KEYINPUT32), .ZN(new_n578));
  INV_X1    g392(.A(KEYINPUT32), .ZN(new_n579));
  NAND3_X1  g393(.A1(new_n575), .A2(new_n579), .A3(new_n576), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n578), .A2(new_n580), .ZN(new_n581));
  OAI21_X1  g395(.A(new_n226), .B1(new_n551), .B2(new_n552), .ZN(new_n582));
  NAND3_X1  g396(.A1(new_n543), .A2(new_n549), .A3(new_n582), .ZN(new_n583));
  AOI21_X1  g397(.A(new_n569), .B1(new_n583), .B2(KEYINPUT28), .ZN(new_n584));
  INV_X1    g398(.A(new_n562), .ZN(new_n585));
  INV_X1    g399(.A(KEYINPUT29), .ZN(new_n586));
  NOR2_X1   g400(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  AOI21_X1  g401(.A(G902), .B1(new_n584), .B2(new_n587), .ZN(new_n588));
  AND2_X1   g402(.A1(new_n574), .A2(new_n562), .ZN(new_n589));
  OAI21_X1  g403(.A(new_n586), .B1(new_n557), .B2(new_n562), .ZN(new_n590));
  OAI21_X1  g404(.A(new_n588), .B1(new_n589), .B2(new_n590), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n591), .A2(G472), .ZN(new_n592));
  AOI21_X1  g406(.A(new_n531), .B1(new_n581), .B2(new_n592), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n488), .A2(new_n593), .ZN(new_n594));
  XNOR2_X1  g408(.A(new_n594), .B(G101), .ZN(G3));
  OAI211_X1 g409(.A(new_n187), .B(new_n486), .C1(new_n294), .C2(new_n295), .ZN(new_n596));
  INV_X1    g410(.A(KEYINPUT33), .ZN(new_n597));
  OR2_X1    g411(.A1(new_n474), .A2(new_n597), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n474), .A2(new_n597), .ZN(new_n599));
  NAND3_X1  g413(.A1(new_n598), .A2(G478), .A3(new_n599), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n475), .A2(new_n476), .ZN(new_n601));
  NOR2_X1   g415(.A1(new_n476), .A2(new_n447), .ZN(new_n602));
  INV_X1    g416(.A(new_n602), .ZN(new_n603));
  NAND3_X1  g417(.A1(new_n600), .A2(new_n601), .A3(new_n603), .ZN(new_n604));
  INV_X1    g418(.A(new_n604), .ZN(new_n605));
  AND3_X1   g419(.A1(new_n438), .A2(new_n442), .A3(new_n439), .ZN(new_n606));
  NOR3_X1   g420(.A1(new_n606), .A2(new_n445), .A3(new_n446), .ZN(new_n607));
  NAND3_X1  g421(.A1(new_n440), .A2(KEYINPUT92), .A3(new_n446), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n451), .A2(new_n452), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  OAI21_X1  g424(.A(new_n605), .B1(new_n607), .B2(new_n610), .ZN(new_n611));
  NOR2_X1   g425(.A1(new_n596), .A2(new_n611), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n575), .A2(new_n447), .ZN(new_n613));
  AOI22_X1  g427(.A1(new_n613), .A2(G472), .B1(new_n576), .B2(new_n575), .ZN(new_n614));
  NOR2_X1   g428(.A1(new_n529), .A2(new_n530), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  NOR2_X1   g430(.A1(new_n616), .A2(new_n382), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n612), .A2(new_n617), .ZN(new_n618));
  XOR2_X1   g432(.A(KEYINPUT34), .B(G104), .Z(new_n619));
  XNOR2_X1  g433(.A(new_n618), .B(new_n619), .ZN(G6));
  INV_X1    g434(.A(new_n478), .ZN(new_n621));
  NAND3_X1  g435(.A1(new_n444), .A2(new_n453), .A3(new_n621), .ZN(new_n622));
  OAI21_X1  g436(.A(KEYINPUT95), .B1(new_n596), .B2(new_n622), .ZN(new_n623));
  INV_X1    g437(.A(new_n187), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n284), .A2(new_n292), .ZN(new_n625));
  INV_X1    g439(.A(new_n293), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  NAND3_X1  g441(.A1(new_n284), .A2(new_n292), .A3(new_n293), .ZN(new_n628));
  AOI21_X1  g442(.A(new_n624), .B1(new_n627), .B2(new_n628), .ZN(new_n629));
  AND3_X1   g443(.A1(new_n444), .A2(new_n453), .A3(new_n621), .ZN(new_n630));
  INV_X1    g444(.A(KEYINPUT95), .ZN(new_n631));
  NAND4_X1  g445(.A1(new_n629), .A2(new_n630), .A3(new_n631), .A4(new_n486), .ZN(new_n632));
  NAND3_X1  g446(.A1(new_n623), .A2(new_n632), .A3(new_n617), .ZN(new_n633));
  XOR2_X1   g447(.A(KEYINPUT35), .B(G107), .Z(new_n634));
  XNOR2_X1  g448(.A(new_n633), .B(new_n634), .ZN(G9));
  NOR2_X1   g449(.A1(new_n515), .A2(KEYINPUT36), .ZN(new_n636));
  XOR2_X1   g450(.A(new_n511), .B(new_n636), .Z(new_n637));
  NOR2_X1   g451(.A1(new_n637), .A2(new_n525), .ZN(new_n638));
  NOR2_X1   g452(.A1(new_n522), .A2(new_n638), .ZN(new_n639));
  INV_X1    g453(.A(new_n639), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n614), .A2(new_n640), .ZN(new_n641));
  INV_X1    g455(.A(KEYINPUT96), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  NAND3_X1  g457(.A1(new_n614), .A2(KEYINPUT96), .A3(new_n640), .ZN(new_n644));
  NAND3_X1  g458(.A1(new_n488), .A2(new_n643), .A3(new_n644), .ZN(new_n645));
  XNOR2_X1  g459(.A(KEYINPUT37), .B(G110), .ZN(new_n646));
  XNOR2_X1  g460(.A(new_n646), .B(KEYINPUT97), .ZN(new_n647));
  XNOR2_X1  g461(.A(new_n645), .B(new_n647), .ZN(G12));
  NOR2_X1   g462(.A1(new_n296), .A2(new_n382), .ZN(new_n649));
  AOI21_X1  g463(.A(new_n639), .B1(new_n581), .B2(new_n592), .ZN(new_n650));
  AND2_X1   g464(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  NAND2_X1  g465(.A1(new_n484), .A2(new_n480), .ZN(new_n652));
  XOR2_X1   g466(.A(new_n652), .B(KEYINPUT98), .Z(new_n653));
  NOR2_X1   g467(.A1(new_n481), .A2(G900), .ZN(new_n654));
  NOR2_X1   g468(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  NOR2_X1   g469(.A1(new_n622), .A2(new_n655), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n651), .A2(new_n656), .ZN(new_n657));
  XNOR2_X1  g471(.A(new_n657), .B(G128), .ZN(G30));
  INV_X1    g472(.A(new_n557), .ZN(new_n659));
  NAND2_X1  g473(.A1(new_n659), .A2(new_n562), .ZN(new_n660));
  OAI211_X1 g474(.A(new_n660), .B(new_n447), .C1(new_n562), .C2(new_n583), .ZN(new_n661));
  AOI21_X1  g475(.A(KEYINPUT99), .B1(new_n661), .B2(G472), .ZN(new_n662));
  AND3_X1   g476(.A1(new_n661), .A2(KEYINPUT99), .A3(G472), .ZN(new_n663));
  OAI21_X1  g477(.A(new_n581), .B1(new_n662), .B2(new_n663), .ZN(new_n664));
  NAND3_X1  g478(.A1(new_n664), .A2(new_n187), .A3(new_n639), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n444), .A2(new_n453), .ZN(new_n666));
  NAND2_X1  g480(.A1(new_n666), .A2(new_n621), .ZN(new_n667));
  NOR2_X1   g481(.A1(new_n665), .A2(new_n667), .ZN(new_n668));
  AND2_X1   g482(.A1(new_n379), .A2(new_n380), .ZN(new_n669));
  NAND2_X1  g483(.A1(new_n361), .A2(new_n373), .ZN(new_n670));
  INV_X1    g484(.A(G469), .ZN(new_n671));
  NAND3_X1  g485(.A1(new_n670), .A2(new_n671), .A3(new_n447), .ZN(new_n672));
  AOI21_X1  g486(.A(new_n300), .B1(new_n669), .B2(new_n672), .ZN(new_n673));
  XOR2_X1   g487(.A(new_n655), .B(KEYINPUT39), .Z(new_n674));
  NAND2_X1  g488(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  OR2_X1    g489(.A1(new_n675), .A2(KEYINPUT40), .ZN(new_n676));
  NAND2_X1  g490(.A1(new_n675), .A2(KEYINPUT40), .ZN(new_n677));
  NAND2_X1  g491(.A1(new_n627), .A2(new_n628), .ZN(new_n678));
  XNOR2_X1  g492(.A(new_n678), .B(KEYINPUT38), .ZN(new_n679));
  NAND4_X1  g493(.A1(new_n668), .A2(new_n676), .A3(new_n677), .A4(new_n679), .ZN(new_n680));
  XNOR2_X1  g494(.A(new_n680), .B(new_n261), .ZN(G45));
  INV_X1    g495(.A(new_n655), .ZN(new_n682));
  OAI211_X1 g496(.A(new_n605), .B(new_n682), .C1(new_n607), .C2(new_n610), .ZN(new_n683));
  INV_X1    g497(.A(new_n683), .ZN(new_n684));
  NAND2_X1  g498(.A1(new_n651), .A2(new_n684), .ZN(new_n685));
  XNOR2_X1  g499(.A(new_n685), .B(G146), .ZN(G48));
  AOI21_X1  g500(.A(new_n372), .B1(new_n377), .B2(new_n362), .ZN(new_n687));
  AND3_X1   g501(.A1(new_n362), .A2(new_n372), .A3(new_n371), .ZN(new_n688));
  OAI21_X1  g502(.A(new_n447), .B1(new_n687), .B2(new_n688), .ZN(new_n689));
  INV_X1    g503(.A(KEYINPUT100), .ZN(new_n690));
  NOR2_X1   g504(.A1(new_n690), .A2(new_n671), .ZN(new_n691));
  NAND2_X1  g505(.A1(new_n689), .A2(new_n691), .ZN(new_n692));
  OAI221_X1 g506(.A(new_n447), .B1(new_n690), .B2(new_n671), .C1(new_n687), .C2(new_n688), .ZN(new_n693));
  NAND3_X1  g507(.A1(new_n692), .A2(new_n693), .A3(new_n301), .ZN(new_n694));
  INV_X1    g508(.A(KEYINPUT101), .ZN(new_n695));
  XNOR2_X1  g509(.A(new_n694), .B(new_n695), .ZN(new_n696));
  NAND3_X1  g510(.A1(new_n696), .A2(new_n593), .A3(new_n612), .ZN(new_n697));
  XNOR2_X1  g511(.A(new_n697), .B(KEYINPUT102), .ZN(new_n698));
  XNOR2_X1  g512(.A(KEYINPUT41), .B(G113), .ZN(new_n699));
  XNOR2_X1  g513(.A(new_n698), .B(new_n699), .ZN(G15));
  NAND4_X1  g514(.A1(new_n696), .A2(new_n593), .A3(new_n623), .A4(new_n632), .ZN(new_n701));
  XNOR2_X1  g515(.A(new_n701), .B(G116), .ZN(G18));
  NOR2_X1   g516(.A1(new_n296), .A2(new_n694), .ZN(new_n703));
  INV_X1    g517(.A(new_n487), .ZN(new_n704));
  NAND3_X1  g518(.A1(new_n703), .A2(new_n704), .A3(new_n650), .ZN(new_n705));
  XNOR2_X1  g519(.A(new_n705), .B(G119), .ZN(G21));
  NOR2_X1   g520(.A1(new_n667), .A2(new_n296), .ZN(new_n707));
  XOR2_X1   g521(.A(new_n576), .B(KEYINPUT103), .Z(new_n708));
  OAI21_X1  g522(.A(new_n568), .B1(new_n562), .B2(new_n584), .ZN(new_n709));
  INV_X1    g523(.A(KEYINPUT104), .ZN(new_n710));
  OAI21_X1  g524(.A(new_n563), .B1(new_n709), .B2(new_n710), .ZN(new_n711));
  OR2_X1    g525(.A1(new_n584), .A2(new_n562), .ZN(new_n712));
  AOI21_X1  g526(.A(KEYINPUT104), .B1(new_n712), .B2(new_n568), .ZN(new_n713));
  OAI21_X1  g527(.A(new_n708), .B1(new_n711), .B2(new_n713), .ZN(new_n714));
  INV_X1    g528(.A(KEYINPUT106), .ZN(new_n715));
  XNOR2_X1  g529(.A(new_n527), .B(new_n715), .ZN(new_n716));
  AOI21_X1  g530(.A(KEYINPUT105), .B1(new_n613), .B2(G472), .ZN(new_n717));
  INV_X1    g531(.A(KEYINPUT105), .ZN(new_n718));
  INV_X1    g532(.A(G472), .ZN(new_n719));
  AOI211_X1 g533(.A(new_n718), .B(new_n719), .C1(new_n575), .C2(new_n447), .ZN(new_n720));
  OAI211_X1 g534(.A(new_n714), .B(new_n716), .C1(new_n717), .C2(new_n720), .ZN(new_n721));
  NOR2_X1   g535(.A1(new_n721), .A2(new_n485), .ZN(new_n722));
  NAND3_X1  g536(.A1(new_n696), .A2(new_n707), .A3(new_n722), .ZN(new_n723));
  XNOR2_X1  g537(.A(new_n723), .B(G122), .ZN(G24));
  OAI211_X1 g538(.A(new_n714), .B(new_n640), .C1(new_n717), .C2(new_n720), .ZN(new_n725));
  INV_X1    g539(.A(new_n725), .ZN(new_n726));
  NAND2_X1  g540(.A1(new_n683), .A2(KEYINPUT107), .ZN(new_n727));
  AOI21_X1  g541(.A(new_n604), .B1(new_n444), .B2(new_n453), .ZN(new_n728));
  INV_X1    g542(.A(KEYINPUT107), .ZN(new_n729));
  NAND3_X1  g543(.A1(new_n728), .A2(new_n729), .A3(new_n682), .ZN(new_n730));
  NAND4_X1  g544(.A1(new_n726), .A2(new_n703), .A3(new_n727), .A4(new_n730), .ZN(new_n731));
  XNOR2_X1  g545(.A(new_n731), .B(G125), .ZN(G27));
  NOR2_X1   g546(.A1(new_n683), .A2(KEYINPUT107), .ZN(new_n733));
  AOI21_X1  g547(.A(new_n729), .B1(new_n728), .B2(new_n682), .ZN(new_n734));
  NOR2_X1   g548(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  NAND3_X1  g549(.A1(new_n627), .A2(new_n187), .A3(new_n628), .ZN(new_n736));
  NOR2_X1   g550(.A1(new_n736), .A2(new_n382), .ZN(new_n737));
  INV_X1    g551(.A(new_n580), .ZN(new_n738));
  AOI21_X1  g552(.A(new_n579), .B1(new_n575), .B2(new_n576), .ZN(new_n739));
  OAI21_X1  g553(.A(new_n592), .B1(new_n738), .B2(new_n739), .ZN(new_n740));
  AND2_X1   g554(.A1(new_n740), .A2(new_n716), .ZN(new_n741));
  NAND4_X1  g555(.A1(new_n735), .A2(KEYINPUT42), .A3(new_n737), .A4(new_n741), .ZN(new_n742));
  INV_X1    g556(.A(KEYINPUT42), .ZN(new_n743));
  NAND4_X1  g557(.A1(new_n737), .A2(new_n727), .A3(new_n593), .A4(new_n730), .ZN(new_n744));
  OAI21_X1  g558(.A(new_n743), .B1(new_n744), .B2(KEYINPUT108), .ZN(new_n745));
  INV_X1    g559(.A(KEYINPUT108), .ZN(new_n746));
  NOR3_X1   g560(.A1(new_n294), .A2(new_n295), .A3(new_n624), .ZN(new_n747));
  AND4_X1   g561(.A1(new_n740), .A2(new_n673), .A3(new_n747), .A4(new_n615), .ZN(new_n748));
  AOI21_X1  g562(.A(new_n746), .B1(new_n735), .B2(new_n748), .ZN(new_n749));
  OAI21_X1  g563(.A(new_n742), .B1(new_n745), .B2(new_n749), .ZN(new_n750));
  INV_X1    g564(.A(KEYINPUT109), .ZN(new_n751));
  NAND2_X1  g565(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  OAI211_X1 g566(.A(new_n742), .B(KEYINPUT109), .C1(new_n745), .C2(new_n749), .ZN(new_n753));
  AND2_X1   g567(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  XNOR2_X1  g568(.A(new_n754), .B(G131), .ZN(G33));
  NAND3_X1  g569(.A1(new_n737), .A2(new_n593), .A3(new_n656), .ZN(new_n756));
  XNOR2_X1  g570(.A(KEYINPUT110), .B(G134), .ZN(new_n757));
  XNOR2_X1  g571(.A(new_n756), .B(new_n757), .ZN(G36));
  NOR2_X1   g572(.A1(new_n607), .A2(new_n610), .ZN(new_n759));
  NAND2_X1  g573(.A1(new_n759), .A2(new_n605), .ZN(new_n760));
  NAND2_X1  g574(.A1(KEYINPUT111), .A2(KEYINPUT43), .ZN(new_n761));
  NAND2_X1  g575(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  XNOR2_X1  g576(.A(KEYINPUT111), .B(KEYINPUT43), .ZN(new_n763));
  NAND3_X1  g577(.A1(new_n759), .A2(new_n605), .A3(new_n763), .ZN(new_n764));
  AOI211_X1 g578(.A(new_n614), .B(new_n639), .C1(new_n762), .C2(new_n764), .ZN(new_n765));
  AND2_X1   g579(.A1(new_n765), .A2(KEYINPUT44), .ZN(new_n766));
  OAI21_X1  g580(.A(new_n747), .B1(new_n765), .B2(KEYINPUT44), .ZN(new_n767));
  NAND2_X1  g581(.A1(new_n376), .A2(new_n378), .ZN(new_n768));
  INV_X1    g582(.A(KEYINPUT45), .ZN(new_n769));
  AOI21_X1  g583(.A(new_n671), .B1(new_n768), .B2(new_n769), .ZN(new_n770));
  OAI21_X1  g584(.A(new_n770), .B1(new_n769), .B2(new_n768), .ZN(new_n771));
  AOI21_X1  g585(.A(KEYINPUT46), .B1(new_n771), .B2(new_n380), .ZN(new_n772));
  NOR2_X1   g586(.A1(new_n772), .A2(new_n374), .ZN(new_n773));
  NAND3_X1  g587(.A1(new_n771), .A2(KEYINPUT46), .A3(new_n380), .ZN(new_n774));
  NAND2_X1  g588(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  NAND3_X1  g589(.A1(new_n775), .A2(new_n301), .A3(new_n674), .ZN(new_n776));
  NOR3_X1   g590(.A1(new_n766), .A2(new_n767), .A3(new_n776), .ZN(new_n777));
  XNOR2_X1  g591(.A(new_n777), .B(new_n323), .ZN(G39));
  NAND2_X1  g592(.A1(new_n775), .A2(new_n301), .ZN(new_n779));
  INV_X1    g593(.A(KEYINPUT47), .ZN(new_n780));
  XNOR2_X1  g594(.A(new_n779), .B(new_n780), .ZN(new_n781));
  NOR4_X1   g595(.A1(new_n740), .A2(new_n683), .A3(new_n736), .A4(new_n615), .ZN(new_n782));
  NAND2_X1  g596(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  XNOR2_X1  g597(.A(new_n783), .B(G140), .ZN(G42));
  INV_X1    g598(.A(new_n781), .ZN(new_n785));
  AND2_X1   g599(.A1(new_n692), .A2(new_n693), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n786), .A2(new_n300), .ZN(new_n787));
  NAND2_X1  g601(.A1(new_n785), .A2(new_n787), .ZN(new_n788));
  NAND2_X1  g602(.A1(new_n762), .A2(new_n764), .ZN(new_n789));
  AND2_X1   g603(.A1(new_n789), .A2(new_n653), .ZN(new_n790));
  INV_X1    g604(.A(new_n721), .ZN(new_n791));
  NAND2_X1  g605(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  INV_X1    g606(.A(new_n792), .ZN(new_n793));
  NAND3_X1  g607(.A1(new_n788), .A2(new_n747), .A3(new_n793), .ZN(new_n794));
  NOR3_X1   g608(.A1(new_n679), .A2(new_n187), .A3(new_n694), .ZN(new_n795));
  NAND2_X1  g609(.A1(new_n793), .A2(new_n795), .ZN(new_n796));
  INV_X1    g610(.A(KEYINPUT50), .ZN(new_n797));
  XNOR2_X1  g611(.A(new_n796), .B(new_n797), .ZN(new_n798));
  AND4_X1   g612(.A1(new_n301), .A2(new_n790), .A3(new_n786), .A4(new_n747), .ZN(new_n799));
  NAND3_X1  g613(.A1(new_n615), .A2(new_n480), .A3(new_n484), .ZN(new_n800));
  NOR4_X1   g614(.A1(new_n664), .A2(new_n800), .A3(new_n736), .A4(new_n694), .ZN(new_n801));
  XOR2_X1   g615(.A(new_n801), .B(KEYINPUT117), .Z(new_n802));
  NOR2_X1   g616(.A1(new_n666), .A2(new_n605), .ZN(new_n803));
  AOI22_X1  g617(.A1(new_n799), .A2(new_n726), .B1(new_n802), .B2(new_n803), .ZN(new_n804));
  NAND3_X1  g618(.A1(new_n794), .A2(new_n798), .A3(new_n804), .ZN(new_n805));
  INV_X1    g619(.A(KEYINPUT51), .ZN(new_n806));
  NAND2_X1  g620(.A1(new_n805), .A2(new_n806), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n799), .A2(new_n741), .ZN(new_n808));
  XOR2_X1   g622(.A(new_n808), .B(KEYINPUT48), .Z(new_n809));
  NAND2_X1  g623(.A1(new_n802), .A2(new_n728), .ZN(new_n810));
  NAND2_X1  g624(.A1(new_n793), .A2(new_n703), .ZN(new_n811));
  NAND3_X1  g625(.A1(new_n810), .A2(new_n811), .A3(new_n484), .ZN(new_n812));
  NOR2_X1   g626(.A1(new_n809), .A2(new_n812), .ZN(new_n813));
  NAND4_X1  g627(.A1(new_n794), .A2(KEYINPUT51), .A3(new_n798), .A4(new_n804), .ZN(new_n814));
  NAND3_X1  g628(.A1(new_n807), .A2(new_n813), .A3(new_n814), .ZN(new_n815));
  NAND4_X1  g629(.A1(new_n701), .A2(new_n697), .A3(new_n723), .A4(new_n705), .ZN(new_n816));
  AOI22_X1  g630(.A1(new_n488), .A2(new_n593), .B1(new_n612), .B2(new_n617), .ZN(new_n817));
  OAI21_X1  g631(.A(KEYINPUT112), .B1(new_n596), .B2(new_n622), .ZN(new_n818));
  INV_X1    g632(.A(KEYINPUT112), .ZN(new_n819));
  NAND4_X1  g633(.A1(new_n629), .A2(new_n630), .A3(new_n819), .A4(new_n486), .ZN(new_n820));
  NAND3_X1  g634(.A1(new_n818), .A2(new_n820), .A3(new_n617), .ZN(new_n821));
  NAND4_X1  g635(.A1(new_n817), .A2(new_n645), .A3(new_n756), .A4(new_n821), .ZN(new_n822));
  INV_X1    g636(.A(new_n737), .ZN(new_n823));
  NAND3_X1  g637(.A1(new_n726), .A2(new_n727), .A3(new_n730), .ZN(new_n824));
  NAND4_X1  g638(.A1(new_n650), .A2(new_n478), .A3(new_n759), .A4(new_n682), .ZN(new_n825));
  AOI21_X1  g639(.A(new_n823), .B1(new_n824), .B2(new_n825), .ZN(new_n826));
  NOR3_X1   g640(.A1(new_n816), .A2(new_n822), .A3(new_n826), .ZN(new_n827));
  AND3_X1   g641(.A1(new_n827), .A2(new_n752), .A3(new_n753), .ZN(new_n828));
  INV_X1    g642(.A(KEYINPUT53), .ZN(new_n829));
  OAI211_X1 g643(.A(new_n649), .B(new_n650), .C1(new_n684), .C2(new_n656), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n639), .A2(new_n682), .ZN(new_n831));
  XNOR2_X1  g645(.A(new_n831), .B(KEYINPUT113), .ZN(new_n832));
  NAND4_X1  g646(.A1(new_n707), .A2(new_n673), .A3(new_n664), .A4(new_n832), .ZN(new_n833));
  NAND3_X1  g647(.A1(new_n731), .A2(new_n830), .A3(new_n833), .ZN(new_n834));
  INV_X1    g648(.A(KEYINPUT52), .ZN(new_n835));
  NAND2_X1  g649(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  NAND4_X1  g650(.A1(new_n731), .A2(new_n830), .A3(new_n833), .A4(KEYINPUT52), .ZN(new_n837));
  NAND2_X1  g651(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  NAND3_X1  g652(.A1(new_n828), .A2(new_n829), .A3(new_n838), .ZN(new_n839));
  AOI21_X1  g653(.A(KEYINPUT114), .B1(new_n836), .B2(new_n837), .ZN(new_n840));
  INV_X1    g654(.A(new_n840), .ZN(new_n841));
  NAND3_X1  g655(.A1(new_n836), .A2(KEYINPUT114), .A3(new_n837), .ZN(new_n842));
  NAND2_X1  g656(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  NAND3_X1  g657(.A1(new_n827), .A2(new_n752), .A3(new_n753), .ZN(new_n844));
  NOR2_X1   g658(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  OAI211_X1 g659(.A(new_n839), .B(KEYINPUT54), .C1(new_n845), .C2(new_n829), .ZN(new_n846));
  INV_X1    g660(.A(new_n816), .ZN(new_n847));
  NAND2_X1  g661(.A1(new_n847), .A2(new_n750), .ZN(new_n848));
  NAND2_X1  g662(.A1(new_n848), .A2(KEYINPUT116), .ZN(new_n849));
  INV_X1    g663(.A(KEYINPUT116), .ZN(new_n850));
  NAND3_X1  g664(.A1(new_n847), .A2(new_n750), .A3(new_n850), .ZN(new_n851));
  NAND2_X1  g665(.A1(new_n849), .A2(new_n851), .ZN(new_n852));
  AND3_X1   g666(.A1(new_n817), .A2(new_n645), .A3(new_n821), .ZN(new_n853));
  INV_X1    g667(.A(KEYINPUT115), .ZN(new_n854));
  INV_X1    g668(.A(new_n826), .ZN(new_n855));
  NAND4_X1  g669(.A1(new_n853), .A2(new_n854), .A3(new_n855), .A4(new_n756), .ZN(new_n856));
  OAI21_X1  g670(.A(KEYINPUT115), .B1(new_n822), .B2(new_n826), .ZN(new_n857));
  AND3_X1   g671(.A1(new_n857), .A2(new_n838), .A3(KEYINPUT53), .ZN(new_n858));
  NAND3_X1  g672(.A1(new_n852), .A2(new_n856), .A3(new_n858), .ZN(new_n859));
  OAI21_X1  g673(.A(new_n829), .B1(new_n843), .B2(new_n844), .ZN(new_n860));
  INV_X1    g674(.A(KEYINPUT54), .ZN(new_n861));
  NAND3_X1  g675(.A1(new_n859), .A2(new_n860), .A3(new_n861), .ZN(new_n862));
  NAND2_X1  g676(.A1(new_n846), .A2(new_n862), .ZN(new_n863));
  OAI22_X1  g677(.A1(new_n815), .A2(new_n863), .B1(G952), .B2(G953), .ZN(new_n864));
  XOR2_X1   g678(.A(new_n786), .B(KEYINPUT49), .Z(new_n865));
  NAND3_X1  g679(.A1(new_n716), .A2(new_n187), .A3(new_n301), .ZN(new_n866));
  OR4_X1    g680(.A1(new_n664), .A2(new_n865), .A3(new_n760), .A4(new_n866), .ZN(new_n867));
  OAI21_X1  g681(.A(new_n864), .B1(new_n679), .B2(new_n867), .ZN(G75));
  AOI21_X1  g682(.A(new_n447), .B1(new_n859), .B2(new_n860), .ZN(new_n869));
  INV_X1    g683(.A(KEYINPUT119), .ZN(new_n870));
  NAND3_X1  g684(.A1(new_n869), .A2(new_n870), .A3(G210), .ZN(new_n871));
  INV_X1    g685(.A(KEYINPUT56), .ZN(new_n872));
  NAND2_X1  g686(.A1(new_n244), .A2(new_n251), .ZN(new_n873));
  XOR2_X1   g687(.A(new_n873), .B(KEYINPUT118), .Z(new_n874));
  XNOR2_X1  g688(.A(new_n874), .B(KEYINPUT55), .ZN(new_n875));
  XNOR2_X1  g689(.A(new_n875), .B(new_n283), .ZN(new_n876));
  NAND3_X1  g690(.A1(new_n871), .A2(new_n872), .A3(new_n876), .ZN(new_n877));
  AOI21_X1  g691(.A(new_n870), .B1(new_n869), .B2(G210), .ZN(new_n878));
  NOR2_X1   g692(.A1(new_n877), .A2(new_n878), .ZN(new_n879));
  NOR2_X1   g693(.A1(new_n302), .A2(G952), .ZN(new_n880));
  INV_X1    g694(.A(new_n880), .ZN(new_n881));
  AOI21_X1  g695(.A(KEYINPUT56), .B1(new_n869), .B2(G210), .ZN(new_n882));
  OAI21_X1  g696(.A(new_n881), .B1(new_n882), .B2(new_n876), .ZN(new_n883));
  NOR2_X1   g697(.A1(new_n879), .A2(new_n883), .ZN(G51));
  INV_X1    g698(.A(new_n842), .ZN(new_n885));
  NOR2_X1   g699(.A1(new_n885), .A2(new_n840), .ZN(new_n886));
  AOI21_X1  g700(.A(KEYINPUT53), .B1(new_n828), .B2(new_n886), .ZN(new_n887));
  NAND4_X1  g701(.A1(new_n856), .A2(new_n857), .A3(KEYINPUT53), .A4(new_n838), .ZN(new_n888));
  AOI21_X1  g702(.A(new_n888), .B1(new_n851), .B2(new_n849), .ZN(new_n889));
  OAI21_X1  g703(.A(KEYINPUT54), .B1(new_n887), .B2(new_n889), .ZN(new_n890));
  INV_X1    g704(.A(KEYINPUT120), .ZN(new_n891));
  NAND3_X1  g705(.A1(new_n890), .A2(new_n891), .A3(new_n862), .ZN(new_n892));
  NAND2_X1  g706(.A1(new_n859), .A2(new_n860), .ZN(new_n893));
  NAND3_X1  g707(.A1(new_n893), .A2(KEYINPUT120), .A3(KEYINPUT54), .ZN(new_n894));
  XOR2_X1   g708(.A(new_n380), .B(KEYINPUT57), .Z(new_n895));
  NAND3_X1  g709(.A1(new_n892), .A2(new_n894), .A3(new_n895), .ZN(new_n896));
  NAND2_X1  g710(.A1(new_n896), .A2(new_n670), .ZN(new_n897));
  INV_X1    g711(.A(new_n869), .ZN(new_n898));
  OR2_X1    g712(.A1(new_n898), .A2(new_n771), .ZN(new_n899));
  AOI21_X1  g713(.A(new_n880), .B1(new_n897), .B2(new_n899), .ZN(G54));
  INV_X1    g714(.A(new_n438), .ZN(new_n901));
  NAND2_X1  g715(.A1(KEYINPUT58), .A2(G475), .ZN(new_n902));
  XOR2_X1   g716(.A(new_n902), .B(KEYINPUT121), .Z(new_n903));
  OAI21_X1  g717(.A(new_n901), .B1(new_n898), .B2(new_n903), .ZN(new_n904));
  NAND2_X1  g718(.A1(new_n904), .A2(new_n881), .ZN(new_n905));
  NOR3_X1   g719(.A1(new_n898), .A2(new_n901), .A3(new_n903), .ZN(new_n906));
  NOR2_X1   g720(.A1(new_n905), .A2(new_n906), .ZN(G60));
  XNOR2_X1  g721(.A(new_n602), .B(KEYINPUT59), .ZN(new_n908));
  AOI21_X1  g722(.A(new_n908), .B1(new_n846), .B2(new_n862), .ZN(new_n909));
  AND2_X1   g723(.A1(new_n598), .A2(new_n599), .ZN(new_n910));
  INV_X1    g724(.A(new_n910), .ZN(new_n911));
  OAI21_X1  g725(.A(new_n881), .B1(new_n909), .B2(new_n911), .ZN(new_n912));
  NOR2_X1   g726(.A1(new_n910), .A2(new_n908), .ZN(new_n913));
  NAND3_X1  g727(.A1(new_n892), .A2(new_n894), .A3(new_n913), .ZN(new_n914));
  INV_X1    g728(.A(KEYINPUT122), .ZN(new_n915));
  NAND2_X1  g729(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  NAND4_X1  g730(.A1(new_n892), .A2(KEYINPUT122), .A3(new_n894), .A4(new_n913), .ZN(new_n917));
  AOI21_X1  g731(.A(new_n912), .B1(new_n916), .B2(new_n917), .ZN(G63));
  INV_X1    g732(.A(KEYINPUT61), .ZN(new_n919));
  NAND2_X1  g733(.A1(G217), .A2(G902), .ZN(new_n920));
  XOR2_X1   g734(.A(new_n920), .B(KEYINPUT60), .Z(new_n921));
  NAND2_X1  g735(.A1(new_n893), .A2(new_n921), .ZN(new_n922));
  NAND2_X1  g736(.A1(new_n922), .A2(new_n523), .ZN(new_n923));
  NAND2_X1  g737(.A1(new_n923), .A2(new_n881), .ZN(new_n924));
  NOR2_X1   g738(.A1(new_n922), .A2(new_n637), .ZN(new_n925));
  OAI21_X1  g739(.A(new_n919), .B1(new_n924), .B2(new_n925), .ZN(new_n926));
  AOI21_X1  g740(.A(new_n880), .B1(new_n922), .B2(new_n523), .ZN(new_n927));
  OAI211_X1 g741(.A(new_n927), .B(KEYINPUT61), .C1(new_n637), .C2(new_n922), .ZN(new_n928));
  NAND2_X1  g742(.A1(new_n926), .A2(new_n928), .ZN(G66));
  INV_X1    g743(.A(G224), .ZN(new_n930));
  OAI21_X1  g744(.A(G953), .B1(new_n483), .B2(new_n930), .ZN(new_n931));
  AND2_X1   g745(.A1(new_n847), .A2(new_n853), .ZN(new_n932));
  OAI21_X1  g746(.A(new_n931), .B1(new_n932), .B2(new_n479), .ZN(new_n933));
  OAI21_X1  g747(.A(new_n874), .B1(G898), .B2(new_n302), .ZN(new_n934));
  XNOR2_X1  g748(.A(new_n933), .B(new_n934), .ZN(G69));
  NOR2_X1   g749(.A1(new_n564), .A2(new_n565), .ZN(new_n936));
  XNOR2_X1  g750(.A(new_n936), .B(new_n430), .ZN(new_n937));
  INV_X1    g751(.A(G227), .ZN(new_n938));
  AOI21_X1  g752(.A(new_n937), .B1(new_n938), .B2(new_n479), .ZN(new_n939));
  OR3_X1    g753(.A1(new_n766), .A2(new_n767), .A3(new_n776), .ZN(new_n940));
  NAND2_X1  g754(.A1(new_n731), .A2(new_n830), .ZN(new_n941));
  INV_X1    g755(.A(new_n941), .ZN(new_n942));
  NAND3_X1  g756(.A1(new_n940), .A2(KEYINPUT124), .A3(new_n942), .ZN(new_n943));
  INV_X1    g757(.A(KEYINPUT124), .ZN(new_n944));
  OAI21_X1  g758(.A(new_n944), .B1(new_n777), .B2(new_n941), .ZN(new_n945));
  NAND2_X1  g759(.A1(new_n943), .A2(new_n945), .ZN(new_n946));
  NAND2_X1  g760(.A1(new_n741), .A2(new_n707), .ZN(new_n947));
  OAI21_X1  g761(.A(new_n756), .B1(new_n776), .B2(new_n947), .ZN(new_n948));
  AOI21_X1  g762(.A(new_n948), .B1(new_n781), .B2(new_n782), .ZN(new_n949));
  AND3_X1   g763(.A1(new_n946), .A2(new_n754), .A3(new_n949), .ZN(new_n950));
  OAI21_X1  g764(.A(new_n939), .B1(new_n950), .B2(new_n479), .ZN(new_n951));
  INV_X1    g765(.A(G900), .ZN(new_n952));
  AOI21_X1  g766(.A(new_n952), .B1(new_n937), .B2(new_n938), .ZN(new_n953));
  NAND2_X1  g767(.A1(new_n611), .A2(new_n622), .ZN(new_n954));
  NAND3_X1  g768(.A1(new_n748), .A2(new_n674), .A3(new_n954), .ZN(new_n955));
  INV_X1    g769(.A(new_n955), .ZN(new_n956));
  NOR2_X1   g770(.A1(new_n777), .A2(new_n956), .ZN(new_n957));
  NAND2_X1  g771(.A1(new_n942), .A2(new_n680), .ZN(new_n958));
  AOI22_X1  g772(.A1(new_n781), .A2(new_n782), .B1(KEYINPUT62), .B2(new_n958), .ZN(new_n959));
  OR2_X1    g773(.A1(new_n958), .A2(KEYINPUT62), .ZN(new_n960));
  NAND3_X1  g774(.A1(new_n957), .A2(new_n959), .A3(new_n960), .ZN(new_n961));
  NAND2_X1  g775(.A1(new_n961), .A2(KEYINPUT123), .ZN(new_n962));
  INV_X1    g776(.A(KEYINPUT123), .ZN(new_n963));
  NAND4_X1  g777(.A1(new_n957), .A2(new_n959), .A3(new_n963), .A4(new_n960), .ZN(new_n964));
  AND2_X1   g778(.A1(new_n962), .A2(new_n964), .ZN(new_n965));
  NAND2_X1  g779(.A1(new_n937), .A2(new_n302), .ZN(new_n966));
  OAI221_X1 g780(.A(new_n951), .B1(new_n302), .B2(new_n953), .C1(new_n965), .C2(new_n966), .ZN(G72));
  NAND2_X1  g781(.A1(G472), .A2(G902), .ZN(new_n968));
  XOR2_X1   g782(.A(new_n968), .B(KEYINPUT63), .Z(new_n969));
  INV_X1    g783(.A(new_n969), .ZN(new_n970));
  NAND2_X1  g784(.A1(new_n659), .A2(new_n585), .ZN(new_n971));
  AOI21_X1  g785(.A(new_n970), .B1(new_n971), .B2(new_n567), .ZN(new_n972));
  OAI211_X1 g786(.A(new_n839), .B(new_n972), .C1(new_n845), .C2(new_n829), .ZN(new_n973));
  NAND3_X1  g787(.A1(new_n962), .A2(new_n932), .A3(new_n964), .ZN(new_n974));
  XOR2_X1   g788(.A(new_n969), .B(KEYINPUT125), .Z(new_n975));
  AND2_X1   g789(.A1(new_n974), .A2(new_n975), .ZN(new_n976));
  OAI211_X1 g790(.A(new_n881), .B(new_n973), .C1(new_n976), .C2(new_n660), .ZN(new_n977));
  NAND2_X1  g791(.A1(new_n557), .A2(new_n585), .ZN(new_n978));
  NAND4_X1  g792(.A1(new_n946), .A2(new_n949), .A3(new_n754), .A4(new_n932), .ZN(new_n979));
  NAND2_X1  g793(.A1(new_n979), .A2(new_n975), .ZN(new_n980));
  NAND2_X1  g794(.A1(new_n980), .A2(KEYINPUT126), .ZN(new_n981));
  INV_X1    g795(.A(KEYINPUT126), .ZN(new_n982));
  NAND3_X1  g796(.A1(new_n979), .A2(new_n982), .A3(new_n975), .ZN(new_n983));
  AOI21_X1  g797(.A(new_n978), .B1(new_n981), .B2(new_n983), .ZN(new_n984));
  NOR2_X1   g798(.A1(new_n977), .A2(new_n984), .ZN(G57));
endmodule


