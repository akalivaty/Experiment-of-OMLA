

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302,
         n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313,
         n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324,
         n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335,
         n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346,
         n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585;

  OR2_X1 U324 ( .A1(n540), .A2(n539), .ZN(n541) );
  NOR2_X1 U325 ( .A1(n544), .A2(n543), .ZN(n545) );
  XNOR2_X1 U326 ( .A(n302), .B(n301), .ZN(n309) );
  XNOR2_X1 U327 ( .A(n333), .B(n292), .ZN(n301) );
  XOR2_X1 U328 ( .A(n429), .B(n428), .Z(n495) );
  AND2_X1 U329 ( .A1(G228GAT), .A2(G233GAT), .ZN(n292) );
  INV_X1 U330 ( .A(KEYINPUT69), .ZN(n336) );
  INV_X1 U331 ( .A(KEYINPUT37), .ZN(n444) );
  XNOR2_X1 U332 ( .A(n337), .B(n336), .ZN(n338) );
  XNOR2_X1 U333 ( .A(n444), .B(KEYINPUT101), .ZN(n445) );
  XNOR2_X1 U334 ( .A(n339), .B(n338), .ZN(n340) );
  XNOR2_X1 U335 ( .A(n446), .B(n445), .ZN(n465) );
  NOR2_X2 U336 ( .A1(n550), .A2(n549), .ZN(n563) );
  XOR2_X1 U337 ( .A(KEYINPUT108), .B(n447), .Z(n496) );
  XOR2_X1 U338 ( .A(KEYINPUT28), .B(n310), .Z(n485) );
  XNOR2_X1 U339 ( .A(n449), .B(n448), .ZN(n450) );
  XNOR2_X1 U340 ( .A(n451), .B(n450), .ZN(G1339GAT) );
  XOR2_X1 U341 ( .A(KEYINPUT22), .B(KEYINPUT90), .Z(n294) );
  XNOR2_X1 U342 ( .A(KEYINPUT89), .B(KEYINPUT24), .ZN(n293) );
  XNOR2_X1 U343 ( .A(n294), .B(n293), .ZN(n298) );
  XOR2_X1 U344 ( .A(G50GAT), .B(G162GAT), .Z(n372) );
  XOR2_X1 U345 ( .A(G78GAT), .B(KEYINPUT23), .Z(n295) );
  XNOR2_X1 U346 ( .A(n372), .B(n295), .ZN(n296) );
  XOR2_X1 U347 ( .A(G22GAT), .B(G155GAT), .Z(n343) );
  XNOR2_X1 U348 ( .A(n296), .B(n343), .ZN(n297) );
  XOR2_X1 U349 ( .A(n298), .B(n297), .Z(n302) );
  XOR2_X1 U350 ( .A(G148GAT), .B(G204GAT), .Z(n300) );
  XNOR2_X1 U351 ( .A(G106GAT), .B(KEYINPUT70), .ZN(n299) );
  XNOR2_X1 U352 ( .A(n300), .B(n299), .ZN(n333) );
  XOR2_X1 U353 ( .A(KEYINPUT87), .B(G218GAT), .Z(n304) );
  XNOR2_X1 U354 ( .A(KEYINPUT21), .B(G211GAT), .ZN(n303) );
  XNOR2_X1 U355 ( .A(n304), .B(n303), .ZN(n305) );
  XOR2_X1 U356 ( .A(G197GAT), .B(n305), .Z(n406) );
  XOR2_X1 U357 ( .A(KEYINPUT88), .B(KEYINPUT3), .Z(n307) );
  XNOR2_X1 U358 ( .A(G141GAT), .B(KEYINPUT2), .ZN(n306) );
  XNOR2_X1 U359 ( .A(n307), .B(n306), .ZN(n385) );
  XNOR2_X1 U360 ( .A(n406), .B(n385), .ZN(n308) );
  XNOR2_X1 U361 ( .A(n309), .B(n308), .ZN(n546) );
  XOR2_X1 U362 ( .A(n546), .B(KEYINPUT66), .Z(n310) );
  XOR2_X1 U363 ( .A(G22GAT), .B(G141GAT), .Z(n312) );
  XNOR2_X1 U364 ( .A(G169GAT), .B(G113GAT), .ZN(n311) );
  XNOR2_X1 U365 ( .A(n312), .B(n311), .ZN(n322) );
  XOR2_X1 U366 ( .A(KEYINPUT29), .B(KEYINPUT30), .Z(n314) );
  XNOR2_X1 U367 ( .A(G197GAT), .B(G8GAT), .ZN(n313) );
  XNOR2_X1 U368 ( .A(n314), .B(n313), .ZN(n318) );
  XOR2_X1 U369 ( .A(G36GAT), .B(G50GAT), .Z(n316) );
  XOR2_X1 U370 ( .A(G15GAT), .B(G1GAT), .Z(n351) );
  XNOR2_X1 U371 ( .A(KEYINPUT67), .B(n351), .ZN(n315) );
  XNOR2_X1 U372 ( .A(n316), .B(n315), .ZN(n317) );
  XOR2_X1 U373 ( .A(n318), .B(n317), .Z(n320) );
  NAND2_X1 U374 ( .A1(G229GAT), .A2(G233GAT), .ZN(n319) );
  XNOR2_X1 U375 ( .A(n320), .B(n319), .ZN(n321) );
  XNOR2_X1 U376 ( .A(n322), .B(n321), .ZN(n326) );
  XOR2_X1 U377 ( .A(KEYINPUT7), .B(KEYINPUT68), .Z(n324) );
  XNOR2_X1 U378 ( .A(G43GAT), .B(G29GAT), .ZN(n323) );
  XNOR2_X1 U379 ( .A(n324), .B(n323), .ZN(n325) );
  XNOR2_X1 U380 ( .A(KEYINPUT8), .B(n325), .ZN(n373) );
  XOR2_X1 U381 ( .A(n326), .B(n373), .Z(n527) );
  INV_X1 U382 ( .A(n527), .ZN(n569) );
  XOR2_X1 U383 ( .A(G57GAT), .B(KEYINPUT13), .Z(n328) );
  XNOR2_X1 U384 ( .A(G71GAT), .B(G78GAT), .ZN(n327) );
  XNOR2_X1 U385 ( .A(n328), .B(n327), .ZN(n344) );
  XNOR2_X1 U386 ( .A(KEYINPUT31), .B(KEYINPUT33), .ZN(n330) );
  AND2_X1 U387 ( .A1(G230GAT), .A2(G233GAT), .ZN(n329) );
  XNOR2_X1 U388 ( .A(n330), .B(n329), .ZN(n331) );
  XOR2_X1 U389 ( .A(n331), .B(KEYINPUT32), .Z(n335) );
  XNOR2_X1 U390 ( .A(G176GAT), .B(G92GAT), .ZN(n332) );
  XNOR2_X1 U391 ( .A(n332), .B(G64GAT), .ZN(n398) );
  XNOR2_X1 U392 ( .A(n333), .B(n398), .ZN(n334) );
  XNOR2_X1 U393 ( .A(n335), .B(n334), .ZN(n339) );
  XOR2_X1 U394 ( .A(G99GAT), .B(G85GAT), .Z(n367) );
  XNOR2_X1 U395 ( .A(G120GAT), .B(n367), .ZN(n337) );
  XOR2_X1 U396 ( .A(n344), .B(n340), .Z(n574) );
  XOR2_X1 U397 ( .A(KEYINPUT41), .B(n574), .Z(n555) );
  INV_X1 U398 ( .A(n555), .ZN(n530) );
  NOR2_X1 U399 ( .A1(n569), .A2(n530), .ZN(n478) );
  XOR2_X1 U400 ( .A(KEYINPUT15), .B(G64GAT), .Z(n342) );
  XNOR2_X1 U401 ( .A(G127GAT), .B(G211GAT), .ZN(n341) );
  XNOR2_X1 U402 ( .A(n342), .B(n341), .ZN(n355) );
  XOR2_X1 U403 ( .A(n344), .B(n343), .Z(n346) );
  NAND2_X1 U404 ( .A1(G231GAT), .A2(G233GAT), .ZN(n345) );
  XNOR2_X1 U405 ( .A(n346), .B(n345), .ZN(n350) );
  XOR2_X1 U406 ( .A(KEYINPUT76), .B(KEYINPUT12), .Z(n348) );
  XNOR2_X1 U407 ( .A(KEYINPUT77), .B(KEYINPUT14), .ZN(n347) );
  XNOR2_X1 U408 ( .A(n348), .B(n347), .ZN(n349) );
  XOR2_X1 U409 ( .A(n350), .B(n349), .Z(n353) );
  XOR2_X1 U410 ( .A(G8GAT), .B(G183GAT), .Z(n400) );
  XNOR2_X1 U411 ( .A(n351), .B(n400), .ZN(n352) );
  XNOR2_X1 U412 ( .A(n353), .B(n352), .ZN(n354) );
  XNOR2_X1 U413 ( .A(n355), .B(n354), .ZN(n578) );
  INV_X1 U414 ( .A(n578), .ZN(n534) );
  XOR2_X1 U415 ( .A(KEYINPUT10), .B(KEYINPUT11), .Z(n357) );
  XNOR2_X1 U416 ( .A(KEYINPUT75), .B(KEYINPUT73), .ZN(n356) );
  XNOR2_X1 U417 ( .A(n357), .B(n356), .ZN(n361) );
  XOR2_X1 U418 ( .A(KEYINPUT65), .B(KEYINPUT72), .Z(n359) );
  XNOR2_X1 U419 ( .A(G134GAT), .B(G92GAT), .ZN(n358) );
  XNOR2_X1 U420 ( .A(n359), .B(n358), .ZN(n360) );
  XOR2_X1 U421 ( .A(n361), .B(n360), .Z(n366) );
  XOR2_X1 U422 ( .A(KEYINPUT9), .B(KEYINPUT71), .Z(n363) );
  NAND2_X1 U423 ( .A1(G232GAT), .A2(G233GAT), .ZN(n362) );
  XNOR2_X1 U424 ( .A(n363), .B(n362), .ZN(n364) );
  XNOR2_X1 U425 ( .A(KEYINPUT74), .B(n364), .ZN(n365) );
  XNOR2_X1 U426 ( .A(n366), .B(n365), .ZN(n371) );
  XOR2_X1 U427 ( .A(G36GAT), .B(G190GAT), .Z(n399) );
  XOR2_X1 U428 ( .A(n367), .B(n399), .Z(n369) );
  XNOR2_X1 U429 ( .A(G218GAT), .B(G106GAT), .ZN(n368) );
  XNOR2_X1 U430 ( .A(n369), .B(n368), .ZN(n370) );
  XOR2_X1 U431 ( .A(n371), .B(n370), .Z(n375) );
  XOR2_X1 U432 ( .A(n373), .B(n372), .Z(n374) );
  XOR2_X1 U433 ( .A(n375), .B(n374), .Z(n562) );
  XOR2_X1 U434 ( .A(KEYINPUT36), .B(n562), .Z(n582) );
  XOR2_X1 U435 ( .A(G155GAT), .B(G148GAT), .Z(n377) );
  XNOR2_X1 U436 ( .A(G29GAT), .B(G1GAT), .ZN(n376) );
  XNOR2_X1 U437 ( .A(n377), .B(n376), .ZN(n381) );
  XOR2_X1 U438 ( .A(KEYINPUT93), .B(KEYINPUT91), .Z(n379) );
  XNOR2_X1 U439 ( .A(G57GAT), .B(KEYINPUT1), .ZN(n378) );
  XNOR2_X1 U440 ( .A(n379), .B(n378), .ZN(n380) );
  XOR2_X1 U441 ( .A(n381), .B(n380), .Z(n387) );
  XOR2_X1 U442 ( .A(G85GAT), .B(G162GAT), .Z(n383) );
  NAND2_X1 U443 ( .A1(G225GAT), .A2(G233GAT), .ZN(n382) );
  XNOR2_X1 U444 ( .A(n383), .B(n382), .ZN(n384) );
  XNOR2_X1 U445 ( .A(n385), .B(n384), .ZN(n386) );
  XNOR2_X1 U446 ( .A(n387), .B(n386), .ZN(n397) );
  XOR2_X1 U447 ( .A(KEYINPUT80), .B(KEYINPUT79), .Z(n389) );
  XNOR2_X1 U448 ( .A(G134GAT), .B(KEYINPUT0), .ZN(n388) );
  XNOR2_X1 U449 ( .A(n389), .B(n388), .ZN(n390) );
  XOR2_X1 U450 ( .A(n390), .B(G127GAT), .Z(n392) );
  XNOR2_X1 U451 ( .A(G113GAT), .B(G120GAT), .ZN(n391) );
  XNOR2_X1 U452 ( .A(n392), .B(n391), .ZN(n425) );
  XOR2_X1 U453 ( .A(KEYINPUT5), .B(KEYINPUT92), .Z(n394) );
  XNOR2_X1 U454 ( .A(KEYINPUT4), .B(KEYINPUT6), .ZN(n393) );
  XNOR2_X1 U455 ( .A(n394), .B(n393), .ZN(n395) );
  XOR2_X1 U456 ( .A(n425), .B(n395), .Z(n396) );
  XNOR2_X1 U457 ( .A(n397), .B(n396), .ZN(n544) );
  XNOR2_X1 U458 ( .A(n399), .B(n398), .ZN(n401) );
  XNOR2_X1 U459 ( .A(n401), .B(n400), .ZN(n405) );
  XOR2_X1 U460 ( .A(KEYINPUT94), .B(KEYINPUT95), .Z(n403) );
  NAND2_X1 U461 ( .A1(G226GAT), .A2(G233GAT), .ZN(n402) );
  XNOR2_X1 U462 ( .A(n403), .B(n402), .ZN(n404) );
  XOR2_X1 U463 ( .A(n405), .B(n404), .Z(n408) );
  XNOR2_X1 U464 ( .A(n406), .B(G204GAT), .ZN(n407) );
  XNOR2_X1 U465 ( .A(n408), .B(n407), .ZN(n412) );
  XOR2_X1 U466 ( .A(KEYINPUT83), .B(KEYINPUT17), .Z(n410) );
  XNOR2_X1 U467 ( .A(KEYINPUT19), .B(KEYINPUT18), .ZN(n409) );
  XNOR2_X1 U468 ( .A(n410), .B(n409), .ZN(n411) );
  XNOR2_X1 U469 ( .A(G169GAT), .B(n411), .ZN(n428) );
  XOR2_X1 U470 ( .A(n412), .B(n428), .Z(n539) );
  XOR2_X1 U471 ( .A(n539), .B(KEYINPUT27), .Z(n436) );
  NAND2_X1 U472 ( .A1(n544), .A2(n436), .ZN(n511) );
  XOR2_X1 U473 ( .A(G71GAT), .B(G183GAT), .Z(n414) );
  XNOR2_X1 U474 ( .A(KEYINPUT85), .B(KEYINPUT82), .ZN(n413) );
  XNOR2_X1 U475 ( .A(n414), .B(n413), .ZN(n418) );
  XOR2_X1 U476 ( .A(G176GAT), .B(KEYINPUT84), .Z(n416) );
  XNOR2_X1 U477 ( .A(G15GAT), .B(KEYINPUT81), .ZN(n415) );
  XNOR2_X1 U478 ( .A(n416), .B(n415), .ZN(n417) );
  XOR2_X1 U479 ( .A(n418), .B(n417), .Z(n427) );
  XOR2_X1 U480 ( .A(KEYINPUT86), .B(G190GAT), .Z(n420) );
  XNOR2_X1 U481 ( .A(G43GAT), .B(G99GAT), .ZN(n419) );
  XNOR2_X1 U482 ( .A(n420), .B(n419), .ZN(n421) );
  XOR2_X1 U483 ( .A(KEYINPUT20), .B(n421), .Z(n423) );
  NAND2_X1 U484 ( .A1(G227GAT), .A2(G233GAT), .ZN(n422) );
  XNOR2_X1 U485 ( .A(n423), .B(n422), .ZN(n424) );
  XNOR2_X1 U486 ( .A(n425), .B(n424), .ZN(n426) );
  XNOR2_X1 U487 ( .A(n427), .B(n426), .ZN(n429) );
  INV_X1 U488 ( .A(n495), .ZN(n550) );
  INV_X1 U489 ( .A(n485), .ZN(n512) );
  NAND2_X1 U490 ( .A1(n550), .A2(n512), .ZN(n430) );
  NOR2_X1 U491 ( .A1(n511), .A2(n430), .ZN(n431) );
  XNOR2_X1 U492 ( .A(n431), .B(KEYINPUT96), .ZN(n442) );
  NOR2_X1 U493 ( .A1(n550), .A2(n539), .ZN(n432) );
  NOR2_X1 U494 ( .A1(n546), .A2(n432), .ZN(n433) );
  XOR2_X1 U495 ( .A(n433), .B(KEYINPUT98), .Z(n434) );
  XNOR2_X1 U496 ( .A(KEYINPUT25), .B(n434), .ZN(n439) );
  NAND2_X1 U497 ( .A1(n546), .A2(n550), .ZN(n435) );
  XOR2_X1 U498 ( .A(n435), .B(KEYINPUT26), .Z(n567) );
  AND2_X1 U499 ( .A1(n567), .A2(n436), .ZN(n437) );
  XOR2_X1 U500 ( .A(KEYINPUT97), .B(n437), .Z(n438) );
  NOR2_X1 U501 ( .A1(n439), .A2(n438), .ZN(n440) );
  NOR2_X1 U502 ( .A1(n544), .A2(n440), .ZN(n441) );
  NOR2_X1 U503 ( .A1(n442), .A2(n441), .ZN(n455) );
  NOR2_X1 U504 ( .A1(n582), .A2(n455), .ZN(n443) );
  NAND2_X1 U505 ( .A1(n534), .A2(n443), .ZN(n446) );
  NAND2_X1 U506 ( .A1(n478), .A2(n465), .ZN(n447) );
  NAND2_X1 U507 ( .A1(n485), .A2(n496), .ZN(n451) );
  XOR2_X1 U508 ( .A(KEYINPUT111), .B(KEYINPUT112), .Z(n449) );
  XNOR2_X1 U509 ( .A(G106GAT), .B(KEYINPUT44), .ZN(n448) );
  NOR2_X1 U510 ( .A1(n527), .A2(n574), .ZN(n466) );
  INV_X1 U511 ( .A(n562), .ZN(n537) );
  NAND2_X1 U512 ( .A1(n578), .A2(n537), .ZN(n452) );
  XNOR2_X1 U513 ( .A(n452), .B(KEYINPUT78), .ZN(n453) );
  XNOR2_X1 U514 ( .A(n453), .B(KEYINPUT16), .ZN(n454) );
  NOR2_X1 U515 ( .A1(n455), .A2(n454), .ZN(n477) );
  AND2_X1 U516 ( .A1(n466), .A2(n477), .ZN(n463) );
  NAND2_X1 U517 ( .A1(n544), .A2(n463), .ZN(n456) );
  XNOR2_X1 U518 ( .A(n456), .B(KEYINPUT34), .ZN(n457) );
  XNOR2_X1 U519 ( .A(G1GAT), .B(n457), .ZN(G1324GAT) );
  XOR2_X1 U520 ( .A(G8GAT), .B(KEYINPUT99), .Z(n459) );
  INV_X1 U521 ( .A(n539), .ZN(n492) );
  NAND2_X1 U522 ( .A1(n463), .A2(n492), .ZN(n458) );
  XNOR2_X1 U523 ( .A(n459), .B(n458), .ZN(G1325GAT) );
  XOR2_X1 U524 ( .A(KEYINPUT100), .B(KEYINPUT35), .Z(n461) );
  NAND2_X1 U525 ( .A1(n463), .A2(n495), .ZN(n460) );
  XNOR2_X1 U526 ( .A(n461), .B(n460), .ZN(n462) );
  XNOR2_X1 U527 ( .A(G15GAT), .B(n462), .ZN(G1326GAT) );
  NAND2_X1 U528 ( .A1(n463), .A2(n485), .ZN(n464) );
  XNOR2_X1 U529 ( .A(n464), .B(G22GAT), .ZN(G1327GAT) );
  XOR2_X1 U530 ( .A(G29GAT), .B(KEYINPUT39), .Z(n470) );
  XOR2_X1 U531 ( .A(KEYINPUT102), .B(KEYINPUT38), .Z(n468) );
  NAND2_X1 U532 ( .A1(n466), .A2(n465), .ZN(n467) );
  XNOR2_X1 U533 ( .A(n468), .B(n467), .ZN(n474) );
  NAND2_X1 U534 ( .A1(n474), .A2(n544), .ZN(n469) );
  XNOR2_X1 U535 ( .A(n470), .B(n469), .ZN(G1328GAT) );
  NAND2_X1 U536 ( .A1(n474), .A2(n492), .ZN(n471) );
  XNOR2_X1 U537 ( .A(n471), .B(G36GAT), .ZN(G1329GAT) );
  NAND2_X1 U538 ( .A1(n495), .A2(n474), .ZN(n472) );
  XNOR2_X1 U539 ( .A(n472), .B(KEYINPUT40), .ZN(n473) );
  XNOR2_X1 U540 ( .A(G43GAT), .B(n473), .ZN(G1330GAT) );
  XOR2_X1 U541 ( .A(G50GAT), .B(KEYINPUT103), .Z(n476) );
  NAND2_X1 U542 ( .A1(n474), .A2(n485), .ZN(n475) );
  XNOR2_X1 U543 ( .A(n476), .B(n475), .ZN(G1331GAT) );
  AND2_X1 U544 ( .A1(n478), .A2(n477), .ZN(n486) );
  NAND2_X1 U545 ( .A1(n544), .A2(n486), .ZN(n481) );
  XNOR2_X1 U546 ( .A(G57GAT), .B(KEYINPUT42), .ZN(n479) );
  XNOR2_X1 U547 ( .A(n479), .B(KEYINPUT104), .ZN(n480) );
  XNOR2_X1 U548 ( .A(n481), .B(n480), .ZN(G1332GAT) );
  XOR2_X1 U549 ( .A(G64GAT), .B(KEYINPUT105), .Z(n483) );
  NAND2_X1 U550 ( .A1(n486), .A2(n492), .ZN(n482) );
  XNOR2_X1 U551 ( .A(n483), .B(n482), .ZN(G1333GAT) );
  NAND2_X1 U552 ( .A1(n495), .A2(n486), .ZN(n484) );
  XNOR2_X1 U553 ( .A(n484), .B(G71GAT), .ZN(G1334GAT) );
  XOR2_X1 U554 ( .A(KEYINPUT43), .B(KEYINPUT107), .Z(n488) );
  NAND2_X1 U555 ( .A1(n486), .A2(n485), .ZN(n487) );
  XNOR2_X1 U556 ( .A(n488), .B(n487), .ZN(n490) );
  XOR2_X1 U557 ( .A(G78GAT), .B(KEYINPUT106), .Z(n489) );
  XNOR2_X1 U558 ( .A(n490), .B(n489), .ZN(G1335GAT) );
  NAND2_X1 U559 ( .A1(n544), .A2(n496), .ZN(n491) );
  XNOR2_X1 U560 ( .A(G85GAT), .B(n491), .ZN(G1336GAT) );
  XOR2_X1 U561 ( .A(G92GAT), .B(KEYINPUT109), .Z(n494) );
  NAND2_X1 U562 ( .A1(n492), .A2(n496), .ZN(n493) );
  XNOR2_X1 U563 ( .A(n494), .B(n493), .ZN(G1337GAT) );
  NAND2_X1 U564 ( .A1(n496), .A2(n495), .ZN(n497) );
  XNOR2_X1 U565 ( .A(n497), .B(KEYINPUT110), .ZN(n498) );
  XNOR2_X1 U566 ( .A(G99GAT), .B(n498), .ZN(G1338GAT) );
  INV_X1 U567 ( .A(KEYINPUT46), .ZN(n500) );
  NAND2_X1 U568 ( .A1(n555), .A2(n569), .ZN(n499) );
  XNOR2_X1 U569 ( .A(n500), .B(n499), .ZN(n503) );
  XOR2_X1 U570 ( .A(n578), .B(KEYINPUT113), .Z(n558) );
  INV_X1 U571 ( .A(n558), .ZN(n501) );
  NAND2_X1 U572 ( .A1(n537), .A2(n501), .ZN(n502) );
  NOR2_X1 U573 ( .A1(n503), .A2(n502), .ZN(n504) );
  XNOR2_X1 U574 ( .A(n504), .B(KEYINPUT47), .ZN(n509) );
  NOR2_X1 U575 ( .A1(n534), .A2(n582), .ZN(n505) );
  XOR2_X1 U576 ( .A(KEYINPUT45), .B(n505), .Z(n506) );
  NOR2_X1 U577 ( .A1(n574), .A2(n506), .ZN(n507) );
  NAND2_X1 U578 ( .A1(n507), .A2(n527), .ZN(n508) );
  NAND2_X1 U579 ( .A1(n509), .A2(n508), .ZN(n510) );
  XOR2_X1 U580 ( .A(KEYINPUT48), .B(n510), .Z(n540) );
  NOR2_X1 U581 ( .A1(n540), .A2(n511), .ZN(n526) );
  NAND2_X1 U582 ( .A1(n526), .A2(n512), .ZN(n513) );
  NOR2_X1 U583 ( .A1(n550), .A2(n513), .ZN(n522) );
  NAND2_X1 U584 ( .A1(n522), .A2(n569), .ZN(n514) );
  XNOR2_X1 U585 ( .A(G113GAT), .B(n514), .ZN(G1340GAT) );
  XOR2_X1 U586 ( .A(KEYINPUT115), .B(KEYINPUT49), .Z(n516) );
  NAND2_X1 U587 ( .A1(n522), .A2(n555), .ZN(n515) );
  XNOR2_X1 U588 ( .A(n516), .B(n515), .ZN(n518) );
  XOR2_X1 U589 ( .A(G120GAT), .B(KEYINPUT114), .Z(n517) );
  XNOR2_X1 U590 ( .A(n518), .B(n517), .ZN(G1341GAT) );
  XOR2_X1 U591 ( .A(KEYINPUT116), .B(KEYINPUT50), .Z(n520) );
  NAND2_X1 U592 ( .A1(n522), .A2(n558), .ZN(n519) );
  XNOR2_X1 U593 ( .A(n520), .B(n519), .ZN(n521) );
  XOR2_X1 U594 ( .A(G127GAT), .B(n521), .Z(G1342GAT) );
  XOR2_X1 U595 ( .A(KEYINPUT117), .B(KEYINPUT51), .Z(n524) );
  NAND2_X1 U596 ( .A1(n522), .A2(n562), .ZN(n523) );
  XNOR2_X1 U597 ( .A(n524), .B(n523), .ZN(n525) );
  XOR2_X1 U598 ( .A(G134GAT), .B(n525), .Z(G1343GAT) );
  NAND2_X1 U599 ( .A1(n526), .A2(n567), .ZN(n536) );
  NOR2_X1 U600 ( .A1(n527), .A2(n536), .ZN(n528) );
  XOR2_X1 U601 ( .A(G141GAT), .B(n528), .Z(n529) );
  XNOR2_X1 U602 ( .A(KEYINPUT118), .B(n529), .ZN(G1344GAT) );
  NOR2_X1 U603 ( .A1(n530), .A2(n536), .ZN(n532) );
  XNOR2_X1 U604 ( .A(KEYINPUT53), .B(KEYINPUT52), .ZN(n531) );
  XNOR2_X1 U605 ( .A(n532), .B(n531), .ZN(n533) );
  XNOR2_X1 U606 ( .A(G148GAT), .B(n533), .ZN(G1345GAT) );
  NOR2_X1 U607 ( .A1(n534), .A2(n536), .ZN(n535) );
  XOR2_X1 U608 ( .A(G155GAT), .B(n535), .Z(G1346GAT) );
  NOR2_X1 U609 ( .A1(n537), .A2(n536), .ZN(n538) );
  XOR2_X1 U610 ( .A(G162GAT), .B(n538), .Z(G1347GAT) );
  XOR2_X1 U611 ( .A(KEYINPUT119), .B(KEYINPUT54), .Z(n542) );
  XNOR2_X1 U612 ( .A(n542), .B(n541), .ZN(n543) );
  XOR2_X1 U613 ( .A(KEYINPUT64), .B(n545), .Z(n566) );
  NOR2_X1 U614 ( .A1(n546), .A2(n566), .ZN(n548) );
  XNOR2_X1 U615 ( .A(KEYINPUT55), .B(KEYINPUT120), .ZN(n547) );
  XNOR2_X1 U616 ( .A(n548), .B(n547), .ZN(n549) );
  NAND2_X1 U617 ( .A1(n563), .A2(n569), .ZN(n551) );
  XNOR2_X1 U618 ( .A(G169GAT), .B(n551), .ZN(G1348GAT) );
  XOR2_X1 U619 ( .A(KEYINPUT57), .B(KEYINPUT122), .Z(n553) );
  XNOR2_X1 U620 ( .A(G176GAT), .B(KEYINPUT56), .ZN(n552) );
  XNOR2_X1 U621 ( .A(n553), .B(n552), .ZN(n554) );
  XOR2_X1 U622 ( .A(KEYINPUT121), .B(n554), .Z(n557) );
  NAND2_X1 U623 ( .A1(n563), .A2(n555), .ZN(n556) );
  XNOR2_X1 U624 ( .A(n557), .B(n556), .ZN(G1349GAT) );
  NAND2_X1 U625 ( .A1(n558), .A2(n563), .ZN(n559) );
  XNOR2_X1 U626 ( .A(n559), .B(G183GAT), .ZN(G1350GAT) );
  XNOR2_X1 U627 ( .A(G190GAT), .B(KEYINPUT58), .ZN(n560) );
  XNOR2_X1 U628 ( .A(n560), .B(KEYINPUT123), .ZN(n561) );
  XOR2_X1 U629 ( .A(KEYINPUT124), .B(n561), .Z(n565) );
  NAND2_X1 U630 ( .A1(n563), .A2(n562), .ZN(n564) );
  XNOR2_X1 U631 ( .A(n565), .B(n564), .ZN(G1351GAT) );
  XOR2_X1 U632 ( .A(G197GAT), .B(KEYINPUT125), .Z(n571) );
  INV_X1 U633 ( .A(n566), .ZN(n568) );
  NAND2_X1 U634 ( .A1(n568), .A2(n567), .ZN(n581) );
  INV_X1 U635 ( .A(n581), .ZN(n579) );
  NAND2_X1 U636 ( .A1(n579), .A2(n569), .ZN(n570) );
  XNOR2_X1 U637 ( .A(n571), .B(n570), .ZN(n573) );
  XOR2_X1 U638 ( .A(KEYINPUT60), .B(KEYINPUT59), .Z(n572) );
  XNOR2_X1 U639 ( .A(n573), .B(n572), .ZN(G1352GAT) );
  XOR2_X1 U640 ( .A(KEYINPUT126), .B(KEYINPUT61), .Z(n576) );
  NAND2_X1 U641 ( .A1(n579), .A2(n574), .ZN(n575) );
  XNOR2_X1 U642 ( .A(n576), .B(n575), .ZN(n577) );
  XNOR2_X1 U643 ( .A(G204GAT), .B(n577), .ZN(G1353GAT) );
  NAND2_X1 U644 ( .A1(n579), .A2(n578), .ZN(n580) );
  XNOR2_X1 U645 ( .A(G211GAT), .B(n580), .ZN(G1354GAT) );
  NOR2_X1 U646 ( .A1(n582), .A2(n581), .ZN(n584) );
  XNOR2_X1 U647 ( .A(KEYINPUT62), .B(KEYINPUT127), .ZN(n583) );
  XNOR2_X1 U648 ( .A(n584), .B(n583), .ZN(n585) );
  XNOR2_X1 U649 ( .A(G218GAT), .B(n585), .ZN(G1355GAT) );
endmodule

