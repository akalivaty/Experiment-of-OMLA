//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 0 1 0 0 1 1 1 1 1 0 1 1 0 1 1 0 0 0 0 1 0 1 0 1 0 1 1 1 0 0 1 1 0 1 1 0 0 1 0 0 0 1 0 0 0 1 0 1 0 1 1 0 0 0 0 0 0 0 1 1 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:34:00 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n437, new_n444, new_n449, new_n453, new_n454, new_n455,
    new_n456, new_n457, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n519, new_n520, new_n521, new_n522, new_n523, new_n524, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n535,
    new_n536, new_n537, new_n538, new_n539, new_n540, new_n541, new_n543,
    new_n545, new_n546, new_n548, new_n549, new_n550, new_n551, new_n552,
    new_n553, new_n554, new_n555, new_n556, new_n557, new_n558, new_n559,
    new_n560, new_n561, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n573, new_n574, new_n575, new_n576, new_n577,
    new_n579, new_n580, new_n581, new_n582, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n601, new_n604,
    new_n605, new_n607, new_n608, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n814, new_n815,
    new_n816, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1101,
    new_n1102, new_n1103;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(new_n436));
  XNOR2_X1  g011(.A(new_n436), .B(KEYINPUT64), .ZN(new_n437));
  INV_X1    g012(.A(new_n437), .ZN(G220));
  XNOR2_X1  g013(.A(KEYINPUT65), .B(G96), .ZN(G221));
  INV_X1    g014(.A(G69), .ZN(G235));
  INV_X1    g015(.A(G120), .ZN(G236));
  XNOR2_X1  g016(.A(KEYINPUT66), .B(G57), .ZN(G237));
  INV_X1    g017(.A(G108), .ZN(G238));
  NAND4_X1  g018(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(new_n444));
  XNOR2_X1  g019(.A(new_n444), .B(KEYINPUT67), .ZN(G158));
  NAND3_X1  g020(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g021(.A(G452), .Z(G391));
  AND2_X1   g022(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g023(.A1(G7), .A2(G661), .ZN(new_n449));
  XOR2_X1   g024(.A(new_n449), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g025(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g026(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g027(.A1(G220), .A2(G218), .A3(G219), .A4(G221), .ZN(new_n453));
  XNOR2_X1  g028(.A(new_n453), .B(KEYINPUT2), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR4_X1   g030(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n456));
  INV_X1    g031(.A(new_n456), .ZN(new_n457));
  NOR2_X1   g032(.A1(new_n455), .A2(new_n457), .ZN(G325));
  INV_X1    g033(.A(G325), .ZN(G261));
  AOI22_X1  g034(.A1(new_n455), .A2(G2106), .B1(G567), .B2(new_n457), .ZN(G319));
  XNOR2_X1  g035(.A(KEYINPUT68), .B(G2105), .ZN(new_n461));
  XNOR2_X1  g036(.A(KEYINPUT3), .B(G2104), .ZN(new_n462));
  NAND3_X1  g037(.A1(new_n461), .A2(new_n462), .A3(G137), .ZN(new_n463));
  INV_X1    g038(.A(G101), .ZN(new_n464));
  INV_X1    g039(.A(G2104), .ZN(new_n465));
  NOR2_X1   g040(.A1(new_n465), .A2(G2105), .ZN(new_n466));
  INV_X1    g041(.A(new_n466), .ZN(new_n467));
  AOI22_X1  g042(.A1(new_n462), .A2(G125), .B1(G113), .B2(G2104), .ZN(new_n468));
  OAI221_X1 g043(.A(new_n463), .B1(new_n464), .B2(new_n467), .C1(new_n468), .C2(new_n461), .ZN(new_n469));
  INV_X1    g044(.A(new_n469), .ZN(G160));
  NAND2_X1  g045(.A1(new_n465), .A2(KEYINPUT3), .ZN(new_n471));
  INV_X1    g046(.A(KEYINPUT3), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n472), .A2(G2104), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n471), .A2(new_n473), .ZN(new_n474));
  NOR2_X1   g049(.A1(new_n474), .A2(new_n461), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n475), .A2(G124), .ZN(new_n476));
  NOR2_X1   g051(.A1(new_n474), .A2(G2105), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n477), .A2(G136), .ZN(new_n478));
  OAI221_X1 g053(.A(G2104), .B1(G100), .B2(G2105), .C1(new_n461), .C2(G112), .ZN(new_n479));
  NAND3_X1  g054(.A1(new_n476), .A2(new_n478), .A3(new_n479), .ZN(new_n480));
  INV_X1    g055(.A(new_n480), .ZN(G162));
  AND2_X1   g056(.A1(KEYINPUT68), .A2(G2105), .ZN(new_n482));
  NOR2_X1   g057(.A1(KEYINPUT68), .A2(G2105), .ZN(new_n483));
  OAI211_X1 g058(.A(new_n471), .B(new_n473), .C1(new_n482), .C2(new_n483), .ZN(new_n484));
  INV_X1    g059(.A(G138), .ZN(new_n485));
  OAI21_X1  g060(.A(KEYINPUT69), .B1(new_n484), .B2(new_n485), .ZN(new_n486));
  INV_X1    g061(.A(KEYINPUT69), .ZN(new_n487));
  NAND4_X1  g062(.A1(new_n461), .A2(new_n462), .A3(new_n487), .A4(G138), .ZN(new_n488));
  NAND3_X1  g063(.A1(new_n486), .A2(KEYINPUT4), .A3(new_n488), .ZN(new_n489));
  OR3_X1    g064(.A1(new_n484), .A2(KEYINPUT4), .A3(new_n485), .ZN(new_n490));
  NAND3_X1  g065(.A1(new_n489), .A2(KEYINPUT70), .A3(new_n490), .ZN(new_n491));
  INV_X1    g066(.A(KEYINPUT70), .ZN(new_n492));
  NAND4_X1  g067(.A1(new_n486), .A2(new_n492), .A3(KEYINPUT4), .A4(new_n488), .ZN(new_n493));
  NAND2_X1  g068(.A1(G114), .A2(G2104), .ZN(new_n494));
  INV_X1    g069(.A(G126), .ZN(new_n495));
  OAI21_X1  g070(.A(new_n494), .B1(new_n474), .B2(new_n495), .ZN(new_n496));
  AOI22_X1  g071(.A1(new_n496), .A2(G2105), .B1(G102), .B2(new_n466), .ZN(new_n497));
  NAND3_X1  g072(.A1(new_n491), .A2(new_n493), .A3(new_n497), .ZN(new_n498));
  INV_X1    g073(.A(new_n498), .ZN(G164));
  AND3_X1   g074(.A1(KEYINPUT71), .A2(KEYINPUT6), .A3(G651), .ZN(new_n500));
  AOI21_X1  g075(.A(KEYINPUT6), .B1(KEYINPUT71), .B2(G651), .ZN(new_n501));
  NOR2_X1   g076(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  INV_X1    g077(.A(G543), .ZN(new_n503));
  NOR2_X1   g078(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n504), .A2(G50), .ZN(new_n505));
  INV_X1    g080(.A(G88), .ZN(new_n506));
  OR2_X1    g081(.A1(new_n500), .A2(new_n501), .ZN(new_n507));
  NAND2_X1  g082(.A1(new_n503), .A2(KEYINPUT5), .ZN(new_n508));
  INV_X1    g083(.A(KEYINPUT5), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n509), .A2(G543), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n508), .A2(new_n510), .ZN(new_n511));
  INV_X1    g086(.A(new_n511), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n507), .A2(new_n512), .ZN(new_n513));
  OAI21_X1  g088(.A(new_n505), .B1(new_n506), .B2(new_n513), .ZN(new_n514));
  AOI22_X1  g089(.A1(new_n512), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n515));
  INV_X1    g090(.A(G651), .ZN(new_n516));
  NOR2_X1   g091(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  NOR2_X1   g092(.A1(new_n514), .A2(new_n517), .ZN(G166));
  NAND2_X1  g093(.A1(new_n504), .A2(G51), .ZN(new_n519));
  NOR2_X1   g094(.A1(new_n502), .A2(new_n511), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n520), .A2(G89), .ZN(new_n521));
  NAND3_X1  g096(.A1(new_n512), .A2(G63), .A3(G651), .ZN(new_n522));
  NAND3_X1  g097(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n523));
  XNOR2_X1  g098(.A(new_n523), .B(KEYINPUT7), .ZN(new_n524));
  NAND4_X1  g099(.A1(new_n519), .A2(new_n521), .A3(new_n522), .A4(new_n524), .ZN(G286));
  INV_X1    g100(.A(G286), .ZN(G168));
  NAND2_X1  g101(.A1(new_n520), .A2(G90), .ZN(new_n527));
  NAND2_X1  g102(.A1(new_n504), .A2(G52), .ZN(new_n528));
  AOI22_X1  g103(.A1(new_n512), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n529));
  OAI211_X1 g104(.A(new_n527), .B(new_n528), .C1(new_n529), .C2(new_n516), .ZN(new_n530));
  INV_X1    g105(.A(KEYINPUT72), .ZN(new_n531));
  OR2_X1    g106(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  NAND2_X1  g107(.A1(new_n530), .A2(new_n531), .ZN(new_n533));
  NAND2_X1  g108(.A1(new_n532), .A2(new_n533), .ZN(G171));
  NAND2_X1  g109(.A1(G68), .A2(G543), .ZN(new_n535));
  INV_X1    g110(.A(G56), .ZN(new_n536));
  OAI21_X1  g111(.A(new_n535), .B1(new_n511), .B2(new_n536), .ZN(new_n537));
  AOI22_X1  g112(.A1(G43), .A2(new_n504), .B1(new_n537), .B2(G651), .ZN(new_n538));
  NAND2_X1  g113(.A1(new_n520), .A2(G81), .ZN(new_n539));
  NAND2_X1  g114(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  INV_X1    g115(.A(new_n540), .ZN(new_n541));
  NAND2_X1  g116(.A1(new_n541), .A2(G860), .ZN(G153));
  AND3_X1   g117(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n543));
  NAND2_X1  g118(.A1(new_n543), .A2(G36), .ZN(G176));
  NAND2_X1  g119(.A1(G1), .A2(G3), .ZN(new_n545));
  XNOR2_X1  g120(.A(new_n545), .B(KEYINPUT8), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n543), .A2(new_n546), .ZN(G188));
  AND2_X1   g122(.A1(new_n520), .A2(KEYINPUT73), .ZN(new_n548));
  NOR2_X1   g123(.A1(new_n520), .A2(KEYINPUT73), .ZN(new_n549));
  OR2_X1    g124(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n550), .A2(G91), .ZN(new_n551));
  AND2_X1   g126(.A1(new_n512), .A2(G65), .ZN(new_n552));
  NAND2_X1  g127(.A1(G78), .A2(G543), .ZN(new_n553));
  XOR2_X1   g128(.A(new_n553), .B(KEYINPUT74), .Z(new_n554));
  OAI21_X1  g129(.A(G651), .B1(new_n552), .B2(new_n554), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n504), .A2(G53), .ZN(new_n556));
  XNOR2_X1  g131(.A(new_n556), .B(KEYINPUT9), .ZN(new_n557));
  NAND3_X1  g132(.A1(new_n551), .A2(new_n555), .A3(new_n557), .ZN(new_n558));
  INV_X1    g133(.A(KEYINPUT75), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  NAND4_X1  g135(.A1(new_n551), .A2(KEYINPUT75), .A3(new_n555), .A4(new_n557), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n560), .A2(new_n561), .ZN(G299));
  INV_X1    g137(.A(G171), .ZN(G301));
  INV_X1    g138(.A(G166), .ZN(G303));
  NAND3_X1  g139(.A1(new_n550), .A2(KEYINPUT76), .A3(G87), .ZN(new_n565));
  OR2_X1    g140(.A1(new_n512), .A2(G74), .ZN(new_n566));
  AOI22_X1  g141(.A1(new_n566), .A2(G651), .B1(G49), .B2(new_n504), .ZN(new_n567));
  INV_X1    g142(.A(KEYINPUT76), .ZN(new_n568));
  NOR2_X1   g143(.A1(new_n548), .A2(new_n549), .ZN(new_n569));
  INV_X1    g144(.A(G87), .ZN(new_n570));
  OAI21_X1  g145(.A(new_n568), .B1(new_n569), .B2(new_n570), .ZN(new_n571));
  NAND3_X1  g146(.A1(new_n565), .A2(new_n567), .A3(new_n571), .ZN(G288));
  NAND2_X1  g147(.A1(G73), .A2(G543), .ZN(new_n573));
  INV_X1    g148(.A(G61), .ZN(new_n574));
  OAI21_X1  g149(.A(new_n573), .B1(new_n511), .B2(new_n574), .ZN(new_n575));
  AOI22_X1  g150(.A1(G48), .A2(new_n504), .B1(new_n575), .B2(G651), .ZN(new_n576));
  INV_X1    g151(.A(G86), .ZN(new_n577));
  OAI21_X1  g152(.A(new_n576), .B1(new_n569), .B2(new_n577), .ZN(G305));
  NAND2_X1  g153(.A1(new_n520), .A2(G85), .ZN(new_n579));
  INV_X1    g154(.A(new_n504), .ZN(new_n580));
  XOR2_X1   g155(.A(KEYINPUT77), .B(G47), .Z(new_n581));
  AOI22_X1  g156(.A1(new_n512), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n582));
  OAI221_X1 g157(.A(new_n579), .B1(new_n580), .B2(new_n581), .C1(new_n516), .C2(new_n582), .ZN(G290));
  INV_X1    g158(.A(G868), .ZN(new_n584));
  NOR2_X1   g159(.A1(G171), .A2(new_n584), .ZN(new_n585));
  INV_X1    g160(.A(KEYINPUT78), .ZN(new_n586));
  NAND2_X1  g161(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  INV_X1    g162(.A(G92), .ZN(new_n588));
  OR3_X1    g163(.A1(new_n569), .A2(KEYINPUT10), .A3(new_n588), .ZN(new_n589));
  NAND2_X1  g164(.A1(G79), .A2(G543), .ZN(new_n590));
  XNOR2_X1  g165(.A(new_n590), .B(KEYINPUT79), .ZN(new_n591));
  INV_X1    g166(.A(G66), .ZN(new_n592));
  OAI21_X1  g167(.A(new_n591), .B1(new_n592), .B2(new_n511), .ZN(new_n593));
  AOI22_X1  g168(.A1(new_n593), .A2(G651), .B1(G54), .B2(new_n504), .ZN(new_n594));
  OAI21_X1  g169(.A(KEYINPUT10), .B1(new_n569), .B2(new_n588), .ZN(new_n595));
  NAND3_X1  g170(.A1(new_n589), .A2(new_n594), .A3(new_n595), .ZN(new_n596));
  XNOR2_X1  g171(.A(new_n596), .B(KEYINPUT80), .ZN(new_n597));
  AOI21_X1  g172(.A(KEYINPUT78), .B1(new_n597), .B2(new_n584), .ZN(new_n598));
  OAI21_X1  g173(.A(new_n587), .B1(new_n598), .B2(new_n585), .ZN(G284));
  OAI21_X1  g174(.A(new_n587), .B1(new_n598), .B2(new_n585), .ZN(G321));
  NAND2_X1  g175(.A1(G299), .A2(new_n584), .ZN(new_n601));
  OAI21_X1  g176(.A(new_n601), .B1(new_n584), .B2(G168), .ZN(G297));
  OAI21_X1  g177(.A(new_n601), .B1(new_n584), .B2(G168), .ZN(G280));
  INV_X1    g178(.A(new_n597), .ZN(new_n604));
  INV_X1    g179(.A(G559), .ZN(new_n605));
  OAI21_X1  g180(.A(new_n604), .B1(new_n605), .B2(G860), .ZN(G148));
  NAND2_X1  g181(.A1(new_n540), .A2(new_n584), .ZN(new_n607));
  NOR2_X1   g182(.A1(new_n597), .A2(G559), .ZN(new_n608));
  OAI21_X1  g183(.A(new_n607), .B1(new_n608), .B2(new_n584), .ZN(G323));
  XNOR2_X1  g184(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NOR2_X1   g185(.A1(new_n461), .A2(G111), .ZN(new_n611));
  XNOR2_X1  g186(.A(new_n611), .B(KEYINPUT84), .ZN(new_n612));
  OAI211_X1 g187(.A(new_n612), .B(G2104), .C1(G99), .C2(G2105), .ZN(new_n613));
  NAND2_X1  g188(.A1(new_n477), .A2(G135), .ZN(new_n614));
  NAND2_X1  g189(.A1(new_n475), .A2(G123), .ZN(new_n615));
  NAND3_X1  g190(.A1(new_n613), .A2(new_n614), .A3(new_n615), .ZN(new_n616));
  INV_X1    g191(.A(new_n616), .ZN(new_n617));
  INV_X1    g192(.A(G2096), .ZN(new_n618));
  AOI22_X1  g193(.A1(new_n617), .A2(new_n618), .B1(KEYINPUT83), .B2(G2100), .ZN(new_n619));
  NAND2_X1  g194(.A1(new_n462), .A2(new_n466), .ZN(new_n620));
  XNOR2_X1  g195(.A(KEYINPUT81), .B(KEYINPUT12), .ZN(new_n621));
  XNOR2_X1  g196(.A(new_n620), .B(new_n621), .ZN(new_n622));
  NOR2_X1   g197(.A1(KEYINPUT83), .A2(G2100), .ZN(new_n623));
  XNOR2_X1  g198(.A(new_n622), .B(new_n623), .ZN(new_n624));
  XOR2_X1   g199(.A(KEYINPUT82), .B(KEYINPUT13), .Z(new_n625));
  XNOR2_X1  g200(.A(new_n624), .B(new_n625), .ZN(new_n626));
  OAI211_X1 g201(.A(new_n619), .B(new_n626), .C1(new_n618), .C2(new_n617), .ZN(G156));
  INV_X1    g202(.A(KEYINPUT85), .ZN(new_n628));
  XNOR2_X1  g203(.A(G2427), .B(G2438), .ZN(new_n629));
  XNOR2_X1  g204(.A(new_n629), .B(G2430), .ZN(new_n630));
  XNOR2_X1  g205(.A(new_n630), .B(KEYINPUT15), .ZN(new_n631));
  INV_X1    g206(.A(G2435), .ZN(new_n632));
  XNOR2_X1  g207(.A(new_n631), .B(new_n632), .ZN(new_n633));
  NAND2_X1  g208(.A1(new_n633), .A2(KEYINPUT14), .ZN(new_n634));
  XNOR2_X1  g209(.A(G2451), .B(G2454), .ZN(new_n635));
  XNOR2_X1  g210(.A(new_n635), .B(KEYINPUT16), .ZN(new_n636));
  NAND2_X1  g211(.A1(new_n634), .A2(new_n636), .ZN(new_n637));
  INV_X1    g212(.A(new_n636), .ZN(new_n638));
  NAND3_X1  g213(.A1(new_n633), .A2(KEYINPUT14), .A3(new_n638), .ZN(new_n639));
  NAND2_X1  g214(.A1(new_n637), .A2(new_n639), .ZN(new_n640));
  XNOR2_X1  g215(.A(G2443), .B(G2446), .ZN(new_n641));
  INV_X1    g216(.A(new_n641), .ZN(new_n642));
  NAND2_X1  g217(.A1(new_n640), .A2(new_n642), .ZN(new_n643));
  NAND3_X1  g218(.A1(new_n637), .A2(new_n641), .A3(new_n639), .ZN(new_n644));
  NAND2_X1  g219(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  XOR2_X1   g220(.A(G1341), .B(G1348), .Z(new_n646));
  OAI21_X1  g221(.A(new_n628), .B1(new_n645), .B2(new_n646), .ZN(new_n647));
  INV_X1    g222(.A(G14), .ZN(new_n648));
  AOI21_X1  g223(.A(new_n648), .B1(new_n645), .B2(new_n646), .ZN(new_n649));
  INV_X1    g224(.A(new_n646), .ZN(new_n650));
  NAND4_X1  g225(.A1(new_n643), .A2(KEYINPUT85), .A3(new_n650), .A4(new_n644), .ZN(new_n651));
  NAND3_X1  g226(.A1(new_n647), .A2(new_n649), .A3(new_n651), .ZN(new_n652));
  INV_X1    g227(.A(new_n652), .ZN(G401));
  XOR2_X1   g228(.A(G2067), .B(G2678), .Z(new_n654));
  INV_X1    g229(.A(new_n654), .ZN(new_n655));
  XNOR2_X1  g230(.A(G2072), .B(G2078), .ZN(new_n656));
  XOR2_X1   g231(.A(G2084), .B(G2090), .Z(new_n657));
  NAND3_X1  g232(.A1(new_n655), .A2(new_n656), .A3(new_n657), .ZN(new_n658));
  XOR2_X1   g233(.A(new_n658), .B(KEYINPUT18), .Z(new_n659));
  XNOR2_X1  g234(.A(new_n656), .B(KEYINPUT86), .ZN(new_n660));
  AOI21_X1  g235(.A(new_n657), .B1(new_n660), .B2(new_n654), .ZN(new_n661));
  XOR2_X1   g236(.A(new_n656), .B(KEYINPUT17), .Z(new_n662));
  OAI21_X1  g237(.A(new_n661), .B1(new_n654), .B2(new_n662), .ZN(new_n663));
  NAND3_X1  g238(.A1(new_n662), .A2(new_n654), .A3(new_n657), .ZN(new_n664));
  NAND3_X1  g239(.A1(new_n659), .A2(new_n663), .A3(new_n664), .ZN(new_n665));
  XNOR2_X1  g240(.A(new_n665), .B(KEYINPUT87), .ZN(new_n666));
  XNOR2_X1  g241(.A(G2096), .B(G2100), .ZN(new_n667));
  XNOR2_X1  g242(.A(new_n666), .B(new_n667), .ZN(new_n668));
  INV_X1    g243(.A(new_n668), .ZN(G227));
  XNOR2_X1  g244(.A(G1961), .B(G1966), .ZN(new_n670));
  XNOR2_X1  g245(.A(new_n670), .B(KEYINPUT88), .ZN(new_n671));
  XOR2_X1   g246(.A(G1956), .B(G2474), .Z(new_n672));
  AND2_X1   g247(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  XOR2_X1   g248(.A(G1971), .B(G1976), .Z(new_n674));
  XNOR2_X1  g249(.A(new_n674), .B(KEYINPUT19), .ZN(new_n675));
  NAND2_X1  g250(.A1(new_n673), .A2(new_n675), .ZN(new_n676));
  INV_X1    g251(.A(KEYINPUT20), .ZN(new_n677));
  NOR2_X1   g252(.A1(new_n671), .A2(new_n672), .ZN(new_n678));
  AOI22_X1  g253(.A1(new_n676), .A2(new_n677), .B1(new_n675), .B2(new_n678), .ZN(new_n679));
  OR3_X1    g254(.A1(new_n673), .A2(new_n678), .A3(new_n675), .ZN(new_n680));
  OAI211_X1 g255(.A(new_n679), .B(new_n680), .C1(new_n677), .C2(new_n676), .ZN(new_n681));
  XNOR2_X1  g256(.A(new_n681), .B(KEYINPUT89), .ZN(new_n682));
  XOR2_X1   g257(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n683));
  XNOR2_X1  g258(.A(G1981), .B(G1986), .ZN(new_n684));
  XNOR2_X1  g259(.A(new_n683), .B(new_n684), .ZN(new_n685));
  XNOR2_X1  g260(.A(new_n682), .B(new_n685), .ZN(new_n686));
  XOR2_X1   g261(.A(G1991), .B(G1996), .Z(new_n687));
  XNOR2_X1  g262(.A(new_n686), .B(new_n687), .ZN(G229));
  INV_X1    g263(.A(KEYINPUT93), .ZN(new_n689));
  NOR2_X1   g264(.A1(new_n689), .A2(KEYINPUT36), .ZN(new_n690));
  INV_X1    g265(.A(new_n690), .ZN(new_n691));
  AOI22_X1  g266(.A1(G119), .A2(new_n475), .B1(new_n477), .B2(G131), .ZN(new_n692));
  NOR2_X1   g267(.A1(new_n461), .A2(G107), .ZN(new_n693));
  OAI21_X1  g268(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n694));
  OAI21_X1  g269(.A(new_n692), .B1(new_n693), .B2(new_n694), .ZN(new_n695));
  NAND2_X1  g270(.A1(new_n695), .A2(G29), .ZN(new_n696));
  INV_X1    g271(.A(G25), .ZN(new_n697));
  OAI21_X1  g272(.A(KEYINPUT90), .B1(new_n697), .B2(G29), .ZN(new_n698));
  OR3_X1    g273(.A1(new_n697), .A2(KEYINPUT90), .A3(G29), .ZN(new_n699));
  NAND3_X1  g274(.A1(new_n696), .A2(new_n698), .A3(new_n699), .ZN(new_n700));
  XNOR2_X1  g275(.A(KEYINPUT35), .B(G1991), .ZN(new_n701));
  XNOR2_X1  g276(.A(new_n700), .B(new_n701), .ZN(new_n702));
  MUX2_X1   g277(.A(G6), .B(G305), .S(G16), .Z(new_n703));
  XNOR2_X1  g278(.A(new_n703), .B(KEYINPUT92), .ZN(new_n704));
  XOR2_X1   g279(.A(KEYINPUT32), .B(G1981), .Z(new_n705));
  XNOR2_X1  g280(.A(new_n704), .B(new_n705), .ZN(new_n706));
  XNOR2_X1  g281(.A(KEYINPUT91), .B(G16), .ZN(new_n707));
  MUX2_X1   g282(.A(G22), .B(G303), .S(new_n707), .Z(new_n708));
  INV_X1    g283(.A(G1971), .ZN(new_n709));
  XNOR2_X1  g284(.A(new_n708), .B(new_n709), .ZN(new_n710));
  NOR2_X1   g285(.A1(G16), .A2(G23), .ZN(new_n711));
  INV_X1    g286(.A(G288), .ZN(new_n712));
  AOI21_X1  g287(.A(new_n711), .B1(new_n712), .B2(G16), .ZN(new_n713));
  XNOR2_X1  g288(.A(KEYINPUT33), .B(G1976), .ZN(new_n714));
  XNOR2_X1  g289(.A(new_n713), .B(new_n714), .ZN(new_n715));
  NAND3_X1  g290(.A1(new_n706), .A2(new_n710), .A3(new_n715), .ZN(new_n716));
  INV_X1    g291(.A(KEYINPUT34), .ZN(new_n717));
  OR2_X1    g292(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  NAND2_X1  g293(.A1(new_n716), .A2(new_n717), .ZN(new_n719));
  AOI21_X1  g294(.A(new_n702), .B1(new_n718), .B2(new_n719), .ZN(new_n720));
  MUX2_X1   g295(.A(G24), .B(G290), .S(new_n707), .Z(new_n721));
  XOR2_X1   g296(.A(new_n721), .B(G1986), .Z(new_n722));
  AOI21_X1  g297(.A(new_n691), .B1(new_n720), .B2(new_n722), .ZN(new_n723));
  INV_X1    g298(.A(new_n723), .ZN(new_n724));
  NAND3_X1  g299(.A1(new_n720), .A2(new_n691), .A3(new_n722), .ZN(new_n725));
  NAND2_X1  g300(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  NAND2_X1  g301(.A1(new_n689), .A2(KEYINPUT36), .ZN(new_n727));
  AOI22_X1  g302(.A1(G129), .A2(new_n475), .B1(new_n477), .B2(G141), .ZN(new_n728));
  NAND2_X1  g303(.A1(new_n466), .A2(G105), .ZN(new_n729));
  NAND3_X1  g304(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n730));
  XOR2_X1   g305(.A(new_n730), .B(KEYINPUT26), .Z(new_n731));
  NAND3_X1  g306(.A1(new_n728), .A2(new_n729), .A3(new_n731), .ZN(new_n732));
  XOR2_X1   g307(.A(new_n732), .B(KEYINPUT97), .Z(new_n733));
  NAND2_X1  g308(.A1(new_n733), .A2(G29), .ZN(new_n734));
  OAI21_X1  g309(.A(new_n734), .B1(G29), .B2(G32), .ZN(new_n735));
  XOR2_X1   g310(.A(KEYINPUT27), .B(G1996), .Z(new_n736));
  INV_X1    g311(.A(new_n736), .ZN(new_n737));
  INV_X1    g312(.A(G29), .ZN(new_n738));
  NAND2_X1  g313(.A1(new_n738), .A2(G33), .ZN(new_n739));
  NAND3_X1  g314(.A1(new_n461), .A2(G103), .A3(G2104), .ZN(new_n740));
  XOR2_X1   g315(.A(new_n740), .B(KEYINPUT25), .Z(new_n741));
  NAND2_X1  g316(.A1(new_n477), .A2(G139), .ZN(new_n742));
  AOI22_X1  g317(.A1(new_n462), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n743));
  OAI211_X1 g318(.A(new_n741), .B(new_n742), .C1(new_n461), .C2(new_n743), .ZN(new_n744));
  INV_X1    g319(.A(new_n744), .ZN(new_n745));
  OAI21_X1  g320(.A(new_n739), .B1(new_n745), .B2(new_n738), .ZN(new_n746));
  AOI22_X1  g321(.A1(new_n735), .A2(new_n737), .B1(G2072), .B2(new_n746), .ZN(new_n747));
  INV_X1    g322(.A(KEYINPUT24), .ZN(new_n748));
  OAI21_X1  g323(.A(new_n738), .B1(new_n748), .B2(G34), .ZN(new_n749));
  INV_X1    g324(.A(KEYINPUT94), .ZN(new_n750));
  OR2_X1    g325(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  NAND2_X1  g326(.A1(new_n748), .A2(G34), .ZN(new_n752));
  NAND2_X1  g327(.A1(new_n749), .A2(new_n750), .ZN(new_n753));
  NAND3_X1  g328(.A1(new_n751), .A2(new_n752), .A3(new_n753), .ZN(new_n754));
  OR2_X1    g329(.A1(new_n754), .A2(KEYINPUT95), .ZN(new_n755));
  NAND2_X1  g330(.A1(new_n754), .A2(KEYINPUT95), .ZN(new_n756));
  OAI211_X1 g331(.A(new_n755), .B(new_n756), .C1(new_n469), .C2(new_n738), .ZN(new_n757));
  INV_X1    g332(.A(G2084), .ZN(new_n758));
  NOR2_X1   g333(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  XOR2_X1   g334(.A(new_n759), .B(KEYINPUT96), .Z(new_n760));
  OAI211_X1 g335(.A(new_n747), .B(new_n760), .C1(G2072), .C2(new_n746), .ZN(new_n761));
  XNOR2_X1  g336(.A(new_n761), .B(KEYINPUT98), .ZN(new_n762));
  INV_X1    g337(.A(G20), .ZN(new_n763));
  NOR2_X1   g338(.A1(new_n707), .A2(new_n763), .ZN(new_n764));
  XNOR2_X1  g339(.A(new_n764), .B(KEYINPUT100), .ZN(new_n765));
  XNOR2_X1  g340(.A(new_n765), .B(KEYINPUT23), .ZN(new_n766));
  AOI21_X1  g341(.A(new_n766), .B1(G299), .B2(G16), .ZN(new_n767));
  XNOR2_X1  g342(.A(new_n767), .B(KEYINPUT101), .ZN(new_n768));
  INV_X1    g343(.A(G1956), .ZN(new_n769));
  XNOR2_X1  g344(.A(new_n768), .B(new_n769), .ZN(new_n770));
  MUX2_X1   g345(.A(G4), .B(new_n597), .S(G16), .Z(new_n771));
  INV_X1    g346(.A(G1348), .ZN(new_n772));
  XNOR2_X1  g347(.A(new_n771), .B(new_n772), .ZN(new_n773));
  XOR2_X1   g348(.A(KEYINPUT31), .B(G11), .Z(new_n774));
  INV_X1    g349(.A(new_n735), .ZN(new_n775));
  AOI21_X1  g350(.A(new_n774), .B1(new_n775), .B2(new_n736), .ZN(new_n776));
  NAND4_X1  g351(.A1(new_n762), .A2(new_n770), .A3(new_n773), .A4(new_n776), .ZN(new_n777));
  NOR2_X1   g352(.A1(G5), .A2(G16), .ZN(new_n778));
  AOI21_X1  g353(.A(new_n778), .B1(G171), .B2(G16), .ZN(new_n779));
  XNOR2_X1  g354(.A(new_n779), .B(G1961), .ZN(new_n780));
  NAND2_X1  g355(.A1(new_n738), .A2(G35), .ZN(new_n781));
  OAI21_X1  g356(.A(new_n781), .B1(G162), .B2(new_n738), .ZN(new_n782));
  XOR2_X1   g357(.A(new_n782), .B(KEYINPUT99), .Z(new_n783));
  XOR2_X1   g358(.A(KEYINPUT29), .B(G2090), .Z(new_n784));
  NAND2_X1  g359(.A1(new_n738), .A2(G26), .ZN(new_n785));
  NAND2_X1  g360(.A1(new_n475), .A2(G128), .ZN(new_n786));
  NAND2_X1  g361(.A1(new_n477), .A2(G140), .ZN(new_n787));
  OAI221_X1 g362(.A(G2104), .B1(G104), .B2(G2105), .C1(new_n461), .C2(G116), .ZN(new_n788));
  NAND3_X1  g363(.A1(new_n786), .A2(new_n787), .A3(new_n788), .ZN(new_n789));
  INV_X1    g364(.A(new_n789), .ZN(new_n790));
  OAI21_X1  g365(.A(new_n785), .B1(new_n790), .B2(new_n738), .ZN(new_n791));
  MUX2_X1   g366(.A(new_n785), .B(new_n791), .S(KEYINPUT28), .Z(new_n792));
  AOI22_X1  g367(.A1(new_n783), .A2(new_n784), .B1(G2067), .B2(new_n792), .ZN(new_n793));
  OAI21_X1  g368(.A(new_n793), .B1(G2067), .B2(new_n792), .ZN(new_n794));
  MUX2_X1   g369(.A(G19), .B(new_n540), .S(new_n707), .Z(new_n795));
  XOR2_X1   g370(.A(new_n795), .B(G1341), .Z(new_n796));
  XNOR2_X1  g371(.A(KEYINPUT30), .B(G28), .ZN(new_n797));
  AOI22_X1  g372(.A1(new_n757), .A2(new_n758), .B1(new_n738), .B2(new_n797), .ZN(new_n798));
  OAI211_X1 g373(.A(new_n796), .B(new_n798), .C1(new_n784), .C2(new_n783), .ZN(new_n799));
  NOR2_X1   g374(.A1(new_n794), .A2(new_n799), .ZN(new_n800));
  MUX2_X1   g375(.A(G21), .B(G286), .S(G16), .Z(new_n801));
  INV_X1    g376(.A(G1966), .ZN(new_n802));
  XNOR2_X1  g377(.A(new_n801), .B(new_n802), .ZN(new_n803));
  NAND2_X1  g378(.A1(new_n738), .A2(G27), .ZN(new_n804));
  OAI21_X1  g379(.A(new_n804), .B1(G164), .B2(new_n738), .ZN(new_n805));
  OR2_X1    g380(.A1(new_n805), .A2(G2078), .ZN(new_n806));
  AOI22_X1  g381(.A1(new_n805), .A2(G2078), .B1(G29), .B2(new_n617), .ZN(new_n807));
  NAND4_X1  g382(.A1(new_n800), .A2(new_n803), .A3(new_n806), .A4(new_n807), .ZN(new_n808));
  NOR3_X1   g383(.A1(new_n777), .A2(new_n780), .A3(new_n808), .ZN(new_n809));
  INV_X1    g384(.A(KEYINPUT102), .ZN(new_n810));
  OR2_X1    g385(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  NAND2_X1  g386(.A1(new_n809), .A2(new_n810), .ZN(new_n812));
  AOI22_X1  g387(.A1(new_n726), .A2(new_n727), .B1(new_n811), .B2(new_n812), .ZN(G311));
  NAND2_X1  g388(.A1(new_n811), .A2(new_n812), .ZN(new_n814));
  INV_X1    g389(.A(new_n725), .ZN(new_n815));
  OAI21_X1  g390(.A(new_n727), .B1(new_n815), .B2(new_n723), .ZN(new_n816));
  NAND2_X1  g391(.A1(new_n814), .A2(new_n816), .ZN(G150));
  NAND2_X1  g392(.A1(new_n520), .A2(G93), .ZN(new_n818));
  NAND2_X1  g393(.A1(new_n504), .A2(G55), .ZN(new_n819));
  AOI22_X1  g394(.A1(new_n512), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n820));
  OAI211_X1 g395(.A(new_n818), .B(new_n819), .C1(new_n820), .C2(new_n516), .ZN(new_n821));
  NAND2_X1  g396(.A1(new_n821), .A2(G860), .ZN(new_n822));
  XOR2_X1   g397(.A(new_n822), .B(KEYINPUT37), .Z(new_n823));
  NAND2_X1  g398(.A1(new_n604), .A2(G559), .ZN(new_n824));
  XNOR2_X1  g399(.A(new_n824), .B(KEYINPUT38), .ZN(new_n825));
  XNOR2_X1  g400(.A(new_n540), .B(new_n821), .ZN(new_n826));
  XOR2_X1   g401(.A(new_n826), .B(KEYINPUT39), .Z(new_n827));
  XNOR2_X1  g402(.A(new_n825), .B(new_n827), .ZN(new_n828));
  OAI21_X1  g403(.A(new_n823), .B1(new_n828), .B2(G860), .ZN(G145));
  XNOR2_X1  g404(.A(new_n480), .B(KEYINPUT103), .ZN(new_n830));
  XNOR2_X1  g405(.A(new_n830), .B(G160), .ZN(new_n831));
  XNOR2_X1  g406(.A(new_n831), .B(new_n616), .ZN(new_n832));
  XNOR2_X1  g407(.A(new_n733), .B(new_n790), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n833), .A2(G164), .ZN(new_n834));
  XNOR2_X1  g409(.A(new_n733), .B(new_n789), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n835), .A2(new_n498), .ZN(new_n836));
  NAND2_X1  g411(.A1(new_n834), .A2(new_n836), .ZN(new_n837));
  INV_X1    g412(.A(KEYINPUT104), .ZN(new_n838));
  AOI21_X1  g413(.A(KEYINPUT105), .B1(new_n745), .B2(new_n838), .ZN(new_n839));
  NAND2_X1  g414(.A1(new_n837), .A2(new_n839), .ZN(new_n840));
  XOR2_X1   g415(.A(new_n695), .B(KEYINPUT106), .Z(new_n841));
  AOI22_X1  g416(.A1(G130), .A2(new_n475), .B1(new_n477), .B2(G142), .ZN(new_n842));
  OAI221_X1 g417(.A(G2104), .B1(G106), .B2(G2105), .C1(new_n461), .C2(G118), .ZN(new_n843));
  NAND2_X1  g418(.A1(new_n842), .A2(new_n843), .ZN(new_n844));
  XNOR2_X1  g419(.A(new_n841), .B(new_n844), .ZN(new_n845));
  XNOR2_X1  g420(.A(new_n845), .B(new_n622), .ZN(new_n846));
  NAND2_X1  g421(.A1(new_n745), .A2(KEYINPUT105), .ZN(new_n847));
  INV_X1    g422(.A(new_n839), .ZN(new_n848));
  NAND4_X1  g423(.A1(new_n834), .A2(new_n836), .A3(new_n847), .A4(new_n848), .ZN(new_n849));
  AND3_X1   g424(.A1(new_n840), .A2(new_n846), .A3(new_n849), .ZN(new_n850));
  AOI21_X1  g425(.A(new_n846), .B1(new_n840), .B2(new_n849), .ZN(new_n851));
  OAI21_X1  g426(.A(new_n832), .B1(new_n850), .B2(new_n851), .ZN(new_n852));
  INV_X1    g427(.A(KEYINPUT107), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  OR3_X1    g429(.A1(new_n850), .A2(new_n851), .A3(new_n832), .ZN(new_n855));
  INV_X1    g430(.A(G37), .ZN(new_n856));
  OAI211_X1 g431(.A(KEYINPUT107), .B(new_n832), .C1(new_n850), .C2(new_n851), .ZN(new_n857));
  NAND4_X1  g432(.A1(new_n854), .A2(new_n855), .A3(new_n856), .A4(new_n857), .ZN(new_n858));
  XNOR2_X1  g433(.A(new_n858), .B(KEYINPUT40), .ZN(G395));
  INV_X1    g434(.A(new_n826), .ZN(new_n860));
  XNOR2_X1  g435(.A(new_n608), .B(new_n860), .ZN(new_n861));
  INV_X1    g436(.A(KEYINPUT108), .ZN(new_n862));
  NAND2_X1  g437(.A1(G299), .A2(new_n862), .ZN(new_n863));
  INV_X1    g438(.A(new_n596), .ZN(new_n864));
  NAND3_X1  g439(.A1(new_n560), .A2(KEYINPUT108), .A3(new_n561), .ZN(new_n865));
  NAND3_X1  g440(.A1(new_n863), .A2(new_n864), .A3(new_n865), .ZN(new_n866));
  NAND3_X1  g441(.A1(G299), .A2(new_n862), .A3(new_n596), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  NAND2_X1  g443(.A1(new_n861), .A2(new_n868), .ZN(new_n869));
  AND3_X1   g444(.A1(new_n866), .A2(KEYINPUT41), .A3(new_n867), .ZN(new_n870));
  AOI21_X1  g445(.A(KEYINPUT41), .B1(new_n866), .B2(new_n867), .ZN(new_n871));
  NOR2_X1   g446(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  OAI21_X1  g447(.A(new_n869), .B1(new_n861), .B2(new_n872), .ZN(new_n873));
  OR2_X1    g448(.A1(new_n873), .A2(KEYINPUT42), .ZN(new_n874));
  XNOR2_X1  g449(.A(G288), .B(G290), .ZN(new_n875));
  XNOR2_X1  g450(.A(G303), .B(G305), .ZN(new_n876));
  XOR2_X1   g451(.A(new_n875), .B(new_n876), .Z(new_n877));
  INV_X1    g452(.A(new_n877), .ZN(new_n878));
  NOR2_X1   g453(.A1(new_n878), .A2(KEYINPUT109), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n873), .A2(KEYINPUT42), .ZN(new_n880));
  AND3_X1   g455(.A1(new_n874), .A2(new_n879), .A3(new_n880), .ZN(new_n881));
  AOI21_X1  g456(.A(new_n879), .B1(new_n874), .B2(new_n880), .ZN(new_n882));
  OAI21_X1  g457(.A(G868), .B1(new_n881), .B2(new_n882), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n821), .A2(new_n584), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n883), .A2(new_n884), .ZN(G295));
  NAND2_X1  g460(.A1(new_n883), .A2(new_n884), .ZN(G331));
  XNOR2_X1  g461(.A(G171), .B(G286), .ZN(new_n887));
  XNOR2_X1  g462(.A(new_n887), .B(new_n826), .ZN(new_n888));
  INV_X1    g463(.A(KEYINPUT41), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n868), .A2(new_n889), .ZN(new_n890));
  NAND3_X1  g465(.A1(new_n866), .A2(KEYINPUT41), .A3(new_n867), .ZN(new_n891));
  AOI21_X1  g466(.A(new_n888), .B1(new_n890), .B2(new_n891), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n868), .A2(new_n888), .ZN(new_n893));
  INV_X1    g468(.A(new_n893), .ZN(new_n894));
  OAI21_X1  g469(.A(new_n878), .B1(new_n892), .B2(new_n894), .ZN(new_n895));
  OAI211_X1 g470(.A(new_n877), .B(new_n893), .C1(new_n872), .C2(new_n888), .ZN(new_n896));
  NAND3_X1  g471(.A1(new_n895), .A2(new_n896), .A3(new_n856), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n897), .A2(KEYINPUT43), .ZN(new_n898));
  INV_X1    g473(.A(KEYINPUT43), .ZN(new_n899));
  NAND4_X1  g474(.A1(new_n895), .A2(new_n896), .A3(new_n899), .A4(new_n856), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n898), .A2(new_n900), .ZN(new_n901));
  XOR2_X1   g476(.A(new_n901), .B(KEYINPUT44), .Z(G397));
  INV_X1    g477(.A(G1384), .ZN(new_n903));
  AND3_X1   g478(.A1(new_n489), .A2(KEYINPUT70), .A3(new_n490), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n493), .A2(new_n497), .ZN(new_n905));
  OAI21_X1  g480(.A(new_n903), .B1(new_n904), .B2(new_n905), .ZN(new_n906));
  INV_X1    g481(.A(KEYINPUT45), .ZN(new_n907));
  AND2_X1   g482(.A1(G160), .A2(G40), .ZN(new_n908));
  NAND3_X1  g483(.A1(new_n906), .A2(new_n907), .A3(new_n908), .ZN(new_n909));
  XNOR2_X1  g484(.A(new_n909), .B(KEYINPUT110), .ZN(new_n910));
  INV_X1    g485(.A(new_n910), .ZN(new_n911));
  NOR2_X1   g486(.A1(new_n909), .A2(G1996), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n912), .A2(new_n733), .ZN(new_n913));
  INV_X1    g488(.A(G2067), .ZN(new_n914));
  XNOR2_X1  g489(.A(new_n789), .B(new_n914), .ZN(new_n915));
  INV_X1    g490(.A(new_n915), .ZN(new_n916));
  INV_X1    g491(.A(new_n733), .ZN(new_n917));
  AOI21_X1  g492(.A(new_n916), .B1(new_n917), .B2(G1996), .ZN(new_n918));
  OAI21_X1  g493(.A(new_n913), .B1(new_n911), .B2(new_n918), .ZN(new_n919));
  OR3_X1    g494(.A1(new_n919), .A2(new_n701), .A3(new_n695), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n790), .A2(new_n914), .ZN(new_n921));
  AOI21_X1  g496(.A(new_n911), .B1(new_n920), .B2(new_n921), .ZN(new_n922));
  XOR2_X1   g497(.A(new_n912), .B(KEYINPUT46), .Z(new_n923));
  OAI21_X1  g498(.A(new_n910), .B1(new_n917), .B2(new_n916), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  XOR2_X1   g500(.A(new_n925), .B(KEYINPUT47), .Z(new_n926));
  XNOR2_X1  g501(.A(new_n695), .B(new_n701), .ZN(new_n927));
  AOI21_X1  g502(.A(new_n919), .B1(new_n927), .B2(new_n910), .ZN(new_n928));
  NOR3_X1   g503(.A1(new_n909), .A2(G1986), .A3(G290), .ZN(new_n929));
  XOR2_X1   g504(.A(new_n929), .B(KEYINPUT48), .Z(new_n930));
  AOI211_X1 g505(.A(new_n922), .B(new_n926), .C1(new_n928), .C2(new_n930), .ZN(new_n931));
  INV_X1    g506(.A(G8), .ZN(new_n932));
  AND2_X1   g507(.A1(new_n493), .A2(new_n497), .ZN(new_n933));
  AOI21_X1  g508(.A(G1384), .B1(new_n933), .B2(new_n491), .ZN(new_n934));
  AOI21_X1  g509(.A(new_n932), .B1(new_n934), .B2(new_n908), .ZN(new_n935));
  OR2_X1    g510(.A1(G305), .A2(G1981), .ZN(new_n936));
  XOR2_X1   g511(.A(KEYINPUT113), .B(G86), .Z(new_n937));
  OAI21_X1  g512(.A(new_n576), .B1(new_n513), .B2(new_n937), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n938), .A2(G1981), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n936), .A2(new_n939), .ZN(new_n940));
  INV_X1    g515(.A(KEYINPUT49), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  NAND3_X1  g517(.A1(new_n936), .A2(KEYINPUT49), .A3(new_n939), .ZN(new_n943));
  NAND3_X1  g518(.A1(new_n942), .A2(new_n943), .A3(new_n935), .ZN(new_n944));
  INV_X1    g519(.A(G1976), .ZN(new_n945));
  AND3_X1   g520(.A1(new_n944), .A2(new_n945), .A3(new_n712), .ZN(new_n946));
  XNOR2_X1  g521(.A(new_n936), .B(KEYINPUT114), .ZN(new_n947));
  OAI21_X1  g522(.A(new_n935), .B1(new_n946), .B2(new_n947), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n906), .A2(KEYINPUT50), .ZN(new_n949));
  INV_X1    g524(.A(KEYINPUT50), .ZN(new_n950));
  NAND3_X1  g525(.A1(new_n498), .A2(new_n950), .A3(new_n903), .ZN(new_n951));
  AND3_X1   g526(.A1(new_n949), .A2(new_n908), .A3(new_n951), .ZN(new_n952));
  INV_X1    g527(.A(G2090), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n906), .A2(new_n907), .ZN(new_n954));
  NAND3_X1  g529(.A1(new_n498), .A2(KEYINPUT45), .A3(new_n903), .ZN(new_n955));
  NAND3_X1  g530(.A1(new_n954), .A2(new_n908), .A3(new_n955), .ZN(new_n956));
  AOI22_X1  g531(.A1(new_n952), .A2(new_n953), .B1(new_n956), .B2(new_n709), .ZN(new_n957));
  OR2_X1    g532(.A1(new_n957), .A2(KEYINPUT111), .ZN(new_n958));
  NAND2_X1  g533(.A1(G303), .A2(G8), .ZN(new_n959));
  XNOR2_X1  g534(.A(new_n959), .B(KEYINPUT55), .ZN(new_n960));
  INV_X1    g535(.A(new_n960), .ZN(new_n961));
  NAND2_X1  g536(.A1(new_n957), .A2(KEYINPUT111), .ZN(new_n962));
  NAND4_X1  g537(.A1(new_n958), .A2(G8), .A3(new_n961), .A4(new_n962), .ZN(new_n963));
  OR3_X1    g538(.A1(G288), .A2(KEYINPUT112), .A3(new_n945), .ZN(new_n964));
  OAI21_X1  g539(.A(KEYINPUT112), .B1(G288), .B2(new_n945), .ZN(new_n965));
  NAND3_X1  g540(.A1(new_n964), .A2(new_n965), .A3(new_n935), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n966), .A2(KEYINPUT52), .ZN(new_n967));
  AOI21_X1  g542(.A(KEYINPUT52), .B1(G288), .B2(new_n945), .ZN(new_n968));
  NAND4_X1  g543(.A1(new_n964), .A2(new_n965), .A3(new_n968), .A4(new_n935), .ZN(new_n969));
  NAND3_X1  g544(.A1(new_n967), .A2(new_n944), .A3(new_n969), .ZN(new_n970));
  OAI21_X1  g545(.A(new_n948), .B1(new_n963), .B2(new_n970), .ZN(new_n971));
  INV_X1    g546(.A(KEYINPUT115), .ZN(new_n972));
  XNOR2_X1  g547(.A(new_n971), .B(new_n972), .ZN(new_n973));
  INV_X1    g548(.A(new_n970), .ZN(new_n974));
  AND2_X1   g549(.A1(new_n963), .A2(new_n974), .ZN(new_n975));
  INV_X1    g550(.A(KEYINPUT116), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n955), .A2(new_n976), .ZN(new_n977));
  NAND3_X1  g552(.A1(new_n934), .A2(KEYINPUT116), .A3(KEYINPUT45), .ZN(new_n978));
  NAND4_X1  g553(.A1(new_n977), .A2(new_n978), .A3(new_n908), .A4(new_n954), .ZN(new_n979));
  AOI22_X1  g554(.A1(new_n802), .A2(new_n979), .B1(new_n952), .B2(new_n758), .ZN(new_n980));
  NOR3_X1   g555(.A1(new_n980), .A2(new_n932), .A3(G286), .ZN(new_n981));
  INV_X1    g556(.A(KEYINPUT63), .ZN(new_n982));
  NAND3_X1  g557(.A1(new_n958), .A2(G8), .A3(new_n962), .ZN(new_n983));
  AOI21_X1  g558(.A(new_n982), .B1(new_n983), .B2(new_n960), .ZN(new_n984));
  NAND3_X1  g559(.A1(new_n975), .A2(new_n981), .A3(new_n984), .ZN(new_n985));
  OAI21_X1  g560(.A(new_n960), .B1(new_n957), .B2(new_n932), .ZN(new_n986));
  NAND4_X1  g561(.A1(new_n963), .A2(new_n974), .A3(new_n986), .A4(new_n981), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n987), .A2(new_n982), .ZN(new_n988));
  NAND2_X1  g563(.A1(new_n985), .A2(new_n988), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n973), .A2(new_n989), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n975), .A2(new_n986), .ZN(new_n991));
  NOR2_X1   g566(.A1(G168), .A2(new_n932), .ZN(new_n992));
  INV_X1    g567(.A(new_n992), .ZN(new_n993));
  NOR2_X1   g568(.A1(new_n980), .A2(new_n993), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n979), .A2(new_n802), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n952), .A2(new_n758), .ZN(new_n996));
  AOI21_X1  g571(.A(new_n932), .B1(new_n995), .B2(new_n996), .ZN(new_n997));
  INV_X1    g572(.A(KEYINPUT121), .ZN(new_n998));
  OAI21_X1  g573(.A(new_n993), .B1(new_n997), .B2(new_n998), .ZN(new_n999));
  NOR3_X1   g574(.A1(new_n980), .A2(KEYINPUT121), .A3(new_n932), .ZN(new_n1000));
  OAI21_X1  g575(.A(KEYINPUT51), .B1(new_n999), .B2(new_n1000), .ZN(new_n1001));
  INV_X1    g576(.A(KEYINPUT122), .ZN(new_n1002));
  AOI21_X1  g577(.A(KEYINPUT51), .B1(new_n997), .B2(new_n1002), .ZN(new_n1003));
  OAI21_X1  g578(.A(KEYINPUT122), .B1(new_n980), .B2(new_n932), .ZN(new_n1004));
  NAND3_X1  g579(.A1(new_n1003), .A2(new_n993), .A3(new_n1004), .ZN(new_n1005));
  AOI21_X1  g580(.A(new_n994), .B1(new_n1001), .B2(new_n1005), .ZN(new_n1006));
  XOR2_X1   g581(.A(KEYINPUT123), .B(G1961), .Z(new_n1007));
  NAND3_X1  g582(.A1(new_n949), .A2(new_n908), .A3(new_n951), .ZN(new_n1008));
  INV_X1    g583(.A(KEYINPUT120), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n1008), .A2(new_n1009), .ZN(new_n1010));
  NAND4_X1  g585(.A1(new_n949), .A2(KEYINPUT120), .A3(new_n908), .A4(new_n951), .ZN(new_n1011));
  AOI21_X1  g586(.A(new_n1007), .B1(new_n1010), .B2(new_n1011), .ZN(new_n1012));
  INV_X1    g587(.A(G2078), .ZN(new_n1013));
  OAI21_X1  g588(.A(new_n908), .B1(new_n934), .B2(KEYINPUT45), .ZN(new_n1014));
  INV_X1    g589(.A(new_n955), .ZN(new_n1015));
  NOR2_X1   g590(.A1(new_n1014), .A2(new_n1015), .ZN(new_n1016));
  INV_X1    g591(.A(KEYINPUT125), .ZN(new_n1017));
  NAND4_X1  g592(.A1(new_n954), .A2(new_n1017), .A3(new_n908), .A4(new_n955), .ZN(new_n1018));
  AOI22_X1  g593(.A1(new_n1013), .A2(new_n1016), .B1(new_n1018), .B2(KEYINPUT53), .ZN(new_n1019));
  INV_X1    g594(.A(KEYINPUT53), .ZN(new_n1020));
  NOR4_X1   g595(.A1(new_n956), .A2(new_n1017), .A3(new_n1020), .A4(G2078), .ZN(new_n1021));
  NOR3_X1   g596(.A1(new_n1012), .A2(new_n1019), .A3(new_n1021), .ZN(new_n1022));
  AOI21_X1  g597(.A(KEYINPUT54), .B1(new_n1022), .B2(G301), .ZN(new_n1023));
  INV_X1    g598(.A(KEYINPUT124), .ZN(new_n1024));
  AOI21_X1  g599(.A(KEYINPUT53), .B1(new_n1016), .B2(new_n1013), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n1013), .A2(KEYINPUT53), .ZN(new_n1026));
  NOR2_X1   g601(.A1(new_n979), .A2(new_n1026), .ZN(new_n1027));
  NOR3_X1   g602(.A1(new_n1012), .A2(new_n1025), .A3(new_n1027), .ZN(new_n1028));
  OAI21_X1  g603(.A(new_n1024), .B1(new_n1028), .B2(G301), .ZN(new_n1029));
  NAND2_X1  g604(.A1(new_n1010), .A2(new_n1011), .ZN(new_n1030));
  INV_X1    g605(.A(new_n1007), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n1030), .A2(new_n1031), .ZN(new_n1032));
  INV_X1    g607(.A(new_n1025), .ZN(new_n1033));
  INV_X1    g608(.A(new_n1027), .ZN(new_n1034));
  NAND3_X1  g609(.A1(new_n1032), .A2(new_n1033), .A3(new_n1034), .ZN(new_n1035));
  NAND3_X1  g610(.A1(new_n1035), .A2(KEYINPUT124), .A3(G171), .ZN(new_n1036));
  NAND3_X1  g611(.A1(new_n1023), .A2(new_n1029), .A3(new_n1036), .ZN(new_n1037));
  NOR2_X1   g612(.A1(new_n1019), .A2(new_n1021), .ZN(new_n1038));
  NAND3_X1  g613(.A1(new_n1038), .A2(G171), .A3(new_n1032), .ZN(new_n1039));
  OAI211_X1 g614(.A(new_n1039), .B(KEYINPUT54), .C1(G171), .C2(new_n1028), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n1037), .A2(new_n1040), .ZN(new_n1041));
  XNOR2_X1  g616(.A(KEYINPUT56), .B(G2072), .ZN(new_n1042));
  AOI22_X1  g617(.A1(new_n1016), .A2(new_n1042), .B1(new_n1008), .B2(new_n769), .ZN(new_n1043));
  NAND2_X1  g618(.A1(KEYINPUT117), .A2(KEYINPUT57), .ZN(new_n1044));
  NOR2_X1   g619(.A1(KEYINPUT117), .A2(KEYINPUT57), .ZN(new_n1045));
  XNOR2_X1  g620(.A(new_n1045), .B(KEYINPUT118), .ZN(new_n1046));
  AND3_X1   g621(.A1(new_n558), .A2(new_n1044), .A3(new_n1046), .ZN(new_n1047));
  AOI21_X1  g622(.A(new_n1046), .B1(new_n558), .B2(new_n1044), .ZN(new_n1048));
  NOR2_X1   g623(.A1(new_n1047), .A2(new_n1048), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n1043), .A2(new_n1049), .ZN(new_n1050));
  AOI21_X1  g625(.A(G1348), .B1(new_n1010), .B2(new_n1011), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n934), .A2(new_n908), .ZN(new_n1052));
  NOR2_X1   g627(.A1(new_n1052), .A2(G2067), .ZN(new_n1053));
  INV_X1    g628(.A(KEYINPUT119), .ZN(new_n1054));
  XNOR2_X1  g629(.A(new_n1053), .B(new_n1054), .ZN(new_n1055));
  OAI211_X1 g630(.A(new_n1050), .B(new_n604), .C1(new_n1051), .C2(new_n1055), .ZN(new_n1056));
  NOR2_X1   g631(.A1(new_n952), .A2(G1956), .ZN(new_n1057));
  INV_X1    g632(.A(new_n1042), .ZN(new_n1058));
  NOR2_X1   g633(.A1(new_n956), .A2(new_n1058), .ZN(new_n1059));
  OAI22_X1  g634(.A1(new_n1057), .A2(new_n1059), .B1(new_n1047), .B2(new_n1048), .ZN(new_n1060));
  AND2_X1   g635(.A1(new_n1056), .A2(new_n1060), .ZN(new_n1061));
  INV_X1    g636(.A(KEYINPUT61), .ZN(new_n1062));
  AND2_X1   g637(.A1(new_n1043), .A2(new_n1049), .ZN(new_n1063));
  NOR2_X1   g638(.A1(new_n1043), .A2(new_n1049), .ZN(new_n1064));
  OAI21_X1  g639(.A(new_n1062), .B1(new_n1063), .B2(new_n1064), .ZN(new_n1065));
  NAND3_X1  g640(.A1(new_n1060), .A2(KEYINPUT61), .A3(new_n1050), .ZN(new_n1066));
  XOR2_X1   g641(.A(KEYINPUT58), .B(G1341), .Z(new_n1067));
  NAND2_X1  g642(.A1(new_n1052), .A2(new_n1067), .ZN(new_n1068));
  OAI21_X1  g643(.A(new_n1068), .B1(new_n956), .B2(G1996), .ZN(new_n1069));
  AND3_X1   g644(.A1(new_n1069), .A2(KEYINPUT59), .A3(new_n541), .ZN(new_n1070));
  AOI21_X1  g645(.A(KEYINPUT59), .B1(new_n1069), .B2(new_n541), .ZN(new_n1071));
  NOR2_X1   g646(.A1(new_n1070), .A2(new_n1071), .ZN(new_n1072));
  NAND3_X1  g647(.A1(new_n1065), .A2(new_n1066), .A3(new_n1072), .ZN(new_n1073));
  INV_X1    g648(.A(new_n1055), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n604), .A2(KEYINPUT60), .ZN(new_n1075));
  INV_X1    g650(.A(new_n1051), .ZN(new_n1076));
  INV_X1    g651(.A(KEYINPUT60), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n597), .A2(new_n1077), .ZN(new_n1078));
  NAND4_X1  g653(.A1(new_n1074), .A2(new_n1075), .A3(new_n1076), .A4(new_n1078), .ZN(new_n1079));
  OAI211_X1 g654(.A(KEYINPUT60), .B(new_n604), .C1(new_n1055), .C2(new_n1051), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1079), .A2(new_n1080), .ZN(new_n1081));
  OAI21_X1  g656(.A(new_n1061), .B1(new_n1073), .B2(new_n1081), .ZN(new_n1082));
  AOI21_X1  g657(.A(new_n1006), .B1(new_n1041), .B2(new_n1082), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n1029), .A2(new_n1036), .ZN(new_n1084));
  INV_X1    g659(.A(KEYINPUT62), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n1084), .A2(new_n1085), .ZN(new_n1086));
  AOI21_X1  g661(.A(new_n991), .B1(new_n1083), .B2(new_n1086), .ZN(new_n1087));
  NAND2_X1  g662(.A1(new_n1084), .A2(KEYINPUT62), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n1006), .A2(new_n1088), .ZN(new_n1089));
  AOI21_X1  g664(.A(new_n990), .B1(new_n1087), .B2(new_n1089), .ZN(new_n1090));
  XOR2_X1   g665(.A(G290), .B(G1986), .Z(new_n1091));
  OAI21_X1  g666(.A(new_n928), .B1(new_n909), .B2(new_n1091), .ZN(new_n1092));
  OAI21_X1  g667(.A(new_n931), .B1(new_n1090), .B2(new_n1092), .ZN(G329));
  assign    G231 = 1'b0;
  NAND3_X1  g668(.A1(new_n652), .A2(G319), .A3(new_n668), .ZN(new_n1095));
  NAND2_X1  g669(.A1(new_n1095), .A2(KEYINPUT126), .ZN(new_n1096));
  INV_X1    g670(.A(KEYINPUT126), .ZN(new_n1097));
  NAND4_X1  g671(.A1(new_n652), .A2(new_n1097), .A3(G319), .A4(new_n668), .ZN(new_n1098));
  AOI21_X1  g672(.A(G229), .B1(new_n1096), .B2(new_n1098), .ZN(new_n1099));
  NAND3_X1  g673(.A1(new_n901), .A2(new_n858), .A3(new_n1099), .ZN(G225));
  NAND2_X1  g674(.A1(G225), .A2(KEYINPUT127), .ZN(new_n1101));
  INV_X1    g675(.A(KEYINPUT127), .ZN(new_n1102));
  NAND4_X1  g676(.A1(new_n901), .A2(new_n1102), .A3(new_n1099), .A4(new_n858), .ZN(new_n1103));
  NAND2_X1  g677(.A1(new_n1101), .A2(new_n1103), .ZN(G308));
endmodule


