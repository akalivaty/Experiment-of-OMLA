//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 1 1 0 0 0 1 1 0 1 1 1 0 0 0 0 1 0 0 0 0 1 0 1 0 0 0 0 0 0 1 1 1 0 1 1 1 0 1 1 1 1 1 1 0 1 0 0 0 1 1 1 0 1 0 0 1 1 0 1 1 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:30:56 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n444, new_n448, new_n452, new_n453, new_n454, new_n455,
    new_n456, new_n457, new_n460, new_n461, new_n462, new_n463, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n528, new_n529, new_n530, new_n531, new_n532,
    new_n533, new_n534, new_n536, new_n537, new_n538, new_n539, new_n540,
    new_n541, new_n542, new_n545, new_n546, new_n547, new_n548, new_n549,
    new_n550, new_n551, new_n552, new_n553, new_n554, new_n555, new_n558,
    new_n559, new_n560, new_n562, new_n563, new_n564, new_n565, new_n566,
    new_n567, new_n568, new_n569, new_n570, new_n571, new_n572, new_n576,
    new_n577, new_n578, new_n580, new_n581, new_n582, new_n583, new_n584,
    new_n585, new_n586, new_n588, new_n589, new_n590, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n604, new_n605, new_n608, new_n610, new_n611, new_n612,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n818, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1193, new_n1194, new_n1195;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  XNOR2_X1  g008(.A(KEYINPUT64), .B(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(new_n436));
  XNOR2_X1  g011(.A(new_n436), .B(KEYINPUT65), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(new_n444));
  XNOR2_X1  g019(.A(new_n444), .B(KEYINPUT66), .ZN(G259));
  BUF_X1    g020(.A(G452), .Z(G391));
  AND2_X1   g021(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XOR2_X1   g023(.A(new_n448), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g024(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g025(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  OR4_X1    g026(.A1(G221), .A2(G220), .A3(G219), .A4(G218), .ZN(new_n452));
  XNOR2_X1  g027(.A(new_n452), .B(KEYINPUT2), .ZN(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  XNOR2_X1  g029(.A(KEYINPUT67), .B(KEYINPUT68), .ZN(new_n455));
  NAND4_X1  g030(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n456));
  XNOR2_X1  g031(.A(new_n455), .B(new_n456), .ZN(new_n457));
  NAND2_X1  g032(.A1(new_n454), .A2(new_n457), .ZN(G261));
  INV_X1    g033(.A(G261), .ZN(G325));
  NAND2_X1  g034(.A1(new_n453), .A2(G2106), .ZN(new_n460));
  INV_X1    g035(.A(G567), .ZN(new_n461));
  OR2_X1    g036(.A1(new_n457), .A2(new_n461), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n460), .A2(new_n462), .ZN(new_n463));
  INV_X1    g038(.A(new_n463), .ZN(G319));
  INV_X1    g039(.A(G2105), .ZN(new_n465));
  XNOR2_X1  g040(.A(KEYINPUT3), .B(G2104), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n466), .A2(G125), .ZN(new_n467));
  NAND2_X1  g042(.A1(G113), .A2(G2104), .ZN(new_n468));
  AOI21_X1  g043(.A(new_n465), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  INV_X1    g044(.A(new_n469), .ZN(new_n470));
  NAND3_X1  g045(.A1(new_n466), .A2(G137), .A3(new_n465), .ZN(new_n471));
  INV_X1    g046(.A(G2104), .ZN(new_n472));
  NOR2_X1   g047(.A1(new_n472), .A2(G2105), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n473), .A2(G101), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n471), .A2(new_n474), .ZN(new_n475));
  INV_X1    g050(.A(new_n475), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n470), .A2(new_n476), .ZN(new_n477));
  INV_X1    g052(.A(new_n477), .ZN(G160));
  OR2_X1    g053(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n479));
  NAND2_X1  g054(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n480));
  AOI21_X1  g055(.A(G2105), .B1(new_n479), .B2(new_n480), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n481), .A2(G136), .ZN(new_n482));
  NOR2_X1   g057(.A1(new_n465), .A2(G112), .ZN(new_n483));
  OAI21_X1  g058(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n484));
  OAI21_X1  g059(.A(new_n482), .B1(new_n483), .B2(new_n484), .ZN(new_n485));
  AOI21_X1  g060(.A(new_n465), .B1(new_n479), .B2(new_n480), .ZN(new_n486));
  XOR2_X1   g061(.A(new_n486), .B(KEYINPUT69), .Z(new_n487));
  AOI21_X1  g062(.A(new_n485), .B1(new_n487), .B2(G124), .ZN(new_n488));
  XOR2_X1   g063(.A(new_n488), .B(KEYINPUT70), .Z(G162));
  INV_X1    g064(.A(G138), .ZN(new_n490));
  NOR2_X1   g065(.A1(new_n490), .A2(G2105), .ZN(new_n491));
  AND2_X1   g066(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n492));
  NOR2_X1   g067(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n493));
  OAI21_X1  g068(.A(new_n491), .B1(new_n492), .B2(new_n493), .ZN(new_n494));
  NAND2_X1  g069(.A1(new_n494), .A2(KEYINPUT71), .ZN(new_n495));
  INV_X1    g070(.A(KEYINPUT71), .ZN(new_n496));
  NAND3_X1  g071(.A1(new_n466), .A2(new_n496), .A3(new_n491), .ZN(new_n497));
  NAND3_X1  g072(.A1(new_n495), .A2(KEYINPUT4), .A3(new_n497), .ZN(new_n498));
  INV_X1    g073(.A(KEYINPUT4), .ZN(new_n499));
  NAND3_X1  g074(.A1(new_n494), .A2(KEYINPUT71), .A3(new_n499), .ZN(new_n500));
  OAI211_X1 g075(.A(G126), .B(G2105), .C1(new_n492), .C2(new_n493), .ZN(new_n501));
  OR2_X1    g076(.A1(G102), .A2(G2105), .ZN(new_n502));
  INV_X1    g077(.A(G114), .ZN(new_n503));
  NAND2_X1  g078(.A1(new_n503), .A2(G2105), .ZN(new_n504));
  NAND3_X1  g079(.A1(new_n502), .A2(new_n504), .A3(G2104), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n501), .A2(new_n505), .ZN(new_n506));
  INV_X1    g081(.A(new_n506), .ZN(new_n507));
  NAND3_X1  g082(.A1(new_n498), .A2(new_n500), .A3(new_n507), .ZN(new_n508));
  INV_X1    g083(.A(new_n508), .ZN(G164));
  INV_X1    g084(.A(G543), .ZN(new_n510));
  NAND2_X1  g085(.A1(KEYINPUT72), .A2(G651), .ZN(new_n511));
  INV_X1    g086(.A(KEYINPUT6), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  NAND3_X1  g088(.A1(KEYINPUT72), .A2(KEYINPUT6), .A3(G651), .ZN(new_n514));
  AOI21_X1  g089(.A(new_n510), .B1(new_n513), .B2(new_n514), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n515), .A2(G50), .ZN(new_n516));
  INV_X1    g091(.A(G88), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n513), .A2(new_n514), .ZN(new_n518));
  OR2_X1    g093(.A1(KEYINPUT5), .A2(G543), .ZN(new_n519));
  NAND2_X1  g094(.A1(KEYINPUT5), .A2(G543), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n518), .A2(new_n521), .ZN(new_n522));
  OAI21_X1  g097(.A(new_n516), .B1(new_n517), .B2(new_n522), .ZN(new_n523));
  AOI22_X1  g098(.A1(new_n521), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n524));
  INV_X1    g099(.A(G651), .ZN(new_n525));
  NOR2_X1   g100(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  NOR2_X1   g101(.A1(new_n523), .A2(new_n526), .ZN(G166));
  NAND2_X1  g102(.A1(new_n515), .A2(G51), .ZN(new_n528));
  NAND3_X1  g103(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n529));
  XNOR2_X1  g104(.A(new_n529), .B(KEYINPUT7), .ZN(new_n530));
  NAND3_X1  g105(.A1(new_n521), .A2(G63), .A3(G651), .ZN(new_n531));
  NAND3_X1  g106(.A1(new_n528), .A2(new_n530), .A3(new_n531), .ZN(new_n532));
  AOI22_X1  g107(.A1(new_n513), .A2(new_n514), .B1(new_n519), .B2(new_n520), .ZN(new_n533));
  AND2_X1   g108(.A1(new_n533), .A2(G89), .ZN(new_n534));
  NOR2_X1   g109(.A1(new_n532), .A2(new_n534), .ZN(G168));
  NAND2_X1  g110(.A1(G77), .A2(G543), .ZN(new_n536));
  AND2_X1   g111(.A1(new_n519), .A2(new_n520), .ZN(new_n537));
  INV_X1    g112(.A(G64), .ZN(new_n538));
  OAI21_X1  g113(.A(new_n536), .B1(new_n537), .B2(new_n538), .ZN(new_n539));
  NAND2_X1  g114(.A1(new_n539), .A2(G651), .ZN(new_n540));
  NAND2_X1  g115(.A1(new_n515), .A2(G52), .ZN(new_n541));
  NAND2_X1  g116(.A1(new_n533), .A2(G90), .ZN(new_n542));
  NAND3_X1  g117(.A1(new_n540), .A2(new_n541), .A3(new_n542), .ZN(G301));
  INV_X1    g118(.A(G301), .ZN(G171));
  INV_X1    g119(.A(G56), .ZN(new_n545));
  INV_X1    g120(.A(G68), .ZN(new_n546));
  OAI22_X1  g121(.A1(new_n537), .A2(new_n545), .B1(new_n546), .B2(new_n510), .ZN(new_n547));
  NAND2_X1  g122(.A1(new_n547), .A2(KEYINPUT73), .ZN(new_n548));
  INV_X1    g123(.A(KEYINPUT73), .ZN(new_n549));
  OAI221_X1 g124(.A(new_n549), .B1(new_n546), .B2(new_n510), .C1(new_n537), .C2(new_n545), .ZN(new_n550));
  NAND3_X1  g125(.A1(new_n548), .A2(G651), .A3(new_n550), .ZN(new_n551));
  XNOR2_X1  g126(.A(KEYINPUT74), .B(G43), .ZN(new_n552));
  AOI22_X1  g127(.A1(new_n533), .A2(G81), .B1(new_n515), .B2(new_n552), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n551), .A2(new_n553), .ZN(new_n554));
  INV_X1    g129(.A(new_n554), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n555), .A2(G860), .ZN(G153));
  NAND4_X1  g131(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g132(.A1(G1), .A2(G3), .ZN(new_n558));
  XNOR2_X1  g133(.A(new_n558), .B(KEYINPUT75), .ZN(new_n559));
  XNOR2_X1  g134(.A(new_n559), .B(KEYINPUT8), .ZN(new_n560));
  NAND4_X1  g135(.A1(G319), .A2(G483), .A3(G661), .A4(new_n560), .ZN(G188));
  INV_X1    g136(.A(new_n514), .ZN(new_n562));
  AOI21_X1  g137(.A(KEYINPUT6), .B1(KEYINPUT72), .B2(G651), .ZN(new_n563));
  OAI211_X1 g138(.A(G53), .B(G543), .C1(new_n562), .C2(new_n563), .ZN(new_n564));
  INV_X1    g139(.A(KEYINPUT76), .ZN(new_n565));
  OAI21_X1  g140(.A(new_n564), .B1(new_n565), .B2(KEYINPUT9), .ZN(new_n566));
  XOR2_X1   g141(.A(KEYINPUT76), .B(KEYINPUT9), .Z(new_n567));
  NAND3_X1  g142(.A1(new_n515), .A2(G53), .A3(new_n567), .ZN(new_n568));
  AND2_X1   g143(.A1(new_n566), .A2(new_n568), .ZN(new_n569));
  AOI22_X1  g144(.A1(new_n521), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n570));
  INV_X1    g145(.A(G91), .ZN(new_n571));
  OAI22_X1  g146(.A1(new_n570), .A2(new_n525), .B1(new_n522), .B2(new_n571), .ZN(new_n572));
  OR2_X1    g147(.A1(new_n569), .A2(new_n572), .ZN(G299));
  INV_X1    g148(.A(G168), .ZN(G286));
  INV_X1    g149(.A(G166), .ZN(G303));
  OR2_X1    g150(.A1(new_n521), .A2(G74), .ZN(new_n576));
  AOI22_X1  g151(.A1(new_n576), .A2(G651), .B1(new_n533), .B2(G87), .ZN(new_n577));
  NAND2_X1  g152(.A1(new_n515), .A2(G49), .ZN(new_n578));
  NAND2_X1  g153(.A1(new_n577), .A2(new_n578), .ZN(G288));
  NAND2_X1  g154(.A1(G73), .A2(G543), .ZN(new_n580));
  XNOR2_X1  g155(.A(new_n580), .B(KEYINPUT77), .ZN(new_n581));
  INV_X1    g156(.A(G61), .ZN(new_n582));
  AOI21_X1  g157(.A(new_n582), .B1(new_n519), .B2(new_n520), .ZN(new_n583));
  OAI21_X1  g158(.A(G651), .B1(new_n581), .B2(new_n583), .ZN(new_n584));
  NAND3_X1  g159(.A1(new_n518), .A2(G48), .A3(G543), .ZN(new_n585));
  NAND2_X1  g160(.A1(new_n533), .A2(G86), .ZN(new_n586));
  NAND3_X1  g161(.A1(new_n584), .A2(new_n585), .A3(new_n586), .ZN(G305));
  NAND2_X1  g162(.A1(new_n533), .A2(G85), .ZN(new_n588));
  NAND2_X1  g163(.A1(new_n515), .A2(G47), .ZN(new_n589));
  AOI22_X1  g164(.A1(new_n521), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n590));
  OAI211_X1 g165(.A(new_n588), .B(new_n589), .C1(new_n525), .C2(new_n590), .ZN(G290));
  INV_X1    g166(.A(G868), .ZN(new_n592));
  NOR2_X1   g167(.A1(G301), .A2(new_n592), .ZN(new_n593));
  NAND2_X1  g168(.A1(new_n533), .A2(G92), .ZN(new_n594));
  XOR2_X1   g169(.A(new_n594), .B(KEYINPUT10), .Z(new_n595));
  NAND2_X1  g170(.A1(G79), .A2(G543), .ZN(new_n596));
  INV_X1    g171(.A(G66), .ZN(new_n597));
  OAI21_X1  g172(.A(new_n596), .B1(new_n537), .B2(new_n597), .ZN(new_n598));
  AOI22_X1  g173(.A1(new_n598), .A2(G651), .B1(G54), .B2(new_n515), .ZN(new_n599));
  NAND2_X1  g174(.A1(new_n595), .A2(new_n599), .ZN(new_n600));
  XNOR2_X1  g175(.A(new_n600), .B(KEYINPUT78), .ZN(new_n601));
  AOI21_X1  g176(.A(new_n593), .B1(new_n601), .B2(new_n592), .ZN(G284));
  AOI21_X1  g177(.A(new_n593), .B1(new_n601), .B2(new_n592), .ZN(G321));
  NAND2_X1  g178(.A1(G286), .A2(G868), .ZN(new_n604));
  NOR2_X1   g179(.A1(new_n569), .A2(new_n572), .ZN(new_n605));
  OAI21_X1  g180(.A(new_n604), .B1(G868), .B2(new_n605), .ZN(G297));
  XOR2_X1   g181(.A(G297), .B(KEYINPUT79), .Z(G280));
  INV_X1    g182(.A(G559), .ZN(new_n608));
  OAI21_X1  g183(.A(new_n601), .B1(new_n608), .B2(G860), .ZN(G148));
  NOR2_X1   g184(.A1(new_n554), .A2(G868), .ZN(new_n610));
  NAND2_X1  g185(.A1(new_n601), .A2(new_n608), .ZN(new_n611));
  XNOR2_X1  g186(.A(new_n611), .B(KEYINPUT80), .ZN(new_n612));
  AOI21_X1  g187(.A(new_n610), .B1(new_n612), .B2(G868), .ZN(G323));
  XNOR2_X1  g188(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g189(.A1(new_n466), .A2(new_n473), .ZN(new_n615));
  XOR2_X1   g190(.A(new_n615), .B(KEYINPUT12), .Z(new_n616));
  XOR2_X1   g191(.A(KEYINPUT81), .B(KEYINPUT13), .Z(new_n617));
  XNOR2_X1  g192(.A(new_n616), .B(new_n617), .ZN(new_n618));
  XNOR2_X1  g193(.A(KEYINPUT82), .B(G2100), .ZN(new_n619));
  NAND2_X1  g194(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  XOR2_X1   g195(.A(new_n620), .B(KEYINPUT83), .Z(new_n621));
  NAND2_X1  g196(.A1(new_n481), .A2(G135), .ZN(new_n622));
  XOR2_X1   g197(.A(new_n622), .B(KEYINPUT84), .Z(new_n623));
  NAND2_X1  g198(.A1(new_n487), .A2(G123), .ZN(new_n624));
  OR2_X1    g199(.A1(G99), .A2(G2105), .ZN(new_n625));
  OAI211_X1 g200(.A(new_n625), .B(G2104), .C1(G111), .C2(new_n465), .ZN(new_n626));
  NAND3_X1  g201(.A1(new_n623), .A2(new_n624), .A3(new_n626), .ZN(new_n627));
  NAND2_X1  g202(.A1(new_n627), .A2(G2096), .ZN(new_n628));
  OR2_X1    g203(.A1(new_n627), .A2(G2096), .ZN(new_n629));
  OR2_X1    g204(.A1(new_n618), .A2(new_n619), .ZN(new_n630));
  NAND4_X1  g205(.A1(new_n621), .A2(new_n628), .A3(new_n629), .A4(new_n630), .ZN(G156));
  XNOR2_X1  g206(.A(KEYINPUT15), .B(G2435), .ZN(new_n632));
  XNOR2_X1  g207(.A(new_n632), .B(G2438), .ZN(new_n633));
  XNOR2_X1  g208(.A(G2427), .B(G2430), .ZN(new_n634));
  XNOR2_X1  g209(.A(new_n634), .B(KEYINPUT86), .ZN(new_n635));
  NAND2_X1  g210(.A1(new_n633), .A2(new_n635), .ZN(new_n636));
  NAND2_X1  g211(.A1(new_n636), .A2(KEYINPUT14), .ZN(new_n637));
  XNOR2_X1  g212(.A(new_n637), .B(KEYINPUT87), .ZN(new_n638));
  OAI21_X1  g213(.A(new_n638), .B1(new_n633), .B2(new_n635), .ZN(new_n639));
  XNOR2_X1  g214(.A(G2443), .B(G2446), .ZN(new_n640));
  XNOR2_X1  g215(.A(new_n639), .B(new_n640), .ZN(new_n641));
  XNOR2_X1  g216(.A(G1341), .B(G1348), .ZN(new_n642));
  XNOR2_X1  g217(.A(KEYINPUT85), .B(KEYINPUT16), .ZN(new_n643));
  XOR2_X1   g218(.A(new_n642), .B(new_n643), .Z(new_n644));
  XNOR2_X1  g219(.A(new_n641), .B(new_n644), .ZN(new_n645));
  XNOR2_X1  g220(.A(G2451), .B(G2454), .ZN(new_n646));
  XNOR2_X1  g221(.A(new_n646), .B(KEYINPUT88), .ZN(new_n647));
  NAND2_X1  g222(.A1(new_n645), .A2(new_n647), .ZN(new_n648));
  NAND2_X1  g223(.A1(new_n648), .A2(G14), .ZN(new_n649));
  NOR2_X1   g224(.A1(new_n645), .A2(new_n647), .ZN(new_n650));
  NOR2_X1   g225(.A1(new_n649), .A2(new_n650), .ZN(G401));
  XOR2_X1   g226(.A(G2072), .B(G2078), .Z(new_n652));
  XOR2_X1   g227(.A(G2084), .B(G2090), .Z(new_n653));
  XNOR2_X1  g228(.A(G2067), .B(G2678), .ZN(new_n654));
  NAND2_X1  g229(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  AOI21_X1  g230(.A(new_n652), .B1(new_n655), .B2(KEYINPUT18), .ZN(new_n656));
  XNOR2_X1  g231(.A(new_n656), .B(KEYINPUT89), .ZN(new_n657));
  XNOR2_X1  g232(.A(new_n657), .B(G2100), .ZN(new_n658));
  INV_X1    g233(.A(KEYINPUT18), .ZN(new_n659));
  NAND2_X1  g234(.A1(new_n655), .A2(KEYINPUT17), .ZN(new_n660));
  NOR2_X1   g235(.A1(new_n653), .A2(new_n654), .ZN(new_n661));
  OAI21_X1  g236(.A(new_n659), .B1(new_n660), .B2(new_n661), .ZN(new_n662));
  XOR2_X1   g237(.A(new_n662), .B(G2096), .Z(new_n663));
  XNOR2_X1  g238(.A(new_n658), .B(new_n663), .ZN(G227));
  XOR2_X1   g239(.A(G1971), .B(G1976), .Z(new_n665));
  XNOR2_X1  g240(.A(new_n665), .B(KEYINPUT19), .ZN(new_n666));
  XOR2_X1   g241(.A(G1956), .B(G2474), .Z(new_n667));
  XOR2_X1   g242(.A(G1961), .B(G1966), .Z(new_n668));
  AND2_X1   g243(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  NAND2_X1  g244(.A1(new_n666), .A2(new_n669), .ZN(new_n670));
  XNOR2_X1  g245(.A(new_n670), .B(KEYINPUT20), .ZN(new_n671));
  NOR2_X1   g246(.A1(new_n667), .A2(new_n668), .ZN(new_n672));
  NOR3_X1   g247(.A1(new_n666), .A2(new_n669), .A3(new_n672), .ZN(new_n673));
  AOI21_X1  g248(.A(new_n673), .B1(new_n666), .B2(new_n672), .ZN(new_n674));
  NAND2_X1  g249(.A1(new_n671), .A2(new_n674), .ZN(new_n675));
  XNOR2_X1  g250(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n676));
  XOR2_X1   g251(.A(new_n675), .B(new_n676), .Z(new_n677));
  XOR2_X1   g252(.A(G1991), .B(G1996), .Z(new_n678));
  INV_X1    g253(.A(new_n678), .ZN(new_n679));
  XNOR2_X1  g254(.A(new_n677), .B(new_n679), .ZN(new_n680));
  XNOR2_X1  g255(.A(G1981), .B(G1986), .ZN(new_n681));
  AND2_X1   g256(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  NOR2_X1   g257(.A1(new_n680), .A2(new_n681), .ZN(new_n683));
  OR2_X1    g258(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  INV_X1    g259(.A(new_n684), .ZN(G229));
  NOR2_X1   g260(.A1(G29), .A2(G35), .ZN(new_n686));
  AOI21_X1  g261(.A(new_n686), .B1(G162), .B2(G29), .ZN(new_n687));
  XOR2_X1   g262(.A(new_n687), .B(KEYINPUT29), .Z(new_n688));
  INV_X1    g263(.A(G2090), .ZN(new_n689));
  OR2_X1    g264(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  INV_X1    g265(.A(G16), .ZN(new_n691));
  NAND2_X1  g266(.A1(new_n691), .A2(G5), .ZN(new_n692));
  OAI21_X1  g267(.A(new_n692), .B1(G171), .B2(new_n691), .ZN(new_n693));
  XNOR2_X1  g268(.A(new_n693), .B(G1961), .ZN(new_n694));
  INV_X1    g269(.A(G34), .ZN(new_n695));
  AOI21_X1  g270(.A(G29), .B1(new_n695), .B2(KEYINPUT24), .ZN(new_n696));
  OAI21_X1  g271(.A(new_n696), .B1(KEYINPUT24), .B2(new_n695), .ZN(new_n697));
  INV_X1    g272(.A(G29), .ZN(new_n698));
  OAI21_X1  g273(.A(new_n697), .B1(new_n477), .B2(new_n698), .ZN(new_n699));
  XNOR2_X1  g274(.A(new_n699), .B(G2084), .ZN(new_n700));
  OR2_X1    g275(.A1(new_n627), .A2(new_n698), .ZN(new_n701));
  INV_X1    g276(.A(G28), .ZN(new_n702));
  OR2_X1    g277(.A1(new_n702), .A2(KEYINPUT30), .ZN(new_n703));
  AOI21_X1  g278(.A(G29), .B1(new_n702), .B2(KEYINPUT30), .ZN(new_n704));
  OR2_X1    g279(.A1(KEYINPUT31), .A2(G11), .ZN(new_n705));
  NAND2_X1  g280(.A1(KEYINPUT31), .A2(G11), .ZN(new_n706));
  AOI22_X1  g281(.A1(new_n703), .A2(new_n704), .B1(new_n705), .B2(new_n706), .ZN(new_n707));
  AND3_X1   g282(.A1(new_n700), .A2(new_n701), .A3(new_n707), .ZN(new_n708));
  AND2_X1   g283(.A1(new_n698), .A2(G33), .ZN(new_n709));
  NAND3_X1  g284(.A1(new_n465), .A2(G103), .A3(G2104), .ZN(new_n710));
  XNOR2_X1  g285(.A(new_n710), .B(KEYINPUT25), .ZN(new_n711));
  NAND2_X1  g286(.A1(new_n466), .A2(G127), .ZN(new_n712));
  NAND2_X1  g287(.A1(G115), .A2(G2104), .ZN(new_n713));
  AOI21_X1  g288(.A(new_n465), .B1(new_n712), .B2(new_n713), .ZN(new_n714));
  AOI211_X1 g289(.A(new_n711), .B(new_n714), .C1(G139), .C2(new_n481), .ZN(new_n715));
  INV_X1    g290(.A(KEYINPUT96), .ZN(new_n716));
  XNOR2_X1  g291(.A(new_n715), .B(new_n716), .ZN(new_n717));
  AOI21_X1  g292(.A(new_n709), .B1(new_n717), .B2(G29), .ZN(new_n718));
  INV_X1    g293(.A(new_n718), .ZN(new_n719));
  OAI21_X1  g294(.A(new_n708), .B1(new_n719), .B2(G2072), .ZN(new_n720));
  AOI211_X1 g295(.A(new_n694), .B(new_n720), .C1(G2072), .C2(new_n719), .ZN(new_n721));
  NAND2_X1  g296(.A1(new_n688), .A2(new_n689), .ZN(new_n722));
  NAND2_X1  g297(.A1(new_n691), .A2(G20), .ZN(new_n723));
  XOR2_X1   g298(.A(new_n723), .B(KEYINPUT23), .Z(new_n724));
  AOI21_X1  g299(.A(new_n724), .B1(G299), .B2(G16), .ZN(new_n725));
  XNOR2_X1  g300(.A(new_n725), .B(G1956), .ZN(new_n726));
  NAND2_X1  g301(.A1(new_n691), .A2(G21), .ZN(new_n727));
  OAI21_X1  g302(.A(new_n727), .B1(G168), .B2(new_n691), .ZN(new_n728));
  OR2_X1    g303(.A1(new_n728), .A2(G1966), .ZN(new_n729));
  NOR2_X1   g304(.A1(G164), .A2(new_n698), .ZN(new_n730));
  AOI21_X1  g305(.A(new_n730), .B1(G27), .B2(new_n698), .ZN(new_n731));
  INV_X1    g306(.A(G2078), .ZN(new_n732));
  OR2_X1    g307(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  AOI22_X1  g308(.A1(new_n731), .A2(new_n732), .B1(G1966), .B2(new_n728), .ZN(new_n734));
  AND4_X1   g309(.A1(new_n726), .A2(new_n729), .A3(new_n733), .A4(new_n734), .ZN(new_n735));
  NAND4_X1  g310(.A1(new_n690), .A2(new_n721), .A3(new_n722), .A4(new_n735), .ZN(new_n736));
  NAND2_X1  g311(.A1(new_n698), .A2(G26), .ZN(new_n737));
  XOR2_X1   g312(.A(new_n737), .B(KEYINPUT28), .Z(new_n738));
  NAND2_X1  g313(.A1(new_n487), .A2(G128), .ZN(new_n739));
  NOR2_X1   g314(.A1(G104), .A2(G2105), .ZN(new_n740));
  XNOR2_X1  g315(.A(new_n740), .B(KEYINPUT94), .ZN(new_n741));
  INV_X1    g316(.A(G116), .ZN(new_n742));
  AOI21_X1  g317(.A(new_n472), .B1(new_n742), .B2(G2105), .ZN(new_n743));
  AOI22_X1  g318(.A1(new_n741), .A2(new_n743), .B1(G140), .B2(new_n481), .ZN(new_n744));
  NAND2_X1  g319(.A1(new_n739), .A2(new_n744), .ZN(new_n745));
  AOI21_X1  g320(.A(new_n738), .B1(new_n745), .B2(G29), .ZN(new_n746));
  XNOR2_X1  g321(.A(new_n746), .B(KEYINPUT95), .ZN(new_n747));
  XNOR2_X1  g322(.A(new_n747), .B(G2067), .ZN(new_n748));
  NAND2_X1  g323(.A1(new_n691), .A2(G4), .ZN(new_n749));
  OAI21_X1  g324(.A(new_n749), .B1(new_n601), .B2(new_n691), .ZN(new_n750));
  NAND2_X1  g325(.A1(new_n750), .A2(G1348), .ZN(new_n751));
  INV_X1    g326(.A(G19), .ZN(new_n752));
  OR3_X1    g327(.A1(new_n752), .A2(KEYINPUT92), .A3(G16), .ZN(new_n753));
  OAI21_X1  g328(.A(KEYINPUT92), .B1(new_n752), .B2(G16), .ZN(new_n754));
  OAI211_X1 g329(.A(new_n753), .B(new_n754), .C1(new_n555), .C2(new_n691), .ZN(new_n755));
  XOR2_X1   g330(.A(new_n755), .B(KEYINPUT93), .Z(new_n756));
  OAI211_X1 g331(.A(new_n748), .B(new_n751), .C1(G1341), .C2(new_n756), .ZN(new_n757));
  XNOR2_X1  g332(.A(KEYINPUT27), .B(G1996), .ZN(new_n758));
  XNOR2_X1  g333(.A(new_n758), .B(KEYINPUT99), .ZN(new_n759));
  AND2_X1   g334(.A1(new_n698), .A2(G32), .ZN(new_n760));
  NAND2_X1  g335(.A1(new_n481), .A2(G141), .ZN(new_n761));
  XNOR2_X1  g336(.A(new_n761), .B(KEYINPUT97), .ZN(new_n762));
  NAND3_X1  g337(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n763));
  INV_X1    g338(.A(KEYINPUT26), .ZN(new_n764));
  OR2_X1    g339(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  NAND2_X1  g340(.A1(new_n763), .A2(new_n764), .ZN(new_n766));
  AOI22_X1  g341(.A1(new_n765), .A2(new_n766), .B1(G105), .B2(new_n473), .ZN(new_n767));
  INV_X1    g342(.A(G129), .ZN(new_n768));
  XNOR2_X1  g343(.A(new_n486), .B(KEYINPUT69), .ZN(new_n769));
  OAI211_X1 g344(.A(new_n762), .B(new_n767), .C1(new_n768), .C2(new_n769), .ZN(new_n770));
  INV_X1    g345(.A(KEYINPUT98), .ZN(new_n771));
  OR2_X1    g346(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  NAND2_X1  g347(.A1(new_n770), .A2(new_n771), .ZN(new_n773));
  NAND2_X1  g348(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  AOI21_X1  g349(.A(new_n760), .B1(new_n774), .B2(G29), .ZN(new_n775));
  AOI22_X1  g350(.A1(new_n756), .A2(G1341), .B1(new_n759), .B2(new_n775), .ZN(new_n776));
  OAI221_X1 g351(.A(new_n776), .B1(G1348), .B2(new_n750), .C1(new_n759), .C2(new_n775), .ZN(new_n777));
  NOR3_X1   g352(.A1(new_n736), .A2(new_n757), .A3(new_n777), .ZN(new_n778));
  INV_X1    g353(.A(new_n778), .ZN(new_n779));
  INV_X1    g354(.A(KEYINPUT36), .ZN(new_n780));
  MUX2_X1   g355(.A(G6), .B(G305), .S(G16), .Z(new_n781));
  XNOR2_X1  g356(.A(new_n781), .B(KEYINPUT32), .ZN(new_n782));
  INV_X1    g357(.A(G1981), .ZN(new_n783));
  XNOR2_X1  g358(.A(new_n782), .B(new_n783), .ZN(new_n784));
  NAND2_X1  g359(.A1(new_n691), .A2(G22), .ZN(new_n785));
  OAI21_X1  g360(.A(new_n785), .B1(G166), .B2(new_n691), .ZN(new_n786));
  XOR2_X1   g361(.A(new_n786), .B(G1971), .Z(new_n787));
  OR2_X1    g362(.A1(new_n787), .A2(KEYINPUT90), .ZN(new_n788));
  NAND2_X1  g363(.A1(new_n691), .A2(G23), .ZN(new_n789));
  AND2_X1   g364(.A1(new_n577), .A2(new_n578), .ZN(new_n790));
  OAI21_X1  g365(.A(new_n789), .B1(new_n790), .B2(new_n691), .ZN(new_n791));
  XOR2_X1   g366(.A(KEYINPUT33), .B(G1976), .Z(new_n792));
  XNOR2_X1  g367(.A(new_n791), .B(new_n792), .ZN(new_n793));
  AOI21_X1  g368(.A(new_n793), .B1(new_n787), .B2(KEYINPUT90), .ZN(new_n794));
  NAND3_X1  g369(.A1(new_n784), .A2(new_n788), .A3(new_n794), .ZN(new_n795));
  OR2_X1    g370(.A1(new_n795), .A2(KEYINPUT91), .ZN(new_n796));
  NAND2_X1  g371(.A1(new_n795), .A2(KEYINPUT91), .ZN(new_n797));
  AOI21_X1  g372(.A(KEYINPUT34), .B1(new_n796), .B2(new_n797), .ZN(new_n798));
  NAND2_X1  g373(.A1(new_n481), .A2(G131), .ZN(new_n799));
  NOR2_X1   g374(.A1(new_n465), .A2(G107), .ZN(new_n800));
  OAI21_X1  g375(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n801));
  INV_X1    g376(.A(G119), .ZN(new_n802));
  OAI221_X1 g377(.A(new_n799), .B1(new_n800), .B2(new_n801), .C1(new_n769), .C2(new_n802), .ZN(new_n803));
  MUX2_X1   g378(.A(G25), .B(new_n803), .S(G29), .Z(new_n804));
  XOR2_X1   g379(.A(KEYINPUT35), .B(G1991), .Z(new_n805));
  INV_X1    g380(.A(new_n805), .ZN(new_n806));
  XNOR2_X1  g381(.A(new_n804), .B(new_n806), .ZN(new_n807));
  MUX2_X1   g382(.A(G24), .B(G290), .S(G16), .Z(new_n808));
  XNOR2_X1  g383(.A(new_n808), .B(G1986), .ZN(new_n809));
  NOR2_X1   g384(.A1(new_n807), .A2(new_n809), .ZN(new_n810));
  INV_X1    g385(.A(new_n810), .ZN(new_n811));
  NOR2_X1   g386(.A1(new_n798), .A2(new_n811), .ZN(new_n812));
  NAND3_X1  g387(.A1(new_n796), .A2(new_n797), .A3(KEYINPUT34), .ZN(new_n813));
  AOI21_X1  g388(.A(new_n780), .B1(new_n812), .B2(new_n813), .ZN(new_n814));
  INV_X1    g389(.A(new_n814), .ZN(new_n815));
  NAND3_X1  g390(.A1(new_n812), .A2(new_n780), .A3(new_n813), .ZN(new_n816));
  AOI21_X1  g391(.A(new_n779), .B1(new_n815), .B2(new_n816), .ZN(G311));
  INV_X1    g392(.A(new_n816), .ZN(new_n818));
  OAI21_X1  g393(.A(new_n778), .B1(new_n818), .B2(new_n814), .ZN(G150));
  NAND2_X1  g394(.A1(new_n601), .A2(G559), .ZN(new_n820));
  XNOR2_X1  g395(.A(new_n820), .B(KEYINPUT38), .ZN(new_n821));
  NAND2_X1  g396(.A1(G80), .A2(G543), .ZN(new_n822));
  INV_X1    g397(.A(G67), .ZN(new_n823));
  OAI21_X1  g398(.A(new_n822), .B1(new_n537), .B2(new_n823), .ZN(new_n824));
  AOI22_X1  g399(.A1(new_n824), .A2(G651), .B1(G93), .B2(new_n533), .ZN(new_n825));
  NAND2_X1  g400(.A1(new_n515), .A2(G55), .ZN(new_n826));
  NAND2_X1  g401(.A1(new_n825), .A2(new_n826), .ZN(new_n827));
  NAND2_X1  g402(.A1(new_n554), .A2(new_n827), .ZN(new_n828));
  NAND4_X1  g403(.A1(new_n551), .A2(new_n553), .A3(new_n826), .A4(new_n825), .ZN(new_n829));
  NAND2_X1  g404(.A1(new_n828), .A2(new_n829), .ZN(new_n830));
  XNOR2_X1  g405(.A(new_n821), .B(new_n830), .ZN(new_n831));
  INV_X1    g406(.A(KEYINPUT39), .ZN(new_n832));
  AOI21_X1  g407(.A(G860), .B1(new_n831), .B2(new_n832), .ZN(new_n833));
  OAI21_X1  g408(.A(new_n833), .B1(new_n832), .B2(new_n831), .ZN(new_n834));
  NAND2_X1  g409(.A1(new_n827), .A2(G860), .ZN(new_n835));
  XOR2_X1   g410(.A(new_n835), .B(KEYINPUT37), .Z(new_n836));
  NAND2_X1  g411(.A1(new_n834), .A2(new_n836), .ZN(G145));
  XNOR2_X1  g412(.A(G162), .B(new_n477), .ZN(new_n838));
  XNOR2_X1  g413(.A(new_n838), .B(new_n627), .ZN(new_n839));
  INV_X1    g414(.A(new_n839), .ZN(new_n840));
  XNOR2_X1  g415(.A(new_n717), .B(new_n508), .ZN(new_n841));
  OAI21_X1  g416(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n842));
  INV_X1    g417(.A(G118), .ZN(new_n843));
  AOI21_X1  g418(.A(new_n842), .B1(new_n843), .B2(G2105), .ZN(new_n844));
  AOI21_X1  g419(.A(new_n844), .B1(new_n481), .B2(G142), .ZN(new_n845));
  INV_X1    g420(.A(G130), .ZN(new_n846));
  OAI21_X1  g421(.A(new_n845), .B1(new_n769), .B2(new_n846), .ZN(new_n847));
  XNOR2_X1  g422(.A(new_n847), .B(new_n616), .ZN(new_n848));
  XNOR2_X1  g423(.A(new_n848), .B(new_n803), .ZN(new_n849));
  XNOR2_X1  g424(.A(new_n841), .B(new_n849), .ZN(new_n850));
  XNOR2_X1  g425(.A(new_n774), .B(new_n745), .ZN(new_n851));
  XNOR2_X1  g426(.A(KEYINPUT100), .B(KEYINPUT101), .ZN(new_n852));
  OR2_X1    g427(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n851), .A2(new_n852), .ZN(new_n854));
  NAND3_X1  g429(.A1(new_n850), .A2(new_n853), .A3(new_n854), .ZN(new_n855));
  INV_X1    g430(.A(new_n855), .ZN(new_n856));
  AOI21_X1  g431(.A(new_n850), .B1(new_n853), .B2(new_n854), .ZN(new_n857));
  OAI21_X1  g432(.A(new_n840), .B1(new_n856), .B2(new_n857), .ZN(new_n858));
  INV_X1    g433(.A(G37), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n853), .A2(new_n854), .ZN(new_n860));
  XOR2_X1   g435(.A(new_n841), .B(new_n849), .Z(new_n861));
  NAND2_X1  g436(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  NAND3_X1  g437(.A1(new_n862), .A2(new_n839), .A3(new_n855), .ZN(new_n863));
  NAND3_X1  g438(.A1(new_n858), .A2(new_n859), .A3(new_n863), .ZN(new_n864));
  XNOR2_X1  g439(.A(new_n864), .B(KEYINPUT40), .ZN(G395));
  XOR2_X1   g440(.A(new_n830), .B(KEYINPUT102), .Z(new_n866));
  XNOR2_X1  g441(.A(new_n612), .B(new_n866), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n600), .A2(new_n605), .ZN(new_n868));
  NAND3_X1  g443(.A1(G299), .A2(new_n595), .A3(new_n599), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  INV_X1    g445(.A(KEYINPUT41), .ZN(new_n871));
  XNOR2_X1  g446(.A(new_n870), .B(new_n871), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n867), .A2(new_n872), .ZN(new_n873));
  XOR2_X1   g448(.A(G166), .B(G305), .Z(new_n874));
  OR2_X1    g449(.A1(G288), .A2(G290), .ZN(new_n875));
  INV_X1    g450(.A(KEYINPUT103), .ZN(new_n876));
  NAND2_X1  g451(.A1(G288), .A2(G290), .ZN(new_n877));
  NAND3_X1  g452(.A1(new_n875), .A2(new_n876), .A3(new_n877), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n874), .A2(new_n878), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n875), .A2(new_n877), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n880), .A2(KEYINPUT103), .ZN(new_n881));
  MUX2_X1   g456(.A(new_n874), .B(new_n879), .S(new_n881), .Z(new_n882));
  XNOR2_X1  g457(.A(new_n882), .B(KEYINPUT42), .ZN(new_n883));
  OR2_X1    g458(.A1(new_n612), .A2(new_n866), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n612), .A2(new_n866), .ZN(new_n885));
  NAND3_X1  g460(.A1(new_n884), .A2(new_n885), .A3(new_n870), .ZN(new_n886));
  AND3_X1   g461(.A1(new_n873), .A2(new_n883), .A3(new_n886), .ZN(new_n887));
  AOI21_X1  g462(.A(new_n883), .B1(new_n873), .B2(new_n886), .ZN(new_n888));
  OAI21_X1  g463(.A(G868), .B1(new_n887), .B2(new_n888), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n827), .A2(new_n592), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n889), .A2(new_n890), .ZN(G295));
  NAND2_X1  g466(.A1(new_n889), .A2(new_n890), .ZN(G331));
  INV_X1    g467(.A(KEYINPUT44), .ZN(new_n893));
  INV_X1    g468(.A(KEYINPUT43), .ZN(new_n894));
  INV_X1    g469(.A(KEYINPUT106), .ZN(new_n895));
  NAND2_X1  g470(.A1(G301), .A2(KEYINPUT104), .ZN(new_n896));
  INV_X1    g471(.A(KEYINPUT104), .ZN(new_n897));
  NAND4_X1  g472(.A1(new_n540), .A2(new_n897), .A3(new_n541), .A4(new_n542), .ZN(new_n898));
  AND3_X1   g473(.A1(new_n896), .A2(G168), .A3(new_n898), .ZN(new_n899));
  AOI21_X1  g474(.A(G168), .B1(new_n896), .B2(new_n898), .ZN(new_n900));
  OAI21_X1  g475(.A(new_n830), .B1(new_n899), .B2(new_n900), .ZN(new_n901));
  INV_X1    g476(.A(new_n901), .ZN(new_n902));
  NOR3_X1   g477(.A1(new_n830), .A2(new_n899), .A3(new_n900), .ZN(new_n903));
  NOR2_X1   g478(.A1(new_n870), .A2(new_n871), .ZN(new_n904));
  AOI21_X1  g479(.A(KEYINPUT41), .B1(new_n868), .B2(new_n869), .ZN(new_n905));
  OAI22_X1  g480(.A1(new_n902), .A2(new_n903), .B1(new_n904), .B2(new_n905), .ZN(new_n906));
  INV_X1    g481(.A(KEYINPUT105), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n901), .A2(new_n907), .ZN(new_n908));
  NOR2_X1   g483(.A1(new_n899), .A2(new_n900), .ZN(new_n909));
  INV_X1    g484(.A(new_n830), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  OAI211_X1 g486(.A(new_n830), .B(KEYINPUT105), .C1(new_n899), .C2(new_n900), .ZN(new_n912));
  NAND4_X1  g487(.A1(new_n908), .A2(new_n911), .A3(new_n870), .A4(new_n912), .ZN(new_n913));
  AND2_X1   g488(.A1(new_n906), .A2(new_n913), .ZN(new_n914));
  OAI211_X1 g489(.A(new_n895), .B(new_n859), .C1(new_n914), .C2(new_n882), .ZN(new_n915));
  NAND3_X1  g490(.A1(new_n882), .A2(new_n906), .A3(new_n913), .ZN(new_n916));
  AND2_X1   g491(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  AOI21_X1  g492(.A(new_n882), .B1(new_n906), .B2(new_n913), .ZN(new_n918));
  OAI21_X1  g493(.A(KEYINPUT106), .B1(new_n918), .B2(G37), .ZN(new_n919));
  AOI21_X1  g494(.A(new_n894), .B1(new_n917), .B2(new_n919), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n916), .A2(new_n859), .ZN(new_n921));
  INV_X1    g496(.A(new_n921), .ZN(new_n922));
  NAND3_X1  g497(.A1(new_n908), .A2(new_n911), .A3(new_n912), .ZN(new_n923));
  AND3_X1   g498(.A1(new_n923), .A2(KEYINPUT107), .A3(new_n872), .ZN(new_n924));
  AOI21_X1  g499(.A(KEYINPUT107), .B1(new_n923), .B2(new_n872), .ZN(new_n925));
  AND3_X1   g500(.A1(new_n911), .A2(new_n870), .A3(new_n901), .ZN(new_n926));
  NOR3_X1   g501(.A1(new_n924), .A2(new_n925), .A3(new_n926), .ZN(new_n927));
  OAI21_X1  g502(.A(new_n922), .B1(new_n927), .B2(new_n882), .ZN(new_n928));
  NOR2_X1   g503(.A1(new_n928), .A2(KEYINPUT43), .ZN(new_n929));
  OAI21_X1  g504(.A(new_n893), .B1(new_n920), .B2(new_n929), .ZN(new_n930));
  INV_X1    g505(.A(KEYINPUT108), .ZN(new_n931));
  AOI21_X1  g506(.A(new_n893), .B1(new_n928), .B2(KEYINPUT43), .ZN(new_n932));
  NAND4_X1  g507(.A1(new_n915), .A2(new_n919), .A3(new_n894), .A4(new_n916), .ZN(new_n933));
  AOI21_X1  g508(.A(new_n931), .B1(new_n932), .B2(new_n933), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n923), .A2(new_n872), .ZN(new_n935));
  INV_X1    g510(.A(KEYINPUT107), .ZN(new_n936));
  AOI21_X1  g511(.A(new_n926), .B1(new_n935), .B2(new_n936), .ZN(new_n937));
  NAND3_X1  g512(.A1(new_n923), .A2(KEYINPUT107), .A3(new_n872), .ZN(new_n938));
  AOI21_X1  g513(.A(new_n882), .B1(new_n937), .B2(new_n938), .ZN(new_n939));
  OAI21_X1  g514(.A(KEYINPUT43), .B1(new_n939), .B2(new_n921), .ZN(new_n940));
  AND4_X1   g515(.A1(new_n931), .A2(new_n940), .A3(new_n933), .A4(KEYINPUT44), .ZN(new_n941));
  OAI21_X1  g516(.A(new_n930), .B1(new_n934), .B2(new_n941), .ZN(G397));
  INV_X1    g517(.A(KEYINPUT45), .ZN(new_n943));
  AOI21_X1  g518(.A(new_n496), .B1(new_n466), .B2(new_n491), .ZN(new_n944));
  AOI21_X1  g519(.A(new_n506), .B1(new_n499), .B2(new_n944), .ZN(new_n945));
  AOI21_X1  g520(.A(G1384), .B1(new_n945), .B2(new_n498), .ZN(new_n946));
  INV_X1    g521(.A(KEYINPUT109), .ZN(new_n947));
  OAI21_X1  g522(.A(new_n943), .B1(new_n946), .B2(new_n947), .ZN(new_n948));
  INV_X1    g523(.A(G1384), .ZN(new_n949));
  AND3_X1   g524(.A1(new_n495), .A2(KEYINPUT4), .A3(new_n497), .ZN(new_n950));
  NAND3_X1  g525(.A1(new_n500), .A2(new_n505), .A3(new_n501), .ZN(new_n951));
  OAI21_X1  g526(.A(new_n949), .B1(new_n950), .B2(new_n951), .ZN(new_n952));
  NOR2_X1   g527(.A1(new_n952), .A2(KEYINPUT109), .ZN(new_n953));
  NAND3_X1  g528(.A1(new_n470), .A2(new_n476), .A3(G40), .ZN(new_n954));
  NOR3_X1   g529(.A1(new_n948), .A2(new_n953), .A3(new_n954), .ZN(new_n955));
  INV_X1    g530(.A(new_n955), .ZN(new_n956));
  OR2_X1    g531(.A1(new_n745), .A2(G2067), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n745), .A2(G2067), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n957), .A2(new_n958), .ZN(new_n959));
  INV_X1    g534(.A(new_n959), .ZN(new_n960));
  XNOR2_X1  g535(.A(new_n803), .B(new_n805), .ZN(new_n961));
  INV_X1    g536(.A(G1996), .ZN(new_n962));
  NOR2_X1   g537(.A1(new_n774), .A2(new_n962), .ZN(new_n963));
  AOI21_X1  g538(.A(G1996), .B1(new_n772), .B2(new_n773), .ZN(new_n964));
  OAI211_X1 g539(.A(new_n960), .B(new_n961), .C1(new_n963), .C2(new_n964), .ZN(new_n965));
  INV_X1    g540(.A(new_n965), .ZN(new_n966));
  XOR2_X1   g541(.A(G290), .B(G1986), .Z(new_n967));
  AOI21_X1  g542(.A(new_n956), .B1(new_n966), .B2(new_n967), .ZN(new_n968));
  INV_X1    g543(.A(G40), .ZN(new_n969));
  NOR3_X1   g544(.A1(new_n469), .A2(new_n475), .A3(new_n969), .ZN(new_n970));
  NAND3_X1  g545(.A1(new_n970), .A2(new_n949), .A3(new_n508), .ZN(new_n971));
  NAND3_X1  g546(.A1(new_n577), .A2(G1976), .A3(new_n578), .ZN(new_n972));
  NAND3_X1  g547(.A1(new_n971), .A2(G8), .A3(new_n972), .ZN(new_n973));
  NOR2_X1   g548(.A1(new_n790), .A2(G1976), .ZN(new_n974));
  OR3_X1    g549(.A1(new_n973), .A2(KEYINPUT52), .A3(new_n974), .ZN(new_n975));
  INV_X1    g550(.A(G86), .ZN(new_n976));
  OAI21_X1  g551(.A(new_n585), .B1(new_n522), .B2(new_n976), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n521), .A2(G61), .ZN(new_n978));
  INV_X1    g553(.A(KEYINPUT77), .ZN(new_n979));
  XNOR2_X1  g554(.A(new_n580), .B(new_n979), .ZN(new_n980));
  AOI21_X1  g555(.A(new_n525), .B1(new_n978), .B2(new_n980), .ZN(new_n981));
  OAI21_X1  g556(.A(G1981), .B1(new_n977), .B2(new_n981), .ZN(new_n982));
  INV_X1    g557(.A(KEYINPUT113), .ZN(new_n983));
  NAND4_X1  g558(.A1(new_n584), .A2(new_n586), .A3(new_n783), .A4(new_n585), .ZN(new_n984));
  NAND3_X1  g559(.A1(new_n982), .A2(new_n983), .A3(new_n984), .ZN(new_n985));
  NAND3_X1  g560(.A1(G305), .A2(KEYINPUT113), .A3(G1981), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n985), .A2(new_n986), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n987), .A2(KEYINPUT49), .ZN(new_n988));
  INV_X1    g563(.A(G8), .ZN(new_n989));
  AOI21_X1  g564(.A(new_n989), .B1(new_n946), .B2(new_n970), .ZN(new_n990));
  INV_X1    g565(.A(KEYINPUT49), .ZN(new_n991));
  NAND3_X1  g566(.A1(new_n985), .A2(new_n991), .A3(new_n986), .ZN(new_n992));
  NAND3_X1  g567(.A1(new_n988), .A2(new_n990), .A3(new_n992), .ZN(new_n993));
  AOI21_X1  g568(.A(KEYINPUT112), .B1(new_n973), .B2(KEYINPUT52), .ZN(new_n994));
  AND3_X1   g569(.A1(new_n973), .A2(KEYINPUT112), .A3(KEYINPUT52), .ZN(new_n995));
  OAI211_X1 g570(.A(new_n975), .B(new_n993), .C1(new_n994), .C2(new_n995), .ZN(new_n996));
  NOR2_X1   g571(.A1(KEYINPUT50), .A2(G1384), .ZN(new_n997));
  OAI21_X1  g572(.A(new_n997), .B1(new_n950), .B2(new_n951), .ZN(new_n998));
  INV_X1    g573(.A(KEYINPUT111), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n998), .A2(new_n999), .ZN(new_n1000));
  NAND3_X1  g575(.A1(new_n508), .A2(KEYINPUT111), .A3(new_n997), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n1000), .A2(new_n1001), .ZN(new_n1002));
  AOI21_X1  g577(.A(new_n954), .B1(new_n952), .B2(KEYINPUT50), .ZN(new_n1003));
  NAND3_X1  g578(.A1(new_n1002), .A2(new_n689), .A3(new_n1003), .ZN(new_n1004));
  XNOR2_X1  g579(.A(KEYINPUT110), .B(G1971), .ZN(new_n1005));
  INV_X1    g580(.A(new_n1005), .ZN(new_n1006));
  OAI21_X1  g581(.A(new_n970), .B1(new_n946), .B2(KEYINPUT45), .ZN(new_n1007));
  NAND3_X1  g582(.A1(new_n508), .A2(KEYINPUT45), .A3(new_n949), .ZN(new_n1008));
  INV_X1    g583(.A(new_n1008), .ZN(new_n1009));
  OAI21_X1  g584(.A(new_n1006), .B1(new_n1007), .B2(new_n1009), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n1004), .A2(new_n1010), .ZN(new_n1011));
  NAND3_X1  g586(.A1(G303), .A2(KEYINPUT55), .A3(G8), .ZN(new_n1012));
  INV_X1    g587(.A(new_n1012), .ZN(new_n1013));
  AOI21_X1  g588(.A(KEYINPUT55), .B1(G303), .B2(G8), .ZN(new_n1014));
  OR2_X1    g589(.A1(new_n1013), .A2(new_n1014), .ZN(new_n1015));
  NAND3_X1  g590(.A1(new_n1011), .A2(new_n1015), .A3(G8), .ZN(new_n1016));
  XOR2_X1   g591(.A(new_n984), .B(KEYINPUT114), .Z(new_n1017));
  NOR2_X1   g592(.A1(G288), .A2(G1976), .ZN(new_n1018));
  XNOR2_X1  g593(.A(new_n1018), .B(KEYINPUT115), .ZN(new_n1019));
  AOI21_X1  g594(.A(new_n1017), .B1(new_n993), .B2(new_n1019), .ZN(new_n1020));
  INV_X1    g595(.A(new_n990), .ZN(new_n1021));
  OAI22_X1  g596(.A1(new_n996), .A2(new_n1016), .B1(new_n1020), .B2(new_n1021), .ZN(new_n1022));
  INV_X1    g597(.A(KEYINPUT63), .ZN(new_n1023));
  INV_X1    g598(.A(KEYINPUT50), .ZN(new_n1024));
  OAI211_X1 g599(.A(new_n970), .B(new_n998), .C1(new_n946), .C2(new_n1024), .ZN(new_n1025));
  NOR2_X1   g600(.A1(new_n1025), .A2(G2090), .ZN(new_n1026));
  AOI21_X1  g601(.A(new_n954), .B1(new_n952), .B2(new_n943), .ZN(new_n1027));
  AOI21_X1  g602(.A(new_n1005), .B1(new_n1027), .B2(new_n1008), .ZN(new_n1028));
  OAI21_X1  g603(.A(G8), .B1(new_n1026), .B2(new_n1028), .ZN(new_n1029));
  NOR2_X1   g604(.A1(new_n1013), .A2(new_n1014), .ZN(new_n1030));
  NAND2_X1  g605(.A1(new_n1029), .A2(new_n1030), .ZN(new_n1031));
  NOR3_X1   g606(.A1(new_n973), .A2(KEYINPUT52), .A3(new_n974), .ZN(new_n1032));
  AND2_X1   g607(.A1(new_n992), .A2(new_n990), .ZN(new_n1033));
  AOI21_X1  g608(.A(new_n1032), .B1(new_n1033), .B2(new_n988), .ZN(new_n1034));
  INV_X1    g609(.A(new_n994), .ZN(new_n1035));
  NAND3_X1  g610(.A1(new_n973), .A2(KEYINPUT112), .A3(KEYINPUT52), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n1035), .A2(new_n1036), .ZN(new_n1037));
  NAND4_X1  g612(.A1(new_n1031), .A2(new_n1016), .A3(new_n1034), .A4(new_n1037), .ZN(new_n1038));
  INV_X1    g613(.A(G2084), .ZN(new_n1039));
  AOI21_X1  g614(.A(KEYINPUT111), .B1(new_n508), .B2(new_n997), .ZN(new_n1040));
  INV_X1    g615(.A(new_n997), .ZN(new_n1041));
  AOI211_X1 g616(.A(new_n999), .B(new_n1041), .C1(new_n945), .C2(new_n498), .ZN(new_n1042));
  OAI211_X1 g617(.A(new_n1003), .B(new_n1039), .C1(new_n1040), .C2(new_n1042), .ZN(new_n1043));
  INV_X1    g618(.A(G1966), .ZN(new_n1044));
  OAI21_X1  g619(.A(new_n1044), .B1(new_n1007), .B2(new_n1009), .ZN(new_n1045));
  NAND2_X1  g620(.A1(new_n1043), .A2(new_n1045), .ZN(new_n1046));
  NAND2_X1  g621(.A1(G168), .A2(G8), .ZN(new_n1047));
  INV_X1    g622(.A(new_n1047), .ZN(new_n1048));
  AOI21_X1  g623(.A(KEYINPUT116), .B1(new_n1046), .B2(new_n1048), .ZN(new_n1049));
  INV_X1    g624(.A(KEYINPUT116), .ZN(new_n1050));
  AOI211_X1 g625(.A(new_n1050), .B(new_n1047), .C1(new_n1043), .C2(new_n1045), .ZN(new_n1051));
  NOR2_X1   g626(.A1(new_n1049), .A2(new_n1051), .ZN(new_n1052));
  OAI21_X1  g627(.A(new_n1023), .B1(new_n1038), .B2(new_n1052), .ZN(new_n1053));
  AND3_X1   g628(.A1(new_n1016), .A2(new_n1034), .A3(new_n1037), .ZN(new_n1054));
  NAND2_X1  g629(.A1(new_n1046), .A2(new_n1048), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n1055), .A2(new_n1050), .ZN(new_n1056));
  NAND3_X1  g631(.A1(new_n1046), .A2(KEYINPUT116), .A3(new_n1048), .ZN(new_n1057));
  NAND2_X1  g632(.A1(new_n1056), .A2(new_n1057), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n1011), .A2(G8), .ZN(new_n1059));
  AOI21_X1  g634(.A(new_n1023), .B1(new_n1059), .B2(new_n1030), .ZN(new_n1060));
  NAND3_X1  g635(.A1(new_n1054), .A2(new_n1058), .A3(new_n1060), .ZN(new_n1061));
  AOI21_X1  g636(.A(new_n1022), .B1(new_n1053), .B2(new_n1061), .ZN(new_n1062));
  NAND3_X1  g637(.A1(new_n1043), .A2(new_n1045), .A3(G168), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n1063), .A2(G8), .ZN(new_n1064));
  AOI21_X1  g639(.A(G168), .B1(new_n1043), .B2(new_n1045), .ZN(new_n1065));
  OAI21_X1  g640(.A(KEYINPUT51), .B1(new_n1064), .B2(new_n1065), .ZN(new_n1066));
  INV_X1    g641(.A(KEYINPUT51), .ZN(new_n1067));
  NAND3_X1  g642(.A1(new_n1063), .A2(new_n1067), .A3(G8), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n1066), .A2(new_n1068), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n1069), .A2(KEYINPUT62), .ZN(new_n1070));
  INV_X1    g645(.A(KEYINPUT62), .ZN(new_n1071));
  NAND3_X1  g646(.A1(new_n1066), .A2(new_n1071), .A3(new_n1068), .ZN(new_n1072));
  OAI21_X1  g647(.A(new_n1003), .B1(new_n1040), .B2(new_n1042), .ZN(new_n1073));
  INV_X1    g648(.A(G1961), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n952), .A2(new_n943), .ZN(new_n1075));
  NAND4_X1  g650(.A1(new_n1075), .A2(new_n732), .A3(new_n970), .A4(new_n1008), .ZN(new_n1076));
  INV_X1    g651(.A(KEYINPUT53), .ZN(new_n1077));
  AOI22_X1  g652(.A1(new_n1073), .A2(new_n1074), .B1(new_n1076), .B2(new_n1077), .ZN(new_n1078));
  NOR3_X1   g653(.A1(new_n954), .A2(new_n1077), .A3(G2078), .ZN(new_n1079));
  NAND3_X1  g654(.A1(new_n1079), .A2(new_n1075), .A3(new_n1008), .ZN(new_n1080));
  AOI21_X1  g655(.A(G301), .B1(new_n1078), .B2(new_n1080), .ZN(new_n1081));
  INV_X1    g656(.A(new_n1081), .ZN(new_n1082));
  NOR2_X1   g657(.A1(new_n1038), .A2(new_n1082), .ZN(new_n1083));
  NAND3_X1  g658(.A1(new_n1070), .A2(new_n1072), .A3(new_n1083), .ZN(new_n1084));
  AND2_X1   g659(.A1(new_n1062), .A2(new_n1084), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n605), .A2(KEYINPUT57), .ZN(new_n1086));
  AND3_X1   g661(.A1(new_n566), .A2(KEYINPUT118), .A3(new_n568), .ZN(new_n1087));
  AOI21_X1  g662(.A(KEYINPUT118), .B1(new_n566), .B2(new_n568), .ZN(new_n1088));
  NOR3_X1   g663(.A1(new_n1087), .A2(new_n1088), .A3(new_n572), .ZN(new_n1089));
  XNOR2_X1  g664(.A(KEYINPUT117), .B(KEYINPUT57), .ZN(new_n1090));
  INV_X1    g665(.A(new_n1090), .ZN(new_n1091));
  OAI21_X1  g666(.A(new_n1086), .B1(new_n1089), .B2(new_n1091), .ZN(new_n1092));
  INV_X1    g667(.A(G1956), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1025), .A2(new_n1093), .ZN(new_n1094));
  XNOR2_X1  g669(.A(KEYINPUT56), .B(G2072), .ZN(new_n1095));
  NAND3_X1  g670(.A1(new_n1027), .A2(new_n1008), .A3(new_n1095), .ZN(new_n1096));
  AND3_X1   g671(.A1(new_n1092), .A2(new_n1094), .A3(new_n1096), .ZN(new_n1097));
  AOI21_X1  g672(.A(new_n1092), .B1(new_n1094), .B2(new_n1096), .ZN(new_n1098));
  OAI211_X1 g673(.A(KEYINPUT122), .B(KEYINPUT61), .C1(new_n1097), .C2(new_n1098), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n1094), .A2(new_n1096), .ZN(new_n1100));
  INV_X1    g675(.A(new_n1092), .ZN(new_n1101));
  NAND3_X1  g676(.A1(new_n1100), .A2(KEYINPUT122), .A3(new_n1101), .ZN(new_n1102));
  INV_X1    g677(.A(KEYINPUT61), .ZN(new_n1103));
  NAND4_X1  g678(.A1(new_n1092), .A2(new_n1094), .A3(new_n1096), .A4(KEYINPUT122), .ZN(new_n1104));
  NAND3_X1  g679(.A1(new_n1102), .A2(new_n1103), .A3(new_n1104), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n1099), .A2(new_n1105), .ZN(new_n1106));
  NOR2_X1   g681(.A1(new_n971), .A2(G2067), .ZN(new_n1107));
  INV_X1    g682(.A(G1348), .ZN(new_n1108));
  AOI21_X1  g683(.A(new_n1107), .B1(new_n1073), .B2(new_n1108), .ZN(new_n1109));
  AOI21_X1  g684(.A(new_n600), .B1(new_n1109), .B2(KEYINPUT60), .ZN(new_n1110));
  AOI21_X1  g685(.A(G1348), .B1(new_n1002), .B2(new_n1003), .ZN(new_n1111));
  INV_X1    g686(.A(KEYINPUT60), .ZN(new_n1112));
  INV_X1    g687(.A(new_n600), .ZN(new_n1113));
  NOR4_X1   g688(.A1(new_n1111), .A2(new_n1112), .A3(new_n1113), .A4(new_n1107), .ZN(new_n1114));
  OAI22_X1  g689(.A1(new_n1110), .A2(new_n1114), .B1(KEYINPUT60), .B2(new_n1109), .ZN(new_n1115));
  AND2_X1   g690(.A1(new_n555), .A2(KEYINPUT121), .ZN(new_n1116));
  NAND3_X1  g691(.A1(new_n1027), .A2(new_n962), .A3(new_n1008), .ZN(new_n1117));
  XOR2_X1   g692(.A(KEYINPUT58), .B(G1341), .Z(new_n1118));
  NAND2_X1  g693(.A1(new_n971), .A2(new_n1118), .ZN(new_n1119));
  AND3_X1   g694(.A1(new_n1117), .A2(KEYINPUT120), .A3(new_n1119), .ZN(new_n1120));
  AOI21_X1  g695(.A(KEYINPUT120), .B1(new_n1117), .B2(new_n1119), .ZN(new_n1121));
  OAI211_X1 g696(.A(KEYINPUT59), .B(new_n1116), .C1(new_n1120), .C2(new_n1121), .ZN(new_n1122));
  OAI21_X1  g697(.A(new_n1116), .B1(new_n1120), .B2(new_n1121), .ZN(new_n1123));
  INV_X1    g698(.A(KEYINPUT59), .ZN(new_n1124));
  NAND2_X1  g699(.A1(new_n1123), .A2(new_n1124), .ZN(new_n1125));
  NAND4_X1  g700(.A1(new_n1106), .A2(new_n1115), .A3(new_n1122), .A4(new_n1125), .ZN(new_n1126));
  NAND2_X1  g701(.A1(new_n1100), .A2(new_n1101), .ZN(new_n1127));
  OAI21_X1  g702(.A(new_n1113), .B1(new_n1111), .B2(new_n1107), .ZN(new_n1128));
  AOI211_X1 g703(.A(KEYINPUT119), .B(new_n1097), .C1(new_n1127), .C2(new_n1128), .ZN(new_n1129));
  INV_X1    g704(.A(KEYINPUT119), .ZN(new_n1130));
  NAND2_X1  g705(.A1(new_n1128), .A2(new_n1127), .ZN(new_n1131));
  INV_X1    g706(.A(new_n1097), .ZN(new_n1132));
  AOI21_X1  g707(.A(new_n1130), .B1(new_n1131), .B2(new_n1132), .ZN(new_n1133));
  NOR2_X1   g708(.A1(new_n1129), .A2(new_n1133), .ZN(new_n1134));
  NAND2_X1  g709(.A1(new_n1126), .A2(new_n1134), .ZN(new_n1135));
  NOR2_X1   g710(.A1(new_n1042), .A2(new_n1040), .ZN(new_n1136));
  OAI21_X1  g711(.A(new_n970), .B1(new_n946), .B2(new_n1024), .ZN(new_n1137));
  OAI21_X1  g712(.A(new_n1074), .B1(new_n1136), .B2(new_n1137), .ZN(new_n1138));
  NAND2_X1  g713(.A1(new_n1076), .A2(new_n1077), .ZN(new_n1139));
  OAI211_X1 g714(.A(new_n1008), .B(new_n1079), .C1(new_n948), .C2(new_n953), .ZN(new_n1140));
  NAND3_X1  g715(.A1(new_n1138), .A2(new_n1139), .A3(new_n1140), .ZN(new_n1141));
  NAND2_X1  g716(.A1(new_n1141), .A2(G171), .ZN(new_n1142));
  INV_X1    g717(.A(KEYINPUT124), .ZN(new_n1143));
  NAND2_X1  g718(.A1(new_n1142), .A2(new_n1143), .ZN(new_n1144));
  NAND4_X1  g719(.A1(new_n1138), .A2(new_n1139), .A3(G301), .A4(new_n1080), .ZN(new_n1145));
  AND2_X1   g720(.A1(new_n1145), .A2(KEYINPUT54), .ZN(new_n1146));
  NAND3_X1  g721(.A1(new_n1141), .A2(KEYINPUT124), .A3(G171), .ZN(new_n1147));
  NAND3_X1  g722(.A1(new_n1144), .A2(new_n1146), .A3(new_n1147), .ZN(new_n1148));
  INV_X1    g723(.A(new_n1038), .ZN(new_n1149));
  AND3_X1   g724(.A1(new_n1148), .A2(new_n1149), .A3(new_n1069), .ZN(new_n1150));
  INV_X1    g725(.A(KEYINPUT54), .ZN(new_n1151));
  NOR2_X1   g726(.A1(new_n1141), .A2(G171), .ZN(new_n1152));
  OAI21_X1  g727(.A(new_n1151), .B1(new_n1152), .B2(new_n1081), .ZN(new_n1153));
  INV_X1    g728(.A(KEYINPUT123), .ZN(new_n1154));
  NAND2_X1  g729(.A1(new_n1153), .A2(new_n1154), .ZN(new_n1155));
  OAI211_X1 g730(.A(KEYINPUT123), .B(new_n1151), .C1(new_n1152), .C2(new_n1081), .ZN(new_n1156));
  NAND2_X1  g731(.A1(new_n1155), .A2(new_n1156), .ZN(new_n1157));
  NAND3_X1  g732(.A1(new_n1135), .A2(new_n1150), .A3(new_n1157), .ZN(new_n1158));
  AOI21_X1  g733(.A(new_n968), .B1(new_n1085), .B2(new_n1158), .ZN(new_n1159));
  NOR2_X1   g734(.A1(new_n803), .A2(new_n806), .ZN(new_n1160));
  OAI211_X1 g735(.A(new_n960), .B(new_n1160), .C1(new_n963), .C2(new_n964), .ZN(new_n1161));
  AOI21_X1  g736(.A(new_n956), .B1(new_n1161), .B2(new_n957), .ZN(new_n1162));
  INV_X1    g737(.A(KEYINPUT126), .ZN(new_n1163));
  NAND3_X1  g738(.A1(new_n965), .A2(new_n1163), .A3(new_n955), .ZN(new_n1164));
  NOR2_X1   g739(.A1(G290), .A2(G1986), .ZN(new_n1165));
  NAND2_X1  g740(.A1(new_n955), .A2(new_n1165), .ZN(new_n1166));
  XNOR2_X1  g741(.A(new_n1166), .B(KEYINPUT48), .ZN(new_n1167));
  AND2_X1   g742(.A1(new_n1164), .A2(new_n1167), .ZN(new_n1168));
  OAI21_X1  g743(.A(KEYINPUT126), .B1(new_n966), .B2(new_n956), .ZN(new_n1169));
  AOI21_X1  g744(.A(new_n1162), .B1(new_n1168), .B2(new_n1169), .ZN(new_n1170));
  NAND2_X1  g745(.A1(new_n955), .A2(new_n962), .ZN(new_n1171));
  XNOR2_X1  g746(.A(new_n1171), .B(KEYINPUT46), .ZN(new_n1172));
  OAI21_X1  g747(.A(new_n955), .B1(new_n774), .B2(new_n959), .ZN(new_n1173));
  NAND2_X1  g748(.A1(new_n1172), .A2(new_n1173), .ZN(new_n1174));
  INV_X1    g749(.A(KEYINPUT47), .ZN(new_n1175));
  NAND2_X1  g750(.A1(new_n1174), .A2(new_n1175), .ZN(new_n1176));
  INV_X1    g751(.A(KEYINPUT125), .ZN(new_n1177));
  NAND3_X1  g752(.A1(new_n1172), .A2(KEYINPUT47), .A3(new_n1173), .ZN(new_n1178));
  NAND3_X1  g753(.A1(new_n1176), .A2(new_n1177), .A3(new_n1178), .ZN(new_n1179));
  NAND2_X1  g754(.A1(new_n1176), .A2(new_n1178), .ZN(new_n1180));
  NAND2_X1  g755(.A1(new_n1180), .A2(KEYINPUT125), .ZN(new_n1181));
  NAND3_X1  g756(.A1(new_n1170), .A2(new_n1179), .A3(new_n1181), .ZN(new_n1182));
  OAI21_X1  g757(.A(KEYINPUT127), .B1(new_n1159), .B2(new_n1182), .ZN(new_n1183));
  INV_X1    g758(.A(new_n968), .ZN(new_n1184));
  AND3_X1   g759(.A1(new_n1135), .A2(new_n1157), .A3(new_n1150), .ZN(new_n1185));
  NAND2_X1  g760(.A1(new_n1062), .A2(new_n1084), .ZN(new_n1186));
  OAI21_X1  g761(.A(new_n1184), .B1(new_n1185), .B2(new_n1186), .ZN(new_n1187));
  INV_X1    g762(.A(KEYINPUT127), .ZN(new_n1188));
  INV_X1    g763(.A(new_n1182), .ZN(new_n1189));
  NAND3_X1  g764(.A1(new_n1187), .A2(new_n1188), .A3(new_n1189), .ZN(new_n1190));
  NAND2_X1  g765(.A1(new_n1183), .A2(new_n1190), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g766(.A1(G227), .A2(new_n463), .ZN(new_n1193));
  OAI21_X1  g767(.A(new_n1193), .B1(new_n682), .B2(new_n683), .ZN(new_n1194));
  NOR2_X1   g768(.A1(G401), .A2(new_n1194), .ZN(new_n1195));
  OAI211_X1 g769(.A(new_n1195), .B(new_n864), .C1(new_n920), .C2(new_n929), .ZN(G225));
  INV_X1    g770(.A(G225), .ZN(G308));
endmodule


