//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 1 1 1 1 0 0 1 0 0 1 1 0 1 0 0 0 0 0 1 0 0 0 0 1 1 1 0 1 1 1 1 0 0 0 1 1 1 1 0 1 1 1 0 0 1 1 1 1 1 0 1 1 1 0 1 0 1 1 0 0 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:23:14 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n608,
    new_n609, new_n611, new_n612, new_n613, new_n614, new_n615, new_n616,
    new_n617, new_n618, new_n620, new_n621, new_n622, new_n623, new_n624,
    new_n625, new_n626, new_n627, new_n628, new_n629, new_n630, new_n631,
    new_n632, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n653, new_n654,
    new_n655, new_n656, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n667, new_n668, new_n669, new_n670,
    new_n672, new_n673, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n712, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n920,
    new_n921, new_n922, new_n923, new_n924, new_n925, new_n926, new_n927,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n945, new_n946, new_n947, new_n948, new_n949, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n978, new_n979, new_n980,
    new_n981, new_n982, new_n983, new_n984, new_n985, new_n986, new_n987,
    new_n988, new_n989, new_n990;
  INV_X1    g000(.A(G237), .ZN(new_n187));
  INV_X1    g001(.A(G953), .ZN(new_n188));
  NAND3_X1  g002(.A1(new_n187), .A2(new_n188), .A3(G214), .ZN(new_n189));
  INV_X1    g003(.A(G143), .ZN(new_n190));
  NOR2_X1   g004(.A1(new_n189), .A2(new_n190), .ZN(new_n191));
  NOR2_X1   g005(.A1(G237), .A2(G953), .ZN(new_n192));
  AOI21_X1  g006(.A(G143), .B1(new_n192), .B2(G214), .ZN(new_n193));
  OAI21_X1  g007(.A(G131), .B1(new_n191), .B2(new_n193), .ZN(new_n194));
  INV_X1    g008(.A(KEYINPUT17), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n189), .A2(new_n190), .ZN(new_n196));
  INV_X1    g010(.A(G131), .ZN(new_n197));
  NAND3_X1  g011(.A1(new_n192), .A2(G143), .A3(G214), .ZN(new_n198));
  NAND3_X1  g012(.A1(new_n196), .A2(new_n197), .A3(new_n198), .ZN(new_n199));
  NAND3_X1  g013(.A1(new_n194), .A2(new_n195), .A3(new_n199), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n200), .A2(KEYINPUT90), .ZN(new_n201));
  INV_X1    g015(.A(KEYINPUT90), .ZN(new_n202));
  NAND4_X1  g016(.A1(new_n194), .A2(new_n202), .A3(new_n195), .A4(new_n199), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n201), .A2(new_n203), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n196), .A2(new_n198), .ZN(new_n205));
  NAND3_X1  g019(.A1(new_n205), .A2(KEYINPUT17), .A3(G131), .ZN(new_n206));
  XNOR2_X1  g020(.A(new_n206), .B(KEYINPUT89), .ZN(new_n207));
  INV_X1    g021(.A(G140), .ZN(new_n208));
  INV_X1    g022(.A(G125), .ZN(new_n209));
  OAI21_X1  g023(.A(new_n208), .B1(new_n209), .B2(KEYINPUT74), .ZN(new_n210));
  INV_X1    g024(.A(KEYINPUT74), .ZN(new_n211));
  NAND3_X1  g025(.A1(new_n211), .A2(G125), .A3(G140), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n210), .A2(new_n212), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n213), .A2(KEYINPUT16), .ZN(new_n214));
  NOR3_X1   g028(.A1(new_n209), .A2(KEYINPUT16), .A3(G140), .ZN(new_n215));
  INV_X1    g029(.A(new_n215), .ZN(new_n216));
  AOI21_X1  g030(.A(G146), .B1(new_n214), .B2(new_n216), .ZN(new_n217));
  INV_X1    g031(.A(KEYINPUT16), .ZN(new_n218));
  AOI21_X1  g032(.A(new_n218), .B1(new_n210), .B2(new_n212), .ZN(new_n219));
  INV_X1    g033(.A(G146), .ZN(new_n220));
  NOR3_X1   g034(.A1(new_n219), .A2(new_n220), .A3(new_n215), .ZN(new_n221));
  NOR2_X1   g035(.A1(new_n217), .A2(new_n221), .ZN(new_n222));
  NAND3_X1  g036(.A1(new_n204), .A2(new_n207), .A3(new_n222), .ZN(new_n223));
  XNOR2_X1  g037(.A(G113), .B(G122), .ZN(new_n224));
  INV_X1    g038(.A(G104), .ZN(new_n225));
  XNOR2_X1  g039(.A(new_n224), .B(new_n225), .ZN(new_n226));
  NAND2_X1  g040(.A1(KEYINPUT18), .A2(G131), .ZN(new_n227));
  OAI21_X1  g041(.A(new_n227), .B1(new_n205), .B2(KEYINPUT87), .ZN(new_n228));
  INV_X1    g042(.A(KEYINPUT87), .ZN(new_n229));
  INV_X1    g043(.A(new_n227), .ZN(new_n230));
  NAND4_X1  g044(.A1(new_n196), .A2(new_n229), .A3(new_n198), .A4(new_n230), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n228), .A2(new_n231), .ZN(new_n232));
  XNOR2_X1  g046(.A(G125), .B(G140), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n233), .A2(new_n220), .ZN(new_n234));
  NAND3_X1  g048(.A1(new_n210), .A2(G146), .A3(new_n212), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n234), .A2(new_n235), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n232), .A2(new_n236), .ZN(new_n237));
  NAND3_X1  g051(.A1(new_n223), .A2(new_n226), .A3(new_n237), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n194), .A2(new_n199), .ZN(new_n239));
  NAND3_X1  g053(.A1(new_n214), .A2(G146), .A3(new_n216), .ZN(new_n240));
  NOR2_X1   g054(.A1(new_n233), .A2(KEYINPUT19), .ZN(new_n241));
  INV_X1    g055(.A(KEYINPUT19), .ZN(new_n242));
  AOI21_X1  g056(.A(new_n242), .B1(new_n210), .B2(new_n212), .ZN(new_n243));
  OAI21_X1  g057(.A(new_n220), .B1(new_n241), .B2(new_n243), .ZN(new_n244));
  AND3_X1   g058(.A1(new_n239), .A2(new_n240), .A3(new_n244), .ZN(new_n245));
  AOI22_X1  g059(.A1(new_n228), .A2(new_n231), .B1(new_n234), .B2(new_n235), .ZN(new_n246));
  OAI21_X1  g060(.A(KEYINPUT88), .B1(new_n245), .B2(new_n246), .ZN(new_n247));
  INV_X1    g061(.A(new_n226), .ZN(new_n248));
  NAND3_X1  g062(.A1(new_n239), .A2(new_n240), .A3(new_n244), .ZN(new_n249));
  INV_X1    g063(.A(KEYINPUT88), .ZN(new_n250));
  NAND3_X1  g064(.A1(new_n237), .A2(new_n249), .A3(new_n250), .ZN(new_n251));
  NAND3_X1  g065(.A1(new_n247), .A2(new_n248), .A3(new_n251), .ZN(new_n252));
  AOI21_X1  g066(.A(G475), .B1(new_n238), .B2(new_n252), .ZN(new_n253));
  INV_X1    g067(.A(G902), .ZN(new_n254));
  AND3_X1   g068(.A1(new_n253), .A2(KEYINPUT20), .A3(new_n254), .ZN(new_n255));
  AOI21_X1  g069(.A(KEYINPUT20), .B1(new_n253), .B2(new_n254), .ZN(new_n256));
  NOR2_X1   g070(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  AND3_X1   g071(.A1(new_n223), .A2(new_n226), .A3(new_n237), .ZN(new_n258));
  AOI21_X1  g072(.A(new_n226), .B1(new_n223), .B2(new_n237), .ZN(new_n259));
  OAI21_X1  g073(.A(new_n254), .B1(new_n258), .B2(new_n259), .ZN(new_n260));
  INV_X1    g074(.A(KEYINPUT91), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  OAI211_X1 g076(.A(KEYINPUT91), .B(new_n254), .C1(new_n258), .C2(new_n259), .ZN(new_n263));
  NAND3_X1  g077(.A1(new_n262), .A2(G475), .A3(new_n263), .ZN(new_n264));
  XNOR2_X1  g078(.A(KEYINPUT9), .B(G234), .ZN(new_n265));
  INV_X1    g079(.A(new_n265), .ZN(new_n266));
  NAND3_X1  g080(.A1(new_n266), .A2(G217), .A3(new_n188), .ZN(new_n267));
  INV_X1    g081(.A(G116), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n268), .A2(G122), .ZN(new_n269));
  OAI21_X1  g083(.A(KEYINPUT92), .B1(new_n269), .B2(KEYINPUT14), .ZN(new_n270));
  OR2_X1    g084(.A1(new_n268), .A2(G122), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n269), .A2(KEYINPUT14), .ZN(new_n272));
  INV_X1    g086(.A(KEYINPUT92), .ZN(new_n273));
  INV_X1    g087(.A(KEYINPUT14), .ZN(new_n274));
  NAND4_X1  g088(.A1(new_n273), .A2(new_n274), .A3(new_n268), .A4(G122), .ZN(new_n275));
  NAND4_X1  g089(.A1(new_n270), .A2(new_n271), .A3(new_n272), .A4(new_n275), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n276), .A2(G107), .ZN(new_n277));
  INV_X1    g091(.A(G107), .ZN(new_n278));
  AND3_X1   g092(.A1(new_n271), .A2(new_n269), .A3(new_n278), .ZN(new_n279));
  INV_X1    g093(.A(new_n279), .ZN(new_n280));
  XNOR2_X1  g094(.A(G128), .B(G143), .ZN(new_n281));
  INV_X1    g095(.A(G134), .ZN(new_n282));
  XNOR2_X1  g096(.A(new_n281), .B(new_n282), .ZN(new_n283));
  NAND3_X1  g097(.A1(new_n277), .A2(new_n280), .A3(new_n283), .ZN(new_n284));
  INV_X1    g098(.A(new_n284), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n281), .A2(new_n282), .ZN(new_n286));
  AOI21_X1  g100(.A(new_n278), .B1(new_n271), .B2(new_n269), .ZN(new_n287));
  OAI21_X1  g101(.A(new_n286), .B1(new_n279), .B2(new_n287), .ZN(new_n288));
  INV_X1    g102(.A(G128), .ZN(new_n289));
  NOR3_X1   g103(.A1(new_n289), .A2(KEYINPUT13), .A3(G143), .ZN(new_n290));
  AOI211_X1 g104(.A(new_n282), .B(new_n290), .C1(KEYINPUT13), .C2(new_n281), .ZN(new_n291));
  NOR2_X1   g105(.A1(new_n288), .A2(new_n291), .ZN(new_n292));
  OAI21_X1  g106(.A(new_n267), .B1(new_n285), .B2(new_n292), .ZN(new_n293));
  INV_X1    g107(.A(new_n267), .ZN(new_n294));
  OAI211_X1 g108(.A(new_n284), .B(new_n294), .C1(new_n291), .C2(new_n288), .ZN(new_n295));
  NAND3_X1  g109(.A1(new_n293), .A2(KEYINPUT93), .A3(new_n295), .ZN(new_n296));
  INV_X1    g110(.A(KEYINPUT93), .ZN(new_n297));
  OAI211_X1 g111(.A(new_n297), .B(new_n267), .C1(new_n285), .C2(new_n292), .ZN(new_n298));
  NAND3_X1  g112(.A1(new_n296), .A2(new_n254), .A3(new_n298), .ZN(new_n299));
  INV_X1    g113(.A(G478), .ZN(new_n300));
  NOR2_X1   g114(.A1(new_n300), .A2(KEYINPUT15), .ZN(new_n301));
  XOR2_X1   g115(.A(new_n299), .B(new_n301), .Z(new_n302));
  NAND2_X1  g116(.A1(G234), .A2(G237), .ZN(new_n303));
  NAND3_X1  g117(.A1(new_n303), .A2(G952), .A3(new_n188), .ZN(new_n304));
  INV_X1    g118(.A(new_n304), .ZN(new_n305));
  XOR2_X1   g119(.A(KEYINPUT21), .B(G898), .Z(new_n306));
  INV_X1    g120(.A(new_n306), .ZN(new_n307));
  NAND3_X1  g121(.A1(new_n303), .A2(G902), .A3(G953), .ZN(new_n308));
  INV_X1    g122(.A(new_n308), .ZN(new_n309));
  AOI21_X1  g123(.A(new_n305), .B1(new_n307), .B2(new_n309), .ZN(new_n310));
  INV_X1    g124(.A(new_n310), .ZN(new_n311));
  NAND4_X1  g125(.A1(new_n257), .A2(new_n264), .A3(new_n302), .A4(new_n311), .ZN(new_n312));
  INV_X1    g126(.A(KEYINPUT84), .ZN(new_n313));
  INV_X1    g127(.A(G469), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n188), .A2(G227), .ZN(new_n315));
  XNOR2_X1  g129(.A(new_n315), .B(new_n208), .ZN(new_n316));
  XNOR2_X1  g130(.A(new_n316), .B(KEYINPUT80), .ZN(new_n317));
  XNOR2_X1  g131(.A(new_n317), .B(G110), .ZN(new_n318));
  NOR2_X1   g132(.A1(new_n289), .A2(KEYINPUT1), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n220), .A2(G143), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n190), .A2(G146), .ZN(new_n321));
  NAND3_X1  g135(.A1(new_n319), .A2(new_n320), .A3(new_n321), .ZN(new_n322));
  NAND3_X1  g136(.A1(new_n289), .A2(new_n220), .A3(G143), .ZN(new_n323));
  OAI211_X1 g137(.A(new_n190), .B(G146), .C1(new_n289), .C2(KEYINPUT1), .ZN(new_n324));
  NAND3_X1  g138(.A1(new_n322), .A2(new_n323), .A3(new_n324), .ZN(new_n325));
  INV_X1    g139(.A(KEYINPUT83), .ZN(new_n326));
  OAI21_X1  g140(.A(KEYINPUT81), .B1(new_n278), .B2(G104), .ZN(new_n327));
  INV_X1    g141(.A(KEYINPUT81), .ZN(new_n328));
  NAND3_X1  g142(.A1(new_n328), .A2(new_n225), .A3(G107), .ZN(new_n329));
  AND2_X1   g143(.A1(new_n327), .A2(new_n329), .ZN(new_n330));
  INV_X1    g144(.A(G101), .ZN(new_n331));
  OAI21_X1  g145(.A(KEYINPUT3), .B1(new_n225), .B2(G107), .ZN(new_n332));
  INV_X1    g146(.A(KEYINPUT3), .ZN(new_n333));
  NAND3_X1  g147(.A1(new_n333), .A2(new_n278), .A3(G104), .ZN(new_n334));
  NAND4_X1  g148(.A1(new_n330), .A2(new_n331), .A3(new_n332), .A4(new_n334), .ZN(new_n335));
  NOR2_X1   g149(.A1(new_n225), .A2(G107), .ZN(new_n336));
  NOR2_X1   g150(.A1(new_n278), .A2(G104), .ZN(new_n337));
  OAI21_X1  g151(.A(G101), .B1(new_n336), .B2(new_n337), .ZN(new_n338));
  AOI21_X1  g152(.A(new_n326), .B1(new_n335), .B2(new_n338), .ZN(new_n339));
  NAND4_X1  g153(.A1(new_n332), .A2(new_n327), .A3(new_n334), .A4(new_n329), .ZN(new_n340));
  OAI211_X1 g154(.A(new_n326), .B(new_n338), .C1(new_n340), .C2(G101), .ZN(new_n341));
  INV_X1    g155(.A(new_n341), .ZN(new_n342));
  OAI211_X1 g156(.A(KEYINPUT10), .B(new_n325), .C1(new_n339), .C2(new_n342), .ZN(new_n343));
  INV_X1    g157(.A(KEYINPUT4), .ZN(new_n344));
  NAND3_X1  g158(.A1(new_n340), .A2(new_n344), .A3(G101), .ZN(new_n345));
  INV_X1    g159(.A(KEYINPUT82), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n345), .A2(new_n346), .ZN(new_n347));
  NAND4_X1  g161(.A1(new_n340), .A2(KEYINPUT82), .A3(new_n344), .A4(G101), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n347), .A2(new_n348), .ZN(new_n349));
  INV_X1    g163(.A(KEYINPUT64), .ZN(new_n350));
  XNOR2_X1  g164(.A(G143), .B(G146), .ZN(new_n351));
  XNOR2_X1  g165(.A(KEYINPUT0), .B(G128), .ZN(new_n352));
  OAI21_X1  g166(.A(new_n350), .B1(new_n351), .B2(new_n352), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n320), .A2(new_n321), .ZN(new_n354));
  NAND2_X1  g168(.A1(KEYINPUT0), .A2(G128), .ZN(new_n355));
  OR2_X1    g169(.A1(KEYINPUT0), .A2(G128), .ZN(new_n356));
  NAND4_X1  g170(.A1(new_n354), .A2(KEYINPUT64), .A3(new_n355), .A4(new_n356), .ZN(new_n357));
  NAND3_X1  g171(.A1(new_n351), .A2(KEYINPUT0), .A3(G128), .ZN(new_n358));
  NAND3_X1  g172(.A1(new_n353), .A2(new_n357), .A3(new_n358), .ZN(new_n359));
  INV_X1    g173(.A(new_n359), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n340), .A2(G101), .ZN(new_n361));
  NAND3_X1  g175(.A1(new_n335), .A2(KEYINPUT4), .A3(new_n361), .ZN(new_n362));
  NAND3_X1  g176(.A1(new_n349), .A2(new_n360), .A3(new_n362), .ZN(new_n363));
  OAI211_X1 g177(.A(new_n325), .B(new_n338), .C1(G101), .C2(new_n340), .ZN(new_n364));
  INV_X1    g178(.A(KEYINPUT10), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  NAND3_X1  g180(.A1(new_n343), .A2(new_n363), .A3(new_n366), .ZN(new_n367));
  INV_X1    g181(.A(KEYINPUT11), .ZN(new_n368));
  OAI21_X1  g182(.A(new_n368), .B1(new_n282), .B2(G137), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n282), .A2(G137), .ZN(new_n370));
  INV_X1    g184(.A(G137), .ZN(new_n371));
  NAND3_X1  g185(.A1(new_n371), .A2(KEYINPUT11), .A3(G134), .ZN(new_n372));
  NAND3_X1  g186(.A1(new_n369), .A2(new_n370), .A3(new_n372), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n373), .A2(G131), .ZN(new_n374));
  NAND4_X1  g188(.A1(new_n369), .A2(new_n372), .A3(new_n197), .A4(new_n370), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n367), .A2(new_n376), .ZN(new_n377));
  AND2_X1   g191(.A1(new_n374), .A2(new_n375), .ZN(new_n378));
  NAND4_X1  g192(.A1(new_n343), .A2(new_n363), .A3(new_n378), .A4(new_n366), .ZN(new_n379));
  AOI21_X1  g193(.A(new_n318), .B1(new_n377), .B2(new_n379), .ZN(new_n380));
  OAI21_X1  g194(.A(new_n338), .B1(new_n340), .B2(G101), .ZN(new_n381));
  INV_X1    g195(.A(new_n325), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n381), .A2(new_n382), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n383), .A2(new_n364), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n384), .A2(new_n376), .ZN(new_n385));
  INV_X1    g199(.A(KEYINPUT12), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n385), .A2(new_n386), .ZN(new_n387));
  NAND3_X1  g201(.A1(new_n384), .A2(KEYINPUT12), .A3(new_n376), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n387), .A2(new_n388), .ZN(new_n389));
  AND3_X1   g203(.A1(new_n389), .A2(new_n379), .A3(new_n318), .ZN(new_n390));
  OAI211_X1 g204(.A(new_n314), .B(new_n254), .C1(new_n380), .C2(new_n390), .ZN(new_n391));
  NAND2_X1  g205(.A1(G469), .A2(G902), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n389), .A2(new_n379), .ZN(new_n393));
  INV_X1    g207(.A(new_n318), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n393), .A2(new_n394), .ZN(new_n395));
  NAND3_X1  g209(.A1(new_n377), .A2(new_n379), .A3(new_n318), .ZN(new_n396));
  NAND3_X1  g210(.A1(new_n395), .A2(G469), .A3(new_n396), .ZN(new_n397));
  AND3_X1   g211(.A1(new_n391), .A2(new_n392), .A3(new_n397), .ZN(new_n398));
  OAI21_X1  g212(.A(G221), .B1(new_n265), .B2(G902), .ZN(new_n399));
  XOR2_X1   g213(.A(new_n399), .B(KEYINPUT79), .Z(new_n400));
  INV_X1    g214(.A(new_n400), .ZN(new_n401));
  OAI21_X1  g215(.A(new_n313), .B1(new_n398), .B2(new_n401), .ZN(new_n402));
  NAND3_X1  g216(.A1(new_n391), .A2(new_n392), .A3(new_n397), .ZN(new_n403));
  NAND3_X1  g217(.A1(new_n403), .A2(KEYINPUT84), .A3(new_n400), .ZN(new_n404));
  AOI21_X1  g218(.A(new_n312), .B1(new_n402), .B2(new_n404), .ZN(new_n405));
  INV_X1    g219(.A(new_n370), .ZN(new_n406));
  NOR2_X1   g220(.A1(new_n282), .A2(G137), .ZN(new_n407));
  OAI21_X1  g221(.A(G131), .B1(new_n406), .B2(new_n407), .ZN(new_n408));
  NAND3_X1  g222(.A1(new_n325), .A2(new_n375), .A3(new_n408), .ZN(new_n409));
  OAI21_X1  g223(.A(new_n409), .B1(new_n378), .B2(new_n359), .ZN(new_n410));
  INV_X1    g224(.A(G119), .ZN(new_n411));
  OAI21_X1  g225(.A(KEYINPUT65), .B1(new_n411), .B2(G116), .ZN(new_n412));
  INV_X1    g226(.A(KEYINPUT65), .ZN(new_n413));
  NAND3_X1  g227(.A1(new_n413), .A2(new_n268), .A3(G119), .ZN(new_n414));
  AOI22_X1  g228(.A1(new_n412), .A2(new_n414), .B1(G116), .B2(new_n411), .ZN(new_n415));
  XOR2_X1   g229(.A(KEYINPUT2), .B(G113), .Z(new_n416));
  XNOR2_X1  g230(.A(new_n415), .B(new_n416), .ZN(new_n417));
  NOR2_X1   g231(.A1(new_n410), .A2(new_n417), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n410), .A2(KEYINPUT30), .ZN(new_n419));
  INV_X1    g233(.A(KEYINPUT30), .ZN(new_n420));
  OAI211_X1 g234(.A(new_n420), .B(new_n409), .C1(new_n378), .C2(new_n359), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n419), .A2(new_n421), .ZN(new_n422));
  AOI21_X1  g236(.A(new_n418), .B1(new_n422), .B2(new_n417), .ZN(new_n423));
  XNOR2_X1  g237(.A(KEYINPUT26), .B(G101), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n192), .A2(G210), .ZN(new_n425));
  XNOR2_X1  g239(.A(new_n424), .B(new_n425), .ZN(new_n426));
  XNOR2_X1  g240(.A(KEYINPUT66), .B(KEYINPUT27), .ZN(new_n427));
  AND2_X1   g241(.A1(new_n426), .A2(new_n427), .ZN(new_n428));
  NOR2_X1   g242(.A1(new_n426), .A2(new_n427), .ZN(new_n429));
  NOR2_X1   g243(.A1(new_n428), .A2(new_n429), .ZN(new_n430));
  INV_X1    g244(.A(new_n430), .ZN(new_n431));
  NOR2_X1   g245(.A1(new_n423), .A2(new_n431), .ZN(new_n432));
  OR2_X1    g246(.A1(new_n432), .A2(KEYINPUT72), .ZN(new_n433));
  INV_X1    g247(.A(KEYINPUT28), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n410), .A2(new_n417), .ZN(new_n435));
  NAND4_X1  g249(.A1(new_n376), .A2(new_n357), .A3(new_n358), .A4(new_n353), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n415), .A2(new_n416), .ZN(new_n437));
  INV_X1    g251(.A(new_n437), .ZN(new_n438));
  NOR2_X1   g252(.A1(new_n415), .A2(new_n416), .ZN(new_n439));
  NOR2_X1   g253(.A1(new_n438), .A2(new_n439), .ZN(new_n440));
  NAND3_X1  g254(.A1(new_n436), .A2(new_n440), .A3(new_n409), .ZN(new_n441));
  AOI21_X1  g255(.A(new_n434), .B1(new_n435), .B2(new_n441), .ZN(new_n442));
  NOR2_X1   g256(.A1(new_n418), .A2(KEYINPUT28), .ZN(new_n443));
  NOR2_X1   g257(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n430), .A2(KEYINPUT70), .ZN(new_n445));
  INV_X1    g259(.A(KEYINPUT70), .ZN(new_n446));
  OAI21_X1  g260(.A(new_n446), .B1(new_n428), .B2(new_n429), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n445), .A2(new_n447), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n444), .A2(new_n448), .ZN(new_n449));
  INV_X1    g263(.A(KEYINPUT29), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n432), .A2(KEYINPUT72), .ZN(new_n451));
  NAND4_X1  g265(.A1(new_n433), .A2(new_n449), .A3(new_n450), .A4(new_n451), .ZN(new_n452));
  NOR2_X1   g266(.A1(new_n430), .A2(new_n450), .ZN(new_n453));
  AOI21_X1  g267(.A(G902), .B1(new_n444), .B2(new_n453), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n452), .A2(new_n454), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n455), .A2(G472), .ZN(new_n456));
  INV_X1    g270(.A(KEYINPUT67), .ZN(new_n457));
  AOI21_X1  g271(.A(new_n457), .B1(new_n423), .B2(new_n431), .ZN(new_n458));
  AOI21_X1  g272(.A(new_n440), .B1(new_n419), .B2(new_n421), .ZN(new_n459));
  NOR4_X1   g273(.A1(new_n459), .A2(KEYINPUT67), .A3(new_n418), .A4(new_n430), .ZN(new_n460));
  OAI21_X1  g274(.A(KEYINPUT31), .B1(new_n458), .B2(new_n460), .ZN(new_n461));
  INV_X1    g275(.A(new_n421), .ZN(new_n462));
  AOI21_X1  g276(.A(new_n420), .B1(new_n436), .B2(new_n409), .ZN(new_n463));
  OAI21_X1  g277(.A(new_n417), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  XOR2_X1   g278(.A(KEYINPUT68), .B(KEYINPUT31), .Z(new_n465));
  NAND4_X1  g279(.A1(new_n464), .A2(new_n441), .A3(new_n431), .A4(new_n465), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n466), .A2(KEYINPUT69), .ZN(new_n467));
  INV_X1    g281(.A(KEYINPUT69), .ZN(new_n468));
  NAND4_X1  g282(.A1(new_n423), .A2(new_n468), .A3(new_n431), .A4(new_n465), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n467), .A2(new_n469), .ZN(new_n470));
  INV_X1    g284(.A(new_n448), .ZN(new_n471));
  OAI21_X1  g285(.A(new_n471), .B1(new_n442), .B2(new_n443), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n472), .A2(KEYINPUT71), .ZN(new_n473));
  OR3_X1    g287(.A1(new_n444), .A2(KEYINPUT71), .A3(new_n448), .ZN(new_n474));
  NAND4_X1  g288(.A1(new_n461), .A2(new_n470), .A3(new_n473), .A4(new_n474), .ZN(new_n475));
  INV_X1    g289(.A(KEYINPUT32), .ZN(new_n476));
  NOR2_X1   g290(.A1(G472), .A2(G902), .ZN(new_n477));
  AND3_X1   g291(.A1(new_n475), .A2(new_n476), .A3(new_n477), .ZN(new_n478));
  AOI21_X1  g292(.A(new_n476), .B1(new_n475), .B2(new_n477), .ZN(new_n479));
  OAI21_X1  g293(.A(new_n456), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  NAND3_X1  g294(.A1(new_n188), .A2(G221), .A3(G234), .ZN(new_n481));
  XNOR2_X1  g295(.A(new_n481), .B(KEYINPUT76), .ZN(new_n482));
  XNOR2_X1  g296(.A(new_n482), .B(KEYINPUT22), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n483), .A2(new_n371), .ZN(new_n484));
  OR2_X1    g298(.A1(new_n482), .A2(KEYINPUT22), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n482), .A2(KEYINPUT22), .ZN(new_n486));
  NAND3_X1  g300(.A1(new_n485), .A2(G137), .A3(new_n486), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n484), .A2(new_n487), .ZN(new_n488));
  INV_X1    g302(.A(KEYINPUT23), .ZN(new_n489));
  OAI21_X1  g303(.A(new_n489), .B1(new_n411), .B2(G128), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n411), .A2(G128), .ZN(new_n491));
  NAND3_X1  g305(.A1(new_n289), .A2(KEYINPUT23), .A3(G119), .ZN(new_n492));
  NAND3_X1  g306(.A1(new_n490), .A2(new_n491), .A3(new_n492), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n493), .A2(G110), .ZN(new_n494));
  XOR2_X1   g308(.A(KEYINPUT24), .B(G110), .Z(new_n495));
  XNOR2_X1  g309(.A(G119), .B(G128), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  OAI211_X1 g311(.A(new_n494), .B(new_n497), .C1(new_n217), .C2(new_n221), .ZN(new_n498));
  INV_X1    g312(.A(KEYINPUT75), .ZN(new_n499));
  OAI22_X1  g313(.A1(new_n493), .A2(G110), .B1(new_n495), .B2(new_n496), .ZN(new_n500));
  NAND3_X1  g314(.A1(new_n240), .A2(new_n500), .A3(new_n234), .ZN(new_n501));
  AND3_X1   g315(.A1(new_n498), .A2(new_n499), .A3(new_n501), .ZN(new_n502));
  AOI21_X1  g316(.A(new_n499), .B1(new_n498), .B2(new_n501), .ZN(new_n503));
  OAI21_X1  g317(.A(new_n488), .B1(new_n502), .B2(new_n503), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n504), .A2(KEYINPUT77), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n498), .A2(new_n501), .ZN(new_n506));
  OR2_X1    g320(.A1(new_n488), .A2(new_n506), .ZN(new_n507));
  INV_X1    g321(.A(KEYINPUT77), .ZN(new_n508));
  OAI211_X1 g322(.A(new_n488), .B(new_n508), .C1(new_n502), .C2(new_n503), .ZN(new_n509));
  NAND4_X1  g323(.A1(new_n505), .A2(new_n254), .A3(new_n507), .A4(new_n509), .ZN(new_n510));
  INV_X1    g324(.A(KEYINPUT25), .ZN(new_n511));
  XNOR2_X1  g325(.A(new_n510), .B(new_n511), .ZN(new_n512));
  INV_X1    g326(.A(G234), .ZN(new_n513));
  OAI21_X1  g327(.A(G217), .B1(new_n513), .B2(G902), .ZN(new_n514));
  XNOR2_X1  g328(.A(new_n514), .B(KEYINPUT73), .ZN(new_n515));
  NOR2_X1   g329(.A1(new_n515), .A2(G902), .ZN(new_n516));
  XNOR2_X1  g330(.A(new_n516), .B(KEYINPUT78), .ZN(new_n517));
  NAND3_X1  g331(.A1(new_n505), .A2(new_n507), .A3(new_n509), .ZN(new_n518));
  INV_X1    g332(.A(new_n518), .ZN(new_n519));
  AOI22_X1  g333(.A1(new_n512), .A2(new_n515), .B1(new_n517), .B2(new_n519), .ZN(new_n520));
  OAI21_X1  g334(.A(G214), .B1(G237), .B2(G902), .ZN(new_n521));
  INV_X1    g335(.A(new_n521), .ZN(new_n522));
  NOR3_X1   g336(.A1(new_n268), .A2(KEYINPUT5), .A3(G119), .ZN(new_n523));
  AOI21_X1  g337(.A(new_n523), .B1(new_n415), .B2(KEYINPUT5), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n524), .A2(G113), .ZN(new_n525));
  OAI211_X1 g339(.A(new_n437), .B(new_n525), .C1(new_n339), .C2(new_n342), .ZN(new_n526));
  NAND3_X1  g340(.A1(new_n349), .A2(new_n417), .A3(new_n362), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  XOR2_X1   g342(.A(G110), .B(G122), .Z(new_n529));
  NAND2_X1  g343(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  INV_X1    g344(.A(new_n529), .ZN(new_n531));
  NAND3_X1  g345(.A1(new_n526), .A2(new_n527), .A3(new_n531), .ZN(new_n532));
  NAND3_X1  g346(.A1(new_n530), .A2(KEYINPUT6), .A3(new_n532), .ZN(new_n533));
  INV_X1    g347(.A(KEYINPUT6), .ZN(new_n534));
  NAND3_X1  g348(.A1(new_n528), .A2(new_n534), .A3(new_n529), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n325), .A2(new_n209), .ZN(new_n536));
  OAI21_X1  g350(.A(new_n536), .B1(new_n359), .B2(new_n209), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n188), .A2(G224), .ZN(new_n538));
  XNOR2_X1  g352(.A(new_n537), .B(new_n538), .ZN(new_n539));
  NAND3_X1  g353(.A1(new_n533), .A2(new_n535), .A3(new_n539), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n525), .A2(new_n437), .ZN(new_n541));
  INV_X1    g355(.A(KEYINPUT86), .ZN(new_n542));
  OAI21_X1  g356(.A(new_n542), .B1(new_n381), .B2(KEYINPUT85), .ZN(new_n543));
  OR2_X1    g357(.A1(new_n541), .A2(new_n543), .ZN(new_n544));
  OAI211_X1 g358(.A(new_n541), .B(new_n543), .C1(new_n542), .C2(new_n381), .ZN(new_n545));
  OR2_X1    g359(.A1(new_n529), .A2(KEYINPUT8), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n529), .A2(KEYINPUT8), .ZN(new_n547));
  NAND4_X1  g361(.A1(new_n544), .A2(new_n545), .A3(new_n546), .A4(new_n547), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n538), .A2(KEYINPUT7), .ZN(new_n549));
  XNOR2_X1  g363(.A(new_n537), .B(new_n549), .ZN(new_n550));
  NAND3_X1  g364(.A1(new_n548), .A2(new_n532), .A3(new_n550), .ZN(new_n551));
  NAND3_X1  g365(.A1(new_n540), .A2(new_n254), .A3(new_n551), .ZN(new_n552));
  OAI21_X1  g366(.A(G210), .B1(G237), .B2(G902), .ZN(new_n553));
  INV_X1    g367(.A(new_n553), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n552), .A2(new_n554), .ZN(new_n555));
  NAND4_X1  g369(.A1(new_n540), .A2(new_n254), .A3(new_n553), .A4(new_n551), .ZN(new_n556));
  AOI21_X1  g370(.A(new_n522), .B1(new_n555), .B2(new_n556), .ZN(new_n557));
  NAND4_X1  g371(.A1(new_n405), .A2(new_n480), .A3(new_n520), .A4(new_n557), .ZN(new_n558));
  XNOR2_X1  g372(.A(new_n558), .B(G101), .ZN(G3));
  INV_X1    g373(.A(G472), .ZN(new_n560));
  AOI21_X1  g374(.A(new_n560), .B1(new_n475), .B2(new_n254), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n506), .A2(KEYINPUT75), .ZN(new_n562));
  NAND3_X1  g376(.A1(new_n498), .A2(new_n499), .A3(new_n501), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  AOI21_X1  g378(.A(new_n508), .B1(new_n564), .B2(new_n488), .ZN(new_n565));
  INV_X1    g379(.A(new_n509), .ZN(new_n566));
  NOR2_X1   g380(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  NAND4_X1  g381(.A1(new_n567), .A2(new_n511), .A3(new_n254), .A4(new_n507), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n510), .A2(KEYINPUT25), .ZN(new_n569));
  NAND3_X1  g383(.A1(new_n568), .A2(new_n569), .A3(new_n515), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n519), .A2(new_n517), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  INV_X1    g386(.A(new_n477), .ZN(new_n573));
  INV_X1    g387(.A(KEYINPUT31), .ZN(new_n574));
  NAND3_X1  g388(.A1(new_n464), .A2(new_n441), .A3(new_n431), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n575), .A2(KEYINPUT67), .ZN(new_n576));
  NAND3_X1  g390(.A1(new_n423), .A2(new_n457), .A3(new_n431), .ZN(new_n577));
  AOI21_X1  g391(.A(new_n574), .B1(new_n576), .B2(new_n577), .ZN(new_n578));
  NOR2_X1   g392(.A1(new_n472), .A2(KEYINPUT71), .ZN(new_n579));
  NOR2_X1   g393(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  AOI22_X1  g394(.A1(new_n467), .A2(new_n469), .B1(new_n472), .B2(KEYINPUT71), .ZN(new_n581));
  AOI21_X1  g395(.A(new_n573), .B1(new_n580), .B2(new_n581), .ZN(new_n582));
  NOR3_X1   g396(.A1(new_n561), .A2(new_n572), .A3(new_n582), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n402), .A2(new_n404), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n557), .A2(new_n311), .ZN(new_n585));
  INV_X1    g399(.A(new_n585), .ZN(new_n586));
  NAND3_X1  g400(.A1(new_n583), .A2(new_n584), .A3(new_n586), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n257), .A2(new_n264), .ZN(new_n588));
  INV_X1    g402(.A(KEYINPUT33), .ZN(new_n589));
  NAND3_X1  g403(.A1(new_n296), .A2(new_n589), .A3(new_n298), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n590), .A2(KEYINPUT94), .ZN(new_n591));
  INV_X1    g405(.A(KEYINPUT94), .ZN(new_n592));
  NAND4_X1  g406(.A1(new_n296), .A2(new_n592), .A3(new_n589), .A4(new_n298), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n591), .A2(new_n593), .ZN(new_n594));
  NAND3_X1  g408(.A1(new_n293), .A2(KEYINPUT33), .A3(new_n295), .ZN(new_n595));
  NOR2_X1   g409(.A1(new_n300), .A2(G902), .ZN(new_n596));
  NAND3_X1  g410(.A1(new_n594), .A2(new_n595), .A3(new_n596), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n299), .A2(new_n300), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n588), .A2(new_n599), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n600), .A2(KEYINPUT95), .ZN(new_n601));
  INV_X1    g415(.A(KEYINPUT95), .ZN(new_n602));
  NAND3_X1  g416(.A1(new_n588), .A2(new_n599), .A3(new_n602), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n601), .A2(new_n603), .ZN(new_n604));
  NOR2_X1   g418(.A1(new_n587), .A2(new_n604), .ZN(new_n605));
  XNOR2_X1  g419(.A(KEYINPUT34), .B(G104), .ZN(new_n606));
  XNOR2_X1  g420(.A(new_n605), .B(new_n606), .ZN(G6));
  NOR3_X1   g421(.A1(new_n587), .A2(new_n302), .A3(new_n588), .ZN(new_n608));
  XNOR2_X1  g422(.A(KEYINPUT35), .B(G107), .ZN(new_n609));
  XNOR2_X1  g423(.A(new_n608), .B(new_n609), .ZN(G9));
  NOR2_X1   g424(.A1(new_n561), .A2(new_n582), .ZN(new_n611));
  NOR2_X1   g425(.A1(new_n488), .A2(KEYINPUT36), .ZN(new_n612));
  XNOR2_X1  g426(.A(new_n564), .B(new_n612), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n613), .A2(new_n517), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n570), .A2(new_n614), .ZN(new_n615));
  AND2_X1   g429(.A1(new_n615), .A2(new_n557), .ZN(new_n616));
  NAND3_X1  g430(.A1(new_n405), .A2(new_n611), .A3(new_n616), .ZN(new_n617));
  XOR2_X1   g431(.A(new_n617), .B(KEYINPUT37), .Z(new_n618));
  XNOR2_X1  g432(.A(new_n618), .B(G110), .ZN(G12));
  INV_X1    g433(.A(G900), .ZN(new_n620));
  AOI21_X1  g434(.A(new_n305), .B1(new_n309), .B2(new_n620), .ZN(new_n621));
  NOR3_X1   g435(.A1(new_n588), .A2(new_n302), .A3(new_n621), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n480), .A2(new_n622), .ZN(new_n623));
  INV_X1    g437(.A(new_n404), .ZN(new_n624));
  AOI21_X1  g438(.A(KEYINPUT84), .B1(new_n403), .B2(new_n400), .ZN(new_n625));
  OAI211_X1 g439(.A(new_n557), .B(new_n615), .C1(new_n624), .C2(new_n625), .ZN(new_n626));
  OAI21_X1  g440(.A(KEYINPUT96), .B1(new_n623), .B2(new_n626), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n615), .A2(new_n557), .ZN(new_n628));
  AOI21_X1  g442(.A(new_n628), .B1(new_n402), .B2(new_n404), .ZN(new_n629));
  INV_X1    g443(.A(KEYINPUT96), .ZN(new_n630));
  NAND4_X1  g444(.A1(new_n629), .A2(new_n630), .A3(new_n480), .A4(new_n622), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n627), .A2(new_n631), .ZN(new_n632));
  XNOR2_X1  g446(.A(new_n632), .B(G128), .ZN(G30));
  AOI21_X1  g447(.A(new_n302), .B1(new_n257), .B2(new_n264), .ZN(new_n634));
  INV_X1    g448(.A(new_n634), .ZN(new_n635));
  NAND2_X1  g449(.A1(new_n555), .A2(new_n556), .ZN(new_n636));
  XOR2_X1   g450(.A(new_n636), .B(KEYINPUT38), .Z(new_n637));
  INV_X1    g451(.A(KEYINPUT40), .ZN(new_n638));
  XNOR2_X1  g452(.A(new_n621), .B(KEYINPUT39), .ZN(new_n639));
  AOI21_X1  g453(.A(new_n639), .B1(new_n402), .B2(new_n404), .ZN(new_n640));
  AOI211_X1 g454(.A(new_n635), .B(new_n637), .C1(new_n638), .C2(new_n640), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n475), .A2(new_n477), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n642), .A2(KEYINPUT32), .ZN(new_n643));
  NAND3_X1  g457(.A1(new_n475), .A2(new_n476), .A3(new_n477), .ZN(new_n644));
  NAND2_X1  g458(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  AOI21_X1  g459(.A(new_n448), .B1(new_n441), .B2(new_n435), .ZN(new_n646));
  AOI21_X1  g460(.A(new_n646), .B1(new_n576), .B2(new_n577), .ZN(new_n647));
  OAI21_X1  g461(.A(G472), .B1(new_n647), .B2(G902), .ZN(new_n648));
  AOI21_X1  g462(.A(new_n615), .B1(new_n645), .B2(new_n648), .ZN(new_n649));
  OR2_X1    g463(.A1(new_n640), .A2(new_n638), .ZN(new_n650));
  NAND4_X1  g464(.A1(new_n641), .A2(new_n521), .A3(new_n649), .A4(new_n650), .ZN(new_n651));
  XNOR2_X1  g465(.A(new_n651), .B(G143), .ZN(G45));
  INV_X1    g466(.A(new_n621), .ZN(new_n653));
  AND3_X1   g467(.A1(new_n588), .A2(new_n599), .A3(new_n653), .ZN(new_n654));
  NAND3_X1  g468(.A1(new_n629), .A2(new_n480), .A3(new_n654), .ZN(new_n655));
  XNOR2_X1  g469(.A(new_n655), .B(KEYINPUT97), .ZN(new_n656));
  XNOR2_X1  g470(.A(new_n656), .B(new_n220), .ZN(G48));
  OAI21_X1  g471(.A(new_n254), .B1(new_n380), .B2(new_n390), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n658), .A2(G469), .ZN(new_n659));
  AND3_X1   g473(.A1(new_n659), .A2(new_n399), .A3(new_n391), .ZN(new_n660));
  NAND3_X1  g474(.A1(new_n480), .A2(new_n520), .A3(new_n660), .ZN(new_n661));
  NAND3_X1  g475(.A1(new_n586), .A2(new_n601), .A3(new_n603), .ZN(new_n662));
  NOR2_X1   g476(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  XNOR2_X1  g477(.A(KEYINPUT41), .B(G113), .ZN(new_n664));
  XNOR2_X1  g478(.A(new_n664), .B(KEYINPUT98), .ZN(new_n665));
  XNOR2_X1  g479(.A(new_n663), .B(new_n665), .ZN(G15));
  AND2_X1   g480(.A1(new_n257), .A2(new_n264), .ZN(new_n667));
  INV_X1    g481(.A(new_n302), .ZN(new_n668));
  AND4_X1   g482(.A1(new_n557), .A2(new_n667), .A3(new_n311), .A4(new_n668), .ZN(new_n669));
  NAND4_X1  g483(.A1(new_n669), .A2(new_n480), .A3(new_n520), .A4(new_n660), .ZN(new_n670));
  XNOR2_X1  g484(.A(new_n670), .B(G116), .ZN(G18));
  INV_X1    g485(.A(new_n312), .ZN(new_n672));
  NAND4_X1  g486(.A1(new_n480), .A2(new_n672), .A3(new_n616), .A4(new_n660), .ZN(new_n673));
  XNOR2_X1  g487(.A(new_n673), .B(G119), .ZN(G21));
  NAND3_X1  g488(.A1(new_n557), .A2(new_n660), .A3(new_n311), .ZN(new_n675));
  INV_X1    g489(.A(new_n675), .ZN(new_n676));
  INV_X1    g490(.A(KEYINPUT99), .ZN(new_n677));
  INV_X1    g491(.A(new_n472), .ZN(new_n678));
  OAI21_X1  g492(.A(new_n677), .B1(new_n578), .B2(new_n678), .ZN(new_n679));
  NAND3_X1  g493(.A1(new_n461), .A2(KEYINPUT99), .A3(new_n472), .ZN(new_n680));
  NAND3_X1  g494(.A1(new_n679), .A2(new_n680), .A3(new_n470), .ZN(new_n681));
  AOI21_X1  g495(.A(new_n561), .B1(new_n477), .B2(new_n681), .ZN(new_n682));
  NAND4_X1  g496(.A1(new_n676), .A2(new_n682), .A3(new_n520), .A4(new_n634), .ZN(new_n683));
  XNOR2_X1  g497(.A(new_n683), .B(G122), .ZN(G24));
  NAND2_X1  g498(.A1(new_n681), .A2(new_n477), .ZN(new_n685));
  NAND2_X1  g499(.A1(new_n475), .A2(new_n254), .ZN(new_n686));
  NAND2_X1  g500(.A1(new_n686), .A2(G472), .ZN(new_n687));
  NAND4_X1  g501(.A1(new_n654), .A2(new_n685), .A3(new_n687), .A4(new_n615), .ZN(new_n688));
  INV_X1    g502(.A(new_n688), .ZN(new_n689));
  NAND2_X1  g503(.A1(new_n557), .A2(new_n660), .ZN(new_n690));
  INV_X1    g504(.A(new_n690), .ZN(new_n691));
  NAND2_X1  g505(.A1(new_n689), .A2(new_n691), .ZN(new_n692));
  XNOR2_X1  g506(.A(new_n692), .B(G125), .ZN(G27));
  AOI21_X1  g507(.A(new_n560), .B1(new_n452), .B2(new_n454), .ZN(new_n694));
  AOI21_X1  g508(.A(new_n694), .B1(new_n643), .B2(new_n644), .ZN(new_n695));
  OAI21_X1  g509(.A(KEYINPUT100), .B1(new_n695), .B2(new_n572), .ZN(new_n696));
  INV_X1    g510(.A(KEYINPUT100), .ZN(new_n697));
  NAND3_X1  g511(.A1(new_n480), .A2(new_n697), .A3(new_n520), .ZN(new_n698));
  NAND4_X1  g512(.A1(new_n555), .A2(new_n521), .A3(new_n556), .A4(new_n399), .ZN(new_n699));
  NOR2_X1   g513(.A1(new_n699), .A2(new_n398), .ZN(new_n700));
  AND3_X1   g514(.A1(new_n700), .A2(new_n654), .A3(KEYINPUT42), .ZN(new_n701));
  NAND3_X1  g515(.A1(new_n696), .A2(new_n698), .A3(new_n701), .ZN(new_n702));
  NAND4_X1  g516(.A1(new_n480), .A2(new_n520), .A3(new_n654), .A4(new_n700), .ZN(new_n703));
  INV_X1    g517(.A(KEYINPUT42), .ZN(new_n704));
  NAND2_X1  g518(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  NAND2_X1  g519(.A1(new_n702), .A2(new_n705), .ZN(new_n706));
  NAND2_X1  g520(.A1(new_n706), .A2(KEYINPUT101), .ZN(new_n707));
  INV_X1    g521(.A(KEYINPUT101), .ZN(new_n708));
  NAND3_X1  g522(.A1(new_n702), .A2(new_n708), .A3(new_n705), .ZN(new_n709));
  NAND2_X1  g523(.A1(new_n707), .A2(new_n709), .ZN(new_n710));
  XNOR2_X1  g524(.A(new_n710), .B(G131), .ZN(G33));
  NAND4_X1  g525(.A1(new_n480), .A2(new_n520), .A3(new_n622), .A4(new_n700), .ZN(new_n712));
  XNOR2_X1  g526(.A(new_n712), .B(G134), .ZN(G36));
  NOR2_X1   g527(.A1(new_n636), .A2(new_n522), .ZN(new_n714));
  XNOR2_X1  g528(.A(new_n714), .B(KEYINPUT103), .ZN(new_n715));
  INV_X1    g529(.A(new_n599), .ZN(new_n716));
  NOR3_X1   g530(.A1(new_n716), .A2(new_n588), .A3(KEYINPUT43), .ZN(new_n717));
  NAND2_X1  g531(.A1(new_n588), .A2(KEYINPUT102), .ZN(new_n718));
  INV_X1    g532(.A(KEYINPUT102), .ZN(new_n719));
  NAND3_X1  g533(.A1(new_n257), .A2(new_n264), .A3(new_n719), .ZN(new_n720));
  NAND3_X1  g534(.A1(new_n718), .A2(new_n599), .A3(new_n720), .ZN(new_n721));
  AOI21_X1  g535(.A(new_n717), .B1(new_n721), .B2(KEYINPUT43), .ZN(new_n722));
  INV_X1    g536(.A(new_n611), .ZN(new_n723));
  NAND3_X1  g537(.A1(new_n722), .A2(new_n723), .A3(new_n615), .ZN(new_n724));
  INV_X1    g538(.A(KEYINPUT44), .ZN(new_n725));
  OAI21_X1  g539(.A(new_n715), .B1(new_n724), .B2(new_n725), .ZN(new_n726));
  INV_X1    g540(.A(KEYINPUT104), .ZN(new_n727));
  OR2_X1    g541(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  NAND2_X1  g542(.A1(new_n395), .A2(new_n396), .ZN(new_n729));
  XNOR2_X1  g543(.A(new_n729), .B(KEYINPUT45), .ZN(new_n730));
  NAND2_X1  g544(.A1(new_n730), .A2(G469), .ZN(new_n731));
  NAND3_X1  g545(.A1(new_n731), .A2(KEYINPUT46), .A3(new_n392), .ZN(new_n732));
  INV_X1    g546(.A(KEYINPUT46), .ZN(new_n733));
  OAI211_X1 g547(.A(new_n733), .B(G469), .C1(new_n730), .C2(G902), .ZN(new_n734));
  NAND3_X1  g548(.A1(new_n732), .A2(new_n391), .A3(new_n734), .ZN(new_n735));
  NAND2_X1  g549(.A1(new_n735), .A2(new_n399), .ZN(new_n736));
  OR2_X1    g550(.A1(new_n736), .A2(new_n639), .ZN(new_n737));
  AOI21_X1  g551(.A(new_n737), .B1(new_n725), .B2(new_n724), .ZN(new_n738));
  NAND2_X1  g552(.A1(new_n726), .A2(new_n727), .ZN(new_n739));
  NAND3_X1  g553(.A1(new_n728), .A2(new_n738), .A3(new_n739), .ZN(new_n740));
  XNOR2_X1  g554(.A(new_n740), .B(KEYINPUT105), .ZN(new_n741));
  XNOR2_X1  g555(.A(new_n741), .B(G137), .ZN(G39));
  INV_X1    g556(.A(KEYINPUT47), .ZN(new_n743));
  NAND2_X1  g557(.A1(new_n736), .A2(new_n743), .ZN(new_n744));
  NAND3_X1  g558(.A1(new_n735), .A2(KEYINPUT47), .A3(new_n399), .ZN(new_n745));
  NAND2_X1  g559(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  NOR3_X1   g560(.A1(new_n520), .A2(new_n522), .A3(new_n636), .ZN(new_n747));
  NAND4_X1  g561(.A1(new_n746), .A2(new_n695), .A3(new_n654), .A4(new_n747), .ZN(new_n748));
  XNOR2_X1  g562(.A(new_n748), .B(G140), .ZN(G42));
  AND3_X1   g563(.A1(new_n557), .A2(new_n653), .A3(new_n634), .ZN(new_n750));
  NAND4_X1  g564(.A1(new_n649), .A2(new_n399), .A3(new_n403), .A4(new_n750), .ZN(new_n751));
  NAND4_X1  g565(.A1(new_n632), .A2(new_n655), .A3(new_n692), .A4(new_n751), .ZN(new_n752));
  INV_X1    g566(.A(KEYINPUT52), .ZN(new_n753));
  NAND2_X1  g567(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  NAND2_X1  g568(.A1(new_n754), .A2(KEYINPUT109), .ZN(new_n755));
  INV_X1    g569(.A(new_n622), .ZN(new_n756));
  NOR2_X1   g570(.A1(new_n695), .A2(new_n756), .ZN(new_n757));
  AOI21_X1  g571(.A(new_n630), .B1(new_n757), .B2(new_n629), .ZN(new_n758));
  NOR3_X1   g572(.A1(new_n623), .A2(KEYINPUT96), .A3(new_n626), .ZN(new_n759));
  OAI21_X1  g573(.A(new_n692), .B1(new_n758), .B2(new_n759), .ZN(new_n760));
  INV_X1    g574(.A(KEYINPUT108), .ZN(new_n761));
  NAND2_X1  g575(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  AND2_X1   g576(.A1(new_n751), .A2(KEYINPUT52), .ZN(new_n763));
  NAND3_X1  g577(.A1(new_n632), .A2(KEYINPUT108), .A3(new_n692), .ZN(new_n764));
  NAND4_X1  g578(.A1(new_n762), .A2(new_n655), .A3(new_n763), .A4(new_n764), .ZN(new_n765));
  INV_X1    g579(.A(KEYINPUT109), .ZN(new_n766));
  NAND3_X1  g580(.A1(new_n752), .A2(new_n766), .A3(new_n753), .ZN(new_n767));
  NAND3_X1  g581(.A1(new_n755), .A2(new_n765), .A3(new_n767), .ZN(new_n768));
  INV_X1    g582(.A(KEYINPUT53), .ZN(new_n769));
  OAI21_X1  g583(.A(new_n600), .B1(new_n302), .B2(new_n588), .ZN(new_n770));
  NAND4_X1  g584(.A1(new_n583), .A2(new_n584), .A3(new_n586), .A4(new_n770), .ZN(new_n771));
  AND3_X1   g585(.A1(new_n558), .A2(new_n771), .A3(new_n617), .ZN(new_n772));
  NAND4_X1  g586(.A1(new_n685), .A2(new_n687), .A3(new_n520), .A4(new_n634), .ZN(new_n773));
  NOR2_X1   g587(.A1(new_n773), .A2(new_n675), .ZN(new_n774));
  AND3_X1   g588(.A1(new_n480), .A2(new_n520), .A3(new_n660), .ZN(new_n775));
  NOR2_X1   g589(.A1(new_n604), .A2(new_n585), .ZN(new_n776));
  AOI21_X1  g590(.A(new_n774), .B1(new_n775), .B2(new_n776), .ZN(new_n777));
  AND2_X1   g591(.A1(new_n670), .A2(new_n673), .ZN(new_n778));
  NAND3_X1  g592(.A1(new_n772), .A2(new_n777), .A3(new_n778), .ZN(new_n779));
  OAI211_X1 g593(.A(new_n615), .B(new_n653), .C1(new_n624), .C2(new_n625), .ZN(new_n780));
  INV_X1    g594(.A(new_n780), .ZN(new_n781));
  NOR2_X1   g595(.A1(new_n588), .A2(new_n668), .ZN(new_n782));
  NAND4_X1  g596(.A1(new_n781), .A2(new_n480), .A3(new_n782), .A4(new_n714), .ZN(new_n783));
  INV_X1    g597(.A(KEYINPUT106), .ZN(new_n784));
  AOI21_X1  g598(.A(new_n784), .B1(new_n689), .B2(new_n700), .ZN(new_n785));
  INV_X1    g599(.A(new_n700), .ZN(new_n786));
  NOR3_X1   g600(.A1(new_n688), .A2(KEYINPUT106), .A3(new_n786), .ZN(new_n787));
  OAI211_X1 g601(.A(new_n712), .B(new_n783), .C1(new_n785), .C2(new_n787), .ZN(new_n788));
  NOR2_X1   g602(.A1(new_n779), .A2(new_n788), .ZN(new_n789));
  INV_X1    g603(.A(KEYINPUT107), .ZN(new_n790));
  NAND3_X1  g604(.A1(new_n789), .A2(new_n710), .A3(new_n790), .ZN(new_n791));
  AND3_X1   g605(.A1(new_n702), .A2(new_n708), .A3(new_n705), .ZN(new_n792));
  AOI21_X1  g606(.A(new_n708), .B1(new_n702), .B2(new_n705), .ZN(new_n793));
  NOR2_X1   g607(.A1(new_n792), .A2(new_n793), .ZN(new_n794));
  OAI21_X1  g608(.A(new_n683), .B1(new_n661), .B2(new_n662), .ZN(new_n795));
  NAND2_X1  g609(.A1(new_n670), .A2(new_n673), .ZN(new_n796));
  NOR2_X1   g610(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  NAND3_X1  g611(.A1(new_n689), .A2(new_n784), .A3(new_n700), .ZN(new_n798));
  OAI21_X1  g612(.A(KEYINPUT106), .B1(new_n688), .B2(new_n786), .ZN(new_n799));
  NAND2_X1  g613(.A1(new_n798), .A2(new_n799), .ZN(new_n800));
  NAND3_X1  g614(.A1(new_n480), .A2(new_n782), .A3(new_n714), .ZN(new_n801));
  OAI21_X1  g615(.A(new_n712), .B1(new_n801), .B2(new_n780), .ZN(new_n802));
  INV_X1    g616(.A(new_n802), .ZN(new_n803));
  NAND4_X1  g617(.A1(new_n797), .A2(new_n772), .A3(new_n800), .A4(new_n803), .ZN(new_n804));
  OAI21_X1  g618(.A(KEYINPUT107), .B1(new_n794), .B2(new_n804), .ZN(new_n805));
  NAND4_X1  g619(.A1(new_n768), .A2(new_n769), .A3(new_n791), .A4(new_n805), .ZN(new_n806));
  NAND4_X1  g620(.A1(new_n763), .A2(new_n632), .A3(new_n655), .A4(new_n692), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n754), .A2(new_n807), .ZN(new_n808));
  NAND3_X1  g622(.A1(new_n805), .A2(new_n791), .A3(new_n808), .ZN(new_n809));
  NAND2_X1  g623(.A1(new_n809), .A2(KEYINPUT53), .ZN(new_n810));
  NAND3_X1  g624(.A1(new_n806), .A2(new_n810), .A3(KEYINPUT54), .ZN(new_n811));
  NAND2_X1  g625(.A1(new_n809), .A2(new_n769), .ZN(new_n812));
  INV_X1    g626(.A(KEYINPUT54), .ZN(new_n813));
  AND3_X1   g627(.A1(new_n789), .A2(KEYINPUT53), .A3(new_n706), .ZN(new_n814));
  NAND2_X1  g628(.A1(new_n768), .A2(new_n814), .ZN(new_n815));
  NAND3_X1  g629(.A1(new_n812), .A2(new_n813), .A3(new_n815), .ZN(new_n816));
  NAND2_X1  g630(.A1(new_n811), .A2(new_n816), .ZN(new_n817));
  AND3_X1   g631(.A1(new_n685), .A2(new_n520), .A3(new_n687), .ZN(new_n818));
  NAND3_X1  g632(.A1(new_n722), .A2(new_n818), .A3(new_n305), .ZN(new_n819));
  INV_X1    g633(.A(new_n819), .ZN(new_n820));
  INV_X1    g634(.A(KEYINPUT50), .ZN(new_n821));
  NAND2_X1  g635(.A1(new_n821), .A2(KEYINPUT112), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n660), .A2(new_n522), .ZN(new_n823));
  XNOR2_X1  g637(.A(new_n823), .B(KEYINPUT111), .ZN(new_n824));
  INV_X1    g638(.A(new_n824), .ZN(new_n825));
  NAND4_X1  g639(.A1(new_n820), .A2(new_n637), .A3(new_n822), .A4(new_n825), .ZN(new_n826));
  NAND4_X1  g640(.A1(new_n722), .A2(new_n818), .A3(new_n305), .A4(new_n637), .ZN(new_n827));
  OAI211_X1 g641(.A(KEYINPUT112), .B(new_n821), .C1(new_n827), .C2(new_n824), .ZN(new_n828));
  NAND2_X1  g642(.A1(new_n826), .A2(new_n828), .ZN(new_n829));
  NAND2_X1  g643(.A1(new_n659), .A2(new_n391), .ZN(new_n830));
  AND2_X1   g644(.A1(new_n830), .A2(KEYINPUT110), .ZN(new_n831));
  NOR2_X1   g645(.A1(new_n830), .A2(KEYINPUT110), .ZN(new_n832));
  NOR3_X1   g646(.A1(new_n831), .A2(new_n832), .A3(new_n400), .ZN(new_n833));
  OAI211_X1 g647(.A(new_n715), .B(new_n820), .C1(new_n746), .C2(new_n833), .ZN(new_n834));
  NOR3_X1   g648(.A1(new_n699), .A2(new_n304), .A3(new_n830), .ZN(new_n835));
  NAND2_X1  g649(.A1(new_n722), .A2(new_n835), .ZN(new_n836));
  NAND2_X1  g650(.A1(new_n682), .A2(new_n615), .ZN(new_n837));
  NOR2_X1   g651(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  INV_X1    g652(.A(new_n838), .ZN(new_n839));
  NAND3_X1  g653(.A1(new_n645), .A2(new_n520), .A3(new_n648), .ZN(new_n840));
  INV_X1    g654(.A(new_n840), .ZN(new_n841));
  NAND4_X1  g655(.A1(new_n841), .A2(new_n667), .A3(new_n716), .A4(new_n835), .ZN(new_n842));
  AND4_X1   g656(.A1(new_n829), .A2(new_n834), .A3(new_n839), .A4(new_n842), .ZN(new_n843));
  OR2_X1    g657(.A1(new_n843), .A2(KEYINPUT51), .ZN(new_n844));
  AND2_X1   g658(.A1(new_n696), .A2(new_n698), .ZN(new_n845));
  INV_X1    g659(.A(new_n836), .ZN(new_n846));
  NAND2_X1  g660(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  NAND2_X1  g661(.A1(new_n847), .A2(KEYINPUT48), .ZN(new_n848));
  INV_X1    g662(.A(KEYINPUT48), .ZN(new_n849));
  NAND3_X1  g663(.A1(new_n845), .A2(new_n846), .A3(new_n849), .ZN(new_n850));
  NAND2_X1  g664(.A1(new_n848), .A2(new_n850), .ZN(new_n851));
  NAND2_X1  g665(.A1(new_n841), .A2(new_n835), .ZN(new_n852));
  OAI211_X1 g666(.A(G952), .B(new_n188), .C1(new_n852), .C2(new_n604), .ZN(new_n853));
  NAND3_X1  g667(.A1(new_n820), .A2(KEYINPUT115), .A3(new_n691), .ZN(new_n854));
  INV_X1    g668(.A(KEYINPUT115), .ZN(new_n855));
  OAI21_X1  g669(.A(new_n855), .B1(new_n819), .B2(new_n690), .ZN(new_n856));
  AOI21_X1  g670(.A(new_n853), .B1(new_n854), .B2(new_n856), .ZN(new_n857));
  AND3_X1   g671(.A1(new_n851), .A2(new_n857), .A3(KEYINPUT116), .ZN(new_n858));
  AOI21_X1  g672(.A(KEYINPUT116), .B1(new_n851), .B2(new_n857), .ZN(new_n859));
  INV_X1    g673(.A(KEYINPUT114), .ZN(new_n860));
  INV_X1    g674(.A(KEYINPUT113), .ZN(new_n861));
  NAND3_X1  g675(.A1(new_n839), .A2(new_n861), .A3(new_n842), .ZN(new_n862));
  INV_X1    g676(.A(new_n842), .ZN(new_n863));
  OAI21_X1  g677(.A(KEYINPUT113), .B1(new_n863), .B2(new_n838), .ZN(new_n864));
  AND2_X1   g678(.A1(new_n862), .A2(new_n864), .ZN(new_n865));
  AOI21_X1  g679(.A(new_n860), .B1(new_n865), .B2(new_n829), .ZN(new_n866));
  NAND4_X1  g680(.A1(new_n829), .A2(new_n862), .A3(new_n860), .A4(new_n864), .ZN(new_n867));
  NAND3_X1  g681(.A1(new_n867), .A2(KEYINPUT51), .A3(new_n834), .ZN(new_n868));
  OAI221_X1 g682(.A(new_n844), .B1(new_n858), .B2(new_n859), .C1(new_n866), .C2(new_n868), .ZN(new_n869));
  OAI22_X1  g683(.A1(new_n817), .A2(new_n869), .B1(G952), .B2(G953), .ZN(new_n870));
  XNOR2_X1  g684(.A(new_n830), .B(KEYINPUT49), .ZN(new_n871));
  NOR4_X1   g685(.A1(new_n871), .A2(new_n721), .A3(new_n572), .A4(new_n522), .ZN(new_n872));
  AND2_X1   g686(.A1(new_n645), .A2(new_n648), .ZN(new_n873));
  NAND4_X1  g687(.A1(new_n872), .A2(new_n400), .A3(new_n873), .A4(new_n637), .ZN(new_n874));
  NAND2_X1  g688(.A1(new_n870), .A2(new_n874), .ZN(new_n875));
  NAND2_X1  g689(.A1(new_n875), .A2(KEYINPUT117), .ZN(new_n876));
  INV_X1    g690(.A(KEYINPUT117), .ZN(new_n877));
  NAND3_X1  g691(.A1(new_n870), .A2(new_n877), .A3(new_n874), .ZN(new_n878));
  NAND2_X1  g692(.A1(new_n876), .A2(new_n878), .ZN(G75));
  NOR2_X1   g693(.A1(new_n188), .A2(G952), .ZN(new_n880));
  XOR2_X1   g694(.A(new_n880), .B(KEYINPUT120), .Z(new_n881));
  AOI22_X1  g695(.A1(new_n809), .A2(new_n769), .B1(new_n768), .B2(new_n814), .ZN(new_n882));
  NOR2_X1   g696(.A1(new_n882), .A2(new_n254), .ZN(new_n883));
  AOI21_X1  g697(.A(KEYINPUT56), .B1(new_n883), .B2(G210), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n533), .A2(new_n535), .ZN(new_n885));
  XNOR2_X1  g699(.A(new_n885), .B(new_n539), .ZN(new_n886));
  XNOR2_X1  g700(.A(new_n886), .B(KEYINPUT55), .ZN(new_n887));
  OAI21_X1  g701(.A(new_n881), .B1(new_n884), .B2(new_n887), .ZN(new_n888));
  NAND2_X1  g702(.A1(new_n812), .A2(new_n815), .ZN(new_n889));
  INV_X1    g703(.A(KEYINPUT118), .ZN(new_n890));
  NAND3_X1  g704(.A1(new_n889), .A2(new_n890), .A3(G902), .ZN(new_n891));
  OAI21_X1  g705(.A(KEYINPUT118), .B1(new_n882), .B2(new_n254), .ZN(new_n892));
  INV_X1    g706(.A(KEYINPUT119), .ZN(new_n893));
  NAND4_X1  g707(.A1(new_n891), .A2(new_n892), .A3(new_n893), .A4(new_n554), .ZN(new_n894));
  AND2_X1   g708(.A1(new_n894), .A2(new_n887), .ZN(new_n895));
  NAND3_X1  g709(.A1(new_n891), .A2(new_n892), .A3(new_n554), .ZN(new_n896));
  AOI21_X1  g710(.A(KEYINPUT56), .B1(new_n896), .B2(KEYINPUT119), .ZN(new_n897));
  AOI21_X1  g711(.A(new_n888), .B1(new_n895), .B2(new_n897), .ZN(G51));
  NAND2_X1  g712(.A1(new_n889), .A2(KEYINPUT54), .ZN(new_n899));
  INV_X1    g713(.A(KEYINPUT121), .ZN(new_n900));
  NAND3_X1  g714(.A1(new_n899), .A2(new_n900), .A3(new_n816), .ZN(new_n901));
  NAND3_X1  g715(.A1(new_n889), .A2(KEYINPUT121), .A3(KEYINPUT54), .ZN(new_n902));
  XOR2_X1   g716(.A(new_n392), .B(KEYINPUT57), .Z(new_n903));
  NAND3_X1  g717(.A1(new_n901), .A2(new_n902), .A3(new_n903), .ZN(new_n904));
  OR2_X1    g718(.A1(new_n380), .A2(new_n390), .ZN(new_n905));
  NAND2_X1  g719(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  NAND4_X1  g720(.A1(new_n891), .A2(new_n892), .A3(G469), .A4(new_n730), .ZN(new_n907));
  AOI21_X1  g721(.A(new_n880), .B1(new_n906), .B2(new_n907), .ZN(G54));
  INV_X1    g722(.A(new_n880), .ZN(new_n909));
  AND2_X1   g723(.A1(KEYINPUT58), .A2(G475), .ZN(new_n910));
  NAND3_X1  g724(.A1(new_n891), .A2(new_n892), .A3(new_n910), .ZN(new_n911));
  NAND2_X1  g725(.A1(new_n238), .A2(new_n252), .ZN(new_n912));
  INV_X1    g726(.A(new_n912), .ZN(new_n913));
  OAI21_X1  g727(.A(new_n909), .B1(new_n911), .B2(new_n913), .ZN(new_n914));
  NAND2_X1  g728(.A1(new_n911), .A2(new_n913), .ZN(new_n915));
  NAND2_X1  g729(.A1(new_n915), .A2(KEYINPUT122), .ZN(new_n916));
  INV_X1    g730(.A(KEYINPUT122), .ZN(new_n917));
  NAND3_X1  g731(.A1(new_n911), .A2(new_n917), .A3(new_n913), .ZN(new_n918));
  AOI21_X1  g732(.A(new_n914), .B1(new_n916), .B2(new_n918), .ZN(G60));
  NAND2_X1  g733(.A1(G478), .A2(G902), .ZN(new_n920));
  XOR2_X1   g734(.A(new_n920), .B(KEYINPUT59), .Z(new_n921));
  INV_X1    g735(.A(new_n921), .ZN(new_n922));
  AND2_X1   g736(.A1(new_n594), .A2(new_n595), .ZN(new_n923));
  XNOR2_X1  g737(.A(new_n923), .B(KEYINPUT123), .ZN(new_n924));
  AND4_X1   g738(.A1(new_n902), .A2(new_n901), .A3(new_n922), .A4(new_n924), .ZN(new_n925));
  AOI21_X1  g739(.A(new_n921), .B1(new_n811), .B2(new_n816), .ZN(new_n926));
  OAI21_X1  g740(.A(new_n881), .B1(new_n926), .B2(new_n924), .ZN(new_n927));
  NOR2_X1   g741(.A1(new_n925), .A2(new_n927), .ZN(G63));
  INV_X1    g742(.A(KEYINPUT126), .ZN(new_n929));
  XOR2_X1   g743(.A(new_n518), .B(KEYINPUT125), .Z(new_n930));
  NAND2_X1  g744(.A1(G217), .A2(G902), .ZN(new_n931));
  XNOR2_X1  g745(.A(new_n931), .B(KEYINPUT60), .ZN(new_n932));
  OAI211_X1 g746(.A(new_n929), .B(new_n930), .C1(new_n882), .C2(new_n932), .ZN(new_n933));
  AND2_X1   g747(.A1(new_n933), .A2(KEYINPUT61), .ZN(new_n934));
  INV_X1    g748(.A(new_n932), .ZN(new_n935));
  NAND3_X1  g749(.A1(new_n889), .A2(new_n613), .A3(new_n935), .ZN(new_n936));
  OAI21_X1  g750(.A(new_n930), .B1(new_n882), .B2(new_n932), .ZN(new_n937));
  NAND2_X1  g751(.A1(new_n937), .A2(KEYINPUT126), .ZN(new_n938));
  NAND4_X1  g752(.A1(new_n934), .A2(new_n881), .A3(new_n936), .A4(new_n938), .ZN(new_n939));
  NAND2_X1  g753(.A1(new_n936), .A2(KEYINPUT124), .ZN(new_n940));
  INV_X1    g754(.A(KEYINPUT124), .ZN(new_n941));
  NAND4_X1  g755(.A1(new_n889), .A2(new_n941), .A3(new_n613), .A4(new_n935), .ZN(new_n942));
  AND4_X1   g756(.A1(new_n881), .A2(new_n940), .A3(new_n937), .A4(new_n942), .ZN(new_n943));
  OAI21_X1  g757(.A(new_n939), .B1(new_n943), .B2(KEYINPUT61), .ZN(G66));
  INV_X1    g758(.A(G224), .ZN(new_n945));
  OAI21_X1  g759(.A(G953), .B1(new_n307), .B2(new_n945), .ZN(new_n946));
  INV_X1    g760(.A(new_n779), .ZN(new_n947));
  OAI21_X1  g761(.A(new_n946), .B1(new_n947), .B2(G953), .ZN(new_n948));
  OAI21_X1  g762(.A(new_n885), .B1(G898), .B2(new_n188), .ZN(new_n949));
  XNOR2_X1  g763(.A(new_n948), .B(new_n949), .ZN(G69));
  NAND2_X1  g764(.A1(G900), .A2(G953), .ZN(new_n951));
  NAND2_X1  g765(.A1(new_n740), .A2(new_n748), .ZN(new_n952));
  INV_X1    g766(.A(new_n737), .ZN(new_n953));
  AND3_X1   g767(.A1(new_n845), .A2(new_n557), .A3(new_n634), .ZN(new_n954));
  AOI21_X1  g768(.A(new_n952), .B1(new_n953), .B2(new_n954), .ZN(new_n955));
  AND3_X1   g769(.A1(new_n762), .A2(new_n655), .A3(new_n764), .ZN(new_n956));
  AND2_X1   g770(.A1(new_n710), .A2(new_n712), .ZN(new_n957));
  NAND3_X1  g771(.A1(new_n955), .A2(new_n956), .A3(new_n957), .ZN(new_n958));
  OAI21_X1  g772(.A(new_n951), .B1(new_n958), .B2(G953), .ZN(new_n959));
  NOR2_X1   g773(.A1(new_n241), .A2(new_n243), .ZN(new_n960));
  XOR2_X1   g774(.A(new_n422), .B(new_n960), .Z(new_n961));
  NAND2_X1  g775(.A1(new_n959), .A2(new_n961), .ZN(new_n962));
  NOR2_X1   g776(.A1(new_n695), .A2(new_n572), .ZN(new_n963));
  NAND4_X1  g777(.A1(new_n963), .A2(new_n640), .A3(new_n714), .A4(new_n770), .ZN(new_n964));
  AND3_X1   g778(.A1(new_n740), .A2(new_n748), .A3(new_n964), .ZN(new_n965));
  NAND4_X1  g779(.A1(new_n762), .A2(new_n651), .A3(new_n655), .A4(new_n764), .ZN(new_n966));
  INV_X1    g780(.A(KEYINPUT62), .ZN(new_n967));
  AND2_X1   g781(.A1(new_n966), .A2(new_n967), .ZN(new_n968));
  NOR2_X1   g782(.A1(new_n966), .A2(new_n967), .ZN(new_n969));
  OAI21_X1  g783(.A(new_n965), .B1(new_n968), .B2(new_n969), .ZN(new_n970));
  INV_X1    g784(.A(new_n961), .ZN(new_n971));
  NAND3_X1  g785(.A1(new_n970), .A2(new_n188), .A3(new_n971), .ZN(new_n972));
  INV_X1    g786(.A(G227), .ZN(new_n973));
  OAI21_X1  g787(.A(G953), .B1(new_n973), .B2(new_n620), .ZN(new_n974));
  AND3_X1   g788(.A1(new_n962), .A2(new_n972), .A3(new_n974), .ZN(new_n975));
  AOI21_X1  g789(.A(new_n974), .B1(new_n962), .B2(new_n972), .ZN(new_n976));
  NOR2_X1   g790(.A1(new_n975), .A2(new_n976), .ZN(G72));
  NAND2_X1  g791(.A1(G472), .A2(G902), .ZN(new_n978));
  XOR2_X1   g792(.A(new_n978), .B(KEYINPUT63), .Z(new_n979));
  OAI211_X1 g793(.A(new_n433), .B(new_n451), .C1(new_n458), .C2(new_n460), .ZN(new_n980));
  NAND4_X1  g794(.A1(new_n806), .A2(new_n810), .A3(new_n979), .A4(new_n980), .ZN(new_n981));
  NAND2_X1  g795(.A1(new_n981), .A2(new_n909), .ZN(new_n982));
  INV_X1    g796(.A(new_n423), .ZN(new_n983));
  NAND4_X1  g797(.A1(new_n955), .A2(new_n947), .A3(new_n956), .A4(new_n957), .ZN(new_n984));
  AOI211_X1 g798(.A(new_n983), .B(new_n431), .C1(new_n984), .C2(new_n979), .ZN(new_n985));
  OAI21_X1  g799(.A(new_n979), .B1(new_n970), .B2(new_n779), .ZN(new_n986));
  NAND3_X1  g800(.A1(new_n986), .A2(new_n983), .A3(new_n431), .ZN(new_n987));
  NAND2_X1  g801(.A1(new_n987), .A2(KEYINPUT127), .ZN(new_n988));
  INV_X1    g802(.A(KEYINPUT127), .ZN(new_n989));
  NAND4_X1  g803(.A1(new_n986), .A2(new_n989), .A3(new_n983), .A4(new_n431), .ZN(new_n990));
  AOI211_X1 g804(.A(new_n982), .B(new_n985), .C1(new_n988), .C2(new_n990), .ZN(G57));
endmodule


