//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 1 1 0 1 0 0 1 0 1 0 0 1 1 1 0 0 1 0 0 1 0 1 0 1 0 0 1 1 0 1 0 0 1 1 1 1 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 0 1 1 0 0 1 1 0 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:42:31 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n203, new_n204, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n603, new_n604, new_n605,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n701, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n818, new_n819, new_n820,
    new_n821, new_n822, new_n823, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n983,
    new_n984, new_n985, new_n986, new_n987, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1015, new_n1016,
    new_n1017, new_n1018, new_n1019, new_n1020, new_n1021, new_n1022,
    new_n1023, new_n1024, new_n1025, new_n1026, new_n1027, new_n1028,
    new_n1029, new_n1030, new_n1031, new_n1032, new_n1033, new_n1034,
    new_n1035, new_n1036, new_n1037, new_n1038, new_n1039, new_n1041,
    new_n1042, new_n1043, new_n1044, new_n1045, new_n1046, new_n1047,
    new_n1048, new_n1049, new_n1050, new_n1051, new_n1052, new_n1053,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1105, new_n1106, new_n1107, new_n1108,
    new_n1109, new_n1110, new_n1111, new_n1112, new_n1113, new_n1114,
    new_n1115, new_n1116, new_n1117, new_n1118, new_n1119, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1161, new_n1162, new_n1163,
    new_n1164, new_n1165, new_n1166, new_n1167, new_n1168, new_n1169,
    new_n1170, new_n1171, new_n1172, new_n1173, new_n1174, new_n1175,
    new_n1176, new_n1177, new_n1178, new_n1179, new_n1180, new_n1181,
    new_n1182, new_n1183, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1194, new_n1195,
    new_n1197, new_n1198, new_n1199, new_n1200, new_n1201, new_n1202,
    new_n1203, new_n1204, new_n1205, new_n1206, new_n1207, new_n1208,
    new_n1209, new_n1210, new_n1211, new_n1212, new_n1213, new_n1214,
    new_n1215, new_n1216, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1261, new_n1262, new_n1263,
    new_n1264, new_n1265;
  NOR4_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .A4(G77), .ZN(G353));
  OAI21_X1  g0001(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0002(.A(G1), .ZN(new_n203));
  INV_X1    g0003(.A(G20), .ZN(new_n204));
  NOR2_X1   g0004(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  INV_X1    g0005(.A(new_n205), .ZN(new_n206));
  NOR2_X1   g0006(.A1(new_n206), .A2(G13), .ZN(new_n207));
  OAI211_X1 g0007(.A(new_n207), .B(G250), .C1(G257), .C2(G264), .ZN(new_n208));
  XOR2_X1   g0008(.A(new_n208), .B(KEYINPUT0), .Z(new_n209));
  INV_X1    g0009(.A(G77), .ZN(new_n210));
  INV_X1    g0010(.A(G244), .ZN(new_n211));
  NOR2_X1   g0011(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  AOI22_X1  g0012(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n213));
  NAND2_X1  g0013(.A1(G107), .A2(G264), .ZN(new_n214));
  INV_X1    g0014(.A(G68), .ZN(new_n215));
  INV_X1    g0015(.A(G238), .ZN(new_n216));
  OAI211_X1 g0016(.A(new_n213), .B(new_n214), .C1(new_n215), .C2(new_n216), .ZN(new_n217));
  AOI211_X1 g0017(.A(new_n212), .B(new_n217), .C1(G116), .C2(G270), .ZN(new_n218));
  INV_X1    g0018(.A(G50), .ZN(new_n219));
  INV_X1    g0019(.A(G226), .ZN(new_n220));
  OAI21_X1  g0020(.A(new_n218), .B1(new_n219), .B2(new_n220), .ZN(new_n221));
  AOI21_X1  g0021(.A(new_n221), .B1(G58), .B2(G232), .ZN(new_n222));
  AOI211_X1 g0022(.A(new_n205), .B(new_n222), .C1(KEYINPUT64), .C2(KEYINPUT1), .ZN(new_n223));
  NOR2_X1   g0023(.A1(KEYINPUT64), .A2(KEYINPUT1), .ZN(new_n224));
  XNOR2_X1  g0024(.A(new_n223), .B(new_n224), .ZN(new_n225));
  NAND2_X1  g0025(.A1(G1), .A2(G13), .ZN(new_n226));
  NOR2_X1   g0026(.A1(new_n226), .A2(new_n204), .ZN(new_n227));
  NOR2_X1   g0027(.A1(G58), .A2(G68), .ZN(new_n228));
  INV_X1    g0028(.A(new_n228), .ZN(new_n229));
  NAND2_X1  g0029(.A1(new_n229), .A2(G50), .ZN(new_n230));
  INV_X1    g0030(.A(new_n230), .ZN(new_n231));
  AOI211_X1 g0031(.A(new_n209), .B(new_n225), .C1(new_n227), .C2(new_n231), .ZN(G361));
  XNOR2_X1  g0032(.A(G250), .B(G257), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n233), .B(G264), .ZN(new_n234));
  XOR2_X1   g0034(.A(new_n234), .B(G270), .Z(new_n235));
  XOR2_X1   g0035(.A(G238), .B(G244), .Z(new_n236));
  XNOR2_X1  g0036(.A(KEYINPUT65), .B(KEYINPUT2), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XOR2_X1   g0038(.A(G226), .B(G232), .Z(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XOR2_X1   g0040(.A(new_n235), .B(new_n240), .Z(G358));
  XOR2_X1   g0041(.A(G68), .B(G77), .Z(new_n242));
  XNOR2_X1  g0042(.A(G50), .B(G58), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XOR2_X1   g0044(.A(G107), .B(G116), .Z(new_n245));
  XNOR2_X1  g0045(.A(G87), .B(G97), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n245), .B(new_n246), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n244), .B(new_n247), .ZN(G351));
  INV_X1    g0048(.A(G33), .ZN(new_n249));
  INV_X1    g0049(.A(G41), .ZN(new_n250));
  OAI211_X1 g0050(.A(G1), .B(G13), .C1(new_n249), .C2(new_n250), .ZN(new_n251));
  INV_X1    g0051(.A(new_n251), .ZN(new_n252));
  INV_X1    g0052(.A(G1698), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n253), .A2(G257), .ZN(new_n254));
  NAND2_X1  g0054(.A1(G264), .A2(G1698), .ZN(new_n255));
  AND2_X1   g0055(.A1(KEYINPUT3), .A2(G33), .ZN(new_n256));
  NOR2_X1   g0056(.A1(KEYINPUT3), .A2(G33), .ZN(new_n257));
  OAI211_X1 g0057(.A(new_n254), .B(new_n255), .C1(new_n256), .C2(new_n257), .ZN(new_n258));
  INV_X1    g0058(.A(KEYINPUT3), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n259), .A2(new_n249), .ZN(new_n260));
  INV_X1    g0060(.A(G303), .ZN(new_n261));
  NAND2_X1  g0061(.A1(KEYINPUT3), .A2(G33), .ZN(new_n262));
  NAND3_X1  g0062(.A1(new_n260), .A2(new_n261), .A3(new_n262), .ZN(new_n263));
  AND3_X1   g0063(.A1(new_n252), .A2(new_n258), .A3(new_n263), .ZN(new_n264));
  INV_X1    g0064(.A(KEYINPUT81), .ZN(new_n265));
  NOR2_X1   g0065(.A1(new_n250), .A2(KEYINPUT5), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n203), .A2(G45), .ZN(new_n267));
  OAI21_X1  g0067(.A(new_n265), .B1(new_n266), .B2(new_n267), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n250), .A2(KEYINPUT5), .ZN(new_n269));
  INV_X1    g0069(.A(KEYINPUT5), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n270), .A2(G41), .ZN(new_n271));
  NAND4_X1  g0071(.A1(new_n271), .A2(KEYINPUT81), .A3(new_n203), .A4(G45), .ZN(new_n272));
  AND4_X1   g0072(.A1(G274), .A2(new_n268), .A3(new_n269), .A4(new_n272), .ZN(new_n273));
  AOI21_X1  g0073(.A(new_n264), .B1(new_n273), .B2(new_n251), .ZN(new_n274));
  NAND3_X1  g0074(.A1(new_n268), .A2(new_n269), .A3(new_n272), .ZN(new_n275));
  NAND3_X1  g0075(.A1(new_n275), .A2(G270), .A3(new_n251), .ZN(new_n276));
  INV_X1    g0076(.A(KEYINPUT82), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  NAND4_X1  g0078(.A1(new_n275), .A2(KEYINPUT82), .A3(G270), .A4(new_n251), .ZN(new_n279));
  NAND3_X1  g0079(.A1(new_n274), .A2(new_n278), .A3(new_n279), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n280), .A2(KEYINPUT83), .ZN(new_n281));
  INV_X1    g0081(.A(G169), .ZN(new_n282));
  NAND2_X1  g0082(.A1(G33), .A2(G283), .ZN(new_n283));
  INV_X1    g0083(.A(G97), .ZN(new_n284));
  OAI211_X1 g0084(.A(new_n283), .B(new_n204), .C1(G33), .C2(new_n284), .ZN(new_n285));
  NAND3_X1  g0085(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n286), .A2(new_n226), .ZN(new_n287));
  OAI211_X1 g0087(.A(new_n285), .B(new_n287), .C1(new_n204), .C2(G116), .ZN(new_n288));
  INV_X1    g0088(.A(KEYINPUT20), .ZN(new_n289));
  OR2_X1    g0089(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n288), .A2(new_n289), .ZN(new_n291));
  INV_X1    g0091(.A(G13), .ZN(new_n292));
  NOR3_X1   g0092(.A1(new_n292), .A2(new_n204), .A3(G1), .ZN(new_n293));
  AOI211_X1 g0093(.A(new_n287), .B(new_n293), .C1(new_n203), .C2(G33), .ZN(new_n294));
  AOI22_X1  g0094(.A1(new_n290), .A2(new_n291), .B1(new_n294), .B2(G116), .ZN(new_n295));
  INV_X1    g0095(.A(G116), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n293), .A2(new_n296), .ZN(new_n297));
  AOI21_X1  g0097(.A(new_n282), .B1(new_n295), .B2(new_n297), .ZN(new_n298));
  INV_X1    g0098(.A(KEYINPUT83), .ZN(new_n299));
  NAND4_X1  g0099(.A1(new_n274), .A2(new_n278), .A3(new_n299), .A4(new_n279), .ZN(new_n300));
  NAND3_X1  g0100(.A1(new_n281), .A2(new_n298), .A3(new_n300), .ZN(new_n301));
  INV_X1    g0101(.A(KEYINPUT21), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  INV_X1    g0103(.A(G179), .ZN(new_n304));
  NOR2_X1   g0104(.A1(new_n280), .A2(new_n304), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n295), .A2(new_n297), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n305), .A2(new_n306), .ZN(new_n307));
  NAND4_X1  g0107(.A1(new_n281), .A2(new_n298), .A3(KEYINPUT21), .A4(new_n300), .ZN(new_n308));
  NAND3_X1  g0108(.A1(new_n303), .A2(new_n307), .A3(new_n308), .ZN(new_n309));
  AND3_X1   g0109(.A1(new_n281), .A2(G200), .A3(new_n300), .ZN(new_n310));
  INV_X1    g0110(.A(G190), .ZN(new_n311));
  AOI21_X1  g0111(.A(new_n311), .B1(new_n281), .B2(new_n300), .ZN(new_n312));
  NOR3_X1   g0112(.A1(new_n310), .A2(new_n312), .A3(new_n306), .ZN(new_n313));
  NOR2_X1   g0113(.A1(new_n309), .A2(new_n313), .ZN(new_n314));
  OAI211_X1 g0114(.A(new_n204), .B(G87), .C1(new_n256), .C2(new_n257), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n315), .A2(KEYINPUT22), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n260), .A2(new_n262), .ZN(new_n317));
  INV_X1    g0117(.A(KEYINPUT22), .ZN(new_n318));
  NAND4_X1  g0118(.A1(new_n317), .A2(new_n318), .A3(new_n204), .A4(G87), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n316), .A2(new_n319), .ZN(new_n320));
  INV_X1    g0120(.A(KEYINPUT24), .ZN(new_n321));
  INV_X1    g0121(.A(KEYINPUT84), .ZN(new_n322));
  OAI21_X1  g0122(.A(new_n322), .B1(new_n204), .B2(G107), .ZN(new_n323));
  INV_X1    g0123(.A(KEYINPUT23), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n323), .A2(new_n324), .ZN(new_n325));
  NAND3_X1  g0125(.A1(new_n204), .A2(G33), .A3(G116), .ZN(new_n326));
  OAI211_X1 g0126(.A(new_n322), .B(KEYINPUT23), .C1(new_n204), .C2(G107), .ZN(new_n327));
  AND3_X1   g0127(.A1(new_n325), .A2(new_n326), .A3(new_n327), .ZN(new_n328));
  AND3_X1   g0128(.A1(new_n320), .A2(new_n321), .A3(new_n328), .ZN(new_n329));
  AOI21_X1  g0129(.A(new_n321), .B1(new_n320), .B2(new_n328), .ZN(new_n330));
  OAI21_X1  g0130(.A(new_n287), .B1(new_n329), .B2(new_n330), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n294), .A2(G107), .ZN(new_n332));
  INV_X1    g0132(.A(G107), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n293), .A2(new_n333), .ZN(new_n334));
  XOR2_X1   g0134(.A(new_n334), .B(KEYINPUT25), .Z(new_n335));
  NAND3_X1  g0135(.A1(new_n331), .A2(new_n332), .A3(new_n335), .ZN(new_n336));
  INV_X1    g0136(.A(new_n336), .ZN(new_n337));
  INV_X1    g0137(.A(KEYINPUT87), .ZN(new_n338));
  OAI211_X1 g0138(.A(G250), .B(new_n253), .C1(new_n256), .C2(new_n257), .ZN(new_n339));
  INV_X1    g0139(.A(KEYINPUT85), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  NAND4_X1  g0141(.A1(new_n317), .A2(KEYINPUT85), .A3(G250), .A4(new_n253), .ZN(new_n342));
  NAND2_X1  g0142(.A1(G33), .A2(G294), .ZN(new_n343));
  NAND3_X1  g0143(.A1(new_n317), .A2(G257), .A3(G1698), .ZN(new_n344));
  NAND4_X1  g0144(.A1(new_n341), .A2(new_n342), .A3(new_n343), .A4(new_n344), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n345), .A2(new_n252), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n273), .A2(new_n251), .ZN(new_n347));
  NAND3_X1  g0147(.A1(new_n275), .A2(G264), .A3(new_n251), .ZN(new_n348));
  NAND3_X1  g0148(.A1(new_n346), .A2(new_n347), .A3(new_n348), .ZN(new_n349));
  NOR2_X1   g0149(.A1(new_n349), .A2(new_n311), .ZN(new_n350));
  INV_X1    g0150(.A(new_n350), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n349), .A2(G200), .ZN(new_n352));
  NAND4_X1  g0152(.A1(new_n337), .A2(new_n338), .A3(new_n351), .A4(new_n352), .ZN(new_n353));
  NAND4_X1  g0153(.A1(new_n352), .A2(new_n332), .A3(new_n331), .A4(new_n335), .ZN(new_n354));
  OAI21_X1  g0154(.A(KEYINPUT87), .B1(new_n354), .B2(new_n350), .ZN(new_n355));
  INV_X1    g0155(.A(KEYINPUT86), .ZN(new_n356));
  AND2_X1   g0156(.A1(new_n275), .A2(new_n251), .ZN(new_n357));
  AOI22_X1  g0157(.A1(new_n357), .A2(G264), .B1(new_n345), .B2(new_n252), .ZN(new_n358));
  AOI21_X1  g0158(.A(new_n282), .B1(new_n358), .B2(new_n347), .ZN(new_n359));
  NOR2_X1   g0159(.A1(new_n349), .A2(new_n304), .ZN(new_n360));
  OAI21_X1  g0160(.A(new_n356), .B1(new_n359), .B2(new_n360), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n349), .A2(G169), .ZN(new_n362));
  OAI211_X1 g0162(.A(new_n362), .B(KEYINPUT86), .C1(new_n304), .C2(new_n349), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n361), .A2(new_n363), .ZN(new_n364));
  AOI22_X1  g0164(.A1(new_n353), .A2(new_n355), .B1(new_n364), .B2(new_n336), .ZN(new_n365));
  INV_X1    g0165(.A(KEYINPUT4), .ZN(new_n366));
  NOR2_X1   g0166(.A1(new_n366), .A2(G1698), .ZN(new_n367));
  OAI211_X1 g0167(.A(new_n367), .B(G244), .C1(new_n257), .C2(new_n256), .ZN(new_n368));
  AOI21_X1  g0168(.A(new_n211), .B1(new_n260), .B2(new_n262), .ZN(new_n369));
  OAI211_X1 g0169(.A(new_n368), .B(new_n283), .C1(new_n369), .C2(KEYINPUT4), .ZN(new_n370));
  OAI21_X1  g0170(.A(G250), .B1(new_n256), .B2(new_n257), .ZN(new_n371));
  AOI21_X1  g0171(.A(new_n253), .B1(new_n371), .B2(KEYINPUT4), .ZN(new_n372));
  OAI21_X1  g0172(.A(KEYINPUT80), .B1(new_n370), .B2(new_n372), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n371), .A2(KEYINPUT4), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n374), .A2(G1698), .ZN(new_n375));
  OAI21_X1  g0175(.A(G244), .B1(new_n256), .B2(new_n257), .ZN(new_n376));
  AOI22_X1  g0176(.A1(new_n376), .A2(new_n366), .B1(G33), .B2(G283), .ZN(new_n377));
  INV_X1    g0177(.A(KEYINPUT80), .ZN(new_n378));
  NAND4_X1  g0178(.A1(new_n375), .A2(new_n377), .A3(new_n378), .A4(new_n368), .ZN(new_n379));
  NAND3_X1  g0179(.A1(new_n373), .A2(new_n379), .A3(new_n252), .ZN(new_n380));
  AOI22_X1  g0180(.A1(new_n357), .A2(G257), .B1(new_n251), .B2(new_n273), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n380), .A2(new_n381), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n382), .A2(new_n282), .ZN(new_n383));
  INV_X1    g0183(.A(new_n287), .ZN(new_n384));
  INV_X1    g0184(.A(KEYINPUT6), .ZN(new_n385));
  NOR2_X1   g0185(.A1(new_n284), .A2(new_n333), .ZN(new_n386));
  NOR2_X1   g0186(.A1(G97), .A2(G107), .ZN(new_n387));
  OAI21_X1  g0187(.A(new_n385), .B1(new_n386), .B2(new_n387), .ZN(new_n388));
  NAND3_X1  g0188(.A1(new_n333), .A2(KEYINPUT6), .A3(G97), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n388), .A2(new_n389), .ZN(new_n390));
  NOR2_X1   g0190(.A1(G20), .A2(G33), .ZN(new_n391));
  AOI22_X1  g0191(.A1(new_n390), .A2(G20), .B1(G77), .B2(new_n391), .ZN(new_n392));
  NAND3_X1  g0192(.A1(new_n260), .A2(new_n204), .A3(new_n262), .ZN(new_n393));
  INV_X1    g0193(.A(KEYINPUT7), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n393), .A2(new_n394), .ZN(new_n395));
  NAND4_X1  g0195(.A1(new_n260), .A2(KEYINPUT7), .A3(new_n204), .A4(new_n262), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n395), .A2(new_n396), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n397), .A2(G107), .ZN(new_n398));
  AOI21_X1  g0198(.A(new_n384), .B1(new_n392), .B2(new_n398), .ZN(new_n399));
  AND2_X1   g0199(.A1(new_n294), .A2(G97), .ZN(new_n400));
  INV_X1    g0200(.A(new_n293), .ZN(new_n401));
  NOR2_X1   g0201(.A1(new_n401), .A2(G97), .ZN(new_n402));
  OR3_X1    g0202(.A1(new_n399), .A2(new_n400), .A3(new_n402), .ZN(new_n403));
  NAND3_X1  g0203(.A1(new_n380), .A2(new_n381), .A3(new_n304), .ZN(new_n404));
  NAND3_X1  g0204(.A1(new_n383), .A2(new_n403), .A3(new_n404), .ZN(new_n405));
  NOR3_X1   g0205(.A1(new_n399), .A2(new_n400), .A3(new_n402), .ZN(new_n406));
  NAND3_X1  g0206(.A1(new_n380), .A2(new_n381), .A3(G190), .ZN(new_n407));
  AND2_X1   g0207(.A1(new_n380), .A2(new_n381), .ZN(new_n408));
  INV_X1    g0208(.A(G200), .ZN(new_n409));
  OAI211_X1 g0209(.A(new_n406), .B(new_n407), .C1(new_n408), .C2(new_n409), .ZN(new_n410));
  AND2_X1   g0210(.A1(new_n405), .A2(new_n410), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n216), .A2(new_n253), .ZN(new_n412));
  OAI211_X1 g0212(.A(new_n317), .B(new_n412), .C1(G244), .C2(new_n253), .ZN(new_n413));
  NAND2_X1  g0213(.A1(G33), .A2(G116), .ZN(new_n414));
  AOI21_X1  g0214(.A(new_n251), .B1(new_n413), .B2(new_n414), .ZN(new_n415));
  AOI21_X1  g0215(.A(G250), .B1(new_n203), .B2(G45), .ZN(new_n416));
  NOR2_X1   g0216(.A1(new_n267), .A2(G274), .ZN(new_n417));
  NOR3_X1   g0217(.A1(new_n252), .A2(new_n416), .A3(new_n417), .ZN(new_n418));
  OR2_X1    g0218(.A1(new_n415), .A2(new_n418), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n419), .A2(G200), .ZN(new_n420));
  NOR2_X1   g0220(.A1(new_n415), .A2(new_n418), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n421), .A2(G190), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n294), .A2(G87), .ZN(new_n423));
  NAND3_X1  g0223(.A1(new_n317), .A2(new_n204), .A3(G68), .ZN(new_n424));
  INV_X1    g0224(.A(G87), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n387), .A2(new_n425), .ZN(new_n426));
  NAND2_X1  g0226(.A1(G33), .A2(G97), .ZN(new_n427));
  INV_X1    g0227(.A(new_n427), .ZN(new_n428));
  OAI211_X1 g0228(.A(new_n426), .B(KEYINPUT19), .C1(new_n428), .C2(G20), .ZN(new_n429));
  NOR2_X1   g0229(.A1(new_n427), .A2(G20), .ZN(new_n430));
  OAI211_X1 g0230(.A(new_n424), .B(new_n429), .C1(KEYINPUT19), .C2(new_n430), .ZN(new_n431));
  XOR2_X1   g0231(.A(KEYINPUT15), .B(G87), .Z(new_n432));
  INV_X1    g0232(.A(new_n432), .ZN(new_n433));
  AOI22_X1  g0233(.A1(new_n431), .A2(new_n287), .B1(new_n293), .B2(new_n433), .ZN(new_n434));
  NAND4_X1  g0234(.A1(new_n420), .A2(new_n422), .A3(new_n423), .A4(new_n434), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n419), .A2(new_n282), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n421), .A2(new_n304), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n294), .A2(new_n432), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n434), .A2(new_n438), .ZN(new_n439));
  NAND3_X1  g0239(.A1(new_n436), .A2(new_n437), .A3(new_n439), .ZN(new_n440));
  AND2_X1   g0240(.A1(new_n435), .A2(new_n440), .ZN(new_n441));
  NAND4_X1  g0241(.A1(new_n314), .A2(new_n365), .A3(new_n411), .A4(new_n441), .ZN(new_n442));
  INV_X1    g0242(.A(KEYINPUT14), .ZN(new_n443));
  NOR2_X1   g0243(.A1(new_n443), .A2(KEYINPUT72), .ZN(new_n444));
  OAI211_X1 g0244(.A(G232), .B(G1698), .C1(new_n256), .C2(new_n257), .ZN(new_n445));
  INV_X1    g0245(.A(KEYINPUT68), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  NAND4_X1  g0247(.A1(new_n317), .A2(KEYINPUT68), .A3(G232), .A4(G1698), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n447), .A2(new_n448), .ZN(new_n449));
  OAI211_X1 g0249(.A(G226), .B(new_n253), .C1(new_n256), .C2(new_n257), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n450), .A2(KEYINPUT67), .ZN(new_n451));
  INV_X1    g0251(.A(KEYINPUT67), .ZN(new_n452));
  NAND4_X1  g0252(.A1(new_n317), .A2(new_n452), .A3(G226), .A4(new_n253), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n451), .A2(new_n453), .ZN(new_n454));
  NAND3_X1  g0254(.A1(new_n449), .A2(new_n454), .A3(new_n427), .ZN(new_n455));
  INV_X1    g0255(.A(KEYINPUT69), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n455), .A2(new_n456), .ZN(new_n457));
  AOI21_X1  g0257(.A(new_n428), .B1(new_n447), .B2(new_n448), .ZN(new_n458));
  NAND3_X1  g0258(.A1(new_n458), .A2(KEYINPUT69), .A3(new_n454), .ZN(new_n459));
  NAND3_X1  g0259(.A1(new_n457), .A2(new_n252), .A3(new_n459), .ZN(new_n460));
  INV_X1    g0260(.A(KEYINPUT13), .ZN(new_n461));
  OAI21_X1  g0261(.A(new_n203), .B1(G41), .B2(G45), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n251), .A2(new_n462), .ZN(new_n463));
  XNOR2_X1  g0263(.A(new_n463), .B(KEYINPUT71), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n464), .A2(G238), .ZN(new_n465));
  INV_X1    g0265(.A(G274), .ZN(new_n466));
  OR2_X1    g0266(.A1(new_n462), .A2(new_n466), .ZN(new_n467));
  XOR2_X1   g0267(.A(new_n467), .B(KEYINPUT70), .Z(new_n468));
  AND2_X1   g0268(.A1(new_n465), .A2(new_n468), .ZN(new_n469));
  AND3_X1   g0269(.A1(new_n460), .A2(new_n461), .A3(new_n469), .ZN(new_n470));
  AOI21_X1  g0270(.A(new_n461), .B1(new_n460), .B2(new_n469), .ZN(new_n471));
  NOR2_X1   g0271(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  AOI21_X1  g0272(.A(new_n444), .B1(new_n472), .B2(G179), .ZN(new_n473));
  OAI21_X1  g0273(.A(G169), .B1(new_n470), .B2(new_n471), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n443), .A2(KEYINPUT72), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  INV_X1    g0276(.A(new_n475), .ZN(new_n477));
  OAI211_X1 g0277(.A(G169), .B(new_n477), .C1(new_n470), .C2(new_n471), .ZN(new_n478));
  NAND3_X1  g0278(.A1(new_n473), .A2(new_n476), .A3(new_n478), .ZN(new_n479));
  INV_X1    g0279(.A(new_n391), .ZN(new_n480));
  OAI22_X1  g0280(.A1(new_n480), .A2(new_n219), .B1(new_n204), .B2(G68), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n204), .A2(G33), .ZN(new_n482));
  NOR2_X1   g0282(.A1(new_n482), .A2(new_n210), .ZN(new_n483));
  OAI21_X1  g0283(.A(new_n287), .B1(new_n481), .B2(new_n483), .ZN(new_n484));
  XNOR2_X1  g0284(.A(new_n484), .B(KEYINPUT11), .ZN(new_n485));
  OR3_X1    g0285(.A1(new_n401), .A2(KEYINPUT12), .A3(G68), .ZN(new_n486));
  OAI21_X1  g0286(.A(KEYINPUT12), .B1(new_n401), .B2(G68), .ZN(new_n487));
  OAI21_X1  g0287(.A(new_n384), .B1(G1), .B2(new_n204), .ZN(new_n488));
  INV_X1    g0288(.A(new_n488), .ZN(new_n489));
  AOI22_X1  g0289(.A1(new_n486), .A2(new_n487), .B1(new_n489), .B2(G68), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n485), .A2(new_n490), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n479), .A2(new_n491), .ZN(new_n492));
  OAI21_X1  g0292(.A(G200), .B1(new_n470), .B2(new_n471), .ZN(new_n493));
  INV_X1    g0293(.A(new_n491), .ZN(new_n494));
  AND3_X1   g0294(.A1(new_n458), .A2(KEYINPUT69), .A3(new_n454), .ZN(new_n495));
  AOI21_X1  g0295(.A(KEYINPUT69), .B1(new_n458), .B2(new_n454), .ZN(new_n496));
  NOR3_X1   g0296(.A1(new_n495), .A2(new_n496), .A3(new_n251), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n465), .A2(new_n468), .ZN(new_n498));
  OAI21_X1  g0298(.A(KEYINPUT13), .B1(new_n497), .B2(new_n498), .ZN(new_n499));
  NAND3_X1  g0299(.A1(new_n460), .A2(new_n461), .A3(new_n469), .ZN(new_n500));
  NAND3_X1  g0300(.A1(new_n499), .A2(G190), .A3(new_n500), .ZN(new_n501));
  AND3_X1   g0301(.A1(new_n493), .A2(new_n494), .A3(new_n501), .ZN(new_n502));
  INV_X1    g0302(.A(new_n502), .ZN(new_n503));
  XNOR2_X1  g0303(.A(KEYINPUT8), .B(G58), .ZN(new_n504));
  INV_X1    g0304(.A(new_n504), .ZN(new_n505));
  AOI22_X1  g0305(.A1(new_n505), .A2(new_n391), .B1(G20), .B2(G77), .ZN(new_n506));
  OAI21_X1  g0306(.A(new_n506), .B1(new_n482), .B2(new_n433), .ZN(new_n507));
  AOI22_X1  g0307(.A1(new_n507), .A2(new_n287), .B1(new_n210), .B2(new_n293), .ZN(new_n508));
  OAI21_X1  g0308(.A(new_n508), .B1(new_n210), .B2(new_n488), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n253), .A2(G232), .ZN(new_n510));
  OAI211_X1 g0310(.A(new_n317), .B(new_n510), .C1(new_n216), .C2(new_n253), .ZN(new_n511));
  OAI211_X1 g0311(.A(new_n511), .B(new_n252), .C1(G107), .C2(new_n317), .ZN(new_n512));
  OAI211_X1 g0312(.A(new_n512), .B(new_n467), .C1(new_n211), .C2(new_n463), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n513), .A2(new_n282), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n509), .A2(new_n514), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n515), .A2(KEYINPUT66), .ZN(new_n516));
  INV_X1    g0316(.A(KEYINPUT66), .ZN(new_n517));
  NAND3_X1  g0317(.A1(new_n509), .A2(new_n517), .A3(new_n514), .ZN(new_n518));
  OAI211_X1 g0318(.A(new_n516), .B(new_n518), .C1(G179), .C2(new_n513), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n513), .A2(G200), .ZN(new_n520));
  OAI21_X1  g0320(.A(new_n520), .B1(new_n311), .B2(new_n513), .ZN(new_n521));
  OR2_X1    g0321(.A1(new_n521), .A2(new_n509), .ZN(new_n522));
  NAND4_X1  g0322(.A1(new_n492), .A2(new_n503), .A3(new_n519), .A4(new_n522), .ZN(new_n523));
  INV_X1    g0323(.A(KEYINPUT79), .ZN(new_n524));
  AOI21_X1  g0324(.A(KEYINPUT74), .B1(new_n397), .B2(G68), .ZN(new_n525));
  INV_X1    g0325(.A(KEYINPUT74), .ZN(new_n526));
  AOI211_X1 g0326(.A(new_n526), .B(new_n215), .C1(new_n395), .C2(new_n396), .ZN(new_n527));
  XNOR2_X1  g0327(.A(G58), .B(G68), .ZN(new_n528));
  AOI22_X1  g0328(.A1(new_n528), .A2(G20), .B1(G159), .B2(new_n391), .ZN(new_n529));
  INV_X1    g0329(.A(new_n529), .ZN(new_n530));
  NOR3_X1   g0330(.A1(new_n525), .A2(new_n527), .A3(new_n530), .ZN(new_n531));
  OAI21_X1  g0331(.A(KEYINPUT75), .B1(new_n531), .B2(KEYINPUT16), .ZN(new_n532));
  INV_X1    g0332(.A(new_n396), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n533), .A2(KEYINPUT73), .ZN(new_n534));
  OAI211_X1 g0334(.A(G68), .B(new_n534), .C1(new_n397), .C2(KEYINPUT73), .ZN(new_n535));
  NAND3_X1  g0335(.A1(new_n535), .A2(KEYINPUT16), .A3(new_n529), .ZN(new_n536));
  AND2_X1   g0336(.A1(new_n536), .A2(new_n287), .ZN(new_n537));
  NOR2_X1   g0337(.A1(new_n256), .A2(new_n257), .ZN(new_n538));
  AOI21_X1  g0338(.A(KEYINPUT7), .B1(new_n538), .B2(new_n204), .ZN(new_n539));
  OAI21_X1  g0339(.A(G68), .B1(new_n539), .B2(new_n533), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n540), .A2(new_n526), .ZN(new_n541));
  NAND3_X1  g0341(.A1(new_n397), .A2(KEYINPUT74), .A3(G68), .ZN(new_n542));
  NAND3_X1  g0342(.A1(new_n541), .A2(new_n529), .A3(new_n542), .ZN(new_n543));
  INV_X1    g0343(.A(KEYINPUT75), .ZN(new_n544));
  INV_X1    g0344(.A(KEYINPUT16), .ZN(new_n545));
  NAND3_X1  g0345(.A1(new_n543), .A2(new_n544), .A3(new_n545), .ZN(new_n546));
  NAND3_X1  g0346(.A1(new_n532), .A2(new_n537), .A3(new_n546), .ZN(new_n547));
  NOR2_X1   g0347(.A1(new_n505), .A2(new_n293), .ZN(new_n548));
  AOI21_X1  g0348(.A(new_n548), .B1(new_n488), .B2(new_n505), .ZN(new_n549));
  INV_X1    g0349(.A(new_n549), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n547), .A2(new_n550), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n220), .A2(G1698), .ZN(new_n552));
  OAI221_X1 g0352(.A(new_n552), .B1(G223), .B2(G1698), .C1(new_n256), .C2(new_n257), .ZN(new_n553));
  INV_X1    g0353(.A(new_n553), .ZN(new_n554));
  NAND2_X1  g0354(.A1(G33), .A2(G87), .ZN(new_n555));
  XNOR2_X1  g0355(.A(new_n555), .B(KEYINPUT76), .ZN(new_n556));
  OAI21_X1  g0356(.A(new_n252), .B1(new_n554), .B2(new_n556), .ZN(new_n557));
  NAND3_X1  g0357(.A1(new_n251), .A2(G232), .A3(new_n462), .ZN(new_n558));
  NAND3_X1  g0358(.A1(new_n557), .A2(new_n467), .A3(new_n558), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n559), .A2(G169), .ZN(new_n560));
  NAND4_X1  g0360(.A1(new_n557), .A2(G179), .A3(new_n467), .A4(new_n558), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  XNOR2_X1  g0362(.A(new_n562), .B(KEYINPUT77), .ZN(new_n563));
  AOI21_X1  g0363(.A(KEYINPUT18), .B1(new_n551), .B2(new_n563), .ZN(new_n564));
  INV_X1    g0364(.A(new_n564), .ZN(new_n565));
  NAND3_X1  g0365(.A1(new_n551), .A2(new_n563), .A3(KEYINPUT18), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n559), .A2(new_n409), .ZN(new_n568));
  OAI21_X1  g0368(.A(new_n568), .B1(G190), .B2(new_n559), .ZN(new_n569));
  NAND3_X1  g0369(.A1(new_n547), .A2(new_n550), .A3(new_n569), .ZN(new_n570));
  NAND2_X1  g0370(.A1(KEYINPUT78), .A2(KEYINPUT17), .ZN(new_n571));
  INV_X1    g0371(.A(new_n571), .ZN(new_n572));
  NOR2_X1   g0372(.A1(KEYINPUT78), .A2(KEYINPUT17), .ZN(new_n573));
  NOR2_X1   g0373(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n570), .A2(new_n574), .ZN(new_n575));
  NAND4_X1  g0375(.A1(new_n547), .A2(new_n572), .A3(new_n550), .A4(new_n569), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  INV_X1    g0377(.A(new_n577), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n253), .A2(G222), .ZN(new_n579));
  INV_X1    g0379(.A(G223), .ZN(new_n580));
  OAI211_X1 g0380(.A(new_n317), .B(new_n579), .C1(new_n580), .C2(new_n253), .ZN(new_n581));
  OAI211_X1 g0381(.A(new_n581), .B(new_n252), .C1(G77), .C2(new_n317), .ZN(new_n582));
  OAI211_X1 g0382(.A(new_n582), .B(new_n467), .C1(new_n220), .C2(new_n463), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n583), .A2(new_n282), .ZN(new_n584));
  OAI21_X1  g0384(.A(G20), .B1(new_n229), .B2(G50), .ZN(new_n585));
  INV_X1    g0385(.A(G150), .ZN(new_n586));
  OAI221_X1 g0386(.A(new_n585), .B1(new_n586), .B2(new_n480), .C1(new_n482), .C2(new_n504), .ZN(new_n587));
  AOI22_X1  g0387(.A1(new_n587), .A2(new_n287), .B1(new_n219), .B2(new_n293), .ZN(new_n588));
  OAI21_X1  g0388(.A(new_n588), .B1(new_n219), .B2(new_n488), .ZN(new_n589));
  OAI211_X1 g0389(.A(new_n584), .B(new_n589), .C1(G179), .C2(new_n583), .ZN(new_n590));
  INV_X1    g0390(.A(new_n590), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n583), .A2(G200), .ZN(new_n592));
  INV_X1    g0392(.A(KEYINPUT9), .ZN(new_n593));
  OAI221_X1 g0393(.A(new_n592), .B1(new_n311), .B2(new_n583), .C1(new_n589), .C2(new_n593), .ZN(new_n594));
  AND2_X1   g0394(.A1(new_n589), .A2(new_n593), .ZN(new_n595));
  OR3_X1    g0395(.A1(new_n594), .A2(KEYINPUT10), .A3(new_n595), .ZN(new_n596));
  OAI21_X1  g0396(.A(KEYINPUT10), .B1(new_n594), .B2(new_n595), .ZN(new_n597));
  AOI21_X1  g0397(.A(new_n591), .B1(new_n596), .B2(new_n597), .ZN(new_n598));
  NAND3_X1  g0398(.A1(new_n567), .A2(new_n578), .A3(new_n598), .ZN(new_n599));
  OR3_X1    g0399(.A1(new_n523), .A2(new_n524), .A3(new_n599), .ZN(new_n600));
  OAI21_X1  g0400(.A(new_n524), .B1(new_n523), .B2(new_n599), .ZN(new_n601));
  AOI21_X1  g0401(.A(new_n442), .B1(new_n600), .B2(new_n601), .ZN(G372));
  NAND2_X1  g0402(.A1(new_n600), .A2(new_n601), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n353), .A2(new_n355), .ZN(new_n604));
  OAI21_X1  g0404(.A(new_n336), .B1(new_n359), .B2(new_n360), .ZN(new_n605));
  NAND4_X1  g0405(.A1(new_n303), .A2(new_n605), .A3(new_n307), .A4(new_n308), .ZN(new_n606));
  NAND3_X1  g0406(.A1(new_n420), .A2(new_n434), .A3(new_n423), .ZN(new_n607));
  AND2_X1   g0407(.A1(new_n607), .A2(KEYINPUT88), .ZN(new_n608));
  NOR2_X1   g0408(.A1(new_n607), .A2(KEYINPUT88), .ZN(new_n609));
  OAI21_X1  g0409(.A(new_n422), .B1(new_n608), .B2(new_n609), .ZN(new_n610));
  NAND4_X1  g0410(.A1(new_n604), .A2(new_n606), .A3(new_n610), .A4(new_n411), .ZN(new_n611));
  INV_X1    g0411(.A(KEYINPUT26), .ZN(new_n612));
  INV_X1    g0412(.A(KEYINPUT89), .ZN(new_n613));
  AND2_X1   g0413(.A1(new_n405), .A2(new_n613), .ZN(new_n614));
  NOR2_X1   g0414(.A1(new_n405), .A2(new_n613), .ZN(new_n615));
  OAI211_X1 g0415(.A(new_n610), .B(new_n612), .C1(new_n614), .C2(new_n615), .ZN(new_n616));
  INV_X1    g0416(.A(new_n440), .ZN(new_n617));
  INV_X1    g0417(.A(new_n405), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n618), .A2(new_n441), .ZN(new_n619));
  AOI21_X1  g0419(.A(new_n617), .B1(new_n619), .B2(KEYINPUT26), .ZN(new_n620));
  NAND3_X1  g0420(.A1(new_n611), .A2(new_n616), .A3(new_n620), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n603), .A2(new_n621), .ZN(new_n622));
  AOI211_X1 g0422(.A(new_n502), .B(new_n577), .C1(new_n492), .C2(new_n519), .ZN(new_n623));
  AOI22_X1  g0423(.A1(new_n547), .A2(new_n550), .B1(new_n560), .B2(new_n561), .ZN(new_n624));
  XNOR2_X1  g0424(.A(new_n624), .B(KEYINPUT18), .ZN(new_n625));
  INV_X1    g0425(.A(new_n625), .ZN(new_n626));
  OR2_X1    g0426(.A1(new_n623), .A2(new_n626), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n596), .A2(new_n597), .ZN(new_n628));
  AOI21_X1  g0428(.A(new_n591), .B1(new_n627), .B2(new_n628), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n622), .A2(new_n629), .ZN(G369));
  INV_X1    g0430(.A(new_n306), .ZN(new_n631));
  NOR2_X1   g0431(.A1(new_n292), .A2(G20), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n632), .A2(new_n203), .ZN(new_n633));
  OR2_X1    g0433(.A1(new_n633), .A2(KEYINPUT27), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n633), .A2(KEYINPUT27), .ZN(new_n635));
  NAND3_X1  g0435(.A1(new_n634), .A2(G213), .A3(new_n635), .ZN(new_n636));
  INV_X1    g0436(.A(G343), .ZN(new_n637));
  NOR2_X1   g0437(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  INV_X1    g0438(.A(new_n638), .ZN(new_n639));
  OAI21_X1  g0439(.A(new_n314), .B1(new_n631), .B2(new_n639), .ZN(new_n640));
  NAND3_X1  g0440(.A1(new_n309), .A2(new_n306), .A3(new_n638), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  INV_X1    g0442(.A(new_n642), .ZN(new_n643));
  INV_X1    g0443(.A(G330), .ZN(new_n644));
  NOR2_X1   g0444(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  AOI21_X1  g0445(.A(new_n337), .B1(new_n361), .B2(new_n363), .ZN(new_n646));
  INV_X1    g0446(.A(new_n646), .ZN(new_n647));
  OAI211_X1 g0447(.A(new_n647), .B(new_n604), .C1(new_n337), .C2(new_n639), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n646), .A2(new_n638), .ZN(new_n649));
  AND3_X1   g0449(.A1(new_n648), .A2(KEYINPUT90), .A3(new_n649), .ZN(new_n650));
  AOI21_X1  g0450(.A(KEYINPUT90), .B1(new_n648), .B2(new_n649), .ZN(new_n651));
  OR2_X1    g0451(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n645), .A2(new_n652), .ZN(new_n653));
  XNOR2_X1  g0453(.A(new_n653), .B(KEYINPUT91), .ZN(new_n654));
  INV_X1    g0454(.A(new_n654), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n309), .A2(new_n639), .ZN(new_n656));
  INV_X1    g0456(.A(new_n656), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n652), .A2(new_n657), .ZN(new_n658));
  OR2_X1    g0458(.A1(new_n605), .A2(new_n638), .ZN(new_n659));
  AND2_X1   g0459(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n655), .A2(new_n660), .ZN(G399));
  INV_X1    g0461(.A(new_n207), .ZN(new_n662));
  NOR2_X1   g0462(.A1(new_n662), .A2(G41), .ZN(new_n663));
  INV_X1    g0463(.A(new_n663), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n664), .A2(G1), .ZN(new_n665));
  NAND3_X1  g0465(.A1(new_n387), .A2(new_n425), .A3(new_n296), .ZN(new_n666));
  OAI22_X1  g0466(.A1(new_n665), .A2(new_n666), .B1(new_n230), .B2(new_n664), .ZN(new_n667));
  XNOR2_X1  g0467(.A(new_n667), .B(KEYINPUT28), .ZN(new_n668));
  INV_X1    g0468(.A(KEYINPUT93), .ZN(new_n669));
  INV_X1    g0469(.A(KEYINPUT30), .ZN(new_n670));
  AOI21_X1  g0470(.A(new_n419), .B1(new_n669), .B2(new_n670), .ZN(new_n671));
  NAND4_X1  g0471(.A1(new_n305), .A2(new_n408), .A3(new_n671), .A4(new_n358), .ZN(new_n672));
  AOI21_X1  g0472(.A(new_n669), .B1(KEYINPUT92), .B2(new_n670), .ZN(new_n673));
  XOR2_X1   g0473(.A(new_n672), .B(new_n673), .Z(new_n674));
  AND3_X1   g0474(.A1(new_n382), .A2(new_n304), .A3(new_n349), .ZN(new_n675));
  AND4_X1   g0475(.A1(new_n419), .A2(new_n675), .A3(new_n281), .A4(new_n300), .ZN(new_n676));
  OAI21_X1  g0476(.A(new_n638), .B1(new_n674), .B2(new_n676), .ZN(new_n677));
  OR2_X1    g0477(.A1(new_n677), .A2(KEYINPUT31), .ZN(new_n678));
  OAI211_X1 g0478(.A(KEYINPUT31), .B(new_n677), .C1(new_n442), .C2(new_n638), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  NOR2_X1   g0480(.A1(new_n680), .A2(new_n644), .ZN(new_n681));
  NAND3_X1  g0481(.A1(new_n618), .A2(new_n612), .A3(new_n441), .ZN(new_n682));
  NAND3_X1  g0482(.A1(new_n604), .A2(new_n610), .A3(new_n411), .ZN(new_n683));
  NOR2_X1   g0483(.A1(new_n309), .A2(new_n646), .ZN(new_n684));
  OAI211_X1 g0484(.A(new_n440), .B(new_n682), .C1(new_n683), .C2(new_n684), .ZN(new_n685));
  OR2_X1    g0485(.A1(new_n614), .A2(new_n615), .ZN(new_n686));
  AOI21_X1  g0486(.A(new_n612), .B1(new_n686), .B2(new_n610), .ZN(new_n687));
  OAI21_X1  g0487(.A(new_n639), .B1(new_n685), .B2(new_n687), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n688), .A2(KEYINPUT96), .ZN(new_n689));
  INV_X1    g0489(.A(KEYINPUT96), .ZN(new_n690));
  OAI211_X1 g0490(.A(new_n690), .B(new_n639), .C1(new_n685), .C2(new_n687), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n689), .A2(new_n691), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n692), .A2(KEYINPUT29), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n621), .A2(new_n639), .ZN(new_n694));
  INV_X1    g0494(.A(KEYINPUT94), .ZN(new_n695));
  XNOR2_X1  g0495(.A(new_n694), .B(new_n695), .ZN(new_n696));
  XOR2_X1   g0496(.A(KEYINPUT95), .B(KEYINPUT29), .Z(new_n697));
  NAND2_X1  g0497(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  AOI21_X1  g0498(.A(new_n681), .B1(new_n693), .B2(new_n698), .ZN(new_n699));
  OAI21_X1  g0499(.A(new_n668), .B1(new_n699), .B2(G1), .ZN(G364));
  NOR2_X1   g0500(.A1(G13), .A2(G33), .ZN(new_n701));
  INV_X1    g0501(.A(new_n701), .ZN(new_n702));
  NOR2_X1   g0502(.A1(new_n702), .A2(G20), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n643), .A2(new_n703), .ZN(new_n704));
  OAI21_X1  g0504(.A(G20), .B1(KEYINPUT98), .B2(G169), .ZN(new_n705));
  AOI21_X1  g0505(.A(new_n705), .B1(KEYINPUT98), .B2(G169), .ZN(new_n706));
  NOR2_X1   g0506(.A1(new_n706), .A2(new_n226), .ZN(new_n707));
  OR2_X1    g0507(.A1(new_n707), .A2(KEYINPUT99), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n707), .A2(KEYINPUT99), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  NOR2_X1   g0510(.A1(new_n710), .A2(new_n703), .ZN(new_n711));
  XNOR2_X1  g0511(.A(new_n711), .B(KEYINPUT100), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n207), .A2(new_n317), .ZN(new_n713));
  XNOR2_X1  g0513(.A(new_n713), .B(KEYINPUT97), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n714), .A2(G355), .ZN(new_n715));
  INV_X1    g0515(.A(G45), .ZN(new_n716));
  NOR2_X1   g0516(.A1(new_n244), .A2(new_n716), .ZN(new_n717));
  NOR2_X1   g0517(.A1(new_n662), .A2(new_n317), .ZN(new_n718));
  OAI21_X1  g0518(.A(new_n718), .B1(G45), .B2(new_n230), .ZN(new_n719));
  OAI221_X1 g0519(.A(new_n715), .B1(G116), .B2(new_n207), .C1(new_n717), .C2(new_n719), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n712), .A2(new_n720), .ZN(new_n721));
  AOI21_X1  g0521(.A(new_n665), .B1(G45), .B2(new_n632), .ZN(new_n722));
  INV_X1    g0522(.A(G58), .ZN(new_n723));
  NOR2_X1   g0523(.A1(new_n204), .A2(new_n304), .ZN(new_n724));
  INV_X1    g0524(.A(KEYINPUT101), .ZN(new_n725));
  NAND2_X1  g0525(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  OAI21_X1  g0526(.A(KEYINPUT101), .B1(new_n204), .B2(new_n304), .ZN(new_n727));
  NOR2_X1   g0527(.A1(new_n311), .A2(G200), .ZN(new_n728));
  NAND3_X1  g0528(.A1(new_n726), .A2(new_n727), .A3(new_n728), .ZN(new_n729));
  NOR2_X1   g0529(.A1(G190), .A2(G200), .ZN(new_n730));
  NAND3_X1  g0530(.A1(new_n726), .A2(new_n730), .A3(new_n727), .ZN(new_n731));
  OAI22_X1  g0531(.A1(new_n723), .A2(new_n729), .B1(new_n731), .B2(new_n210), .ZN(new_n732));
  NAND2_X1  g0532(.A1(new_n724), .A2(G200), .ZN(new_n733));
  NOR2_X1   g0533(.A1(new_n733), .A2(G190), .ZN(new_n734));
  AOI21_X1  g0534(.A(new_n732), .B1(G68), .B2(new_n734), .ZN(new_n735));
  NOR2_X1   g0535(.A1(new_n204), .A2(G179), .ZN(new_n736));
  NAND3_X1  g0536(.A1(new_n736), .A2(G190), .A3(G200), .ZN(new_n737));
  INV_X1    g0537(.A(KEYINPUT102), .ZN(new_n738));
  OR2_X1    g0538(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n737), .A2(new_n738), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  NOR2_X1   g0541(.A1(new_n741), .A2(new_n425), .ZN(new_n742));
  INV_X1    g0542(.A(new_n742), .ZN(new_n743));
  NOR2_X1   g0543(.A1(new_n733), .A2(new_n311), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n744), .A2(G50), .ZN(new_n745));
  NAND2_X1  g0545(.A1(new_n736), .A2(new_n730), .ZN(new_n746));
  INV_X1    g0546(.A(new_n746), .ZN(new_n747));
  NAND3_X1  g0547(.A1(new_n747), .A2(KEYINPUT32), .A3(G159), .ZN(new_n748));
  INV_X1    g0548(.A(KEYINPUT32), .ZN(new_n749));
  INV_X1    g0549(.A(G159), .ZN(new_n750));
  OAI21_X1  g0550(.A(new_n749), .B1(new_n746), .B2(new_n750), .ZN(new_n751));
  NAND3_X1  g0551(.A1(new_n736), .A2(new_n311), .A3(G200), .ZN(new_n752));
  INV_X1    g0552(.A(new_n752), .ZN(new_n753));
  AOI22_X1  g0553(.A1(new_n748), .A2(new_n751), .B1(G107), .B2(new_n753), .ZN(new_n754));
  NAND4_X1  g0554(.A1(new_n735), .A2(new_n743), .A3(new_n745), .A4(new_n754), .ZN(new_n755));
  AOI21_X1  g0555(.A(new_n204), .B1(new_n728), .B2(new_n304), .ZN(new_n756));
  INV_X1    g0556(.A(new_n756), .ZN(new_n757));
  AOI211_X1 g0557(.A(new_n538), .B(new_n755), .C1(G97), .C2(new_n757), .ZN(new_n758));
  AOI22_X1  g0558(.A1(new_n744), .A2(G326), .B1(G329), .B2(new_n747), .ZN(new_n759));
  INV_X1    g0559(.A(G322), .ZN(new_n760));
  OAI221_X1 g0560(.A(new_n759), .B1(new_n760), .B2(new_n729), .C1(new_n741), .C2(new_n261), .ZN(new_n761));
  INV_X1    g0561(.A(G294), .ZN(new_n762));
  INV_X1    g0562(.A(new_n734), .ZN(new_n763));
  XOR2_X1   g0563(.A(KEYINPUT33), .B(G317), .Z(new_n764));
  OAI221_X1 g0564(.A(new_n538), .B1(new_n756), .B2(new_n762), .C1(new_n763), .C2(new_n764), .ZN(new_n765));
  INV_X1    g0565(.A(G311), .ZN(new_n766));
  NOR2_X1   g0566(.A1(new_n731), .A2(new_n766), .ZN(new_n767));
  INV_X1    g0567(.A(G283), .ZN(new_n768));
  NOR2_X1   g0568(.A1(new_n752), .A2(new_n768), .ZN(new_n769));
  NOR4_X1   g0569(.A1(new_n761), .A2(new_n765), .A3(new_n767), .A4(new_n769), .ZN(new_n770));
  OAI21_X1  g0570(.A(new_n710), .B1(new_n758), .B2(new_n770), .ZN(new_n771));
  NAND4_X1  g0571(.A1(new_n704), .A2(new_n721), .A3(new_n722), .A4(new_n771), .ZN(new_n772));
  XNOR2_X1  g0572(.A(new_n642), .B(G330), .ZN(new_n773));
  OAI21_X1  g0573(.A(new_n772), .B1(new_n722), .B2(new_n773), .ZN(G396));
  NAND2_X1  g0574(.A1(new_n509), .A2(new_n638), .ZN(new_n775));
  NAND3_X1  g0575(.A1(new_n519), .A2(new_n522), .A3(new_n775), .ZN(new_n776));
  OAI21_X1  g0576(.A(new_n776), .B1(new_n519), .B2(new_n775), .ZN(new_n777));
  INV_X1    g0577(.A(new_n777), .ZN(new_n778));
  NAND2_X1  g0578(.A1(new_n778), .A2(new_n701), .ZN(new_n779));
  NOR2_X1   g0579(.A1(new_n710), .A2(new_n701), .ZN(new_n780));
  NAND2_X1  g0580(.A1(new_n780), .A2(new_n210), .ZN(new_n781));
  NOR2_X1   g0581(.A1(new_n752), .A2(new_n215), .ZN(new_n782));
  AOI211_X1 g0582(.A(new_n538), .B(new_n782), .C1(G132), .C2(new_n747), .ZN(new_n783));
  OAI221_X1 g0583(.A(new_n783), .B1(new_n219), .B2(new_n741), .C1(new_n723), .C2(new_n756), .ZN(new_n784));
  XOR2_X1   g0584(.A(new_n784), .B(KEYINPUT104), .Z(new_n785));
  INV_X1    g0585(.A(new_n729), .ZN(new_n786));
  AOI22_X1  g0586(.A1(new_n786), .A2(G143), .B1(G150), .B2(new_n734), .ZN(new_n787));
  INV_X1    g0587(.A(G137), .ZN(new_n788));
  INV_X1    g0588(.A(new_n744), .ZN(new_n789));
  OAI221_X1 g0589(.A(new_n787), .B1(new_n788), .B2(new_n789), .C1(new_n750), .C2(new_n731), .ZN(new_n790));
  XOR2_X1   g0590(.A(new_n790), .B(KEYINPUT34), .Z(new_n791));
  NOR2_X1   g0591(.A1(new_n785), .A2(new_n791), .ZN(new_n792));
  INV_X1    g0592(.A(new_n741), .ZN(new_n793));
  NAND2_X1  g0593(.A1(new_n753), .A2(G87), .ZN(new_n794));
  OAI21_X1  g0594(.A(new_n794), .B1(new_n766), .B2(new_n746), .ZN(new_n795));
  INV_X1    g0595(.A(KEYINPUT103), .ZN(new_n796));
  AOI22_X1  g0596(.A1(new_n793), .A2(G107), .B1(new_n795), .B2(new_n796), .ZN(new_n797));
  OAI21_X1  g0597(.A(new_n797), .B1(new_n796), .B2(new_n795), .ZN(new_n798));
  AOI22_X1  g0598(.A1(new_n734), .A2(G283), .B1(new_n757), .B2(G97), .ZN(new_n799));
  OAI211_X1 g0599(.A(new_n799), .B(new_n538), .C1(new_n261), .C2(new_n789), .ZN(new_n800));
  NOR2_X1   g0600(.A1(new_n729), .A2(new_n762), .ZN(new_n801));
  NOR2_X1   g0601(.A1(new_n731), .A2(new_n296), .ZN(new_n802));
  NOR4_X1   g0602(.A1(new_n798), .A2(new_n800), .A3(new_n801), .A4(new_n802), .ZN(new_n803));
  OAI21_X1  g0603(.A(new_n710), .B1(new_n792), .B2(new_n803), .ZN(new_n804));
  NAND4_X1  g0604(.A1(new_n779), .A2(new_n722), .A3(new_n781), .A4(new_n804), .ZN(new_n805));
  XOR2_X1   g0605(.A(new_n805), .B(KEYINPUT105), .Z(new_n806));
  AND2_X1   g0606(.A1(new_n696), .A2(new_n778), .ZN(new_n807));
  INV_X1    g0607(.A(KEYINPUT106), .ZN(new_n808));
  NAND2_X1  g0608(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  NAND3_X1  g0609(.A1(new_n621), .A2(new_n639), .A3(new_n777), .ZN(new_n810));
  NAND2_X1  g0610(.A1(new_n810), .A2(KEYINPUT106), .ZN(new_n811));
  OAI21_X1  g0611(.A(new_n809), .B1(new_n807), .B2(new_n811), .ZN(new_n812));
  INV_X1    g0612(.A(new_n681), .ZN(new_n813));
  XNOR2_X1  g0613(.A(new_n812), .B(new_n813), .ZN(new_n814));
  INV_X1    g0614(.A(new_n722), .ZN(new_n815));
  AOI21_X1  g0615(.A(new_n806), .B1(new_n814), .B2(new_n815), .ZN(new_n816));
  INV_X1    g0616(.A(new_n816), .ZN(G384));
  INV_X1    g0617(.A(KEYINPUT40), .ZN(new_n818));
  NOR2_X1   g0618(.A1(new_n494), .A2(new_n639), .ZN(new_n819));
  AOI211_X1 g0619(.A(new_n819), .B(new_n502), .C1(new_n479), .C2(new_n491), .ZN(new_n820));
  AND3_X1   g0620(.A1(new_n479), .A2(new_n491), .A3(new_n638), .ZN(new_n821));
  OAI21_X1  g0621(.A(KEYINPUT108), .B1(new_n820), .B2(new_n821), .ZN(new_n822));
  INV_X1    g0622(.A(new_n819), .ZN(new_n823));
  NAND3_X1  g0623(.A1(new_n492), .A2(new_n503), .A3(new_n823), .ZN(new_n824));
  INV_X1    g0624(.A(KEYINPUT108), .ZN(new_n825));
  NAND3_X1  g0625(.A1(new_n479), .A2(new_n491), .A3(new_n638), .ZN(new_n826));
  NAND3_X1  g0626(.A1(new_n824), .A2(new_n825), .A3(new_n826), .ZN(new_n827));
  NAND2_X1  g0627(.A1(new_n822), .A2(new_n827), .ZN(new_n828));
  INV_X1    g0628(.A(new_n680), .ZN(new_n829));
  NAND3_X1  g0629(.A1(new_n828), .A2(new_n829), .A3(new_n777), .ZN(new_n830));
  INV_X1    g0630(.A(KEYINPUT37), .ZN(new_n831));
  NAND2_X1  g0631(.A1(new_n551), .A2(new_n563), .ZN(new_n832));
  INV_X1    g0632(.A(new_n636), .ZN(new_n833));
  AND3_X1   g0633(.A1(new_n543), .A2(new_n544), .A3(new_n545), .ZN(new_n834));
  AOI21_X1  g0634(.A(new_n544), .B1(new_n543), .B2(new_n545), .ZN(new_n835));
  NAND2_X1  g0635(.A1(new_n536), .A2(new_n287), .ZN(new_n836));
  NOR3_X1   g0636(.A1(new_n834), .A2(new_n835), .A3(new_n836), .ZN(new_n837));
  OAI21_X1  g0637(.A(new_n833), .B1(new_n837), .B2(new_n549), .ZN(new_n838));
  AND4_X1   g0638(.A1(new_n831), .A2(new_n832), .A3(new_n838), .A4(new_n570), .ZN(new_n839));
  AOI21_X1  g0639(.A(KEYINPUT16), .B1(new_n535), .B2(new_n529), .ZN(new_n840));
  OAI21_X1  g0640(.A(new_n550), .B1(new_n836), .B2(new_n840), .ZN(new_n841));
  NAND2_X1  g0641(.A1(new_n841), .A2(new_n562), .ZN(new_n842));
  NAND2_X1  g0642(.A1(new_n570), .A2(new_n842), .ZN(new_n843));
  INV_X1    g0643(.A(KEYINPUT109), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  NAND3_X1  g0645(.A1(new_n570), .A2(KEYINPUT109), .A3(new_n842), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n841), .A2(new_n833), .ZN(new_n847));
  NAND3_X1  g0647(.A1(new_n845), .A2(new_n846), .A3(new_n847), .ZN(new_n848));
  AOI21_X1  g0648(.A(new_n839), .B1(new_n848), .B2(KEYINPUT37), .ZN(new_n849));
  AOI21_X1  g0649(.A(new_n847), .B1(new_n567), .B2(new_n578), .ZN(new_n850));
  INV_X1    g0650(.A(KEYINPUT38), .ZN(new_n851));
  NOR3_X1   g0651(.A1(new_n849), .A2(new_n850), .A3(new_n851), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n846), .A2(new_n847), .ZN(new_n853));
  AOI21_X1  g0653(.A(KEYINPUT109), .B1(new_n570), .B2(new_n842), .ZN(new_n854));
  OAI21_X1  g0654(.A(KEYINPUT37), .B1(new_n853), .B2(new_n854), .ZN(new_n855));
  AND2_X1   g0655(.A1(new_n838), .A2(new_n570), .ZN(new_n856));
  NAND3_X1  g0656(.A1(new_n856), .A2(new_n831), .A3(new_n832), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n855), .A2(new_n857), .ZN(new_n858));
  AND3_X1   g0658(.A1(new_n551), .A2(KEYINPUT18), .A3(new_n563), .ZN(new_n859));
  NOR2_X1   g0659(.A1(new_n859), .A2(new_n564), .ZN(new_n860));
  OAI211_X1 g0660(.A(new_n833), .B(new_n841), .C1(new_n860), .C2(new_n577), .ZN(new_n861));
  AOI21_X1  g0661(.A(KEYINPUT38), .B1(new_n858), .B2(new_n861), .ZN(new_n862));
  NOR2_X1   g0662(.A1(new_n852), .A2(new_n862), .ZN(new_n863));
  OAI21_X1  g0663(.A(new_n818), .B1(new_n830), .B2(new_n863), .ZN(new_n864));
  INV_X1    g0664(.A(new_n624), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n856), .A2(new_n865), .ZN(new_n866));
  AOI21_X1  g0666(.A(new_n839), .B1(new_n866), .B2(KEYINPUT37), .ZN(new_n867));
  AOI21_X1  g0667(.A(new_n838), .B1(new_n625), .B2(new_n578), .ZN(new_n868));
  OAI21_X1  g0668(.A(new_n851), .B1(new_n867), .B2(new_n868), .ZN(new_n869));
  NAND3_X1  g0669(.A1(new_n858), .A2(KEYINPUT38), .A3(new_n861), .ZN(new_n870));
  AOI21_X1  g0670(.A(new_n818), .B1(new_n869), .B2(new_n870), .ZN(new_n871));
  NAND4_X1  g0671(.A1(new_n871), .A2(new_n829), .A3(new_n777), .A4(new_n828), .ZN(new_n872));
  NAND3_X1  g0672(.A1(new_n864), .A2(G330), .A3(new_n872), .ZN(new_n873));
  NAND3_X1  g0673(.A1(new_n603), .A2(G330), .A3(new_n829), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  NAND4_X1  g0675(.A1(new_n864), .A2(new_n603), .A3(new_n829), .A4(new_n872), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  NOR2_X1   g0677(.A1(new_n519), .A2(new_n638), .ZN(new_n878));
  INV_X1    g0678(.A(new_n878), .ZN(new_n879));
  AND3_X1   g0679(.A1(new_n810), .A2(KEYINPUT107), .A3(new_n879), .ZN(new_n880));
  AOI21_X1  g0680(.A(KEYINPUT107), .B1(new_n810), .B2(new_n879), .ZN(new_n881));
  NOR3_X1   g0681(.A1(new_n820), .A2(KEYINPUT108), .A3(new_n821), .ZN(new_n882));
  AOI21_X1  g0682(.A(new_n825), .B1(new_n824), .B2(new_n826), .ZN(new_n883));
  OAI22_X1  g0683(.A1(new_n880), .A2(new_n881), .B1(new_n882), .B2(new_n883), .ZN(new_n884));
  OAI22_X1  g0684(.A1(new_n884), .A2(new_n863), .B1(new_n625), .B2(new_n833), .ZN(new_n885));
  INV_X1    g0685(.A(KEYINPUT39), .ZN(new_n886));
  NAND3_X1  g0686(.A1(new_n869), .A2(new_n870), .A3(new_n886), .ZN(new_n887));
  OAI21_X1  g0687(.A(new_n851), .B1(new_n849), .B2(new_n850), .ZN(new_n888));
  AOI21_X1  g0688(.A(new_n886), .B1(new_n888), .B2(new_n870), .ZN(new_n889));
  INV_X1    g0689(.A(KEYINPUT110), .ZN(new_n890));
  OAI21_X1  g0690(.A(new_n887), .B1(new_n889), .B2(new_n890), .ZN(new_n891));
  NAND4_X1  g0691(.A1(new_n869), .A2(new_n870), .A3(KEYINPUT110), .A4(new_n886), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  NAND3_X1  g0693(.A1(new_n479), .A2(new_n491), .A3(new_n639), .ZN(new_n894));
  INV_X1    g0694(.A(new_n894), .ZN(new_n895));
  AOI21_X1  g0695(.A(new_n885), .B1(new_n893), .B2(new_n895), .ZN(new_n896));
  XNOR2_X1  g0696(.A(new_n877), .B(new_n896), .ZN(new_n897));
  NAND3_X1  g0697(.A1(new_n693), .A2(new_n698), .A3(new_n603), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n898), .A2(new_n629), .ZN(new_n899));
  XNOR2_X1  g0699(.A(new_n897), .B(new_n899), .ZN(new_n900));
  OAI21_X1  g0700(.A(new_n900), .B1(new_n203), .B2(new_n632), .ZN(new_n901));
  AOI21_X1  g0701(.A(new_n296), .B1(new_n390), .B2(KEYINPUT35), .ZN(new_n902));
  OAI211_X1 g0702(.A(new_n902), .B(new_n227), .C1(KEYINPUT35), .C2(new_n390), .ZN(new_n903));
  XNOR2_X1  g0703(.A(new_n903), .B(KEYINPUT36), .ZN(new_n904));
  OAI21_X1  g0704(.A(G77), .B1(new_n723), .B2(new_n215), .ZN(new_n905));
  OAI22_X1  g0705(.A1(new_n230), .A2(new_n905), .B1(G50), .B2(new_n215), .ZN(new_n906));
  NAND3_X1  g0706(.A1(new_n906), .A2(G1), .A3(new_n292), .ZN(new_n907));
  NAND3_X1  g0707(.A1(new_n901), .A2(new_n904), .A3(new_n907), .ZN(G367));
  OAI21_X1  g0708(.A(new_n411), .B1(new_n406), .B2(new_n639), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n618), .A2(new_n638), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  NAND3_X1  g0711(.A1(new_n652), .A2(new_n657), .A3(new_n911), .ZN(new_n912));
  OR2_X1    g0712(.A1(new_n912), .A2(KEYINPUT42), .ZN(new_n913));
  OAI21_X1  g0713(.A(new_n405), .B1(new_n909), .B2(new_n647), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n914), .A2(new_n639), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n912), .A2(KEYINPUT42), .ZN(new_n916));
  NAND3_X1  g0716(.A1(new_n913), .A2(new_n915), .A3(new_n916), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n434), .A2(new_n423), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n918), .A2(new_n638), .ZN(new_n919));
  INV_X1    g0719(.A(new_n610), .ZN(new_n920));
  OAI21_X1  g0720(.A(new_n919), .B1(new_n920), .B2(new_n617), .ZN(new_n921));
  OAI21_X1  g0721(.A(new_n921), .B1(new_n617), .B2(new_n919), .ZN(new_n922));
  INV_X1    g0722(.A(KEYINPUT43), .ZN(new_n923));
  OR2_X1    g0723(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n917), .A2(new_n924), .ZN(new_n925));
  NAND3_X1  g0725(.A1(new_n925), .A2(new_n923), .A3(new_n922), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n922), .A2(new_n923), .ZN(new_n927));
  NAND3_X1  g0727(.A1(new_n917), .A2(new_n927), .A3(new_n924), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n926), .A2(new_n928), .ZN(new_n929));
  INV_X1    g0729(.A(new_n911), .ZN(new_n930));
  NOR2_X1   g0730(.A1(new_n655), .A2(new_n930), .ZN(new_n931));
  XNOR2_X1  g0731(.A(new_n929), .B(new_n931), .ZN(new_n932));
  XNOR2_X1  g0732(.A(new_n663), .B(KEYINPUT41), .ZN(new_n933));
  INV_X1    g0733(.A(new_n933), .ZN(new_n934));
  OAI21_X1  g0734(.A(KEYINPUT111), .B1(new_n660), .B2(new_n911), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n658), .A2(new_n659), .ZN(new_n936));
  INV_X1    g0736(.A(KEYINPUT111), .ZN(new_n937));
  NAND3_X1  g0737(.A1(new_n936), .A2(new_n937), .A3(new_n930), .ZN(new_n938));
  NAND3_X1  g0738(.A1(new_n935), .A2(KEYINPUT44), .A3(new_n938), .ZN(new_n939));
  INV_X1    g0739(.A(KEYINPUT44), .ZN(new_n940));
  AOI21_X1  g0740(.A(new_n937), .B1(new_n936), .B2(new_n930), .ZN(new_n941));
  AOI211_X1 g0741(.A(KEYINPUT111), .B(new_n911), .C1(new_n658), .C2(new_n659), .ZN(new_n942));
  OAI21_X1  g0742(.A(new_n940), .B1(new_n941), .B2(new_n942), .ZN(new_n943));
  NAND3_X1  g0743(.A1(new_n658), .A2(new_n659), .A3(new_n911), .ZN(new_n944));
  INV_X1    g0744(.A(KEYINPUT45), .ZN(new_n945));
  XNOR2_X1  g0745(.A(new_n944), .B(new_n945), .ZN(new_n946));
  NAND3_X1  g0746(.A1(new_n939), .A2(new_n943), .A3(new_n946), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n947), .A2(new_n654), .ZN(new_n948));
  NAND4_X1  g0748(.A1(new_n939), .A2(new_n943), .A3(new_n655), .A4(new_n946), .ZN(new_n949));
  NOR2_X1   g0749(.A1(new_n645), .A2(new_n657), .ZN(new_n950));
  XNOR2_X1  g0750(.A(new_n950), .B(new_n652), .ZN(new_n951));
  AND2_X1   g0751(.A1(new_n951), .A2(new_n699), .ZN(new_n952));
  NAND3_X1  g0752(.A1(new_n948), .A2(new_n949), .A3(new_n952), .ZN(new_n953));
  AOI21_X1  g0753(.A(new_n934), .B1(new_n953), .B2(new_n699), .ZN(new_n954));
  AOI21_X1  g0754(.A(new_n203), .B1(new_n632), .B2(G45), .ZN(new_n955));
  INV_X1    g0755(.A(new_n955), .ZN(new_n956));
  OAI21_X1  g0756(.A(new_n932), .B1(new_n954), .B2(new_n956), .ZN(new_n957));
  OAI22_X1  g0757(.A1(new_n756), .A2(new_n215), .B1(new_n746), .B2(new_n788), .ZN(new_n958));
  INV_X1    g0758(.A(new_n731), .ZN(new_n959));
  AOI211_X1 g0759(.A(new_n538), .B(new_n958), .C1(G50), .C2(new_n959), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n734), .A2(G159), .ZN(new_n961));
  NOR2_X1   g0761(.A1(new_n752), .A2(new_n210), .ZN(new_n962));
  AOI21_X1  g0762(.A(new_n962), .B1(G143), .B2(new_n744), .ZN(new_n963));
  AND3_X1   g0763(.A1(new_n960), .A2(new_n961), .A3(new_n963), .ZN(new_n964));
  OAI221_X1 g0764(.A(new_n964), .B1(new_n723), .B2(new_n741), .C1(new_n586), .C2(new_n729), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n793), .A2(G116), .ZN(new_n966));
  XNOR2_X1  g0766(.A(new_n966), .B(KEYINPUT46), .ZN(new_n967));
  NOR2_X1   g0767(.A1(new_n752), .A2(new_n284), .ZN(new_n968));
  XOR2_X1   g0768(.A(KEYINPUT112), .B(G317), .Z(new_n969));
  AOI211_X1 g0769(.A(new_n317), .B(new_n968), .C1(new_n747), .C2(new_n969), .ZN(new_n970));
  AOI22_X1  g0770(.A1(new_n959), .A2(G283), .B1(G311), .B2(new_n744), .ZN(new_n971));
  AND3_X1   g0771(.A1(new_n967), .A2(new_n970), .A3(new_n971), .ZN(new_n972));
  OAI221_X1 g0772(.A(new_n972), .B1(new_n762), .B2(new_n763), .C1(new_n261), .C2(new_n729), .ZN(new_n973));
  NOR2_X1   g0773(.A1(new_n756), .A2(new_n333), .ZN(new_n974));
  OAI21_X1  g0774(.A(new_n965), .B1(new_n973), .B2(new_n974), .ZN(new_n975));
  XNOR2_X1  g0775(.A(new_n975), .B(KEYINPUT47), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n976), .A2(new_n710), .ZN(new_n977));
  AOI21_X1  g0777(.A(new_n815), .B1(new_n922), .B2(new_n703), .ZN(new_n978));
  INV_X1    g0778(.A(new_n718), .ZN(new_n979));
  OAI221_X1 g0779(.A(new_n711), .B1(new_n207), .B2(new_n433), .C1(new_n235), .C2(new_n979), .ZN(new_n980));
  NAND3_X1  g0780(.A1(new_n977), .A2(new_n978), .A3(new_n980), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n957), .A2(new_n981), .ZN(G387));
  INV_X1    g0782(.A(new_n712), .ZN(new_n983));
  AOI21_X1  g0783(.A(new_n979), .B1(new_n240), .B2(G45), .ZN(new_n984));
  AND2_X1   g0784(.A1(new_n714), .A2(new_n666), .ZN(new_n985));
  NOR2_X1   g0785(.A1(new_n504), .A2(G50), .ZN(new_n986));
  XNOR2_X1  g0786(.A(new_n986), .B(KEYINPUT50), .ZN(new_n987));
  OAI211_X1 g0787(.A(new_n987), .B(new_n716), .C1(new_n215), .C2(new_n210), .ZN(new_n988));
  OAI22_X1  g0788(.A1(new_n984), .A2(new_n985), .B1(new_n666), .B2(new_n988), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n662), .A2(new_n333), .ZN(new_n990));
  AOI21_X1  g0790(.A(new_n983), .B1(new_n989), .B2(new_n990), .ZN(new_n991));
  NOR2_X1   g0791(.A1(new_n731), .A2(new_n215), .ZN(new_n992));
  NOR2_X1   g0792(.A1(new_n741), .A2(new_n210), .ZN(new_n993));
  AOI211_X1 g0793(.A(new_n992), .B(new_n993), .C1(G159), .C2(new_n744), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n757), .A2(new_n432), .ZN(new_n995));
  OAI21_X1  g0795(.A(new_n995), .B1(new_n586), .B2(new_n746), .ZN(new_n996));
  AOI211_X1 g0796(.A(new_n968), .B(new_n996), .C1(G50), .C2(new_n786), .ZN(new_n997));
  NAND2_X1  g0797(.A1(new_n734), .A2(new_n505), .ZN(new_n998));
  NAND4_X1  g0798(.A1(new_n994), .A2(new_n997), .A3(new_n317), .A4(new_n998), .ZN(new_n999));
  AOI22_X1  g0799(.A1(new_n959), .A2(G303), .B1(G322), .B2(new_n744), .ZN(new_n1000));
  OAI21_X1  g0800(.A(new_n1000), .B1(new_n766), .B2(new_n763), .ZN(new_n1001));
  AOI21_X1  g0801(.A(new_n1001), .B1(new_n786), .B2(new_n969), .ZN(new_n1002));
  XOR2_X1   g0802(.A(new_n1002), .B(KEYINPUT48), .Z(new_n1003));
  OAI221_X1 g0803(.A(new_n1003), .B1(new_n768), .B2(new_n756), .C1(new_n762), .C2(new_n741), .ZN(new_n1004));
  XOR2_X1   g0804(.A(new_n1004), .B(KEYINPUT49), .Z(new_n1005));
  AOI21_X1  g0805(.A(new_n317), .B1(new_n747), .B2(G326), .ZN(new_n1006));
  OAI21_X1  g0806(.A(new_n1006), .B1(new_n296), .B2(new_n752), .ZN(new_n1007));
  OAI21_X1  g0807(.A(new_n999), .B1(new_n1005), .B2(new_n1007), .ZN(new_n1008));
  AOI211_X1 g0808(.A(new_n815), .B(new_n991), .C1(new_n1008), .C2(new_n710), .ZN(new_n1009));
  INV_X1    g0809(.A(new_n703), .ZN(new_n1010));
  OR2_X1    g0810(.A1(new_n652), .A2(new_n1010), .ZN(new_n1011));
  AOI22_X1  g0811(.A1(new_n956), .A2(new_n951), .B1(new_n1009), .B2(new_n1011), .ZN(new_n1012));
  OAI21_X1  g0812(.A(new_n663), .B1(new_n951), .B2(new_n699), .ZN(new_n1013));
  OAI21_X1  g0813(.A(new_n1012), .B1(new_n1013), .B2(new_n952), .ZN(G393));
  NAND3_X1  g0814(.A1(new_n948), .A2(new_n956), .A3(new_n949), .ZN(new_n1015));
  NAND2_X1  g0815(.A1(new_n930), .A2(new_n703), .ZN(new_n1016));
  AOI22_X1  g0816(.A1(new_n786), .A2(G311), .B1(G317), .B2(new_n744), .ZN(new_n1017));
  XNOR2_X1  g0817(.A(new_n1017), .B(KEYINPUT52), .ZN(new_n1018));
  NOR2_X1   g0818(.A1(new_n1018), .A2(new_n317), .ZN(new_n1019));
  OAI221_X1 g0819(.A(new_n1019), .B1(new_n762), .B2(new_n731), .C1(new_n760), .C2(new_n746), .ZN(new_n1020));
  NOR2_X1   g0820(.A1(new_n763), .A2(new_n261), .ZN(new_n1021));
  NOR2_X1   g0821(.A1(new_n756), .A2(new_n296), .ZN(new_n1022));
  OAI22_X1  g0822(.A1(new_n741), .A2(new_n768), .B1(new_n333), .B2(new_n752), .ZN(new_n1023));
  NOR4_X1   g0823(.A1(new_n1020), .A2(new_n1021), .A3(new_n1022), .A4(new_n1023), .ZN(new_n1024));
  OAI22_X1  g0824(.A1(new_n789), .A2(new_n586), .B1(new_n750), .B2(new_n729), .ZN(new_n1025));
  XNOR2_X1  g0825(.A(new_n1025), .B(KEYINPUT51), .ZN(new_n1026));
  OAI221_X1 g0826(.A(new_n1026), .B1(new_n210), .B2(new_n756), .C1(new_n504), .C2(new_n731), .ZN(new_n1027));
  NOR2_X1   g0827(.A1(new_n741), .A2(new_n215), .ZN(new_n1028));
  NAND2_X1  g0828(.A1(new_n747), .A2(G143), .ZN(new_n1029));
  OAI211_X1 g0829(.A(new_n794), .B(new_n1029), .C1(new_n763), .C2(new_n219), .ZN(new_n1030));
  NOR4_X1   g0830(.A1(new_n1027), .A2(new_n538), .A3(new_n1028), .A4(new_n1030), .ZN(new_n1031));
  OAI21_X1  g0831(.A(new_n710), .B1(new_n1024), .B2(new_n1031), .ZN(new_n1032));
  INV_X1    g0832(.A(new_n711), .ZN(new_n1033));
  OAI22_X1  g0833(.A1(new_n979), .A2(new_n247), .B1(new_n284), .B2(new_n207), .ZN(new_n1034));
  OAI21_X1  g0834(.A(new_n722), .B1(new_n1033), .B2(new_n1034), .ZN(new_n1035));
  XNOR2_X1  g0835(.A(new_n1035), .B(KEYINPUT113), .ZN(new_n1036));
  NAND3_X1  g0836(.A1(new_n1016), .A2(new_n1032), .A3(new_n1036), .ZN(new_n1037));
  NAND2_X1  g0837(.A1(new_n953), .A2(new_n663), .ZN(new_n1038));
  AOI21_X1  g0838(.A(new_n952), .B1(new_n948), .B2(new_n949), .ZN(new_n1039));
  OAI211_X1 g0839(.A(new_n1015), .B(new_n1037), .C1(new_n1038), .C2(new_n1039), .ZN(G390));
  AND3_X1   g0840(.A1(new_n898), .A2(new_n874), .A3(new_n629), .ZN(new_n1041));
  NAND4_X1  g0841(.A1(new_n678), .A2(new_n679), .A3(G330), .A4(new_n777), .ZN(new_n1042));
  INV_X1    g0842(.A(new_n1042), .ZN(new_n1043));
  NOR2_X1   g0843(.A1(new_n1043), .A2(new_n828), .ZN(new_n1044));
  NOR2_X1   g0844(.A1(new_n882), .A2(new_n883), .ZN(new_n1045));
  NOR2_X1   g0845(.A1(new_n1045), .A2(new_n1042), .ZN(new_n1046));
  OAI22_X1  g0846(.A1(new_n1044), .A2(new_n1046), .B1(new_n881), .B2(new_n880), .ZN(new_n1047));
  AOI21_X1  g0847(.A(new_n878), .B1(new_n692), .B2(new_n777), .ZN(new_n1048));
  NAND3_X1  g0848(.A1(new_n681), .A2(new_n777), .A3(new_n828), .ZN(new_n1049));
  NAND2_X1  g0849(.A1(new_n1045), .A2(new_n1042), .ZN(new_n1050));
  NAND3_X1  g0850(.A1(new_n1048), .A2(new_n1049), .A3(new_n1050), .ZN(new_n1051));
  NAND2_X1  g0851(.A1(new_n1047), .A2(new_n1051), .ZN(new_n1052));
  INV_X1    g0852(.A(KEYINPUT114), .ZN(new_n1053));
  NAND2_X1  g0853(.A1(new_n884), .A2(new_n894), .ZN(new_n1054));
  NAND3_X1  g0854(.A1(new_n1054), .A2(new_n891), .A3(new_n892), .ZN(new_n1055));
  AOI21_X1  g0855(.A(new_n895), .B1(new_n869), .B2(new_n870), .ZN(new_n1056));
  OAI21_X1  g0856(.A(new_n1056), .B1(new_n1048), .B2(new_n1045), .ZN(new_n1057));
  AOI211_X1 g0857(.A(new_n1053), .B(new_n1046), .C1(new_n1055), .C2(new_n1057), .ZN(new_n1058));
  NAND2_X1  g0858(.A1(new_n1049), .A2(KEYINPUT114), .ZN(new_n1059));
  NAND2_X1  g0859(.A1(new_n1046), .A2(new_n1053), .ZN(new_n1060));
  NAND4_X1  g0860(.A1(new_n1055), .A2(new_n1057), .A3(new_n1059), .A4(new_n1060), .ZN(new_n1061));
  INV_X1    g0861(.A(new_n1061), .ZN(new_n1062));
  OAI211_X1 g0862(.A(new_n1041), .B(new_n1052), .C1(new_n1058), .C2(new_n1062), .ZN(new_n1063));
  NAND2_X1  g0863(.A1(new_n1055), .A2(new_n1057), .ZN(new_n1064));
  NAND3_X1  g0864(.A1(new_n1064), .A2(KEYINPUT114), .A3(new_n1049), .ZN(new_n1065));
  NAND2_X1  g0865(.A1(new_n1052), .A2(new_n1041), .ZN(new_n1066));
  NAND3_X1  g0866(.A1(new_n1065), .A2(new_n1066), .A3(new_n1061), .ZN(new_n1067));
  NAND3_X1  g0867(.A1(new_n1063), .A2(new_n663), .A3(new_n1067), .ZN(new_n1068));
  INV_X1    g0868(.A(KEYINPUT117), .ZN(new_n1069));
  AOI21_X1  g0869(.A(new_n955), .B1(new_n1065), .B2(new_n1061), .ZN(new_n1070));
  INV_X1    g0870(.A(new_n892), .ZN(new_n1071));
  OAI21_X1  g0871(.A(KEYINPUT39), .B1(new_n852), .B2(new_n862), .ZN(new_n1072));
  NAND2_X1  g0872(.A1(new_n1072), .A2(KEYINPUT110), .ZN(new_n1073));
  AOI21_X1  g0873(.A(new_n1071), .B1(new_n1073), .B2(new_n887), .ZN(new_n1074));
  NAND2_X1  g0874(.A1(new_n1074), .A2(new_n701), .ZN(new_n1075));
  OAI21_X1  g0875(.A(new_n317), .B1(new_n752), .B2(new_n219), .ZN(new_n1076));
  XNOR2_X1  g0876(.A(new_n1076), .B(KEYINPUT115), .ZN(new_n1077));
  XOR2_X1   g0877(.A(KEYINPUT54), .B(G143), .Z(new_n1078));
  NAND2_X1  g0878(.A1(new_n959), .A2(new_n1078), .ZN(new_n1079));
  INV_X1    g0879(.A(G125), .ZN(new_n1080));
  OAI221_X1 g0880(.A(new_n1079), .B1(new_n1080), .B2(new_n746), .C1(new_n750), .C2(new_n756), .ZN(new_n1081));
  AOI211_X1 g0881(.A(new_n1077), .B(new_n1081), .C1(G132), .C2(new_n786), .ZN(new_n1082));
  NOR2_X1   g0882(.A1(new_n741), .A2(new_n586), .ZN(new_n1083));
  XNOR2_X1  g0883(.A(new_n1083), .B(KEYINPUT53), .ZN(new_n1084));
  NAND2_X1  g0884(.A1(new_n734), .A2(G137), .ZN(new_n1085));
  NAND3_X1  g0885(.A1(new_n1082), .A2(new_n1084), .A3(new_n1085), .ZN(new_n1086));
  AOI21_X1  g0886(.A(new_n1086), .B1(G128), .B2(new_n744), .ZN(new_n1087));
  AOI211_X1 g0887(.A(new_n782), .B(new_n742), .C1(G294), .C2(new_n747), .ZN(new_n1088));
  OAI22_X1  g0888(.A1(new_n729), .A2(new_n296), .B1(new_n210), .B2(new_n756), .ZN(new_n1089));
  AOI211_X1 g0889(.A(new_n317), .B(new_n1089), .C1(G283), .C2(new_n744), .ZN(new_n1090));
  OAI211_X1 g0890(.A(new_n1088), .B(new_n1090), .C1(new_n284), .C2(new_n731), .ZN(new_n1091));
  AOI21_X1  g0891(.A(new_n1091), .B1(G107), .B2(new_n734), .ZN(new_n1092));
  OAI21_X1  g0892(.A(new_n710), .B1(new_n1087), .B2(new_n1092), .ZN(new_n1093));
  INV_X1    g0893(.A(new_n780), .ZN(new_n1094));
  OAI211_X1 g0894(.A(new_n1093), .B(new_n722), .C1(new_n505), .C2(new_n1094), .ZN(new_n1095));
  XOR2_X1   g0895(.A(new_n1095), .B(KEYINPUT116), .Z(new_n1096));
  NAND2_X1  g0896(.A1(new_n1075), .A2(new_n1096), .ZN(new_n1097));
  INV_X1    g0897(.A(new_n1097), .ZN(new_n1098));
  OAI21_X1  g0898(.A(new_n1069), .B1(new_n1070), .B2(new_n1098), .ZN(new_n1099));
  OAI21_X1  g0899(.A(new_n956), .B1(new_n1058), .B2(new_n1062), .ZN(new_n1100));
  NAND3_X1  g0900(.A1(new_n1100), .A2(KEYINPUT117), .A3(new_n1097), .ZN(new_n1101));
  AND3_X1   g0901(.A1(new_n1099), .A2(new_n1101), .A3(KEYINPUT118), .ZN(new_n1102));
  AOI21_X1  g0902(.A(KEYINPUT118), .B1(new_n1099), .B2(new_n1101), .ZN(new_n1103));
  OAI21_X1  g0903(.A(new_n1068), .B1(new_n1102), .B2(new_n1103), .ZN(G378));
  XOR2_X1   g0904(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1105));
  XNOR2_X1  g0905(.A(new_n598), .B(new_n1105), .ZN(new_n1106));
  NAND2_X1  g0906(.A1(new_n589), .A2(new_n833), .ZN(new_n1107));
  XNOR2_X1  g0907(.A(new_n1106), .B(new_n1107), .ZN(new_n1108));
  INV_X1    g0908(.A(new_n1108), .ZN(new_n1109));
  NAND2_X1  g0909(.A1(new_n873), .A2(new_n1109), .ZN(new_n1110));
  INV_X1    g0910(.A(KEYINPUT121), .ZN(new_n1111));
  NAND2_X1  g0911(.A1(new_n1110), .A2(new_n1111), .ZN(new_n1112));
  NAND4_X1  g0912(.A1(new_n864), .A2(G330), .A3(new_n872), .A4(new_n1108), .ZN(new_n1113));
  AND2_X1   g0913(.A1(new_n896), .A2(new_n1113), .ZN(new_n1114));
  NOR2_X1   g0914(.A1(new_n896), .A2(new_n1113), .ZN(new_n1115));
  OAI21_X1  g0915(.A(new_n1112), .B1(new_n1114), .B2(new_n1115), .ZN(new_n1116));
  INV_X1    g0916(.A(new_n1113), .ZN(new_n1117));
  INV_X1    g0917(.A(new_n885), .ZN(new_n1118));
  OAI21_X1  g0918(.A(new_n1118), .B1(new_n1074), .B2(new_n894), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n1117), .A2(new_n1119), .ZN(new_n1120));
  NAND2_X1  g0920(.A1(new_n896), .A2(new_n1113), .ZN(new_n1121));
  AOI21_X1  g0921(.A(KEYINPUT121), .B1(new_n873), .B2(new_n1109), .ZN(new_n1122));
  NAND3_X1  g0922(.A1(new_n1120), .A2(new_n1121), .A3(new_n1122), .ZN(new_n1123));
  NAND3_X1  g0923(.A1(new_n1116), .A2(new_n956), .A3(new_n1123), .ZN(new_n1124));
  OAI21_X1  g0924(.A(new_n250), .B1(new_n789), .B2(new_n296), .ZN(new_n1125));
  AOI21_X1  g0925(.A(new_n993), .B1(new_n432), .B2(new_n959), .ZN(new_n1126));
  OAI221_X1 g0926(.A(new_n1126), .B1(new_n284), .B2(new_n763), .C1(new_n333), .C2(new_n729), .ZN(new_n1127));
  AOI211_X1 g0927(.A(new_n1125), .B(new_n1127), .C1(G68), .C2(new_n757), .ZN(new_n1128));
  OAI21_X1  g0928(.A(new_n1128), .B1(new_n768), .B2(new_n746), .ZN(new_n1129));
  NOR2_X1   g0929(.A1(new_n752), .A2(new_n723), .ZN(new_n1130));
  NOR3_X1   g0930(.A1(new_n1129), .A2(new_n317), .A3(new_n1130), .ZN(new_n1131));
  XOR2_X1   g0931(.A(KEYINPUT119), .B(KEYINPUT58), .Z(new_n1132));
  XNOR2_X1  g0932(.A(new_n1131), .B(new_n1132), .ZN(new_n1133));
  OAI21_X1  g0933(.A(new_n219), .B1(new_n256), .B2(G41), .ZN(new_n1134));
  AOI21_X1  g0934(.A(G33), .B1(new_n753), .B2(G159), .ZN(new_n1135));
  NAND2_X1  g0935(.A1(new_n747), .A2(G124), .ZN(new_n1136));
  NAND3_X1  g0936(.A1(new_n1135), .A2(new_n250), .A3(new_n1136), .ZN(new_n1137));
  XOR2_X1   g0937(.A(new_n1137), .B(KEYINPUT120), .Z(new_n1138));
  NOR2_X1   g0938(.A1(new_n756), .A2(new_n586), .ZN(new_n1139));
  INV_X1    g0939(.A(G132), .ZN(new_n1140));
  OAI22_X1  g0940(.A1(new_n763), .A2(new_n1140), .B1(new_n788), .B2(new_n731), .ZN(new_n1141));
  AOI211_X1 g0941(.A(new_n1139), .B(new_n1141), .C1(new_n793), .C2(new_n1078), .ZN(new_n1142));
  OAI21_X1  g0942(.A(new_n1142), .B1(new_n1080), .B2(new_n789), .ZN(new_n1143));
  AOI21_X1  g0943(.A(new_n1143), .B1(G128), .B2(new_n786), .ZN(new_n1144));
  XOR2_X1   g0944(.A(new_n1144), .B(KEYINPUT59), .Z(new_n1145));
  OAI211_X1 g0945(.A(new_n1133), .B(new_n1134), .C1(new_n1138), .C2(new_n1145), .ZN(new_n1146));
  AOI22_X1  g0946(.A1(new_n1146), .A2(new_n710), .B1(new_n219), .B2(new_n780), .ZN(new_n1147));
  OAI211_X1 g0947(.A(new_n1147), .B(new_n722), .C1(new_n702), .C2(new_n1108), .ZN(new_n1148));
  AND2_X1   g0948(.A1(new_n1124), .A2(new_n1148), .ZN(new_n1149));
  AOI21_X1  g0949(.A(new_n1066), .B1(new_n1065), .B2(new_n1061), .ZN(new_n1150));
  INV_X1    g0950(.A(new_n1041), .ZN(new_n1151));
  OAI211_X1 g0951(.A(new_n1116), .B(new_n1123), .C1(new_n1150), .C2(new_n1151), .ZN(new_n1152));
  INV_X1    g0952(.A(KEYINPUT57), .ZN(new_n1153));
  OAI21_X1  g0953(.A(new_n663), .B1(new_n1152), .B2(new_n1153), .ZN(new_n1154));
  AND3_X1   g0954(.A1(new_n1120), .A2(new_n1121), .A3(new_n1122), .ZN(new_n1155));
  AOI21_X1  g0955(.A(new_n1122), .B1(new_n1120), .B2(new_n1121), .ZN(new_n1156));
  NOR2_X1   g0956(.A1(new_n1155), .A2(new_n1156), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n1063), .A2(new_n1041), .ZN(new_n1158));
  AOI21_X1  g0958(.A(KEYINPUT57), .B1(new_n1157), .B2(new_n1158), .ZN(new_n1159));
  OAI21_X1  g0959(.A(new_n1149), .B1(new_n1154), .B2(new_n1159), .ZN(G375));
  OR2_X1    g0960(.A1(new_n1052), .A2(new_n1041), .ZN(new_n1161));
  XOR2_X1   g0961(.A(new_n933), .B(KEYINPUT122), .Z(new_n1162));
  INV_X1    g0962(.A(new_n1162), .ZN(new_n1163));
  NAND3_X1  g0963(.A1(new_n1161), .A2(new_n1066), .A3(new_n1163), .ZN(new_n1164));
  NOR2_X1   g0964(.A1(new_n828), .A2(new_n702), .ZN(new_n1165));
  NOR2_X1   g0965(.A1(new_n1094), .A2(G68), .ZN(new_n1166));
  AOI22_X1  g0966(.A1(new_n786), .A2(G137), .B1(new_n734), .B2(new_n1078), .ZN(new_n1167));
  OAI21_X1  g0967(.A(new_n1167), .B1(new_n1140), .B2(new_n789), .ZN(new_n1168));
  XOR2_X1   g0968(.A(new_n1168), .B(KEYINPUT124), .Z(new_n1169));
  AOI211_X1 g0969(.A(new_n1130), .B(new_n1169), .C1(G159), .C2(new_n793), .ZN(new_n1170));
  NAND2_X1  g0970(.A1(new_n747), .A2(G128), .ZN(new_n1171));
  NAND2_X1  g0971(.A1(new_n959), .A2(G150), .ZN(new_n1172));
  AOI21_X1  g0972(.A(new_n538), .B1(new_n757), .B2(G50), .ZN(new_n1173));
  NAND4_X1  g0973(.A1(new_n1170), .A2(new_n1171), .A3(new_n1172), .A4(new_n1173), .ZN(new_n1174));
  OAI21_X1  g0974(.A(new_n995), .B1(new_n768), .B2(new_n729), .ZN(new_n1175));
  XNOR2_X1  g0975(.A(new_n1175), .B(KEYINPUT123), .ZN(new_n1176));
  OAI22_X1  g0976(.A1(new_n741), .A2(new_n284), .B1(new_n762), .B2(new_n789), .ZN(new_n1177));
  OAI221_X1 g0977(.A(new_n538), .B1(new_n210), .B2(new_n752), .C1(new_n763), .C2(new_n296), .ZN(new_n1178));
  NOR3_X1   g0978(.A1(new_n1176), .A2(new_n1177), .A3(new_n1178), .ZN(new_n1179));
  OAI221_X1 g0979(.A(new_n1179), .B1(new_n333), .B2(new_n731), .C1(new_n261), .C2(new_n746), .ZN(new_n1180));
  AOI22_X1  g0980(.A1(new_n1174), .A2(new_n1180), .B1(new_n708), .B2(new_n709), .ZN(new_n1181));
  NOR4_X1   g0981(.A1(new_n1165), .A2(new_n815), .A3(new_n1166), .A4(new_n1181), .ZN(new_n1182));
  AOI21_X1  g0982(.A(new_n1182), .B1(new_n1052), .B2(new_n956), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n1164), .A2(new_n1183), .ZN(G381));
  NOR2_X1   g0984(.A1(G387), .A2(G390), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n1185), .A2(new_n816), .ZN(new_n1186));
  NOR4_X1   g0986(.A1(new_n1186), .A2(G396), .A3(G393), .A4(G381), .ZN(new_n1187));
  INV_X1    g0987(.A(G375), .ZN(new_n1188));
  INV_X1    g0988(.A(new_n1068), .ZN(new_n1189));
  AOI21_X1  g0989(.A(KEYINPUT117), .B1(new_n1100), .B2(new_n1097), .ZN(new_n1190));
  NOR3_X1   g0990(.A1(new_n1070), .A2(new_n1069), .A3(new_n1098), .ZN(new_n1191));
  NOR3_X1   g0991(.A1(new_n1189), .A2(new_n1190), .A3(new_n1191), .ZN(new_n1192));
  NAND3_X1  g0992(.A1(new_n1187), .A2(new_n1188), .A3(new_n1192), .ZN(G407));
  NOR2_X1   g0993(.A1(new_n1187), .A2(new_n637), .ZN(new_n1194));
  NAND2_X1  g0994(.A1(new_n1188), .A2(new_n1192), .ZN(new_n1195));
  OAI21_X1  g0995(.A(G213), .B1(new_n1194), .B2(new_n1195), .ZN(G409));
  INV_X1    g0996(.A(KEYINPUT126), .ZN(new_n1197));
  INV_X1    g0997(.A(G213), .ZN(new_n1198));
  NOR2_X1   g0998(.A1(new_n1198), .A2(G343), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n1199), .A2(G2897), .ZN(new_n1200));
  INV_X1    g1000(.A(new_n1200), .ZN(new_n1201));
  INV_X1    g1001(.A(KEYINPUT60), .ZN(new_n1202));
  AOI21_X1  g1002(.A(new_n664), .B1(new_n1161), .B2(new_n1202), .ZN(new_n1203));
  NAND4_X1  g1003(.A1(new_n1151), .A2(KEYINPUT60), .A3(new_n1047), .A4(new_n1051), .ZN(new_n1204));
  NAND3_X1  g1004(.A1(new_n1203), .A2(new_n1066), .A3(new_n1204), .ZN(new_n1205));
  NAND3_X1  g1005(.A1(new_n1205), .A2(G384), .A3(new_n1183), .ZN(new_n1206));
  INV_X1    g1006(.A(new_n1206), .ZN(new_n1207));
  AOI21_X1  g1007(.A(G384), .B1(new_n1205), .B2(new_n1183), .ZN(new_n1208));
  OAI21_X1  g1008(.A(new_n1201), .B1(new_n1207), .B2(new_n1208), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(new_n1205), .A2(new_n1183), .ZN(new_n1210));
  NAND2_X1  g1010(.A1(new_n1210), .A2(new_n816), .ZN(new_n1211));
  NAND3_X1  g1011(.A1(new_n1211), .A2(new_n1206), .A3(new_n1200), .ZN(new_n1212));
  NAND2_X1  g1012(.A1(new_n1209), .A2(new_n1212), .ZN(new_n1213));
  OAI211_X1 g1013(.A(new_n1124), .B(new_n1148), .C1(new_n1152), .C2(new_n1162), .ZN(new_n1214));
  NAND2_X1  g1014(.A1(new_n1192), .A2(new_n1214), .ZN(new_n1215));
  INV_X1    g1015(.A(KEYINPUT118), .ZN(new_n1216));
  OAI21_X1  g1016(.A(new_n1216), .B1(new_n1190), .B2(new_n1191), .ZN(new_n1217));
  NAND3_X1  g1017(.A1(new_n1099), .A2(new_n1101), .A3(KEYINPUT118), .ZN(new_n1218));
  AOI21_X1  g1018(.A(new_n1189), .B1(new_n1217), .B2(new_n1218), .ZN(new_n1219));
  OAI21_X1  g1019(.A(new_n1215), .B1(G375), .B2(new_n1219), .ZN(new_n1220));
  INV_X1    g1020(.A(new_n1199), .ZN(new_n1221));
  AOI21_X1  g1021(.A(new_n1213), .B1(new_n1220), .B2(new_n1221), .ZN(new_n1222));
  OAI21_X1  g1022(.A(new_n1197), .B1(new_n1222), .B2(KEYINPUT61), .ZN(new_n1223));
  INV_X1    g1023(.A(KEYINPUT61), .ZN(new_n1224));
  NAND3_X1  g1024(.A1(new_n1157), .A2(KEYINPUT57), .A3(new_n1158), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(new_n1152), .A2(new_n1153), .ZN(new_n1226));
  NAND3_X1  g1026(.A1(new_n1225), .A2(new_n1226), .A3(new_n663), .ZN(new_n1227));
  NAND3_X1  g1027(.A1(G378), .A2(new_n1149), .A3(new_n1227), .ZN(new_n1228));
  AOI21_X1  g1028(.A(new_n1199), .B1(new_n1228), .B2(new_n1215), .ZN(new_n1229));
  OAI211_X1 g1029(.A(KEYINPUT126), .B(new_n1224), .C1(new_n1229), .C2(new_n1213), .ZN(new_n1230));
  NOR2_X1   g1030(.A1(new_n1207), .A2(new_n1208), .ZN(new_n1231));
  NAND3_X1  g1031(.A1(new_n1220), .A2(new_n1221), .A3(new_n1231), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(new_n1232), .A2(KEYINPUT62), .ZN(new_n1233));
  INV_X1    g1033(.A(KEYINPUT62), .ZN(new_n1234));
  NAND3_X1  g1034(.A1(new_n1229), .A2(new_n1234), .A3(new_n1231), .ZN(new_n1235));
  NAND4_X1  g1035(.A1(new_n1223), .A2(new_n1230), .A3(new_n1233), .A4(new_n1235), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(G387), .A2(G390), .ZN(new_n1237));
  INV_X1    g1037(.A(new_n1037), .ZN(new_n1238));
  INV_X1    g1038(.A(new_n1038), .ZN(new_n1239));
  INV_X1    g1039(.A(new_n1039), .ZN(new_n1240));
  AOI21_X1  g1040(.A(new_n1238), .B1(new_n1239), .B2(new_n1240), .ZN(new_n1241));
  NAND4_X1  g1041(.A1(new_n1241), .A2(new_n957), .A3(new_n981), .A4(new_n1015), .ZN(new_n1242));
  AOI21_X1  g1042(.A(KEYINPUT125), .B1(new_n1237), .B2(new_n1242), .ZN(new_n1243));
  XNOR2_X1  g1043(.A(G393), .B(G396), .ZN(new_n1244));
  NOR2_X1   g1044(.A1(new_n1243), .A2(new_n1244), .ZN(new_n1245));
  INV_X1    g1045(.A(KEYINPUT125), .ZN(new_n1246));
  AOI22_X1  g1046(.A1(new_n1241), .A2(new_n1015), .B1(new_n957), .B2(new_n981), .ZN(new_n1247));
  OAI21_X1  g1047(.A(new_n1246), .B1(new_n1185), .B2(new_n1247), .ZN(new_n1248));
  NAND3_X1  g1048(.A1(new_n1237), .A2(KEYINPUT125), .A3(new_n1242), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n1248), .A2(new_n1249), .ZN(new_n1250));
  AOI21_X1  g1050(.A(new_n1245), .B1(new_n1250), .B2(new_n1244), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n1236), .A2(new_n1251), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(new_n1250), .A2(new_n1244), .ZN(new_n1253));
  INV_X1    g1053(.A(new_n1245), .ZN(new_n1254));
  NAND2_X1  g1054(.A1(new_n1253), .A2(new_n1254), .ZN(new_n1255));
  NAND3_X1  g1055(.A1(new_n1229), .A2(KEYINPUT63), .A3(new_n1231), .ZN(new_n1256));
  INV_X1    g1056(.A(KEYINPUT63), .ZN(new_n1257));
  OAI21_X1  g1057(.A(new_n1232), .B1(new_n1222), .B2(new_n1257), .ZN(new_n1258));
  NAND4_X1  g1058(.A1(new_n1255), .A2(new_n1224), .A3(new_n1256), .A4(new_n1258), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(new_n1252), .A2(new_n1259), .ZN(G405));
  INV_X1    g1060(.A(new_n1228), .ZN(new_n1261));
  AND2_X1   g1061(.A1(G375), .A2(new_n1192), .ZN(new_n1262));
  OR3_X1    g1062(.A1(new_n1261), .A2(new_n1262), .A3(new_n1231), .ZN(new_n1263));
  OAI21_X1  g1063(.A(new_n1231), .B1(new_n1261), .B2(new_n1262), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(new_n1263), .A2(new_n1264), .ZN(new_n1265));
  XNOR2_X1  g1065(.A(new_n1265), .B(new_n1251), .ZN(G402));
endmodule


