//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 1 1 1 1 0 0 0 0 0 0 1 0 1 1 1 1 0 1 0 0 1 1 1 0 0 0 1 1 0 0 0 1 0 0 1 1 0 1 1 1 1 1 1 0 0 0 0 1 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:34:17 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n447, new_n449, new_n452, new_n453, new_n454, new_n455,
    new_n458, new_n459, new_n460, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n524, new_n525, new_n526,
    new_n527, new_n528, new_n529, new_n530, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n538, new_n539, new_n540, new_n541, new_n542,
    new_n545, new_n546, new_n548, new_n549, new_n550, new_n551, new_n552,
    new_n553, new_n554, new_n555, new_n556, new_n557, new_n558, new_n559,
    new_n560, new_n561, new_n565, new_n566, new_n567, new_n569, new_n570,
    new_n571, new_n572, new_n573, new_n574, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n596, new_n597, new_n600, new_n602, new_n603, new_n604, new_n605,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n824,
    new_n825, new_n826, new_n827, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n898,
    new_n899, new_n900, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1125, new_n1126;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  XOR2_X1   g002(.A(KEYINPUT64), .B(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  XOR2_X1   g012(.A(KEYINPUT65), .B(G69), .Z(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  XOR2_X1   g015(.A(KEYINPUT66), .B(G108), .Z(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  XNOR2_X1  g020(.A(KEYINPUT67), .B(KEYINPUT1), .ZN(new_n446));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XNOR2_X1  g022(.A(new_n446), .B(new_n447), .ZN(G223));
  INV_X1    g023(.A(new_n447), .ZN(new_n449));
  NAND2_X1  g024(.A1(new_n449), .A2(G567), .ZN(G234));
  NAND2_X1  g025(.A1(new_n449), .A2(G2106), .ZN(G217));
  NOR4_X1   g026(.A1(G238), .A2(G235), .A3(G237), .A4(G236), .ZN(new_n452));
  XOR2_X1   g027(.A(new_n452), .B(KEYINPUT68), .Z(new_n453));
  NOR4_X1   g028(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n454));
  XOR2_X1   g029(.A(new_n454), .B(KEYINPUT2), .Z(new_n455));
  NOR2_X1   g030(.A1(new_n453), .A2(new_n455), .ZN(G325));
  INV_X1    g031(.A(G325), .ZN(G261));
  NAND2_X1  g032(.A1(new_n453), .A2(G567), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n455), .A2(G2106), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  INV_X1    g035(.A(new_n460), .ZN(G319));
  INV_X1    g036(.A(G2105), .ZN(new_n462));
  AND2_X1   g037(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n463));
  NOR2_X1   g038(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n464));
  OAI21_X1  g039(.A(KEYINPUT69), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  INV_X1    g040(.A(KEYINPUT3), .ZN(new_n466));
  INV_X1    g041(.A(G2104), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  INV_X1    g043(.A(KEYINPUT69), .ZN(new_n469));
  NAND2_X1  g044(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n470));
  NAND3_X1  g045(.A1(new_n468), .A2(new_n469), .A3(new_n470), .ZN(new_n471));
  NAND3_X1  g046(.A1(new_n465), .A2(new_n471), .A3(G125), .ZN(new_n472));
  NAND2_X1  g047(.A1(G113), .A2(G2104), .ZN(new_n473));
  AOI21_X1  g048(.A(new_n462), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n462), .A2(G2104), .ZN(new_n475));
  INV_X1    g050(.A(new_n475), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n476), .A2(G101), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n468), .A2(new_n470), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n478), .A2(new_n462), .ZN(new_n479));
  INV_X1    g054(.A(G137), .ZN(new_n480));
  OAI21_X1  g055(.A(new_n477), .B1(new_n479), .B2(new_n480), .ZN(new_n481));
  NOR2_X1   g056(.A1(new_n474), .A2(new_n481), .ZN(G160));
  AOI21_X1  g057(.A(new_n462), .B1(new_n468), .B2(new_n470), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n483), .A2(G124), .ZN(new_n484));
  NOR2_X1   g059(.A1(new_n462), .A2(G112), .ZN(new_n485));
  OAI21_X1  g060(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n486));
  OAI21_X1  g061(.A(new_n484), .B1(new_n485), .B2(new_n486), .ZN(new_n487));
  INV_X1    g062(.A(new_n479), .ZN(new_n488));
  AOI21_X1  g063(.A(new_n487), .B1(G136), .B2(new_n488), .ZN(new_n489));
  XNOR2_X1  g064(.A(new_n489), .B(KEYINPUT70), .ZN(G162));
  INV_X1    g065(.A(G138), .ZN(new_n491));
  NOR3_X1   g066(.A1(new_n491), .A2(KEYINPUT4), .A3(G2105), .ZN(new_n492));
  NAND3_X1  g067(.A1(new_n465), .A2(new_n471), .A3(new_n492), .ZN(new_n493));
  INV_X1    g068(.A(KEYINPUT71), .ZN(new_n494));
  NAND2_X1  g069(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  NAND4_X1  g070(.A1(new_n465), .A2(new_n471), .A3(KEYINPUT71), .A4(new_n492), .ZN(new_n496));
  NAND3_X1  g071(.A1(new_n478), .A2(G138), .A3(new_n462), .ZN(new_n497));
  NAND2_X1  g072(.A1(new_n497), .A2(KEYINPUT4), .ZN(new_n498));
  NAND3_X1  g073(.A1(new_n495), .A2(new_n496), .A3(new_n498), .ZN(new_n499));
  OAI21_X1  g074(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n500));
  INV_X1    g075(.A(G114), .ZN(new_n501));
  AOI21_X1  g076(.A(new_n500), .B1(new_n501), .B2(G2105), .ZN(new_n502));
  AOI21_X1  g077(.A(new_n502), .B1(new_n483), .B2(G126), .ZN(new_n503));
  AND3_X1   g078(.A1(new_n499), .A2(KEYINPUT72), .A3(new_n503), .ZN(new_n504));
  AOI21_X1  g079(.A(KEYINPUT72), .B1(new_n499), .B2(new_n503), .ZN(new_n505));
  NOR2_X1   g080(.A1(new_n504), .A2(new_n505), .ZN(G164));
  OR2_X1    g081(.A1(KEYINPUT5), .A2(G543), .ZN(new_n507));
  NAND2_X1  g082(.A1(KEYINPUT5), .A2(G543), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  AOI22_X1  g084(.A1(new_n509), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n510));
  INV_X1    g085(.A(G651), .ZN(new_n511));
  NOR2_X1   g086(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  INV_X1    g087(.A(G543), .ZN(new_n513));
  OR2_X1    g088(.A1(KEYINPUT6), .A2(G651), .ZN(new_n514));
  NAND2_X1  g089(.A1(KEYINPUT6), .A2(G651), .ZN(new_n515));
  AOI21_X1  g090(.A(new_n513), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n516), .A2(G50), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n514), .A2(new_n515), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n518), .A2(new_n509), .ZN(new_n519));
  INV_X1    g094(.A(G88), .ZN(new_n520));
  OAI21_X1  g095(.A(new_n517), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  OR2_X1    g096(.A1(new_n512), .A2(new_n521), .ZN(G303));
  INV_X1    g097(.A(G303), .ZN(G166));
  NAND3_X1  g098(.A1(new_n509), .A2(G63), .A3(G651), .ZN(new_n524));
  XOR2_X1   g099(.A(new_n524), .B(KEYINPUT73), .Z(new_n525));
  NAND2_X1  g100(.A1(new_n516), .A2(G51), .ZN(new_n526));
  NAND3_X1  g101(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n527));
  XNOR2_X1  g102(.A(new_n527), .B(KEYINPUT7), .ZN(new_n528));
  XNOR2_X1  g103(.A(KEYINPUT74), .B(G89), .ZN(new_n529));
  OAI211_X1 g104(.A(new_n526), .B(new_n528), .C1(new_n519), .C2(new_n529), .ZN(new_n530));
  NOR2_X1   g105(.A1(new_n525), .A2(new_n530), .ZN(G168));
  AOI22_X1  g106(.A1(new_n509), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n532));
  NOR2_X1   g107(.A1(new_n532), .A2(new_n511), .ZN(new_n533));
  NAND2_X1  g108(.A1(new_n516), .A2(G52), .ZN(new_n534));
  INV_X1    g109(.A(G90), .ZN(new_n535));
  OAI21_X1  g110(.A(new_n534), .B1(new_n519), .B2(new_n535), .ZN(new_n536));
  NOR2_X1   g111(.A1(new_n533), .A2(new_n536), .ZN(G171));
  AOI22_X1  g112(.A1(new_n509), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n538));
  OR2_X1    g113(.A1(new_n538), .A2(new_n511), .ZN(new_n539));
  AND2_X1   g114(.A1(new_n518), .A2(new_n509), .ZN(new_n540));
  AOI22_X1  g115(.A1(new_n540), .A2(G81), .B1(G43), .B2(new_n516), .ZN(new_n541));
  AND2_X1   g116(.A1(new_n539), .A2(new_n541), .ZN(new_n542));
  NAND2_X1  g117(.A1(new_n542), .A2(G860), .ZN(G153));
  NAND4_X1  g118(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g119(.A1(G1), .A2(G3), .ZN(new_n545));
  XNOR2_X1  g120(.A(new_n545), .B(KEYINPUT8), .ZN(new_n546));
  NAND4_X1  g121(.A1(G319), .A2(G483), .A3(G661), .A4(new_n546), .ZN(G188));
  INV_X1    g122(.A(G65), .ZN(new_n548));
  AOI21_X1  g123(.A(new_n548), .B1(new_n507), .B2(new_n508), .ZN(new_n549));
  AND2_X1   g124(.A1(G78), .A2(G543), .ZN(new_n550));
  OAI21_X1  g125(.A(G651), .B1(new_n549), .B2(new_n550), .ZN(new_n551));
  AOI22_X1  g126(.A1(new_n551), .A2(KEYINPUT75), .B1(new_n540), .B2(G91), .ZN(new_n552));
  INV_X1    g127(.A(KEYINPUT9), .ZN(new_n553));
  NAND3_X1  g128(.A1(new_n516), .A2(new_n553), .A3(G53), .ZN(new_n554));
  AND2_X1   g129(.A1(KEYINPUT6), .A2(G651), .ZN(new_n555));
  NOR2_X1   g130(.A1(KEYINPUT6), .A2(G651), .ZN(new_n556));
  OAI211_X1 g131(.A(G53), .B(G543), .C1(new_n555), .C2(new_n556), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n557), .A2(KEYINPUT9), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n554), .A2(new_n558), .ZN(new_n559));
  INV_X1    g134(.A(KEYINPUT75), .ZN(new_n560));
  OAI211_X1 g135(.A(new_n560), .B(G651), .C1(new_n549), .C2(new_n550), .ZN(new_n561));
  NAND3_X1  g136(.A1(new_n552), .A2(new_n559), .A3(new_n561), .ZN(G299));
  INV_X1    g137(.A(G171), .ZN(G301));
  INV_X1    g138(.A(G168), .ZN(G286));
  NAND2_X1  g139(.A1(new_n540), .A2(G87), .ZN(new_n565));
  OAI21_X1  g140(.A(G651), .B1(new_n509), .B2(G74), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n516), .A2(G49), .ZN(new_n567));
  NAND3_X1  g142(.A1(new_n565), .A2(new_n566), .A3(new_n567), .ZN(G288));
  AOI22_X1  g143(.A1(new_n509), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n569));
  NOR2_X1   g144(.A1(new_n569), .A2(new_n511), .ZN(new_n570));
  NAND2_X1  g145(.A1(new_n516), .A2(G48), .ZN(new_n571));
  INV_X1    g146(.A(G86), .ZN(new_n572));
  OAI21_X1  g147(.A(new_n571), .B1(new_n519), .B2(new_n572), .ZN(new_n573));
  NOR2_X1   g148(.A1(new_n570), .A2(new_n573), .ZN(new_n574));
  INV_X1    g149(.A(new_n574), .ZN(G305));
  AND2_X1   g150(.A1(new_n509), .A2(G60), .ZN(new_n576));
  AND2_X1   g151(.A1(G72), .A2(G543), .ZN(new_n577));
  OAI21_X1  g152(.A(G651), .B1(new_n576), .B2(new_n577), .ZN(new_n578));
  INV_X1    g153(.A(KEYINPUT76), .ZN(new_n579));
  NAND2_X1  g154(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  AOI22_X1  g155(.A1(new_n540), .A2(G85), .B1(G47), .B2(new_n516), .ZN(new_n581));
  AND2_X1   g156(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  OR2_X1    g157(.A1(new_n578), .A2(new_n579), .ZN(new_n583));
  NAND2_X1  g158(.A1(new_n582), .A2(new_n583), .ZN(G290));
  NAND2_X1  g159(.A1(G301), .A2(G868), .ZN(new_n585));
  AND3_X1   g160(.A1(new_n518), .A2(new_n509), .A3(G92), .ZN(new_n586));
  XNOR2_X1  g161(.A(new_n586), .B(KEYINPUT10), .ZN(new_n587));
  NAND2_X1  g162(.A1(new_n509), .A2(G66), .ZN(new_n588));
  INV_X1    g163(.A(G79), .ZN(new_n589));
  OAI21_X1  g164(.A(new_n588), .B1(new_n589), .B2(new_n513), .ZN(new_n590));
  AOI22_X1  g165(.A1(new_n590), .A2(G651), .B1(G54), .B2(new_n516), .ZN(new_n591));
  NAND2_X1  g166(.A1(new_n587), .A2(new_n591), .ZN(new_n592));
  INV_X1    g167(.A(new_n592), .ZN(new_n593));
  OAI21_X1  g168(.A(new_n585), .B1(new_n593), .B2(G868), .ZN(G284));
  OAI21_X1  g169(.A(new_n585), .B1(new_n593), .B2(G868), .ZN(G321));
  INV_X1    g170(.A(G868), .ZN(new_n596));
  NAND2_X1  g171(.A1(G299), .A2(new_n596), .ZN(new_n597));
  OAI21_X1  g172(.A(new_n597), .B1(G168), .B2(new_n596), .ZN(G297));
  OAI21_X1  g173(.A(new_n597), .B1(G168), .B2(new_n596), .ZN(G280));
  INV_X1    g174(.A(G559), .ZN(new_n600));
  OAI21_X1  g175(.A(new_n593), .B1(new_n600), .B2(G860), .ZN(G148));
  NAND2_X1  g176(.A1(new_n593), .A2(new_n600), .ZN(new_n602));
  NAND2_X1  g177(.A1(new_n602), .A2(G868), .ZN(new_n603));
  OR2_X1    g178(.A1(new_n603), .A2(KEYINPUT77), .ZN(new_n604));
  NAND2_X1  g179(.A1(new_n603), .A2(KEYINPUT77), .ZN(new_n605));
  OAI211_X1 g180(.A(new_n604), .B(new_n605), .C1(G868), .C2(new_n542), .ZN(G323));
  XNOR2_X1  g181(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g182(.A1(new_n465), .A2(new_n471), .ZN(new_n608));
  NOR2_X1   g183(.A1(new_n608), .A2(new_n475), .ZN(new_n609));
  XNOR2_X1  g184(.A(KEYINPUT78), .B(KEYINPUT12), .ZN(new_n610));
  XNOR2_X1  g185(.A(new_n609), .B(new_n610), .ZN(new_n611));
  XNOR2_X1  g186(.A(new_n611), .B(KEYINPUT13), .ZN(new_n612));
  OR2_X1    g187(.A1(new_n612), .A2(G2100), .ZN(new_n613));
  NAND2_X1  g188(.A1(new_n612), .A2(G2100), .ZN(new_n614));
  NAND2_X1  g189(.A1(new_n483), .A2(G123), .ZN(new_n615));
  NOR2_X1   g190(.A1(new_n462), .A2(G111), .ZN(new_n616));
  OAI21_X1  g191(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n617));
  INV_X1    g192(.A(G135), .ZN(new_n618));
  OAI221_X1 g193(.A(new_n615), .B1(new_n616), .B2(new_n617), .C1(new_n618), .C2(new_n479), .ZN(new_n619));
  XOR2_X1   g194(.A(new_n619), .B(G2096), .Z(new_n620));
  NAND3_X1  g195(.A1(new_n613), .A2(new_n614), .A3(new_n620), .ZN(G156));
  INV_X1    g196(.A(G14), .ZN(new_n622));
  XNOR2_X1  g197(.A(G2427), .B(G2438), .ZN(new_n623));
  XNOR2_X1  g198(.A(new_n623), .B(G2430), .ZN(new_n624));
  XNOR2_X1  g199(.A(KEYINPUT15), .B(G2435), .ZN(new_n625));
  OR2_X1    g200(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  NAND2_X1  g201(.A1(new_n624), .A2(new_n625), .ZN(new_n627));
  NAND3_X1  g202(.A1(new_n626), .A2(KEYINPUT14), .A3(new_n627), .ZN(new_n628));
  XNOR2_X1  g203(.A(G2443), .B(G2446), .ZN(new_n629));
  XNOR2_X1  g204(.A(new_n628), .B(new_n629), .ZN(new_n630));
  XOR2_X1   g205(.A(G2451), .B(G2454), .Z(new_n631));
  XNOR2_X1  g206(.A(new_n631), .B(KEYINPUT16), .ZN(new_n632));
  XNOR2_X1  g207(.A(new_n632), .B(KEYINPUT79), .ZN(new_n633));
  XNOR2_X1  g208(.A(new_n630), .B(new_n633), .ZN(new_n634));
  INV_X1    g209(.A(new_n634), .ZN(new_n635));
  XNOR2_X1  g210(.A(G1341), .B(G1348), .ZN(new_n636));
  NOR2_X1   g211(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  XNOR2_X1  g212(.A(new_n637), .B(KEYINPUT80), .ZN(new_n638));
  AOI211_X1 g213(.A(new_n622), .B(new_n638), .C1(new_n636), .C2(new_n635), .ZN(G401));
  XOR2_X1   g214(.A(KEYINPUT81), .B(KEYINPUT18), .Z(new_n640));
  XOR2_X1   g215(.A(G2084), .B(G2090), .Z(new_n641));
  XNOR2_X1  g216(.A(G2067), .B(G2678), .ZN(new_n642));
  NAND2_X1  g217(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  NAND2_X1  g218(.A1(new_n643), .A2(KEYINPUT17), .ZN(new_n644));
  NOR2_X1   g219(.A1(new_n641), .A2(new_n642), .ZN(new_n645));
  OAI21_X1  g220(.A(new_n640), .B1(new_n644), .B2(new_n645), .ZN(new_n646));
  XOR2_X1   g221(.A(G2072), .B(G2078), .Z(new_n647));
  INV_X1    g222(.A(new_n640), .ZN(new_n648));
  AOI21_X1  g223(.A(new_n647), .B1(new_n643), .B2(new_n648), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n646), .B(new_n649), .ZN(new_n650));
  XNOR2_X1  g225(.A(G2096), .B(G2100), .ZN(new_n651));
  XNOR2_X1  g226(.A(new_n650), .B(new_n651), .ZN(G227));
  XNOR2_X1  g227(.A(G1971), .B(G1976), .ZN(new_n653));
  XNOR2_X1  g228(.A(new_n653), .B(KEYINPUT19), .ZN(new_n654));
  INV_X1    g229(.A(KEYINPUT82), .ZN(new_n655));
  XNOR2_X1  g230(.A(G1956), .B(G2474), .ZN(new_n656));
  INV_X1    g231(.A(new_n656), .ZN(new_n657));
  XNOR2_X1  g232(.A(G1961), .B(G1966), .ZN(new_n658));
  INV_X1    g233(.A(new_n658), .ZN(new_n659));
  NAND2_X1  g234(.A1(new_n657), .A2(new_n659), .ZN(new_n660));
  AOI21_X1  g235(.A(new_n654), .B1(new_n655), .B2(new_n660), .ZN(new_n661));
  OAI21_X1  g236(.A(new_n661), .B1(new_n655), .B2(new_n660), .ZN(new_n662));
  XNOR2_X1  g237(.A(new_n662), .B(KEYINPUT20), .ZN(new_n663));
  NOR2_X1   g238(.A1(new_n657), .A2(new_n659), .ZN(new_n664));
  INV_X1    g239(.A(new_n664), .ZN(new_n665));
  NAND3_X1  g240(.A1(new_n665), .A2(new_n660), .A3(new_n654), .ZN(new_n666));
  OAI211_X1 g241(.A(new_n663), .B(new_n666), .C1(new_n654), .C2(new_n665), .ZN(new_n667));
  XNOR2_X1  g242(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n668));
  XNOR2_X1  g243(.A(new_n667), .B(new_n668), .ZN(new_n669));
  XNOR2_X1  g244(.A(G1991), .B(G1996), .ZN(new_n670));
  XNOR2_X1  g245(.A(new_n669), .B(new_n670), .ZN(new_n671));
  XNOR2_X1  g246(.A(G1981), .B(G1986), .ZN(new_n672));
  XNOR2_X1  g247(.A(new_n671), .B(new_n672), .ZN(G229));
  INV_X1    g248(.A(G16), .ZN(new_n674));
  NAND2_X1  g249(.A1(new_n674), .A2(G22), .ZN(new_n675));
  OAI21_X1  g250(.A(new_n675), .B1(G166), .B2(new_n674), .ZN(new_n676));
  XNOR2_X1  g251(.A(new_n676), .B(G1971), .ZN(new_n677));
  INV_X1    g252(.A(KEYINPUT83), .ZN(new_n678));
  OR2_X1    g253(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  NOR2_X1   g254(.A1(G6), .A2(G16), .ZN(new_n680));
  AOI21_X1  g255(.A(new_n680), .B1(new_n574), .B2(G16), .ZN(new_n681));
  XNOR2_X1  g256(.A(new_n681), .B(KEYINPUT32), .ZN(new_n682));
  INV_X1    g257(.A(G1981), .ZN(new_n683));
  XNOR2_X1  g258(.A(new_n682), .B(new_n683), .ZN(new_n684));
  NAND2_X1  g259(.A1(new_n677), .A2(new_n678), .ZN(new_n685));
  NAND2_X1  g260(.A1(new_n674), .A2(G23), .ZN(new_n686));
  INV_X1    g261(.A(G288), .ZN(new_n687));
  OAI21_X1  g262(.A(new_n686), .B1(new_n687), .B2(new_n674), .ZN(new_n688));
  XNOR2_X1  g263(.A(KEYINPUT33), .B(G1976), .ZN(new_n689));
  XNOR2_X1  g264(.A(new_n688), .B(new_n689), .ZN(new_n690));
  NAND4_X1  g265(.A1(new_n679), .A2(new_n684), .A3(new_n685), .A4(new_n690), .ZN(new_n691));
  OR2_X1    g266(.A1(new_n691), .A2(KEYINPUT34), .ZN(new_n692));
  NAND2_X1  g267(.A1(new_n691), .A2(KEYINPUT34), .ZN(new_n693));
  NAND2_X1  g268(.A1(new_n674), .A2(G24), .ZN(new_n694));
  INV_X1    g269(.A(G290), .ZN(new_n695));
  OAI21_X1  g270(.A(new_n694), .B1(new_n695), .B2(new_n674), .ZN(new_n696));
  INV_X1    g271(.A(G1986), .ZN(new_n697));
  XNOR2_X1  g272(.A(new_n696), .B(new_n697), .ZN(new_n698));
  NAND2_X1  g273(.A1(new_n483), .A2(G119), .ZN(new_n699));
  NOR2_X1   g274(.A1(new_n462), .A2(G107), .ZN(new_n700));
  OAI21_X1  g275(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n701));
  INV_X1    g276(.A(G131), .ZN(new_n702));
  OAI221_X1 g277(.A(new_n699), .B1(new_n700), .B2(new_n701), .C1(new_n702), .C2(new_n479), .ZN(new_n703));
  MUX2_X1   g278(.A(G25), .B(new_n703), .S(G29), .Z(new_n704));
  XOR2_X1   g279(.A(KEYINPUT35), .B(G1991), .Z(new_n705));
  XNOR2_X1  g280(.A(new_n704), .B(new_n705), .ZN(new_n706));
  NAND4_X1  g281(.A1(new_n692), .A2(new_n693), .A3(new_n698), .A4(new_n706), .ZN(new_n707));
  XOR2_X1   g282(.A(KEYINPUT84), .B(KEYINPUT36), .Z(new_n708));
  XNOR2_X1  g283(.A(new_n707), .B(new_n708), .ZN(new_n709));
  NAND2_X1  g284(.A1(new_n488), .A2(G141), .ZN(new_n710));
  XOR2_X1   g285(.A(new_n710), .B(KEYINPUT87), .Z(new_n711));
  NAND2_X1  g286(.A1(new_n483), .A2(G129), .ZN(new_n712));
  XNOR2_X1  g287(.A(new_n712), .B(KEYINPUT88), .ZN(new_n713));
  NAND3_X1  g288(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n714));
  INV_X1    g289(.A(KEYINPUT26), .ZN(new_n715));
  OR2_X1    g290(.A1(new_n714), .A2(new_n715), .ZN(new_n716));
  NAND2_X1  g291(.A1(new_n714), .A2(new_n715), .ZN(new_n717));
  AOI22_X1  g292(.A1(new_n716), .A2(new_n717), .B1(G105), .B2(new_n476), .ZN(new_n718));
  NAND3_X1  g293(.A1(new_n711), .A2(new_n713), .A3(new_n718), .ZN(new_n719));
  XNOR2_X1  g294(.A(new_n719), .B(KEYINPUT89), .ZN(new_n720));
  NAND2_X1  g295(.A1(new_n720), .A2(G29), .ZN(new_n721));
  OAI211_X1 g296(.A(new_n721), .B(KEYINPUT90), .C1(G29), .C2(G32), .ZN(new_n722));
  OAI21_X1  g297(.A(new_n722), .B1(KEYINPUT90), .B2(new_n721), .ZN(new_n723));
  XOR2_X1   g298(.A(KEYINPUT27), .B(G1996), .Z(new_n724));
  XNOR2_X1  g299(.A(new_n723), .B(new_n724), .ZN(new_n725));
  XOR2_X1   g300(.A(KEYINPUT31), .B(G11), .Z(new_n726));
  INV_X1    g301(.A(G29), .ZN(new_n727));
  INV_X1    g302(.A(KEYINPUT30), .ZN(new_n728));
  OAI21_X1  g303(.A(new_n727), .B1(new_n728), .B2(G28), .ZN(new_n729));
  NOR2_X1   g304(.A1(new_n729), .A2(KEYINPUT91), .ZN(new_n730));
  AOI21_X1  g305(.A(new_n730), .B1(new_n728), .B2(G28), .ZN(new_n731));
  NAND2_X1  g306(.A1(new_n729), .A2(KEYINPUT91), .ZN(new_n732));
  AOI21_X1  g307(.A(new_n726), .B1(new_n731), .B2(new_n732), .ZN(new_n733));
  NAND2_X1  g308(.A1(new_n542), .A2(G16), .ZN(new_n734));
  OAI21_X1  g309(.A(new_n734), .B1(G16), .B2(G19), .ZN(new_n735));
  INV_X1    g310(.A(G1341), .ZN(new_n736));
  OAI221_X1 g311(.A(new_n733), .B1(new_n727), .B2(new_n619), .C1(new_n735), .C2(new_n736), .ZN(new_n737));
  AOI21_X1  g312(.A(new_n737), .B1(new_n736), .B2(new_n735), .ZN(new_n738));
  NAND2_X1  g313(.A1(new_n727), .A2(G33), .ZN(new_n739));
  NAND3_X1  g314(.A1(new_n462), .A2(G103), .A3(G2104), .ZN(new_n740));
  XNOR2_X1  g315(.A(new_n740), .B(KEYINPUT25), .ZN(new_n741));
  INV_X1    g316(.A(new_n608), .ZN(new_n742));
  AOI22_X1  g317(.A1(new_n742), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n743));
  NOR2_X1   g318(.A1(new_n743), .A2(new_n462), .ZN(new_n744));
  AOI211_X1 g319(.A(new_n741), .B(new_n744), .C1(G139), .C2(new_n488), .ZN(new_n745));
  OAI21_X1  g320(.A(new_n739), .B1(new_n745), .B2(new_n727), .ZN(new_n746));
  OR2_X1    g321(.A1(new_n746), .A2(G2072), .ZN(new_n747));
  NAND2_X1  g322(.A1(new_n674), .A2(G21), .ZN(new_n748));
  OAI21_X1  g323(.A(new_n748), .B1(G168), .B2(new_n674), .ZN(new_n749));
  OR2_X1    g324(.A1(new_n749), .A2(G1966), .ZN(new_n750));
  NAND2_X1  g325(.A1(new_n727), .A2(G26), .ZN(new_n751));
  XNOR2_X1  g326(.A(new_n751), .B(KEYINPUT28), .ZN(new_n752));
  NAND2_X1  g327(.A1(new_n488), .A2(G140), .ZN(new_n753));
  NAND2_X1  g328(.A1(new_n483), .A2(G128), .ZN(new_n754));
  OR2_X1    g329(.A1(G104), .A2(G2105), .ZN(new_n755));
  OAI211_X1 g330(.A(new_n755), .B(G2104), .C1(G116), .C2(new_n462), .ZN(new_n756));
  NAND3_X1  g331(.A1(new_n753), .A2(new_n754), .A3(new_n756), .ZN(new_n757));
  INV_X1    g332(.A(new_n757), .ZN(new_n758));
  OAI21_X1  g333(.A(new_n752), .B1(new_n758), .B2(new_n727), .ZN(new_n759));
  XNOR2_X1  g334(.A(new_n759), .B(G2067), .ZN(new_n760));
  AOI21_X1  g335(.A(new_n760), .B1(new_n749), .B2(G1966), .ZN(new_n761));
  NAND4_X1  g336(.A1(new_n738), .A2(new_n747), .A3(new_n750), .A4(new_n761), .ZN(new_n762));
  NOR2_X1   g337(.A1(G5), .A2(G16), .ZN(new_n763));
  XOR2_X1   g338(.A(new_n763), .B(KEYINPUT92), .Z(new_n764));
  OAI21_X1  g339(.A(new_n764), .B1(G301), .B2(new_n674), .ZN(new_n765));
  XNOR2_X1  g340(.A(new_n765), .B(KEYINPUT93), .ZN(new_n766));
  INV_X1    g341(.A(G1961), .ZN(new_n767));
  OR2_X1    g342(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  INV_X1    g343(.A(G34), .ZN(new_n769));
  AOI21_X1  g344(.A(G29), .B1(new_n769), .B2(KEYINPUT24), .ZN(new_n770));
  OAI21_X1  g345(.A(new_n770), .B1(KEYINPUT24), .B2(new_n769), .ZN(new_n771));
  INV_X1    g346(.A(G160), .ZN(new_n772));
  OAI21_X1  g347(.A(new_n771), .B1(new_n772), .B2(new_n727), .ZN(new_n773));
  INV_X1    g348(.A(G2084), .ZN(new_n774));
  NAND2_X1  g349(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  NAND2_X1  g350(.A1(new_n766), .A2(new_n767), .ZN(new_n776));
  NAND2_X1  g351(.A1(new_n674), .A2(G4), .ZN(new_n777));
  OAI21_X1  g352(.A(new_n777), .B1(new_n593), .B2(new_n674), .ZN(new_n778));
  INV_X1    g353(.A(G1348), .ZN(new_n779));
  XNOR2_X1  g354(.A(new_n778), .B(new_n779), .ZN(new_n780));
  NAND4_X1  g355(.A1(new_n768), .A2(new_n775), .A3(new_n776), .A4(new_n780), .ZN(new_n781));
  NOR2_X1   g356(.A1(new_n762), .A2(new_n781), .ZN(new_n782));
  NAND2_X1  g357(.A1(new_n746), .A2(G2072), .ZN(new_n783));
  XOR2_X1   g358(.A(new_n783), .B(KEYINPUT86), .Z(new_n784));
  NOR2_X1   g359(.A1(new_n773), .A2(new_n774), .ZN(new_n785));
  XNOR2_X1  g360(.A(new_n785), .B(KEYINPUT85), .ZN(new_n786));
  NAND2_X1  g361(.A1(new_n727), .A2(G27), .ZN(new_n787));
  OAI21_X1  g362(.A(new_n787), .B1(G164), .B2(new_n727), .ZN(new_n788));
  INV_X1    g363(.A(G2078), .ZN(new_n789));
  XNOR2_X1  g364(.A(new_n788), .B(new_n789), .ZN(new_n790));
  NAND4_X1  g365(.A1(new_n782), .A2(new_n784), .A3(new_n786), .A4(new_n790), .ZN(new_n791));
  NAND2_X1  g366(.A1(G299), .A2(G16), .ZN(new_n792));
  XOR2_X1   g367(.A(KEYINPUT94), .B(KEYINPUT23), .Z(new_n793));
  NAND2_X1  g368(.A1(new_n674), .A2(G20), .ZN(new_n794));
  XNOR2_X1  g369(.A(new_n793), .B(new_n794), .ZN(new_n795));
  NAND2_X1  g370(.A1(new_n792), .A2(new_n795), .ZN(new_n796));
  XNOR2_X1  g371(.A(new_n796), .B(G1956), .ZN(new_n797));
  NOR2_X1   g372(.A1(G29), .A2(G35), .ZN(new_n798));
  AOI21_X1  g373(.A(new_n798), .B1(G162), .B2(G29), .ZN(new_n799));
  XNOR2_X1  g374(.A(new_n799), .B(KEYINPUT29), .ZN(new_n800));
  AOI21_X1  g375(.A(new_n797), .B1(new_n800), .B2(G2090), .ZN(new_n801));
  OAI21_X1  g376(.A(new_n801), .B1(G2090), .B2(new_n800), .ZN(new_n802));
  NOR3_X1   g377(.A1(new_n725), .A2(new_n791), .A3(new_n802), .ZN(new_n803));
  NAND2_X1  g378(.A1(new_n709), .A2(new_n803), .ZN(G150));
  INV_X1    g379(.A(G150), .ZN(G311));
  NAND2_X1  g380(.A1(new_n593), .A2(G559), .ZN(new_n806));
  XNOR2_X1  g381(.A(new_n806), .B(KEYINPUT38), .ZN(new_n807));
  AOI22_X1  g382(.A1(new_n509), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n808));
  NOR2_X1   g383(.A1(new_n808), .A2(new_n511), .ZN(new_n809));
  NAND2_X1  g384(.A1(new_n516), .A2(G55), .ZN(new_n810));
  XOR2_X1   g385(.A(KEYINPUT95), .B(G93), .Z(new_n811));
  OAI21_X1  g386(.A(new_n810), .B1(new_n519), .B2(new_n811), .ZN(new_n812));
  NOR2_X1   g387(.A1(new_n809), .A2(new_n812), .ZN(new_n813));
  XNOR2_X1  g388(.A(new_n542), .B(new_n813), .ZN(new_n814));
  XOR2_X1   g389(.A(new_n807), .B(new_n814), .Z(new_n815));
  AND2_X1   g390(.A1(new_n815), .A2(KEYINPUT39), .ZN(new_n816));
  NOR2_X1   g391(.A1(new_n815), .A2(KEYINPUT39), .ZN(new_n817));
  NOR3_X1   g392(.A1(new_n816), .A2(new_n817), .A3(G860), .ZN(new_n818));
  OAI21_X1  g393(.A(G860), .B1(new_n812), .B2(new_n809), .ZN(new_n819));
  XNOR2_X1  g394(.A(new_n819), .B(KEYINPUT97), .ZN(new_n820));
  XNOR2_X1  g395(.A(new_n820), .B(KEYINPUT96), .ZN(new_n821));
  XNOR2_X1  g396(.A(new_n821), .B(KEYINPUT37), .ZN(new_n822));
  OR2_X1    g397(.A1(new_n818), .A2(new_n822), .ZN(G145));
  MUX2_X1   g398(.A(new_n719), .B(new_n720), .S(new_n745), .Z(new_n824));
  NAND2_X1  g399(.A1(new_n499), .A2(new_n503), .ZN(new_n825));
  XNOR2_X1  g400(.A(new_n825), .B(new_n758), .ZN(new_n826));
  XOR2_X1   g401(.A(new_n824), .B(new_n826), .Z(new_n827));
  AOI22_X1  g402(.A1(new_n488), .A2(G142), .B1(G130), .B2(new_n483), .ZN(new_n828));
  OAI21_X1  g403(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n829));
  INV_X1    g404(.A(G118), .ZN(new_n830));
  AOI22_X1  g405(.A1(new_n829), .A2(KEYINPUT98), .B1(new_n830), .B2(G2105), .ZN(new_n831));
  OAI21_X1  g406(.A(new_n831), .B1(KEYINPUT98), .B2(new_n829), .ZN(new_n832));
  NAND2_X1  g407(.A1(new_n828), .A2(new_n832), .ZN(new_n833));
  XNOR2_X1  g408(.A(new_n833), .B(new_n703), .ZN(new_n834));
  XNOR2_X1  g409(.A(new_n834), .B(new_n611), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n827), .A2(new_n835), .ZN(new_n836));
  XNOR2_X1  g411(.A(new_n824), .B(new_n826), .ZN(new_n837));
  INV_X1    g412(.A(new_n835), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n837), .A2(new_n838), .ZN(new_n839));
  XNOR2_X1  g414(.A(G160), .B(new_n619), .ZN(new_n840));
  XNOR2_X1  g415(.A(G162), .B(new_n840), .ZN(new_n841));
  NAND3_X1  g416(.A1(new_n836), .A2(new_n839), .A3(new_n841), .ZN(new_n842));
  XNOR2_X1  g417(.A(new_n842), .B(KEYINPUT99), .ZN(new_n843));
  NAND2_X1  g418(.A1(new_n838), .A2(KEYINPUT100), .ZN(new_n844));
  OR2_X1    g419(.A1(new_n837), .A2(new_n844), .ZN(new_n845));
  AOI21_X1  g420(.A(new_n841), .B1(new_n837), .B2(new_n844), .ZN(new_n846));
  AOI21_X1  g421(.A(G37), .B1(new_n845), .B2(new_n846), .ZN(new_n847));
  NAND2_X1  g422(.A1(new_n843), .A2(new_n847), .ZN(new_n848));
  XNOR2_X1  g423(.A(new_n848), .B(KEYINPUT40), .ZN(G395));
  XNOR2_X1  g424(.A(G305), .B(G303), .ZN(new_n850));
  XNOR2_X1  g425(.A(G290), .B(G288), .ZN(new_n851));
  AOI21_X1  g426(.A(new_n850), .B1(new_n851), .B2(KEYINPUT103), .ZN(new_n852));
  NOR2_X1   g427(.A1(new_n851), .A2(KEYINPUT103), .ZN(new_n853));
  XNOR2_X1  g428(.A(new_n852), .B(new_n853), .ZN(new_n854));
  XOR2_X1   g429(.A(new_n854), .B(KEYINPUT42), .Z(new_n855));
  XOR2_X1   g430(.A(new_n592), .B(G299), .Z(new_n856));
  INV_X1    g431(.A(KEYINPUT41), .ZN(new_n857));
  XNOR2_X1  g432(.A(new_n856), .B(new_n857), .ZN(new_n858));
  NAND2_X1  g433(.A1(new_n856), .A2(new_n857), .ZN(new_n859));
  MUX2_X1   g434(.A(new_n858), .B(new_n859), .S(KEYINPUT102), .Z(new_n860));
  XOR2_X1   g435(.A(new_n814), .B(KEYINPUT101), .Z(new_n861));
  XNOR2_X1  g436(.A(new_n861), .B(new_n602), .ZN(new_n862));
  MUX2_X1   g437(.A(new_n860), .B(new_n856), .S(new_n862), .Z(new_n863));
  OAI21_X1  g438(.A(new_n855), .B1(new_n863), .B2(KEYINPUT104), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n863), .A2(KEYINPUT104), .ZN(new_n865));
  NAND2_X1  g440(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  NAND3_X1  g441(.A1(new_n863), .A2(new_n855), .A3(KEYINPUT104), .ZN(new_n867));
  AOI21_X1  g442(.A(new_n596), .B1(new_n866), .B2(new_n867), .ZN(new_n868));
  NOR2_X1   g443(.A1(new_n813), .A2(G868), .ZN(new_n869));
  OR3_X1    g444(.A1(new_n868), .A2(KEYINPUT105), .A3(new_n869), .ZN(new_n870));
  OAI21_X1  g445(.A(KEYINPUT105), .B1(new_n868), .B2(new_n869), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n870), .A2(new_n871), .ZN(G295));
  OR2_X1    g447(.A1(new_n868), .A2(new_n869), .ZN(G331));
  XNOR2_X1  g448(.A(G168), .B(G171), .ZN(new_n874));
  OR2_X1    g449(.A1(new_n874), .A2(new_n814), .ZN(new_n875));
  XOR2_X1   g450(.A(new_n875), .B(KEYINPUT106), .Z(new_n876));
  NAND2_X1  g451(.A1(new_n874), .A2(new_n814), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  AND2_X1   g453(.A1(new_n877), .A2(new_n856), .ZN(new_n879));
  AOI22_X1  g454(.A1(new_n878), .A2(new_n858), .B1(new_n875), .B2(new_n879), .ZN(new_n880));
  NOR2_X1   g455(.A1(new_n880), .A2(new_n854), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n875), .A2(new_n877), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n860), .A2(new_n882), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n876), .A2(new_n879), .ZN(new_n884));
  AND3_X1   g459(.A1(new_n883), .A2(new_n854), .A3(new_n884), .ZN(new_n885));
  NOR3_X1   g460(.A1(new_n881), .A2(G37), .A3(new_n885), .ZN(new_n886));
  AND2_X1   g461(.A1(new_n886), .A2(KEYINPUT43), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n883), .A2(new_n884), .ZN(new_n888));
  NOR2_X1   g463(.A1(new_n854), .A2(KEYINPUT107), .ZN(new_n889));
  OR2_X1    g464(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  AOI21_X1  g465(.A(G37), .B1(new_n888), .B2(new_n889), .ZN(new_n891));
  AOI21_X1  g466(.A(KEYINPUT43), .B1(new_n890), .B2(new_n891), .ZN(new_n892));
  OAI21_X1  g467(.A(KEYINPUT44), .B1(new_n887), .B2(new_n892), .ZN(new_n893));
  INV_X1    g468(.A(KEYINPUT43), .ZN(new_n894));
  AOI21_X1  g469(.A(new_n894), .B1(new_n890), .B2(new_n891), .ZN(new_n895));
  AOI21_X1  g470(.A(new_n895), .B1(new_n894), .B2(new_n886), .ZN(new_n896));
  OAI21_X1  g471(.A(new_n893), .B1(new_n896), .B2(KEYINPUT44), .ZN(G397));
  AOI21_X1  g472(.A(G1384), .B1(new_n499), .B2(new_n503), .ZN(new_n898));
  XNOR2_X1  g473(.A(KEYINPUT108), .B(KEYINPUT45), .ZN(new_n899));
  INV_X1    g474(.A(new_n899), .ZN(new_n900));
  NOR2_X1   g475(.A1(new_n898), .A2(new_n900), .ZN(new_n901));
  XOR2_X1   g476(.A(KEYINPUT109), .B(G40), .Z(new_n902));
  NOR3_X1   g477(.A1(new_n474), .A2(new_n481), .A3(new_n902), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n901), .A2(new_n903), .ZN(new_n904));
  XNOR2_X1  g479(.A(new_n757), .B(G2067), .ZN(new_n905));
  AND2_X1   g480(.A1(new_n719), .A2(G1996), .ZN(new_n906));
  INV_X1    g481(.A(G1996), .ZN(new_n907));
  AOI211_X1 g482(.A(new_n905), .B(new_n906), .C1(new_n720), .C2(new_n907), .ZN(new_n908));
  INV_X1    g483(.A(new_n705), .ZN(new_n909));
  NOR2_X1   g484(.A1(new_n703), .A2(new_n909), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n908), .A2(new_n910), .ZN(new_n911));
  INV_X1    g486(.A(G2067), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n758), .A2(new_n912), .ZN(new_n913));
  AOI21_X1  g488(.A(new_n904), .B1(new_n911), .B2(new_n913), .ZN(new_n914));
  XOR2_X1   g489(.A(new_n914), .B(KEYINPUT127), .Z(new_n915));
  INV_X1    g490(.A(new_n904), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n916), .A2(new_n907), .ZN(new_n917));
  XNOR2_X1  g492(.A(new_n917), .B(KEYINPUT46), .ZN(new_n918));
  OAI21_X1  g493(.A(new_n916), .B1(new_n719), .B2(new_n905), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  XNOR2_X1  g495(.A(new_n920), .B(KEYINPUT47), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n695), .A2(new_n697), .ZN(new_n922));
  XNOR2_X1  g497(.A(new_n922), .B(KEYINPUT110), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n923), .A2(new_n916), .ZN(new_n924));
  INV_X1    g499(.A(new_n924), .ZN(new_n925));
  XNOR2_X1  g500(.A(new_n703), .B(new_n705), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n908), .A2(new_n926), .ZN(new_n927));
  AOI22_X1  g502(.A1(KEYINPUT48), .A2(new_n925), .B1(new_n927), .B2(new_n916), .ZN(new_n928));
  OAI21_X1  g503(.A(new_n928), .B1(KEYINPUT48), .B2(new_n925), .ZN(new_n929));
  AND3_X1   g504(.A1(new_n915), .A2(new_n921), .A3(new_n929), .ZN(new_n930));
  INV_X1    g505(.A(new_n903), .ZN(new_n931));
  AOI21_X1  g506(.A(new_n931), .B1(KEYINPUT45), .B2(new_n898), .ZN(new_n932));
  INV_X1    g507(.A(KEYINPUT72), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n825), .A2(new_n933), .ZN(new_n934));
  NAND3_X1  g509(.A1(new_n499), .A2(KEYINPUT72), .A3(new_n503), .ZN(new_n935));
  AOI21_X1  g510(.A(G1384), .B1(new_n934), .B2(new_n935), .ZN(new_n936));
  OAI21_X1  g511(.A(new_n932), .B1(new_n936), .B2(new_n900), .ZN(new_n937));
  INV_X1    g512(.A(G1971), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  INV_X1    g514(.A(KEYINPUT50), .ZN(new_n940));
  AOI21_X1  g515(.A(new_n931), .B1(new_n940), .B2(new_n898), .ZN(new_n941));
  OAI21_X1  g516(.A(new_n941), .B1(new_n936), .B2(new_n940), .ZN(new_n942));
  OAI21_X1  g517(.A(new_n939), .B1(G2090), .B2(new_n942), .ZN(new_n943));
  NAND2_X1  g518(.A1(G303), .A2(G8), .ZN(new_n944));
  XOR2_X1   g519(.A(new_n944), .B(KEYINPUT55), .Z(new_n945));
  NAND3_X1  g520(.A1(new_n943), .A2(G8), .A3(new_n945), .ZN(new_n946));
  INV_X1    g521(.A(KEYINPUT52), .ZN(new_n947));
  INV_X1    g522(.A(G1384), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n825), .A2(new_n948), .ZN(new_n949));
  NOR2_X1   g524(.A1(new_n949), .A2(new_n931), .ZN(new_n950));
  XNOR2_X1  g525(.A(KEYINPUT111), .B(G8), .ZN(new_n951));
  NOR2_X1   g526(.A1(new_n950), .A2(new_n951), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n687), .A2(G1976), .ZN(new_n953));
  OR2_X1    g528(.A1(new_n687), .A2(G1976), .ZN(new_n954));
  AND4_X1   g529(.A1(new_n947), .A2(new_n952), .A3(new_n953), .A4(new_n954), .ZN(new_n955));
  NOR2_X1   g530(.A1(G305), .A2(G1981), .ZN(new_n956));
  INV_X1    g531(.A(KEYINPUT49), .ZN(new_n957));
  NOR2_X1   g532(.A1(new_n574), .A2(new_n683), .ZN(new_n958));
  OR3_X1    g533(.A1(new_n956), .A2(new_n957), .A3(new_n958), .ZN(new_n959));
  OAI21_X1  g534(.A(new_n957), .B1(new_n956), .B2(new_n958), .ZN(new_n960));
  AND3_X1   g535(.A1(new_n959), .A2(new_n952), .A3(new_n960), .ZN(new_n961));
  AOI21_X1  g536(.A(new_n947), .B1(new_n952), .B2(new_n953), .ZN(new_n962));
  NOR3_X1   g537(.A1(new_n955), .A2(new_n961), .A3(new_n962), .ZN(new_n963));
  AOI21_X1  g538(.A(new_n931), .B1(new_n949), .B2(KEYINPUT50), .ZN(new_n964));
  OAI21_X1  g539(.A(new_n948), .B1(new_n504), .B2(new_n505), .ZN(new_n965));
  OAI21_X1  g540(.A(new_n964), .B1(new_n965), .B2(KEYINPUT50), .ZN(new_n966));
  OR2_X1    g541(.A1(new_n966), .A2(G2090), .ZN(new_n967));
  AOI21_X1  g542(.A(new_n951), .B1(new_n967), .B2(new_n939), .ZN(new_n968));
  OAI211_X1 g543(.A(new_n946), .B(new_n963), .C1(new_n945), .C2(new_n968), .ZN(new_n969));
  INV_X1    g544(.A(KEYINPUT53), .ZN(new_n970));
  OAI21_X1  g545(.A(new_n970), .B1(new_n937), .B2(G2078), .ZN(new_n971));
  INV_X1    g546(.A(KEYINPUT118), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n942), .A2(new_n972), .ZN(new_n973));
  OAI211_X1 g548(.A(KEYINPUT118), .B(new_n941), .C1(new_n936), .C2(new_n940), .ZN(new_n974));
  NAND3_X1  g549(.A1(new_n973), .A2(new_n767), .A3(new_n974), .ZN(new_n975));
  OAI21_X1  g550(.A(new_n903), .B1(new_n898), .B2(KEYINPUT45), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n976), .A2(KEYINPUT112), .ZN(new_n977));
  INV_X1    g552(.A(KEYINPUT112), .ZN(new_n978));
  OAI211_X1 g553(.A(new_n978), .B(new_n903), .C1(new_n898), .C2(KEYINPUT45), .ZN(new_n979));
  OAI211_X1 g554(.A(new_n948), .B(new_n900), .C1(new_n504), .C2(new_n505), .ZN(new_n980));
  NAND3_X1  g555(.A1(new_n977), .A2(new_n979), .A3(new_n980), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n789), .A2(KEYINPUT53), .ZN(new_n982));
  OR2_X1    g557(.A1(new_n981), .A2(new_n982), .ZN(new_n983));
  AND3_X1   g558(.A1(new_n975), .A2(KEYINPUT125), .A3(new_n983), .ZN(new_n984));
  AOI21_X1  g559(.A(KEYINPUT125), .B1(new_n975), .B2(new_n983), .ZN(new_n985));
  OAI211_X1 g560(.A(G301), .B(new_n971), .C1(new_n984), .C2(new_n985), .ZN(new_n986));
  INV_X1    g561(.A(KEYINPUT54), .ZN(new_n987));
  AND2_X1   g562(.A1(new_n898), .A2(KEYINPUT45), .ZN(new_n988));
  NAND3_X1  g563(.A1(new_n789), .A2(KEYINPUT53), .A3(G40), .ZN(new_n989));
  OR4_X1    g564(.A1(new_n772), .A2(new_n988), .A3(new_n901), .A4(new_n989), .ZN(new_n990));
  NAND3_X1  g565(.A1(new_n975), .A2(new_n971), .A3(new_n990), .ZN(new_n991));
  AOI21_X1  g566(.A(new_n987), .B1(new_n991), .B2(G171), .ZN(new_n992));
  AOI21_X1  g567(.A(new_n969), .B1(new_n986), .B2(new_n992), .ZN(new_n993));
  INV_X1    g568(.A(new_n951), .ZN(new_n994));
  INV_X1    g569(.A(G1966), .ZN(new_n995));
  AND2_X1   g570(.A1(new_n981), .A2(new_n995), .ZN(new_n996));
  OAI211_X1 g571(.A(new_n774), .B(new_n941), .C1(new_n936), .C2(new_n940), .ZN(new_n997));
  INV_X1    g572(.A(new_n997), .ZN(new_n998));
  OAI21_X1  g573(.A(new_n994), .B1(new_n996), .B2(new_n998), .ZN(new_n999));
  NOR2_X1   g574(.A1(G168), .A2(new_n951), .ZN(new_n1000));
  NOR2_X1   g575(.A1(new_n1000), .A2(KEYINPUT51), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n999), .A2(new_n1001), .ZN(new_n1002));
  INV_X1    g577(.A(G8), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n981), .A2(new_n995), .ZN(new_n1004));
  AOI21_X1  g579(.A(new_n1003), .B1(new_n1004), .B2(new_n997), .ZN(new_n1005));
  OAI21_X1  g580(.A(KEYINPUT51), .B1(new_n1005), .B2(new_n1000), .ZN(new_n1006));
  OAI21_X1  g581(.A(new_n903), .B1(new_n949), .B2(KEYINPUT50), .ZN(new_n1007));
  AOI21_X1  g582(.A(new_n1007), .B1(KEYINPUT50), .B2(new_n965), .ZN(new_n1008));
  AOI22_X1  g583(.A1(new_n774), .A2(new_n1008), .B1(new_n981), .B2(new_n995), .ZN(new_n1009));
  NOR3_X1   g584(.A1(new_n1009), .A2(G168), .A3(new_n951), .ZN(new_n1010));
  OAI21_X1  g585(.A(new_n1002), .B1(new_n1006), .B2(new_n1010), .ZN(new_n1011));
  NOR2_X1   g586(.A1(new_n1011), .A2(KEYINPUT124), .ZN(new_n1012));
  INV_X1    g587(.A(KEYINPUT124), .ZN(new_n1013));
  OAI211_X1 g588(.A(G286), .B(new_n994), .C1(new_n996), .C2(new_n998), .ZN(new_n1014));
  OAI211_X1 g589(.A(new_n1014), .B(KEYINPUT51), .C1(new_n1000), .C2(new_n1005), .ZN(new_n1015));
  AOI21_X1  g590(.A(new_n1013), .B1(new_n1015), .B2(new_n1002), .ZN(new_n1016));
  OAI21_X1  g591(.A(new_n993), .B1(new_n1012), .B2(new_n1016), .ZN(new_n1017));
  INV_X1    g592(.A(new_n1017), .ZN(new_n1018));
  AOI21_X1  g593(.A(new_n553), .B1(new_n516), .B2(G53), .ZN(new_n1019));
  NOR2_X1   g594(.A1(new_n557), .A2(KEYINPUT9), .ZN(new_n1020));
  OAI21_X1  g595(.A(KEYINPUT114), .B1(new_n1019), .B2(new_n1020), .ZN(new_n1021));
  INV_X1    g596(.A(KEYINPUT114), .ZN(new_n1022));
  NAND3_X1  g597(.A1(new_n554), .A2(new_n558), .A3(new_n1022), .ZN(new_n1023));
  NAND4_X1  g598(.A1(new_n552), .A2(new_n1021), .A3(new_n561), .A4(new_n1023), .ZN(new_n1024));
  INV_X1    g599(.A(KEYINPUT57), .ZN(new_n1025));
  NAND3_X1  g600(.A1(new_n1024), .A2(KEYINPUT115), .A3(new_n1025), .ZN(new_n1026));
  NAND4_X1  g601(.A1(new_n552), .A2(KEYINPUT57), .A3(new_n559), .A4(new_n561), .ZN(new_n1027));
  NAND2_X1  g602(.A1(new_n1026), .A2(new_n1027), .ZN(new_n1028));
  AOI21_X1  g603(.A(KEYINPUT115), .B1(new_n1024), .B2(new_n1025), .ZN(new_n1029));
  OAI21_X1  g604(.A(KEYINPUT116), .B1(new_n1028), .B2(new_n1029), .ZN(new_n1030));
  NAND2_X1  g605(.A1(new_n1024), .A2(new_n1025), .ZN(new_n1031));
  INV_X1    g606(.A(KEYINPUT115), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n1031), .A2(new_n1032), .ZN(new_n1033));
  INV_X1    g608(.A(KEYINPUT116), .ZN(new_n1034));
  NAND4_X1  g609(.A1(new_n1033), .A2(new_n1034), .A3(new_n1027), .A4(new_n1026), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n1030), .A2(new_n1035), .ZN(new_n1036));
  INV_X1    g611(.A(G1956), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n966), .A2(new_n1037), .ZN(new_n1038));
  XNOR2_X1  g613(.A(KEYINPUT56), .B(G2072), .ZN(new_n1039));
  OAI211_X1 g614(.A(new_n932), .B(new_n1039), .C1(new_n936), .C2(new_n900), .ZN(new_n1040));
  NAND3_X1  g615(.A1(new_n1036), .A2(new_n1038), .A3(new_n1040), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n1041), .A2(KEYINPUT117), .ZN(new_n1042));
  INV_X1    g617(.A(KEYINPUT117), .ZN(new_n1043));
  NAND4_X1  g618(.A1(new_n1036), .A2(new_n1038), .A3(new_n1043), .A4(new_n1040), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n1042), .A2(new_n1044), .ZN(new_n1045));
  NAND2_X1  g620(.A1(new_n1038), .A2(new_n1040), .ZN(new_n1046));
  INV_X1    g621(.A(KEYINPUT119), .ZN(new_n1047));
  AOI21_X1  g622(.A(new_n1036), .B1(new_n1046), .B2(new_n1047), .ZN(new_n1048));
  NAND3_X1  g623(.A1(new_n1038), .A2(KEYINPUT119), .A3(new_n1040), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n1048), .A2(new_n1049), .ZN(new_n1050));
  INV_X1    g625(.A(new_n1050), .ZN(new_n1051));
  NAND3_X1  g626(.A1(new_n973), .A2(new_n779), .A3(new_n974), .ZN(new_n1052));
  NAND2_X1  g627(.A1(new_n950), .A2(new_n912), .ZN(new_n1053));
  AOI21_X1  g628(.A(new_n592), .B1(new_n1052), .B2(new_n1053), .ZN(new_n1054));
  OAI21_X1  g629(.A(new_n1045), .B1(new_n1051), .B2(new_n1054), .ZN(new_n1055));
  OR2_X1    g630(.A1(new_n1041), .A2(KEYINPUT122), .ZN(new_n1056));
  INV_X1    g631(.A(KEYINPUT61), .ZN(new_n1057));
  AOI21_X1  g632(.A(new_n1057), .B1(new_n1041), .B2(KEYINPUT122), .ZN(new_n1058));
  NAND3_X1  g633(.A1(new_n1050), .A2(new_n1056), .A3(new_n1058), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n1052), .A2(new_n1053), .ZN(new_n1060));
  INV_X1    g635(.A(KEYINPUT60), .ZN(new_n1061));
  NAND2_X1  g636(.A1(new_n1060), .A2(new_n1061), .ZN(new_n1062));
  NAND3_X1  g637(.A1(new_n1052), .A2(KEYINPUT60), .A3(new_n1053), .ZN(new_n1063));
  NAND3_X1  g638(.A1(new_n1062), .A2(new_n593), .A3(new_n1063), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n1059), .A2(new_n1064), .ZN(new_n1065));
  NAND4_X1  g640(.A1(new_n1052), .A2(KEYINPUT60), .A3(new_n592), .A4(new_n1053), .ZN(new_n1066));
  OR2_X1    g641(.A1(KEYINPUT121), .A2(KEYINPUT59), .ZN(new_n1067));
  XNOR2_X1  g642(.A(KEYINPUT120), .B(KEYINPUT58), .ZN(new_n1068));
  XNOR2_X1  g643(.A(new_n1068), .B(new_n736), .ZN(new_n1069));
  OAI21_X1  g644(.A(new_n1069), .B1(new_n949), .B2(new_n931), .ZN(new_n1070));
  OAI21_X1  g645(.A(new_n1070), .B1(new_n937), .B2(G1996), .ZN(new_n1071));
  AOI21_X1  g646(.A(new_n1067), .B1(new_n1071), .B2(new_n542), .ZN(new_n1072));
  AND2_X1   g647(.A1(new_n1071), .A2(new_n542), .ZN(new_n1073));
  XOR2_X1   g648(.A(KEYINPUT121), .B(KEYINPUT59), .Z(new_n1074));
  AOI21_X1  g649(.A(new_n1072), .B1(new_n1073), .B2(new_n1074), .ZN(new_n1075));
  AOI21_X1  g650(.A(new_n1036), .B1(new_n1038), .B2(new_n1040), .ZN(new_n1076));
  AOI21_X1  g651(.A(new_n1076), .B1(new_n1042), .B2(new_n1044), .ZN(new_n1077));
  OAI211_X1 g652(.A(new_n1066), .B(new_n1075), .C1(new_n1077), .C2(KEYINPUT61), .ZN(new_n1078));
  OAI21_X1  g653(.A(new_n1055), .B1(new_n1065), .B2(new_n1078), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n1079), .A2(KEYINPUT123), .ZN(new_n1080));
  OAI21_X1  g655(.A(new_n971), .B1(new_n984), .B2(new_n985), .ZN(new_n1081));
  AND2_X1   g656(.A1(new_n1081), .A2(G171), .ZN(new_n1082));
  NOR2_X1   g657(.A1(new_n991), .A2(G171), .ZN(new_n1083));
  OAI21_X1  g658(.A(new_n987), .B1(new_n1082), .B2(new_n1083), .ZN(new_n1084));
  INV_X1    g659(.A(KEYINPUT123), .ZN(new_n1085));
  OAI211_X1 g660(.A(new_n1085), .B(new_n1055), .C1(new_n1065), .C2(new_n1078), .ZN(new_n1086));
  NAND4_X1  g661(.A1(new_n1018), .A2(new_n1080), .A3(new_n1084), .A4(new_n1086), .ZN(new_n1087));
  NAND2_X1  g662(.A1(new_n943), .A2(G8), .ZN(new_n1088));
  INV_X1    g663(.A(KEYINPUT113), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n1088), .A2(new_n1089), .ZN(new_n1090));
  INV_X1    g665(.A(new_n945), .ZN(new_n1091));
  NAND3_X1  g666(.A1(new_n943), .A2(KEYINPUT113), .A3(G8), .ZN(new_n1092));
  NAND3_X1  g667(.A1(new_n1090), .A2(new_n1091), .A3(new_n1092), .ZN(new_n1093));
  AND3_X1   g668(.A1(new_n946), .A2(new_n963), .A3(KEYINPUT63), .ZN(new_n1094));
  NOR2_X1   g669(.A1(new_n999), .A2(G286), .ZN(new_n1095));
  NAND3_X1  g670(.A1(new_n1093), .A2(new_n1094), .A3(new_n1095), .ZN(new_n1096));
  INV_X1    g671(.A(KEYINPUT63), .ZN(new_n1097));
  OR2_X1    g672(.A1(new_n999), .A2(G286), .ZN(new_n1098));
  OAI21_X1  g673(.A(new_n1097), .B1(new_n969), .B2(new_n1098), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n1096), .A2(new_n1099), .ZN(new_n1100));
  NOR3_X1   g675(.A1(new_n961), .A2(G1976), .A3(G288), .ZN(new_n1101));
  OR2_X1    g676(.A1(new_n1101), .A2(new_n956), .ZN(new_n1102));
  NOR2_X1   g677(.A1(new_n1088), .A2(new_n1091), .ZN(new_n1103));
  AOI22_X1  g678(.A1(new_n952), .A2(new_n1102), .B1(new_n1103), .B2(new_n963), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n1100), .A2(new_n1104), .ZN(new_n1105));
  INV_X1    g680(.A(new_n969), .ZN(new_n1106));
  NAND3_X1  g681(.A1(new_n1106), .A2(G171), .A3(new_n1081), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n1011), .A2(KEYINPUT124), .ZN(new_n1108));
  NAND3_X1  g683(.A1(new_n1015), .A2(new_n1013), .A3(new_n1002), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n1108), .A2(new_n1109), .ZN(new_n1110));
  AOI21_X1  g685(.A(new_n1107), .B1(new_n1110), .B2(KEYINPUT62), .ZN(new_n1111));
  INV_X1    g686(.A(KEYINPUT62), .ZN(new_n1112));
  NAND3_X1  g687(.A1(new_n1108), .A2(new_n1112), .A3(new_n1109), .ZN(new_n1113));
  AOI21_X1  g688(.A(new_n1105), .B1(new_n1111), .B2(new_n1113), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n1087), .A2(new_n1114), .ZN(new_n1115));
  INV_X1    g690(.A(new_n927), .ZN(new_n1116));
  AOI21_X1  g691(.A(new_n923), .B1(G1986), .B2(G290), .ZN(new_n1117));
  AOI21_X1  g692(.A(new_n904), .B1(new_n1116), .B2(new_n1117), .ZN(new_n1118));
  INV_X1    g693(.A(new_n1118), .ZN(new_n1119));
  AOI21_X1  g694(.A(KEYINPUT126), .B1(new_n1115), .B2(new_n1119), .ZN(new_n1120));
  INV_X1    g695(.A(KEYINPUT126), .ZN(new_n1121));
  AOI211_X1 g696(.A(new_n1121), .B(new_n1118), .C1(new_n1087), .C2(new_n1114), .ZN(new_n1122));
  OAI21_X1  g697(.A(new_n930), .B1(new_n1120), .B2(new_n1122), .ZN(G329));
  assign    G231 = 1'b0;
  NOR4_X1   g698(.A1(G401), .A2(G229), .A3(new_n460), .A4(G227), .ZN(new_n1125));
  NAND2_X1  g699(.A1(new_n848), .A2(new_n1125), .ZN(new_n1126));
  NOR2_X1   g700(.A1(new_n1126), .A2(new_n896), .ZN(G308));
  OR2_X1    g701(.A1(new_n1126), .A2(new_n896), .ZN(G225));
endmodule


