//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 0 1 0 1 1 1 1 0 1 0 1 1 0 1 1 0 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 0 0 0 0 0 0 1 1 1 1 1 1 0 0 1 0 1 1 0 0 1 1 0 1 0 1 1 0 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:30:01 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n443, new_n444, new_n446, new_n450, new_n451, new_n455,
    new_n456, new_n457, new_n458, new_n461, new_n462, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n530, new_n531, new_n532,
    new_n533, new_n534, new_n535, new_n536, new_n537, new_n538, new_n539,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n548, new_n549,
    new_n550, new_n551, new_n552, new_n553, new_n556, new_n557, new_n559,
    new_n560, new_n561, new_n562, new_n564, new_n566, new_n567, new_n568,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n576, new_n577,
    new_n578, new_n579, new_n580, new_n581, new_n582, new_n584, new_n585,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n599, new_n602, new_n604, new_n605,
    new_n607, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n652,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1125, new_n1126, new_n1127, new_n1128;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  XOR2_X1   g003(.A(KEYINPUT64), .B(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  XNOR2_X1  g011(.A(KEYINPUT65), .B(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  XNOR2_X1  g013(.A(KEYINPUT66), .B(G120), .ZN(G236));
  XOR2_X1   g014(.A(KEYINPUT67), .B(G57), .Z(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  INV_X1    g016(.A(G2072), .ZN(new_n442));
  INV_X1    g017(.A(G2078), .ZN(new_n443));
  NOR2_X1   g018(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  NAND3_X1  g019(.A1(new_n444), .A2(G2084), .A3(G2090), .ZN(G158));
  NAND3_X1  g020(.A1(G2), .A2(G15), .A3(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT68), .Z(G259));
  BUF_X1    g022(.A(G452), .Z(G391));
  AND2_X1   g023(.A1(G94), .A2(G452), .ZN(G173));
  XNOR2_X1  g024(.A(KEYINPUT69), .B(KEYINPUT1), .ZN(new_n450));
  AND2_X1   g025(.A1(G7), .A2(G661), .ZN(new_n451));
  XNOR2_X1  g026(.A(new_n450), .B(new_n451), .ZN(G223));
  NAND2_X1  g027(.A1(new_n451), .A2(G567), .ZN(G234));
  NAND2_X1  g028(.A1(new_n451), .A2(G2106), .ZN(G217));
  OR4_X1    g029(.A1(G218), .A2(G220), .A3(G221), .A4(G219), .ZN(new_n455));
  XOR2_X1   g030(.A(new_n455), .B(KEYINPUT2), .Z(new_n456));
  NOR4_X1   g031(.A1(G237), .A2(G236), .A3(G235), .A4(G238), .ZN(new_n457));
  NAND2_X1  g032(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  XNOR2_X1  g033(.A(new_n458), .B(KEYINPUT70), .ZN(G261));
  INV_X1    g034(.A(G261), .ZN(G325));
  INV_X1    g035(.A(new_n456), .ZN(new_n461));
  INV_X1    g036(.A(new_n457), .ZN(new_n462));
  AOI22_X1  g037(.A1(new_n461), .A2(G2106), .B1(G567), .B2(new_n462), .ZN(G319));
  INV_X1    g038(.A(G2105), .ZN(new_n464));
  AND2_X1   g039(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n465));
  NOR2_X1   g040(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n466));
  OAI211_X1 g041(.A(G137), .B(new_n464), .C1(new_n465), .C2(new_n466), .ZN(new_n467));
  INV_X1    g042(.A(G101), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n464), .A2(G2104), .ZN(new_n469));
  OAI21_X1  g044(.A(new_n467), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  OAI21_X1  g045(.A(G125), .B1(new_n465), .B2(new_n466), .ZN(new_n471));
  INV_X1    g046(.A(KEYINPUT71), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  OAI211_X1 g048(.A(KEYINPUT71), .B(G125), .C1(new_n465), .C2(new_n466), .ZN(new_n474));
  NAND2_X1  g049(.A1(G113), .A2(G2104), .ZN(new_n475));
  NAND3_X1  g050(.A1(new_n473), .A2(new_n474), .A3(new_n475), .ZN(new_n476));
  AOI21_X1  g051(.A(new_n470), .B1(new_n476), .B2(G2105), .ZN(G160));
  OR2_X1    g052(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n478));
  NAND2_X1  g053(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n480), .A2(G2105), .ZN(new_n481));
  XNOR2_X1  g056(.A(new_n481), .B(KEYINPUT73), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n482), .A2(G124), .ZN(new_n483));
  OAI21_X1  g058(.A(KEYINPUT74), .B1(G100), .B2(G2105), .ZN(new_n484));
  INV_X1    g059(.A(new_n484), .ZN(new_n485));
  NOR3_X1   g060(.A1(KEYINPUT74), .A2(G100), .A3(G2105), .ZN(new_n486));
  OAI221_X1 g061(.A(G2104), .B1(G112), .B2(new_n464), .C1(new_n485), .C2(new_n486), .ZN(new_n487));
  INV_X1    g062(.A(G136), .ZN(new_n488));
  AOI21_X1  g063(.A(G2105), .B1(new_n478), .B2(new_n479), .ZN(new_n489));
  INV_X1    g064(.A(KEYINPUT72), .ZN(new_n490));
  OR2_X1    g065(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  NAND2_X1  g066(.A1(new_n489), .A2(new_n490), .ZN(new_n492));
  NAND2_X1  g067(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  OAI211_X1 g068(.A(new_n483), .B(new_n487), .C1(new_n488), .C2(new_n493), .ZN(new_n494));
  XNOR2_X1  g069(.A(new_n494), .B(KEYINPUT75), .ZN(G162));
  NAND2_X1  g070(.A1(G126), .A2(G2105), .ZN(new_n496));
  INV_X1    g071(.A(new_n496), .ZN(new_n497));
  OAI21_X1  g072(.A(new_n497), .B1(new_n465), .B2(new_n466), .ZN(new_n498));
  INV_X1    g073(.A(G102), .ZN(new_n499));
  NAND2_X1  g074(.A1(new_n499), .A2(new_n464), .ZN(new_n500));
  INV_X1    g075(.A(G114), .ZN(new_n501));
  NAND2_X1  g076(.A1(new_n501), .A2(G2105), .ZN(new_n502));
  NAND3_X1  g077(.A1(new_n500), .A2(new_n502), .A3(G2104), .ZN(new_n503));
  NAND2_X1  g078(.A1(new_n498), .A2(new_n503), .ZN(new_n504));
  OAI211_X1 g079(.A(G138), .B(new_n464), .C1(new_n465), .C2(new_n466), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n505), .A2(KEYINPUT4), .ZN(new_n506));
  INV_X1    g081(.A(KEYINPUT4), .ZN(new_n507));
  NAND4_X1  g082(.A1(new_n480), .A2(new_n507), .A3(G138), .A4(new_n464), .ZN(new_n508));
  AOI21_X1  g083(.A(new_n504), .B1(new_n506), .B2(new_n508), .ZN(G164));
  INV_X1    g084(.A(KEYINPUT5), .ZN(new_n510));
  OAI21_X1  g085(.A(KEYINPUT77), .B1(new_n510), .B2(G543), .ZN(new_n511));
  INV_X1    g086(.A(KEYINPUT77), .ZN(new_n512));
  INV_X1    g087(.A(G543), .ZN(new_n513));
  NAND3_X1  g088(.A1(new_n512), .A2(new_n513), .A3(KEYINPUT5), .ZN(new_n514));
  AOI22_X1  g089(.A1(new_n511), .A2(new_n514), .B1(new_n510), .B2(G543), .ZN(new_n515));
  INV_X1    g090(.A(G651), .ZN(new_n516));
  OAI21_X1  g091(.A(KEYINPUT76), .B1(new_n516), .B2(KEYINPUT6), .ZN(new_n517));
  INV_X1    g092(.A(KEYINPUT76), .ZN(new_n518));
  INV_X1    g093(.A(KEYINPUT6), .ZN(new_n519));
  NAND3_X1  g094(.A1(new_n518), .A2(new_n519), .A3(G651), .ZN(new_n520));
  AOI22_X1  g095(.A1(new_n517), .A2(new_n520), .B1(KEYINPUT6), .B2(new_n516), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n515), .A2(new_n521), .ZN(new_n522));
  INV_X1    g097(.A(G88), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n521), .A2(G543), .ZN(new_n524));
  INV_X1    g099(.A(G50), .ZN(new_n525));
  OAI22_X1  g100(.A1(new_n522), .A2(new_n523), .B1(new_n524), .B2(new_n525), .ZN(new_n526));
  AOI22_X1  g101(.A1(new_n515), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n527));
  NOR2_X1   g102(.A1(new_n527), .A2(new_n516), .ZN(new_n528));
  NOR2_X1   g103(.A1(new_n526), .A2(new_n528), .ZN(G166));
  AND2_X1   g104(.A1(new_n515), .A2(new_n521), .ZN(new_n530));
  NAND2_X1  g105(.A1(new_n530), .A2(G89), .ZN(new_n531));
  AND2_X1   g106(.A1(new_n521), .A2(G543), .ZN(new_n532));
  XOR2_X1   g107(.A(KEYINPUT78), .B(G51), .Z(new_n533));
  NAND2_X1  g108(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  AND2_X1   g109(.A1(G63), .A2(G651), .ZN(new_n535));
  NAND3_X1  g110(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n536));
  NAND2_X1  g111(.A1(new_n536), .A2(KEYINPUT7), .ZN(new_n537));
  OR2_X1    g112(.A1(new_n536), .A2(KEYINPUT7), .ZN(new_n538));
  AOI22_X1  g113(.A1(new_n515), .A2(new_n535), .B1(new_n537), .B2(new_n538), .ZN(new_n539));
  NAND3_X1  g114(.A1(new_n531), .A2(new_n534), .A3(new_n539), .ZN(G286));
  INV_X1    g115(.A(G286), .ZN(G168));
  INV_X1    g116(.A(G90), .ZN(new_n542));
  INV_X1    g117(.A(G52), .ZN(new_n543));
  OAI22_X1  g118(.A1(new_n522), .A2(new_n542), .B1(new_n524), .B2(new_n543), .ZN(new_n544));
  AOI22_X1  g119(.A1(new_n515), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n545));
  NOR2_X1   g120(.A1(new_n545), .A2(new_n516), .ZN(new_n546));
  NOR2_X1   g121(.A1(new_n544), .A2(new_n546), .ZN(G171));
  INV_X1    g122(.A(G81), .ZN(new_n548));
  INV_X1    g123(.A(G43), .ZN(new_n549));
  OAI22_X1  g124(.A1(new_n522), .A2(new_n548), .B1(new_n524), .B2(new_n549), .ZN(new_n550));
  AOI22_X1  g125(.A1(new_n515), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n551));
  NOR2_X1   g126(.A1(new_n551), .A2(new_n516), .ZN(new_n552));
  NOR2_X1   g127(.A1(new_n550), .A2(new_n552), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n553), .A2(G860), .ZN(G153));
  NAND4_X1  g129(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g130(.A1(G1), .A2(G3), .ZN(new_n556));
  XNOR2_X1  g131(.A(new_n556), .B(KEYINPUT8), .ZN(new_n557));
  NAND4_X1  g132(.A1(G319), .A2(G483), .A3(G661), .A4(new_n557), .ZN(G188));
  NAND4_X1  g133(.A1(new_n521), .A2(KEYINPUT79), .A3(G53), .A4(G543), .ZN(new_n559));
  XNOR2_X1  g134(.A(new_n559), .B(KEYINPUT9), .ZN(new_n560));
  NAND2_X1  g135(.A1(new_n530), .A2(G91), .ZN(new_n561));
  AOI22_X1  g136(.A1(new_n515), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n562));
  OAI211_X1 g137(.A(new_n560), .B(new_n561), .C1(new_n516), .C2(new_n562), .ZN(G299));
  XNOR2_X1  g138(.A(G171), .B(KEYINPUT80), .ZN(new_n564));
  INV_X1    g139(.A(new_n564), .ZN(G301));
  INV_X1    g140(.A(KEYINPUT81), .ZN(new_n566));
  NAND2_X1  g141(.A1(G166), .A2(new_n566), .ZN(new_n567));
  OAI21_X1  g142(.A(KEYINPUT81), .B1(new_n526), .B2(new_n528), .ZN(new_n568));
  AND2_X1   g143(.A1(new_n567), .A2(new_n568), .ZN(G303));
  NAND2_X1  g144(.A1(new_n530), .A2(G87), .ZN(new_n570));
  NAND2_X1  g145(.A1(new_n532), .A2(G49), .ZN(new_n571));
  OAI21_X1  g146(.A(G651), .B1(new_n515), .B2(G74), .ZN(new_n572));
  NAND3_X1  g147(.A1(new_n570), .A2(new_n571), .A3(new_n572), .ZN(new_n573));
  XNOR2_X1  g148(.A(new_n573), .B(KEYINPUT82), .ZN(new_n574));
  INV_X1    g149(.A(new_n574), .ZN(G288));
  INV_X1    g150(.A(G86), .ZN(new_n576));
  INV_X1    g151(.A(G48), .ZN(new_n577));
  OAI22_X1  g152(.A1(new_n522), .A2(new_n576), .B1(new_n524), .B2(new_n577), .ZN(new_n578));
  NAND2_X1  g153(.A1(new_n515), .A2(G61), .ZN(new_n579));
  NAND2_X1  g154(.A1(G73), .A2(G543), .ZN(new_n580));
  XNOR2_X1  g155(.A(new_n580), .B(KEYINPUT83), .ZN(new_n581));
  AOI21_X1  g156(.A(new_n516), .B1(new_n579), .B2(new_n581), .ZN(new_n582));
  OR2_X1    g157(.A1(new_n578), .A2(new_n582), .ZN(G305));
  AOI22_X1  g158(.A1(G85), .A2(new_n530), .B1(new_n532), .B2(G47), .ZN(new_n584));
  AOI22_X1  g159(.A1(new_n515), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n585));
  OAI21_X1  g160(.A(new_n584), .B1(new_n516), .B2(new_n585), .ZN(G290));
  INV_X1    g161(.A(G868), .ZN(new_n587));
  NOR2_X1   g162(.A1(G301), .A2(new_n587), .ZN(new_n588));
  NAND2_X1  g163(.A1(new_n532), .A2(G54), .ZN(new_n589));
  AOI22_X1  g164(.A1(new_n515), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n590));
  NAND2_X1  g165(.A1(new_n530), .A2(G92), .ZN(new_n591));
  INV_X1    g166(.A(KEYINPUT10), .ZN(new_n592));
  NOR2_X1   g167(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  AOI21_X1  g168(.A(KEYINPUT10), .B1(new_n530), .B2(G92), .ZN(new_n594));
  OAI221_X1 g169(.A(new_n589), .B1(new_n516), .B2(new_n590), .C1(new_n593), .C2(new_n594), .ZN(new_n595));
  XOR2_X1   g170(.A(new_n595), .B(KEYINPUT84), .Z(new_n596));
  AOI21_X1  g171(.A(new_n588), .B1(new_n596), .B2(new_n587), .ZN(G284));
  AOI21_X1  g172(.A(new_n588), .B1(new_n596), .B2(new_n587), .ZN(G321));
  NAND2_X1  g173(.A1(G299), .A2(new_n587), .ZN(new_n599));
  OAI21_X1  g174(.A(new_n599), .B1(new_n587), .B2(G168), .ZN(G297));
  OAI21_X1  g175(.A(new_n599), .B1(new_n587), .B2(G168), .ZN(G280));
  INV_X1    g176(.A(G559), .ZN(new_n602));
  OAI21_X1  g177(.A(new_n596), .B1(new_n602), .B2(G860), .ZN(G148));
  NAND2_X1  g178(.A1(new_n596), .A2(new_n602), .ZN(new_n604));
  NAND2_X1  g179(.A1(new_n604), .A2(G868), .ZN(new_n605));
  OAI21_X1  g180(.A(new_n605), .B1(G868), .B2(new_n553), .ZN(G323));
  XNOR2_X1  g181(.A(KEYINPUT85), .B(KEYINPUT11), .ZN(new_n607));
  XNOR2_X1  g182(.A(G323), .B(new_n607), .ZN(G282));
  AND2_X1   g183(.A1(new_n482), .A2(G123), .ZN(new_n609));
  OR2_X1    g184(.A1(G99), .A2(G2105), .ZN(new_n610));
  OAI211_X1 g185(.A(new_n610), .B(G2104), .C1(G111), .C2(new_n464), .ZN(new_n611));
  INV_X1    g186(.A(G135), .ZN(new_n612));
  OAI21_X1  g187(.A(new_n611), .B1(new_n493), .B2(new_n612), .ZN(new_n613));
  NOR2_X1   g188(.A1(new_n609), .A2(new_n613), .ZN(new_n614));
  XNOR2_X1  g189(.A(KEYINPUT86), .B(G2096), .ZN(new_n615));
  OR2_X1    g190(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  NAND2_X1  g191(.A1(new_n614), .A2(new_n615), .ZN(new_n617));
  NAND3_X1  g192(.A1(new_n464), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n618));
  XNOR2_X1  g193(.A(new_n618), .B(KEYINPUT12), .ZN(new_n619));
  XNOR2_X1  g194(.A(new_n619), .B(KEYINPUT13), .ZN(new_n620));
  XNOR2_X1  g195(.A(new_n620), .B(G2100), .ZN(new_n621));
  NAND3_X1  g196(.A1(new_n616), .A2(new_n617), .A3(new_n621), .ZN(G156));
  XOR2_X1   g197(.A(G2451), .B(G2454), .Z(new_n623));
  XNOR2_X1  g198(.A(new_n623), .B(KEYINPUT16), .ZN(new_n624));
  XNOR2_X1  g199(.A(G1341), .B(G1348), .ZN(new_n625));
  XNOR2_X1  g200(.A(new_n624), .B(new_n625), .ZN(new_n626));
  INV_X1    g201(.A(KEYINPUT14), .ZN(new_n627));
  XNOR2_X1  g202(.A(G2427), .B(G2438), .ZN(new_n628));
  XNOR2_X1  g203(.A(new_n628), .B(G2430), .ZN(new_n629));
  XNOR2_X1  g204(.A(KEYINPUT15), .B(G2435), .ZN(new_n630));
  AOI21_X1  g205(.A(new_n627), .B1(new_n629), .B2(new_n630), .ZN(new_n631));
  OAI21_X1  g206(.A(new_n631), .B1(new_n630), .B2(new_n629), .ZN(new_n632));
  XOR2_X1   g207(.A(new_n626), .B(new_n632), .Z(new_n633));
  XNOR2_X1  g208(.A(G2443), .B(G2446), .ZN(new_n634));
  OR2_X1    g209(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  NAND2_X1  g210(.A1(new_n633), .A2(new_n634), .ZN(new_n636));
  NAND3_X1  g211(.A1(new_n635), .A2(new_n636), .A3(G14), .ZN(new_n637));
  XNOR2_X1  g212(.A(new_n637), .B(KEYINPUT87), .ZN(G401));
  XOR2_X1   g213(.A(G2084), .B(G2090), .Z(new_n639));
  XNOR2_X1  g214(.A(new_n639), .B(KEYINPUT88), .ZN(new_n640));
  XNOR2_X1  g215(.A(G2067), .B(G2678), .ZN(new_n641));
  NAND2_X1  g216(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  AND2_X1   g217(.A1(new_n642), .A2(KEYINPUT17), .ZN(new_n643));
  OR2_X1    g218(.A1(new_n640), .A2(new_n641), .ZN(new_n644));
  AOI21_X1  g219(.A(KEYINPUT18), .B1(new_n643), .B2(new_n644), .ZN(new_n645));
  XNOR2_X1  g220(.A(G2096), .B(G2100), .ZN(new_n646));
  XNOR2_X1  g221(.A(new_n645), .B(new_n646), .ZN(new_n647));
  XOR2_X1   g222(.A(G2072), .B(G2078), .Z(new_n648));
  AOI21_X1  g223(.A(new_n648), .B1(new_n642), .B2(KEYINPUT18), .ZN(new_n649));
  XOR2_X1   g224(.A(new_n649), .B(KEYINPUT89), .Z(new_n650));
  XNOR2_X1  g225(.A(new_n647), .B(new_n650), .ZN(G227));
  XOR2_X1   g226(.A(G1971), .B(G1976), .Z(new_n652));
  XNOR2_X1  g227(.A(new_n652), .B(KEYINPUT19), .ZN(new_n653));
  XNOR2_X1  g228(.A(G1956), .B(G2474), .ZN(new_n654));
  XNOR2_X1  g229(.A(G1961), .B(G1966), .ZN(new_n655));
  NOR2_X1   g230(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  AND2_X1   g231(.A1(new_n654), .A2(new_n655), .ZN(new_n657));
  NOR3_X1   g232(.A1(new_n653), .A2(new_n656), .A3(new_n657), .ZN(new_n658));
  NAND2_X1  g233(.A1(new_n653), .A2(new_n656), .ZN(new_n659));
  XOR2_X1   g234(.A(new_n659), .B(KEYINPUT20), .Z(new_n660));
  AOI211_X1 g235(.A(new_n658), .B(new_n660), .C1(new_n653), .C2(new_n657), .ZN(new_n661));
  XNOR2_X1  g236(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n662));
  XNOR2_X1  g237(.A(new_n661), .B(new_n662), .ZN(new_n663));
  XNOR2_X1  g238(.A(G1991), .B(G1996), .ZN(new_n664));
  XNOR2_X1  g239(.A(new_n663), .B(new_n664), .ZN(new_n665));
  XNOR2_X1  g240(.A(G1981), .B(G1986), .ZN(new_n666));
  XNOR2_X1  g241(.A(new_n665), .B(new_n666), .ZN(new_n667));
  INV_X1    g242(.A(new_n667), .ZN(G229));
  NAND3_X1  g243(.A1(new_n464), .A2(G103), .A3(G2104), .ZN(new_n669));
  XOR2_X1   g244(.A(new_n669), .B(KEYINPUT25), .Z(new_n670));
  AOI22_X1  g245(.A1(new_n480), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n671));
  OAI21_X1  g246(.A(new_n670), .B1(new_n671), .B2(new_n464), .ZN(new_n672));
  INV_X1    g247(.A(new_n493), .ZN(new_n673));
  AOI21_X1  g248(.A(new_n672), .B1(new_n673), .B2(G139), .ZN(new_n674));
  XNOR2_X1  g249(.A(new_n674), .B(KEYINPUT99), .ZN(new_n675));
  MUX2_X1   g250(.A(G33), .B(new_n675), .S(G29), .Z(new_n676));
  XNOR2_X1  g251(.A(new_n676), .B(KEYINPUT100), .ZN(new_n677));
  OR2_X1    g252(.A1(new_n677), .A2(new_n442), .ZN(new_n678));
  NAND2_X1  g253(.A1(new_n677), .A2(new_n442), .ZN(new_n679));
  NAND3_X1  g254(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n680));
  XOR2_X1   g255(.A(new_n680), .B(KEYINPUT26), .Z(new_n681));
  INV_X1    g256(.A(G105), .ZN(new_n682));
  OAI21_X1  g257(.A(new_n681), .B1(new_n682), .B2(new_n469), .ZN(new_n683));
  AOI21_X1  g258(.A(new_n683), .B1(new_n482), .B2(G129), .ZN(new_n684));
  NAND2_X1  g259(.A1(new_n673), .A2(G141), .ZN(new_n685));
  NAND2_X1  g260(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  INV_X1    g261(.A(new_n686), .ZN(new_n687));
  INV_X1    g262(.A(G29), .ZN(new_n688));
  NOR2_X1   g263(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  AOI21_X1  g264(.A(new_n689), .B1(new_n688), .B2(G32), .ZN(new_n690));
  XNOR2_X1  g265(.A(KEYINPUT27), .B(G1996), .ZN(new_n691));
  INV_X1    g266(.A(KEYINPUT24), .ZN(new_n692));
  OAI21_X1  g267(.A(new_n688), .B1(new_n692), .B2(G34), .ZN(new_n693));
  AOI21_X1  g268(.A(new_n693), .B1(new_n692), .B2(G34), .ZN(new_n694));
  AOI21_X1  g269(.A(new_n694), .B1(G160), .B2(G29), .ZN(new_n695));
  AOI22_X1  g270(.A1(new_n690), .A2(new_n691), .B1(new_n695), .B2(G2084), .ZN(new_n696));
  AND3_X1   g271(.A1(new_n678), .A2(new_n679), .A3(new_n696), .ZN(new_n697));
  NOR2_X1   g272(.A1(new_n697), .A2(KEYINPUT101), .ZN(new_n698));
  NAND2_X1  g273(.A1(new_n688), .A2(G35), .ZN(new_n699));
  OAI21_X1  g274(.A(new_n699), .B1(G162), .B2(new_n688), .ZN(new_n700));
  XNOR2_X1  g275(.A(new_n700), .B(KEYINPUT29), .ZN(new_n701));
  NOR2_X1   g276(.A1(new_n701), .A2(G2090), .ZN(new_n702));
  NAND2_X1  g277(.A1(new_n688), .A2(G26), .ZN(new_n703));
  XNOR2_X1  g278(.A(new_n703), .B(KEYINPUT28), .ZN(new_n704));
  OR2_X1    g279(.A1(G104), .A2(G2105), .ZN(new_n705));
  OAI211_X1 g280(.A(new_n705), .B(G2104), .C1(G116), .C2(new_n464), .ZN(new_n706));
  XOR2_X1   g281(.A(new_n706), .B(KEYINPUT97), .Z(new_n707));
  AOI21_X1  g282(.A(new_n707), .B1(G128), .B2(new_n482), .ZN(new_n708));
  NAND2_X1  g283(.A1(new_n673), .A2(G140), .ZN(new_n709));
  NAND2_X1  g284(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  INV_X1    g285(.A(new_n710), .ZN(new_n711));
  OAI21_X1  g286(.A(new_n704), .B1(new_n711), .B2(new_n688), .ZN(new_n712));
  XNOR2_X1  g287(.A(KEYINPUT98), .B(G2067), .ZN(new_n713));
  INV_X1    g288(.A(new_n713), .ZN(new_n714));
  INV_X1    g289(.A(G16), .ZN(new_n715));
  NAND2_X1  g290(.A1(new_n715), .A2(G5), .ZN(new_n716));
  OAI21_X1  g291(.A(new_n716), .B1(G171), .B2(new_n715), .ZN(new_n717));
  OAI22_X1  g292(.A1(new_n712), .A2(new_n714), .B1(G1961), .B2(new_n717), .ZN(new_n718));
  XNOR2_X1  g293(.A(KEYINPUT90), .B(G16), .ZN(new_n719));
  NOR2_X1   g294(.A1(new_n553), .A2(new_n719), .ZN(new_n720));
  AOI21_X1  g295(.A(new_n720), .B1(G19), .B2(new_n719), .ZN(new_n721));
  XOR2_X1   g296(.A(KEYINPUT96), .B(G1341), .Z(new_n722));
  INV_X1    g297(.A(new_n722), .ZN(new_n723));
  AOI22_X1  g298(.A1(new_n721), .A2(new_n723), .B1(G1961), .B2(new_n717), .ZN(new_n724));
  OAI221_X1 g299(.A(new_n724), .B1(new_n723), .B2(new_n721), .C1(new_n690), .C2(new_n691), .ZN(new_n725));
  AOI211_X1 g300(.A(new_n718), .B(new_n725), .C1(new_n712), .C2(new_n714), .ZN(new_n726));
  NAND2_X1  g301(.A1(new_n715), .A2(G4), .ZN(new_n727));
  OAI21_X1  g302(.A(new_n727), .B1(new_n596), .B2(new_n715), .ZN(new_n728));
  XOR2_X1   g303(.A(KEYINPUT95), .B(G1348), .Z(new_n729));
  XNOR2_X1  g304(.A(new_n728), .B(new_n729), .ZN(new_n730));
  XNOR2_X1  g305(.A(KEYINPUT31), .B(G11), .ZN(new_n731));
  XNOR2_X1  g306(.A(new_n731), .B(KEYINPUT102), .ZN(new_n732));
  INV_X1    g307(.A(G28), .ZN(new_n733));
  OR2_X1    g308(.A1(new_n733), .A2(KEYINPUT30), .ZN(new_n734));
  AOI21_X1  g309(.A(G29), .B1(new_n733), .B2(KEYINPUT30), .ZN(new_n735));
  AOI21_X1  g310(.A(new_n732), .B1(new_n734), .B2(new_n735), .ZN(new_n736));
  INV_X1    g311(.A(new_n614), .ZN(new_n737));
  NOR2_X1   g312(.A1(new_n737), .A2(new_n688), .ZN(new_n738));
  INV_X1    g313(.A(KEYINPUT103), .ZN(new_n739));
  OAI221_X1 g314(.A(new_n736), .B1(G2084), .B2(new_n695), .C1(new_n738), .C2(new_n739), .ZN(new_n740));
  NOR2_X1   g315(.A1(G164), .A2(new_n688), .ZN(new_n741));
  AOI21_X1  g316(.A(new_n741), .B1(G27), .B2(new_n688), .ZN(new_n742));
  NAND2_X1  g317(.A1(new_n742), .A2(new_n443), .ZN(new_n743));
  INV_X1    g318(.A(new_n738), .ZN(new_n744));
  OAI21_X1  g319(.A(new_n743), .B1(new_n744), .B2(KEYINPUT103), .ZN(new_n745));
  NAND2_X1  g320(.A1(new_n715), .A2(G21), .ZN(new_n746));
  OAI21_X1  g321(.A(new_n746), .B1(G168), .B2(new_n715), .ZN(new_n747));
  XNOR2_X1  g322(.A(new_n747), .B(G1966), .ZN(new_n748));
  NOR2_X1   g323(.A1(new_n742), .A2(new_n443), .ZN(new_n749));
  NOR4_X1   g324(.A1(new_n740), .A2(new_n745), .A3(new_n748), .A4(new_n749), .ZN(new_n750));
  NAND3_X1  g325(.A1(new_n726), .A2(new_n730), .A3(new_n750), .ZN(new_n751));
  NOR3_X1   g326(.A1(new_n698), .A2(new_n702), .A3(new_n751), .ZN(new_n752));
  NAND2_X1  g327(.A1(new_n701), .A2(G2090), .ZN(new_n753));
  XOR2_X1   g328(.A(KEYINPUT104), .B(KEYINPUT23), .Z(new_n754));
  XNOR2_X1  g329(.A(new_n754), .B(KEYINPUT105), .ZN(new_n755));
  NAND2_X1  g330(.A1(new_n719), .A2(G20), .ZN(new_n756));
  XNOR2_X1  g331(.A(new_n755), .B(new_n756), .ZN(new_n757));
  AOI21_X1  g332(.A(new_n757), .B1(G299), .B2(G16), .ZN(new_n758));
  AND2_X1   g333(.A1(new_n758), .A2(G1956), .ZN(new_n759));
  NOR2_X1   g334(.A1(new_n758), .A2(G1956), .ZN(new_n760));
  OAI21_X1  g335(.A(new_n753), .B1(new_n759), .B2(new_n760), .ZN(new_n761));
  OR2_X1    g336(.A1(new_n761), .A2(KEYINPUT106), .ZN(new_n762));
  NAND2_X1  g337(.A1(new_n697), .A2(KEYINPUT101), .ZN(new_n763));
  NAND2_X1  g338(.A1(new_n761), .A2(KEYINPUT106), .ZN(new_n764));
  NAND4_X1  g339(.A1(new_n752), .A2(new_n762), .A3(new_n763), .A4(new_n764), .ZN(new_n765));
  INV_X1    g340(.A(new_n719), .ZN(new_n766));
  NOR2_X1   g341(.A1(new_n766), .A2(G24), .ZN(new_n767));
  XNOR2_X1  g342(.A(G290), .B(KEYINPUT91), .ZN(new_n768));
  AOI21_X1  g343(.A(new_n767), .B1(new_n768), .B2(new_n766), .ZN(new_n769));
  XNOR2_X1  g344(.A(new_n769), .B(KEYINPUT92), .ZN(new_n770));
  INV_X1    g345(.A(G1986), .ZN(new_n771));
  XNOR2_X1  g346(.A(new_n770), .B(new_n771), .ZN(new_n772));
  NAND2_X1  g347(.A1(new_n688), .A2(G25), .ZN(new_n773));
  INV_X1    g348(.A(G131), .ZN(new_n774));
  NOR2_X1   g349(.A1(new_n464), .A2(G107), .ZN(new_n775));
  OAI21_X1  g350(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n776));
  OAI22_X1  g351(.A1(new_n493), .A2(new_n774), .B1(new_n775), .B2(new_n776), .ZN(new_n777));
  AOI21_X1  g352(.A(new_n777), .B1(G119), .B2(new_n482), .ZN(new_n778));
  OAI21_X1  g353(.A(new_n773), .B1(new_n778), .B2(new_n688), .ZN(new_n779));
  XOR2_X1   g354(.A(KEYINPUT35), .B(G1991), .Z(new_n780));
  XOR2_X1   g355(.A(new_n779), .B(new_n780), .Z(new_n781));
  NAND2_X1  g356(.A1(new_n715), .A2(G6), .ZN(new_n782));
  NOR2_X1   g357(.A1(new_n578), .A2(new_n582), .ZN(new_n783));
  OAI21_X1  g358(.A(new_n782), .B1(new_n783), .B2(new_n715), .ZN(new_n784));
  XOR2_X1   g359(.A(new_n784), .B(KEYINPUT93), .Z(new_n785));
  XNOR2_X1  g360(.A(KEYINPUT32), .B(G1981), .ZN(new_n786));
  INV_X1    g361(.A(new_n786), .ZN(new_n787));
  OR2_X1    g362(.A1(new_n785), .A2(new_n787), .ZN(new_n788));
  NAND2_X1  g363(.A1(new_n785), .A2(new_n787), .ZN(new_n789));
  NOR2_X1   g364(.A1(new_n766), .A2(G22), .ZN(new_n790));
  AOI21_X1  g365(.A(new_n790), .B1(G166), .B2(new_n766), .ZN(new_n791));
  INV_X1    g366(.A(G1971), .ZN(new_n792));
  XNOR2_X1  g367(.A(new_n791), .B(new_n792), .ZN(new_n793));
  NAND2_X1  g368(.A1(new_n715), .A2(G23), .ZN(new_n794));
  INV_X1    g369(.A(new_n573), .ZN(new_n795));
  OAI21_X1  g370(.A(new_n794), .B1(new_n795), .B2(new_n715), .ZN(new_n796));
  XNOR2_X1  g371(.A(KEYINPUT33), .B(G1976), .ZN(new_n797));
  XNOR2_X1  g372(.A(new_n796), .B(new_n797), .ZN(new_n798));
  NAND4_X1  g373(.A1(new_n788), .A2(new_n789), .A3(new_n793), .A4(new_n798), .ZN(new_n799));
  AOI21_X1  g374(.A(new_n781), .B1(new_n799), .B2(KEYINPUT34), .ZN(new_n800));
  OAI211_X1 g375(.A(new_n772), .B(new_n800), .C1(KEYINPUT34), .C2(new_n799), .ZN(new_n801));
  XNOR2_X1  g376(.A(KEYINPUT94), .B(KEYINPUT36), .ZN(new_n802));
  XNOR2_X1  g377(.A(new_n801), .B(new_n802), .ZN(new_n803));
  NOR2_X1   g378(.A1(new_n765), .A2(new_n803), .ZN(G311));
  INV_X1    g379(.A(G311), .ZN(G150));
  NAND2_X1  g380(.A1(new_n596), .A2(G559), .ZN(new_n806));
  INV_X1    g381(.A(G93), .ZN(new_n807));
  INV_X1    g382(.A(G55), .ZN(new_n808));
  OAI22_X1  g383(.A1(new_n522), .A2(new_n807), .B1(new_n524), .B2(new_n808), .ZN(new_n809));
  AOI22_X1  g384(.A1(new_n515), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n810));
  NOR2_X1   g385(.A1(new_n810), .A2(new_n516), .ZN(new_n811));
  OR2_X1    g386(.A1(new_n809), .A2(new_n811), .ZN(new_n812));
  INV_X1    g387(.A(KEYINPUT108), .ZN(new_n813));
  AOI21_X1  g388(.A(new_n553), .B1(new_n812), .B2(new_n813), .ZN(new_n814));
  OAI21_X1  g389(.A(new_n814), .B1(new_n813), .B2(new_n812), .ZN(new_n815));
  INV_X1    g390(.A(new_n812), .ZN(new_n816));
  NAND3_X1  g391(.A1(new_n816), .A2(KEYINPUT108), .A3(new_n553), .ZN(new_n817));
  NAND2_X1  g392(.A1(new_n815), .A2(new_n817), .ZN(new_n818));
  XNOR2_X1  g393(.A(new_n806), .B(new_n818), .ZN(new_n819));
  XOR2_X1   g394(.A(KEYINPUT107), .B(KEYINPUT38), .Z(new_n820));
  XNOR2_X1  g395(.A(new_n819), .B(new_n820), .ZN(new_n821));
  OR2_X1    g396(.A1(new_n821), .A2(KEYINPUT39), .ZN(new_n822));
  INV_X1    g397(.A(G860), .ZN(new_n823));
  NAND2_X1  g398(.A1(new_n821), .A2(KEYINPUT39), .ZN(new_n824));
  NAND3_X1  g399(.A1(new_n822), .A2(new_n823), .A3(new_n824), .ZN(new_n825));
  NAND2_X1  g400(.A1(new_n812), .A2(G860), .ZN(new_n826));
  XOR2_X1   g401(.A(new_n826), .B(KEYINPUT37), .Z(new_n827));
  NAND2_X1  g402(.A1(new_n825), .A2(new_n827), .ZN(G145));
  AOI21_X1  g403(.A(new_n496), .B1(new_n478), .B2(new_n479), .ZN(new_n829));
  NOR2_X1   g404(.A1(new_n464), .A2(G114), .ZN(new_n830));
  OAI21_X1  g405(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n831));
  NOR2_X1   g406(.A1(new_n830), .A2(new_n831), .ZN(new_n832));
  OAI21_X1  g407(.A(KEYINPUT109), .B1(new_n829), .B2(new_n832), .ZN(new_n833));
  INV_X1    g408(.A(KEYINPUT109), .ZN(new_n834));
  NAND3_X1  g409(.A1(new_n498), .A2(new_n503), .A3(new_n834), .ZN(new_n835));
  AOI21_X1  g410(.A(new_n507), .B1(new_n489), .B2(G138), .ZN(new_n836));
  NOR2_X1   g411(.A1(new_n505), .A2(KEYINPUT4), .ZN(new_n837));
  OAI211_X1 g412(.A(new_n833), .B(new_n835), .C1(new_n836), .C2(new_n837), .ZN(new_n838));
  XNOR2_X1  g413(.A(new_n710), .B(new_n838), .ZN(new_n839));
  XNOR2_X1  g414(.A(new_n839), .B(new_n686), .ZN(new_n840));
  MUX2_X1   g415(.A(new_n675), .B(new_n674), .S(new_n840), .Z(new_n841));
  XNOR2_X1  g416(.A(new_n778), .B(KEYINPUT110), .ZN(new_n842));
  XNOR2_X1  g417(.A(new_n842), .B(new_n619), .ZN(new_n843));
  NAND2_X1  g418(.A1(new_n673), .A2(G142), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n482), .A2(G130), .ZN(new_n845));
  NOR2_X1   g420(.A1(new_n464), .A2(G118), .ZN(new_n846));
  OAI21_X1  g421(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n847));
  OAI211_X1 g422(.A(new_n844), .B(new_n845), .C1(new_n846), .C2(new_n847), .ZN(new_n848));
  XOR2_X1   g423(.A(new_n843), .B(new_n848), .Z(new_n849));
  AND2_X1   g424(.A1(new_n841), .A2(new_n849), .ZN(new_n850));
  NOR2_X1   g425(.A1(new_n841), .A2(new_n849), .ZN(new_n851));
  XNOR2_X1  g426(.A(new_n614), .B(G160), .ZN(new_n852));
  XOR2_X1   g427(.A(new_n852), .B(G162), .Z(new_n853));
  OR3_X1    g428(.A1(new_n850), .A2(new_n851), .A3(new_n853), .ZN(new_n854));
  XNOR2_X1  g429(.A(new_n841), .B(new_n849), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n855), .A2(new_n853), .ZN(new_n856));
  INV_X1    g431(.A(G37), .ZN(new_n857));
  NAND3_X1  g432(.A1(new_n854), .A2(new_n856), .A3(new_n857), .ZN(new_n858));
  XNOR2_X1  g433(.A(new_n858), .B(KEYINPUT40), .ZN(G395));
  NOR2_X1   g434(.A1(new_n812), .A2(G868), .ZN(new_n860));
  XNOR2_X1  g435(.A(G290), .B(new_n783), .ZN(new_n861));
  XNOR2_X1  g436(.A(G166), .B(new_n573), .ZN(new_n862));
  XOR2_X1   g437(.A(new_n861), .B(new_n862), .Z(new_n863));
  AND2_X1   g438(.A1(KEYINPUT111), .A2(KEYINPUT42), .ZN(new_n864));
  NOR2_X1   g439(.A1(KEYINPUT111), .A2(KEYINPUT42), .ZN(new_n865));
  OAI21_X1  g440(.A(new_n863), .B1(new_n864), .B2(new_n865), .ZN(new_n866));
  OAI21_X1  g441(.A(new_n866), .B1(new_n863), .B2(new_n865), .ZN(new_n867));
  XNOR2_X1  g442(.A(new_n604), .B(new_n818), .ZN(new_n868));
  XNOR2_X1  g443(.A(new_n595), .B(G299), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  XNOR2_X1  g445(.A(new_n869), .B(KEYINPUT41), .ZN(new_n871));
  OAI21_X1  g446(.A(new_n870), .B1(new_n871), .B2(new_n868), .ZN(new_n872));
  INV_X1    g447(.A(KEYINPUT112), .ZN(new_n873));
  AOI21_X1  g448(.A(new_n867), .B1(new_n872), .B2(new_n873), .ZN(new_n874));
  NOR2_X1   g449(.A1(new_n872), .A2(new_n873), .ZN(new_n875));
  XOR2_X1   g450(.A(new_n874), .B(new_n875), .Z(new_n876));
  AOI21_X1  g451(.A(new_n860), .B1(new_n876), .B2(G868), .ZN(G295));
  AOI21_X1  g452(.A(new_n860), .B1(new_n876), .B2(G868), .ZN(G331));
  INV_X1    g453(.A(KEYINPUT44), .ZN(new_n879));
  NOR2_X1   g454(.A1(G168), .A2(G171), .ZN(new_n880));
  AOI21_X1  g455(.A(new_n880), .B1(new_n564), .B2(G168), .ZN(new_n881));
  OR2_X1    g456(.A1(new_n818), .A2(new_n881), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n818), .A2(new_n881), .ZN(new_n883));
  NAND3_X1  g458(.A1(new_n871), .A2(new_n882), .A3(new_n883), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n882), .A2(new_n883), .ZN(new_n885));
  INV_X1    g460(.A(new_n869), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n884), .A2(new_n887), .ZN(new_n888));
  INV_X1    g463(.A(KEYINPUT113), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  AND2_X1   g465(.A1(new_n882), .A2(new_n883), .ZN(new_n891));
  AOI21_X1  g466(.A(new_n889), .B1(new_n891), .B2(new_n871), .ZN(new_n892));
  INV_X1    g467(.A(new_n892), .ZN(new_n893));
  NAND3_X1  g468(.A1(new_n890), .A2(KEYINPUT114), .A3(new_n893), .ZN(new_n894));
  INV_X1    g469(.A(KEYINPUT114), .ZN(new_n895));
  AOI21_X1  g470(.A(KEYINPUT113), .B1(new_n884), .B2(new_n887), .ZN(new_n896));
  OAI21_X1  g471(.A(new_n895), .B1(new_n896), .B2(new_n892), .ZN(new_n897));
  NAND3_X1  g472(.A1(new_n894), .A2(new_n897), .A3(new_n863), .ZN(new_n898));
  INV_X1    g473(.A(KEYINPUT43), .ZN(new_n899));
  INV_X1    g474(.A(new_n863), .ZN(new_n900));
  NAND3_X1  g475(.A1(new_n890), .A2(new_n900), .A3(new_n893), .ZN(new_n901));
  NAND4_X1  g476(.A1(new_n898), .A2(new_n899), .A3(new_n857), .A4(new_n901), .ZN(new_n902));
  AOI21_X1  g477(.A(G37), .B1(new_n888), .B2(new_n863), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n901), .A2(new_n903), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n904), .A2(KEYINPUT43), .ZN(new_n905));
  AOI21_X1  g480(.A(new_n879), .B1(new_n902), .B2(new_n905), .ZN(new_n906));
  AND3_X1   g481(.A1(new_n901), .A2(new_n899), .A3(new_n903), .ZN(new_n907));
  NAND3_X1  g482(.A1(new_n898), .A2(new_n857), .A3(new_n901), .ZN(new_n908));
  AOI21_X1  g483(.A(new_n907), .B1(new_n908), .B2(KEYINPUT43), .ZN(new_n909));
  AOI21_X1  g484(.A(new_n906), .B1(new_n909), .B2(new_n879), .ZN(G397));
  XOR2_X1   g485(.A(KEYINPUT115), .B(G1384), .Z(new_n911));
  NAND2_X1  g486(.A1(new_n838), .A2(new_n911), .ZN(new_n912));
  XNOR2_X1  g487(.A(KEYINPUT116), .B(KEYINPUT45), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  NAND2_X1  g489(.A1(G160), .A2(G40), .ZN(new_n915));
  NOR2_X1   g490(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  INV_X1    g491(.A(new_n916), .ZN(new_n917));
  INV_X1    g492(.A(G2067), .ZN(new_n918));
  XNOR2_X1  g493(.A(new_n710), .B(new_n918), .ZN(new_n919));
  INV_X1    g494(.A(G1996), .ZN(new_n920));
  XNOR2_X1  g495(.A(new_n686), .B(new_n920), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n919), .A2(new_n921), .ZN(new_n922));
  XNOR2_X1  g497(.A(new_n778), .B(new_n780), .ZN(new_n923));
  NOR2_X1   g498(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  XNOR2_X1  g499(.A(G290), .B(new_n771), .ZN(new_n925));
  AOI21_X1  g500(.A(new_n917), .B1(new_n924), .B2(new_n925), .ZN(new_n926));
  INV_X1    g501(.A(KEYINPUT50), .ZN(new_n927));
  INV_X1    g502(.A(G1384), .ZN(new_n928));
  NAND3_X1  g503(.A1(new_n838), .A2(new_n927), .A3(new_n928), .ZN(new_n929));
  INV_X1    g504(.A(G40), .ZN(new_n930));
  AOI211_X1 g505(.A(new_n930), .B(new_n470), .C1(new_n476), .C2(G2105), .ZN(new_n931));
  INV_X1    g506(.A(G2084), .ZN(new_n932));
  OAI21_X1  g507(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n933));
  NAND4_X1  g508(.A1(new_n929), .A2(new_n931), .A3(new_n932), .A4(new_n933), .ZN(new_n934));
  XNOR2_X1  g509(.A(new_n934), .B(KEYINPUT119), .ZN(new_n935));
  AOI21_X1  g510(.A(KEYINPUT45), .B1(new_n838), .B2(new_n928), .ZN(new_n936));
  OAI21_X1  g511(.A(KEYINPUT118), .B1(new_n936), .B2(new_n915), .ZN(new_n937));
  INV_X1    g512(.A(KEYINPUT118), .ZN(new_n938));
  AND3_X1   g513(.A1(new_n498), .A2(new_n503), .A3(new_n834), .ZN(new_n939));
  AOI21_X1  g514(.A(new_n834), .B1(new_n498), .B2(new_n503), .ZN(new_n940));
  NOR2_X1   g515(.A1(new_n939), .A2(new_n940), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n506), .A2(new_n508), .ZN(new_n942));
  AOI21_X1  g517(.A(G1384), .B1(new_n941), .B2(new_n942), .ZN(new_n943));
  OAI211_X1 g518(.A(new_n938), .B(new_n931), .C1(new_n943), .C2(KEYINPUT45), .ZN(new_n944));
  OR3_X1    g519(.A1(G164), .A2(G1384), .A3(new_n913), .ZN(new_n945));
  NAND3_X1  g520(.A1(new_n937), .A2(new_n944), .A3(new_n945), .ZN(new_n946));
  INV_X1    g521(.A(G1966), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n935), .A2(new_n948), .ZN(new_n949));
  INV_X1    g524(.A(G8), .ZN(new_n950));
  NOR2_X1   g525(.A1(G168), .A2(new_n950), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n949), .A2(new_n951), .ZN(new_n952));
  AOI21_X1  g527(.A(new_n950), .B1(new_n935), .B2(new_n948), .ZN(new_n953));
  NOR3_X1   g528(.A1(new_n953), .A2(KEYINPUT51), .A3(new_n951), .ZN(new_n954));
  INV_X1    g529(.A(new_n954), .ZN(new_n955));
  INV_X1    g530(.A(KEYINPUT51), .ZN(new_n956));
  AOI21_X1  g531(.A(new_n951), .B1(new_n953), .B2(KEYINPUT123), .ZN(new_n957));
  INV_X1    g532(.A(new_n945), .ZN(new_n958));
  NOR2_X1   g533(.A1(new_n936), .A2(new_n915), .ZN(new_n959));
  AOI21_X1  g534(.A(new_n958), .B1(new_n959), .B2(new_n938), .ZN(new_n960));
  AOI21_X1  g535(.A(G1966), .B1(new_n960), .B2(new_n937), .ZN(new_n961));
  INV_X1    g536(.A(KEYINPUT119), .ZN(new_n962));
  XNOR2_X1  g537(.A(new_n934), .B(new_n962), .ZN(new_n963));
  OAI21_X1  g538(.A(G8), .B1(new_n961), .B2(new_n963), .ZN(new_n964));
  INV_X1    g539(.A(KEYINPUT123), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n964), .A2(new_n965), .ZN(new_n966));
  AOI21_X1  g541(.A(new_n956), .B1(new_n957), .B2(new_n966), .ZN(new_n967));
  OAI21_X1  g542(.A(new_n955), .B1(new_n967), .B2(KEYINPUT124), .ZN(new_n968));
  OAI211_X1 g543(.A(KEYINPUT123), .B(G8), .C1(new_n961), .C2(new_n963), .ZN(new_n969));
  INV_X1    g544(.A(new_n951), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n969), .A2(new_n970), .ZN(new_n971));
  NOR2_X1   g546(.A1(new_n953), .A2(KEYINPUT123), .ZN(new_n972));
  OAI21_X1  g547(.A(KEYINPUT51), .B1(new_n971), .B2(new_n972), .ZN(new_n973));
  INV_X1    g548(.A(KEYINPUT124), .ZN(new_n974));
  NOR2_X1   g549(.A1(new_n973), .A2(new_n974), .ZN(new_n975));
  OAI21_X1  g550(.A(new_n952), .B1(new_n968), .B2(new_n975), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n976), .A2(KEYINPUT62), .ZN(new_n977));
  INV_X1    g552(.A(KEYINPUT62), .ZN(new_n978));
  OAI211_X1 g553(.A(new_n978), .B(new_n952), .C1(new_n968), .C2(new_n975), .ZN(new_n979));
  INV_X1    g554(.A(KEYINPUT49), .ZN(new_n980));
  INV_X1    g555(.A(G1981), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n783), .A2(new_n981), .ZN(new_n982));
  INV_X1    g557(.A(new_n982), .ZN(new_n983));
  NOR2_X1   g558(.A1(new_n783), .A2(new_n981), .ZN(new_n984));
  OAI21_X1  g559(.A(new_n980), .B1(new_n983), .B2(new_n984), .ZN(new_n985));
  NAND2_X1  g560(.A1(G305), .A2(G1981), .ZN(new_n986));
  NAND3_X1  g561(.A1(new_n986), .A2(KEYINPUT49), .A3(new_n982), .ZN(new_n987));
  AND2_X1   g562(.A1(new_n943), .A2(new_n931), .ZN(new_n988));
  NOR2_X1   g563(.A1(new_n988), .A2(new_n950), .ZN(new_n989));
  NAND3_X1  g564(.A1(new_n985), .A2(new_n987), .A3(new_n989), .ZN(new_n990));
  INV_X1    g565(.A(KEYINPUT117), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n990), .A2(new_n991), .ZN(new_n992));
  NAND4_X1  g567(.A1(new_n985), .A2(new_n987), .A3(KEYINPUT117), .A4(new_n989), .ZN(new_n993));
  NAND2_X1  g568(.A1(new_n992), .A2(new_n993), .ZN(new_n994));
  INV_X1    g569(.A(KEYINPUT52), .ZN(new_n995));
  OAI21_X1  g570(.A(new_n995), .B1(new_n574), .B2(G1976), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n795), .A2(G1976), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n989), .A2(new_n997), .ZN(new_n998));
  NOR2_X1   g573(.A1(new_n996), .A2(new_n998), .ZN(new_n999));
  AOI21_X1  g574(.A(new_n995), .B1(new_n989), .B2(new_n997), .ZN(new_n1000));
  NOR2_X1   g575(.A1(new_n999), .A2(new_n1000), .ZN(new_n1001));
  NAND3_X1  g576(.A1(new_n567), .A2(G8), .A3(new_n568), .ZN(new_n1002));
  XNOR2_X1  g577(.A(new_n1002), .B(KEYINPUT55), .ZN(new_n1003));
  OR3_X1    g578(.A1(G164), .A2(KEYINPUT50), .A3(G1384), .ZN(new_n1004));
  OAI211_X1 g579(.A(new_n1004), .B(new_n931), .C1(new_n927), .C2(new_n943), .ZN(new_n1005));
  NOR2_X1   g580(.A1(new_n1005), .A2(G2090), .ZN(new_n1006));
  NAND3_X1  g581(.A1(new_n838), .A2(KEYINPUT45), .A3(new_n911), .ZN(new_n1007));
  OAI21_X1  g582(.A(new_n913), .B1(G164), .B2(G1384), .ZN(new_n1008));
  NAND3_X1  g583(.A1(new_n1007), .A2(new_n931), .A3(new_n1008), .ZN(new_n1009));
  AOI21_X1  g584(.A(new_n1006), .B1(new_n792), .B2(new_n1009), .ZN(new_n1010));
  OAI21_X1  g585(.A(new_n1003), .B1(new_n1010), .B2(new_n950), .ZN(new_n1011));
  INV_X1    g586(.A(KEYINPUT55), .ZN(new_n1012));
  XNOR2_X1  g587(.A(new_n1002), .B(new_n1012), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n1009), .A2(new_n792), .ZN(new_n1014));
  NAND3_X1  g589(.A1(new_n929), .A2(new_n931), .A3(new_n933), .ZN(new_n1015));
  OAI21_X1  g590(.A(new_n1014), .B1(G2090), .B2(new_n1015), .ZN(new_n1016));
  NAND3_X1  g591(.A1(new_n1013), .A2(new_n1016), .A3(G8), .ZN(new_n1017));
  NAND4_X1  g592(.A1(new_n994), .A2(new_n1001), .A3(new_n1011), .A4(new_n1017), .ZN(new_n1018));
  OR2_X1    g593(.A1(new_n1009), .A2(G2078), .ZN(new_n1019));
  INV_X1    g594(.A(KEYINPUT53), .ZN(new_n1020));
  INV_X1    g595(.A(G1961), .ZN(new_n1021));
  AOI22_X1  g596(.A1(new_n1019), .A2(new_n1020), .B1(new_n1021), .B2(new_n1015), .ZN(new_n1022));
  NOR2_X1   g597(.A1(new_n1020), .A2(G2078), .ZN(new_n1023));
  NAND3_X1  g598(.A1(new_n960), .A2(new_n937), .A3(new_n1023), .ZN(new_n1024));
  AOI21_X1  g599(.A(G301), .B1(new_n1022), .B2(new_n1024), .ZN(new_n1025));
  INV_X1    g600(.A(new_n1025), .ZN(new_n1026));
  NOR2_X1   g601(.A1(new_n1018), .A2(new_n1026), .ZN(new_n1027));
  NAND3_X1  g602(.A1(new_n977), .A2(new_n979), .A3(new_n1027), .ZN(new_n1028));
  INV_X1    g603(.A(KEYINPUT63), .ZN(new_n1029));
  NOR2_X1   g604(.A1(new_n964), .A2(G286), .ZN(new_n1030));
  INV_X1    g605(.A(new_n1030), .ZN(new_n1031));
  OAI21_X1  g606(.A(new_n1029), .B1(new_n1018), .B2(new_n1031), .ZN(new_n1032));
  AND2_X1   g607(.A1(new_n994), .A2(new_n1001), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n1016), .A2(G8), .ZN(new_n1034));
  AOI21_X1  g609(.A(new_n1029), .B1(new_n1003), .B2(new_n1034), .ZN(new_n1035));
  NAND4_X1  g610(.A1(new_n1033), .A2(new_n1017), .A3(new_n1030), .A4(new_n1035), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n1032), .A2(new_n1036), .ZN(new_n1037));
  NOR2_X1   g612(.A1(G288), .A2(G1976), .ZN(new_n1038));
  AOI21_X1  g613(.A(new_n983), .B1(new_n994), .B2(new_n1038), .ZN(new_n1039));
  INV_X1    g614(.A(new_n989), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n994), .A2(new_n1001), .ZN(new_n1041));
  OAI22_X1  g616(.A1(new_n1039), .A2(new_n1040), .B1(new_n1041), .B2(new_n1017), .ZN(new_n1042));
  INV_X1    g617(.A(new_n1042), .ZN(new_n1043));
  NAND2_X1  g618(.A1(new_n1037), .A2(new_n1043), .ZN(new_n1044));
  OR2_X1    g619(.A1(G299), .A2(KEYINPUT57), .ZN(new_n1045));
  NAND2_X1  g620(.A1(G299), .A2(KEYINPUT57), .ZN(new_n1046));
  INV_X1    g621(.A(G1956), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n1005), .A2(new_n1047), .ZN(new_n1048));
  XNOR2_X1  g623(.A(KEYINPUT56), .B(G2072), .ZN(new_n1049));
  NAND4_X1  g624(.A1(new_n1007), .A2(new_n931), .A3(new_n1008), .A4(new_n1049), .ZN(new_n1050));
  AOI22_X1  g625(.A1(new_n1045), .A2(new_n1046), .B1(new_n1048), .B2(new_n1050), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n988), .A2(new_n918), .ZN(new_n1052));
  INV_X1    g627(.A(G1348), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n1015), .A2(new_n1053), .ZN(new_n1054));
  AND2_X1   g629(.A1(new_n1052), .A2(new_n1054), .ZN(new_n1055));
  NOR2_X1   g630(.A1(new_n1055), .A2(new_n595), .ZN(new_n1056));
  NAND4_X1  g631(.A1(new_n1045), .A2(new_n1046), .A3(new_n1048), .A4(new_n1050), .ZN(new_n1057));
  AOI21_X1  g632(.A(new_n1051), .B1(new_n1056), .B2(new_n1057), .ZN(new_n1058));
  INV_X1    g633(.A(KEYINPUT61), .ZN(new_n1059));
  INV_X1    g634(.A(new_n1057), .ZN(new_n1060));
  OAI21_X1  g635(.A(new_n1059), .B1(new_n1060), .B2(new_n1051), .ZN(new_n1061));
  NAND2_X1  g636(.A1(new_n1045), .A2(new_n1046), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n1048), .A2(new_n1050), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n1062), .A2(new_n1063), .ZN(new_n1064));
  NAND3_X1  g639(.A1(new_n1064), .A2(KEYINPUT61), .A3(new_n1057), .ZN(new_n1065));
  AND3_X1   g640(.A1(new_n1052), .A2(new_n595), .A3(new_n1054), .ZN(new_n1066));
  OAI21_X1  g641(.A(KEYINPUT60), .B1(new_n1056), .B2(new_n1066), .ZN(new_n1067));
  NOR2_X1   g642(.A1(new_n595), .A2(KEYINPUT60), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n1055), .A2(new_n1068), .ZN(new_n1069));
  NAND4_X1  g644(.A1(new_n1061), .A2(new_n1065), .A3(new_n1067), .A4(new_n1069), .ZN(new_n1070));
  NAND4_X1  g645(.A1(new_n1007), .A2(new_n931), .A3(new_n920), .A4(new_n1008), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n1071), .A2(KEYINPUT120), .ZN(new_n1072));
  XOR2_X1   g647(.A(KEYINPUT121), .B(KEYINPUT58), .Z(new_n1073));
  XOR2_X1   g648(.A(new_n1073), .B(G1341), .Z(new_n1074));
  OAI21_X1  g649(.A(new_n1072), .B1(new_n988), .B2(new_n1074), .ZN(new_n1075));
  NOR2_X1   g650(.A1(new_n1071), .A2(KEYINPUT120), .ZN(new_n1076));
  OAI21_X1  g651(.A(new_n553), .B1(new_n1075), .B2(new_n1076), .ZN(new_n1077));
  NOR2_X1   g652(.A1(KEYINPUT122), .A2(KEYINPUT59), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n1077), .A2(new_n1078), .ZN(new_n1079));
  OAI221_X1 g654(.A(new_n553), .B1(KEYINPUT122), .B2(KEYINPUT59), .C1(new_n1075), .C2(new_n1076), .ZN(new_n1080));
  AOI22_X1  g655(.A1(new_n1079), .A2(new_n1080), .B1(KEYINPUT122), .B2(KEYINPUT59), .ZN(new_n1081));
  OAI21_X1  g656(.A(new_n1058), .B1(new_n1070), .B2(new_n1081), .ZN(new_n1082));
  INV_X1    g657(.A(new_n1018), .ZN(new_n1083));
  INV_X1    g658(.A(KEYINPUT54), .ZN(new_n1084));
  NAND4_X1  g659(.A1(new_n914), .A2(new_n931), .A3(new_n1007), .A4(new_n1023), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n1022), .A2(new_n1085), .ZN(new_n1086));
  OAI211_X1 g661(.A(new_n1026), .B(new_n1084), .C1(new_n564), .C2(new_n1086), .ZN(new_n1087));
  NAND2_X1  g662(.A1(new_n1086), .A2(G171), .ZN(new_n1088));
  NAND3_X1  g663(.A1(new_n1022), .A2(G301), .A3(new_n1024), .ZN(new_n1089));
  AND2_X1   g664(.A1(new_n1088), .A2(new_n1089), .ZN(new_n1090));
  OAI21_X1  g665(.A(new_n1087), .B1(new_n1090), .B2(new_n1084), .ZN(new_n1091));
  NAND3_X1  g666(.A1(new_n1082), .A2(new_n1083), .A3(new_n1091), .ZN(new_n1092));
  INV_X1    g667(.A(new_n1092), .ZN(new_n1093));
  AOI21_X1  g668(.A(new_n1044), .B1(new_n1093), .B2(new_n976), .ZN(new_n1094));
  AOI21_X1  g669(.A(new_n926), .B1(new_n1028), .B2(new_n1094), .ZN(new_n1095));
  AOI21_X1  g670(.A(new_n917), .B1(new_n919), .B2(new_n687), .ZN(new_n1096));
  OAI21_X1  g671(.A(KEYINPUT46), .B1(new_n917), .B2(G1996), .ZN(new_n1097));
  OR3_X1    g672(.A1(new_n917), .A2(KEYINPUT46), .A3(G1996), .ZN(new_n1098));
  AOI21_X1  g673(.A(new_n1096), .B1(new_n1097), .B2(new_n1098), .ZN(new_n1099));
  XNOR2_X1  g674(.A(new_n1099), .B(KEYINPUT47), .ZN(new_n1100));
  NOR3_X1   g675(.A1(new_n917), .A2(G1986), .A3(G290), .ZN(new_n1101));
  XOR2_X1   g676(.A(KEYINPUT125), .B(KEYINPUT48), .Z(new_n1102));
  XNOR2_X1  g677(.A(new_n1102), .B(KEYINPUT126), .ZN(new_n1103));
  XNOR2_X1  g678(.A(new_n1101), .B(new_n1103), .ZN(new_n1104));
  OAI21_X1  g679(.A(new_n1104), .B1(new_n924), .B2(new_n917), .ZN(new_n1105));
  AND4_X1   g680(.A1(new_n780), .A2(new_n919), .A3(new_n778), .A4(new_n921), .ZN(new_n1106));
  AOI21_X1  g681(.A(new_n1106), .B1(new_n918), .B2(new_n711), .ZN(new_n1107));
  OAI21_X1  g682(.A(new_n1105), .B1(new_n1107), .B2(new_n917), .ZN(new_n1108));
  NOR2_X1   g683(.A1(new_n1100), .A2(new_n1108), .ZN(new_n1109));
  INV_X1    g684(.A(new_n1109), .ZN(new_n1110));
  OAI21_X1  g685(.A(KEYINPUT127), .B1(new_n1095), .B2(new_n1110), .ZN(new_n1111));
  INV_X1    g686(.A(KEYINPUT127), .ZN(new_n1112));
  AOI21_X1  g687(.A(new_n1042), .B1(new_n1032), .B2(new_n1036), .ZN(new_n1113));
  INV_X1    g688(.A(new_n952), .ZN(new_n1114));
  AOI21_X1  g689(.A(new_n954), .B1(new_n973), .B2(new_n974), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n967), .A2(KEYINPUT124), .ZN(new_n1116));
  AOI21_X1  g691(.A(new_n1114), .B1(new_n1115), .B2(new_n1116), .ZN(new_n1117));
  OAI21_X1  g692(.A(new_n1113), .B1(new_n1117), .B2(new_n1092), .ZN(new_n1118));
  INV_X1    g693(.A(new_n1027), .ZN(new_n1119));
  AOI21_X1  g694(.A(new_n1119), .B1(new_n976), .B2(KEYINPUT62), .ZN(new_n1120));
  AOI21_X1  g695(.A(new_n1118), .B1(new_n979), .B2(new_n1120), .ZN(new_n1121));
  OAI211_X1 g696(.A(new_n1112), .B(new_n1109), .C1(new_n1121), .C2(new_n926), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n1111), .A2(new_n1122), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g698(.A(G319), .ZN(new_n1125));
  NOR3_X1   g699(.A1(G401), .A2(new_n1125), .A3(G227), .ZN(new_n1126));
  AND2_X1   g700(.A1(new_n667), .A2(new_n1126), .ZN(new_n1127));
  NAND2_X1  g701(.A1(new_n858), .A2(new_n1127), .ZN(new_n1128));
  NOR2_X1   g702(.A1(new_n1128), .A2(new_n909), .ZN(G308));
  OR2_X1    g703(.A1(new_n1128), .A2(new_n909), .ZN(G225));
endmodule


