//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 1 1 1 0 0 0 1 1 1 0 1 1 1 0 1 1 1 1 0 1 0 0 1 1 1 0 1 1 0 0 0 1 1 1 0 1 1 0 0 0 1 1 0 0 1 0 0 0 1 1 1 0 1 1 0 1 0 1 1 1 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:29:55 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n443, new_n446, new_n448, new_n452, new_n453, new_n454, new_n457,
    new_n458, new_n459, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n527, new_n528, new_n529, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n544, new_n545, new_n546, new_n547, new_n548, new_n549,
    new_n552, new_n553, new_n554, new_n556, new_n557, new_n558, new_n559,
    new_n560, new_n561, new_n562, new_n563, new_n564, new_n565, new_n566,
    new_n570, new_n571, new_n572, new_n573, new_n575, new_n576, new_n577,
    new_n578, new_n579, new_n580, new_n581, new_n582, new_n583, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n606, new_n609, new_n610, new_n612,
    new_n613, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1217, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1234, new_n1235, new_n1236;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  XNOR2_X1  g003(.A(KEYINPUT64), .B(G1083), .ZN(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  XNOR2_X1  g008(.A(KEYINPUT65), .B(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(new_n443));
  XNOR2_X1  g018(.A(new_n443), .B(KEYINPUT66), .ZN(G259));
  XNOR2_X1  g019(.A(KEYINPUT67), .B(G452), .ZN(G391));
  NAND2_X1  g020(.A1(G94), .A2(G452), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT68), .Z(G173));
  NAND2_X1  g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XOR2_X1   g023(.A(new_n448), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g024(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g025(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g026(.A1(G218), .A2(G220), .A3(G221), .A4(G219), .ZN(new_n452));
  XOR2_X1   g027(.A(new_n452), .B(KEYINPUT2), .Z(new_n453));
  NAND4_X1  g028(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n454));
  NOR2_X1   g029(.A1(new_n453), .A2(new_n454), .ZN(G325));
  INV_X1    g030(.A(G325), .ZN(G261));
  NAND2_X1  g031(.A1(new_n453), .A2(G2106), .ZN(new_n457));
  NAND2_X1  g032(.A1(new_n454), .A2(G567), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  INV_X1    g034(.A(new_n459), .ZN(G319));
  INV_X1    g035(.A(G125), .ZN(new_n461));
  OR2_X1    g036(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n462));
  NAND2_X1  g037(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n463));
  AOI21_X1  g038(.A(new_n461), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  AND2_X1   g039(.A1(G113), .A2(G2104), .ZN(new_n465));
  OAI21_X1  g040(.A(G2105), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  INV_X1    g041(.A(G2105), .ZN(new_n467));
  AND3_X1   g042(.A1(new_n467), .A2(G101), .A3(G2104), .ZN(new_n468));
  AOI21_X1  g043(.A(G2105), .B1(new_n462), .B2(new_n463), .ZN(new_n469));
  AOI21_X1  g044(.A(new_n468), .B1(new_n469), .B2(G137), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n466), .A2(new_n470), .ZN(new_n471));
  INV_X1    g046(.A(new_n471), .ZN(G160));
  NAND2_X1  g047(.A1(new_n469), .A2(KEYINPUT69), .ZN(new_n473));
  INV_X1    g048(.A(KEYINPUT69), .ZN(new_n474));
  AND2_X1   g049(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n475));
  NOR2_X1   g050(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n476));
  NOR2_X1   g051(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  OAI21_X1  g052(.A(new_n474), .B1(new_n477), .B2(G2105), .ZN(new_n478));
  AND2_X1   g053(.A1(new_n473), .A2(new_n478), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n479), .A2(G136), .ZN(new_n480));
  OAI21_X1  g055(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n481));
  INV_X1    g056(.A(G112), .ZN(new_n482));
  AOI21_X1  g057(.A(new_n481), .B1(new_n482), .B2(G2105), .ZN(new_n483));
  NOR2_X1   g058(.A1(new_n477), .A2(new_n467), .ZN(new_n484));
  AOI21_X1  g059(.A(new_n483), .B1(new_n484), .B2(G124), .ZN(new_n485));
  NAND2_X1  g060(.A1(new_n480), .A2(new_n485), .ZN(new_n486));
  INV_X1    g061(.A(new_n486), .ZN(G162));
  OAI21_X1  g062(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n488));
  INV_X1    g063(.A(G114), .ZN(new_n489));
  AOI21_X1  g064(.A(new_n488), .B1(new_n489), .B2(G2105), .ZN(new_n490));
  AND2_X1   g065(.A1(G126), .A2(G2105), .ZN(new_n491));
  OAI21_X1  g066(.A(new_n491), .B1(new_n475), .B2(new_n476), .ZN(new_n492));
  INV_X1    g067(.A(KEYINPUT70), .ZN(new_n493));
  NAND2_X1  g068(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  OAI211_X1 g069(.A(KEYINPUT70), .B(new_n491), .C1(new_n475), .C2(new_n476), .ZN(new_n495));
  AOI21_X1  g070(.A(new_n490), .B1(new_n494), .B2(new_n495), .ZN(new_n496));
  OAI211_X1 g071(.A(G138), .B(new_n467), .C1(new_n475), .C2(new_n476), .ZN(new_n497));
  NAND2_X1  g072(.A1(new_n497), .A2(KEYINPUT4), .ZN(new_n498));
  XNOR2_X1  g073(.A(KEYINPUT3), .B(G2104), .ZN(new_n499));
  INV_X1    g074(.A(KEYINPUT4), .ZN(new_n500));
  NAND4_X1  g075(.A1(new_n499), .A2(new_n500), .A3(G138), .A4(new_n467), .ZN(new_n501));
  NAND2_X1  g076(.A1(new_n498), .A2(new_n501), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n496), .A2(new_n502), .ZN(new_n503));
  INV_X1    g078(.A(new_n503), .ZN(G164));
  INV_X1    g079(.A(G62), .ZN(new_n505));
  OR2_X1    g080(.A1(KEYINPUT5), .A2(G543), .ZN(new_n506));
  NAND2_X1  g081(.A1(KEYINPUT5), .A2(G543), .ZN(new_n507));
  AOI21_X1  g082(.A(new_n505), .B1(new_n506), .B2(new_n507), .ZN(new_n508));
  AND2_X1   g083(.A1(G75), .A2(G543), .ZN(new_n509));
  OAI21_X1  g084(.A(G651), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n506), .A2(new_n507), .ZN(new_n511));
  OR2_X1    g086(.A1(KEYINPUT6), .A2(G651), .ZN(new_n512));
  NAND2_X1  g087(.A1(KEYINPUT6), .A2(G651), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  XNOR2_X1  g089(.A(KEYINPUT72), .B(G88), .ZN(new_n515));
  NAND3_X1  g090(.A1(new_n511), .A2(new_n514), .A3(new_n515), .ZN(new_n516));
  INV_X1    g091(.A(G543), .ZN(new_n517));
  AOI21_X1  g092(.A(new_n517), .B1(new_n512), .B2(new_n513), .ZN(new_n518));
  AOI21_X1  g093(.A(KEYINPUT71), .B1(new_n518), .B2(G50), .ZN(new_n519));
  AND2_X1   g094(.A1(KEYINPUT6), .A2(G651), .ZN(new_n520));
  NOR2_X1   g095(.A1(KEYINPUT6), .A2(G651), .ZN(new_n521));
  OAI211_X1 g096(.A(G50), .B(G543), .C1(new_n520), .C2(new_n521), .ZN(new_n522));
  INV_X1    g097(.A(KEYINPUT71), .ZN(new_n523));
  NOR2_X1   g098(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  OAI211_X1 g099(.A(new_n510), .B(new_n516), .C1(new_n519), .C2(new_n524), .ZN(G303));
  INV_X1    g100(.A(G303), .ZN(G166));
  NAND3_X1  g101(.A1(new_n511), .A2(G63), .A3(G651), .ZN(new_n527));
  NAND2_X1  g102(.A1(new_n518), .A2(G51), .ZN(new_n528));
  NAND3_X1  g103(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n529));
  XNOR2_X1  g104(.A(new_n529), .B(KEYINPUT7), .ZN(new_n530));
  NAND2_X1  g105(.A1(new_n511), .A2(new_n514), .ZN(new_n531));
  INV_X1    g106(.A(G89), .ZN(new_n532));
  OAI21_X1  g107(.A(new_n530), .B1(new_n531), .B2(new_n532), .ZN(new_n533));
  OAI211_X1 g108(.A(new_n527), .B(new_n528), .C1(new_n533), .C2(KEYINPUT73), .ZN(new_n534));
  AND2_X1   g109(.A1(new_n533), .A2(KEYINPUT73), .ZN(new_n535));
  NOR2_X1   g110(.A1(new_n534), .A2(new_n535), .ZN(G168));
  AOI22_X1  g111(.A1(new_n511), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n537));
  INV_X1    g112(.A(G651), .ZN(new_n538));
  NOR2_X1   g113(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  NAND2_X1  g114(.A1(new_n518), .A2(G52), .ZN(new_n540));
  INV_X1    g115(.A(G90), .ZN(new_n541));
  OAI21_X1  g116(.A(new_n540), .B1(new_n531), .B2(new_n541), .ZN(new_n542));
  NOR2_X1   g117(.A1(new_n539), .A2(new_n542), .ZN(G171));
  AOI22_X1  g118(.A1(new_n511), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n544));
  NOR2_X1   g119(.A1(new_n544), .A2(new_n538), .ZN(new_n545));
  NAND2_X1  g120(.A1(new_n518), .A2(G43), .ZN(new_n546));
  INV_X1    g121(.A(G81), .ZN(new_n547));
  OAI21_X1  g122(.A(new_n546), .B1(new_n531), .B2(new_n547), .ZN(new_n548));
  NOR2_X1   g123(.A1(new_n545), .A2(new_n548), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n549), .A2(G860), .ZN(G153));
  NAND4_X1  g125(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g126(.A1(G1), .A2(G3), .ZN(new_n552));
  XNOR2_X1  g127(.A(new_n552), .B(KEYINPUT74), .ZN(new_n553));
  XNOR2_X1  g128(.A(new_n553), .B(KEYINPUT8), .ZN(new_n554));
  NAND4_X1  g129(.A1(G319), .A2(G483), .A3(G661), .A4(new_n554), .ZN(G188));
  NAND2_X1  g130(.A1(new_n518), .A2(G53), .ZN(new_n556));
  XNOR2_X1  g131(.A(new_n556), .B(KEYINPUT9), .ZN(new_n557));
  NAND2_X1  g132(.A1(G78), .A2(G543), .ZN(new_n558));
  INV_X1    g133(.A(new_n507), .ZN(new_n559));
  NOR2_X1   g134(.A1(KEYINPUT5), .A2(G543), .ZN(new_n560));
  NOR2_X1   g135(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  INV_X1    g136(.A(G65), .ZN(new_n562));
  OAI21_X1  g137(.A(new_n558), .B1(new_n561), .B2(new_n562), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n563), .A2(G651), .ZN(new_n564));
  AND2_X1   g139(.A1(new_n511), .A2(new_n514), .ZN(new_n565));
  NAND2_X1  g140(.A1(new_n565), .A2(G91), .ZN(new_n566));
  NAND3_X1  g141(.A1(new_n557), .A2(new_n564), .A3(new_n566), .ZN(G299));
  INV_X1    g142(.A(G171), .ZN(G301));
  INV_X1    g143(.A(G168), .ZN(G286));
  OAI21_X1  g144(.A(G651), .B1(new_n511), .B2(G74), .ZN(new_n570));
  INV_X1    g145(.A(G87), .ZN(new_n571));
  INV_X1    g146(.A(G49), .ZN(new_n572));
  INV_X1    g147(.A(new_n518), .ZN(new_n573));
  OAI221_X1 g148(.A(new_n570), .B1(new_n531), .B2(new_n571), .C1(new_n572), .C2(new_n573), .ZN(G288));
  NAND2_X1  g149(.A1(G73), .A2(G543), .ZN(new_n575));
  INV_X1    g150(.A(G61), .ZN(new_n576));
  AOI21_X1  g151(.A(new_n576), .B1(new_n506), .B2(new_n507), .ZN(new_n577));
  INV_X1    g152(.A(KEYINPUT75), .ZN(new_n578));
  OAI21_X1  g153(.A(new_n575), .B1(new_n577), .B2(new_n578), .ZN(new_n579));
  OAI211_X1 g154(.A(new_n578), .B(G61), .C1(new_n559), .C2(new_n560), .ZN(new_n580));
  INV_X1    g155(.A(new_n580), .ZN(new_n581));
  OAI21_X1  g156(.A(G651), .B1(new_n579), .B2(new_n581), .ZN(new_n582));
  AOI22_X1  g157(.A1(new_n565), .A2(G86), .B1(G48), .B2(new_n518), .ZN(new_n583));
  NAND2_X1  g158(.A1(new_n582), .A2(new_n583), .ZN(G305));
  AOI22_X1  g159(.A1(new_n511), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n585));
  NOR2_X1   g160(.A1(new_n585), .A2(new_n538), .ZN(new_n586));
  NAND2_X1  g161(.A1(new_n518), .A2(G47), .ZN(new_n587));
  INV_X1    g162(.A(G85), .ZN(new_n588));
  OAI21_X1  g163(.A(new_n587), .B1(new_n531), .B2(new_n588), .ZN(new_n589));
  NOR2_X1   g164(.A1(new_n586), .A2(new_n589), .ZN(new_n590));
  INV_X1    g165(.A(new_n590), .ZN(G290));
  NAND3_X1  g166(.A1(new_n565), .A2(KEYINPUT10), .A3(G92), .ZN(new_n592));
  INV_X1    g167(.A(KEYINPUT10), .ZN(new_n593));
  INV_X1    g168(.A(G92), .ZN(new_n594));
  OAI21_X1  g169(.A(new_n593), .B1(new_n531), .B2(new_n594), .ZN(new_n595));
  NAND2_X1  g170(.A1(new_n592), .A2(new_n595), .ZN(new_n596));
  NAND2_X1  g171(.A1(G79), .A2(G543), .ZN(new_n597));
  XOR2_X1   g172(.A(KEYINPUT76), .B(G66), .Z(new_n598));
  OAI21_X1  g173(.A(new_n597), .B1(new_n598), .B2(new_n561), .ZN(new_n599));
  AOI22_X1  g174(.A1(new_n599), .A2(G651), .B1(G54), .B2(new_n518), .ZN(new_n600));
  NAND2_X1  g175(.A1(new_n596), .A2(new_n600), .ZN(new_n601));
  INV_X1    g176(.A(G868), .ZN(new_n602));
  NAND2_X1  g177(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  OAI21_X1  g178(.A(new_n603), .B1(new_n602), .B2(G171), .ZN(G284));
  OAI21_X1  g179(.A(new_n603), .B1(new_n602), .B2(G171), .ZN(G321));
  NAND2_X1  g180(.A1(G299), .A2(new_n602), .ZN(new_n606));
  OAI21_X1  g181(.A(new_n606), .B1(G168), .B2(new_n602), .ZN(G280));
  XNOR2_X1  g182(.A(G280), .B(KEYINPUT77), .ZN(G297));
  AND2_X1   g183(.A1(new_n596), .A2(new_n600), .ZN(new_n609));
  INV_X1    g184(.A(G559), .ZN(new_n610));
  OAI21_X1  g185(.A(new_n609), .B1(new_n610), .B2(G860), .ZN(G148));
  NAND2_X1  g186(.A1(new_n609), .A2(new_n610), .ZN(new_n612));
  NAND2_X1  g187(.A1(new_n612), .A2(G868), .ZN(new_n613));
  OAI21_X1  g188(.A(new_n613), .B1(G868), .B2(new_n549), .ZN(G323));
  XNOR2_X1  g189(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g190(.A1(new_n484), .A2(G123), .ZN(new_n616));
  NOR2_X1   g191(.A1(new_n467), .A2(G111), .ZN(new_n617));
  OAI21_X1  g192(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n618));
  NAND2_X1  g193(.A1(new_n473), .A2(new_n478), .ZN(new_n619));
  INV_X1    g194(.A(G135), .ZN(new_n620));
  OAI221_X1 g195(.A(new_n616), .B1(new_n617), .B2(new_n618), .C1(new_n619), .C2(new_n620), .ZN(new_n621));
  XNOR2_X1  g196(.A(new_n621), .B(KEYINPUT79), .ZN(new_n622));
  INV_X1    g197(.A(new_n622), .ZN(new_n623));
  OR2_X1    g198(.A1(new_n623), .A2(G2096), .ZN(new_n624));
  NAND2_X1  g199(.A1(new_n623), .A2(G2096), .ZN(new_n625));
  NAND3_X1  g200(.A1(new_n467), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n626));
  XNOR2_X1  g201(.A(new_n626), .B(KEYINPUT12), .ZN(new_n627));
  XNOR2_X1  g202(.A(new_n627), .B(G2100), .ZN(new_n628));
  XNOR2_X1  g203(.A(KEYINPUT78), .B(KEYINPUT13), .ZN(new_n629));
  XNOR2_X1  g204(.A(new_n628), .B(new_n629), .ZN(new_n630));
  NAND3_X1  g205(.A1(new_n624), .A2(new_n625), .A3(new_n630), .ZN(G156));
  INV_X1    g206(.A(KEYINPUT14), .ZN(new_n632));
  XNOR2_X1  g207(.A(G2427), .B(G2438), .ZN(new_n633));
  XNOR2_X1  g208(.A(new_n633), .B(G2430), .ZN(new_n634));
  XNOR2_X1  g209(.A(KEYINPUT15), .B(G2435), .ZN(new_n635));
  AOI21_X1  g210(.A(new_n632), .B1(new_n634), .B2(new_n635), .ZN(new_n636));
  OAI21_X1  g211(.A(new_n636), .B1(new_n635), .B2(new_n634), .ZN(new_n637));
  XNOR2_X1  g212(.A(G2451), .B(G2454), .ZN(new_n638));
  XNOR2_X1  g213(.A(new_n638), .B(KEYINPUT16), .ZN(new_n639));
  XNOR2_X1  g214(.A(G1341), .B(G1348), .ZN(new_n640));
  XNOR2_X1  g215(.A(new_n639), .B(new_n640), .ZN(new_n641));
  XNOR2_X1  g216(.A(new_n637), .B(new_n641), .ZN(new_n642));
  XNOR2_X1  g217(.A(G2443), .B(G2446), .ZN(new_n643));
  NAND2_X1  g218(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  NAND2_X1  g219(.A1(new_n644), .A2(G14), .ZN(new_n645));
  NOR2_X1   g220(.A1(new_n642), .A2(new_n643), .ZN(new_n646));
  NOR2_X1   g221(.A1(new_n645), .A2(new_n646), .ZN(G401));
  INV_X1    g222(.A(KEYINPUT18), .ZN(new_n648));
  XOR2_X1   g223(.A(G2084), .B(G2090), .Z(new_n649));
  XNOR2_X1  g224(.A(G2067), .B(G2678), .ZN(new_n650));
  NAND2_X1  g225(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  NAND2_X1  g226(.A1(new_n651), .A2(KEYINPUT17), .ZN(new_n652));
  NOR2_X1   g227(.A1(new_n649), .A2(new_n650), .ZN(new_n653));
  OAI21_X1  g228(.A(new_n648), .B1(new_n652), .B2(new_n653), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n654), .B(G2100), .ZN(new_n655));
  XOR2_X1   g230(.A(G2072), .B(G2078), .Z(new_n656));
  AOI21_X1  g231(.A(new_n656), .B1(new_n651), .B2(KEYINPUT18), .ZN(new_n657));
  XNOR2_X1  g232(.A(new_n657), .B(G2096), .ZN(new_n658));
  XNOR2_X1  g233(.A(new_n655), .B(new_n658), .ZN(G227));
  XNOR2_X1  g234(.A(G1981), .B(G1986), .ZN(new_n660));
  INV_X1    g235(.A(new_n660), .ZN(new_n661));
  XOR2_X1   g236(.A(G1956), .B(G2474), .Z(new_n662));
  XOR2_X1   g237(.A(G1961), .B(G1966), .Z(new_n663));
  NAND2_X1  g238(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  OR2_X1    g239(.A1(new_n664), .A2(KEYINPUT80), .ZN(new_n665));
  XOR2_X1   g240(.A(G1971), .B(G1976), .Z(new_n666));
  XNOR2_X1  g241(.A(new_n666), .B(KEYINPUT19), .ZN(new_n667));
  NAND2_X1  g242(.A1(new_n664), .A2(KEYINPUT80), .ZN(new_n668));
  NAND3_X1  g243(.A1(new_n665), .A2(new_n667), .A3(new_n668), .ZN(new_n669));
  XNOR2_X1  g244(.A(new_n669), .B(KEYINPUT81), .ZN(new_n670));
  INV_X1    g245(.A(KEYINPUT20), .ZN(new_n671));
  NAND2_X1  g246(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  OR2_X1    g247(.A1(new_n669), .A2(KEYINPUT81), .ZN(new_n673));
  NAND2_X1  g248(.A1(new_n669), .A2(KEYINPUT81), .ZN(new_n674));
  NAND3_X1  g249(.A1(new_n673), .A2(KEYINPUT20), .A3(new_n674), .ZN(new_n675));
  NOR2_X1   g250(.A1(new_n662), .A2(new_n663), .ZN(new_n676));
  NAND2_X1  g251(.A1(new_n667), .A2(new_n676), .ZN(new_n677));
  XNOR2_X1  g252(.A(new_n677), .B(KEYINPUT82), .ZN(new_n678));
  INV_X1    g253(.A(new_n664), .ZN(new_n679));
  OR3_X1    g254(.A1(new_n667), .A2(new_n679), .A3(new_n676), .ZN(new_n680));
  NAND4_X1  g255(.A1(new_n672), .A2(new_n675), .A3(new_n678), .A4(new_n680), .ZN(new_n681));
  XNOR2_X1  g256(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n682));
  XNOR2_X1  g257(.A(new_n681), .B(new_n682), .ZN(new_n683));
  XOR2_X1   g258(.A(G1991), .B(G1996), .Z(new_n684));
  INV_X1    g259(.A(new_n684), .ZN(new_n685));
  NOR2_X1   g260(.A1(new_n683), .A2(new_n685), .ZN(new_n686));
  INV_X1    g261(.A(new_n682), .ZN(new_n687));
  XNOR2_X1  g262(.A(new_n681), .B(new_n687), .ZN(new_n688));
  NOR2_X1   g263(.A1(new_n688), .A2(new_n684), .ZN(new_n689));
  OAI21_X1  g264(.A(new_n661), .B1(new_n686), .B2(new_n689), .ZN(new_n690));
  NAND2_X1  g265(.A1(new_n688), .A2(new_n684), .ZN(new_n691));
  NAND2_X1  g266(.A1(new_n683), .A2(new_n685), .ZN(new_n692));
  NAND3_X1  g267(.A1(new_n691), .A2(new_n692), .A3(new_n660), .ZN(new_n693));
  AND2_X1   g268(.A1(new_n690), .A2(new_n693), .ZN(G229));
  MUX2_X1   g269(.A(G6), .B(G305), .S(G16), .Z(new_n695));
  XNOR2_X1  g270(.A(KEYINPUT32), .B(G1981), .ZN(new_n696));
  XOR2_X1   g271(.A(new_n695), .B(new_n696), .Z(new_n697));
  INV_X1    g272(.A(G16), .ZN(new_n698));
  NAND2_X1  g273(.A1(new_n698), .A2(G22), .ZN(new_n699));
  OAI21_X1  g274(.A(new_n699), .B1(G166), .B2(new_n698), .ZN(new_n700));
  INV_X1    g275(.A(G1971), .ZN(new_n701));
  XNOR2_X1  g276(.A(new_n700), .B(new_n701), .ZN(new_n702));
  NAND2_X1  g277(.A1(new_n698), .A2(G23), .ZN(new_n703));
  INV_X1    g278(.A(G288), .ZN(new_n704));
  OAI21_X1  g279(.A(new_n703), .B1(new_n704), .B2(new_n698), .ZN(new_n705));
  XNOR2_X1  g280(.A(KEYINPUT33), .B(G1976), .ZN(new_n706));
  XNOR2_X1  g281(.A(new_n705), .B(new_n706), .ZN(new_n707));
  NAND3_X1  g282(.A1(new_n697), .A2(new_n702), .A3(new_n707), .ZN(new_n708));
  NAND2_X1  g283(.A1(new_n708), .A2(KEYINPUT34), .ZN(new_n709));
  XNOR2_X1  g284(.A(new_n709), .B(KEYINPUT83), .ZN(new_n710));
  NAND2_X1  g285(.A1(new_n479), .A2(G131), .ZN(new_n711));
  OAI21_X1  g286(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n712));
  INV_X1    g287(.A(G107), .ZN(new_n713));
  AOI21_X1  g288(.A(new_n712), .B1(new_n713), .B2(G2105), .ZN(new_n714));
  AOI21_X1  g289(.A(new_n714), .B1(new_n484), .B2(G119), .ZN(new_n715));
  NAND2_X1  g290(.A1(new_n711), .A2(new_n715), .ZN(new_n716));
  INV_X1    g291(.A(new_n716), .ZN(new_n717));
  NAND2_X1  g292(.A1(new_n717), .A2(G29), .ZN(new_n718));
  OAI21_X1  g293(.A(new_n718), .B1(G25), .B2(G29), .ZN(new_n719));
  XOR2_X1   g294(.A(KEYINPUT35), .B(G1991), .Z(new_n720));
  AND2_X1   g295(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  NOR2_X1   g296(.A1(new_n590), .A2(new_n698), .ZN(new_n722));
  AOI21_X1  g297(.A(new_n722), .B1(new_n698), .B2(G24), .ZN(new_n723));
  INV_X1    g298(.A(new_n723), .ZN(new_n724));
  AND2_X1   g299(.A1(new_n724), .A2(G1986), .ZN(new_n725));
  NOR2_X1   g300(.A1(new_n719), .A2(new_n720), .ZN(new_n726));
  NOR2_X1   g301(.A1(new_n724), .A2(G1986), .ZN(new_n727));
  NOR4_X1   g302(.A1(new_n721), .A2(new_n725), .A3(new_n726), .A4(new_n727), .ZN(new_n728));
  OAI211_X1 g303(.A(new_n710), .B(new_n728), .C1(KEYINPUT34), .C2(new_n708), .ZN(new_n729));
  XOR2_X1   g304(.A(new_n729), .B(KEYINPUT36), .Z(new_n730));
  INV_X1    g305(.A(G29), .ZN(new_n731));
  NAND2_X1  g306(.A1(new_n731), .A2(G35), .ZN(new_n732));
  XOR2_X1   g307(.A(new_n732), .B(KEYINPUT90), .Z(new_n733));
  AOI21_X1  g308(.A(new_n733), .B1(new_n486), .B2(G29), .ZN(new_n734));
  XNOR2_X1  g309(.A(new_n734), .B(KEYINPUT29), .ZN(new_n735));
  INV_X1    g310(.A(G2090), .ZN(new_n736));
  NOR2_X1   g311(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  XOR2_X1   g312(.A(new_n737), .B(KEYINPUT91), .Z(new_n738));
  XNOR2_X1  g313(.A(KEYINPUT27), .B(G1996), .ZN(new_n739));
  NAND3_X1  g314(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n740));
  XNOR2_X1  g315(.A(new_n740), .B(KEYINPUT86), .ZN(new_n741));
  XNOR2_X1  g316(.A(new_n741), .B(KEYINPUT26), .ZN(new_n742));
  NAND2_X1  g317(.A1(new_n484), .A2(G129), .ZN(new_n743));
  NAND3_X1  g318(.A1(new_n467), .A2(G105), .A3(G2104), .ZN(new_n744));
  XNOR2_X1  g319(.A(new_n744), .B(KEYINPUT85), .ZN(new_n745));
  AND3_X1   g320(.A1(new_n742), .A2(new_n743), .A3(new_n745), .ZN(new_n746));
  NAND3_X1  g321(.A1(new_n479), .A2(KEYINPUT84), .A3(G141), .ZN(new_n747));
  INV_X1    g322(.A(KEYINPUT84), .ZN(new_n748));
  INV_X1    g323(.A(G141), .ZN(new_n749));
  OAI21_X1  g324(.A(new_n748), .B1(new_n619), .B2(new_n749), .ZN(new_n750));
  NAND2_X1  g325(.A1(new_n747), .A2(new_n750), .ZN(new_n751));
  NAND3_X1  g326(.A1(new_n746), .A2(new_n751), .A3(KEYINPUT87), .ZN(new_n752));
  INV_X1    g327(.A(new_n752), .ZN(new_n753));
  AOI21_X1  g328(.A(KEYINPUT87), .B1(new_n746), .B2(new_n751), .ZN(new_n754));
  NOR2_X1   g329(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  NAND2_X1  g330(.A1(new_n755), .A2(G29), .ZN(new_n756));
  OAI21_X1  g331(.A(new_n756), .B1(G29), .B2(G32), .ZN(new_n757));
  AOI21_X1  g332(.A(new_n738), .B1(new_n739), .B2(new_n757), .ZN(new_n758));
  INV_X1    g333(.A(G34), .ZN(new_n759));
  AOI21_X1  g334(.A(G29), .B1(new_n759), .B2(KEYINPUT24), .ZN(new_n760));
  OAI21_X1  g335(.A(new_n760), .B1(KEYINPUT24), .B2(new_n759), .ZN(new_n761));
  OAI21_X1  g336(.A(new_n761), .B1(new_n471), .B2(new_n731), .ZN(new_n762));
  INV_X1    g337(.A(G2084), .ZN(new_n763));
  NOR2_X1   g338(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  NOR2_X1   g339(.A1(G171), .A2(new_n698), .ZN(new_n765));
  AOI21_X1  g340(.A(new_n765), .B1(G5), .B2(new_n698), .ZN(new_n766));
  INV_X1    g341(.A(G1961), .ZN(new_n767));
  NOR2_X1   g342(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  INV_X1    g343(.A(G1341), .ZN(new_n769));
  NAND2_X1  g344(.A1(new_n549), .A2(G16), .ZN(new_n770));
  OAI21_X1  g345(.A(new_n770), .B1(G16), .B2(G19), .ZN(new_n771));
  AOI211_X1 g346(.A(new_n764), .B(new_n768), .C1(new_n769), .C2(new_n771), .ZN(new_n772));
  INV_X1    g347(.A(G28), .ZN(new_n773));
  OR2_X1    g348(.A1(new_n773), .A2(KEYINPUT30), .ZN(new_n774));
  AOI21_X1  g349(.A(G29), .B1(new_n773), .B2(KEYINPUT30), .ZN(new_n775));
  OR2_X1    g350(.A1(KEYINPUT31), .A2(G11), .ZN(new_n776));
  NAND2_X1  g351(.A1(KEYINPUT31), .A2(G11), .ZN(new_n777));
  AOI22_X1  g352(.A1(new_n774), .A2(new_n775), .B1(new_n776), .B2(new_n777), .ZN(new_n778));
  OAI21_X1  g353(.A(new_n778), .B1(new_n771), .B2(new_n769), .ZN(new_n779));
  NOR2_X1   g354(.A1(new_n609), .A2(new_n698), .ZN(new_n780));
  AOI21_X1  g355(.A(new_n780), .B1(G4), .B2(new_n698), .ZN(new_n781));
  INV_X1    g356(.A(G1348), .ZN(new_n782));
  AOI21_X1  g357(.A(new_n779), .B1(new_n781), .B2(new_n782), .ZN(new_n783));
  NAND2_X1  g358(.A1(new_n698), .A2(G20), .ZN(new_n784));
  XNOR2_X1  g359(.A(new_n784), .B(KEYINPUT23), .ZN(new_n785));
  INV_X1    g360(.A(KEYINPUT9), .ZN(new_n786));
  XNOR2_X1  g361(.A(new_n556), .B(new_n786), .ZN(new_n787));
  NAND2_X1  g362(.A1(new_n564), .A2(new_n566), .ZN(new_n788));
  NOR2_X1   g363(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  OAI21_X1  g364(.A(new_n785), .B1(new_n789), .B2(new_n698), .ZN(new_n790));
  XOR2_X1   g365(.A(KEYINPUT92), .B(G1956), .Z(new_n791));
  XNOR2_X1  g366(.A(new_n790), .B(new_n791), .ZN(new_n792));
  NAND2_X1  g367(.A1(new_n731), .A2(G27), .ZN(new_n793));
  OAI21_X1  g368(.A(new_n793), .B1(G164), .B2(new_n731), .ZN(new_n794));
  XOR2_X1   g369(.A(KEYINPUT89), .B(G2078), .Z(new_n795));
  XNOR2_X1  g370(.A(new_n794), .B(new_n795), .ZN(new_n796));
  NAND4_X1  g371(.A1(new_n772), .A2(new_n783), .A3(new_n792), .A4(new_n796), .ZN(new_n797));
  NAND2_X1  g372(.A1(new_n731), .A2(G26), .ZN(new_n798));
  XOR2_X1   g373(.A(new_n798), .B(KEYINPUT28), .Z(new_n799));
  NAND2_X1  g374(.A1(new_n484), .A2(G128), .ZN(new_n800));
  NOR2_X1   g375(.A1(new_n467), .A2(G116), .ZN(new_n801));
  OAI21_X1  g376(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n802));
  INV_X1    g377(.A(G140), .ZN(new_n803));
  OAI221_X1 g378(.A(new_n800), .B1(new_n801), .B2(new_n802), .C1(new_n619), .C2(new_n803), .ZN(new_n804));
  AOI21_X1  g379(.A(new_n799), .B1(new_n804), .B2(G29), .ZN(new_n805));
  INV_X1    g380(.A(G2067), .ZN(new_n806));
  XNOR2_X1  g381(.A(new_n805), .B(new_n806), .ZN(new_n807));
  NAND2_X1  g382(.A1(new_n698), .A2(G21), .ZN(new_n808));
  OAI21_X1  g383(.A(new_n808), .B1(G168), .B2(new_n698), .ZN(new_n809));
  XNOR2_X1  g384(.A(new_n809), .B(G1966), .ZN(new_n810));
  OR2_X1    g385(.A1(new_n781), .A2(new_n782), .ZN(new_n811));
  NAND2_X1  g386(.A1(new_n735), .A2(new_n736), .ZN(new_n812));
  NAND2_X1  g387(.A1(new_n731), .A2(G33), .ZN(new_n813));
  NAND3_X1  g388(.A1(new_n467), .A2(G103), .A3(G2104), .ZN(new_n814));
  XOR2_X1   g389(.A(new_n814), .B(KEYINPUT25), .Z(new_n815));
  AOI22_X1  g390(.A1(new_n499), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n816));
  OAI21_X1  g391(.A(new_n815), .B1(new_n816), .B2(new_n467), .ZN(new_n817));
  AOI21_X1  g392(.A(new_n817), .B1(new_n479), .B2(G139), .ZN(new_n818));
  OAI21_X1  g393(.A(new_n813), .B1(new_n818), .B2(new_n731), .ZN(new_n819));
  XOR2_X1   g394(.A(new_n819), .B(G2072), .Z(new_n820));
  NAND2_X1  g395(.A1(new_n622), .A2(G29), .ZN(new_n821));
  NAND4_X1  g396(.A1(new_n811), .A2(new_n812), .A3(new_n820), .A4(new_n821), .ZN(new_n822));
  NOR4_X1   g397(.A1(new_n797), .A2(new_n807), .A3(new_n810), .A4(new_n822), .ZN(new_n823));
  AOI22_X1  g398(.A1(new_n766), .A2(new_n767), .B1(new_n763), .B2(new_n762), .ZN(new_n824));
  OAI21_X1  g399(.A(new_n824), .B1(new_n757), .B2(new_n739), .ZN(new_n825));
  NAND2_X1  g400(.A1(new_n825), .A2(KEYINPUT88), .ZN(new_n826));
  OR2_X1    g401(.A1(new_n825), .A2(KEYINPUT88), .ZN(new_n827));
  NAND4_X1  g402(.A1(new_n758), .A2(new_n823), .A3(new_n826), .A4(new_n827), .ZN(new_n828));
  NOR2_X1   g403(.A1(new_n730), .A2(new_n828), .ZN(G311));
  INV_X1    g404(.A(G311), .ZN(G150));
  NAND2_X1  g405(.A1(new_n609), .A2(G559), .ZN(new_n831));
  XNOR2_X1  g406(.A(new_n831), .B(KEYINPUT38), .ZN(new_n832));
  AOI22_X1  g407(.A1(new_n511), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n833));
  OR2_X1    g408(.A1(new_n833), .A2(new_n538), .ZN(new_n834));
  NAND2_X1  g409(.A1(new_n518), .A2(G55), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n565), .A2(G93), .ZN(new_n836));
  NAND4_X1  g411(.A1(new_n549), .A2(new_n834), .A3(new_n835), .A4(new_n836), .ZN(new_n837));
  INV_X1    g412(.A(G93), .ZN(new_n838));
  OAI221_X1 g413(.A(new_n835), .B1(new_n531), .B2(new_n838), .C1(new_n833), .C2(new_n538), .ZN(new_n839));
  OAI21_X1  g414(.A(new_n839), .B1(new_n545), .B2(new_n548), .ZN(new_n840));
  NAND2_X1  g415(.A1(new_n837), .A2(new_n840), .ZN(new_n841));
  XNOR2_X1  g416(.A(new_n832), .B(new_n841), .ZN(new_n842));
  INV_X1    g417(.A(KEYINPUT39), .ZN(new_n843));
  AOI21_X1  g418(.A(G860), .B1(new_n842), .B2(new_n843), .ZN(new_n844));
  OAI21_X1  g419(.A(new_n844), .B1(new_n843), .B2(new_n842), .ZN(new_n845));
  XNOR2_X1  g420(.A(new_n845), .B(KEYINPUT93), .ZN(new_n846));
  NAND2_X1  g421(.A1(new_n839), .A2(G860), .ZN(new_n847));
  XOR2_X1   g422(.A(new_n847), .B(KEYINPUT37), .Z(new_n848));
  NAND2_X1  g423(.A1(new_n846), .A2(new_n848), .ZN(G145));
  NAND2_X1  g424(.A1(G162), .A2(G160), .ZN(new_n850));
  INV_X1    g425(.A(KEYINPUT94), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n486), .A2(new_n471), .ZN(new_n852));
  NAND3_X1  g427(.A1(new_n850), .A2(new_n851), .A3(new_n852), .ZN(new_n853));
  INV_X1    g428(.A(new_n853), .ZN(new_n854));
  AOI21_X1  g429(.A(new_n851), .B1(new_n850), .B2(new_n852), .ZN(new_n855));
  OAI21_X1  g430(.A(new_n623), .B1(new_n854), .B2(new_n855), .ZN(new_n856));
  INV_X1    g431(.A(new_n855), .ZN(new_n857));
  NAND3_X1  g432(.A1(new_n857), .A2(new_n622), .A3(new_n853), .ZN(new_n858));
  NAND2_X1  g433(.A1(new_n856), .A2(new_n858), .ZN(new_n859));
  INV_X1    g434(.A(new_n859), .ZN(new_n860));
  XNOR2_X1  g435(.A(new_n804), .B(new_n503), .ZN(new_n861));
  INV_X1    g436(.A(new_n861), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n746), .A2(new_n751), .ZN(new_n863));
  NOR2_X1   g438(.A1(new_n863), .A2(new_n818), .ZN(new_n864));
  INV_X1    g439(.A(new_n864), .ZN(new_n865));
  INV_X1    g440(.A(new_n818), .ZN(new_n866));
  OAI211_X1 g441(.A(new_n862), .B(new_n865), .C1(new_n755), .C2(new_n866), .ZN(new_n867));
  INV_X1    g442(.A(KEYINPUT87), .ZN(new_n868));
  NAND2_X1  g443(.A1(new_n863), .A2(new_n868), .ZN(new_n869));
  AOI21_X1  g444(.A(new_n866), .B1(new_n869), .B2(new_n752), .ZN(new_n870));
  OAI21_X1  g445(.A(new_n861), .B1(new_n870), .B2(new_n864), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n867), .A2(new_n871), .ZN(new_n872));
  OAI21_X1  g447(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n873));
  INV_X1    g448(.A(KEYINPUT95), .ZN(new_n874));
  OR2_X1    g449(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  INV_X1    g450(.A(G118), .ZN(new_n876));
  AOI22_X1  g451(.A1(new_n873), .A2(new_n874), .B1(new_n876), .B2(G2105), .ZN(new_n877));
  AOI22_X1  g452(.A1(new_n484), .A2(G130), .B1(new_n875), .B2(new_n877), .ZN(new_n878));
  INV_X1    g453(.A(G142), .ZN(new_n879));
  OAI21_X1  g454(.A(new_n878), .B1(new_n619), .B2(new_n879), .ZN(new_n880));
  XNOR2_X1  g455(.A(new_n880), .B(new_n627), .ZN(new_n881));
  XNOR2_X1  g456(.A(new_n881), .B(new_n716), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n882), .A2(KEYINPUT97), .ZN(new_n883));
  AOI21_X1  g458(.A(new_n860), .B1(new_n872), .B2(new_n883), .ZN(new_n884));
  OR2_X1    g459(.A1(new_n872), .A2(new_n883), .ZN(new_n885));
  AOI21_X1  g460(.A(G37), .B1(new_n884), .B2(new_n885), .ZN(new_n886));
  INV_X1    g461(.A(new_n882), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n872), .A2(new_n887), .ZN(new_n888));
  NAND3_X1  g463(.A1(new_n867), .A2(new_n871), .A3(new_n882), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  AOI21_X1  g465(.A(KEYINPUT96), .B1(new_n890), .B2(new_n860), .ZN(new_n891));
  INV_X1    g466(.A(KEYINPUT96), .ZN(new_n892));
  AOI211_X1 g467(.A(new_n892), .B(new_n859), .C1(new_n888), .C2(new_n889), .ZN(new_n893));
  OAI21_X1  g468(.A(new_n886), .B1(new_n891), .B2(new_n893), .ZN(new_n894));
  XNOR2_X1  g469(.A(KEYINPUT98), .B(KEYINPUT40), .ZN(new_n895));
  XNOR2_X1  g470(.A(new_n894), .B(new_n895), .ZN(G395));
  NAND2_X1  g471(.A1(new_n839), .A2(new_n602), .ZN(new_n897));
  XOR2_X1   g472(.A(new_n841), .B(new_n612), .Z(new_n898));
  OAI21_X1  g473(.A(KEYINPUT99), .B1(new_n789), .B2(new_n601), .ZN(new_n899));
  INV_X1    g474(.A(KEYINPUT99), .ZN(new_n900));
  NAND3_X1  g475(.A1(new_n609), .A2(G299), .A3(new_n900), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n899), .A2(new_n901), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n789), .A2(new_n601), .ZN(new_n903));
  AND2_X1   g478(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  NOR2_X1   g479(.A1(new_n898), .A2(new_n904), .ZN(new_n905));
  INV_X1    g480(.A(KEYINPUT41), .ZN(new_n906));
  AND2_X1   g481(.A1(new_n899), .A2(new_n901), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n903), .A2(KEYINPUT100), .ZN(new_n908));
  INV_X1    g483(.A(KEYINPUT100), .ZN(new_n909));
  NAND3_X1  g484(.A1(new_n789), .A2(new_n909), .A3(new_n601), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n908), .A2(new_n910), .ZN(new_n911));
  OAI21_X1  g486(.A(new_n906), .B1(new_n907), .B2(new_n911), .ZN(new_n912));
  INV_X1    g487(.A(KEYINPUT101), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  NAND3_X1  g489(.A1(new_n902), .A2(new_n908), .A3(new_n910), .ZN(new_n915));
  NAND3_X1  g490(.A1(new_n915), .A2(KEYINPUT101), .A3(new_n906), .ZN(new_n916));
  NAND3_X1  g491(.A1(new_n902), .A2(KEYINPUT41), .A3(new_n903), .ZN(new_n917));
  NAND3_X1  g492(.A1(new_n914), .A2(new_n916), .A3(new_n917), .ZN(new_n918));
  AOI21_X1  g493(.A(new_n905), .B1(new_n918), .B2(new_n898), .ZN(new_n919));
  XNOR2_X1  g494(.A(G305), .B(G288), .ZN(new_n920));
  XNOR2_X1  g495(.A(new_n590), .B(G303), .ZN(new_n921));
  XNOR2_X1  g496(.A(new_n920), .B(new_n921), .ZN(new_n922));
  XOR2_X1   g497(.A(new_n922), .B(KEYINPUT42), .Z(new_n923));
  XOR2_X1   g498(.A(new_n919), .B(new_n923), .Z(new_n924));
  OAI21_X1  g499(.A(new_n897), .B1(new_n924), .B2(new_n602), .ZN(G295));
  XNOR2_X1  g500(.A(G295), .B(KEYINPUT102), .ZN(G331));
  AND3_X1   g501(.A1(new_n837), .A2(new_n840), .A3(G301), .ZN(new_n927));
  AOI21_X1  g502(.A(G301), .B1(new_n837), .B2(new_n840), .ZN(new_n928));
  OAI21_X1  g503(.A(G286), .B1(new_n927), .B2(new_n928), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n841), .A2(G171), .ZN(new_n930));
  NAND3_X1  g505(.A1(new_n837), .A2(new_n840), .A3(G301), .ZN(new_n931));
  NAND3_X1  g506(.A1(new_n930), .A2(G168), .A3(new_n931), .ZN(new_n932));
  AND2_X1   g507(.A1(new_n929), .A2(new_n932), .ZN(new_n933));
  NAND4_X1  g508(.A1(new_n914), .A2(new_n916), .A3(new_n917), .A4(new_n933), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n929), .A2(new_n932), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n935), .A2(new_n904), .ZN(new_n936));
  AND3_X1   g511(.A1(new_n934), .A2(new_n922), .A3(new_n936), .ZN(new_n937));
  AOI21_X1  g512(.A(new_n922), .B1(new_n934), .B2(new_n936), .ZN(new_n938));
  NOR3_X1   g513(.A1(new_n937), .A2(new_n938), .A3(G37), .ZN(new_n939));
  XNOR2_X1  g514(.A(KEYINPUT103), .B(KEYINPUT43), .ZN(new_n940));
  OAI21_X1  g515(.A(KEYINPUT104), .B1(new_n939), .B2(new_n940), .ZN(new_n941));
  NAND3_X1  g516(.A1(new_n929), .A2(new_n932), .A3(KEYINPUT41), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n942), .A2(new_n904), .ZN(new_n943));
  NAND4_X1  g518(.A1(new_n915), .A2(new_n929), .A3(new_n932), .A4(KEYINPUT41), .ZN(new_n944));
  AND3_X1   g519(.A1(new_n943), .A2(new_n944), .A3(new_n922), .ZN(new_n945));
  INV_X1    g520(.A(new_n940), .ZN(new_n946));
  NOR4_X1   g521(.A1(new_n938), .A2(new_n945), .A3(G37), .A4(new_n946), .ZN(new_n947));
  INV_X1    g522(.A(KEYINPUT105), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n934), .A2(new_n936), .ZN(new_n950));
  INV_X1    g525(.A(new_n922), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n950), .A2(new_n951), .ZN(new_n952));
  INV_X1    g527(.A(G37), .ZN(new_n953));
  NAND3_X1  g528(.A1(new_n934), .A2(new_n922), .A3(new_n936), .ZN(new_n954));
  NAND3_X1  g529(.A1(new_n952), .A2(new_n953), .A3(new_n954), .ZN(new_n955));
  INV_X1    g530(.A(KEYINPUT104), .ZN(new_n956));
  NAND3_X1  g531(.A1(new_n955), .A2(new_n956), .A3(new_n946), .ZN(new_n957));
  INV_X1    g532(.A(new_n945), .ZN(new_n958));
  NAND4_X1  g533(.A1(new_n952), .A2(new_n953), .A3(new_n958), .A4(new_n940), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n959), .A2(KEYINPUT105), .ZN(new_n960));
  NAND4_X1  g535(.A1(new_n941), .A2(new_n949), .A3(new_n957), .A4(new_n960), .ZN(new_n961));
  NOR2_X1   g536(.A1(new_n961), .A2(KEYINPUT44), .ZN(new_n962));
  AOI21_X1  g537(.A(G37), .B1(new_n950), .B2(new_n951), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n963), .A2(new_n958), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n964), .A2(KEYINPUT43), .ZN(new_n965));
  INV_X1    g540(.A(KEYINPUT106), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n965), .A2(new_n966), .ZN(new_n967));
  NAND3_X1  g542(.A1(new_n964), .A2(KEYINPUT106), .A3(KEYINPUT43), .ZN(new_n968));
  OAI211_X1 g543(.A(new_n967), .B(new_n968), .C1(new_n955), .C2(new_n946), .ZN(new_n969));
  AOI21_X1  g544(.A(new_n962), .B1(KEYINPUT44), .B2(new_n969), .ZN(G397));
  INV_X1    g545(.A(G1966), .ZN(new_n971));
  INV_X1    g546(.A(KEYINPUT45), .ZN(new_n972));
  NOR2_X1   g547(.A1(new_n972), .A2(G1384), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n503), .A2(new_n973), .ZN(new_n974));
  NAND3_X1  g549(.A1(new_n466), .A2(new_n470), .A3(G40), .ZN(new_n975));
  INV_X1    g550(.A(new_n975), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n974), .A2(new_n976), .ZN(new_n977));
  AOI21_X1  g552(.A(G1384), .B1(new_n496), .B2(new_n502), .ZN(new_n978));
  NOR2_X1   g553(.A1(new_n978), .A2(KEYINPUT45), .ZN(new_n979));
  OAI211_X1 g554(.A(KEYINPUT114), .B(new_n971), .C1(new_n977), .C2(new_n979), .ZN(new_n980));
  INV_X1    g555(.A(G1384), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n503), .A2(new_n981), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n982), .A2(KEYINPUT50), .ZN(new_n983));
  INV_X1    g558(.A(KEYINPUT50), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n978), .A2(new_n984), .ZN(new_n985));
  NAND4_X1  g560(.A1(new_n983), .A2(new_n763), .A3(new_n976), .A4(new_n985), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n980), .A2(new_n986), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n982), .A2(new_n972), .ZN(new_n988));
  AOI21_X1  g563(.A(new_n975), .B1(new_n503), .B2(new_n973), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n988), .A2(new_n989), .ZN(new_n990));
  AOI21_X1  g565(.A(KEYINPUT114), .B1(new_n990), .B2(new_n971), .ZN(new_n991));
  OAI211_X1 g566(.A(KEYINPUT118), .B(G8), .C1(new_n987), .C2(new_n991), .ZN(new_n992));
  NAND2_X1  g567(.A1(G286), .A2(G8), .ZN(new_n993));
  NAND2_X1  g568(.A1(new_n992), .A2(new_n993), .ZN(new_n994));
  OAI21_X1  g569(.A(new_n971), .B1(new_n977), .B2(new_n979), .ZN(new_n995));
  INV_X1    g570(.A(KEYINPUT114), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n995), .A2(new_n996), .ZN(new_n997));
  NAND3_X1  g572(.A1(new_n997), .A2(new_n986), .A3(new_n980), .ZN(new_n998));
  AOI21_X1  g573(.A(KEYINPUT118), .B1(new_n998), .B2(G8), .ZN(new_n999));
  OAI21_X1  g574(.A(KEYINPUT51), .B1(new_n994), .B2(new_n999), .ZN(new_n1000));
  INV_X1    g575(.A(KEYINPUT119), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n1000), .A2(new_n1001), .ZN(new_n1002));
  OAI211_X1 g577(.A(KEYINPUT119), .B(KEYINPUT51), .C1(new_n994), .C2(new_n999), .ZN(new_n1003));
  NOR2_X1   g578(.A1(new_n987), .A2(new_n991), .ZN(new_n1004));
  INV_X1    g579(.A(G8), .ZN(new_n1005));
  NOR2_X1   g580(.A1(new_n1004), .A2(new_n1005), .ZN(new_n1006));
  INV_X1    g581(.A(KEYINPUT51), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n993), .A2(new_n1007), .ZN(new_n1008));
  NOR2_X1   g583(.A1(new_n1006), .A2(new_n1008), .ZN(new_n1009));
  INV_X1    g584(.A(new_n1009), .ZN(new_n1010));
  NAND3_X1  g585(.A1(new_n1002), .A2(new_n1003), .A3(new_n1010), .ZN(new_n1011));
  NOR2_X1   g586(.A1(new_n1004), .A2(new_n993), .ZN(new_n1012));
  INV_X1    g587(.A(new_n1012), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n1011), .A2(new_n1013), .ZN(new_n1014));
  NAND3_X1  g589(.A1(new_n1014), .A2(KEYINPUT124), .A3(KEYINPUT62), .ZN(new_n1015));
  INV_X1    g590(.A(KEYINPUT124), .ZN(new_n1016));
  AOI21_X1  g591(.A(new_n1009), .B1(new_n1000), .B2(new_n1001), .ZN(new_n1017));
  AOI21_X1  g592(.A(new_n1012), .B1(new_n1017), .B2(new_n1003), .ZN(new_n1018));
  INV_X1    g593(.A(KEYINPUT62), .ZN(new_n1019));
  OAI21_X1  g594(.A(new_n1016), .B1(new_n1018), .B2(new_n1019), .ZN(new_n1020));
  INV_X1    g595(.A(KEYINPUT55), .ZN(new_n1021));
  NAND2_X1  g596(.A1(G303), .A2(G8), .ZN(new_n1022));
  INV_X1    g597(.A(KEYINPUT110), .ZN(new_n1023));
  AOI21_X1  g598(.A(new_n1021), .B1(new_n1022), .B2(new_n1023), .ZN(new_n1024));
  INV_X1    g599(.A(KEYINPUT111), .ZN(new_n1025));
  NAND4_X1  g600(.A1(G303), .A2(KEYINPUT110), .A3(new_n1025), .A4(G8), .ZN(new_n1026));
  NAND3_X1  g601(.A1(G303), .A2(KEYINPUT110), .A3(G8), .ZN(new_n1027));
  NAND2_X1  g602(.A1(new_n1027), .A2(KEYINPUT111), .ZN(new_n1028));
  AND3_X1   g603(.A1(new_n1024), .A2(new_n1026), .A3(new_n1028), .ZN(new_n1029));
  NAND2_X1  g604(.A1(new_n1022), .A2(new_n1023), .ZN(new_n1030));
  AOI22_X1  g605(.A1(new_n1028), .A2(new_n1026), .B1(new_n1030), .B2(KEYINPUT55), .ZN(new_n1031));
  NOR2_X1   g606(.A1(new_n1029), .A2(new_n1031), .ZN(new_n1032));
  AOI21_X1  g607(.A(new_n975), .B1(new_n982), .B2(KEYINPUT50), .ZN(new_n1033));
  NAND3_X1  g608(.A1(new_n1033), .A2(new_n736), .A3(new_n985), .ZN(new_n1034));
  OAI21_X1  g609(.A(new_n701), .B1(new_n977), .B2(new_n979), .ZN(new_n1035));
  AOI21_X1  g610(.A(new_n1005), .B1(new_n1034), .B2(new_n1035), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n1032), .A2(new_n1036), .ZN(new_n1037));
  OAI21_X1  g612(.A(KEYINPUT113), .B1(new_n1032), .B2(new_n1036), .ZN(new_n1038));
  AOI21_X1  g613(.A(new_n1005), .B1(new_n978), .B2(new_n976), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n704), .A2(G1976), .ZN(new_n1040));
  INV_X1    g615(.A(G1976), .ZN(new_n1041));
  AOI21_X1  g616(.A(KEYINPUT52), .B1(G288), .B2(new_n1041), .ZN(new_n1042));
  NAND3_X1  g617(.A1(new_n1039), .A2(new_n1040), .A3(new_n1042), .ZN(new_n1043));
  AND2_X1   g618(.A1(new_n1039), .A2(new_n1040), .ZN(new_n1044));
  INV_X1    g619(.A(KEYINPUT52), .ZN(new_n1045));
  OAI21_X1  g620(.A(new_n1043), .B1(new_n1044), .B2(new_n1045), .ZN(new_n1046));
  OAI21_X1  g621(.A(G61), .B1(new_n559), .B2(new_n560), .ZN(new_n1047));
  AOI22_X1  g622(.A1(new_n1047), .A2(KEYINPUT75), .B1(G73), .B2(G543), .ZN(new_n1048));
  AOI21_X1  g623(.A(new_n538), .B1(new_n1048), .B2(new_n580), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n518), .A2(G48), .ZN(new_n1050));
  INV_X1    g625(.A(G86), .ZN(new_n1051));
  OAI21_X1  g626(.A(new_n1050), .B1(new_n531), .B2(new_n1051), .ZN(new_n1052));
  OAI21_X1  g627(.A(G1981), .B1(new_n1049), .B2(new_n1052), .ZN(new_n1053));
  INV_X1    g628(.A(G1981), .ZN(new_n1054));
  NAND3_X1  g629(.A1(new_n582), .A2(new_n1054), .A3(new_n583), .ZN(new_n1055));
  INV_X1    g630(.A(KEYINPUT112), .ZN(new_n1056));
  NAND3_X1  g631(.A1(new_n1053), .A2(new_n1055), .A3(new_n1056), .ZN(new_n1057));
  INV_X1    g632(.A(KEYINPUT49), .ZN(new_n1058));
  NAND3_X1  g633(.A1(G305), .A2(KEYINPUT112), .A3(G1981), .ZN(new_n1059));
  NAND3_X1  g634(.A1(new_n1057), .A2(new_n1058), .A3(new_n1059), .ZN(new_n1060));
  AND2_X1   g635(.A1(new_n1060), .A2(new_n1039), .ZN(new_n1061));
  NAND2_X1  g636(.A1(new_n1057), .A2(new_n1059), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n1062), .A2(KEYINPUT49), .ZN(new_n1063));
  AOI21_X1  g638(.A(new_n1046), .B1(new_n1061), .B2(new_n1063), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n1028), .A2(new_n1026), .ZN(new_n1065));
  INV_X1    g640(.A(new_n1024), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n1065), .A2(new_n1066), .ZN(new_n1067));
  NAND3_X1  g642(.A1(new_n1024), .A2(new_n1026), .A3(new_n1028), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n1067), .A2(new_n1068), .ZN(new_n1069));
  OAI21_X1  g644(.A(new_n976), .B1(new_n978), .B2(new_n984), .ZN(new_n1070));
  AOI211_X1 g645(.A(KEYINPUT50), .B(G1384), .C1(new_n496), .C2(new_n502), .ZN(new_n1071));
  NOR3_X1   g646(.A1(new_n1070), .A2(G2090), .A3(new_n1071), .ZN(new_n1072));
  AOI21_X1  g647(.A(G1971), .B1(new_n988), .B2(new_n989), .ZN(new_n1073));
  OAI21_X1  g648(.A(G8), .B1(new_n1072), .B2(new_n1073), .ZN(new_n1074));
  INV_X1    g649(.A(KEYINPUT113), .ZN(new_n1075));
  NAND3_X1  g650(.A1(new_n1069), .A2(new_n1074), .A3(new_n1075), .ZN(new_n1076));
  AND4_X1   g651(.A1(new_n1037), .A2(new_n1038), .A3(new_n1064), .A4(new_n1076), .ZN(new_n1077));
  INV_X1    g652(.A(G2078), .ZN(new_n1078));
  OAI211_X1 g653(.A(new_n989), .B(new_n1078), .C1(KEYINPUT45), .C2(new_n978), .ZN(new_n1079));
  INV_X1    g654(.A(KEYINPUT53), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1079), .A2(new_n1080), .ZN(new_n1081));
  OAI21_X1  g656(.A(new_n767), .B1(new_n1070), .B2(new_n1071), .ZN(new_n1082));
  NAND4_X1  g657(.A1(new_n988), .A2(KEYINPUT53), .A3(new_n1078), .A4(new_n989), .ZN(new_n1083));
  INV_X1    g658(.A(KEYINPUT120), .ZN(new_n1084));
  AND3_X1   g659(.A1(new_n1082), .A2(new_n1083), .A3(new_n1084), .ZN(new_n1085));
  AOI21_X1  g660(.A(new_n1084), .B1(new_n1082), .B2(new_n1083), .ZN(new_n1086));
  OAI21_X1  g661(.A(new_n1081), .B1(new_n1085), .B2(new_n1086), .ZN(new_n1087));
  NAND3_X1  g662(.A1(new_n1077), .A2(G171), .A3(new_n1087), .ZN(new_n1088));
  AOI21_X1  g663(.A(new_n1088), .B1(new_n1018), .B2(new_n1019), .ZN(new_n1089));
  NAND3_X1  g664(.A1(new_n1015), .A2(new_n1020), .A3(new_n1089), .ZN(new_n1090));
  NAND3_X1  g665(.A1(new_n983), .A2(new_n976), .A3(new_n985), .ZN(new_n1091));
  AOI22_X1  g666(.A1(new_n767), .A2(new_n1091), .B1(new_n1079), .B2(new_n1080), .ZN(new_n1092));
  INV_X1    g667(.A(new_n973), .ZN(new_n1093));
  AOI21_X1  g668(.A(new_n1093), .B1(new_n496), .B2(new_n502), .ZN(new_n1094));
  NAND2_X1  g669(.A1(new_n1078), .A2(KEYINPUT53), .ZN(new_n1095));
  NOR3_X1   g670(.A1(new_n1094), .A2(new_n975), .A3(new_n1095), .ZN(new_n1096));
  AND2_X1   g671(.A1(new_n978), .A2(KEYINPUT107), .ZN(new_n1097));
  OAI21_X1  g672(.A(new_n972), .B1(new_n978), .B2(KEYINPUT107), .ZN(new_n1098));
  OAI21_X1  g673(.A(new_n1096), .B1(new_n1097), .B2(new_n1098), .ZN(new_n1099));
  AOI21_X1  g674(.A(KEYINPUT122), .B1(new_n1092), .B2(new_n1099), .ZN(new_n1100));
  NAND4_X1  g675(.A1(new_n1081), .A2(KEYINPUT122), .A3(new_n1082), .A4(new_n1099), .ZN(new_n1101));
  INV_X1    g676(.A(new_n1101), .ZN(new_n1102));
  OAI21_X1  g677(.A(G171), .B1(new_n1100), .B2(new_n1102), .ZN(new_n1103));
  INV_X1    g678(.A(new_n1081), .ZN(new_n1104));
  AOI21_X1  g679(.A(G1961), .B1(new_n1033), .B2(new_n985), .ZN(new_n1105));
  NOR3_X1   g680(.A1(new_n977), .A2(new_n979), .A3(new_n1095), .ZN(new_n1106));
  OAI21_X1  g681(.A(KEYINPUT120), .B1(new_n1105), .B2(new_n1106), .ZN(new_n1107));
  NAND3_X1  g682(.A1(new_n1082), .A2(new_n1083), .A3(new_n1084), .ZN(new_n1108));
  AOI21_X1  g683(.A(new_n1104), .B1(new_n1107), .B2(new_n1108), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n1109), .A2(G301), .ZN(new_n1110));
  NAND3_X1  g685(.A1(new_n1103), .A2(new_n1110), .A3(KEYINPUT54), .ZN(new_n1111));
  NAND2_X1  g686(.A1(new_n1111), .A2(new_n1077), .ZN(new_n1112));
  NAND3_X1  g687(.A1(new_n1081), .A2(new_n1082), .A3(new_n1099), .ZN(new_n1113));
  NOR2_X1   g688(.A1(new_n1113), .A2(G171), .ZN(new_n1114));
  AOI21_X1  g689(.A(new_n1114), .B1(new_n1087), .B2(G171), .ZN(new_n1115));
  OAI21_X1  g690(.A(KEYINPUT121), .B1(new_n1115), .B2(KEYINPUT54), .ZN(new_n1116));
  NAND3_X1  g691(.A1(new_n1092), .A2(G301), .A3(new_n1099), .ZN(new_n1117));
  OAI21_X1  g692(.A(new_n1117), .B1(new_n1109), .B2(G301), .ZN(new_n1118));
  INV_X1    g693(.A(KEYINPUT121), .ZN(new_n1119));
  INV_X1    g694(.A(KEYINPUT54), .ZN(new_n1120));
  NAND3_X1  g695(.A1(new_n1118), .A2(new_n1119), .A3(new_n1120), .ZN(new_n1121));
  AOI21_X1  g696(.A(new_n1112), .B1(new_n1116), .B2(new_n1121), .ZN(new_n1122));
  INV_X1    g697(.A(KEYINPUT123), .ZN(new_n1123));
  NAND3_X1  g698(.A1(new_n1014), .A2(new_n1122), .A3(new_n1123), .ZN(new_n1124));
  NAND4_X1  g699(.A1(new_n1038), .A2(new_n1064), .A3(new_n1037), .A4(new_n1076), .ZN(new_n1125));
  INV_X1    g700(.A(KEYINPUT122), .ZN(new_n1126));
  NAND2_X1  g701(.A1(new_n1113), .A2(new_n1126), .ZN(new_n1127));
  NAND2_X1  g702(.A1(new_n1127), .A2(new_n1101), .ZN(new_n1128));
  AOI21_X1  g703(.A(new_n1120), .B1(new_n1128), .B2(G171), .ZN(new_n1129));
  AOI21_X1  g704(.A(new_n1125), .B1(new_n1129), .B2(new_n1110), .ZN(new_n1130));
  NOR3_X1   g705(.A1(new_n1115), .A2(KEYINPUT121), .A3(KEYINPUT54), .ZN(new_n1131));
  AOI21_X1  g706(.A(new_n1119), .B1(new_n1118), .B2(new_n1120), .ZN(new_n1132));
  OAI21_X1  g707(.A(new_n1130), .B1(new_n1131), .B2(new_n1132), .ZN(new_n1133));
  OAI21_X1  g708(.A(KEYINPUT123), .B1(new_n1018), .B2(new_n1133), .ZN(new_n1134));
  NOR2_X1   g709(.A1(new_n1070), .A2(new_n1071), .ZN(new_n1135));
  XOR2_X1   g710(.A(KEYINPUT56), .B(G2072), .Z(new_n1136));
  OAI22_X1  g711(.A1(new_n1135), .A2(G1956), .B1(new_n990), .B2(new_n1136), .ZN(new_n1137));
  XOR2_X1   g712(.A(KEYINPUT115), .B(KEYINPUT57), .Z(new_n1138));
  XNOR2_X1  g713(.A(new_n789), .B(new_n1138), .ZN(new_n1139));
  NOR2_X1   g714(.A1(new_n1137), .A2(new_n1139), .ZN(new_n1140));
  INV_X1    g715(.A(new_n1140), .ZN(new_n1141));
  AND2_X1   g716(.A1(new_n1137), .A2(new_n1139), .ZN(new_n1142));
  XNOR2_X1  g717(.A(new_n1142), .B(KEYINPUT116), .ZN(new_n1143));
  NOR2_X1   g718(.A1(new_n982), .A2(new_n975), .ZN(new_n1144));
  NAND2_X1  g719(.A1(new_n1144), .A2(new_n806), .ZN(new_n1145));
  OAI21_X1  g720(.A(new_n1145), .B1(new_n1135), .B2(G1348), .ZN(new_n1146));
  AND2_X1   g721(.A1(new_n1146), .A2(new_n609), .ZN(new_n1147));
  OAI21_X1  g722(.A(new_n1141), .B1(new_n1143), .B2(new_n1147), .ZN(new_n1148));
  NAND2_X1  g723(.A1(new_n1148), .A2(KEYINPUT117), .ZN(new_n1149));
  INV_X1    g724(.A(KEYINPUT117), .ZN(new_n1150));
  OAI211_X1 g725(.A(new_n1150), .B(new_n1141), .C1(new_n1143), .C2(new_n1147), .ZN(new_n1151));
  INV_X1    g726(.A(KEYINPUT61), .ZN(new_n1152));
  NOR3_X1   g727(.A1(new_n1143), .A2(new_n1152), .A3(new_n1140), .ZN(new_n1153));
  NOR3_X1   g728(.A1(new_n1146), .A2(KEYINPUT60), .A3(new_n601), .ZN(new_n1154));
  NOR2_X1   g729(.A1(new_n990), .A2(G1996), .ZN(new_n1155));
  XNOR2_X1  g730(.A(KEYINPUT58), .B(G1341), .ZN(new_n1156));
  NOR2_X1   g731(.A1(new_n1144), .A2(new_n1156), .ZN(new_n1157));
  OAI21_X1  g732(.A(new_n549), .B1(new_n1155), .B2(new_n1157), .ZN(new_n1158));
  OR2_X1    g733(.A1(new_n1158), .A2(KEYINPUT59), .ZN(new_n1159));
  NAND2_X1  g734(.A1(new_n1158), .A2(KEYINPUT59), .ZN(new_n1160));
  AOI21_X1  g735(.A(new_n1154), .B1(new_n1159), .B2(new_n1160), .ZN(new_n1161));
  NOR2_X1   g736(.A1(new_n1146), .A2(new_n609), .ZN(new_n1162));
  OAI21_X1  g737(.A(KEYINPUT60), .B1(new_n1147), .B2(new_n1162), .ZN(new_n1163));
  OAI21_X1  g738(.A(new_n1152), .B1(new_n1142), .B2(new_n1140), .ZN(new_n1164));
  NAND3_X1  g739(.A1(new_n1161), .A2(new_n1163), .A3(new_n1164), .ZN(new_n1165));
  OAI211_X1 g740(.A(new_n1149), .B(new_n1151), .C1(new_n1153), .C2(new_n1165), .ZN(new_n1166));
  NAND3_X1  g741(.A1(new_n1124), .A2(new_n1134), .A3(new_n1166), .ZN(new_n1167));
  INV_X1    g742(.A(new_n1055), .ZN(new_n1168));
  NAND2_X1  g743(.A1(new_n1061), .A2(new_n1063), .ZN(new_n1169));
  NOR2_X1   g744(.A1(G288), .A2(G1976), .ZN(new_n1170));
  AOI21_X1  g745(.A(new_n1168), .B1(new_n1169), .B2(new_n1170), .ZN(new_n1171));
  INV_X1    g746(.A(new_n1039), .ZN(new_n1172));
  INV_X1    g747(.A(new_n1064), .ZN(new_n1173));
  OAI22_X1  g748(.A1(new_n1171), .A2(new_n1172), .B1(new_n1173), .B2(new_n1037), .ZN(new_n1174));
  NAND2_X1  g749(.A1(new_n1006), .A2(G168), .ZN(new_n1175));
  INV_X1    g750(.A(new_n1175), .ZN(new_n1176));
  INV_X1    g751(.A(KEYINPUT63), .ZN(new_n1177));
  AOI21_X1  g752(.A(new_n1177), .B1(new_n1069), .B2(new_n1074), .ZN(new_n1178));
  NAND4_X1  g753(.A1(new_n1176), .A2(new_n1037), .A3(new_n1064), .A4(new_n1178), .ZN(new_n1179));
  OAI21_X1  g754(.A(new_n1177), .B1(new_n1125), .B2(new_n1175), .ZN(new_n1180));
  AOI21_X1  g755(.A(new_n1174), .B1(new_n1179), .B2(new_n1180), .ZN(new_n1181));
  NAND3_X1  g756(.A1(new_n1090), .A2(new_n1167), .A3(new_n1181), .ZN(new_n1182));
  NOR3_X1   g757(.A1(new_n1097), .A2(new_n1098), .A3(new_n975), .ZN(new_n1183));
  INV_X1    g758(.A(new_n1183), .ZN(new_n1184));
  OR2_X1    g759(.A1(new_n1184), .A2(G1996), .ZN(new_n1185));
  XOR2_X1   g760(.A(new_n1185), .B(KEYINPUT108), .Z(new_n1186));
  INV_X1    g761(.A(new_n755), .ZN(new_n1187));
  NOR2_X1   g762(.A1(new_n1186), .A2(new_n1187), .ZN(new_n1188));
  XOR2_X1   g763(.A(new_n590), .B(G1986), .Z(new_n1189));
  AND2_X1   g764(.A1(new_n1183), .A2(new_n1189), .ZN(new_n1190));
  XNOR2_X1  g765(.A(new_n804), .B(G2067), .ZN(new_n1191));
  AOI21_X1  g766(.A(new_n1191), .B1(G1996), .B2(new_n863), .ZN(new_n1192));
  NOR2_X1   g767(.A1(new_n1192), .A2(new_n1184), .ZN(new_n1193));
  XNOR2_X1  g768(.A(new_n716), .B(new_n720), .ZN(new_n1194));
  XOR2_X1   g769(.A(new_n1194), .B(KEYINPUT109), .Z(new_n1195));
  NOR2_X1   g770(.A1(new_n1195), .A2(new_n1184), .ZN(new_n1196));
  NOR4_X1   g771(.A1(new_n1188), .A2(new_n1190), .A3(new_n1193), .A4(new_n1196), .ZN(new_n1197));
  NAND2_X1  g772(.A1(new_n1182), .A2(new_n1197), .ZN(new_n1198));
  NOR3_X1   g773(.A1(new_n1184), .A2(G1986), .A3(G290), .ZN(new_n1199));
  XNOR2_X1  g774(.A(new_n1199), .B(KEYINPUT48), .ZN(new_n1200));
  NOR4_X1   g775(.A1(new_n1188), .A2(new_n1193), .A3(new_n1196), .A4(new_n1200), .ZN(new_n1201));
  OAI21_X1  g776(.A(new_n1183), .B1(new_n1191), .B2(new_n863), .ZN(new_n1202));
  AND2_X1   g777(.A1(new_n1186), .A2(KEYINPUT46), .ZN(new_n1203));
  NOR2_X1   g778(.A1(new_n1186), .A2(KEYINPUT46), .ZN(new_n1204));
  OAI21_X1  g779(.A(new_n1202), .B1(new_n1203), .B2(new_n1204), .ZN(new_n1205));
  NAND2_X1  g780(.A1(new_n1205), .A2(KEYINPUT47), .ZN(new_n1206));
  INV_X1    g781(.A(KEYINPUT47), .ZN(new_n1207));
  OAI211_X1 g782(.A(new_n1207), .B(new_n1202), .C1(new_n1203), .C2(new_n1204), .ZN(new_n1208));
  AOI21_X1  g783(.A(new_n1201), .B1(new_n1206), .B2(new_n1208), .ZN(new_n1209));
  NAND2_X1  g784(.A1(new_n717), .A2(new_n720), .ZN(new_n1210));
  NOR3_X1   g785(.A1(new_n1188), .A2(new_n1193), .A3(new_n1210), .ZN(new_n1211));
  NOR2_X1   g786(.A1(new_n804), .A2(G2067), .ZN(new_n1212));
  OAI21_X1  g787(.A(new_n1183), .B1(new_n1211), .B2(new_n1212), .ZN(new_n1213));
  INV_X1    g788(.A(KEYINPUT125), .ZN(new_n1214));
  NAND2_X1  g789(.A1(new_n1213), .A2(new_n1214), .ZN(new_n1215));
  OAI211_X1 g790(.A(KEYINPUT125), .B(new_n1183), .C1(new_n1211), .C2(new_n1212), .ZN(new_n1216));
  AND3_X1   g791(.A1(new_n1209), .A2(new_n1215), .A3(new_n1216), .ZN(new_n1217));
  NAND2_X1  g792(.A1(new_n1198), .A2(new_n1217), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g793(.A1(G227), .A2(new_n459), .ZN(new_n1220));
  OAI21_X1  g794(.A(new_n1220), .B1(new_n646), .B2(new_n645), .ZN(new_n1221));
  XOR2_X1   g795(.A(new_n1221), .B(KEYINPUT126), .Z(new_n1222));
  AOI21_X1  g796(.A(new_n1222), .B1(new_n690), .B2(new_n693), .ZN(new_n1223));
  NAND2_X1  g797(.A1(new_n894), .A2(new_n1223), .ZN(new_n1224));
  NAND2_X1  g798(.A1(new_n955), .A2(new_n946), .ZN(new_n1225));
  AOI22_X1  g799(.A1(new_n1225), .A2(KEYINPUT104), .B1(new_n948), .B2(new_n947), .ZN(new_n1226));
  AOI21_X1  g800(.A(new_n940), .B1(new_n963), .B2(new_n954), .ZN(new_n1227));
  AOI22_X1  g801(.A1(new_n1227), .A2(new_n956), .B1(new_n959), .B2(KEYINPUT105), .ZN(new_n1228));
  AOI211_X1 g802(.A(KEYINPUT127), .B(new_n1224), .C1(new_n1226), .C2(new_n1228), .ZN(new_n1229));
  INV_X1    g803(.A(KEYINPUT127), .ZN(new_n1230));
  INV_X1    g804(.A(new_n1224), .ZN(new_n1231));
  AOI21_X1  g805(.A(new_n1230), .B1(new_n961), .B2(new_n1231), .ZN(new_n1232));
  NOR2_X1   g806(.A1(new_n1229), .A2(new_n1232), .ZN(G308));
  NAND2_X1  g807(.A1(new_n961), .A2(new_n1231), .ZN(new_n1234));
  NAND2_X1  g808(.A1(new_n1234), .A2(KEYINPUT127), .ZN(new_n1235));
  NAND3_X1  g809(.A1(new_n961), .A2(new_n1230), .A3(new_n1231), .ZN(new_n1236));
  NAND2_X1  g810(.A1(new_n1235), .A2(new_n1236), .ZN(G225));
endmodule


