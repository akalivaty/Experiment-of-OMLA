//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 0 0 0 0 0 1 0 0 1 1 1 1 0 0 0 1 0 0 1 1 0 1 1 1 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 0 1 0 1 0 0 0 0 0 1 1 0 0 1 1 1 1 0 1 0 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:15:14 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n615,
    new_n616, new_n617, new_n618, new_n619, new_n620, new_n622, new_n623,
    new_n624, new_n625, new_n626, new_n627, new_n629, new_n630, new_n631,
    new_n632, new_n633, new_n634, new_n635, new_n636, new_n637, new_n638,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n664, new_n665, new_n666, new_n667, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n684, new_n685,
    new_n686, new_n687, new_n688, new_n689, new_n690, new_n691, new_n692,
    new_n693, new_n694, new_n695, new_n696, new_n698, new_n699, new_n700,
    new_n701, new_n702, new_n703, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n716, new_n717, new_n718, new_n719, new_n720, new_n721, new_n723,
    new_n725, new_n726, new_n727, new_n728, new_n729, new_n730, new_n731,
    new_n732, new_n733, new_n734, new_n735, new_n736, new_n737, new_n738,
    new_n739, new_n740, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n756, new_n757, new_n758, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n811, new_n812, new_n814,
    new_n815, new_n817, new_n818, new_n819, new_n820, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n883, new_n884, new_n885, new_n887, new_n888, new_n889,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n900, new_n901, new_n902, new_n904, new_n905, new_n906,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n938,
    new_n939, new_n940, new_n941, new_n943, new_n944;
  INV_X1    g000(.A(KEYINPUT36), .ZN(new_n202));
  NAND2_X1  g001(.A1(G183gat), .A2(G190gat), .ZN(new_n203));
  INV_X1    g002(.A(new_n203), .ZN(new_n204));
  XNOR2_X1  g003(.A(KEYINPUT27), .B(G183gat), .ZN(new_n205));
  INV_X1    g004(.A(G190gat), .ZN(new_n206));
  NAND2_X1  g005(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  AOI21_X1  g006(.A(new_n204), .B1(new_n207), .B2(KEYINPUT28), .ZN(new_n208));
  OR4_X1    g007(.A1(KEYINPUT66), .A2(KEYINPUT26), .A3(G169gat), .A4(G176gat), .ZN(new_n209));
  INV_X1    g008(.A(G169gat), .ZN(new_n210));
  INV_X1    g009(.A(G176gat), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  OAI21_X1  g011(.A(KEYINPUT26), .B1(new_n212), .B2(KEYINPUT66), .ZN(new_n213));
  NAND2_X1  g012(.A1(G169gat), .A2(G176gat), .ZN(new_n214));
  NAND3_X1  g013(.A1(new_n209), .A2(new_n213), .A3(new_n214), .ZN(new_n215));
  OAI211_X1 g014(.A(new_n208), .B(new_n215), .C1(KEYINPUT28), .C2(new_n207), .ZN(new_n216));
  NAND3_X1  g015(.A1(new_n210), .A2(new_n211), .A3(KEYINPUT23), .ZN(new_n217));
  INV_X1    g016(.A(KEYINPUT23), .ZN(new_n218));
  OAI21_X1  g017(.A(new_n218), .B1(G169gat), .B2(G176gat), .ZN(new_n219));
  NAND3_X1  g018(.A1(new_n217), .A2(new_n219), .A3(new_n214), .ZN(new_n220));
  INV_X1    g019(.A(KEYINPUT64), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  NOR2_X1   g021(.A1(KEYINPUT64), .A2(KEYINPUT25), .ZN(new_n223));
  NOR2_X1   g022(.A1(new_n204), .A2(KEYINPUT24), .ZN(new_n224));
  NAND3_X1  g023(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n225));
  OAI21_X1  g024(.A(new_n225), .B1(G183gat), .B2(G190gat), .ZN(new_n226));
  OAI221_X1 g025(.A(new_n222), .B1(new_n220), .B2(new_n223), .C1(new_n224), .C2(new_n226), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n204), .A2(KEYINPUT65), .ZN(new_n228));
  INV_X1    g027(.A(KEYINPUT65), .ZN(new_n229));
  AOI21_X1  g028(.A(KEYINPUT24), .B1(new_n203), .B2(new_n229), .ZN(new_n230));
  AOI21_X1  g029(.A(new_n226), .B1(new_n228), .B2(new_n230), .ZN(new_n231));
  OAI21_X1  g030(.A(KEYINPUT25), .B1(new_n231), .B2(new_n220), .ZN(new_n232));
  NAND3_X1  g031(.A1(new_n216), .A2(new_n227), .A3(new_n232), .ZN(new_n233));
  INV_X1    g032(.A(G134gat), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n234), .A2(G127gat), .ZN(new_n235));
  INV_X1    g034(.A(G127gat), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n236), .A2(G134gat), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n235), .A2(new_n237), .ZN(new_n238));
  XNOR2_X1  g037(.A(G113gat), .B(G120gat), .ZN(new_n239));
  OAI21_X1  g038(.A(new_n238), .B1(new_n239), .B2(KEYINPUT1), .ZN(new_n240));
  INV_X1    g039(.A(G120gat), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n241), .A2(G113gat), .ZN(new_n242));
  INV_X1    g041(.A(G113gat), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n243), .A2(G120gat), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n242), .A2(new_n244), .ZN(new_n245));
  XNOR2_X1  g044(.A(G127gat), .B(G134gat), .ZN(new_n246));
  INV_X1    g045(.A(KEYINPUT1), .ZN(new_n247));
  NAND3_X1  g046(.A1(new_n245), .A2(new_n246), .A3(new_n247), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n240), .A2(new_n248), .ZN(new_n249));
  XNOR2_X1  g048(.A(new_n249), .B(KEYINPUT67), .ZN(new_n250));
  XNOR2_X1  g049(.A(new_n233), .B(new_n250), .ZN(new_n251));
  NAND2_X1  g050(.A1(G227gat), .A2(G233gat), .ZN(new_n252));
  AND2_X1   g051(.A1(new_n251), .A2(new_n252), .ZN(new_n253));
  XNOR2_X1  g052(.A(KEYINPUT69), .B(KEYINPUT34), .ZN(new_n254));
  INV_X1    g053(.A(new_n254), .ZN(new_n255));
  NOR2_X1   g054(.A1(new_n253), .A2(new_n255), .ZN(new_n256));
  INV_X1    g055(.A(KEYINPUT34), .ZN(new_n257));
  NOR2_X1   g056(.A1(new_n257), .A2(KEYINPUT69), .ZN(new_n258));
  AOI21_X1  g057(.A(new_n256), .B1(new_n253), .B2(new_n258), .ZN(new_n259));
  INV_X1    g058(.A(new_n259), .ZN(new_n260));
  OR2_X1    g059(.A1(new_n251), .A2(new_n252), .ZN(new_n261));
  INV_X1    g060(.A(KEYINPUT33), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  INV_X1    g062(.A(KEYINPUT68), .ZN(new_n264));
  NAND2_X1  g063(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  NAND3_X1  g064(.A1(new_n261), .A2(KEYINPUT68), .A3(new_n262), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n265), .A2(new_n266), .ZN(new_n267));
  NAND2_X1  g066(.A1(new_n261), .A2(KEYINPUT32), .ZN(new_n268));
  XOR2_X1   g067(.A(G71gat), .B(G99gat), .Z(new_n269));
  XNOR2_X1  g068(.A(G15gat), .B(G43gat), .ZN(new_n270));
  XNOR2_X1  g069(.A(new_n269), .B(new_n270), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n268), .A2(new_n271), .ZN(new_n272));
  INV_X1    g071(.A(new_n272), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n267), .A2(new_n273), .ZN(new_n274));
  AOI21_X1  g073(.A(new_n268), .B1(KEYINPUT33), .B2(new_n271), .ZN(new_n275));
  INV_X1    g074(.A(new_n275), .ZN(new_n276));
  AOI21_X1  g075(.A(new_n260), .B1(new_n274), .B2(new_n276), .ZN(new_n277));
  AOI21_X1  g076(.A(new_n272), .B1(new_n265), .B2(new_n266), .ZN(new_n278));
  NOR3_X1   g077(.A1(new_n278), .A2(new_n275), .A3(new_n259), .ZN(new_n279));
  OAI21_X1  g078(.A(new_n202), .B1(new_n277), .B2(new_n279), .ZN(new_n280));
  OAI21_X1  g079(.A(new_n259), .B1(new_n278), .B2(new_n275), .ZN(new_n281));
  NAND3_X1  g080(.A1(new_n274), .A2(new_n276), .A3(new_n260), .ZN(new_n282));
  NAND3_X1  g081(.A1(new_n281), .A2(new_n282), .A3(KEYINPUT36), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n280), .A2(new_n283), .ZN(new_n284));
  INV_X1    g083(.A(KEYINPUT3), .ZN(new_n285));
  XNOR2_X1  g084(.A(G197gat), .B(G204gat), .ZN(new_n286));
  INV_X1    g085(.A(G211gat), .ZN(new_n287));
  INV_X1    g086(.A(G218gat), .ZN(new_n288));
  NOR2_X1   g087(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  OAI21_X1  g088(.A(new_n286), .B1(KEYINPUT22), .B2(new_n289), .ZN(new_n290));
  XNOR2_X1  g089(.A(G211gat), .B(G218gat), .ZN(new_n291));
  XNOR2_X1  g090(.A(new_n290), .B(new_n291), .ZN(new_n292));
  OAI21_X1  g091(.A(new_n285), .B1(new_n292), .B2(KEYINPUT29), .ZN(new_n293));
  OR2_X1    g092(.A1(G141gat), .A2(G148gat), .ZN(new_n294));
  INV_X1    g093(.A(KEYINPUT2), .ZN(new_n295));
  NAND2_X1  g094(.A1(G141gat), .A2(G148gat), .ZN(new_n296));
  NAND3_X1  g095(.A1(new_n294), .A2(new_n295), .A3(new_n296), .ZN(new_n297));
  INV_X1    g096(.A(G162gat), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n298), .A2(G155gat), .ZN(new_n299));
  INV_X1    g098(.A(G155gat), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n300), .A2(G162gat), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n299), .A2(new_n301), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n297), .A2(new_n302), .ZN(new_n303));
  XNOR2_X1  g102(.A(KEYINPUT71), .B(G162gat), .ZN(new_n304));
  AOI21_X1  g103(.A(new_n295), .B1(new_n304), .B2(G155gat), .ZN(new_n305));
  NAND4_X1  g104(.A1(new_n294), .A2(new_n299), .A3(new_n301), .A4(new_n296), .ZN(new_n306));
  OAI21_X1  g105(.A(new_n303), .B1(new_n305), .B2(new_n306), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n293), .A2(new_n307), .ZN(new_n308));
  INV_X1    g107(.A(KEYINPUT73), .ZN(new_n309));
  OAI21_X1  g108(.A(new_n309), .B1(new_n307), .B2(KEYINPUT3), .ZN(new_n310));
  AND2_X1   g109(.A1(KEYINPUT71), .A2(G162gat), .ZN(new_n311));
  NOR2_X1   g110(.A1(KEYINPUT71), .A2(G162gat), .ZN(new_n312));
  OAI21_X1  g111(.A(G155gat), .B1(new_n311), .B2(new_n312), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n313), .A2(KEYINPUT2), .ZN(new_n314));
  AND4_X1   g113(.A1(new_n294), .A2(new_n299), .A3(new_n301), .A4(new_n296), .ZN(new_n315));
  AOI22_X1  g114(.A1(new_n314), .A2(new_n315), .B1(new_n297), .B2(new_n302), .ZN(new_n316));
  NAND3_X1  g115(.A1(new_n316), .A2(KEYINPUT73), .A3(new_n285), .ZN(new_n317));
  AOI21_X1  g116(.A(KEYINPUT29), .B1(new_n310), .B2(new_n317), .ZN(new_n318));
  INV_X1    g117(.A(new_n292), .ZN(new_n319));
  OAI21_X1  g118(.A(new_n308), .B1(new_n318), .B2(new_n319), .ZN(new_n320));
  INV_X1    g119(.A(G22gat), .ZN(new_n321));
  OR2_X1    g120(.A1(new_n320), .A2(new_n321), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n320), .A2(new_n321), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  NAND2_X1  g123(.A1(G228gat), .A2(G233gat), .ZN(new_n325));
  AOI21_X1  g124(.A(KEYINPUT79), .B1(new_n324), .B2(new_n325), .ZN(new_n326));
  NAND4_X1  g125(.A1(new_n322), .A2(G228gat), .A3(G233gat), .A4(new_n323), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n326), .A2(new_n327), .ZN(new_n328));
  XNOR2_X1  g127(.A(G78gat), .B(G106gat), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n328), .A2(new_n329), .ZN(new_n330));
  INV_X1    g129(.A(new_n329), .ZN(new_n331));
  NAND3_X1  g130(.A1(new_n326), .A2(new_n331), .A3(new_n327), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n330), .A2(new_n332), .ZN(new_n333));
  XNOR2_X1  g132(.A(KEYINPUT31), .B(G50gat), .ZN(new_n334));
  INV_X1    g133(.A(new_n334), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n333), .A2(new_n335), .ZN(new_n336));
  NAND3_X1  g135(.A1(new_n330), .A2(new_n334), .A3(new_n332), .ZN(new_n337));
  XNOR2_X1  g136(.A(G8gat), .B(G36gat), .ZN(new_n338));
  XNOR2_X1  g137(.A(G64gat), .B(G92gat), .ZN(new_n339));
  XOR2_X1   g138(.A(new_n338), .B(new_n339), .Z(new_n340));
  INV_X1    g139(.A(new_n340), .ZN(new_n341));
  INV_X1    g140(.A(KEYINPUT70), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n233), .A2(new_n342), .ZN(new_n343));
  NAND4_X1  g142(.A1(new_n216), .A2(new_n227), .A3(KEYINPUT70), .A4(new_n232), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  INV_X1    g144(.A(G226gat), .ZN(new_n346));
  INV_X1    g145(.A(G233gat), .ZN(new_n347));
  NOR2_X1   g146(.A1(new_n346), .A2(new_n347), .ZN(new_n348));
  NOR2_X1   g147(.A1(new_n348), .A2(KEYINPUT29), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n345), .A2(new_n349), .ZN(new_n350));
  INV_X1    g149(.A(new_n348), .ZN(new_n351));
  NOR2_X1   g150(.A1(new_n233), .A2(new_n351), .ZN(new_n352));
  INV_X1    g151(.A(new_n352), .ZN(new_n353));
  AOI21_X1  g152(.A(new_n292), .B1(new_n350), .B2(new_n353), .ZN(new_n354));
  NAND3_X1  g153(.A1(new_n343), .A2(new_n348), .A3(new_n344), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n233), .A2(new_n349), .ZN(new_n356));
  NAND3_X1  g155(.A1(new_n355), .A2(new_n292), .A3(new_n356), .ZN(new_n357));
  INV_X1    g156(.A(new_n357), .ZN(new_n358));
  OAI21_X1  g157(.A(new_n341), .B1(new_n354), .B2(new_n358), .ZN(new_n359));
  AOI21_X1  g158(.A(new_n352), .B1(new_n345), .B2(new_n349), .ZN(new_n360));
  OAI211_X1 g159(.A(new_n357), .B(new_n340), .C1(new_n360), .C2(new_n292), .ZN(new_n361));
  NAND3_X1  g160(.A1(new_n359), .A2(KEYINPUT30), .A3(new_n361), .ZN(new_n362));
  NOR2_X1   g161(.A1(new_n354), .A2(new_n358), .ZN(new_n363));
  INV_X1    g162(.A(KEYINPUT30), .ZN(new_n364));
  NAND3_X1  g163(.A1(new_n363), .A2(new_n364), .A3(new_n340), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n362), .A2(new_n365), .ZN(new_n366));
  NAND2_X1  g165(.A1(G225gat), .A2(G233gat), .ZN(new_n367));
  INV_X1    g166(.A(new_n367), .ZN(new_n368));
  NOR2_X1   g167(.A1(new_n307), .A2(new_n249), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n369), .A2(KEYINPUT4), .ZN(new_n370));
  INV_X1    g169(.A(new_n249), .ZN(new_n371));
  NOR2_X1   g170(.A1(new_n371), .A2(KEYINPUT67), .ZN(new_n372));
  INV_X1    g171(.A(KEYINPUT67), .ZN(new_n373));
  NOR2_X1   g172(.A1(new_n249), .A2(new_n373), .ZN(new_n374));
  NOR3_X1   g173(.A1(new_n372), .A2(new_n307), .A3(new_n374), .ZN(new_n375));
  OAI21_X1  g174(.A(new_n370), .B1(new_n375), .B2(KEYINPUT4), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n310), .A2(new_n317), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n307), .A2(KEYINPUT3), .ZN(new_n378));
  INV_X1    g177(.A(KEYINPUT72), .ZN(new_n379));
  AND3_X1   g178(.A1(new_n245), .A2(new_n246), .A3(new_n247), .ZN(new_n380));
  AOI22_X1  g179(.A1(new_n245), .A2(new_n247), .B1(new_n235), .B2(new_n237), .ZN(new_n381));
  OAI21_X1  g180(.A(new_n379), .B1(new_n380), .B2(new_n381), .ZN(new_n382));
  NAND3_X1  g181(.A1(new_n240), .A2(new_n248), .A3(KEYINPUT72), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n382), .A2(new_n383), .ZN(new_n384));
  NAND3_X1  g183(.A1(new_n377), .A2(new_n378), .A3(new_n384), .ZN(new_n385));
  INV_X1    g184(.A(new_n385), .ZN(new_n386));
  OAI21_X1  g185(.A(new_n368), .B1(new_n376), .B2(new_n386), .ZN(new_n387));
  AND3_X1   g186(.A1(new_n240), .A2(new_n248), .A3(KEYINPUT72), .ZN(new_n388));
  AOI21_X1  g187(.A(KEYINPUT72), .B1(new_n240), .B2(new_n248), .ZN(new_n389));
  OAI21_X1  g188(.A(new_n307), .B1(new_n388), .B2(new_n389), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n371), .A2(new_n316), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n390), .A2(new_n391), .ZN(new_n392));
  OAI211_X1 g191(.A(new_n387), .B(KEYINPUT39), .C1(new_n368), .C2(new_n392), .ZN(new_n393));
  XOR2_X1   g192(.A(G1gat), .B(G29gat), .Z(new_n394));
  XNOR2_X1  g193(.A(G57gat), .B(G85gat), .ZN(new_n395));
  XNOR2_X1  g194(.A(new_n394), .B(new_n395), .ZN(new_n396));
  XNOR2_X1  g195(.A(KEYINPUT76), .B(KEYINPUT0), .ZN(new_n397));
  XNOR2_X1  g196(.A(new_n396), .B(new_n397), .ZN(new_n398));
  OAI211_X1 g197(.A(new_n393), .B(new_n398), .C1(KEYINPUT39), .C2(new_n387), .ZN(new_n399));
  INV_X1    g198(.A(KEYINPUT40), .ZN(new_n400));
  OR2_X1    g199(.A1(new_n399), .A2(new_n400), .ZN(new_n401));
  INV_X1    g200(.A(KEYINPUT74), .ZN(new_n402));
  AOI21_X1  g201(.A(new_n367), .B1(new_n390), .B2(new_n391), .ZN(new_n403));
  INV_X1    g202(.A(KEYINPUT5), .ZN(new_n404));
  OAI21_X1  g203(.A(new_n402), .B1(new_n403), .B2(new_n404), .ZN(new_n405));
  AOI21_X1  g204(.A(new_n316), .B1(new_n382), .B2(new_n383), .ZN(new_n406));
  OAI21_X1  g205(.A(new_n368), .B1(new_n406), .B2(new_n369), .ZN(new_n407));
  NAND3_X1  g206(.A1(new_n407), .A2(KEYINPUT74), .A3(KEYINPUT5), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n405), .A2(new_n408), .ZN(new_n409));
  INV_X1    g208(.A(KEYINPUT75), .ZN(new_n410));
  NAND3_X1  g209(.A1(new_n250), .A2(KEYINPUT4), .A3(new_n316), .ZN(new_n411));
  OR2_X1    g210(.A1(new_n369), .A2(KEYINPUT4), .ZN(new_n412));
  NAND4_X1  g211(.A1(new_n385), .A2(new_n367), .A3(new_n411), .A4(new_n412), .ZN(new_n413));
  AND3_X1   g212(.A1(new_n409), .A2(new_n410), .A3(new_n413), .ZN(new_n414));
  AOI21_X1  g213(.A(new_n410), .B1(new_n409), .B2(new_n413), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n385), .A2(new_n367), .ZN(new_n416));
  OAI211_X1 g215(.A(new_n404), .B(new_n370), .C1(new_n375), .C2(KEYINPUT4), .ZN(new_n417));
  OAI22_X1  g216(.A1(new_n414), .A2(new_n415), .B1(new_n416), .B2(new_n417), .ZN(new_n418));
  INV_X1    g217(.A(new_n398), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n418), .A2(new_n419), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n399), .A2(new_n400), .ZN(new_n421));
  NAND3_X1  g220(.A1(new_n401), .A2(new_n420), .A3(new_n421), .ZN(new_n422));
  OAI211_X1 g221(.A(new_n336), .B(new_n337), .C1(new_n366), .C2(new_n422), .ZN(new_n423));
  NAND3_X1  g222(.A1(new_n418), .A2(KEYINPUT6), .A3(new_n419), .ZN(new_n424));
  INV_X1    g223(.A(KEYINPUT37), .ZN(new_n425));
  AOI21_X1  g224(.A(new_n340), .B1(new_n363), .B2(new_n425), .ZN(new_n426));
  OAI21_X1  g225(.A(new_n426), .B1(new_n425), .B2(new_n363), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n427), .A2(KEYINPUT38), .ZN(new_n428));
  INV_X1    g227(.A(KEYINPUT6), .ZN(new_n429));
  OAI21_X1  g228(.A(new_n398), .B1(new_n417), .B2(new_n416), .ZN(new_n430));
  INV_X1    g229(.A(new_n430), .ZN(new_n431));
  OAI21_X1  g230(.A(new_n431), .B1(new_n414), .B2(new_n415), .ZN(new_n432));
  NAND3_X1  g231(.A1(new_n420), .A2(new_n429), .A3(new_n432), .ZN(new_n433));
  AND2_X1   g232(.A1(new_n355), .A2(new_n356), .ZN(new_n434));
  AOI21_X1  g233(.A(new_n425), .B1(new_n434), .B2(new_n319), .ZN(new_n435));
  OR2_X1    g234(.A1(new_n360), .A2(new_n319), .ZN(new_n436));
  AOI21_X1  g235(.A(KEYINPUT38), .B1(new_n435), .B2(new_n436), .ZN(new_n437));
  AOI22_X1  g236(.A1(new_n426), .A2(new_n437), .B1(new_n363), .B2(new_n340), .ZN(new_n438));
  AND4_X1   g237(.A1(new_n424), .A2(new_n428), .A3(new_n433), .A4(new_n438), .ZN(new_n439));
  OAI21_X1  g238(.A(new_n284), .B1(new_n423), .B2(new_n439), .ZN(new_n440));
  INV_X1    g239(.A(new_n440), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n336), .A2(new_n337), .ZN(new_n442));
  NOR3_X1   g241(.A1(new_n403), .A2(new_n402), .A3(new_n404), .ZN(new_n443));
  AOI21_X1  g242(.A(KEYINPUT74), .B1(new_n407), .B2(KEYINPUT5), .ZN(new_n444));
  OAI21_X1  g243(.A(new_n413), .B1(new_n443), .B2(new_n444), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n445), .A2(KEYINPUT75), .ZN(new_n446));
  NAND3_X1  g245(.A1(new_n409), .A2(new_n410), .A3(new_n413), .ZN(new_n447));
  AOI21_X1  g246(.A(new_n430), .B1(new_n446), .B2(new_n447), .ZN(new_n448));
  OAI21_X1  g247(.A(KEYINPUT77), .B1(new_n448), .B2(KEYINPUT6), .ZN(new_n449));
  INV_X1    g248(.A(KEYINPUT77), .ZN(new_n450));
  NAND3_X1  g249(.A1(new_n432), .A2(new_n450), .A3(new_n429), .ZN(new_n451));
  NAND3_X1  g250(.A1(new_n449), .A2(new_n420), .A3(new_n451), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n452), .A2(new_n424), .ZN(new_n453));
  AOI21_X1  g252(.A(KEYINPUT78), .B1(new_n453), .B2(new_n366), .ZN(new_n454));
  INV_X1    g253(.A(KEYINPUT78), .ZN(new_n455));
  AND2_X1   g254(.A1(new_n362), .A2(new_n365), .ZN(new_n456));
  AOI211_X1 g255(.A(new_n455), .B(new_n456), .C1(new_n452), .C2(new_n424), .ZN(new_n457));
  OAI21_X1  g256(.A(new_n442), .B1(new_n454), .B2(new_n457), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n441), .A2(new_n458), .ZN(new_n459));
  INV_X1    g258(.A(KEYINPUT80), .ZN(new_n460));
  AND3_X1   g259(.A1(new_n281), .A2(new_n282), .A3(new_n366), .ZN(new_n461));
  AOI21_X1  g260(.A(KEYINPUT35), .B1(new_n433), .B2(new_n424), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  OAI21_X1  g262(.A(new_n460), .B1(new_n463), .B2(new_n442), .ZN(new_n464));
  INV_X1    g263(.A(new_n442), .ZN(new_n465));
  NAND4_X1  g264(.A1(new_n465), .A2(KEYINPUT80), .A3(new_n461), .A4(new_n462), .ZN(new_n466));
  AND2_X1   g265(.A1(new_n464), .A2(new_n466), .ZN(new_n467));
  INV_X1    g266(.A(KEYINPUT35), .ZN(new_n468));
  NOR2_X1   g267(.A1(new_n454), .A2(new_n457), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n281), .A2(new_n282), .ZN(new_n470));
  NOR2_X1   g269(.A1(new_n442), .A2(new_n470), .ZN(new_n471));
  AOI21_X1  g270(.A(new_n468), .B1(new_n469), .B2(new_n471), .ZN(new_n472));
  OAI21_X1  g271(.A(new_n459), .B1(new_n467), .B2(new_n472), .ZN(new_n473));
  INV_X1    g272(.A(KEYINPUT92), .ZN(new_n474));
  XNOR2_X1  g273(.A(G134gat), .B(G162gat), .ZN(new_n475));
  NAND2_X1  g274(.A1(G232gat), .A2(G233gat), .ZN(new_n476));
  INV_X1    g275(.A(KEYINPUT41), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  XOR2_X1   g277(.A(new_n475), .B(new_n478), .Z(new_n479));
  XNOR2_X1  g278(.A(G190gat), .B(G218gat), .ZN(new_n480));
  INV_X1    g279(.A(new_n480), .ZN(new_n481));
  OAI22_X1  g280(.A1(new_n481), .A2(KEYINPUT91), .B1(new_n477), .B2(new_n476), .ZN(new_n482));
  XNOR2_X1  g281(.A(KEYINPUT82), .B(G36gat), .ZN(new_n483));
  INV_X1    g282(.A(G29gat), .ZN(new_n484));
  NOR2_X1   g283(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  INV_X1    g284(.A(KEYINPUT84), .ZN(new_n486));
  XNOR2_X1  g285(.A(new_n485), .B(new_n486), .ZN(new_n487));
  INV_X1    g286(.A(KEYINPUT15), .ZN(new_n488));
  NAND2_X1  g287(.A1(G43gat), .A2(G50gat), .ZN(new_n489));
  XOR2_X1   g288(.A(KEYINPUT83), .B(G50gat), .Z(new_n490));
  OAI211_X1 g289(.A(new_n488), .B(new_n489), .C1(new_n490), .C2(G43gat), .ZN(new_n491));
  NOR2_X1   g290(.A1(G29gat), .A2(G36gat), .ZN(new_n492));
  XNOR2_X1  g291(.A(new_n492), .B(KEYINPUT14), .ZN(new_n493));
  OR2_X1    g292(.A1(G43gat), .A2(G50gat), .ZN(new_n494));
  AOI21_X1  g293(.A(new_n488), .B1(new_n494), .B2(new_n489), .ZN(new_n495));
  NOR2_X1   g294(.A1(new_n493), .A2(new_n495), .ZN(new_n496));
  NAND3_X1  g295(.A1(new_n487), .A2(new_n491), .A3(new_n496), .ZN(new_n497));
  OAI21_X1  g296(.A(new_n495), .B1(new_n485), .B2(new_n493), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  INV_X1    g298(.A(KEYINPUT90), .ZN(new_n500));
  NAND2_X1  g299(.A1(G99gat), .A2(G106gat), .ZN(new_n501));
  INV_X1    g300(.A(G85gat), .ZN(new_n502));
  INV_X1    g301(.A(G92gat), .ZN(new_n503));
  AOI22_X1  g302(.A1(KEYINPUT8), .A2(new_n501), .B1(new_n502), .B2(new_n503), .ZN(new_n504));
  NAND2_X1  g303(.A1(KEYINPUT89), .A2(KEYINPUT7), .ZN(new_n505));
  OAI21_X1  g304(.A(new_n505), .B1(new_n502), .B2(new_n503), .ZN(new_n506));
  NAND4_X1  g305(.A1(KEYINPUT89), .A2(KEYINPUT7), .A3(G85gat), .A4(G92gat), .ZN(new_n507));
  NAND3_X1  g306(.A1(new_n504), .A2(new_n506), .A3(new_n507), .ZN(new_n508));
  XNOR2_X1  g307(.A(G99gat), .B(G106gat), .ZN(new_n509));
  INV_X1    g308(.A(new_n509), .ZN(new_n510));
  OAI21_X1  g309(.A(new_n500), .B1(new_n508), .B2(new_n510), .ZN(new_n511));
  AND2_X1   g310(.A1(new_n506), .A2(new_n507), .ZN(new_n512));
  NAND4_X1  g311(.A1(new_n512), .A2(KEYINPUT90), .A3(new_n509), .A4(new_n504), .ZN(new_n513));
  AOI22_X1  g312(.A1(new_n511), .A2(new_n513), .B1(new_n510), .B2(new_n508), .ZN(new_n514));
  AOI21_X1  g313(.A(new_n482), .B1(new_n499), .B2(new_n514), .ZN(new_n515));
  INV_X1    g314(.A(KEYINPUT17), .ZN(new_n516));
  AND3_X1   g315(.A1(new_n497), .A2(new_n516), .A3(new_n498), .ZN(new_n517));
  AOI21_X1  g316(.A(new_n516), .B1(new_n497), .B2(new_n498), .ZN(new_n518));
  NOR2_X1   g317(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  OAI21_X1  g318(.A(new_n515), .B1(new_n519), .B2(new_n514), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n481), .A2(KEYINPUT91), .ZN(new_n521));
  INV_X1    g320(.A(new_n521), .ZN(new_n522));
  OR2_X1    g321(.A1(new_n520), .A2(new_n522), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n520), .A2(new_n522), .ZN(new_n524));
  AOI21_X1  g323(.A(new_n479), .B1(new_n523), .B2(new_n524), .ZN(new_n525));
  INV_X1    g324(.A(new_n525), .ZN(new_n526));
  NAND3_X1  g325(.A1(new_n523), .A2(new_n479), .A3(new_n524), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  INV_X1    g327(.A(new_n528), .ZN(new_n529));
  XNOR2_X1  g328(.A(G57gat), .B(G64gat), .ZN(new_n530));
  AOI21_X1  g329(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n531));
  OR2_X1    g330(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  XNOR2_X1  g331(.A(G71gat), .B(G78gat), .ZN(new_n533));
  XNOR2_X1  g332(.A(new_n532), .B(new_n533), .ZN(new_n534));
  NOR2_X1   g333(.A1(new_n534), .A2(KEYINPUT21), .ZN(new_n535));
  XNOR2_X1  g334(.A(G127gat), .B(G155gat), .ZN(new_n536));
  XOR2_X1   g335(.A(new_n535), .B(new_n536), .Z(new_n537));
  XNOR2_X1  g336(.A(G15gat), .B(G22gat), .ZN(new_n538));
  INV_X1    g337(.A(G1gat), .ZN(new_n539));
  NAND3_X1  g338(.A1(new_n538), .A2(KEYINPUT16), .A3(new_n539), .ZN(new_n540));
  OAI221_X1 g339(.A(new_n540), .B1(KEYINPUT85), .B2(G8gat), .C1(new_n539), .C2(new_n538), .ZN(new_n541));
  NAND2_X1  g340(.A1(KEYINPUT85), .A2(G8gat), .ZN(new_n542));
  XNOR2_X1  g341(.A(new_n541), .B(new_n542), .ZN(new_n543));
  AOI21_X1  g342(.A(new_n543), .B1(KEYINPUT21), .B2(new_n534), .ZN(new_n544));
  XNOR2_X1  g343(.A(new_n537), .B(new_n544), .ZN(new_n545));
  NAND2_X1  g344(.A1(G231gat), .A2(G233gat), .ZN(new_n546));
  XNOR2_X1  g345(.A(new_n546), .B(KEYINPUT88), .ZN(new_n547));
  XOR2_X1   g346(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n548));
  XNOR2_X1  g347(.A(new_n547), .B(new_n548), .ZN(new_n549));
  XNOR2_X1  g348(.A(G183gat), .B(G211gat), .ZN(new_n550));
  XNOR2_X1  g349(.A(new_n549), .B(new_n550), .ZN(new_n551));
  XNOR2_X1  g350(.A(new_n545), .B(new_n551), .ZN(new_n552));
  OAI21_X1  g351(.A(new_n474), .B1(new_n529), .B2(new_n552), .ZN(new_n553));
  INV_X1    g352(.A(new_n552), .ZN(new_n554));
  NAND3_X1  g353(.A1(new_n554), .A2(new_n528), .A3(KEYINPUT92), .ZN(new_n555));
  NAND2_X1  g354(.A1(G230gat), .A2(G233gat), .ZN(new_n556));
  XOR2_X1   g355(.A(new_n556), .B(KEYINPUT94), .Z(new_n557));
  AOI21_X1  g356(.A(new_n509), .B1(new_n508), .B2(KEYINPUT93), .ZN(new_n558));
  OAI21_X1  g357(.A(new_n558), .B1(KEYINPUT93), .B2(new_n508), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n511), .A2(new_n513), .ZN(new_n560));
  NAND3_X1  g359(.A1(new_n534), .A2(new_n559), .A3(new_n560), .ZN(new_n561));
  INV_X1    g360(.A(KEYINPUT10), .ZN(new_n562));
  OAI211_X1 g361(.A(new_n561), .B(new_n562), .C1(new_n514), .C2(new_n534), .ZN(new_n563));
  NAND3_X1  g362(.A1(new_n514), .A2(KEYINPUT10), .A3(new_n534), .ZN(new_n564));
  AOI21_X1  g363(.A(new_n557), .B1(new_n563), .B2(new_n564), .ZN(new_n565));
  INV_X1    g364(.A(new_n565), .ZN(new_n566));
  OAI21_X1  g365(.A(new_n561), .B1(new_n514), .B2(new_n534), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n567), .A2(new_n557), .ZN(new_n568));
  NAND2_X1  g367(.A1(new_n566), .A2(new_n568), .ZN(new_n569));
  XOR2_X1   g368(.A(G120gat), .B(G148gat), .Z(new_n570));
  XNOR2_X1  g369(.A(new_n570), .B(KEYINPUT95), .ZN(new_n571));
  XNOR2_X1  g370(.A(G176gat), .B(G204gat), .ZN(new_n572));
  XOR2_X1   g371(.A(new_n571), .B(new_n572), .Z(new_n573));
  NAND2_X1  g372(.A1(new_n569), .A2(new_n573), .ZN(new_n574));
  INV_X1    g373(.A(new_n573), .ZN(new_n575));
  NAND3_X1  g374(.A1(new_n566), .A2(new_n568), .A3(new_n575), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n574), .A2(new_n576), .ZN(new_n577));
  INV_X1    g376(.A(new_n577), .ZN(new_n578));
  NAND3_X1  g377(.A1(new_n553), .A2(new_n555), .A3(new_n578), .ZN(new_n579));
  INV_X1    g378(.A(new_n543), .ZN(new_n580));
  OAI21_X1  g379(.A(new_n580), .B1(new_n517), .B2(new_n518), .ZN(new_n581));
  NAND2_X1  g380(.A1(G229gat), .A2(G233gat), .ZN(new_n582));
  XOR2_X1   g381(.A(new_n582), .B(KEYINPUT86), .Z(new_n583));
  INV_X1    g382(.A(KEYINPUT87), .ZN(new_n584));
  AOI21_X1  g383(.A(new_n584), .B1(new_n499), .B2(new_n543), .ZN(new_n585));
  AND3_X1   g384(.A1(new_n499), .A2(new_n543), .A3(new_n584), .ZN(new_n586));
  OAI211_X1 g385(.A(new_n581), .B(new_n583), .C1(new_n585), .C2(new_n586), .ZN(new_n587));
  INV_X1    g386(.A(KEYINPUT18), .ZN(new_n588));
  NAND2_X1  g387(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  NAND2_X1  g388(.A1(new_n499), .A2(new_n543), .ZN(new_n590));
  NAND2_X1  g389(.A1(new_n590), .A2(KEYINPUT87), .ZN(new_n591));
  NAND3_X1  g390(.A1(new_n499), .A2(new_n543), .A3(new_n584), .ZN(new_n592));
  NAND2_X1  g391(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  NAND4_X1  g392(.A1(new_n593), .A2(KEYINPUT18), .A3(new_n583), .A4(new_n581), .ZN(new_n594));
  OAI22_X1  g393(.A1(new_n586), .A2(new_n585), .B1(new_n499), .B2(new_n543), .ZN(new_n595));
  XOR2_X1   g394(.A(new_n583), .B(KEYINPUT13), .Z(new_n596));
  NAND2_X1  g395(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  XNOR2_X1  g396(.A(G113gat), .B(G141gat), .ZN(new_n598));
  XNOR2_X1  g397(.A(G169gat), .B(G197gat), .ZN(new_n599));
  XNOR2_X1  g398(.A(new_n598), .B(new_n599), .ZN(new_n600));
  XOR2_X1   g399(.A(KEYINPUT81), .B(KEYINPUT11), .Z(new_n601));
  XNOR2_X1  g400(.A(new_n600), .B(new_n601), .ZN(new_n602));
  XNOR2_X1  g401(.A(new_n602), .B(KEYINPUT12), .ZN(new_n603));
  NAND4_X1  g402(.A1(new_n589), .A2(new_n594), .A3(new_n597), .A4(new_n603), .ZN(new_n604));
  INV_X1    g403(.A(new_n604), .ZN(new_n605));
  AOI22_X1  g404(.A1(new_n587), .A2(new_n588), .B1(new_n595), .B2(new_n596), .ZN(new_n606));
  AOI21_X1  g405(.A(new_n603), .B1(new_n606), .B2(new_n594), .ZN(new_n607));
  NOR2_X1   g406(.A1(new_n605), .A2(new_n607), .ZN(new_n608));
  NOR2_X1   g407(.A1(new_n579), .A2(new_n608), .ZN(new_n609));
  AND2_X1   g408(.A1(new_n473), .A2(new_n609), .ZN(new_n610));
  XNOR2_X1  g409(.A(new_n453), .B(KEYINPUT96), .ZN(new_n611));
  INV_X1    g410(.A(new_n611), .ZN(new_n612));
  NAND2_X1  g411(.A1(new_n610), .A2(new_n612), .ZN(new_n613));
  XNOR2_X1  g412(.A(new_n613), .B(G1gat), .ZN(G1324gat));
  NAND2_X1  g413(.A1(new_n610), .A2(new_n456), .ZN(new_n615));
  XNOR2_X1  g414(.A(KEYINPUT16), .B(G8gat), .ZN(new_n616));
  NOR2_X1   g415(.A1(new_n615), .A2(new_n616), .ZN(new_n617));
  XOR2_X1   g416(.A(new_n617), .B(KEYINPUT42), .Z(new_n618));
  NAND2_X1  g417(.A1(new_n615), .A2(G8gat), .ZN(new_n619));
  XNOR2_X1  g418(.A(new_n619), .B(KEYINPUT97), .ZN(new_n620));
  NAND2_X1  g419(.A1(new_n618), .A2(new_n620), .ZN(G1325gat));
  INV_X1    g420(.A(G15gat), .ZN(new_n622));
  INV_X1    g421(.A(new_n470), .ZN(new_n623));
  NAND3_X1  g422(.A1(new_n610), .A2(new_n622), .A3(new_n623), .ZN(new_n624));
  INV_X1    g423(.A(new_n284), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n610), .A2(new_n625), .ZN(new_n626));
  INV_X1    g425(.A(new_n626), .ZN(new_n627));
  OAI21_X1  g426(.A(new_n624), .B1(new_n627), .B2(new_n622), .ZN(G1326gat));
  INV_X1    g427(.A(KEYINPUT99), .ZN(new_n629));
  NAND3_X1  g428(.A1(new_n473), .A2(new_n442), .A3(new_n609), .ZN(new_n630));
  OR2_X1    g429(.A1(new_n630), .A2(KEYINPUT98), .ZN(new_n631));
  NAND2_X1  g430(.A1(new_n630), .A2(KEYINPUT98), .ZN(new_n632));
  AOI21_X1  g431(.A(new_n629), .B1(new_n631), .B2(new_n632), .ZN(new_n633));
  INV_X1    g432(.A(new_n633), .ZN(new_n634));
  XNOR2_X1  g433(.A(KEYINPUT43), .B(G22gat), .ZN(new_n635));
  NAND3_X1  g434(.A1(new_n631), .A2(new_n629), .A3(new_n632), .ZN(new_n636));
  AND3_X1   g435(.A1(new_n634), .A2(new_n635), .A3(new_n636), .ZN(new_n637));
  AOI21_X1  g436(.A(new_n635), .B1(new_n634), .B2(new_n636), .ZN(new_n638));
  NOR2_X1   g437(.A1(new_n637), .A2(new_n638), .ZN(G1327gat));
  OR2_X1    g438(.A1(new_n467), .A2(new_n472), .ZN(new_n640));
  INV_X1    g439(.A(KEYINPUT101), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n458), .A2(KEYINPUT100), .ZN(new_n642));
  INV_X1    g441(.A(KEYINPUT100), .ZN(new_n643));
  OAI211_X1 g442(.A(new_n643), .B(new_n442), .C1(new_n454), .C2(new_n457), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n642), .A2(new_n644), .ZN(new_n645));
  AOI21_X1  g444(.A(new_n641), .B1(new_n645), .B2(new_n441), .ZN(new_n646));
  AOI211_X1 g445(.A(KEYINPUT101), .B(new_n440), .C1(new_n642), .C2(new_n644), .ZN(new_n647));
  OAI21_X1  g446(.A(new_n640), .B1(new_n646), .B2(new_n647), .ZN(new_n648));
  NOR2_X1   g447(.A1(new_n528), .A2(KEYINPUT44), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n473), .A2(new_n529), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n651), .A2(KEYINPUT44), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n650), .A2(new_n652), .ZN(new_n653));
  NOR3_X1   g452(.A1(new_n554), .A2(new_n608), .A3(new_n577), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  OAI21_X1  g454(.A(G29gat), .B1(new_n655), .B2(new_n611), .ZN(new_n656));
  INV_X1    g455(.A(KEYINPUT45), .ZN(new_n657));
  INV_X1    g456(.A(new_n651), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n658), .A2(new_n654), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n612), .A2(new_n484), .ZN(new_n660));
  OAI21_X1  g459(.A(new_n657), .B1(new_n659), .B2(new_n660), .ZN(new_n661));
  OR3_X1    g460(.A1(new_n659), .A2(new_n657), .A3(new_n660), .ZN(new_n662));
  NAND3_X1  g461(.A1(new_n656), .A2(new_n661), .A3(new_n662), .ZN(G1328gat));
  NAND2_X1  g462(.A1(new_n456), .A2(new_n483), .ZN(new_n664));
  OAI21_X1  g463(.A(KEYINPUT46), .B1(new_n659), .B2(new_n664), .ZN(new_n665));
  OR3_X1    g464(.A1(new_n659), .A2(KEYINPUT46), .A3(new_n664), .ZN(new_n666));
  NOR2_X1   g465(.A1(new_n655), .A2(new_n366), .ZN(new_n667));
  OAI211_X1 g466(.A(new_n665), .B(new_n666), .C1(new_n667), .C2(new_n483), .ZN(G1329gat));
  NAND4_X1  g467(.A1(new_n653), .A2(G43gat), .A3(new_n625), .A4(new_n654), .ZN(new_n669));
  OR2_X1    g468(.A1(KEYINPUT102), .A2(KEYINPUT47), .ZN(new_n670));
  NAND3_X1  g469(.A1(new_n658), .A2(new_n623), .A3(new_n654), .ZN(new_n671));
  INV_X1    g470(.A(G43gat), .ZN(new_n672));
  AOI22_X1  g471(.A1(new_n671), .A2(new_n672), .B1(KEYINPUT102), .B2(KEYINPUT47), .ZN(new_n673));
  AND3_X1   g472(.A1(new_n669), .A2(new_n670), .A3(new_n673), .ZN(new_n674));
  AOI21_X1  g473(.A(new_n670), .B1(new_n669), .B2(new_n673), .ZN(new_n675));
  NOR2_X1   g474(.A1(new_n674), .A2(new_n675), .ZN(G1330gat));
  NAND4_X1  g475(.A1(new_n653), .A2(new_n442), .A3(new_n490), .A4(new_n654), .ZN(new_n677));
  INV_X1    g476(.A(new_n490), .ZN(new_n678));
  OAI21_X1  g477(.A(new_n678), .B1(new_n659), .B2(new_n465), .ZN(new_n679));
  XNOR2_X1  g478(.A(KEYINPUT103), .B(KEYINPUT48), .ZN(new_n680));
  AND3_X1   g479(.A1(new_n677), .A2(new_n679), .A3(new_n680), .ZN(new_n681));
  AOI21_X1  g480(.A(new_n680), .B1(new_n677), .B2(new_n679), .ZN(new_n682));
  NOR2_X1   g481(.A1(new_n681), .A2(new_n682), .ZN(G1331gat));
  INV_X1    g482(.A(new_n555), .ZN(new_n684));
  AOI21_X1  g483(.A(KEYINPUT92), .B1(new_n554), .B2(new_n528), .ZN(new_n685));
  NOR2_X1   g484(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  NAND3_X1  g485(.A1(new_n686), .A2(new_n608), .A3(new_n577), .ZN(new_n687));
  AOI21_X1  g486(.A(new_n440), .B1(new_n642), .B2(new_n644), .ZN(new_n688));
  XNOR2_X1  g487(.A(new_n688), .B(new_n641), .ZN(new_n689));
  AOI21_X1  g488(.A(new_n687), .B1(new_n689), .B2(new_n640), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n612), .A2(KEYINPUT104), .ZN(new_n691));
  INV_X1    g490(.A(KEYINPUT104), .ZN(new_n692));
  NAND2_X1  g491(.A1(new_n611), .A2(new_n692), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n691), .A2(new_n693), .ZN(new_n694));
  INV_X1    g493(.A(new_n694), .ZN(new_n695));
  NAND2_X1  g494(.A1(new_n690), .A2(new_n695), .ZN(new_n696));
  XNOR2_X1  g495(.A(new_n696), .B(G57gat), .ZN(G1332gat));
  INV_X1    g496(.A(new_n687), .ZN(new_n698));
  NAND2_X1  g497(.A1(new_n648), .A2(new_n698), .ZN(new_n699));
  NOR2_X1   g498(.A1(new_n699), .A2(new_n366), .ZN(new_n700));
  NOR2_X1   g499(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n701));
  AND2_X1   g500(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n702));
  OAI21_X1  g501(.A(new_n700), .B1(new_n701), .B2(new_n702), .ZN(new_n703));
  OAI21_X1  g502(.A(new_n703), .B1(new_n700), .B2(new_n701), .ZN(G1333gat));
  XNOR2_X1  g503(.A(KEYINPUT106), .B(KEYINPUT50), .ZN(new_n705));
  INV_X1    g504(.A(new_n705), .ZN(new_n706));
  INV_X1    g505(.A(G71gat), .ZN(new_n707));
  XNOR2_X1  g506(.A(new_n470), .B(KEYINPUT105), .ZN(new_n708));
  INV_X1    g507(.A(new_n708), .ZN(new_n709));
  OAI21_X1  g508(.A(new_n707), .B1(new_n699), .B2(new_n709), .ZN(new_n710));
  INV_X1    g509(.A(KEYINPUT107), .ZN(new_n711));
  NOR2_X1   g510(.A1(new_n284), .A2(new_n707), .ZN(new_n712));
  NAND3_X1  g511(.A1(new_n648), .A2(new_n698), .A3(new_n712), .ZN(new_n713));
  AND3_X1   g512(.A1(new_n710), .A2(new_n711), .A3(new_n713), .ZN(new_n714));
  AOI21_X1  g513(.A(new_n711), .B1(new_n710), .B2(new_n713), .ZN(new_n715));
  OAI21_X1  g514(.A(new_n706), .B1(new_n714), .B2(new_n715), .ZN(new_n716));
  AOI21_X1  g515(.A(G71gat), .B1(new_n690), .B2(new_n708), .ZN(new_n717));
  INV_X1    g516(.A(new_n713), .ZN(new_n718));
  OAI21_X1  g517(.A(KEYINPUT107), .B1(new_n717), .B2(new_n718), .ZN(new_n719));
  NAND3_X1  g518(.A1(new_n710), .A2(new_n711), .A3(new_n713), .ZN(new_n720));
  NAND3_X1  g519(.A1(new_n719), .A2(new_n720), .A3(new_n705), .ZN(new_n721));
  NAND2_X1  g520(.A1(new_n716), .A2(new_n721), .ZN(G1334gat));
  NAND2_X1  g521(.A1(new_n690), .A2(new_n442), .ZN(new_n723));
  XNOR2_X1  g522(.A(new_n723), .B(G78gat), .ZN(G1335gat));
  NAND2_X1  g523(.A1(new_n606), .A2(new_n594), .ZN(new_n725));
  INV_X1    g524(.A(new_n603), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n727), .A2(new_n604), .ZN(new_n728));
  NOR3_X1   g527(.A1(new_n728), .A2(new_n554), .A3(new_n528), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n648), .A2(new_n729), .ZN(new_n730));
  INV_X1    g529(.A(KEYINPUT51), .ZN(new_n731));
  NOR2_X1   g530(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  AOI21_X1  g531(.A(KEYINPUT51), .B1(new_n648), .B2(new_n729), .ZN(new_n733));
  OR2_X1    g532(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  NAND4_X1  g533(.A1(new_n734), .A2(new_n502), .A3(new_n577), .A4(new_n612), .ZN(new_n735));
  NOR2_X1   g534(.A1(new_n728), .A2(new_n554), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n736), .A2(new_n577), .ZN(new_n737));
  AOI21_X1  g536(.A(new_n737), .B1(new_n650), .B2(new_n652), .ZN(new_n738));
  INV_X1    g537(.A(new_n738), .ZN(new_n739));
  OAI21_X1  g538(.A(G85gat), .B1(new_n739), .B2(new_n611), .ZN(new_n740));
  NAND2_X1  g539(.A1(new_n735), .A2(new_n740), .ZN(G1336gat));
  INV_X1    g540(.A(KEYINPUT109), .ZN(new_n742));
  AOI21_X1  g541(.A(KEYINPUT51), .B1(new_n730), .B2(new_n742), .ZN(new_n743));
  AOI211_X1 g542(.A(KEYINPUT109), .B(new_n731), .C1(new_n648), .C2(new_n729), .ZN(new_n744));
  NOR3_X1   g543(.A1(new_n366), .A2(new_n578), .A3(G92gat), .ZN(new_n745));
  XOR2_X1   g544(.A(new_n745), .B(KEYINPUT108), .Z(new_n746));
  NOR3_X1   g545(.A1(new_n743), .A2(new_n744), .A3(new_n746), .ZN(new_n747));
  AOI21_X1  g546(.A(new_n503), .B1(new_n738), .B2(new_n456), .ZN(new_n748));
  OAI21_X1  g547(.A(KEYINPUT52), .B1(new_n747), .B2(new_n748), .ZN(new_n749));
  OAI21_X1  g548(.A(new_n745), .B1(new_n732), .B2(new_n733), .ZN(new_n750));
  INV_X1    g549(.A(KEYINPUT52), .ZN(new_n751));
  AOI22_X1  g550(.A1(new_n648), .A2(new_n649), .B1(new_n651), .B2(KEYINPUT44), .ZN(new_n752));
  NOR3_X1   g551(.A1(new_n752), .A2(new_n366), .A3(new_n737), .ZN(new_n753));
  OAI211_X1 g552(.A(new_n750), .B(new_n751), .C1(new_n753), .C2(new_n503), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n749), .A2(new_n754), .ZN(G1337gat));
  NOR3_X1   g554(.A1(new_n470), .A2(G99gat), .A3(new_n578), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n734), .A2(new_n756), .ZN(new_n757));
  OAI21_X1  g556(.A(G99gat), .B1(new_n739), .B2(new_n284), .ZN(new_n758));
  NAND2_X1  g557(.A1(new_n757), .A2(new_n758), .ZN(G1338gat));
  NOR3_X1   g558(.A1(new_n465), .A2(G106gat), .A3(new_n578), .ZN(new_n760));
  INV_X1    g559(.A(new_n760), .ZN(new_n761));
  NOR3_X1   g560(.A1(new_n743), .A2(new_n744), .A3(new_n761), .ZN(new_n762));
  INV_X1    g561(.A(G106gat), .ZN(new_n763));
  AOI21_X1  g562(.A(new_n763), .B1(new_n738), .B2(new_n442), .ZN(new_n764));
  OAI21_X1  g563(.A(KEYINPUT53), .B1(new_n762), .B2(new_n764), .ZN(new_n765));
  OAI21_X1  g564(.A(new_n760), .B1(new_n732), .B2(new_n733), .ZN(new_n766));
  INV_X1    g565(.A(KEYINPUT53), .ZN(new_n767));
  NOR3_X1   g566(.A1(new_n752), .A2(new_n465), .A3(new_n737), .ZN(new_n768));
  OAI211_X1 g567(.A(new_n766), .B(new_n767), .C1(new_n768), .C2(new_n763), .ZN(new_n769));
  NAND2_X1  g568(.A1(new_n765), .A2(new_n769), .ZN(G1339gat));
  INV_X1    g569(.A(KEYINPUT110), .ZN(new_n771));
  OAI21_X1  g570(.A(new_n771), .B1(new_n579), .B2(new_n728), .ZN(new_n772));
  NAND4_X1  g571(.A1(new_n686), .A2(KEYINPUT110), .A3(new_n608), .A4(new_n578), .ZN(new_n773));
  NAND2_X1  g572(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  NAND3_X1  g573(.A1(new_n563), .A2(new_n557), .A3(new_n564), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n775), .A2(KEYINPUT111), .ZN(new_n776));
  INV_X1    g575(.A(KEYINPUT111), .ZN(new_n777));
  NAND4_X1  g576(.A1(new_n563), .A2(new_n777), .A3(new_n557), .A4(new_n564), .ZN(new_n778));
  NAND4_X1  g577(.A1(new_n776), .A2(new_n566), .A3(KEYINPUT54), .A4(new_n778), .ZN(new_n779));
  INV_X1    g578(.A(KEYINPUT54), .ZN(new_n780));
  AOI21_X1  g579(.A(new_n575), .B1(new_n565), .B2(new_n780), .ZN(new_n781));
  NAND3_X1  g580(.A1(new_n779), .A2(KEYINPUT55), .A3(new_n781), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n782), .A2(new_n576), .ZN(new_n783));
  AOI21_X1  g582(.A(KEYINPUT55), .B1(new_n779), .B2(new_n781), .ZN(new_n784));
  NOR2_X1   g583(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  NOR2_X1   g584(.A1(new_n595), .A2(new_n596), .ZN(new_n786));
  AOI21_X1  g585(.A(new_n583), .B1(new_n593), .B2(new_n581), .ZN(new_n787));
  OAI21_X1  g586(.A(new_n602), .B1(new_n786), .B2(new_n787), .ZN(new_n788));
  AND2_X1   g587(.A1(new_n604), .A2(new_n788), .ZN(new_n789));
  AND4_X1   g588(.A1(new_n527), .A2(new_n785), .A3(new_n526), .A4(new_n789), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n789), .A2(new_n577), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n779), .A2(new_n781), .ZN(new_n792));
  INV_X1    g591(.A(KEYINPUT55), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n792), .A2(new_n793), .ZN(new_n794));
  NAND3_X1  g593(.A1(new_n794), .A2(new_n576), .A3(new_n782), .ZN(new_n795));
  OAI21_X1  g594(.A(new_n791), .B1(new_n608), .B2(new_n795), .ZN(new_n796));
  AOI21_X1  g595(.A(new_n790), .B1(new_n528), .B2(new_n796), .ZN(new_n797));
  OR2_X1    g596(.A1(new_n797), .A2(new_n554), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n774), .A2(new_n798), .ZN(new_n799));
  NAND4_X1  g598(.A1(new_n799), .A2(new_n465), .A3(new_n461), .A4(new_n612), .ZN(new_n800));
  NOR3_X1   g599(.A1(new_n800), .A2(new_n243), .A3(new_n608), .ZN(new_n801));
  NOR2_X1   g600(.A1(new_n797), .A2(new_n554), .ZN(new_n802));
  AOI21_X1  g601(.A(new_n802), .B1(new_n772), .B2(new_n773), .ZN(new_n803));
  NOR2_X1   g602(.A1(new_n803), .A2(new_n694), .ZN(new_n804));
  AOI21_X1  g603(.A(KEYINPUT112), .B1(new_n804), .B2(new_n471), .ZN(new_n805));
  NOR2_X1   g604(.A1(new_n805), .A2(new_n456), .ZN(new_n806));
  NAND3_X1  g605(.A1(new_n804), .A2(KEYINPUT112), .A3(new_n471), .ZN(new_n807));
  AND2_X1   g606(.A1(new_n806), .A2(new_n807), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n808), .A2(new_n728), .ZN(new_n809));
  AOI21_X1  g608(.A(new_n801), .B1(new_n809), .B2(new_n243), .ZN(G1340gat));
  NOR3_X1   g609(.A1(new_n800), .A2(new_n241), .A3(new_n578), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n808), .A2(new_n577), .ZN(new_n812));
  AOI21_X1  g611(.A(new_n811), .B1(new_n812), .B2(new_n241), .ZN(G1341gat));
  NAND3_X1  g612(.A1(new_n808), .A2(new_n236), .A3(new_n554), .ZN(new_n814));
  OAI21_X1  g613(.A(G127gat), .B1(new_n800), .B2(new_n552), .ZN(new_n815));
  NAND2_X1  g614(.A1(new_n814), .A2(new_n815), .ZN(G1342gat));
  NAND4_X1  g615(.A1(new_n806), .A2(new_n234), .A3(new_n529), .A4(new_n807), .ZN(new_n817));
  OR2_X1    g616(.A1(new_n817), .A2(KEYINPUT56), .ZN(new_n818));
  OAI21_X1  g617(.A(G134gat), .B1(new_n800), .B2(new_n528), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n817), .A2(KEYINPUT56), .ZN(new_n820));
  NAND3_X1  g619(.A1(new_n818), .A2(new_n819), .A3(new_n820), .ZN(G1343gat));
  INV_X1    g620(.A(KEYINPUT116), .ZN(new_n822));
  NOR2_X1   g621(.A1(new_n625), .A2(new_n456), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n823), .A2(new_n612), .ZN(new_n824));
  INV_X1    g623(.A(new_n824), .ZN(new_n825));
  INV_X1    g624(.A(KEYINPUT57), .ZN(new_n826));
  NOR2_X1   g625(.A1(new_n465), .A2(new_n826), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n796), .A2(KEYINPUT113), .ZN(new_n828));
  INV_X1    g627(.A(KEYINPUT113), .ZN(new_n829));
  OAI211_X1 g628(.A(new_n791), .B(new_n829), .C1(new_n608), .C2(new_n795), .ZN(new_n830));
  NAND3_X1  g629(.A1(new_n828), .A2(new_n528), .A3(new_n830), .ZN(new_n831));
  INV_X1    g630(.A(KEYINPUT114), .ZN(new_n832));
  AOI21_X1  g631(.A(new_n790), .B1(new_n831), .B2(new_n832), .ZN(new_n833));
  NAND4_X1  g632(.A1(new_n828), .A2(KEYINPUT114), .A3(new_n528), .A4(new_n830), .ZN(new_n834));
  AOI21_X1  g633(.A(new_n554), .B1(new_n833), .B2(new_n834), .ZN(new_n835));
  INV_X1    g634(.A(new_n774), .ZN(new_n836));
  OAI211_X1 g635(.A(KEYINPUT115), .B(new_n827), .C1(new_n835), .C2(new_n836), .ZN(new_n837));
  OAI21_X1  g636(.A(new_n826), .B1(new_n803), .B2(new_n465), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n837), .A2(new_n838), .ZN(new_n839));
  AOI22_X1  g638(.A1(new_n785), .A2(new_n728), .B1(new_n577), .B2(new_n789), .ZN(new_n840));
  OAI21_X1  g639(.A(new_n528), .B1(new_n840), .B2(new_n829), .ZN(new_n841));
  INV_X1    g640(.A(new_n830), .ZN(new_n842));
  OAI21_X1  g641(.A(new_n832), .B1(new_n841), .B2(new_n842), .ZN(new_n843));
  INV_X1    g642(.A(new_n790), .ZN(new_n844));
  NAND3_X1  g643(.A1(new_n843), .A2(new_n844), .A3(new_n834), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n845), .A2(new_n552), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n846), .A2(new_n774), .ZN(new_n847));
  AOI21_X1  g646(.A(KEYINPUT115), .B1(new_n847), .B2(new_n827), .ZN(new_n848));
  OAI211_X1 g647(.A(new_n728), .B(new_n825), .C1(new_n839), .C2(new_n848), .ZN(new_n849));
  AOI21_X1  g648(.A(new_n822), .B1(new_n849), .B2(G141gat), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n284), .A2(new_n442), .ZN(new_n851));
  NOR2_X1   g650(.A1(new_n851), .A2(new_n456), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n804), .A2(new_n852), .ZN(new_n853));
  NOR3_X1   g652(.A1(new_n853), .A2(G141gat), .A3(new_n608), .ZN(new_n854));
  AOI21_X1  g653(.A(new_n854), .B1(new_n849), .B2(G141gat), .ZN(new_n855));
  NOR3_X1   g654(.A1(new_n850), .A2(new_n855), .A3(KEYINPUT58), .ZN(new_n856));
  INV_X1    g655(.A(KEYINPUT58), .ZN(new_n857));
  AOI221_X4 g656(.A(new_n854), .B1(new_n822), .B2(new_n857), .C1(new_n849), .C2(G141gat), .ZN(new_n858));
  NOR2_X1   g657(.A1(new_n856), .A2(new_n858), .ZN(G1344gat));
  NOR3_X1   g658(.A1(new_n853), .A2(G148gat), .A3(new_n578), .ZN(new_n860));
  XNOR2_X1  g659(.A(new_n860), .B(KEYINPUT117), .ZN(new_n861));
  INV_X1    g660(.A(G148gat), .ZN(new_n862));
  NOR2_X1   g661(.A1(new_n862), .A2(KEYINPUT59), .ZN(new_n863));
  OAI21_X1  g662(.A(new_n825), .B1(new_n839), .B2(new_n848), .ZN(new_n864));
  OAI21_X1  g663(.A(new_n863), .B1(new_n864), .B2(new_n578), .ZN(new_n865));
  INV_X1    g664(.A(KEYINPUT118), .ZN(new_n866));
  NAND2_X1  g665(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  NAND3_X1  g666(.A1(new_n799), .A2(KEYINPUT57), .A3(new_n442), .ZN(new_n868));
  INV_X1    g667(.A(new_n831), .ZN(new_n869));
  OAI21_X1  g668(.A(new_n552), .B1(new_n869), .B2(new_n790), .ZN(new_n870));
  NAND3_X1  g669(.A1(new_n686), .A2(new_n608), .A3(new_n578), .ZN(new_n871));
  AOI21_X1  g670(.A(new_n465), .B1(new_n870), .B2(new_n871), .ZN(new_n872));
  OAI21_X1  g671(.A(new_n868), .B1(new_n872), .B2(KEYINPUT57), .ZN(new_n873));
  OAI21_X1  g672(.A(new_n577), .B1(new_n824), .B2(KEYINPUT119), .ZN(new_n874));
  AOI21_X1  g673(.A(new_n874), .B1(KEYINPUT119), .B2(new_n824), .ZN(new_n875));
  NAND3_X1  g674(.A1(new_n873), .A2(new_n875), .A3(KEYINPUT120), .ZN(new_n876));
  NAND2_X1  g675(.A1(new_n876), .A2(G148gat), .ZN(new_n877));
  AOI21_X1  g676(.A(KEYINPUT120), .B1(new_n873), .B2(new_n875), .ZN(new_n878));
  OAI21_X1  g677(.A(KEYINPUT59), .B1(new_n877), .B2(new_n878), .ZN(new_n879));
  NAND2_X1  g678(.A1(new_n867), .A2(new_n879), .ZN(new_n880));
  NOR2_X1   g679(.A1(new_n865), .A2(new_n866), .ZN(new_n881));
  OAI21_X1  g680(.A(new_n861), .B1(new_n880), .B2(new_n881), .ZN(G1345gat));
  OAI21_X1  g681(.A(G155gat), .B1(new_n864), .B2(new_n552), .ZN(new_n883));
  INV_X1    g682(.A(new_n853), .ZN(new_n884));
  NAND3_X1  g683(.A1(new_n884), .A2(new_n300), .A3(new_n554), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n883), .A2(new_n885), .ZN(G1346gat));
  AOI21_X1  g685(.A(new_n304), .B1(new_n884), .B2(new_n529), .ZN(new_n887));
  INV_X1    g686(.A(new_n864), .ZN(new_n888));
  AND2_X1   g687(.A1(new_n529), .A2(new_n304), .ZN(new_n889));
  AOI21_X1  g688(.A(new_n887), .B1(new_n888), .B2(new_n889), .ZN(G1347gat));
  NOR2_X1   g689(.A1(new_n803), .A2(new_n612), .ZN(new_n891));
  AND3_X1   g690(.A1(new_n891), .A2(new_n456), .A3(new_n471), .ZN(new_n892));
  AOI21_X1  g691(.A(G169gat), .B1(new_n892), .B2(new_n728), .ZN(new_n893));
  NOR3_X1   g692(.A1(new_n803), .A2(new_n442), .A3(new_n709), .ZN(new_n894));
  NAND2_X1  g693(.A1(new_n694), .A2(new_n456), .ZN(new_n895));
  INV_X1    g694(.A(new_n895), .ZN(new_n896));
  NAND2_X1  g695(.A1(new_n894), .A2(new_n896), .ZN(new_n897));
  NOR3_X1   g696(.A1(new_n897), .A2(new_n210), .A3(new_n608), .ZN(new_n898));
  NOR2_X1   g697(.A1(new_n893), .A2(new_n898), .ZN(G1348gat));
  AOI21_X1  g698(.A(G176gat), .B1(new_n892), .B2(new_n577), .ZN(new_n900));
  XNOR2_X1  g699(.A(new_n900), .B(KEYINPUT121), .ZN(new_n901));
  NOR3_X1   g700(.A1(new_n897), .A2(new_n211), .A3(new_n578), .ZN(new_n902));
  NOR2_X1   g701(.A1(new_n901), .A2(new_n902), .ZN(G1349gat));
  NAND3_X1  g702(.A1(new_n892), .A2(new_n205), .A3(new_n554), .ZN(new_n904));
  OAI21_X1  g703(.A(G183gat), .B1(new_n897), .B2(new_n552), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  XNOR2_X1  g705(.A(new_n906), .B(KEYINPUT60), .ZN(G1350gat));
  NAND3_X1  g706(.A1(new_n892), .A2(new_n206), .A3(new_n529), .ZN(new_n908));
  NAND3_X1  g707(.A1(new_n894), .A2(new_n529), .A3(new_n896), .ZN(new_n909));
  XNOR2_X1  g708(.A(KEYINPUT122), .B(KEYINPUT61), .ZN(new_n910));
  AND3_X1   g709(.A1(new_n909), .A2(G190gat), .A3(new_n910), .ZN(new_n911));
  AOI21_X1  g710(.A(new_n910), .B1(new_n909), .B2(G190gat), .ZN(new_n912));
  OAI21_X1  g711(.A(new_n908), .B1(new_n911), .B2(new_n912), .ZN(G1351gat));
  INV_X1    g712(.A(G197gat), .ZN(new_n914));
  NOR2_X1   g713(.A1(new_n895), .A2(new_n625), .ZN(new_n915));
  AND2_X1   g714(.A1(new_n873), .A2(new_n915), .ZN(new_n916));
  NAND2_X1  g715(.A1(new_n916), .A2(new_n728), .ZN(new_n917));
  AOI21_X1  g716(.A(new_n914), .B1(new_n917), .B2(KEYINPUT124), .ZN(new_n918));
  OAI21_X1  g717(.A(new_n918), .B1(KEYINPUT124), .B2(new_n917), .ZN(new_n919));
  NOR2_X1   g718(.A1(new_n851), .A2(new_n366), .ZN(new_n920));
  NAND2_X1  g719(.A1(new_n891), .A2(new_n920), .ZN(new_n921));
  XOR2_X1   g720(.A(new_n921), .B(KEYINPUT123), .Z(new_n922));
  NAND3_X1  g721(.A1(new_n922), .A2(new_n914), .A3(new_n728), .ZN(new_n923));
  NAND2_X1  g722(.A1(new_n919), .A2(new_n923), .ZN(G1352gat));
  INV_X1    g723(.A(G204gat), .ZN(new_n925));
  NAND2_X1  g724(.A1(new_n916), .A2(new_n577), .ZN(new_n926));
  AOI21_X1  g725(.A(new_n925), .B1(new_n926), .B2(KEYINPUT127), .ZN(new_n927));
  OAI21_X1  g726(.A(new_n927), .B1(KEYINPUT127), .B2(new_n926), .ZN(new_n928));
  NAND4_X1  g727(.A1(new_n891), .A2(new_n925), .A3(new_n577), .A4(new_n920), .ZN(new_n929));
  INV_X1    g728(.A(KEYINPUT125), .ZN(new_n930));
  OR2_X1    g729(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  NAND2_X1  g730(.A1(new_n929), .A2(new_n930), .ZN(new_n932));
  NAND2_X1  g731(.A1(new_n931), .A2(new_n932), .ZN(new_n933));
  OAI21_X1  g732(.A(new_n933), .B1(KEYINPUT126), .B2(KEYINPUT62), .ZN(new_n934));
  XNOR2_X1  g733(.A(KEYINPUT126), .B(KEYINPUT62), .ZN(new_n935));
  NAND3_X1  g734(.A1(new_n931), .A2(new_n932), .A3(new_n935), .ZN(new_n936));
  NAND3_X1  g735(.A1(new_n928), .A2(new_n934), .A3(new_n936), .ZN(G1353gat));
  NAND3_X1  g736(.A1(new_n922), .A2(new_n287), .A3(new_n554), .ZN(new_n938));
  NAND2_X1  g737(.A1(new_n916), .A2(new_n554), .ZN(new_n939));
  AND3_X1   g738(.A1(new_n939), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n940));
  AOI21_X1  g739(.A(KEYINPUT63), .B1(new_n939), .B2(G211gat), .ZN(new_n941));
  OAI21_X1  g740(.A(new_n938), .B1(new_n940), .B2(new_n941), .ZN(G1354gat));
  NAND3_X1  g741(.A1(new_n922), .A2(new_n288), .A3(new_n529), .ZN(new_n943));
  AND2_X1   g742(.A1(new_n916), .A2(new_n529), .ZN(new_n944));
  OAI21_X1  g743(.A(new_n943), .B1(new_n288), .B2(new_n944), .ZN(G1355gat));
endmodule


