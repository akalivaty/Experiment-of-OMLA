//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 1 0 0 0 1 1 0 1 1 1 1 1 0 1 0 0 0 1 1 1 0 0 0 0 1 1 1 1 0 0 0 0 0 0 0 0 0 1 0 0 0 1 1 1 0 1 1 0 1 0 1 0 1 1 0 0 1 1 0 0 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:25:07 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n703,
    new_n704, new_n705, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n719,
    new_n720, new_n721, new_n722, new_n724, new_n725, new_n727, new_n728,
    new_n729, new_n730, new_n731, new_n732, new_n733, new_n734, new_n736,
    new_n737, new_n738, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n758, new_n759,
    new_n760, new_n761, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n784, new_n785, new_n786, new_n787, new_n788, new_n789,
    new_n790, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n912, new_n913, new_n914, new_n915, new_n916, new_n917,
    new_n918, new_n919, new_n920, new_n921, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n938, new_n939, new_n940, new_n941,
    new_n942, new_n943, new_n944, new_n945, new_n946, new_n947, new_n948,
    new_n950, new_n951, new_n952, new_n953, new_n954, new_n955, new_n956,
    new_n957, new_n958, new_n959, new_n960, new_n961, new_n962, new_n963,
    new_n964, new_n965, new_n966, new_n967, new_n968, new_n969, new_n970,
    new_n971, new_n972, new_n974, new_n975, new_n976, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018;
  INV_X1    g000(.A(KEYINPUT70), .ZN(new_n187));
  XOR2_X1   g001(.A(KEYINPUT68), .B(KEYINPUT28), .Z(new_n188));
  INV_X1    g002(.A(KEYINPUT11), .ZN(new_n189));
  INV_X1    g003(.A(G134), .ZN(new_n190));
  OAI21_X1  g004(.A(new_n189), .B1(new_n190), .B2(G137), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n190), .A2(G137), .ZN(new_n192));
  INV_X1    g006(.A(G137), .ZN(new_n193));
  NAND3_X1  g007(.A1(new_n193), .A2(KEYINPUT11), .A3(G134), .ZN(new_n194));
  NAND3_X1  g008(.A1(new_n191), .A2(new_n192), .A3(new_n194), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n195), .A2(G131), .ZN(new_n196));
  INV_X1    g010(.A(G131), .ZN(new_n197));
  NAND4_X1  g011(.A1(new_n191), .A2(new_n194), .A3(new_n197), .A4(new_n192), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n196), .A2(new_n198), .ZN(new_n199));
  INV_X1    g013(.A(KEYINPUT66), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n199), .A2(new_n200), .ZN(new_n201));
  INV_X1    g015(.A(G146), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n202), .A2(G143), .ZN(new_n203));
  XNOR2_X1  g017(.A(KEYINPUT64), .B(G146), .ZN(new_n204));
  OAI21_X1  g018(.A(new_n203), .B1(new_n204), .B2(G143), .ZN(new_n205));
  AND2_X1   g019(.A1(KEYINPUT0), .A2(G128), .ZN(new_n206));
  NOR2_X1   g020(.A1(KEYINPUT0), .A2(G128), .ZN(new_n207));
  NOR2_X1   g021(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  NOR2_X1   g022(.A1(new_n202), .A2(G143), .ZN(new_n209));
  AOI21_X1  g023(.A(new_n209), .B1(new_n204), .B2(G143), .ZN(new_n210));
  AOI22_X1  g024(.A1(new_n205), .A2(new_n208), .B1(new_n210), .B2(new_n206), .ZN(new_n211));
  NAND3_X1  g025(.A1(new_n196), .A2(KEYINPUT66), .A3(new_n198), .ZN(new_n212));
  NAND3_X1  g026(.A1(new_n201), .A2(new_n211), .A3(new_n212), .ZN(new_n213));
  INV_X1    g027(.A(G113), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n214), .A2(KEYINPUT2), .ZN(new_n215));
  INV_X1    g029(.A(KEYINPUT2), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n216), .A2(G113), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n215), .A2(new_n217), .ZN(new_n218));
  XNOR2_X1  g032(.A(G116), .B(G119), .ZN(new_n219));
  XNOR2_X1  g033(.A(new_n218), .B(new_n219), .ZN(new_n220));
  INV_X1    g034(.A(new_n220), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n202), .A2(KEYINPUT64), .ZN(new_n222));
  INV_X1    g036(.A(KEYINPUT64), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n223), .A2(G146), .ZN(new_n224));
  NAND3_X1  g038(.A1(new_n222), .A2(new_n224), .A3(G143), .ZN(new_n225));
  INV_X1    g039(.A(new_n209), .ZN(new_n226));
  XNOR2_X1  g040(.A(KEYINPUT65), .B(KEYINPUT1), .ZN(new_n227));
  NAND4_X1  g041(.A1(new_n225), .A2(G128), .A3(new_n226), .A4(new_n227), .ZN(new_n228));
  INV_X1    g042(.A(G128), .ZN(new_n229));
  INV_X1    g043(.A(KEYINPUT1), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n230), .A2(KEYINPUT65), .ZN(new_n231));
  INV_X1    g045(.A(KEYINPUT65), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n232), .A2(KEYINPUT1), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n231), .A2(new_n233), .ZN(new_n234));
  AOI21_X1  g048(.A(new_n229), .B1(new_n225), .B2(new_n234), .ZN(new_n235));
  INV_X1    g049(.A(new_n203), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n222), .A2(new_n224), .ZN(new_n237));
  INV_X1    g051(.A(G143), .ZN(new_n238));
  AOI21_X1  g052(.A(new_n236), .B1(new_n237), .B2(new_n238), .ZN(new_n239));
  OAI21_X1  g053(.A(new_n228), .B1(new_n235), .B2(new_n239), .ZN(new_n240));
  INV_X1    g054(.A(new_n192), .ZN(new_n241));
  NOR2_X1   g055(.A1(new_n190), .A2(G137), .ZN(new_n242));
  OAI21_X1  g056(.A(G131), .B1(new_n241), .B2(new_n242), .ZN(new_n243));
  AND2_X1   g057(.A1(new_n243), .A2(new_n198), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n240), .A2(new_n244), .ZN(new_n245));
  AND3_X1   g059(.A1(new_n213), .A2(new_n221), .A3(new_n245), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n211), .A2(new_n199), .ZN(new_n247));
  AOI21_X1  g061(.A(new_n221), .B1(new_n247), .B2(new_n245), .ZN(new_n248));
  OAI21_X1  g062(.A(new_n188), .B1(new_n246), .B2(new_n248), .ZN(new_n249));
  NOR2_X1   g063(.A1(G237), .A2(G953), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n250), .A2(G210), .ZN(new_n251));
  XNOR2_X1  g065(.A(new_n251), .B(KEYINPUT27), .ZN(new_n252));
  XNOR2_X1  g066(.A(KEYINPUT26), .B(G101), .ZN(new_n253));
  XNOR2_X1  g067(.A(new_n252), .B(new_n253), .ZN(new_n254));
  NAND3_X1  g068(.A1(new_n213), .A2(new_n221), .A3(new_n245), .ZN(new_n255));
  INV_X1    g069(.A(KEYINPUT28), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  NAND3_X1  g071(.A1(new_n249), .A2(new_n254), .A3(new_n257), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n258), .A2(KEYINPUT69), .ZN(new_n259));
  INV_X1    g073(.A(KEYINPUT69), .ZN(new_n260));
  NAND4_X1  g074(.A1(new_n249), .A2(new_n260), .A3(new_n254), .A4(new_n257), .ZN(new_n261));
  INV_X1    g075(.A(KEYINPUT30), .ZN(new_n262));
  AND2_X1   g076(.A1(new_n240), .A2(new_n244), .ZN(new_n263));
  NAND3_X1  g077(.A1(new_n225), .A2(new_n206), .A3(new_n226), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n205), .A2(new_n208), .ZN(new_n265));
  AND3_X1   g079(.A1(new_n199), .A2(new_n264), .A3(new_n265), .ZN(new_n266));
  OAI21_X1  g080(.A(new_n262), .B1(new_n263), .B2(new_n266), .ZN(new_n267));
  NAND3_X1  g081(.A1(new_n213), .A2(KEYINPUT30), .A3(new_n245), .ZN(new_n268));
  NAND3_X1  g082(.A1(new_n267), .A2(new_n268), .A3(new_n220), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n269), .A2(new_n255), .ZN(new_n270));
  INV_X1    g084(.A(new_n254), .ZN(new_n271));
  AOI21_X1  g085(.A(KEYINPUT29), .B1(new_n270), .B2(new_n271), .ZN(new_n272));
  NAND3_X1  g086(.A1(new_n259), .A2(new_n261), .A3(new_n272), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n213), .A2(new_n245), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n274), .A2(new_n220), .ZN(new_n275));
  AOI21_X1  g089(.A(new_n256), .B1(new_n275), .B2(new_n255), .ZN(new_n276));
  INV_X1    g090(.A(new_n257), .ZN(new_n277));
  NOR2_X1   g091(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  AND2_X1   g092(.A1(new_n254), .A2(KEYINPUT29), .ZN(new_n279));
  AOI21_X1  g093(.A(G902), .B1(new_n278), .B2(new_n279), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n273), .A2(new_n280), .ZN(new_n281));
  AOI21_X1  g095(.A(new_n187), .B1(new_n281), .B2(G472), .ZN(new_n282));
  INV_X1    g096(.A(G472), .ZN(new_n283));
  AOI211_X1 g097(.A(KEYINPUT70), .B(new_n283), .C1(new_n273), .C2(new_n280), .ZN(new_n284));
  INV_X1    g098(.A(new_n188), .ZN(new_n285));
  INV_X1    g099(.A(new_n248), .ZN(new_n286));
  AOI21_X1  g100(.A(new_n285), .B1(new_n286), .B2(new_n255), .ZN(new_n287));
  OAI21_X1  g101(.A(new_n271), .B1(new_n287), .B2(new_n277), .ZN(new_n288));
  INV_X1    g102(.A(KEYINPUT31), .ZN(new_n289));
  NAND4_X1  g103(.A1(new_n269), .A2(new_n289), .A3(new_n254), .A4(new_n255), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n288), .A2(new_n290), .ZN(new_n291));
  NAND3_X1  g105(.A1(new_n269), .A2(new_n254), .A3(new_n255), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n292), .A2(KEYINPUT31), .ZN(new_n293));
  INV_X1    g107(.A(KEYINPUT67), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n293), .A2(new_n294), .ZN(new_n295));
  NAND3_X1  g109(.A1(new_n292), .A2(KEYINPUT67), .A3(KEYINPUT31), .ZN(new_n296));
  AOI21_X1  g110(.A(new_n291), .B1(new_n295), .B2(new_n296), .ZN(new_n297));
  NOR2_X1   g111(.A1(G472), .A2(G902), .ZN(new_n298));
  INV_X1    g112(.A(new_n298), .ZN(new_n299));
  NOR3_X1   g113(.A1(new_n297), .A2(KEYINPUT32), .A3(new_n299), .ZN(new_n300));
  INV_X1    g114(.A(KEYINPUT32), .ZN(new_n301));
  AND3_X1   g115(.A1(new_n292), .A2(KEYINPUT67), .A3(KEYINPUT31), .ZN(new_n302));
  AOI21_X1  g116(.A(KEYINPUT67), .B1(new_n292), .B2(KEYINPUT31), .ZN(new_n303));
  OAI211_X1 g117(.A(new_n288), .B(new_n290), .C1(new_n302), .C2(new_n303), .ZN(new_n304));
  AOI21_X1  g118(.A(new_n301), .B1(new_n304), .B2(new_n298), .ZN(new_n305));
  OAI22_X1  g119(.A1(new_n282), .A2(new_n284), .B1(new_n300), .B2(new_n305), .ZN(new_n306));
  XNOR2_X1  g120(.A(KEYINPUT22), .B(G137), .ZN(new_n307));
  INV_X1    g121(.A(G953), .ZN(new_n308));
  NAND3_X1  g122(.A1(new_n308), .A2(G221), .A3(G234), .ZN(new_n309));
  XNOR2_X1  g123(.A(new_n307), .B(new_n309), .ZN(new_n310));
  XOR2_X1   g124(.A(G119), .B(G128), .Z(new_n311));
  XNOR2_X1  g125(.A(KEYINPUT24), .B(G110), .ZN(new_n312));
  NOR2_X1   g126(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  INV_X1    g127(.A(G110), .ZN(new_n314));
  OAI211_X1 g128(.A(new_n229), .B(G119), .C1(KEYINPUT72), .C2(KEYINPUT23), .ZN(new_n315));
  INV_X1    g129(.A(KEYINPUT23), .ZN(new_n316));
  INV_X1    g130(.A(G119), .ZN(new_n317));
  AOI21_X1  g131(.A(new_n316), .B1(new_n317), .B2(G128), .ZN(new_n318));
  INV_X1    g132(.A(KEYINPUT72), .ZN(new_n319));
  OAI21_X1  g133(.A(new_n319), .B1(new_n317), .B2(G128), .ZN(new_n320));
  OAI21_X1  g134(.A(new_n315), .B1(new_n318), .B2(new_n320), .ZN(new_n321));
  INV_X1    g135(.A(KEYINPUT73), .ZN(new_n322));
  AOI21_X1  g136(.A(new_n314), .B1(new_n321), .B2(new_n322), .ZN(new_n323));
  OAI211_X1 g137(.A(KEYINPUT73), .B(new_n315), .C1(new_n318), .C2(new_n320), .ZN(new_n324));
  AOI21_X1  g138(.A(new_n313), .B1(new_n323), .B2(new_n324), .ZN(new_n325));
  INV_X1    g139(.A(G140), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n326), .A2(G125), .ZN(new_n327));
  INV_X1    g141(.A(G125), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n328), .A2(G140), .ZN(new_n329));
  NAND3_X1  g143(.A1(new_n327), .A2(new_n329), .A3(KEYINPUT16), .ZN(new_n330));
  INV_X1    g144(.A(KEYINPUT16), .ZN(new_n331));
  NAND3_X1  g145(.A1(new_n331), .A2(new_n326), .A3(G125), .ZN(new_n332));
  INV_X1    g146(.A(KEYINPUT74), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  NAND4_X1  g148(.A1(new_n331), .A2(new_n326), .A3(KEYINPUT74), .A4(G125), .ZN(new_n335));
  NAND3_X1  g149(.A1(new_n330), .A2(new_n334), .A3(new_n335), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n336), .A2(new_n202), .ZN(new_n337));
  NAND4_X1  g151(.A1(new_n330), .A2(new_n334), .A3(G146), .A4(new_n335), .ZN(new_n338));
  NAND3_X1  g152(.A1(new_n337), .A2(KEYINPUT75), .A3(new_n338), .ZN(new_n339));
  INV_X1    g153(.A(KEYINPUT75), .ZN(new_n340));
  NAND3_X1  g154(.A1(new_n336), .A2(new_n340), .A3(new_n202), .ZN(new_n341));
  NAND3_X1  g155(.A1(new_n325), .A2(new_n339), .A3(new_n341), .ZN(new_n342));
  XNOR2_X1  g156(.A(G125), .B(G140), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n204), .A2(new_n343), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n311), .A2(new_n312), .ZN(new_n345));
  OAI211_X1 g159(.A(new_n314), .B(new_n315), .C1(new_n318), .C2(new_n320), .ZN(new_n346));
  INV_X1    g160(.A(KEYINPUT76), .ZN(new_n347));
  AND3_X1   g161(.A1(new_n345), .A2(new_n346), .A3(new_n347), .ZN(new_n348));
  AOI21_X1  g162(.A(new_n347), .B1(new_n345), .B2(new_n346), .ZN(new_n349));
  OAI211_X1 g163(.A(new_n338), .B(new_n344), .C1(new_n348), .C2(new_n349), .ZN(new_n350));
  AOI21_X1  g164(.A(new_n310), .B1(new_n342), .B2(new_n350), .ZN(new_n351));
  INV_X1    g165(.A(new_n351), .ZN(new_n352));
  NAND3_X1  g166(.A1(new_n342), .A2(new_n350), .A3(new_n310), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n352), .A2(new_n353), .ZN(new_n354));
  INV_X1    g168(.A(G234), .ZN(new_n355));
  OAI21_X1  g169(.A(G217), .B1(new_n355), .B2(G902), .ZN(new_n356));
  INV_X1    g170(.A(G902), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  NOR2_X1   g172(.A1(new_n354), .A2(new_n358), .ZN(new_n359));
  INV_X1    g173(.A(KEYINPUT77), .ZN(new_n360));
  NAND3_X1  g174(.A1(new_n352), .A2(new_n357), .A3(new_n353), .ZN(new_n361));
  INV_X1    g175(.A(KEYINPUT25), .ZN(new_n362));
  AOI21_X1  g176(.A(new_n360), .B1(new_n361), .B2(new_n362), .ZN(new_n363));
  OAI21_X1  g177(.A(new_n363), .B1(new_n362), .B2(new_n361), .ZN(new_n364));
  NAND3_X1  g178(.A1(new_n361), .A2(new_n360), .A3(new_n362), .ZN(new_n365));
  XNOR2_X1  g179(.A(new_n356), .B(KEYINPUT71), .ZN(new_n366));
  INV_X1    g180(.A(new_n366), .ZN(new_n367));
  AND2_X1   g181(.A1(new_n365), .A2(new_n367), .ZN(new_n368));
  AOI21_X1  g182(.A(new_n359), .B1(new_n364), .B2(new_n368), .ZN(new_n369));
  INV_X1    g183(.A(G469), .ZN(new_n370));
  INV_X1    g184(.A(G104), .ZN(new_n371));
  OAI21_X1  g185(.A(KEYINPUT3), .B1(new_n371), .B2(G107), .ZN(new_n372));
  INV_X1    g186(.A(KEYINPUT3), .ZN(new_n373));
  INV_X1    g187(.A(G107), .ZN(new_n374));
  NAND3_X1  g188(.A1(new_n373), .A2(new_n374), .A3(G104), .ZN(new_n375));
  INV_X1    g189(.A(G101), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n371), .A2(G107), .ZN(new_n377));
  NAND4_X1  g191(.A1(new_n372), .A2(new_n375), .A3(new_n376), .A4(new_n377), .ZN(new_n378));
  NOR2_X1   g192(.A1(new_n374), .A2(G104), .ZN(new_n379));
  NOR2_X1   g193(.A1(new_n371), .A2(G107), .ZN(new_n380));
  OAI21_X1  g194(.A(G101), .B1(new_n379), .B2(new_n380), .ZN(new_n381));
  AND2_X1   g195(.A1(new_n378), .A2(new_n381), .ZN(new_n382));
  AND4_X1   g196(.A1(G128), .A2(new_n225), .A3(new_n226), .A4(new_n227), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n203), .A2(KEYINPUT1), .ZN(new_n384));
  AOI22_X1  g198(.A1(new_n225), .A2(new_n226), .B1(new_n384), .B2(G128), .ZN(new_n385));
  OAI21_X1  g199(.A(new_n382), .B1(new_n383), .B2(new_n385), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n378), .A2(new_n381), .ZN(new_n387));
  OAI211_X1 g201(.A(new_n387), .B(new_n228), .C1(new_n235), .C2(new_n239), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n386), .A2(new_n388), .ZN(new_n389));
  INV_X1    g203(.A(new_n212), .ZN(new_n390));
  AOI21_X1  g204(.A(KEYINPUT66), .B1(new_n196), .B2(new_n198), .ZN(new_n391));
  NOR2_X1   g205(.A1(new_n390), .A2(new_n391), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n389), .A2(new_n392), .ZN(new_n393));
  INV_X1    g207(.A(KEYINPUT12), .ZN(new_n394));
  AOI21_X1  g208(.A(new_n394), .B1(new_n196), .B2(new_n198), .ZN(new_n395));
  AOI22_X1  g209(.A1(new_n393), .A2(new_n394), .B1(new_n389), .B2(new_n395), .ZN(new_n396));
  INV_X1    g210(.A(KEYINPUT10), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n386), .A2(new_n397), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n387), .A2(KEYINPUT79), .ZN(new_n399));
  INV_X1    g213(.A(KEYINPUT79), .ZN(new_n400));
  NAND3_X1  g214(.A1(new_n378), .A2(new_n381), .A3(new_n400), .ZN(new_n401));
  NAND4_X1  g215(.A1(new_n240), .A2(KEYINPUT10), .A3(new_n399), .A4(new_n401), .ZN(new_n402));
  NAND3_X1  g216(.A1(new_n372), .A2(new_n375), .A3(new_n377), .ZN(new_n403));
  INV_X1    g217(.A(KEYINPUT4), .ZN(new_n404));
  NAND3_X1  g218(.A1(new_n403), .A2(new_n404), .A3(G101), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n403), .A2(G101), .ZN(new_n406));
  NAND3_X1  g220(.A1(new_n406), .A2(KEYINPUT4), .A3(new_n378), .ZN(new_n407));
  NAND3_X1  g221(.A1(new_n211), .A2(new_n405), .A3(new_n407), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n201), .A2(new_n212), .ZN(new_n409));
  NAND4_X1  g223(.A1(new_n398), .A2(new_n402), .A3(new_n408), .A4(new_n409), .ZN(new_n410));
  XNOR2_X1  g224(.A(G110), .B(G140), .ZN(new_n411));
  AND2_X1   g225(.A1(new_n308), .A2(G227), .ZN(new_n412));
  XNOR2_X1  g226(.A(new_n411), .B(new_n412), .ZN(new_n413));
  INV_X1    g227(.A(new_n413), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n410), .A2(new_n414), .ZN(new_n415));
  NOR2_X1   g229(.A1(new_n396), .A2(new_n415), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n407), .A2(new_n405), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n265), .A2(new_n264), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n225), .A2(new_n226), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n384), .A2(G128), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  AOI21_X1  g235(.A(new_n387), .B1(new_n421), .B2(new_n228), .ZN(new_n422));
  OAI22_X1  g236(.A1(new_n417), .A2(new_n418), .B1(new_n422), .B2(KEYINPUT10), .ZN(new_n423));
  INV_X1    g237(.A(new_n402), .ZN(new_n424));
  OAI21_X1  g238(.A(new_n392), .B1(new_n423), .B2(new_n424), .ZN(new_n425));
  AOI21_X1  g239(.A(new_n414), .B1(new_n425), .B2(new_n410), .ZN(new_n426));
  OAI211_X1 g240(.A(new_n370), .B(new_n357), .C1(new_n416), .C2(new_n426), .ZN(new_n427));
  INV_X1    g241(.A(new_n410), .ZN(new_n428));
  OAI21_X1  g242(.A(new_n413), .B1(new_n396), .B2(new_n428), .ZN(new_n429));
  NAND3_X1  g243(.A1(new_n425), .A2(new_n410), .A3(new_n414), .ZN(new_n430));
  NAND3_X1  g244(.A1(new_n429), .A2(G469), .A3(new_n430), .ZN(new_n431));
  NOR2_X1   g245(.A1(new_n370), .A2(new_n357), .ZN(new_n432));
  INV_X1    g246(.A(new_n432), .ZN(new_n433));
  NAND3_X1  g247(.A1(new_n427), .A2(new_n431), .A3(new_n433), .ZN(new_n434));
  XOR2_X1   g248(.A(KEYINPUT9), .B(G234), .Z(new_n435));
  XNOR2_X1  g249(.A(new_n435), .B(KEYINPUT78), .ZN(new_n436));
  OAI21_X1  g250(.A(G221), .B1(new_n436), .B2(G902), .ZN(new_n437));
  AND3_X1   g251(.A1(new_n434), .A2(KEYINPUT80), .A3(new_n437), .ZN(new_n438));
  OAI21_X1  g252(.A(G214), .B1(G237), .B2(G902), .ZN(new_n439));
  OAI21_X1  g253(.A(G210), .B1(G237), .B2(G902), .ZN(new_n440));
  XNOR2_X1  g254(.A(G110), .B(G122), .ZN(new_n441));
  INV_X1    g255(.A(new_n441), .ZN(new_n442));
  AND3_X1   g256(.A1(new_n407), .A2(new_n220), .A3(new_n405), .ZN(new_n443));
  AND3_X1   g257(.A1(new_n378), .A2(new_n381), .A3(new_n400), .ZN(new_n444));
  AOI21_X1  g258(.A(new_n400), .B1(new_n378), .B2(new_n381), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n218), .A2(new_n219), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n317), .A2(G116), .ZN(new_n447));
  INV_X1    g261(.A(G116), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n448), .A2(G119), .ZN(new_n449));
  AND3_X1   g263(.A1(new_n447), .A2(new_n449), .A3(KEYINPUT5), .ZN(new_n450));
  OAI21_X1  g264(.A(G113), .B1(new_n447), .B2(KEYINPUT5), .ZN(new_n451));
  OAI21_X1  g265(.A(new_n446), .B1(new_n450), .B2(new_n451), .ZN(new_n452));
  NOR3_X1   g266(.A1(new_n444), .A2(new_n445), .A3(new_n452), .ZN(new_n453));
  OAI21_X1  g267(.A(new_n442), .B1(new_n443), .B2(new_n453), .ZN(new_n454));
  INV_X1    g268(.A(new_n452), .ZN(new_n455));
  NAND3_X1  g269(.A1(new_n455), .A2(new_n399), .A3(new_n401), .ZN(new_n456));
  NAND3_X1  g270(.A1(new_n407), .A2(new_n220), .A3(new_n405), .ZN(new_n457));
  NAND3_X1  g271(.A1(new_n456), .A2(new_n457), .A3(new_n441), .ZN(new_n458));
  NAND3_X1  g272(.A1(new_n454), .A2(KEYINPUT6), .A3(new_n458), .ZN(new_n459));
  INV_X1    g273(.A(KEYINPUT6), .ZN(new_n460));
  OAI211_X1 g274(.A(new_n460), .B(new_n442), .C1(new_n443), .C2(new_n453), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n240), .A2(new_n328), .ZN(new_n462));
  NAND3_X1  g276(.A1(new_n265), .A2(G125), .A3(new_n264), .ZN(new_n463));
  XNOR2_X1  g277(.A(KEYINPUT81), .B(G224), .ZN(new_n464));
  OR2_X1    g278(.A1(new_n464), .A2(G953), .ZN(new_n465));
  AND3_X1   g279(.A1(new_n462), .A2(new_n463), .A3(new_n465), .ZN(new_n466));
  AOI21_X1  g280(.A(new_n465), .B1(new_n462), .B2(new_n463), .ZN(new_n467));
  NOR2_X1   g281(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  AND3_X1   g282(.A1(new_n459), .A2(new_n461), .A3(new_n468), .ZN(new_n469));
  INV_X1    g283(.A(KEYINPUT83), .ZN(new_n470));
  AND2_X1   g284(.A1(new_n465), .A2(KEYINPUT7), .ZN(new_n471));
  AOI22_X1  g285(.A1(new_n204), .A2(G143), .B1(new_n231), .B2(new_n233), .ZN(new_n472));
  OAI21_X1  g286(.A(new_n205), .B1(new_n472), .B2(new_n229), .ZN(new_n473));
  AOI21_X1  g287(.A(G125), .B1(new_n473), .B2(new_n228), .ZN(new_n474));
  AND3_X1   g288(.A1(new_n265), .A2(G125), .A3(new_n264), .ZN(new_n475));
  OAI21_X1  g289(.A(new_n471), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  XOR2_X1   g290(.A(KEYINPUT82), .B(KEYINPUT7), .Z(new_n477));
  NAND2_X1  g291(.A1(new_n465), .A2(new_n477), .ZN(new_n478));
  NAND3_X1  g292(.A1(new_n462), .A2(new_n463), .A3(new_n478), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n455), .A2(new_n387), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n382), .A2(new_n452), .ZN(new_n481));
  XNOR2_X1  g295(.A(new_n441), .B(KEYINPUT8), .ZN(new_n482));
  NAND3_X1  g296(.A1(new_n480), .A2(new_n481), .A3(new_n482), .ZN(new_n483));
  NAND4_X1  g297(.A1(new_n476), .A2(new_n458), .A3(new_n479), .A4(new_n483), .ZN(new_n484));
  AOI21_X1  g298(.A(new_n470), .B1(new_n484), .B2(new_n357), .ZN(new_n485));
  NOR2_X1   g299(.A1(new_n469), .A2(new_n485), .ZN(new_n486));
  NAND3_X1  g300(.A1(new_n484), .A2(new_n470), .A3(new_n357), .ZN(new_n487));
  AOI21_X1  g301(.A(new_n440), .B1(new_n486), .B2(new_n487), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n484), .A2(new_n357), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n489), .A2(KEYINPUT83), .ZN(new_n490));
  NAND3_X1  g304(.A1(new_n459), .A2(new_n461), .A3(new_n468), .ZN(new_n491));
  NAND4_X1  g305(.A1(new_n490), .A2(new_n440), .A3(new_n487), .A4(new_n491), .ZN(new_n492));
  INV_X1    g306(.A(new_n492), .ZN(new_n493));
  OAI21_X1  g307(.A(new_n439), .B1(new_n488), .B2(new_n493), .ZN(new_n494));
  AOI21_X1  g308(.A(KEYINPUT80), .B1(new_n434), .B2(new_n437), .ZN(new_n495));
  NOR3_X1   g309(.A1(new_n438), .A2(new_n494), .A3(new_n495), .ZN(new_n496));
  INV_X1    g310(.A(KEYINPUT20), .ZN(new_n497));
  AND3_X1   g311(.A1(new_n250), .A2(G143), .A3(G214), .ZN(new_n498));
  AOI21_X1  g312(.A(G143), .B1(new_n250), .B2(G214), .ZN(new_n499));
  NOR2_X1   g313(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  INV_X1    g314(.A(KEYINPUT18), .ZN(new_n501));
  NOR2_X1   g315(.A1(new_n501), .A2(new_n197), .ZN(new_n502));
  INV_X1    g316(.A(new_n502), .ZN(new_n503));
  OAI21_X1  g317(.A(KEYINPUT84), .B1(new_n500), .B2(new_n503), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n250), .A2(G214), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n505), .A2(new_n238), .ZN(new_n506));
  NAND3_X1  g320(.A1(new_n250), .A2(G143), .A3(G214), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  INV_X1    g322(.A(KEYINPUT84), .ZN(new_n509));
  NAND3_X1  g323(.A1(new_n508), .A2(new_n509), .A3(new_n502), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n504), .A2(new_n510), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n500), .A2(new_n503), .ZN(new_n512));
  OAI21_X1  g326(.A(new_n344), .B1(new_n202), .B2(new_n343), .ZN(new_n513));
  NAND3_X1  g327(.A1(new_n511), .A2(new_n512), .A3(new_n513), .ZN(new_n514));
  XNOR2_X1  g328(.A(G113), .B(G122), .ZN(new_n515));
  XNOR2_X1  g329(.A(KEYINPUT86), .B(G104), .ZN(new_n516));
  XOR2_X1   g330(.A(new_n515), .B(new_n516), .Z(new_n517));
  INV_X1    g331(.A(new_n517), .ZN(new_n518));
  INV_X1    g332(.A(KEYINPUT87), .ZN(new_n519));
  NAND3_X1  g333(.A1(new_n339), .A2(new_n519), .A3(new_n341), .ZN(new_n520));
  OAI21_X1  g334(.A(G131), .B1(new_n498), .B2(new_n499), .ZN(new_n521));
  INV_X1    g335(.A(KEYINPUT17), .ZN(new_n522));
  NOR2_X1   g336(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  NAND3_X1  g337(.A1(new_n506), .A2(new_n197), .A3(new_n507), .ZN(new_n524));
  AND2_X1   g338(.A1(new_n521), .A2(new_n524), .ZN(new_n525));
  AOI21_X1  g339(.A(new_n523), .B1(new_n525), .B2(new_n522), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n520), .A2(new_n526), .ZN(new_n527));
  AOI21_X1  g341(.A(new_n519), .B1(new_n339), .B2(new_n341), .ZN(new_n528));
  OAI211_X1 g342(.A(new_n514), .B(new_n518), .C1(new_n527), .C2(new_n528), .ZN(new_n529));
  INV_X1    g343(.A(new_n338), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n343), .A2(KEYINPUT85), .ZN(new_n531));
  INV_X1    g345(.A(KEYINPUT19), .ZN(new_n532));
  XNOR2_X1  g346(.A(new_n531), .B(new_n532), .ZN(new_n533));
  AOI211_X1 g347(.A(new_n530), .B(new_n525), .C1(new_n204), .C2(new_n533), .ZN(new_n534));
  INV_X1    g348(.A(new_n514), .ZN(new_n535));
  OAI21_X1  g349(.A(new_n517), .B1(new_n534), .B2(new_n535), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n529), .A2(new_n536), .ZN(new_n537));
  NOR2_X1   g351(.A1(G475), .A2(G902), .ZN(new_n538));
  XNOR2_X1  g352(.A(new_n538), .B(KEYINPUT88), .ZN(new_n539));
  INV_X1    g353(.A(new_n539), .ZN(new_n540));
  AOI21_X1  g354(.A(new_n497), .B1(new_n537), .B2(new_n540), .ZN(new_n541));
  AOI211_X1 g355(.A(KEYINPUT20), .B(new_n539), .C1(new_n529), .C2(new_n536), .ZN(new_n542));
  OAI21_X1  g356(.A(new_n514), .B1(new_n527), .B2(new_n528), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n543), .A2(new_n517), .ZN(new_n544));
  AOI21_X1  g358(.A(G902), .B1(new_n544), .B2(new_n529), .ZN(new_n545));
  INV_X1    g359(.A(G475), .ZN(new_n546));
  OAI22_X1  g360(.A1(new_n541), .A2(new_n542), .B1(new_n545), .B2(new_n546), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n308), .A2(G952), .ZN(new_n548));
  AOI21_X1  g362(.A(new_n548), .B1(G234), .B2(G237), .ZN(new_n549));
  INV_X1    g363(.A(new_n549), .ZN(new_n550));
  NAND2_X1  g364(.A1(G234), .A2(G237), .ZN(new_n551));
  NAND3_X1  g365(.A1(new_n551), .A2(G902), .A3(G953), .ZN(new_n552));
  XNOR2_X1  g366(.A(new_n552), .B(KEYINPUT92), .ZN(new_n553));
  XNOR2_X1  g367(.A(KEYINPUT21), .B(G898), .ZN(new_n554));
  INV_X1    g368(.A(new_n554), .ZN(new_n555));
  OAI21_X1  g369(.A(new_n550), .B1(new_n553), .B2(new_n555), .ZN(new_n556));
  INV_X1    g370(.A(KEYINPUT91), .ZN(new_n557));
  INV_X1    g371(.A(G217), .ZN(new_n558));
  NOR3_X1   g372(.A1(new_n436), .A2(new_n558), .A3(G953), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n448), .A2(G122), .ZN(new_n560));
  INV_X1    g374(.A(KEYINPUT14), .ZN(new_n561));
  OAI21_X1  g375(.A(new_n561), .B1(new_n448), .B2(G122), .ZN(new_n562));
  NAND3_X1  g376(.A1(new_n561), .A2(new_n448), .A3(G122), .ZN(new_n563));
  INV_X1    g377(.A(KEYINPUT90), .ZN(new_n564));
  AOI22_X1  g378(.A1(new_n560), .A2(new_n562), .B1(new_n563), .B2(new_n564), .ZN(new_n565));
  OR2_X1    g379(.A1(new_n563), .A2(new_n564), .ZN(new_n566));
  AOI21_X1  g380(.A(new_n374), .B1(new_n565), .B2(new_n566), .ZN(new_n567));
  OR2_X1    g381(.A1(new_n448), .A2(G122), .ZN(new_n568));
  NAND3_X1  g382(.A1(new_n568), .A2(new_n560), .A3(new_n374), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n238), .A2(G128), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n229), .A2(G143), .ZN(new_n571));
  AND3_X1   g385(.A1(new_n570), .A2(new_n571), .A3(new_n190), .ZN(new_n572));
  AOI21_X1  g386(.A(new_n190), .B1(new_n570), .B2(new_n571), .ZN(new_n573));
  OAI21_X1  g387(.A(new_n569), .B1(new_n572), .B2(new_n573), .ZN(new_n574));
  OR2_X1    g388(.A1(new_n567), .A2(new_n574), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n568), .A2(new_n560), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n576), .A2(G107), .ZN(new_n577));
  AOI21_X1  g391(.A(new_n572), .B1(new_n577), .B2(new_n569), .ZN(new_n578));
  INV_X1    g392(.A(KEYINPUT13), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n570), .A2(new_n579), .ZN(new_n580));
  NAND3_X1  g394(.A1(new_n238), .A2(KEYINPUT13), .A3(G128), .ZN(new_n581));
  NAND3_X1  g395(.A1(new_n580), .A2(new_n581), .A3(new_n571), .ZN(new_n582));
  AND3_X1   g396(.A1(new_n582), .A2(KEYINPUT89), .A3(G134), .ZN(new_n583));
  AOI21_X1  g397(.A(KEYINPUT89), .B1(new_n582), .B2(G134), .ZN(new_n584));
  OAI21_X1  g398(.A(new_n578), .B1(new_n583), .B2(new_n584), .ZN(new_n585));
  NAND3_X1  g399(.A1(new_n559), .A2(new_n575), .A3(new_n585), .ZN(new_n586));
  INV_X1    g400(.A(new_n586), .ZN(new_n587));
  AOI21_X1  g401(.A(new_n559), .B1(new_n585), .B2(new_n575), .ZN(new_n588));
  OAI211_X1 g402(.A(new_n557), .B(new_n357), .C1(new_n587), .C2(new_n588), .ZN(new_n589));
  INV_X1    g403(.A(G478), .ZN(new_n590));
  NOR2_X1   g404(.A1(new_n590), .A2(KEYINPUT15), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n589), .A2(new_n591), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n575), .A2(new_n585), .ZN(new_n593));
  INV_X1    g407(.A(new_n559), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  AOI21_X1  g409(.A(G902), .B1(new_n595), .B2(new_n586), .ZN(new_n596));
  NOR2_X1   g410(.A1(new_n596), .A2(new_n557), .ZN(new_n597));
  NOR2_X1   g411(.A1(new_n592), .A2(new_n597), .ZN(new_n598));
  NOR3_X1   g412(.A1(new_n596), .A2(new_n557), .A3(new_n591), .ZN(new_n599));
  OAI21_X1  g413(.A(new_n556), .B1(new_n598), .B2(new_n599), .ZN(new_n600));
  NOR2_X1   g414(.A1(new_n547), .A2(new_n600), .ZN(new_n601));
  NAND4_X1  g415(.A1(new_n306), .A2(new_n369), .A3(new_n496), .A4(new_n601), .ZN(new_n602));
  XNOR2_X1  g416(.A(new_n602), .B(G101), .ZN(G3));
  OAI21_X1  g417(.A(G472), .B1(new_n297), .B2(G902), .ZN(new_n604));
  OAI21_X1  g418(.A(new_n604), .B1(new_n299), .B2(new_n297), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n434), .A2(new_n437), .ZN(new_n606));
  INV_X1    g420(.A(KEYINPUT80), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  NAND3_X1  g422(.A1(new_n434), .A2(KEYINPUT80), .A3(new_n437), .ZN(new_n609));
  NAND3_X1  g423(.A1(new_n608), .A2(new_n369), .A3(new_n609), .ZN(new_n610));
  NOR2_X1   g424(.A1(new_n605), .A2(new_n610), .ZN(new_n611));
  XNOR2_X1  g425(.A(new_n611), .B(KEYINPUT93), .ZN(new_n612));
  NOR2_X1   g426(.A1(new_n587), .A2(new_n588), .ZN(new_n613));
  INV_X1    g427(.A(KEYINPUT33), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  OAI21_X1  g429(.A(KEYINPUT33), .B1(new_n587), .B2(new_n588), .ZN(new_n616));
  NAND3_X1  g430(.A1(new_n615), .A2(G478), .A3(new_n616), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n596), .A2(new_n590), .ZN(new_n618));
  NAND2_X1  g432(.A1(G478), .A2(G902), .ZN(new_n619));
  NAND3_X1  g433(.A1(new_n617), .A2(new_n618), .A3(new_n619), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n537), .A2(new_n540), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n621), .A2(KEYINPUT20), .ZN(new_n622));
  NAND3_X1  g436(.A1(new_n537), .A2(new_n497), .A3(new_n540), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  OR2_X1    g438(.A1(new_n545), .A2(new_n546), .ZN(new_n625));
  AOI21_X1  g439(.A(new_n620), .B1(new_n624), .B2(new_n625), .ZN(new_n626));
  NAND3_X1  g440(.A1(new_n490), .A2(new_n487), .A3(new_n491), .ZN(new_n627));
  INV_X1    g441(.A(new_n440), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n629), .A2(new_n492), .ZN(new_n630));
  NAND3_X1  g444(.A1(new_n630), .A2(new_n439), .A3(new_n556), .ZN(new_n631));
  INV_X1    g445(.A(new_n631), .ZN(new_n632));
  NAND3_X1  g446(.A1(new_n612), .A2(new_n626), .A3(new_n632), .ZN(new_n633));
  XNOR2_X1  g447(.A(new_n633), .B(KEYINPUT94), .ZN(new_n634));
  XNOR2_X1  g448(.A(KEYINPUT34), .B(G104), .ZN(new_n635));
  XNOR2_X1  g449(.A(new_n634), .B(new_n635), .ZN(G6));
  OAI21_X1  g450(.A(KEYINPUT91), .B1(new_n613), .B2(G902), .ZN(new_n637));
  NAND3_X1  g451(.A1(new_n637), .A2(new_n589), .A3(new_n591), .ZN(new_n638));
  INV_X1    g452(.A(new_n599), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  NOR2_X1   g454(.A1(new_n547), .A2(new_n640), .ZN(new_n641));
  NAND3_X1  g455(.A1(new_n612), .A2(new_n632), .A3(new_n641), .ZN(new_n642));
  XOR2_X1   g456(.A(KEYINPUT35), .B(G107), .Z(new_n643));
  XNOR2_X1  g457(.A(new_n642), .B(new_n643), .ZN(G9));
  NAND2_X1  g458(.A1(new_n304), .A2(new_n357), .ZN(new_n645));
  AOI22_X1  g459(.A1(new_n645), .A2(G472), .B1(new_n298), .B2(new_n304), .ZN(new_n646));
  AND3_X1   g460(.A1(new_n342), .A2(new_n350), .A3(new_n310), .ZN(new_n647));
  NOR3_X1   g461(.A1(new_n647), .A2(new_n351), .A3(G902), .ZN(new_n648));
  OAI21_X1  g462(.A(KEYINPUT77), .B1(new_n648), .B2(KEYINPUT25), .ZN(new_n649));
  NOR2_X1   g463(.A1(new_n361), .A2(new_n362), .ZN(new_n650));
  OAI211_X1 g464(.A(new_n365), .B(new_n367), .C1(new_n649), .C2(new_n650), .ZN(new_n651));
  NAND2_X1  g465(.A1(new_n342), .A2(new_n350), .ZN(new_n652));
  INV_X1    g466(.A(new_n310), .ZN(new_n653));
  NOR2_X1   g467(.A1(new_n653), .A2(KEYINPUT36), .ZN(new_n654));
  XNOR2_X1  g468(.A(new_n652), .B(new_n654), .ZN(new_n655));
  NAND3_X1  g469(.A1(new_n655), .A2(new_n357), .A3(new_n356), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n651), .A2(new_n656), .ZN(new_n657));
  INV_X1    g471(.A(KEYINPUT95), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  NAND3_X1  g473(.A1(new_n651), .A2(KEYINPUT95), .A3(new_n656), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  NAND4_X1  g475(.A1(new_n496), .A2(new_n601), .A3(new_n646), .A4(new_n661), .ZN(new_n662));
  XNOR2_X1  g476(.A(new_n662), .B(KEYINPUT96), .ZN(new_n663));
  XNOR2_X1  g477(.A(KEYINPUT37), .B(G110), .ZN(new_n664));
  XNOR2_X1  g478(.A(new_n663), .B(new_n664), .ZN(G12));
  INV_X1    g479(.A(new_n439), .ZN(new_n666));
  AOI21_X1  g480(.A(new_n666), .B1(new_n629), .B2(new_n492), .ZN(new_n667));
  OAI21_X1  g481(.A(KEYINPUT97), .B1(new_n553), .B2(G900), .ZN(new_n668));
  NAND2_X1  g482(.A1(new_n668), .A2(new_n550), .ZN(new_n669));
  NOR3_X1   g483(.A1(new_n553), .A2(KEYINPUT97), .A3(G900), .ZN(new_n670));
  NOR2_X1   g484(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  XNOR2_X1  g485(.A(new_n671), .B(KEYINPUT98), .ZN(new_n672));
  INV_X1    g486(.A(new_n672), .ZN(new_n673));
  NOR3_X1   g487(.A1(new_n547), .A2(new_n640), .A3(new_n673), .ZN(new_n674));
  AND4_X1   g488(.A1(new_n667), .A2(new_n608), .A3(new_n674), .A4(new_n609), .ZN(new_n675));
  NAND3_X1  g489(.A1(new_n675), .A2(new_n306), .A3(new_n661), .ZN(new_n676));
  XNOR2_X1  g490(.A(new_n676), .B(G128), .ZN(G30));
  XNOR2_X1  g491(.A(KEYINPUT100), .B(KEYINPUT39), .ZN(new_n678));
  XNOR2_X1  g492(.A(new_n672), .B(new_n678), .ZN(new_n679));
  NOR3_X1   g493(.A1(new_n438), .A2(new_n495), .A3(new_n679), .ZN(new_n680));
  XNOR2_X1  g494(.A(new_n680), .B(KEYINPUT101), .ZN(new_n681));
  OR2_X1    g495(.A1(new_n681), .A2(KEYINPUT40), .ZN(new_n682));
  NAND2_X1  g496(.A1(new_n681), .A2(KEYINPUT40), .ZN(new_n683));
  OAI21_X1  g497(.A(KEYINPUT32), .B1(new_n297), .B2(new_n299), .ZN(new_n684));
  NAND3_X1  g498(.A1(new_n304), .A2(new_n301), .A3(new_n298), .ZN(new_n685));
  NAND2_X1  g499(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  NAND3_X1  g500(.A1(new_n275), .A2(new_n271), .A3(new_n255), .ZN(new_n687));
  NAND2_X1  g501(.A1(new_n687), .A2(new_n357), .ZN(new_n688));
  AOI21_X1  g502(.A(new_n271), .B1(new_n269), .B2(new_n255), .ZN(new_n689));
  OAI21_X1  g503(.A(G472), .B1(new_n688), .B2(new_n689), .ZN(new_n690));
  XOR2_X1   g504(.A(new_n690), .B(KEYINPUT99), .Z(new_n691));
  NAND2_X1  g505(.A1(new_n686), .A2(new_n691), .ZN(new_n692));
  AND3_X1   g506(.A1(new_n651), .A2(KEYINPUT95), .A3(new_n656), .ZN(new_n693));
  AOI21_X1  g507(.A(KEYINPUT95), .B1(new_n651), .B2(new_n656), .ZN(new_n694));
  NOR2_X1   g508(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  NOR2_X1   g509(.A1(new_n640), .A2(new_n666), .ZN(new_n696));
  NAND3_X1  g510(.A1(new_n695), .A2(new_n547), .A3(new_n696), .ZN(new_n697));
  XNOR2_X1  g511(.A(new_n630), .B(KEYINPUT38), .ZN(new_n698));
  INV_X1    g512(.A(new_n698), .ZN(new_n699));
  NOR2_X1   g513(.A1(new_n697), .A2(new_n699), .ZN(new_n700));
  NAND4_X1  g514(.A1(new_n682), .A2(new_n683), .A3(new_n692), .A4(new_n700), .ZN(new_n701));
  XNOR2_X1  g515(.A(new_n701), .B(G143), .ZN(G45));
  INV_X1    g516(.A(new_n620), .ZN(new_n703));
  AND3_X1   g517(.A1(new_n547), .A2(new_n703), .A3(new_n672), .ZN(new_n704));
  NAND4_X1  g518(.A1(new_n306), .A2(new_n496), .A3(new_n661), .A4(new_n704), .ZN(new_n705));
  XNOR2_X1  g519(.A(new_n705), .B(G146), .ZN(G48));
  OAI21_X1  g520(.A(new_n357), .B1(new_n416), .B2(new_n426), .ZN(new_n707));
  NAND2_X1  g521(.A1(new_n707), .A2(G469), .ZN(new_n708));
  NAND3_X1  g522(.A1(new_n708), .A2(new_n437), .A3(new_n427), .ZN(new_n709));
  INV_X1    g523(.A(KEYINPUT102), .ZN(new_n710));
  NAND2_X1  g524(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  NAND4_X1  g525(.A1(new_n708), .A2(KEYINPUT102), .A3(new_n437), .A4(new_n427), .ZN(new_n712));
  NAND3_X1  g526(.A1(new_n711), .A2(new_n369), .A3(new_n712), .ZN(new_n713));
  NAND3_X1  g527(.A1(new_n626), .A2(new_n667), .A3(new_n556), .ZN(new_n714));
  NOR2_X1   g528(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  NAND2_X1  g529(.A1(new_n715), .A2(new_n306), .ZN(new_n716));
  XNOR2_X1  g530(.A(KEYINPUT41), .B(G113), .ZN(new_n717));
  XNOR2_X1  g531(.A(new_n716), .B(new_n717), .ZN(G15));
  NAND3_X1  g532(.A1(new_n641), .A2(new_n667), .A3(new_n556), .ZN(new_n719));
  NOR2_X1   g533(.A1(new_n713), .A2(new_n719), .ZN(new_n720));
  NAND2_X1  g534(.A1(new_n720), .A2(new_n306), .ZN(new_n721));
  XNOR2_X1  g535(.A(KEYINPUT103), .B(G116), .ZN(new_n722));
  XNOR2_X1  g536(.A(new_n721), .B(new_n722), .ZN(G18));
  AND4_X1   g537(.A1(new_n667), .A2(new_n711), .A3(new_n601), .A4(new_n712), .ZN(new_n724));
  NAND3_X1  g538(.A1(new_n306), .A2(new_n724), .A3(new_n661), .ZN(new_n725));
  XNOR2_X1  g539(.A(new_n725), .B(G119), .ZN(G21));
  OAI211_X1 g540(.A(new_n293), .B(new_n290), .C1(new_n278), .C2(new_n254), .ZN(new_n727));
  NAND2_X1  g541(.A1(new_n727), .A2(new_n298), .ZN(new_n728));
  AND3_X1   g542(.A1(new_n604), .A2(new_n728), .A3(new_n369), .ZN(new_n729));
  AND3_X1   g543(.A1(new_n711), .A2(new_n556), .A3(new_n712), .ZN(new_n730));
  NAND3_X1  g544(.A1(new_n696), .A2(new_n630), .A3(new_n547), .ZN(new_n731));
  INV_X1    g545(.A(new_n731), .ZN(new_n732));
  NAND3_X1  g546(.A1(new_n729), .A2(new_n730), .A3(new_n732), .ZN(new_n733));
  XOR2_X1   g547(.A(KEYINPUT104), .B(G122), .Z(new_n734));
  XNOR2_X1  g548(.A(new_n733), .B(new_n734), .ZN(G24));
  OAI211_X1 g549(.A(new_n604), .B(new_n728), .C1(new_n693), .C2(new_n694), .ZN(new_n736));
  NAND4_X1  g550(.A1(new_n704), .A2(new_n667), .A3(new_n711), .A4(new_n712), .ZN(new_n737));
  NOR2_X1   g551(.A1(new_n736), .A2(new_n737), .ZN(new_n738));
  XNOR2_X1  g552(.A(new_n738), .B(new_n328), .ZN(G27));
  INV_X1    g553(.A(new_n369), .ZN(new_n740));
  NAND2_X1  g554(.A1(new_n281), .A2(G472), .ZN(new_n741));
  NAND2_X1  g555(.A1(new_n741), .A2(KEYINPUT70), .ZN(new_n742));
  NAND3_X1  g556(.A1(new_n281), .A2(new_n187), .A3(G472), .ZN(new_n743));
  NAND2_X1  g557(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  AOI21_X1  g558(.A(new_n740), .B1(new_n744), .B2(new_n686), .ZN(new_n745));
  NAND3_X1  g559(.A1(new_n629), .A2(new_n439), .A3(new_n492), .ZN(new_n746));
  INV_X1    g560(.A(KEYINPUT105), .ZN(new_n747));
  NAND2_X1  g561(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  NAND4_X1  g562(.A1(new_n629), .A2(KEYINPUT105), .A3(new_n439), .A4(new_n492), .ZN(new_n749));
  AND3_X1   g563(.A1(new_n434), .A2(new_n437), .A3(new_n672), .ZN(new_n750));
  AND4_X1   g564(.A1(new_n626), .A2(new_n748), .A3(new_n749), .A4(new_n750), .ZN(new_n751));
  NAND2_X1  g565(.A1(new_n745), .A2(new_n751), .ZN(new_n752));
  INV_X1    g566(.A(KEYINPUT42), .ZN(new_n753));
  NAND2_X1  g567(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  NAND3_X1  g568(.A1(new_n745), .A2(KEYINPUT42), .A3(new_n751), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  XNOR2_X1  g570(.A(new_n756), .B(G131), .ZN(G33));
  NAND2_X1  g571(.A1(new_n748), .A2(new_n749), .ZN(new_n758));
  INV_X1    g572(.A(new_n758), .ZN(new_n759));
  NOR4_X1   g573(.A1(new_n606), .A2(new_n547), .A3(new_n640), .A4(new_n673), .ZN(new_n760));
  NAND4_X1  g574(.A1(new_n306), .A2(new_n759), .A3(new_n369), .A4(new_n760), .ZN(new_n761));
  XNOR2_X1  g575(.A(new_n761), .B(G134), .ZN(G36));
  AND2_X1   g576(.A1(new_n429), .A2(new_n430), .ZN(new_n763));
  AND2_X1   g577(.A1(new_n763), .A2(KEYINPUT45), .ZN(new_n764));
  OAI21_X1  g578(.A(G469), .B1(new_n763), .B2(KEYINPUT45), .ZN(new_n765));
  NOR2_X1   g579(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  NOR2_X1   g580(.A1(new_n766), .A2(new_n432), .ZN(new_n767));
  OR2_X1    g581(.A1(new_n767), .A2(KEYINPUT46), .ZN(new_n768));
  NAND2_X1  g582(.A1(new_n767), .A2(KEYINPUT46), .ZN(new_n769));
  NAND3_X1  g583(.A1(new_n768), .A2(new_n427), .A3(new_n769), .ZN(new_n770));
  NAND2_X1  g584(.A1(new_n770), .A2(new_n437), .ZN(new_n771));
  NOR3_X1   g585(.A1(new_n771), .A2(new_n679), .A3(new_n758), .ZN(new_n772));
  NAND3_X1  g586(.A1(new_n703), .A2(new_n624), .A3(new_n625), .ZN(new_n773));
  INV_X1    g587(.A(KEYINPUT43), .ZN(new_n774));
  OAI21_X1  g588(.A(new_n773), .B1(KEYINPUT106), .B2(new_n774), .ZN(new_n775));
  XNOR2_X1  g589(.A(KEYINPUT106), .B(KEYINPUT43), .ZN(new_n776));
  OAI21_X1  g590(.A(new_n775), .B1(new_n773), .B2(new_n776), .ZN(new_n777));
  NAND3_X1  g591(.A1(new_n777), .A2(new_n605), .A3(new_n661), .ZN(new_n778));
  INV_X1    g592(.A(KEYINPUT44), .ZN(new_n779));
  OR2_X1    g593(.A1(new_n778), .A2(new_n779), .ZN(new_n780));
  NAND2_X1  g594(.A1(new_n778), .A2(new_n779), .ZN(new_n781));
  NAND3_X1  g595(.A1(new_n772), .A2(new_n780), .A3(new_n781), .ZN(new_n782));
  XNOR2_X1  g596(.A(new_n782), .B(G137), .ZN(G39));
  INV_X1    g597(.A(KEYINPUT47), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n771), .A2(new_n784), .ZN(new_n785));
  NAND3_X1  g599(.A1(new_n770), .A2(KEYINPUT47), .A3(new_n437), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  NAND2_X1  g601(.A1(new_n704), .A2(new_n740), .ZN(new_n788));
  NOR3_X1   g602(.A1(new_n306), .A2(new_n758), .A3(new_n788), .ZN(new_n789));
  NAND2_X1  g603(.A1(new_n787), .A2(new_n789), .ZN(new_n790));
  XNOR2_X1  g604(.A(new_n790), .B(G140), .ZN(G42));
  NAND2_X1  g605(.A1(new_n777), .A2(new_n549), .ZN(new_n792));
  INV_X1    g606(.A(new_n792), .ZN(new_n793));
  NAND2_X1  g607(.A1(new_n711), .A2(new_n712), .ZN(new_n794));
  NOR3_X1   g608(.A1(new_n698), .A2(new_n439), .A3(new_n794), .ZN(new_n795));
  NAND3_X1  g609(.A1(new_n793), .A2(new_n729), .A3(new_n795), .ZN(new_n796));
  XOR2_X1   g610(.A(new_n796), .B(KEYINPUT50), .Z(new_n797));
  OR2_X1    g611(.A1(new_n758), .A2(new_n794), .ZN(new_n798));
  NOR4_X1   g612(.A1(new_n798), .A2(new_n740), .A3(new_n692), .A4(new_n550), .ZN(new_n799));
  NOR2_X1   g613(.A1(new_n547), .A2(new_n703), .ZN(new_n800));
  NOR2_X1   g614(.A1(new_n792), .A2(new_n798), .ZN(new_n801));
  INV_X1    g615(.A(new_n736), .ZN(new_n802));
  AOI22_X1  g616(.A1(new_n799), .A2(new_n800), .B1(new_n801), .B2(new_n802), .ZN(new_n803));
  NAND2_X1  g617(.A1(new_n708), .A2(new_n427), .ZN(new_n804));
  NOR2_X1   g618(.A1(new_n804), .A2(new_n437), .ZN(new_n805));
  NOR2_X1   g619(.A1(new_n787), .A2(new_n805), .ZN(new_n806));
  NAND3_X1  g620(.A1(new_n793), .A2(new_n729), .A3(new_n759), .ZN(new_n807));
  OAI211_X1 g621(.A(new_n797), .B(new_n803), .C1(new_n806), .C2(new_n807), .ZN(new_n808));
  INV_X1    g622(.A(KEYINPUT51), .ZN(new_n809));
  OR2_X1    g623(.A1(new_n808), .A2(new_n809), .ZN(new_n810));
  NOR2_X1   g624(.A1(new_n794), .A2(new_n494), .ZN(new_n811));
  NAND3_X1  g625(.A1(new_n793), .A2(new_n811), .A3(new_n729), .ZN(new_n812));
  XNOR2_X1  g626(.A(new_n812), .B(KEYINPUT111), .ZN(new_n813));
  INV_X1    g627(.A(KEYINPUT112), .ZN(new_n814));
  AOI21_X1  g628(.A(new_n548), .B1(new_n799), .B2(new_n626), .ZN(new_n815));
  AND3_X1   g629(.A1(new_n813), .A2(new_n814), .A3(new_n815), .ZN(new_n816));
  AOI21_X1  g630(.A(new_n814), .B1(new_n813), .B2(new_n815), .ZN(new_n817));
  NAND2_X1  g631(.A1(new_n801), .A2(new_n745), .ZN(new_n818));
  INV_X1    g632(.A(KEYINPUT48), .ZN(new_n819));
  XNOR2_X1  g633(.A(new_n818), .B(new_n819), .ZN(new_n820));
  NOR3_X1   g634(.A1(new_n816), .A2(new_n817), .A3(new_n820), .ZN(new_n821));
  NAND2_X1  g635(.A1(new_n808), .A2(new_n809), .ZN(new_n822));
  NAND3_X1  g636(.A1(new_n810), .A2(new_n821), .A3(new_n822), .ZN(new_n823));
  INV_X1    g637(.A(KEYINPUT113), .ZN(new_n824));
  NAND2_X1  g638(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  NAND4_X1  g639(.A1(new_n810), .A2(KEYINPUT113), .A3(new_n821), .A4(new_n822), .ZN(new_n826));
  NAND2_X1  g640(.A1(new_n825), .A2(new_n826), .ZN(new_n827));
  AND2_X1   g641(.A1(new_n602), .A2(new_n725), .ZN(new_n828));
  AND2_X1   g642(.A1(new_n716), .A2(new_n662), .ZN(new_n829));
  AND2_X1   g643(.A1(new_n721), .A2(new_n733), .ZN(new_n830));
  INV_X1    g644(.A(KEYINPUT107), .ZN(new_n831));
  NAND2_X1  g645(.A1(new_n547), .A2(new_n703), .ZN(new_n832));
  OAI21_X1  g646(.A(new_n831), .B1(new_n631), .B2(new_n832), .ZN(new_n833));
  OAI21_X1  g647(.A(KEYINPUT108), .B1(new_n547), .B2(new_n640), .ZN(new_n834));
  NOR2_X1   g648(.A1(new_n598), .A2(new_n599), .ZN(new_n835));
  INV_X1    g649(.A(KEYINPUT108), .ZN(new_n836));
  NAND4_X1  g650(.A1(new_n624), .A2(new_n835), .A3(new_n625), .A4(new_n836), .ZN(new_n837));
  NAND4_X1  g651(.A1(new_n834), .A2(new_n837), .A3(new_n667), .A4(new_n556), .ZN(new_n838));
  NAND4_X1  g652(.A1(new_n626), .A2(new_n667), .A3(KEYINPUT107), .A4(new_n556), .ZN(new_n839));
  NAND3_X1  g653(.A1(new_n833), .A2(new_n838), .A3(new_n839), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n840), .A2(new_n611), .ZN(new_n841));
  NAND4_X1  g655(.A1(new_n828), .A2(new_n829), .A3(new_n830), .A4(new_n841), .ZN(new_n842));
  NAND4_X1  g656(.A1(new_n748), .A2(new_n750), .A3(new_n626), .A4(new_n749), .ZN(new_n843));
  NOR2_X1   g657(.A1(new_n736), .A2(new_n843), .ZN(new_n844));
  AOI21_X1  g658(.A(new_n695), .B1(new_n744), .B2(new_n686), .ZN(new_n845));
  NAND4_X1  g659(.A1(new_n624), .A2(new_n625), .A3(new_n640), .A4(new_n672), .ZN(new_n846));
  INV_X1    g660(.A(new_n846), .ZN(new_n847));
  NAND3_X1  g661(.A1(new_n847), .A2(new_n608), .A3(new_n609), .ZN(new_n848));
  NOR2_X1   g662(.A1(new_n848), .A2(new_n758), .ZN(new_n849));
  AOI21_X1  g663(.A(new_n844), .B1(new_n845), .B2(new_n849), .ZN(new_n850));
  AOI21_X1  g664(.A(KEYINPUT42), .B1(new_n745), .B2(new_n751), .ZN(new_n851));
  AND4_X1   g665(.A1(KEYINPUT42), .A2(new_n751), .A3(new_n306), .A4(new_n369), .ZN(new_n852));
  OAI211_X1 g666(.A(new_n761), .B(new_n850), .C1(new_n851), .C2(new_n852), .ZN(new_n853));
  INV_X1    g667(.A(KEYINPUT53), .ZN(new_n854));
  NOR3_X1   g668(.A1(new_n842), .A2(new_n853), .A3(new_n854), .ZN(new_n855));
  AOI21_X1  g669(.A(new_n738), .B1(new_n845), .B2(new_n675), .ZN(new_n856));
  NOR4_X1   g670(.A1(new_n731), .A2(new_n606), .A3(new_n657), .A4(new_n673), .ZN(new_n857));
  NAND2_X1  g671(.A1(new_n857), .A2(new_n692), .ZN(new_n858));
  NAND4_X1  g672(.A1(new_n856), .A2(KEYINPUT52), .A3(new_n705), .A4(new_n858), .ZN(new_n859));
  AND2_X1   g673(.A1(new_n604), .A2(new_n728), .ZN(new_n860));
  NAND4_X1  g674(.A1(new_n811), .A2(new_n860), .A3(new_n661), .A4(new_n704), .ZN(new_n861));
  NAND4_X1  g675(.A1(new_n676), .A2(new_n705), .A3(new_n861), .A4(new_n858), .ZN(new_n862));
  INV_X1    g676(.A(KEYINPUT52), .ZN(new_n863));
  NAND2_X1  g677(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  NAND2_X1  g678(.A1(new_n859), .A2(new_n864), .ZN(new_n865));
  NAND2_X1  g679(.A1(new_n865), .A2(KEYINPUT110), .ZN(new_n866));
  INV_X1    g680(.A(KEYINPUT110), .ZN(new_n867));
  NAND3_X1  g681(.A1(new_n859), .A2(new_n864), .A3(new_n867), .ZN(new_n868));
  NAND3_X1  g682(.A1(new_n855), .A2(new_n866), .A3(new_n868), .ZN(new_n869));
  INV_X1    g683(.A(KEYINPUT54), .ZN(new_n870));
  AND2_X1   g684(.A1(new_n859), .A2(new_n864), .ZN(new_n871));
  INV_X1    g685(.A(KEYINPUT109), .ZN(new_n872));
  OAI21_X1  g686(.A(new_n872), .B1(new_n842), .B2(new_n853), .ZN(new_n873));
  NOR3_X1   g687(.A1(new_n438), .A2(new_n846), .A3(new_n495), .ZN(new_n874));
  NAND4_X1  g688(.A1(new_n306), .A2(new_n759), .A3(new_n661), .A4(new_n874), .ZN(new_n875));
  NAND2_X1  g689(.A1(new_n802), .A2(new_n751), .ZN(new_n876));
  NAND3_X1  g690(.A1(new_n761), .A2(new_n875), .A3(new_n876), .ZN(new_n877));
  AOI21_X1  g691(.A(new_n877), .B1(new_n754), .B2(new_n755), .ZN(new_n878));
  NAND4_X1  g692(.A1(new_n716), .A2(new_n721), .A3(new_n662), .A4(new_n733), .ZN(new_n879));
  NAND2_X1  g693(.A1(new_n602), .A2(new_n725), .ZN(new_n880));
  AND2_X1   g694(.A1(new_n840), .A2(new_n611), .ZN(new_n881));
  NOR3_X1   g695(.A1(new_n879), .A2(new_n880), .A3(new_n881), .ZN(new_n882));
  NAND3_X1  g696(.A1(new_n878), .A2(new_n882), .A3(KEYINPUT109), .ZN(new_n883));
  AOI21_X1  g697(.A(new_n871), .B1(new_n873), .B2(new_n883), .ZN(new_n884));
  OAI211_X1 g698(.A(new_n869), .B(new_n870), .C1(new_n884), .C2(KEYINPUT53), .ZN(new_n885));
  NOR3_X1   g699(.A1(new_n842), .A2(new_n853), .A3(new_n872), .ZN(new_n886));
  AOI21_X1  g700(.A(KEYINPUT109), .B1(new_n878), .B2(new_n882), .ZN(new_n887));
  OAI21_X1  g701(.A(new_n854), .B1(new_n886), .B2(new_n887), .ZN(new_n888));
  AND3_X1   g702(.A1(new_n859), .A2(new_n864), .A3(new_n867), .ZN(new_n889));
  AOI21_X1  g703(.A(new_n867), .B1(new_n859), .B2(new_n864), .ZN(new_n890));
  NOR2_X1   g704(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  INV_X1    g705(.A(new_n891), .ZN(new_n892));
  OAI22_X1  g706(.A1(new_n888), .A2(new_n892), .B1(new_n884), .B2(new_n854), .ZN(new_n893));
  OAI21_X1  g707(.A(new_n885), .B1(new_n893), .B2(new_n870), .ZN(new_n894));
  OAI22_X1  g708(.A1(new_n827), .A2(new_n894), .B1(G952), .B2(G953), .ZN(new_n895));
  XNOR2_X1  g709(.A(new_n804), .B(KEYINPUT49), .ZN(new_n896));
  NAND3_X1  g710(.A1(new_n369), .A2(new_n439), .A3(new_n437), .ZN(new_n897));
  OR4_X1    g711(.A1(new_n698), .A2(new_n896), .A3(new_n773), .A4(new_n897), .ZN(new_n898));
  OAI21_X1  g712(.A(new_n895), .B1(new_n692), .B2(new_n898), .ZN(G75));
  INV_X1    g713(.A(KEYINPUT118), .ZN(new_n900));
  OAI21_X1  g714(.A(new_n869), .B1(new_n884), .B2(KEYINPUT53), .ZN(new_n901));
  AND2_X1   g715(.A1(new_n901), .A2(G902), .ZN(new_n902));
  NAND2_X1  g716(.A1(new_n902), .A2(G210), .ZN(new_n903));
  NAND2_X1  g717(.A1(new_n459), .A2(new_n461), .ZN(new_n904));
  XOR2_X1   g718(.A(new_n904), .B(new_n468), .Z(new_n905));
  XNOR2_X1  g719(.A(KEYINPUT114), .B(KEYINPUT55), .ZN(new_n906));
  XNOR2_X1  g720(.A(new_n905), .B(new_n906), .ZN(new_n907));
  XOR2_X1   g721(.A(KEYINPUT115), .B(KEYINPUT56), .Z(new_n908));
  NOR2_X1   g722(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  NAND2_X1  g723(.A1(new_n903), .A2(new_n909), .ZN(new_n910));
  NOR2_X1   g724(.A1(new_n308), .A2(G952), .ZN(new_n911));
  XNOR2_X1  g725(.A(new_n911), .B(KEYINPUT116), .ZN(new_n912));
  XNOR2_X1  g726(.A(new_n912), .B(KEYINPUT117), .ZN(new_n913));
  NAND2_X1  g727(.A1(new_n910), .A2(new_n913), .ZN(new_n914));
  AOI21_X1  g728(.A(KEYINPUT56), .B1(new_n902), .B2(G210), .ZN(new_n915));
  INV_X1    g729(.A(new_n907), .ZN(new_n916));
  NOR2_X1   g730(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  OAI21_X1  g731(.A(new_n900), .B1(new_n914), .B2(new_n917), .ZN(new_n918));
  INV_X1    g732(.A(new_n913), .ZN(new_n919));
  AOI21_X1  g733(.A(new_n919), .B1(new_n903), .B2(new_n909), .ZN(new_n920));
  OAI211_X1 g734(.A(new_n920), .B(KEYINPUT118), .C1(new_n916), .C2(new_n915), .ZN(new_n921));
  NAND2_X1  g735(.A1(new_n918), .A2(new_n921), .ZN(G51));
  NAND2_X1  g736(.A1(new_n901), .A2(KEYINPUT54), .ZN(new_n923));
  NAND2_X1  g737(.A1(new_n923), .A2(new_n885), .ZN(new_n924));
  XNOR2_X1  g738(.A(new_n432), .B(KEYINPUT57), .ZN(new_n925));
  NAND2_X1  g739(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  OAI21_X1  g740(.A(new_n926), .B1(new_n426), .B2(new_n416), .ZN(new_n927));
  NAND2_X1  g741(.A1(new_n902), .A2(new_n766), .ZN(new_n928));
  AOI21_X1  g742(.A(new_n912), .B1(new_n927), .B2(new_n928), .ZN(G54));
  NAND4_X1  g743(.A1(new_n902), .A2(KEYINPUT58), .A3(G475), .A4(new_n537), .ZN(new_n930));
  INV_X1    g744(.A(KEYINPUT119), .ZN(new_n931));
  OR2_X1    g745(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  NAND2_X1  g746(.A1(new_n930), .A2(new_n931), .ZN(new_n933));
  NAND3_X1  g747(.A1(new_n902), .A2(KEYINPUT58), .A3(G475), .ZN(new_n934));
  INV_X1    g748(.A(new_n537), .ZN(new_n935));
  AOI21_X1  g749(.A(new_n912), .B1(new_n934), .B2(new_n935), .ZN(new_n936));
  AND3_X1   g750(.A1(new_n932), .A2(new_n933), .A3(new_n936), .ZN(G60));
  NAND2_X1  g751(.A1(new_n615), .A2(new_n616), .ZN(new_n938));
  XOR2_X1   g752(.A(new_n938), .B(KEYINPUT120), .Z(new_n939));
  XNOR2_X1  g753(.A(new_n619), .B(KEYINPUT59), .ZN(new_n940));
  AND2_X1   g754(.A1(new_n939), .A2(new_n940), .ZN(new_n941));
  AOI21_X1  g755(.A(new_n919), .B1(new_n924), .B2(new_n941), .ZN(new_n942));
  INV_X1    g756(.A(new_n942), .ZN(new_n943));
  AOI21_X1  g757(.A(new_n939), .B1(new_n894), .B2(new_n940), .ZN(new_n944));
  OAI21_X1  g758(.A(KEYINPUT121), .B1(new_n943), .B2(new_n944), .ZN(new_n945));
  INV_X1    g759(.A(KEYINPUT121), .ZN(new_n946));
  AND2_X1   g760(.A1(new_n894), .A2(new_n940), .ZN(new_n947));
  OAI211_X1 g761(.A(new_n942), .B(new_n946), .C1(new_n947), .C2(new_n939), .ZN(new_n948));
  NAND2_X1  g762(.A1(new_n945), .A2(new_n948), .ZN(G63));
  XNOR2_X1  g763(.A(KEYINPUT122), .B(KEYINPUT60), .ZN(new_n950));
  NOR2_X1   g764(.A1(new_n558), .A2(new_n357), .ZN(new_n951));
  XNOR2_X1  g765(.A(new_n950), .B(new_n951), .ZN(new_n952));
  AND3_X1   g766(.A1(new_n901), .A2(KEYINPUT123), .A3(new_n952), .ZN(new_n953));
  AOI21_X1  g767(.A(KEYINPUT123), .B1(new_n901), .B2(new_n952), .ZN(new_n954));
  OAI21_X1  g768(.A(new_n655), .B1(new_n953), .B2(new_n954), .ZN(new_n955));
  INV_X1    g769(.A(KEYINPUT123), .ZN(new_n956));
  OAI21_X1  g770(.A(new_n865), .B1(new_n886), .B2(new_n887), .ZN(new_n957));
  AOI22_X1  g771(.A1(new_n957), .A2(new_n854), .B1(new_n891), .B2(new_n855), .ZN(new_n958));
  INV_X1    g772(.A(new_n952), .ZN(new_n959));
  OAI21_X1  g773(.A(new_n956), .B1(new_n958), .B2(new_n959), .ZN(new_n960));
  NAND3_X1  g774(.A1(new_n901), .A2(KEYINPUT123), .A3(new_n952), .ZN(new_n961));
  NAND3_X1  g775(.A1(new_n960), .A2(new_n354), .A3(new_n961), .ZN(new_n962));
  AND3_X1   g776(.A1(new_n955), .A2(new_n962), .A3(new_n913), .ZN(new_n963));
  INV_X1    g777(.A(KEYINPUT61), .ZN(new_n964));
  INV_X1    g778(.A(new_n655), .ZN(new_n965));
  AOI21_X1  g779(.A(new_n965), .B1(new_n960), .B2(new_n961), .ZN(new_n966));
  INV_X1    g780(.A(KEYINPUT124), .ZN(new_n967));
  OAI21_X1  g781(.A(new_n964), .B1(new_n966), .B2(new_n967), .ZN(new_n968));
  NAND2_X1  g782(.A1(new_n963), .A2(new_n968), .ZN(new_n969));
  AOI21_X1  g783(.A(KEYINPUT61), .B1(new_n955), .B2(KEYINPUT124), .ZN(new_n970));
  NAND3_X1  g784(.A1(new_n955), .A2(new_n962), .A3(new_n913), .ZN(new_n971));
  NAND2_X1  g785(.A1(new_n970), .A2(new_n971), .ZN(new_n972));
  NAND2_X1  g786(.A1(new_n969), .A2(new_n972), .ZN(G66));
  OAI21_X1  g787(.A(G953), .B1(new_n464), .B2(new_n554), .ZN(new_n974));
  OAI21_X1  g788(.A(new_n974), .B1(new_n882), .B2(G953), .ZN(new_n975));
  OAI21_X1  g789(.A(new_n904), .B1(G898), .B2(new_n308), .ZN(new_n976));
  XNOR2_X1  g790(.A(new_n975), .B(new_n976), .ZN(G69));
  INV_X1    g791(.A(new_n745), .ZN(new_n978));
  OR4_X1    g792(.A1(new_n978), .A2(new_n771), .A3(new_n679), .A4(new_n731), .ZN(new_n979));
  AND3_X1   g793(.A1(new_n979), .A2(new_n790), .A3(new_n761), .ZN(new_n980));
  AND2_X1   g794(.A1(new_n856), .A2(new_n705), .ZN(new_n981));
  AND2_X1   g795(.A1(new_n782), .A2(new_n756), .ZN(new_n982));
  NAND3_X1  g796(.A1(new_n980), .A2(new_n981), .A3(new_n982), .ZN(new_n983));
  INV_X1    g797(.A(KEYINPUT126), .ZN(new_n984));
  NAND2_X1  g798(.A1(new_n983), .A2(new_n984), .ZN(new_n985));
  NAND4_X1  g799(.A1(new_n980), .A2(KEYINPUT126), .A3(new_n981), .A4(new_n982), .ZN(new_n986));
  NAND3_X1  g800(.A1(new_n985), .A2(new_n308), .A3(new_n986), .ZN(new_n987));
  NAND2_X1  g801(.A1(new_n267), .A2(new_n268), .ZN(new_n988));
  XNOR2_X1  g802(.A(new_n988), .B(new_n533), .ZN(new_n989));
  AOI21_X1  g803(.A(new_n989), .B1(G900), .B2(G953), .ZN(new_n990));
  AND2_X1   g804(.A1(new_n987), .A2(new_n990), .ZN(new_n991));
  AOI21_X1  g805(.A(new_n308), .B1(G227), .B2(G900), .ZN(new_n992));
  INV_X1    g806(.A(KEYINPUT125), .ZN(new_n993));
  AOI21_X1  g807(.A(new_n626), .B1(new_n834), .B2(new_n837), .ZN(new_n994));
  OR4_X1    g808(.A1(new_n978), .A2(new_n681), .A3(new_n758), .A4(new_n994), .ZN(new_n995));
  NAND3_X1  g809(.A1(new_n790), .A2(new_n782), .A3(new_n995), .ZN(new_n996));
  NAND2_X1  g810(.A1(new_n701), .A2(new_n981), .ZN(new_n997));
  AOI21_X1  g811(.A(new_n996), .B1(KEYINPUT62), .B2(new_n997), .ZN(new_n998));
  OR2_X1    g812(.A1(new_n997), .A2(KEYINPUT62), .ZN(new_n999));
  AOI21_X1  g813(.A(G953), .B1(new_n998), .B2(new_n999), .ZN(new_n1000));
  INV_X1    g814(.A(new_n989), .ZN(new_n1001));
  OAI21_X1  g815(.A(new_n993), .B1(new_n1000), .B2(new_n1001), .ZN(new_n1002));
  OR3_X1    g816(.A1(new_n991), .A2(new_n992), .A3(new_n1002), .ZN(new_n1003));
  OAI21_X1  g817(.A(new_n992), .B1(new_n991), .B2(new_n1002), .ZN(new_n1004));
  NAND2_X1  g818(.A1(new_n1003), .A2(new_n1004), .ZN(G72));
  NAND3_X1  g819(.A1(new_n985), .A2(new_n882), .A3(new_n986), .ZN(new_n1006));
  NAND2_X1  g820(.A1(G472), .A2(G902), .ZN(new_n1007));
  XOR2_X1   g821(.A(new_n1007), .B(KEYINPUT63), .Z(new_n1008));
  AOI211_X1 g822(.A(new_n254), .B(new_n270), .C1(new_n1006), .C2(new_n1008), .ZN(new_n1009));
  NAND2_X1  g823(.A1(new_n270), .A2(new_n254), .ZN(new_n1010));
  NAND3_X1  g824(.A1(new_n998), .A2(new_n882), .A3(new_n999), .ZN(new_n1011));
  AOI21_X1  g825(.A(new_n1010), .B1(new_n1011), .B2(new_n1008), .ZN(new_n1012));
  INV_X1    g826(.A(KEYINPUT127), .ZN(new_n1013));
  NAND2_X1  g827(.A1(new_n292), .A2(new_n1013), .ZN(new_n1014));
  NAND2_X1  g828(.A1(new_n270), .A2(new_n271), .ZN(new_n1015));
  XNOR2_X1  g829(.A(new_n1014), .B(new_n1015), .ZN(new_n1016));
  NAND2_X1  g830(.A1(new_n1016), .A2(new_n1008), .ZN(new_n1017));
  NOR2_X1   g831(.A1(new_n893), .A2(new_n1017), .ZN(new_n1018));
  NOR4_X1   g832(.A1(new_n1009), .A2(new_n1012), .A3(new_n912), .A4(new_n1018), .ZN(G57));
endmodule


