

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n523, n524, n525, n526,
         n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537,
         n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
         n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559,
         n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570,
         n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581,
         n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592,
         n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603,
         n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614,
         n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625,
         n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636,
         n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647,
         n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658,
         n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669,
         n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680,
         n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691,
         n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702,
         n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713,
         n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724,
         n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735,
         n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746,
         n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757,
         n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768,
         n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779,
         n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790,
         n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801,
         n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812,
         n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823,
         n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834,
         n835, n836, n837, n838, n839, n840, n841, n842, n843, n844, n845,
         n846, n847, n848, n849, n850, n851, n852, n853, n854, n855, n856,
         n857, n858, n859, n860, n861, n862, n863, n864, n865, n866, n867,
         n868, n869, n870, n871, n872, n873, n874, n875, n876, n877, n878,
         n879, n880, n881, n882, n883, n884, n885, n886, n887, n888, n889,
         n890, n891, n892, n893, n894, n895, n896, n897, n898, n899, n900,
         n901, n902, n903, n904, n905, n906, n907, n908, n909, n910, n911,
         n912, n913, n914, n915, n916, n917, n918, n919, n920, n921, n922,
         n923, n924, n925, n926, n927, n928, n929, n930, n931, n932, n933,
         n934, n935, n936, n937, n938, n939, n940, n941, n942, n943, n944,
         n945, n946, n947, n948, n949, n950, n951, n952, n953, n954, n955,
         n956, n957, n958, n959, n960, n961, n962, n963, n964, n965, n966,
         n967, n968, n969, n970, n971, n972, n973, n974, n975, n976, n977,
         n978, n979, n980, n981, n982, n983, n984, n985, n986, n987, n988,
         n989, n990, n991, n992, n993, n994, n995, n996, n997, n998, n999,
         n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009,
         n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019,
         n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029,
         n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039,
         n1040;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NAND2_X1 U558 ( .A1(n583), .A2(n582), .ZN(n1000) );
  NOR2_X1 U559 ( .A1(n640), .A2(n530), .ZN(n649) );
  XNOR2_X1 U560 ( .A(KEYINPUT64), .B(n524), .ZN(n654) );
  XNOR2_X2 U561 ( .A(n759), .B(KEYINPUT100), .ZN(n778) );
  XNOR2_X1 U562 ( .A(n550), .B(n549), .ZN(n551) );
  BUF_X1 U563 ( .A(n615), .Z(n616) );
  NOR2_X2 U564 ( .A1(G2104), .A2(n547), .ZN(n902) );
  NOR2_X1 U565 ( .A1(G168), .A2(n729), .ZN(n731) );
  NAND2_X1 U566 ( .A1(n748), .A2(n747), .ZN(n750) );
  INV_X1 U567 ( .A(KEYINPUT102), .ZN(n763) );
  INV_X1 U568 ( .A(KEYINPUT23), .ZN(n549) );
  NOR2_X1 U569 ( .A1(n694), .A2(n1000), .ZN(n702) );
  XNOR2_X1 U570 ( .A(n735), .B(KEYINPUT31), .ZN(n737) );
  AND2_X1 U571 ( .A1(n769), .A2(n768), .ZN(n770) );
  NOR2_X1 U572 ( .A1(n556), .A2(n555), .ZN(n687) );
  INV_X1 U573 ( .A(n724), .ZN(n695) );
  INV_X1 U574 ( .A(KEYINPUT98), .ZN(n730) );
  INV_X1 U575 ( .A(KEYINPUT29), .ZN(n717) );
  INV_X1 U576 ( .A(KEYINPUT99), .ZN(n736) );
  BUF_X1 U577 ( .A(n724), .Z(n741) );
  INV_X1 U578 ( .A(KEYINPUT32), .ZN(n749) );
  INV_X1 U579 ( .A(KEYINPUT104), .ZN(n767) );
  NOR2_X1 U580 ( .A1(n986), .A2(n767), .ZN(n768) );
  NAND2_X1 U581 ( .A1(n688), .A2(n805), .ZN(n724) );
  NOR2_X1 U582 ( .A1(n580), .A2(n579), .ZN(n581) );
  NOR2_X1 U583 ( .A1(G651), .A2(G543), .ZN(n648) );
  XOR2_X1 U584 ( .A(G543), .B(KEYINPUT0), .Z(n640) );
  XNOR2_X1 U585 ( .A(KEYINPUT69), .B(KEYINPUT6), .ZN(n527) );
  XNOR2_X1 U586 ( .A(n528), .B(n527), .ZN(n536) );
  INV_X1 U587 ( .A(G651), .ZN(n530) );
  NOR2_X1 U588 ( .A1(G543), .A2(n530), .ZN(n523) );
  XOR2_X2 U589 ( .A(KEYINPUT1), .B(n523), .Z(n647) );
  NAND2_X1 U590 ( .A1(G63), .A2(n647), .ZN(n526) );
  NOR2_X1 U591 ( .A1(G651), .A2(n640), .ZN(n524) );
  NAND2_X1 U592 ( .A1(G51), .A2(n654), .ZN(n525) );
  NAND2_X1 U593 ( .A1(n526), .A2(n525), .ZN(n528) );
  XNOR2_X1 U594 ( .A(KEYINPUT68), .B(KEYINPUT5), .ZN(n534) );
  NAND2_X1 U595 ( .A1(n648), .A2(G89), .ZN(n529) );
  XNOR2_X1 U596 ( .A(n529), .B(KEYINPUT4), .ZN(n532) );
  NAND2_X1 U597 ( .A1(G76), .A2(n649), .ZN(n531) );
  NAND2_X1 U598 ( .A1(n532), .A2(n531), .ZN(n533) );
  XNOR2_X1 U599 ( .A(n534), .B(n533), .ZN(n535) );
  NAND2_X1 U600 ( .A1(n536), .A2(n535), .ZN(n537) );
  XNOR2_X1 U601 ( .A(KEYINPUT7), .B(n537), .ZN(G168) );
  INV_X2 U602 ( .A(G2105), .ZN(n547) );
  AND2_X1 U603 ( .A1(n547), .A2(G2104), .ZN(n905) );
  NAND2_X1 U604 ( .A1(G102), .A2(n905), .ZN(n541) );
  XNOR2_X1 U605 ( .A(KEYINPUT65), .B(KEYINPUT17), .ZN(n539) );
  NOR2_X1 U606 ( .A1(G2104), .A2(G2105), .ZN(n538) );
  XNOR2_X1 U607 ( .A(n539), .B(n538), .ZN(n615) );
  NAND2_X1 U608 ( .A1(G138), .A2(n615), .ZN(n540) );
  NAND2_X1 U609 ( .A1(n541), .A2(n540), .ZN(n546) );
  INV_X1 U610 ( .A(G2104), .ZN(n542) );
  NOR2_X2 U611 ( .A1(n542), .A2(n547), .ZN(n901) );
  NAND2_X1 U612 ( .A1(G114), .A2(n901), .ZN(n544) );
  NAND2_X1 U613 ( .A1(G126), .A2(n902), .ZN(n543) );
  NAND2_X1 U614 ( .A1(n544), .A2(n543), .ZN(n545) );
  NOR2_X1 U615 ( .A1(n546), .A2(n545), .ZN(G164) );
  AND2_X1 U616 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U617 ( .A(G132), .ZN(G219) );
  INV_X1 U618 ( .A(G82), .ZN(G220) );
  INV_X1 U619 ( .A(G120), .ZN(G236) );
  INV_X1 U620 ( .A(G69), .ZN(G235) );
  INV_X1 U621 ( .A(G108), .ZN(G238) );
  NAND2_X1 U622 ( .A1(n901), .A2(G113), .ZN(n552) );
  AND2_X1 U623 ( .A1(n547), .A2(G101), .ZN(n548) );
  NAND2_X1 U624 ( .A1(n548), .A2(G2104), .ZN(n550) );
  NAND2_X1 U625 ( .A1(n552), .A2(n551), .ZN(n556) );
  NAND2_X1 U626 ( .A1(G125), .A2(n902), .ZN(n554) );
  NAND2_X1 U627 ( .A1(G137), .A2(n615), .ZN(n553) );
  NAND2_X1 U628 ( .A1(n554), .A2(n553), .ZN(n555) );
  BUF_X1 U629 ( .A(n687), .Z(G160) );
  NAND2_X1 U630 ( .A1(G64), .A2(n647), .ZN(n558) );
  NAND2_X1 U631 ( .A1(G52), .A2(n654), .ZN(n557) );
  NAND2_X1 U632 ( .A1(n558), .A2(n557), .ZN(n563) );
  NAND2_X1 U633 ( .A1(G90), .A2(n648), .ZN(n560) );
  NAND2_X1 U634 ( .A1(G77), .A2(n649), .ZN(n559) );
  NAND2_X1 U635 ( .A1(n560), .A2(n559), .ZN(n561) );
  XOR2_X1 U636 ( .A(KEYINPUT9), .B(n561), .Z(n562) );
  NOR2_X1 U637 ( .A1(n563), .A2(n562), .ZN(G171) );
  NAND2_X1 U638 ( .A1(G75), .A2(n649), .ZN(n565) );
  NAND2_X1 U639 ( .A1(G50), .A2(n654), .ZN(n564) );
  NAND2_X1 U640 ( .A1(n565), .A2(n564), .ZN(n571) );
  NAND2_X1 U641 ( .A1(G62), .A2(n647), .ZN(n566) );
  XNOR2_X1 U642 ( .A(n566), .B(KEYINPUT76), .ZN(n569) );
  NAND2_X1 U643 ( .A1(G88), .A2(n648), .ZN(n567) );
  XOR2_X1 U644 ( .A(KEYINPUT77), .B(n567), .Z(n568) );
  NAND2_X1 U645 ( .A1(n569), .A2(n568), .ZN(n570) );
  NOR2_X1 U646 ( .A1(n571), .A2(n570), .ZN(G166) );
  XOR2_X1 U647 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U648 ( .A1(G7), .A2(G661), .ZN(n572) );
  XNOR2_X1 U649 ( .A(n572), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U650 ( .A(G223), .ZN(n844) );
  NAND2_X1 U651 ( .A1(n844), .A2(G567), .ZN(n573) );
  XOR2_X1 U652 ( .A(KEYINPUT11), .B(n573), .Z(G234) );
  NAND2_X1 U653 ( .A1(n647), .A2(G56), .ZN(n574) );
  XOR2_X1 U654 ( .A(KEYINPUT14), .B(n574), .Z(n580) );
  NAND2_X1 U655 ( .A1(n648), .A2(G81), .ZN(n575) );
  XNOR2_X1 U656 ( .A(n575), .B(KEYINPUT12), .ZN(n577) );
  NAND2_X1 U657 ( .A1(G68), .A2(n649), .ZN(n576) );
  NAND2_X1 U658 ( .A1(n577), .A2(n576), .ZN(n578) );
  XOR2_X1 U659 ( .A(KEYINPUT13), .B(n578), .Z(n579) );
  XNOR2_X1 U660 ( .A(n581), .B(KEYINPUT66), .ZN(n583) );
  NAND2_X1 U661 ( .A1(G43), .A2(n654), .ZN(n582) );
  INV_X1 U662 ( .A(n1000), .ZN(n584) );
  XOR2_X1 U663 ( .A(G860), .B(KEYINPUT67), .Z(n604) );
  NAND2_X1 U664 ( .A1(n584), .A2(n604), .ZN(G153) );
  INV_X1 U665 ( .A(G171), .ZN(G301) );
  NAND2_X1 U666 ( .A1(G868), .A2(G301), .ZN(n593) );
  NAND2_X1 U667 ( .A1(G92), .A2(n648), .ZN(n586) );
  NAND2_X1 U668 ( .A1(G79), .A2(n649), .ZN(n585) );
  NAND2_X1 U669 ( .A1(n586), .A2(n585), .ZN(n590) );
  NAND2_X1 U670 ( .A1(G66), .A2(n647), .ZN(n588) );
  NAND2_X1 U671 ( .A1(G54), .A2(n654), .ZN(n587) );
  NAND2_X1 U672 ( .A1(n588), .A2(n587), .ZN(n589) );
  NOR2_X1 U673 ( .A1(n590), .A2(n589), .ZN(n591) );
  XOR2_X1 U674 ( .A(KEYINPUT15), .B(n591), .Z(n701) );
  INV_X1 U675 ( .A(n701), .ZN(n995) );
  INV_X1 U676 ( .A(G868), .ZN(n665) );
  NAND2_X1 U677 ( .A1(n995), .A2(n665), .ZN(n592) );
  NAND2_X1 U678 ( .A1(n593), .A2(n592), .ZN(G284) );
  NAND2_X1 U679 ( .A1(G65), .A2(n647), .ZN(n595) );
  NAND2_X1 U680 ( .A1(G53), .A2(n654), .ZN(n594) );
  NAND2_X1 U681 ( .A1(n595), .A2(n594), .ZN(n599) );
  NAND2_X1 U682 ( .A1(G91), .A2(n648), .ZN(n597) );
  NAND2_X1 U683 ( .A1(G78), .A2(n649), .ZN(n596) );
  NAND2_X1 U684 ( .A1(n597), .A2(n596), .ZN(n598) );
  NOR2_X1 U685 ( .A1(n599), .A2(n598), .ZN(n711) );
  INV_X1 U686 ( .A(n711), .ZN(G299) );
  NOR2_X1 U687 ( .A1(G868), .A2(G299), .ZN(n600) );
  XNOR2_X1 U688 ( .A(n600), .B(KEYINPUT70), .ZN(n602) );
  NOR2_X1 U689 ( .A1(n665), .A2(G286), .ZN(n601) );
  NOR2_X1 U690 ( .A1(n602), .A2(n601), .ZN(G297) );
  INV_X1 U691 ( .A(G559), .ZN(n603) );
  NOR2_X1 U692 ( .A1(n604), .A2(n603), .ZN(n605) );
  NOR2_X1 U693 ( .A1(n995), .A2(n605), .ZN(n606) );
  XOR2_X1 U694 ( .A(KEYINPUT16), .B(n606), .Z(G148) );
  NOR2_X1 U695 ( .A1(n995), .A2(n665), .ZN(n607) );
  XNOR2_X1 U696 ( .A(n607), .B(KEYINPUT71), .ZN(n608) );
  NOR2_X1 U697 ( .A1(G559), .A2(n608), .ZN(n610) );
  NOR2_X1 U698 ( .A1(G868), .A2(n1000), .ZN(n609) );
  NOR2_X1 U699 ( .A1(n610), .A2(n609), .ZN(G282) );
  NAND2_X1 U700 ( .A1(G123), .A2(n902), .ZN(n611) );
  XNOR2_X1 U701 ( .A(n611), .B(KEYINPUT18), .ZN(n614) );
  NAND2_X1 U702 ( .A1(G111), .A2(n901), .ZN(n612) );
  XNOR2_X1 U703 ( .A(n612), .B(KEYINPUT72), .ZN(n613) );
  NAND2_X1 U704 ( .A1(n614), .A2(n613), .ZN(n620) );
  NAND2_X1 U705 ( .A1(G99), .A2(n905), .ZN(n618) );
  NAND2_X1 U706 ( .A1(G135), .A2(n616), .ZN(n617) );
  NAND2_X1 U707 ( .A1(n618), .A2(n617), .ZN(n619) );
  NOR2_X1 U708 ( .A1(n620), .A2(n619), .ZN(n941) );
  XNOR2_X1 U709 ( .A(G2096), .B(n941), .ZN(n622) );
  INV_X1 U710 ( .A(G2100), .ZN(n621) );
  NAND2_X1 U711 ( .A1(n622), .A2(n621), .ZN(G156) );
  NAND2_X1 U712 ( .A1(G67), .A2(n647), .ZN(n624) );
  NAND2_X1 U713 ( .A1(G55), .A2(n654), .ZN(n623) );
  NAND2_X1 U714 ( .A1(n624), .A2(n623), .ZN(n628) );
  NAND2_X1 U715 ( .A1(G93), .A2(n648), .ZN(n626) );
  NAND2_X1 U716 ( .A1(G80), .A2(n649), .ZN(n625) );
  NAND2_X1 U717 ( .A1(n626), .A2(n625), .ZN(n627) );
  NOR2_X1 U718 ( .A1(n628), .A2(n627), .ZN(n666) );
  NAND2_X1 U719 ( .A1(n701), .A2(G559), .ZN(n663) );
  XNOR2_X1 U720 ( .A(n1000), .B(n663), .ZN(n629) );
  NOR2_X1 U721 ( .A1(G860), .A2(n629), .ZN(n630) );
  XOR2_X1 U722 ( .A(KEYINPUT73), .B(n630), .Z(n631) );
  XNOR2_X1 U723 ( .A(n666), .B(n631), .ZN(G145) );
  NAND2_X1 U724 ( .A1(G73), .A2(n649), .ZN(n632) );
  XOR2_X1 U725 ( .A(KEYINPUT2), .B(n632), .Z(n637) );
  NAND2_X1 U726 ( .A1(G86), .A2(n648), .ZN(n634) );
  NAND2_X1 U727 ( .A1(G61), .A2(n647), .ZN(n633) );
  NAND2_X1 U728 ( .A1(n634), .A2(n633), .ZN(n635) );
  XOR2_X1 U729 ( .A(KEYINPUT75), .B(n635), .Z(n636) );
  NOR2_X1 U730 ( .A1(n637), .A2(n636), .ZN(n639) );
  NAND2_X1 U731 ( .A1(G48), .A2(n654), .ZN(n638) );
  NAND2_X1 U732 ( .A1(n639), .A2(n638), .ZN(G305) );
  NAND2_X1 U733 ( .A1(G87), .A2(n640), .ZN(n641) );
  XNOR2_X1 U734 ( .A(n641), .B(KEYINPUT74), .ZN(n646) );
  NAND2_X1 U735 ( .A1(G651), .A2(G74), .ZN(n643) );
  NAND2_X1 U736 ( .A1(G49), .A2(n654), .ZN(n642) );
  NAND2_X1 U737 ( .A1(n643), .A2(n642), .ZN(n644) );
  NOR2_X1 U738 ( .A1(n647), .A2(n644), .ZN(n645) );
  NAND2_X1 U739 ( .A1(n646), .A2(n645), .ZN(G288) );
  AND2_X1 U740 ( .A1(n647), .A2(G60), .ZN(n653) );
  NAND2_X1 U741 ( .A1(G85), .A2(n648), .ZN(n651) );
  NAND2_X1 U742 ( .A1(G72), .A2(n649), .ZN(n650) );
  NAND2_X1 U743 ( .A1(n651), .A2(n650), .ZN(n652) );
  NOR2_X1 U744 ( .A1(n653), .A2(n652), .ZN(n656) );
  NAND2_X1 U745 ( .A1(G47), .A2(n654), .ZN(n655) );
  NAND2_X1 U746 ( .A1(n656), .A2(n655), .ZN(G290) );
  XNOR2_X1 U747 ( .A(G166), .B(n666), .ZN(n659) );
  XNOR2_X1 U748 ( .A(KEYINPUT19), .B(G305), .ZN(n657) );
  XNOR2_X1 U749 ( .A(n657), .B(G288), .ZN(n658) );
  XNOR2_X1 U750 ( .A(n659), .B(n658), .ZN(n660) );
  XNOR2_X1 U751 ( .A(n711), .B(n660), .ZN(n661) );
  XNOR2_X1 U752 ( .A(n661), .B(G290), .ZN(n662) );
  XNOR2_X1 U753 ( .A(n1000), .B(n662), .ZN(n916) );
  XOR2_X1 U754 ( .A(n916), .B(n663), .Z(n664) );
  NOR2_X1 U755 ( .A1(n665), .A2(n664), .ZN(n668) );
  NOR2_X1 U756 ( .A1(G868), .A2(n666), .ZN(n667) );
  NOR2_X1 U757 ( .A1(n668), .A2(n667), .ZN(n669) );
  XOR2_X1 U758 ( .A(KEYINPUT78), .B(n669), .Z(G295) );
  NAND2_X1 U759 ( .A1(G2084), .A2(G2078), .ZN(n670) );
  XNOR2_X1 U760 ( .A(n670), .B(KEYINPUT20), .ZN(n671) );
  XNOR2_X1 U761 ( .A(KEYINPUT79), .B(n671), .ZN(n672) );
  NAND2_X1 U762 ( .A1(n672), .A2(G2090), .ZN(n673) );
  XNOR2_X1 U763 ( .A(n673), .B(KEYINPUT80), .ZN(n674) );
  XNOR2_X1 U764 ( .A(KEYINPUT21), .B(n674), .ZN(n675) );
  NAND2_X1 U765 ( .A1(n675), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U766 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U767 ( .A1(G235), .A2(G236), .ZN(n676) );
  XOR2_X1 U768 ( .A(KEYINPUT82), .B(n676), .Z(n677) );
  NOR2_X1 U769 ( .A1(G238), .A2(n677), .ZN(n678) );
  NAND2_X1 U770 ( .A1(G57), .A2(n678), .ZN(n849) );
  NAND2_X1 U771 ( .A1(n849), .A2(G567), .ZN(n684) );
  NOR2_X1 U772 ( .A1(G220), .A2(G219), .ZN(n679) );
  XOR2_X1 U773 ( .A(KEYINPUT22), .B(n679), .Z(n680) );
  NOR2_X1 U774 ( .A1(G218), .A2(n680), .ZN(n681) );
  XOR2_X1 U775 ( .A(KEYINPUT81), .B(n681), .Z(n682) );
  NAND2_X1 U776 ( .A1(G96), .A2(n682), .ZN(n850) );
  NAND2_X1 U777 ( .A1(n850), .A2(G2106), .ZN(n683) );
  NAND2_X1 U778 ( .A1(n684), .A2(n683), .ZN(n851) );
  NAND2_X1 U779 ( .A1(G483), .A2(G661), .ZN(n685) );
  NOR2_X1 U780 ( .A1(n851), .A2(n685), .ZN(n686) );
  XOR2_X1 U781 ( .A(KEYINPUT83), .B(n686), .Z(n847) );
  NAND2_X1 U782 ( .A1(n847), .A2(G36), .ZN(G176) );
  INV_X1 U783 ( .A(G166), .ZN(G303) );
  INV_X1 U784 ( .A(KEYINPUT95), .ZN(n693) );
  NAND2_X1 U785 ( .A1(n687), .A2(G40), .ZN(n804) );
  XNOR2_X1 U786 ( .A(KEYINPUT91), .B(n804), .ZN(n688) );
  NOR2_X1 U787 ( .A1(G164), .A2(G1384), .ZN(n805) );
  NAND2_X1 U788 ( .A1(G1996), .A2(n695), .ZN(n689) );
  XNOR2_X1 U789 ( .A(n689), .B(KEYINPUT26), .ZN(n691) );
  NAND2_X1 U790 ( .A1(G1341), .A2(n741), .ZN(n690) );
  NAND2_X1 U791 ( .A1(n691), .A2(n690), .ZN(n692) );
  XNOR2_X1 U792 ( .A(n693), .B(n692), .ZN(n694) );
  NAND2_X1 U793 ( .A1(n702), .A2(n701), .ZN(n700) );
  BUF_X1 U794 ( .A(n695), .Z(n696) );
  NOR2_X1 U795 ( .A1(n696), .A2(G1348), .ZN(n698) );
  NOR2_X1 U796 ( .A1(G2067), .A2(n741), .ZN(n697) );
  NOR2_X1 U797 ( .A1(n698), .A2(n697), .ZN(n699) );
  NAND2_X1 U798 ( .A1(n700), .A2(n699), .ZN(n704) );
  OR2_X1 U799 ( .A1(n702), .A2(n701), .ZN(n703) );
  NAND2_X1 U800 ( .A1(n704), .A2(n703), .ZN(n705) );
  XNOR2_X1 U801 ( .A(n705), .B(KEYINPUT96), .ZN(n710) );
  NAND2_X1 U802 ( .A1(n696), .A2(G2072), .ZN(n706) );
  XNOR2_X1 U803 ( .A(n706), .B(KEYINPUT27), .ZN(n708) );
  INV_X1 U804 ( .A(G1956), .ZN(n961) );
  NOR2_X1 U805 ( .A1(n961), .A2(n696), .ZN(n707) );
  NOR2_X1 U806 ( .A1(n708), .A2(n707), .ZN(n712) );
  NAND2_X1 U807 ( .A1(n712), .A2(n711), .ZN(n709) );
  NAND2_X1 U808 ( .A1(n710), .A2(n709), .ZN(n716) );
  NOR2_X1 U809 ( .A1(n712), .A2(n711), .ZN(n714) );
  XOR2_X1 U810 ( .A(KEYINPUT28), .B(KEYINPUT94), .Z(n713) );
  XNOR2_X1 U811 ( .A(n714), .B(n713), .ZN(n715) );
  NAND2_X1 U812 ( .A1(n716), .A2(n715), .ZN(n718) );
  XNOR2_X1 U813 ( .A(n718), .B(n717), .ZN(n723) );
  NOR2_X1 U814 ( .A1(n696), .A2(G1961), .ZN(n719) );
  XOR2_X1 U815 ( .A(KEYINPUT93), .B(n719), .Z(n721) );
  XOR2_X1 U816 ( .A(G2078), .B(KEYINPUT25), .Z(n1023) );
  NOR2_X1 U817 ( .A1(n1023), .A2(n741), .ZN(n720) );
  NOR2_X1 U818 ( .A1(n721), .A2(n720), .ZN(n732) );
  OR2_X1 U819 ( .A1(n732), .A2(G301), .ZN(n722) );
  NAND2_X1 U820 ( .A1(n723), .A2(n722), .ZN(n739) );
  NOR2_X1 U821 ( .A1(G2084), .A2(n741), .ZN(n751) );
  NAND2_X2 U822 ( .A1(G8), .A2(n724), .ZN(n783) );
  NOR2_X1 U823 ( .A1(n783), .A2(G1966), .ZN(n725) );
  XNOR2_X1 U824 ( .A(n725), .B(KEYINPUT92), .ZN(n753) );
  NOR2_X1 U825 ( .A1(n751), .A2(n753), .ZN(n726) );
  NAND2_X1 U826 ( .A1(n726), .A2(G8), .ZN(n728) );
  XOR2_X1 U827 ( .A(KEYINPUT30), .B(KEYINPUT97), .Z(n727) );
  XNOR2_X1 U828 ( .A(n728), .B(n727), .ZN(n729) );
  XNOR2_X1 U829 ( .A(n731), .B(n730), .ZN(n734) );
  NAND2_X1 U830 ( .A1(G301), .A2(n732), .ZN(n733) );
  NAND2_X1 U831 ( .A1(n734), .A2(n733), .ZN(n735) );
  XNOR2_X1 U832 ( .A(n737), .B(n736), .ZN(n738) );
  NAND2_X1 U833 ( .A1(n739), .A2(n738), .ZN(n752) );
  AND2_X1 U834 ( .A1(G286), .A2(G8), .ZN(n740) );
  NAND2_X1 U835 ( .A1(n752), .A2(n740), .ZN(n748) );
  INV_X1 U836 ( .A(G8), .ZN(n746) );
  NOR2_X1 U837 ( .A1(G1971), .A2(n783), .ZN(n743) );
  NOR2_X1 U838 ( .A1(G2090), .A2(n741), .ZN(n742) );
  NOR2_X1 U839 ( .A1(n743), .A2(n742), .ZN(n744) );
  NAND2_X1 U840 ( .A1(n744), .A2(G303), .ZN(n745) );
  OR2_X1 U841 ( .A1(n746), .A2(n745), .ZN(n747) );
  XNOR2_X1 U842 ( .A(n750), .B(n749), .ZN(n758) );
  NAND2_X1 U843 ( .A1(G8), .A2(n751), .ZN(n756) );
  INV_X1 U844 ( .A(n752), .ZN(n754) );
  NOR2_X1 U845 ( .A1(n754), .A2(n753), .ZN(n755) );
  NAND2_X1 U846 ( .A1(n756), .A2(n755), .ZN(n757) );
  NAND2_X1 U847 ( .A1(n758), .A2(n757), .ZN(n759) );
  NOR2_X1 U848 ( .A1(G1976), .A2(G288), .ZN(n985) );
  NOR2_X1 U849 ( .A1(G1971), .A2(G303), .ZN(n760) );
  XOR2_X1 U850 ( .A(n760), .B(KEYINPUT101), .Z(n761) );
  NOR2_X1 U851 ( .A1(n985), .A2(n761), .ZN(n762) );
  NAND2_X1 U852 ( .A1(n778), .A2(n762), .ZN(n764) );
  XNOR2_X1 U853 ( .A(n764), .B(n763), .ZN(n765) );
  NOR2_X1 U854 ( .A1(n765), .A2(n783), .ZN(n769) );
  NAND2_X1 U855 ( .A1(G288), .A2(G1976), .ZN(n766) );
  XNOR2_X1 U856 ( .A(n766), .B(KEYINPUT103), .ZN(n986) );
  NOR2_X1 U857 ( .A1(KEYINPUT33), .A2(n770), .ZN(n774) );
  XNOR2_X1 U858 ( .A(n985), .B(KEYINPUT104), .ZN(n771) );
  NAND2_X1 U859 ( .A1(n771), .A2(KEYINPUT33), .ZN(n772) );
  NOR2_X1 U860 ( .A1(n783), .A2(n772), .ZN(n773) );
  NOR2_X1 U861 ( .A1(n774), .A2(n773), .ZN(n775) );
  XOR2_X1 U862 ( .A(G1981), .B(G305), .Z(n1003) );
  NAND2_X1 U863 ( .A1(n775), .A2(n1003), .ZN(n776) );
  XNOR2_X1 U864 ( .A(n776), .B(KEYINPUT105), .ZN(n832) );
  NOR2_X1 U865 ( .A1(G2090), .A2(G303), .ZN(n777) );
  NAND2_X1 U866 ( .A1(G8), .A2(n777), .ZN(n779) );
  NAND2_X1 U867 ( .A1(n779), .A2(n778), .ZN(n780) );
  AND2_X1 U868 ( .A1(n780), .A2(n783), .ZN(n785) );
  NOR2_X1 U869 ( .A1(G1981), .A2(G305), .ZN(n781) );
  XOR2_X1 U870 ( .A(n781), .B(KEYINPUT24), .Z(n782) );
  NOR2_X1 U871 ( .A1(n783), .A2(n782), .ZN(n784) );
  OR2_X1 U872 ( .A1(n785), .A2(n784), .ZN(n830) );
  NAND2_X1 U873 ( .A1(G129), .A2(n902), .ZN(n792) );
  NAND2_X1 U874 ( .A1(G141), .A2(n616), .ZN(n787) );
  NAND2_X1 U875 ( .A1(G117), .A2(n901), .ZN(n786) );
  NAND2_X1 U876 ( .A1(n787), .A2(n786), .ZN(n790) );
  NAND2_X1 U877 ( .A1(n905), .A2(G105), .ZN(n788) );
  XOR2_X1 U878 ( .A(KEYINPUT38), .B(n788), .Z(n789) );
  NOR2_X1 U879 ( .A1(n790), .A2(n789), .ZN(n791) );
  NAND2_X1 U880 ( .A1(n792), .A2(n791), .ZN(n793) );
  XNOR2_X1 U881 ( .A(n793), .B(KEYINPUT90), .ZN(n880) );
  NOR2_X1 U882 ( .A1(G1996), .A2(n880), .ZN(n936) );
  NAND2_X1 U883 ( .A1(G95), .A2(n905), .ZN(n795) );
  NAND2_X1 U884 ( .A1(G131), .A2(n616), .ZN(n794) );
  NAND2_X1 U885 ( .A1(n795), .A2(n794), .ZN(n796) );
  XOR2_X1 U886 ( .A(KEYINPUT88), .B(n796), .Z(n798) );
  NAND2_X1 U887 ( .A1(n901), .A2(G107), .ZN(n797) );
  NAND2_X1 U888 ( .A1(n798), .A2(n797), .ZN(n801) );
  NAND2_X1 U889 ( .A1(G119), .A2(n902), .ZN(n799) );
  XNOR2_X1 U890 ( .A(KEYINPUT87), .B(n799), .ZN(n800) );
  NOR2_X1 U891 ( .A1(n801), .A2(n800), .ZN(n884) );
  XNOR2_X1 U892 ( .A(KEYINPUT89), .B(G1991), .ZN(n1015) );
  NOR2_X1 U893 ( .A1(n884), .A2(n1015), .ZN(n803) );
  AND2_X1 U894 ( .A1(n880), .A2(G1996), .ZN(n802) );
  NOR2_X1 U895 ( .A1(n803), .A2(n802), .ZN(n943) );
  NOR2_X1 U896 ( .A1(n805), .A2(n804), .ZN(n836) );
  INV_X1 U897 ( .A(n836), .ZN(n806) );
  NOR2_X1 U898 ( .A1(n943), .A2(n806), .ZN(n833) );
  AND2_X1 U899 ( .A1(n1015), .A2(n884), .ZN(n945) );
  NOR2_X1 U900 ( .A1(G1986), .A2(G290), .ZN(n807) );
  NOR2_X1 U901 ( .A1(n945), .A2(n807), .ZN(n808) );
  XNOR2_X1 U902 ( .A(n808), .B(KEYINPUT106), .ZN(n809) );
  NOR2_X1 U903 ( .A1(n833), .A2(n809), .ZN(n810) );
  NOR2_X1 U904 ( .A1(n936), .A2(n810), .ZN(n811) );
  XNOR2_X1 U905 ( .A(n811), .B(KEYINPUT39), .ZN(n824) );
  XNOR2_X1 U906 ( .A(G2067), .B(KEYINPUT37), .ZN(n812) );
  XOR2_X1 U907 ( .A(n812), .B(KEYINPUT84), .Z(n825) );
  NAND2_X1 U908 ( .A1(G116), .A2(n901), .ZN(n814) );
  NAND2_X1 U909 ( .A1(G128), .A2(n902), .ZN(n813) );
  NAND2_X1 U910 ( .A1(n814), .A2(n813), .ZN(n815) );
  XOR2_X1 U911 ( .A(KEYINPUT35), .B(n815), .Z(n822) );
  XNOR2_X1 U912 ( .A(KEYINPUT85), .B(KEYINPUT86), .ZN(n816) );
  XNOR2_X1 U913 ( .A(n816), .B(KEYINPUT34), .ZN(n820) );
  NAND2_X1 U914 ( .A1(G104), .A2(n905), .ZN(n818) );
  NAND2_X1 U915 ( .A1(G140), .A2(n616), .ZN(n817) );
  NAND2_X1 U916 ( .A1(n818), .A2(n817), .ZN(n819) );
  XOR2_X1 U917 ( .A(n820), .B(n819), .Z(n821) );
  NOR2_X1 U918 ( .A1(n822), .A2(n821), .ZN(n823) );
  XOR2_X1 U919 ( .A(KEYINPUT36), .B(n823), .Z(n881) );
  AND2_X1 U920 ( .A1(n825), .A2(n881), .ZN(n939) );
  NAND2_X1 U921 ( .A1(n836), .A2(n939), .ZN(n835) );
  NAND2_X1 U922 ( .A1(n824), .A2(n835), .ZN(n827) );
  NOR2_X1 U923 ( .A1(n825), .A2(n881), .ZN(n826) );
  XNOR2_X1 U924 ( .A(n826), .B(KEYINPUT107), .ZN(n952) );
  NAND2_X1 U925 ( .A1(n827), .A2(n952), .ZN(n828) );
  NAND2_X1 U926 ( .A1(n828), .A2(n836), .ZN(n840) );
  INV_X1 U927 ( .A(n840), .ZN(n829) );
  OR2_X1 U928 ( .A1(n830), .A2(n829), .ZN(n831) );
  NOR2_X1 U929 ( .A1(n832), .A2(n831), .ZN(n842) );
  INV_X1 U930 ( .A(n833), .ZN(n834) );
  AND2_X1 U931 ( .A1(n835), .A2(n834), .ZN(n838) );
  XNOR2_X1 U932 ( .A(G1986), .B(G290), .ZN(n991) );
  NAND2_X1 U933 ( .A1(n991), .A2(n836), .ZN(n837) );
  NAND2_X1 U934 ( .A1(n838), .A2(n837), .ZN(n839) );
  AND2_X1 U935 ( .A1(n840), .A2(n839), .ZN(n841) );
  NOR2_X1 U936 ( .A1(n842), .A2(n841), .ZN(n843) );
  XNOR2_X1 U937 ( .A(n843), .B(KEYINPUT40), .ZN(G329) );
  NAND2_X1 U938 ( .A1(G2106), .A2(n844), .ZN(G217) );
  AND2_X1 U939 ( .A1(G15), .A2(G2), .ZN(n845) );
  NAND2_X1 U940 ( .A1(G661), .A2(n845), .ZN(G259) );
  NAND2_X1 U941 ( .A1(G3), .A2(G1), .ZN(n846) );
  NAND2_X1 U942 ( .A1(n847), .A2(n846), .ZN(n848) );
  XNOR2_X1 U943 ( .A(KEYINPUT108), .B(n848), .ZN(G188) );
  NOR2_X1 U944 ( .A1(n850), .A2(n849), .ZN(G325) );
  XNOR2_X1 U945 ( .A(KEYINPUT109), .B(G325), .ZN(G261) );
  INV_X1 U947 ( .A(G96), .ZN(G221) );
  INV_X1 U948 ( .A(n851), .ZN(G319) );
  XOR2_X1 U949 ( .A(KEYINPUT110), .B(KEYINPUT112), .Z(n853) );
  XNOR2_X1 U950 ( .A(G2678), .B(G2096), .ZN(n852) );
  XNOR2_X1 U951 ( .A(n853), .B(n852), .ZN(n854) );
  XOR2_X1 U952 ( .A(n854), .B(KEYINPUT111), .Z(n856) );
  XNOR2_X1 U953 ( .A(G2067), .B(G2072), .ZN(n855) );
  XNOR2_X1 U954 ( .A(n856), .B(n855), .ZN(n860) );
  XOR2_X1 U955 ( .A(G2100), .B(G2084), .Z(n858) );
  XNOR2_X1 U956 ( .A(G2090), .B(G2078), .ZN(n857) );
  XNOR2_X1 U957 ( .A(n858), .B(n857), .ZN(n859) );
  XOR2_X1 U958 ( .A(n860), .B(n859), .Z(n862) );
  XNOR2_X1 U959 ( .A(KEYINPUT42), .B(KEYINPUT43), .ZN(n861) );
  XNOR2_X1 U960 ( .A(n862), .B(n861), .ZN(G227) );
  XOR2_X1 U961 ( .A(G1981), .B(G1956), .Z(n864) );
  XNOR2_X1 U962 ( .A(G1991), .B(G1961), .ZN(n863) );
  XNOR2_X1 U963 ( .A(n864), .B(n863), .ZN(n868) );
  XOR2_X1 U964 ( .A(G1976), .B(G1971), .Z(n866) );
  XNOR2_X1 U965 ( .A(G1986), .B(G1966), .ZN(n865) );
  XNOR2_X1 U966 ( .A(n866), .B(n865), .ZN(n867) );
  XOR2_X1 U967 ( .A(n868), .B(n867), .Z(n870) );
  XNOR2_X1 U968 ( .A(KEYINPUT113), .B(G2474), .ZN(n869) );
  XNOR2_X1 U969 ( .A(n870), .B(n869), .ZN(n871) );
  XNOR2_X1 U970 ( .A(KEYINPUT41), .B(n871), .ZN(n872) );
  XOR2_X1 U971 ( .A(n872), .B(G1996), .Z(G229) );
  NAND2_X1 U972 ( .A1(G124), .A2(n902), .ZN(n873) );
  XNOR2_X1 U973 ( .A(n873), .B(KEYINPUT44), .ZN(n875) );
  NAND2_X1 U974 ( .A1(n901), .A2(G112), .ZN(n874) );
  NAND2_X1 U975 ( .A1(n875), .A2(n874), .ZN(n879) );
  NAND2_X1 U976 ( .A1(G100), .A2(n905), .ZN(n877) );
  NAND2_X1 U977 ( .A1(G136), .A2(n616), .ZN(n876) );
  NAND2_X1 U978 ( .A1(n877), .A2(n876), .ZN(n878) );
  NOR2_X1 U979 ( .A1(n879), .A2(n878), .ZN(G162) );
  XOR2_X1 U980 ( .A(G162), .B(n880), .Z(n883) );
  XNOR2_X1 U981 ( .A(G160), .B(n881), .ZN(n882) );
  XNOR2_X1 U982 ( .A(n883), .B(n882), .ZN(n887) );
  XNOR2_X1 U983 ( .A(G164), .B(n884), .ZN(n885) );
  XNOR2_X1 U984 ( .A(n885), .B(n941), .ZN(n886) );
  XOR2_X1 U985 ( .A(n887), .B(n886), .Z(n892) );
  XOR2_X1 U986 ( .A(KEYINPUT48), .B(KEYINPUT117), .Z(n889) );
  XNOR2_X1 U987 ( .A(KEYINPUT118), .B(KEYINPUT116), .ZN(n888) );
  XNOR2_X1 U988 ( .A(n889), .B(n888), .ZN(n890) );
  XNOR2_X1 U989 ( .A(KEYINPUT46), .B(n890), .ZN(n891) );
  XNOR2_X1 U990 ( .A(n892), .B(n891), .ZN(n914) );
  NAND2_X1 U991 ( .A1(G103), .A2(n905), .ZN(n894) );
  NAND2_X1 U992 ( .A1(G139), .A2(n616), .ZN(n893) );
  NAND2_X1 U993 ( .A1(n894), .A2(n893), .ZN(n900) );
  NAND2_X1 U994 ( .A1(n901), .A2(G115), .ZN(n895) );
  XOR2_X1 U995 ( .A(KEYINPUT115), .B(n895), .Z(n897) );
  NAND2_X1 U996 ( .A1(n902), .A2(G127), .ZN(n896) );
  NAND2_X1 U997 ( .A1(n897), .A2(n896), .ZN(n898) );
  XOR2_X1 U998 ( .A(KEYINPUT47), .B(n898), .Z(n899) );
  NOR2_X1 U999 ( .A1(n900), .A2(n899), .ZN(n948) );
  NAND2_X1 U1000 ( .A1(G118), .A2(n901), .ZN(n904) );
  NAND2_X1 U1001 ( .A1(G130), .A2(n902), .ZN(n903) );
  NAND2_X1 U1002 ( .A1(n904), .A2(n903), .ZN(n911) );
  NAND2_X1 U1003 ( .A1(G106), .A2(n905), .ZN(n907) );
  NAND2_X1 U1004 ( .A1(G142), .A2(n616), .ZN(n906) );
  NAND2_X1 U1005 ( .A1(n907), .A2(n906), .ZN(n908) );
  XOR2_X1 U1006 ( .A(KEYINPUT45), .B(n908), .Z(n909) );
  XNOR2_X1 U1007 ( .A(KEYINPUT114), .B(n909), .ZN(n910) );
  NOR2_X1 U1008 ( .A1(n911), .A2(n910), .ZN(n912) );
  XNOR2_X1 U1009 ( .A(n948), .B(n912), .ZN(n913) );
  XNOR2_X1 U1010 ( .A(n914), .B(n913), .ZN(n915) );
  NOR2_X1 U1011 ( .A1(G37), .A2(n915), .ZN(G395) );
  XNOR2_X1 U1012 ( .A(G286), .B(n995), .ZN(n917) );
  XNOR2_X1 U1013 ( .A(n917), .B(n916), .ZN(n918) );
  XNOR2_X1 U1014 ( .A(n918), .B(G171), .ZN(n919) );
  NOR2_X1 U1015 ( .A1(G37), .A2(n919), .ZN(G397) );
  XOR2_X1 U1016 ( .A(G2451), .B(G2430), .Z(n921) );
  XNOR2_X1 U1017 ( .A(G2438), .B(G2443), .ZN(n920) );
  XNOR2_X1 U1018 ( .A(n921), .B(n920), .ZN(n927) );
  XOR2_X1 U1019 ( .A(G2435), .B(G2454), .Z(n923) );
  XNOR2_X1 U1020 ( .A(G1341), .B(G1348), .ZN(n922) );
  XNOR2_X1 U1021 ( .A(n923), .B(n922), .ZN(n925) );
  XOR2_X1 U1022 ( .A(G2446), .B(G2427), .Z(n924) );
  XNOR2_X1 U1023 ( .A(n925), .B(n924), .ZN(n926) );
  XOR2_X1 U1024 ( .A(n927), .B(n926), .Z(n928) );
  NAND2_X1 U1025 ( .A1(G14), .A2(n928), .ZN(n934) );
  NAND2_X1 U1026 ( .A1(G319), .A2(n934), .ZN(n931) );
  NOR2_X1 U1027 ( .A1(G227), .A2(G229), .ZN(n929) );
  XNOR2_X1 U1028 ( .A(KEYINPUT49), .B(n929), .ZN(n930) );
  NOR2_X1 U1029 ( .A1(n931), .A2(n930), .ZN(n933) );
  NOR2_X1 U1030 ( .A1(G395), .A2(G397), .ZN(n932) );
  NAND2_X1 U1031 ( .A1(n933), .A2(n932), .ZN(G225) );
  INV_X1 U1032 ( .A(G225), .ZN(G308) );
  INV_X1 U1033 ( .A(G57), .ZN(G237) );
  INV_X1 U1034 ( .A(n934), .ZN(G401) );
  XOR2_X1 U1035 ( .A(G2090), .B(G162), .Z(n935) );
  NOR2_X1 U1036 ( .A1(n936), .A2(n935), .ZN(n937) );
  XNOR2_X1 U1037 ( .A(n937), .B(KEYINPUT51), .ZN(n938) );
  NOR2_X1 U1038 ( .A1(n939), .A2(n938), .ZN(n947) );
  XOR2_X1 U1039 ( .A(G2084), .B(G160), .Z(n940) );
  NOR2_X1 U1040 ( .A1(n941), .A2(n940), .ZN(n942) );
  NAND2_X1 U1041 ( .A1(n943), .A2(n942), .ZN(n944) );
  NOR2_X1 U1042 ( .A1(n945), .A2(n944), .ZN(n946) );
  NAND2_X1 U1043 ( .A1(n947), .A2(n946), .ZN(n955) );
  XOR2_X1 U1044 ( .A(G2072), .B(n948), .Z(n950) );
  XOR2_X1 U1045 ( .A(G164), .B(G2078), .Z(n949) );
  NOR2_X1 U1046 ( .A1(n950), .A2(n949), .ZN(n951) );
  XNOR2_X1 U1047 ( .A(n951), .B(KEYINPUT50), .ZN(n953) );
  NAND2_X1 U1048 ( .A1(n953), .A2(n952), .ZN(n954) );
  NOR2_X1 U1049 ( .A1(n955), .A2(n954), .ZN(n956) );
  XOR2_X1 U1050 ( .A(KEYINPUT52), .B(n956), .Z(n957) );
  NOR2_X1 U1051 ( .A1(KEYINPUT55), .A2(n957), .ZN(n958) );
  XNOR2_X1 U1052 ( .A(KEYINPUT119), .B(n958), .ZN(n959) );
  NAND2_X1 U1053 ( .A1(n959), .A2(G29), .ZN(n1014) );
  XNOR2_X1 U1054 ( .A(G21), .B(G1966), .ZN(n960) );
  XNOR2_X1 U1055 ( .A(n960), .B(KEYINPUT127), .ZN(n973) );
  XNOR2_X1 U1056 ( .A(G20), .B(n961), .ZN(n965) );
  XNOR2_X1 U1057 ( .A(G1341), .B(G19), .ZN(n963) );
  XNOR2_X1 U1058 ( .A(G1981), .B(G6), .ZN(n962) );
  NOR2_X1 U1059 ( .A1(n963), .A2(n962), .ZN(n964) );
  NAND2_X1 U1060 ( .A1(n965), .A2(n964), .ZN(n968) );
  XOR2_X1 U1061 ( .A(KEYINPUT59), .B(G1348), .Z(n966) );
  XNOR2_X1 U1062 ( .A(G4), .B(n966), .ZN(n967) );
  NOR2_X1 U1063 ( .A1(n968), .A2(n967), .ZN(n969) );
  XOR2_X1 U1064 ( .A(KEYINPUT60), .B(n969), .Z(n971) );
  XNOR2_X1 U1065 ( .A(G1961), .B(G5), .ZN(n970) );
  NOR2_X1 U1066 ( .A1(n971), .A2(n970), .ZN(n972) );
  NAND2_X1 U1067 ( .A1(n973), .A2(n972), .ZN(n980) );
  XNOR2_X1 U1068 ( .A(G1971), .B(G22), .ZN(n975) );
  XNOR2_X1 U1069 ( .A(G23), .B(G1976), .ZN(n974) );
  NOR2_X1 U1070 ( .A1(n975), .A2(n974), .ZN(n977) );
  XOR2_X1 U1071 ( .A(G1986), .B(G24), .Z(n976) );
  NAND2_X1 U1072 ( .A1(n977), .A2(n976), .ZN(n978) );
  XNOR2_X1 U1073 ( .A(KEYINPUT58), .B(n978), .ZN(n979) );
  NOR2_X1 U1074 ( .A1(n980), .A2(n979), .ZN(n981) );
  XNOR2_X1 U1075 ( .A(KEYINPUT61), .B(n981), .ZN(n983) );
  INV_X1 U1076 ( .A(G16), .ZN(n982) );
  NAND2_X1 U1077 ( .A1(n983), .A2(n982), .ZN(n984) );
  NAND2_X1 U1078 ( .A1(n984), .A2(G11), .ZN(n1012) );
  XNOR2_X1 U1079 ( .A(KEYINPUT56), .B(G16), .ZN(n1009) );
  XNOR2_X1 U1080 ( .A(G166), .B(G1971), .ZN(n988) );
  NOR2_X1 U1081 ( .A1(n986), .A2(n985), .ZN(n987) );
  NAND2_X1 U1082 ( .A1(n988), .A2(n987), .ZN(n989) );
  XOR2_X1 U1083 ( .A(KEYINPUT124), .B(n989), .Z(n993) );
  XNOR2_X1 U1084 ( .A(G1956), .B(G299), .ZN(n990) );
  NOR2_X1 U1085 ( .A1(n991), .A2(n990), .ZN(n992) );
  NAND2_X1 U1086 ( .A1(n993), .A2(n992), .ZN(n994) );
  XNOR2_X1 U1087 ( .A(n994), .B(KEYINPUT125), .ZN(n999) );
  XNOR2_X1 U1088 ( .A(G301), .B(G1961), .ZN(n997) );
  XNOR2_X1 U1089 ( .A(n995), .B(G1348), .ZN(n996) );
  NOR2_X1 U1090 ( .A1(n997), .A2(n996), .ZN(n998) );
  NAND2_X1 U1091 ( .A1(n999), .A2(n998), .ZN(n1002) );
  XNOR2_X1 U1092 ( .A(n1000), .B(G1341), .ZN(n1001) );
  NOR2_X1 U1093 ( .A1(n1002), .A2(n1001), .ZN(n1007) );
  XNOR2_X1 U1094 ( .A(G1966), .B(G168), .ZN(n1004) );
  NAND2_X1 U1095 ( .A1(n1004), .A2(n1003), .ZN(n1005) );
  XNOR2_X1 U1096 ( .A(n1005), .B(KEYINPUT57), .ZN(n1006) );
  NAND2_X1 U1097 ( .A1(n1007), .A2(n1006), .ZN(n1008) );
  NAND2_X1 U1098 ( .A1(n1009), .A2(n1008), .ZN(n1010) );
  XOR2_X1 U1099 ( .A(KEYINPUT126), .B(n1010), .Z(n1011) );
  NOR2_X1 U1100 ( .A1(n1012), .A2(n1011), .ZN(n1013) );
  NAND2_X1 U1101 ( .A1(n1014), .A2(n1013), .ZN(n1039) );
  XOR2_X1 U1102 ( .A(G2090), .B(G35), .Z(n1032) );
  XOR2_X1 U1103 ( .A(n1015), .B(KEYINPUT120), .Z(n1016) );
  XNOR2_X1 U1104 ( .A(n1016), .B(G25), .ZN(n1021) );
  XNOR2_X1 U1105 ( .A(G2067), .B(G26), .ZN(n1018) );
  XNOR2_X1 U1106 ( .A(G2072), .B(G33), .ZN(n1017) );
  NOR2_X1 U1107 ( .A1(n1018), .A2(n1017), .ZN(n1019) );
  XNOR2_X1 U1108 ( .A(n1019), .B(KEYINPUT121), .ZN(n1020) );
  NOR2_X1 U1109 ( .A1(n1021), .A2(n1020), .ZN(n1028) );
  XOR2_X1 U1110 ( .A(G32), .B(G1996), .Z(n1022) );
  NAND2_X1 U1111 ( .A1(n1022), .A2(G28), .ZN(n1026) );
  XNOR2_X1 U1112 ( .A(KEYINPUT122), .B(n1023), .ZN(n1024) );
  XNOR2_X1 U1113 ( .A(G27), .B(n1024), .ZN(n1025) );
  NOR2_X1 U1114 ( .A1(n1026), .A2(n1025), .ZN(n1027) );
  NAND2_X1 U1115 ( .A1(n1028), .A2(n1027), .ZN(n1029) );
  XOR2_X1 U1116 ( .A(KEYINPUT123), .B(n1029), .Z(n1030) );
  XNOR2_X1 U1117 ( .A(n1030), .B(KEYINPUT53), .ZN(n1031) );
  NAND2_X1 U1118 ( .A1(n1032), .A2(n1031), .ZN(n1035) );
  XNOR2_X1 U1119 ( .A(G34), .B(G2084), .ZN(n1033) );
  XNOR2_X1 U1120 ( .A(KEYINPUT54), .B(n1033), .ZN(n1034) );
  NOR2_X1 U1121 ( .A1(n1035), .A2(n1034), .ZN(n1036) );
  XOR2_X1 U1122 ( .A(KEYINPUT55), .B(n1036), .Z(n1037) );
  NOR2_X1 U1123 ( .A1(G29), .A2(n1037), .ZN(n1038) );
  NOR2_X1 U1124 ( .A1(n1039), .A2(n1038), .ZN(n1040) );
  XNOR2_X1 U1125 ( .A(n1040), .B(KEYINPUT62), .ZN(G311) );
  INV_X1 U1126 ( .A(G311), .ZN(G150) );
endmodule

