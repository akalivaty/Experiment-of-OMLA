//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 0 1 1 0 0 0 0 1 1 1 1 0 0 1 0 0 1 0 1 1 0 0 0 1 1 1 0 1 0 0 0 1 0 0 1 0 0 0 1 1 0 1 0 0 1 1 1 1 1 0 0 0 1 0 1 0 1 0 0 1 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:32:00 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n456, new_n457,
    new_n458, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n525,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n531, new_n532,
    new_n533, new_n534, new_n535, new_n536, new_n538, new_n539, new_n540,
    new_n541, new_n542, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n553, new_n554, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n571, new_n572, new_n574, new_n575, new_n576,
    new_n578, new_n579, new_n580, new_n581, new_n582, new_n583, new_n584,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n620, new_n623, new_n625, new_n626,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n854, new_n855, new_n856,
    new_n857, new_n858, new_n859, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1183, new_n1184,
    new_n1185, new_n1186, new_n1187, new_n1188, new_n1189, new_n1190,
    new_n1191, new_n1192, new_n1193, new_n1194, new_n1195, new_n1196,
    new_n1198, new_n1199, new_n1200;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  XOR2_X1   g008(.A(KEYINPUT64), .B(G44), .Z(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G218), .A2(G220), .A3(G221), .A4(G219), .ZN(new_n450));
  XOR2_X1   g025(.A(new_n450), .B(KEYINPUT2), .Z(new_n451));
  NOR4_X1   g026(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n452));
  INV_X1    g027(.A(new_n452), .ZN(new_n453));
  NOR2_X1   g028(.A1(new_n451), .A2(new_n453), .ZN(G325));
  XOR2_X1   g029(.A(G325), .B(KEYINPUT65), .Z(G261));
  NAND2_X1  g030(.A1(new_n451), .A2(G2106), .ZN(new_n456));
  NAND2_X1  g031(.A1(new_n453), .A2(G567), .ZN(new_n457));
  NAND2_X1  g032(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  INV_X1    g033(.A(new_n458), .ZN(G319));
  INV_X1    g034(.A(KEYINPUT67), .ZN(new_n460));
  INV_X1    g035(.A(KEYINPUT3), .ZN(new_n461));
  OAI21_X1  g036(.A(new_n460), .B1(new_n461), .B2(G2104), .ZN(new_n462));
  INV_X1    g037(.A(G2104), .ZN(new_n463));
  NAND3_X1  g038(.A1(new_n463), .A2(KEYINPUT67), .A3(KEYINPUT3), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n461), .A2(G2104), .ZN(new_n465));
  NAND4_X1  g040(.A1(new_n462), .A2(new_n464), .A3(G137), .A4(new_n465), .ZN(new_n466));
  NAND2_X1  g041(.A1(G101), .A2(G2104), .ZN(new_n467));
  AOI21_X1  g042(.A(G2105), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n463), .A2(KEYINPUT3), .ZN(new_n469));
  NAND3_X1  g044(.A1(new_n469), .A2(new_n465), .A3(G125), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n470), .A2(KEYINPUT66), .ZN(new_n471));
  INV_X1    g046(.A(KEYINPUT66), .ZN(new_n472));
  NAND4_X1  g047(.A1(new_n469), .A2(new_n465), .A3(new_n472), .A4(G125), .ZN(new_n473));
  NAND2_X1  g048(.A1(G113), .A2(G2104), .ZN(new_n474));
  NAND3_X1  g049(.A1(new_n471), .A2(new_n473), .A3(new_n474), .ZN(new_n475));
  AOI21_X1  g050(.A(new_n468), .B1(new_n475), .B2(G2105), .ZN(G160));
  NAND4_X1  g051(.A1(new_n462), .A2(new_n464), .A3(G2105), .A4(new_n465), .ZN(new_n477));
  INV_X1    g052(.A(G124), .ZN(new_n478));
  NOR2_X1   g053(.A1(G100), .A2(G2105), .ZN(new_n479));
  INV_X1    g054(.A(G2105), .ZN(new_n480));
  OAI21_X1  g055(.A(G2104), .B1(new_n480), .B2(G112), .ZN(new_n481));
  OAI22_X1  g056(.A1(new_n477), .A2(new_n478), .B1(new_n479), .B2(new_n481), .ZN(new_n482));
  AND4_X1   g057(.A1(new_n480), .A2(new_n462), .A3(new_n465), .A4(new_n464), .ZN(new_n483));
  AOI21_X1  g058(.A(new_n482), .B1(new_n483), .B2(G136), .ZN(G162));
  INV_X1    g059(.A(G138), .ZN(new_n485));
  NOR2_X1   g060(.A1(new_n485), .A2(G2105), .ZN(new_n486));
  NAND3_X1  g061(.A1(new_n486), .A2(new_n469), .A3(new_n465), .ZN(new_n487));
  INV_X1    g062(.A(KEYINPUT4), .ZN(new_n488));
  NAND2_X1  g063(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  AND3_X1   g064(.A1(new_n480), .A2(KEYINPUT4), .A3(G138), .ZN(new_n490));
  NAND4_X1  g065(.A1(new_n490), .A2(new_n462), .A3(new_n465), .A4(new_n464), .ZN(new_n491));
  INV_X1    g066(.A(G126), .ZN(new_n492));
  OAI211_X1 g067(.A(new_n489), .B(new_n491), .C1(new_n492), .C2(new_n477), .ZN(new_n493));
  OAI21_X1  g068(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n494));
  INV_X1    g069(.A(KEYINPUT69), .ZN(new_n495));
  XNOR2_X1  g070(.A(KEYINPUT68), .B(G114), .ZN(new_n496));
  OAI21_X1  g071(.A(new_n495), .B1(new_n496), .B2(new_n480), .ZN(new_n497));
  INV_X1    g072(.A(KEYINPUT68), .ZN(new_n498));
  NOR2_X1   g073(.A1(new_n498), .A2(G114), .ZN(new_n499));
  INV_X1    g074(.A(G114), .ZN(new_n500));
  NOR2_X1   g075(.A1(new_n500), .A2(KEYINPUT68), .ZN(new_n501));
  OAI211_X1 g076(.A(KEYINPUT69), .B(G2105), .C1(new_n499), .C2(new_n501), .ZN(new_n502));
  AOI21_X1  g077(.A(new_n494), .B1(new_n497), .B2(new_n502), .ZN(new_n503));
  NOR2_X1   g078(.A1(new_n493), .A2(new_n503), .ZN(G164));
  XNOR2_X1  g079(.A(KEYINPUT6), .B(G651), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n505), .A2(G543), .ZN(new_n506));
  INV_X1    g081(.A(G50), .ZN(new_n507));
  INV_X1    g082(.A(G651), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n508), .A2(KEYINPUT6), .ZN(new_n509));
  INV_X1    g084(.A(KEYINPUT6), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n510), .A2(G651), .ZN(new_n511));
  AND2_X1   g086(.A1(KEYINPUT5), .A2(G543), .ZN(new_n512));
  NOR2_X1   g087(.A1(KEYINPUT5), .A2(G543), .ZN(new_n513));
  OAI211_X1 g088(.A(new_n509), .B(new_n511), .C1(new_n512), .C2(new_n513), .ZN(new_n514));
  INV_X1    g089(.A(G88), .ZN(new_n515));
  OAI22_X1  g090(.A1(new_n506), .A2(new_n507), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n516), .A2(KEYINPUT70), .ZN(new_n517));
  INV_X1    g092(.A(KEYINPUT70), .ZN(new_n518));
  OAI221_X1 g093(.A(new_n518), .B1(new_n514), .B2(new_n515), .C1(new_n506), .C2(new_n507), .ZN(new_n519));
  NAND2_X1  g094(.A1(G75), .A2(G543), .ZN(new_n520));
  NOR2_X1   g095(.A1(new_n512), .A2(new_n513), .ZN(new_n521));
  INV_X1    g096(.A(G62), .ZN(new_n522));
  OAI21_X1  g097(.A(new_n520), .B1(new_n521), .B2(new_n522), .ZN(new_n523));
  AOI22_X1  g098(.A1(new_n517), .A2(new_n519), .B1(G651), .B2(new_n523), .ZN(G166));
  OR2_X1    g099(.A1(KEYINPUT5), .A2(G543), .ZN(new_n525));
  NAND2_X1  g100(.A1(KEYINPUT5), .A2(G543), .ZN(new_n526));
  NAND2_X1  g101(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  NAND3_X1  g102(.A1(new_n527), .A2(G63), .A3(G651), .ZN(new_n528));
  INV_X1    g103(.A(G51), .ZN(new_n529));
  OAI21_X1  g104(.A(new_n528), .B1(new_n506), .B2(new_n529), .ZN(new_n530));
  NAND3_X1  g105(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n531));
  XNOR2_X1  g106(.A(new_n531), .B(KEYINPUT7), .ZN(new_n532));
  INV_X1    g107(.A(G89), .ZN(new_n533));
  OAI21_X1  g108(.A(new_n532), .B1(new_n533), .B2(new_n514), .ZN(new_n534));
  OR3_X1    g109(.A1(new_n530), .A2(new_n534), .A3(KEYINPUT71), .ZN(new_n535));
  OAI21_X1  g110(.A(KEYINPUT71), .B1(new_n530), .B2(new_n534), .ZN(new_n536));
  NAND2_X1  g111(.A1(new_n535), .A2(new_n536), .ZN(G168));
  AOI22_X1  g112(.A1(new_n527), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n538));
  NOR2_X1   g113(.A1(new_n538), .A2(new_n508), .ZN(new_n539));
  INV_X1    g114(.A(G52), .ZN(new_n540));
  INV_X1    g115(.A(G90), .ZN(new_n541));
  OAI22_X1  g116(.A1(new_n506), .A2(new_n540), .B1(new_n514), .B2(new_n541), .ZN(new_n542));
  NOR2_X1   g117(.A1(new_n539), .A2(new_n542), .ZN(G171));
  AOI22_X1  g118(.A1(new_n527), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n544));
  NOR2_X1   g119(.A1(new_n544), .A2(new_n508), .ZN(new_n545));
  INV_X1    g120(.A(G43), .ZN(new_n546));
  INV_X1    g121(.A(G81), .ZN(new_n547));
  OAI22_X1  g122(.A1(new_n506), .A2(new_n546), .B1(new_n514), .B2(new_n547), .ZN(new_n548));
  OR2_X1    g123(.A1(new_n545), .A2(new_n548), .ZN(new_n549));
  INV_X1    g124(.A(new_n549), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n550), .A2(G860), .ZN(G153));
  NAND4_X1  g126(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g127(.A1(G1), .A2(G3), .ZN(new_n553));
  XNOR2_X1  g128(.A(new_n553), .B(KEYINPUT8), .ZN(new_n554));
  NAND4_X1  g129(.A1(G319), .A2(G483), .A3(G661), .A4(new_n554), .ZN(G188));
  AND2_X1   g130(.A1(new_n527), .A2(G65), .ZN(new_n556));
  NAND2_X1  g131(.A1(G78), .A2(G543), .ZN(new_n557));
  XOR2_X1   g132(.A(new_n557), .B(KEYINPUT73), .Z(new_n558));
  OAI21_X1  g133(.A(G651), .B1(new_n556), .B2(new_n558), .ZN(new_n559));
  INV_X1    g134(.A(G53), .ZN(new_n560));
  NOR2_X1   g135(.A1(new_n560), .A2(KEYINPUT72), .ZN(new_n561));
  NAND3_X1  g136(.A1(new_n505), .A2(G543), .A3(new_n561), .ZN(new_n562));
  INV_X1    g137(.A(KEYINPUT9), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  NAND4_X1  g139(.A1(new_n505), .A2(KEYINPUT9), .A3(G543), .A4(new_n561), .ZN(new_n565));
  INV_X1    g140(.A(new_n514), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n566), .A2(G91), .ZN(new_n567));
  NAND4_X1  g142(.A1(new_n559), .A2(new_n564), .A3(new_n565), .A4(new_n567), .ZN(G299));
  INV_X1    g143(.A(G171), .ZN(G301));
  INV_X1    g144(.A(G168), .ZN(G286));
  NAND2_X1  g145(.A1(new_n517), .A2(new_n519), .ZN(new_n571));
  NAND2_X1  g146(.A1(new_n523), .A2(G651), .ZN(new_n572));
  NAND2_X1  g147(.A1(new_n571), .A2(new_n572), .ZN(G303));
  NAND2_X1  g148(.A1(new_n566), .A2(G87), .ZN(new_n574));
  OAI21_X1  g149(.A(G651), .B1(new_n527), .B2(G74), .ZN(new_n575));
  NAND3_X1  g150(.A1(new_n505), .A2(G49), .A3(G543), .ZN(new_n576));
  NAND3_X1  g151(.A1(new_n574), .A2(new_n575), .A3(new_n576), .ZN(G288));
  INV_X1    g152(.A(G61), .ZN(new_n578));
  AOI21_X1  g153(.A(new_n578), .B1(new_n525), .B2(new_n526), .ZN(new_n579));
  NAND2_X1  g154(.A1(G73), .A2(G543), .ZN(new_n580));
  INV_X1    g155(.A(new_n580), .ZN(new_n581));
  OAI21_X1  g156(.A(G651), .B1(new_n579), .B2(new_n581), .ZN(new_n582));
  NAND3_X1  g157(.A1(new_n527), .A2(new_n505), .A3(G86), .ZN(new_n583));
  NAND3_X1  g158(.A1(new_n505), .A2(G48), .A3(G543), .ZN(new_n584));
  NAND3_X1  g159(.A1(new_n582), .A2(new_n583), .A3(new_n584), .ZN(G305));
  INV_X1    g160(.A(G47), .ZN(new_n586));
  INV_X1    g161(.A(G85), .ZN(new_n587));
  OAI22_X1  g162(.A1(new_n506), .A2(new_n586), .B1(new_n514), .B2(new_n587), .ZN(new_n588));
  XOR2_X1   g163(.A(new_n588), .B(KEYINPUT76), .Z(new_n589));
  INV_X1    g164(.A(G60), .ZN(new_n590));
  INV_X1    g165(.A(G72), .ZN(new_n591));
  INV_X1    g166(.A(G543), .ZN(new_n592));
  OAI22_X1  g167(.A1(new_n521), .A2(new_n590), .B1(new_n591), .B2(new_n592), .ZN(new_n593));
  INV_X1    g168(.A(KEYINPUT74), .ZN(new_n594));
  NAND2_X1  g169(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  OAI221_X1 g170(.A(KEYINPUT74), .B1(new_n591), .B2(new_n592), .C1(new_n521), .C2(new_n590), .ZN(new_n596));
  NAND3_X1  g171(.A1(new_n595), .A2(G651), .A3(new_n596), .ZN(new_n597));
  INV_X1    g172(.A(KEYINPUT75), .ZN(new_n598));
  OR2_X1    g173(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  NAND2_X1  g174(.A1(new_n597), .A2(new_n598), .ZN(new_n600));
  NAND3_X1  g175(.A1(new_n589), .A2(new_n599), .A3(new_n600), .ZN(new_n601));
  INV_X1    g176(.A(KEYINPUT77), .ZN(new_n602));
  OR2_X1    g177(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  NAND2_X1  g178(.A1(new_n601), .A2(new_n602), .ZN(new_n604));
  NAND2_X1  g179(.A1(new_n603), .A2(new_n604), .ZN(G290));
  NAND2_X1  g180(.A1(G301), .A2(G868), .ZN(new_n606));
  NAND2_X1  g181(.A1(new_n566), .A2(G92), .ZN(new_n607));
  XOR2_X1   g182(.A(new_n607), .B(KEYINPUT10), .Z(new_n608));
  AOI22_X1  g183(.A1(new_n527), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n609));
  NOR2_X1   g184(.A1(new_n609), .A2(new_n508), .ZN(new_n610));
  NAND3_X1  g185(.A1(new_n505), .A2(KEYINPUT78), .A3(G543), .ZN(new_n611));
  INV_X1    g186(.A(G54), .ZN(new_n612));
  INV_X1    g187(.A(KEYINPUT78), .ZN(new_n613));
  AOI21_X1  g188(.A(new_n612), .B1(new_n506), .B2(new_n613), .ZN(new_n614));
  AOI21_X1  g189(.A(new_n610), .B1(new_n611), .B2(new_n614), .ZN(new_n615));
  NAND2_X1  g190(.A1(new_n608), .A2(new_n615), .ZN(new_n616));
  INV_X1    g191(.A(new_n616), .ZN(new_n617));
  OAI21_X1  g192(.A(new_n606), .B1(new_n617), .B2(G868), .ZN(G284));
  OAI21_X1  g193(.A(new_n606), .B1(new_n617), .B2(G868), .ZN(G321));
  NOR2_X1   g194(.A1(G299), .A2(G868), .ZN(new_n620));
  AOI21_X1  g195(.A(new_n620), .B1(G168), .B2(G868), .ZN(G297));
  AOI21_X1  g196(.A(new_n620), .B1(G168), .B2(G868), .ZN(G280));
  INV_X1    g197(.A(G559), .ZN(new_n623));
  OAI21_X1  g198(.A(new_n617), .B1(new_n623), .B2(G860), .ZN(G148));
  NAND2_X1  g199(.A1(new_n617), .A2(new_n623), .ZN(new_n625));
  NAND2_X1  g200(.A1(new_n625), .A2(G868), .ZN(new_n626));
  OAI21_X1  g201(.A(new_n626), .B1(G868), .B2(new_n550), .ZN(G323));
  XNOR2_X1  g202(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g203(.A1(new_n483), .A2(G135), .ZN(new_n629));
  XNOR2_X1  g204(.A(new_n629), .B(KEYINPUT79), .ZN(new_n630));
  INV_X1    g205(.A(new_n477), .ZN(new_n631));
  NAND2_X1  g206(.A1(new_n631), .A2(G123), .ZN(new_n632));
  NOR2_X1   g207(.A1(G99), .A2(G2105), .ZN(new_n633));
  OAI21_X1  g208(.A(G2104), .B1(new_n480), .B2(G111), .ZN(new_n634));
  OAI211_X1 g209(.A(new_n630), .B(new_n632), .C1(new_n633), .C2(new_n634), .ZN(new_n635));
  XNOR2_X1  g210(.A(new_n635), .B(KEYINPUT80), .ZN(new_n636));
  INV_X1    g211(.A(G2096), .ZN(new_n637));
  OR2_X1    g212(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  NAND2_X1  g213(.A1(new_n636), .A2(new_n637), .ZN(new_n639));
  NAND3_X1  g214(.A1(new_n480), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n640));
  XNOR2_X1  g215(.A(new_n640), .B(KEYINPUT12), .ZN(new_n641));
  XNOR2_X1  g216(.A(new_n641), .B(KEYINPUT13), .ZN(new_n642));
  XNOR2_X1  g217(.A(new_n642), .B(G2100), .ZN(new_n643));
  NAND3_X1  g218(.A1(new_n638), .A2(new_n639), .A3(new_n643), .ZN(G156));
  XNOR2_X1  g219(.A(G2427), .B(G2438), .ZN(new_n645));
  XNOR2_X1  g220(.A(new_n645), .B(G2430), .ZN(new_n646));
  XNOR2_X1  g221(.A(KEYINPUT15), .B(G2435), .ZN(new_n647));
  OR2_X1    g222(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  NAND2_X1  g223(.A1(new_n646), .A2(new_n647), .ZN(new_n649));
  NAND3_X1  g224(.A1(new_n648), .A2(KEYINPUT14), .A3(new_n649), .ZN(new_n650));
  XNOR2_X1  g225(.A(G2451), .B(G2454), .ZN(new_n651));
  XNOR2_X1  g226(.A(new_n651), .B(KEYINPUT16), .ZN(new_n652));
  XNOR2_X1  g227(.A(new_n650), .B(new_n652), .ZN(new_n653));
  XNOR2_X1  g228(.A(G2443), .B(G2446), .ZN(new_n654));
  OR2_X1    g229(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  XNOR2_X1  g230(.A(G1341), .B(G1348), .ZN(new_n656));
  INV_X1    g231(.A(new_n656), .ZN(new_n657));
  NAND2_X1  g232(.A1(new_n653), .A2(new_n654), .ZN(new_n658));
  NAND3_X1  g233(.A1(new_n655), .A2(new_n657), .A3(new_n658), .ZN(new_n659));
  NAND2_X1  g234(.A1(new_n659), .A2(G14), .ZN(new_n660));
  INV_X1    g235(.A(KEYINPUT81), .ZN(new_n661));
  INV_X1    g236(.A(new_n654), .ZN(new_n662));
  XNOR2_X1  g237(.A(new_n653), .B(new_n662), .ZN(new_n663));
  OAI21_X1  g238(.A(new_n661), .B1(new_n663), .B2(new_n657), .ZN(new_n664));
  NAND2_X1  g239(.A1(new_n655), .A2(new_n658), .ZN(new_n665));
  NAND3_X1  g240(.A1(new_n665), .A2(KEYINPUT81), .A3(new_n656), .ZN(new_n666));
  AOI21_X1  g241(.A(new_n660), .B1(new_n664), .B2(new_n666), .ZN(G401));
  XOR2_X1   g242(.A(G2084), .B(G2090), .Z(new_n668));
  XNOR2_X1  g243(.A(G2067), .B(G2678), .ZN(new_n669));
  NAND2_X1  g244(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  INV_X1    g245(.A(new_n668), .ZN(new_n671));
  XOR2_X1   g246(.A(G2072), .B(G2078), .Z(new_n672));
  NAND2_X1  g247(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  XNOR2_X1  g248(.A(new_n672), .B(KEYINPUT17), .ZN(new_n674));
  NOR2_X1   g249(.A1(new_n668), .A2(new_n669), .ZN(new_n675));
  OAI221_X1 g250(.A(new_n670), .B1(new_n669), .B2(new_n673), .C1(new_n674), .C2(new_n675), .ZN(new_n676));
  NOR2_X1   g251(.A1(new_n670), .A2(new_n672), .ZN(new_n677));
  XNOR2_X1  g252(.A(new_n677), .B(KEYINPUT18), .ZN(new_n678));
  NAND2_X1  g253(.A1(new_n676), .A2(new_n678), .ZN(new_n679));
  XNOR2_X1  g254(.A(new_n679), .B(new_n637), .ZN(new_n680));
  XNOR2_X1  g255(.A(new_n680), .B(G2100), .ZN(G227));
  XNOR2_X1  g256(.A(G1971), .B(G1976), .ZN(new_n682));
  INV_X1    g257(.A(KEYINPUT19), .ZN(new_n683));
  XNOR2_X1  g258(.A(new_n682), .B(new_n683), .ZN(new_n684));
  XOR2_X1   g259(.A(G1956), .B(G2474), .Z(new_n685));
  XOR2_X1   g260(.A(G1961), .B(G1966), .Z(new_n686));
  AND2_X1   g261(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  NAND2_X1  g262(.A1(new_n684), .A2(new_n687), .ZN(new_n688));
  INV_X1    g263(.A(KEYINPUT20), .ZN(new_n689));
  XNOR2_X1  g264(.A(new_n688), .B(new_n689), .ZN(new_n690));
  NOR2_X1   g265(.A1(new_n685), .A2(new_n686), .ZN(new_n691));
  NOR2_X1   g266(.A1(new_n687), .A2(new_n691), .ZN(new_n692));
  MUX2_X1   g267(.A(new_n692), .B(new_n691), .S(new_n684), .Z(new_n693));
  NOR2_X1   g268(.A1(new_n690), .A2(new_n693), .ZN(new_n694));
  INV_X1    g269(.A(G1986), .ZN(new_n695));
  XNOR2_X1  g270(.A(new_n694), .B(new_n695), .ZN(new_n696));
  XNOR2_X1  g271(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n697));
  XNOR2_X1  g272(.A(new_n696), .B(new_n697), .ZN(new_n698));
  XNOR2_X1  g273(.A(G1991), .B(G1996), .ZN(new_n699));
  INV_X1    g274(.A(G1981), .ZN(new_n700));
  XNOR2_X1  g275(.A(new_n699), .B(new_n700), .ZN(new_n701));
  XNOR2_X1  g276(.A(new_n698), .B(new_n701), .ZN(new_n702));
  INV_X1    g277(.A(new_n702), .ZN(G229));
  INV_X1    g278(.A(G119), .ZN(new_n704));
  NOR2_X1   g279(.A1(G95), .A2(G2105), .ZN(new_n705));
  OAI21_X1  g280(.A(G2104), .B1(new_n480), .B2(G107), .ZN(new_n706));
  OAI22_X1  g281(.A1(new_n477), .A2(new_n704), .B1(new_n705), .B2(new_n706), .ZN(new_n707));
  AOI21_X1  g282(.A(new_n707), .B1(new_n483), .B2(G131), .ZN(new_n708));
  XOR2_X1   g283(.A(new_n708), .B(KEYINPUT82), .Z(new_n709));
  MUX2_X1   g284(.A(G25), .B(new_n709), .S(G29), .Z(new_n710));
  XOR2_X1   g285(.A(KEYINPUT35), .B(G1991), .Z(new_n711));
  XNOR2_X1  g286(.A(new_n711), .B(KEYINPUT83), .ZN(new_n712));
  XNOR2_X1  g287(.A(new_n710), .B(new_n712), .ZN(new_n713));
  INV_X1    g288(.A(G16), .ZN(new_n714));
  NAND2_X1  g289(.A1(new_n714), .A2(G24), .ZN(new_n715));
  INV_X1    g290(.A(G290), .ZN(new_n716));
  OAI21_X1  g291(.A(new_n715), .B1(new_n716), .B2(new_n714), .ZN(new_n717));
  AOI21_X1  g292(.A(new_n713), .B1(G1986), .B2(new_n717), .ZN(new_n718));
  OAI21_X1  g293(.A(new_n718), .B1(G1986), .B2(new_n717), .ZN(new_n719));
  INV_X1    g294(.A(KEYINPUT87), .ZN(new_n720));
  NAND2_X1  g295(.A1(new_n720), .A2(KEYINPUT36), .ZN(new_n721));
  XNOR2_X1  g296(.A(new_n721), .B(KEYINPUT88), .ZN(new_n722));
  INV_X1    g297(.A(new_n722), .ZN(new_n723));
  NOR2_X1   g298(.A1(G16), .A2(G23), .ZN(new_n724));
  XOR2_X1   g299(.A(new_n724), .B(KEYINPUT85), .Z(new_n725));
  INV_X1    g300(.A(KEYINPUT86), .ZN(new_n726));
  NAND2_X1  g301(.A1(G288), .A2(new_n726), .ZN(new_n727));
  NAND4_X1  g302(.A1(new_n574), .A2(KEYINPUT86), .A3(new_n575), .A4(new_n576), .ZN(new_n728));
  NAND2_X1  g303(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  OAI21_X1  g304(.A(new_n725), .B1(new_n729), .B2(new_n714), .ZN(new_n730));
  XOR2_X1   g305(.A(KEYINPUT33), .B(G1976), .Z(new_n731));
  XNOR2_X1  g306(.A(new_n730), .B(new_n731), .ZN(new_n732));
  NAND2_X1  g307(.A1(new_n714), .A2(G22), .ZN(new_n733));
  OAI21_X1  g308(.A(new_n733), .B1(G166), .B2(new_n714), .ZN(new_n734));
  OR2_X1    g309(.A1(new_n734), .A2(G1971), .ZN(new_n735));
  NAND2_X1  g310(.A1(new_n714), .A2(G6), .ZN(new_n736));
  NAND2_X1  g311(.A1(new_n583), .A2(new_n584), .ZN(new_n737));
  OAI21_X1  g312(.A(G61), .B1(new_n512), .B2(new_n513), .ZN(new_n738));
  AOI21_X1  g313(.A(new_n508), .B1(new_n738), .B2(new_n580), .ZN(new_n739));
  NOR2_X1   g314(.A1(new_n737), .A2(new_n739), .ZN(new_n740));
  OAI21_X1  g315(.A(new_n736), .B1(new_n740), .B2(new_n714), .ZN(new_n741));
  XOR2_X1   g316(.A(KEYINPUT32), .B(G1981), .Z(new_n742));
  XNOR2_X1  g317(.A(new_n742), .B(KEYINPUT84), .ZN(new_n743));
  XNOR2_X1  g318(.A(new_n741), .B(new_n743), .ZN(new_n744));
  NAND2_X1  g319(.A1(new_n734), .A2(G1971), .ZN(new_n745));
  NAND4_X1  g320(.A1(new_n732), .A2(new_n735), .A3(new_n744), .A4(new_n745), .ZN(new_n746));
  XNOR2_X1  g321(.A(new_n746), .B(KEYINPUT34), .ZN(new_n747));
  NOR3_X1   g322(.A1(new_n719), .A2(new_n723), .A3(new_n747), .ZN(new_n748));
  INV_X1    g323(.A(G29), .ZN(new_n749));
  NAND2_X1  g324(.A1(new_n749), .A2(G33), .ZN(new_n750));
  NAND2_X1  g325(.A1(new_n483), .A2(G139), .ZN(new_n751));
  NAND3_X1  g326(.A1(new_n480), .A2(G103), .A3(G2104), .ZN(new_n752));
  XOR2_X1   g327(.A(new_n752), .B(KEYINPUT25), .Z(new_n753));
  AND2_X1   g328(.A1(new_n469), .A2(new_n465), .ZN(new_n754));
  AOI22_X1  g329(.A1(new_n754), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n755));
  OAI211_X1 g330(.A(new_n751), .B(new_n753), .C1(new_n480), .C2(new_n755), .ZN(new_n756));
  XNOR2_X1  g331(.A(new_n756), .B(KEYINPUT91), .ZN(new_n757));
  INV_X1    g332(.A(new_n757), .ZN(new_n758));
  OAI21_X1  g333(.A(new_n750), .B1(new_n758), .B2(new_n749), .ZN(new_n759));
  XNOR2_X1  g334(.A(new_n759), .B(G2072), .ZN(new_n760));
  NAND2_X1  g335(.A1(new_n749), .A2(G32), .ZN(new_n761));
  NAND2_X1  g336(.A1(new_n631), .A2(G129), .ZN(new_n762));
  NAND3_X1  g337(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n763));
  XOR2_X1   g338(.A(new_n763), .B(KEYINPUT26), .Z(new_n764));
  NAND3_X1  g339(.A1(new_n480), .A2(G105), .A3(G2104), .ZN(new_n765));
  XOR2_X1   g340(.A(new_n765), .B(KEYINPUT92), .Z(new_n766));
  NAND3_X1  g341(.A1(new_n762), .A2(new_n764), .A3(new_n766), .ZN(new_n767));
  AND2_X1   g342(.A1(new_n483), .A2(G141), .ZN(new_n768));
  NOR2_X1   g343(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  XOR2_X1   g344(.A(new_n769), .B(KEYINPUT93), .Z(new_n770));
  INV_X1    g345(.A(new_n770), .ZN(new_n771));
  OAI21_X1  g346(.A(new_n761), .B1(new_n771), .B2(new_n749), .ZN(new_n772));
  INV_X1    g347(.A(new_n772), .ZN(new_n773));
  XNOR2_X1  g348(.A(KEYINPUT27), .B(G1996), .ZN(new_n774));
  AOI21_X1  g349(.A(new_n760), .B1(new_n773), .B2(new_n774), .ZN(new_n775));
  NAND2_X1  g350(.A1(new_n749), .A2(G35), .ZN(new_n776));
  OAI21_X1  g351(.A(new_n776), .B1(G162), .B2(new_n749), .ZN(new_n777));
  XOR2_X1   g352(.A(new_n777), .B(KEYINPUT29), .Z(new_n778));
  INV_X1    g353(.A(G2090), .ZN(new_n779));
  NOR2_X1   g354(.A1(new_n778), .A2(new_n779), .ZN(new_n780));
  XNOR2_X1  g355(.A(new_n780), .B(KEYINPUT95), .ZN(new_n781));
  INV_X1    g356(.A(new_n774), .ZN(new_n782));
  AOI22_X1  g357(.A1(new_n772), .A2(new_n782), .B1(new_n778), .B2(new_n779), .ZN(new_n783));
  NAND3_X1  g358(.A1(new_n775), .A2(new_n781), .A3(new_n783), .ZN(new_n784));
  INV_X1    g359(.A(new_n784), .ZN(new_n785));
  NAND2_X1  g360(.A1(new_n631), .A2(G128), .ZN(new_n786));
  NAND2_X1  g361(.A1(new_n483), .A2(G140), .ZN(new_n787));
  NOR2_X1   g362(.A1(G104), .A2(G2105), .ZN(new_n788));
  OAI21_X1  g363(.A(G2104), .B1(new_n480), .B2(G116), .ZN(new_n789));
  OAI211_X1 g364(.A(new_n786), .B(new_n787), .C1(new_n788), .C2(new_n789), .ZN(new_n790));
  NAND2_X1  g365(.A1(new_n790), .A2(G29), .ZN(new_n791));
  XNOR2_X1  g366(.A(new_n791), .B(KEYINPUT90), .ZN(new_n792));
  NAND2_X1  g367(.A1(new_n749), .A2(G26), .ZN(new_n793));
  XNOR2_X1  g368(.A(new_n793), .B(KEYINPUT28), .ZN(new_n794));
  NAND2_X1  g369(.A1(new_n792), .A2(new_n794), .ZN(new_n795));
  INV_X1    g370(.A(G2067), .ZN(new_n796));
  XNOR2_X1  g371(.A(new_n795), .B(new_n796), .ZN(new_n797));
  NAND2_X1  g372(.A1(new_n616), .A2(G16), .ZN(new_n798));
  NAND2_X1  g373(.A1(new_n714), .A2(G4), .ZN(new_n799));
  NAND2_X1  g374(.A1(new_n798), .A2(new_n799), .ZN(new_n800));
  INV_X1    g375(.A(new_n800), .ZN(new_n801));
  INV_X1    g376(.A(G1348), .ZN(new_n802));
  NAND2_X1  g377(.A1(new_n714), .A2(G21), .ZN(new_n803));
  OAI21_X1  g378(.A(new_n803), .B1(G168), .B2(new_n714), .ZN(new_n804));
  XNOR2_X1  g379(.A(KEYINPUT94), .B(G1966), .ZN(new_n805));
  INV_X1    g380(.A(new_n805), .ZN(new_n806));
  AOI22_X1  g381(.A1(new_n801), .A2(new_n802), .B1(new_n804), .B2(new_n806), .ZN(new_n807));
  NAND2_X1  g382(.A1(new_n749), .A2(G27), .ZN(new_n808));
  OAI21_X1  g383(.A(new_n808), .B1(G164), .B2(new_n749), .ZN(new_n809));
  INV_X1    g384(.A(G2078), .ZN(new_n810));
  XNOR2_X1  g385(.A(new_n809), .B(new_n810), .ZN(new_n811));
  NOR2_X1   g386(.A1(new_n804), .A2(new_n806), .ZN(new_n812));
  INV_X1    g387(.A(KEYINPUT24), .ZN(new_n813));
  INV_X1    g388(.A(G34), .ZN(new_n814));
  AOI21_X1  g389(.A(G29), .B1(new_n813), .B2(new_n814), .ZN(new_n815));
  OAI21_X1  g390(.A(new_n815), .B1(new_n813), .B2(new_n814), .ZN(new_n816));
  OAI21_X1  g391(.A(new_n816), .B1(G160), .B2(new_n749), .ZN(new_n817));
  AOI21_X1  g392(.A(new_n812), .B1(G2084), .B2(new_n817), .ZN(new_n818));
  NOR2_X1   g393(.A1(new_n817), .A2(G2084), .ZN(new_n819));
  AOI21_X1  g394(.A(new_n819), .B1(new_n800), .B2(G1348), .ZN(new_n820));
  NAND4_X1  g395(.A1(new_n807), .A2(new_n811), .A3(new_n818), .A4(new_n820), .ZN(new_n821));
  INV_X1    g396(.A(new_n821), .ZN(new_n822));
  NAND2_X1  g397(.A1(new_n714), .A2(G19), .ZN(new_n823));
  OAI21_X1  g398(.A(new_n823), .B1(new_n550), .B2(new_n714), .ZN(new_n824));
  INV_X1    g399(.A(KEYINPUT89), .ZN(new_n825));
  XNOR2_X1  g400(.A(new_n824), .B(new_n825), .ZN(new_n826));
  XNOR2_X1  g401(.A(new_n826), .B(G1341), .ZN(new_n827));
  NAND2_X1  g402(.A1(new_n636), .A2(G29), .ZN(new_n828));
  NOR2_X1   g403(.A1(G171), .A2(new_n714), .ZN(new_n829));
  AOI21_X1  g404(.A(new_n829), .B1(G5), .B2(new_n714), .ZN(new_n830));
  INV_X1    g405(.A(G1961), .ZN(new_n831));
  AND2_X1   g406(.A1(new_n830), .A2(new_n831), .ZN(new_n832));
  NOR2_X1   g407(.A1(new_n830), .A2(new_n831), .ZN(new_n833));
  INV_X1    g408(.A(KEYINPUT30), .ZN(new_n834));
  AND2_X1   g409(.A1(new_n834), .A2(G28), .ZN(new_n835));
  OAI21_X1  g410(.A(new_n749), .B1(new_n834), .B2(G28), .ZN(new_n836));
  AND2_X1   g411(.A1(KEYINPUT31), .A2(G11), .ZN(new_n837));
  NOR2_X1   g412(.A1(KEYINPUT31), .A2(G11), .ZN(new_n838));
  OAI22_X1  g413(.A1(new_n835), .A2(new_n836), .B1(new_n837), .B2(new_n838), .ZN(new_n839));
  NOR3_X1   g414(.A1(new_n832), .A2(new_n833), .A3(new_n839), .ZN(new_n840));
  XOR2_X1   g415(.A(KEYINPUT96), .B(KEYINPUT23), .Z(new_n841));
  NAND2_X1  g416(.A1(new_n714), .A2(G20), .ZN(new_n842));
  XNOR2_X1  g417(.A(new_n841), .B(new_n842), .ZN(new_n843));
  INV_X1    g418(.A(G299), .ZN(new_n844));
  OAI21_X1  g419(.A(new_n843), .B1(new_n844), .B2(new_n714), .ZN(new_n845));
  INV_X1    g420(.A(G1956), .ZN(new_n846));
  XNOR2_X1  g421(.A(new_n845), .B(new_n846), .ZN(new_n847));
  AND3_X1   g422(.A1(new_n828), .A2(new_n840), .A3(new_n847), .ZN(new_n848));
  AND3_X1   g423(.A1(new_n822), .A2(new_n827), .A3(new_n848), .ZN(new_n849));
  NAND4_X1  g424(.A1(new_n785), .A2(KEYINPUT97), .A3(new_n797), .A4(new_n849), .ZN(new_n850));
  INV_X1    g425(.A(KEYINPUT97), .ZN(new_n851));
  NAND4_X1  g426(.A1(new_n822), .A2(new_n797), .A3(new_n827), .A4(new_n848), .ZN(new_n852));
  OAI21_X1  g427(.A(new_n851), .B1(new_n784), .B2(new_n852), .ZN(new_n853));
  AOI21_X1  g428(.A(new_n748), .B1(new_n850), .B2(new_n853), .ZN(new_n854));
  OAI21_X1  g429(.A(new_n723), .B1(new_n719), .B2(new_n747), .ZN(new_n855));
  AOI21_X1  g430(.A(KEYINPUT98), .B1(new_n854), .B2(new_n855), .ZN(new_n856));
  NAND2_X1  g431(.A1(new_n850), .A2(new_n853), .ZN(new_n857));
  OR3_X1    g432(.A1(new_n719), .A2(new_n723), .A3(new_n747), .ZN(new_n858));
  AND4_X1   g433(.A1(KEYINPUT98), .A2(new_n857), .A3(new_n855), .A4(new_n858), .ZN(new_n859));
  NOR2_X1   g434(.A1(new_n856), .A2(new_n859), .ZN(G311));
  NAND2_X1  g435(.A1(new_n854), .A2(new_n855), .ZN(G150));
  NOR2_X1   g436(.A1(new_n616), .A2(new_n623), .ZN(new_n862));
  XNOR2_X1  g437(.A(new_n862), .B(KEYINPUT38), .ZN(new_n863));
  INV_X1    g438(.A(G55), .ZN(new_n864));
  INV_X1    g439(.A(G93), .ZN(new_n865));
  OAI22_X1  g440(.A1(new_n506), .A2(new_n864), .B1(new_n514), .B2(new_n865), .ZN(new_n866));
  INV_X1    g441(.A(KEYINPUT100), .ZN(new_n867));
  XNOR2_X1  g442(.A(new_n866), .B(new_n867), .ZN(new_n868));
  INV_X1    g443(.A(KEYINPUT101), .ZN(new_n869));
  NAND2_X1  g444(.A1(G80), .A2(G543), .ZN(new_n870));
  INV_X1    g445(.A(G67), .ZN(new_n871));
  OAI21_X1  g446(.A(new_n870), .B1(new_n521), .B2(new_n871), .ZN(new_n872));
  AOI21_X1  g447(.A(new_n508), .B1(new_n872), .B2(KEYINPUT99), .ZN(new_n873));
  OAI21_X1  g448(.A(new_n873), .B1(KEYINPUT99), .B2(new_n872), .ZN(new_n874));
  NAND3_X1  g449(.A1(new_n868), .A2(new_n869), .A3(new_n874), .ZN(new_n875));
  INV_X1    g450(.A(new_n875), .ZN(new_n876));
  AOI21_X1  g451(.A(new_n869), .B1(new_n868), .B2(new_n874), .ZN(new_n877));
  OAI21_X1  g452(.A(new_n549), .B1(new_n876), .B2(new_n877), .ZN(new_n878));
  INV_X1    g453(.A(new_n877), .ZN(new_n879));
  NAND3_X1  g454(.A1(new_n879), .A2(new_n550), .A3(new_n875), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n878), .A2(new_n880), .ZN(new_n881));
  XNOR2_X1  g456(.A(new_n863), .B(new_n881), .ZN(new_n882));
  INV_X1    g457(.A(KEYINPUT39), .ZN(new_n883));
  AOI21_X1  g458(.A(G860), .B1(new_n882), .B2(new_n883), .ZN(new_n884));
  OAI21_X1  g459(.A(new_n884), .B1(new_n883), .B2(new_n882), .ZN(new_n885));
  XOR2_X1   g460(.A(new_n885), .B(KEYINPUT102), .Z(new_n886));
  NAND2_X1  g461(.A1(new_n868), .A2(new_n874), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n887), .A2(G860), .ZN(new_n888));
  XOR2_X1   g463(.A(new_n888), .B(KEYINPUT37), .Z(new_n889));
  NAND2_X1  g464(.A1(new_n886), .A2(new_n889), .ZN(G145));
  XNOR2_X1  g465(.A(new_n636), .B(G160), .ZN(new_n891));
  XNOR2_X1  g466(.A(new_n891), .B(G162), .ZN(new_n892));
  INV_X1    g467(.A(new_n892), .ZN(new_n893));
  XNOR2_X1  g468(.A(G164), .B(new_n790), .ZN(new_n894));
  INV_X1    g469(.A(KEYINPUT103), .ZN(new_n895));
  AND2_X1   g470(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  NOR2_X1   g471(.A1(new_n894), .A2(new_n895), .ZN(new_n897));
  OR3_X1    g472(.A1(new_n896), .A2(new_n897), .A3(new_n770), .ZN(new_n898));
  OAI21_X1  g473(.A(new_n770), .B1(new_n896), .B2(new_n897), .ZN(new_n899));
  NAND3_X1  g474(.A1(new_n898), .A2(new_n758), .A3(new_n899), .ZN(new_n900));
  AOI21_X1  g475(.A(new_n758), .B1(new_n769), .B2(new_n894), .ZN(new_n901));
  OAI21_X1  g476(.A(new_n901), .B1(new_n769), .B2(new_n894), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n900), .A2(new_n902), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n631), .A2(G130), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n483), .A2(G142), .ZN(new_n905));
  NOR2_X1   g480(.A1(G106), .A2(G2105), .ZN(new_n906));
  OAI21_X1  g481(.A(G2104), .B1(new_n480), .B2(G118), .ZN(new_n907));
  OAI211_X1 g482(.A(new_n904), .B(new_n905), .C1(new_n906), .C2(new_n907), .ZN(new_n908));
  XNOR2_X1  g483(.A(new_n908), .B(KEYINPUT104), .ZN(new_n909));
  XNOR2_X1  g484(.A(new_n909), .B(new_n641), .ZN(new_n910));
  XNOR2_X1  g485(.A(new_n910), .B(new_n708), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n903), .A2(new_n911), .ZN(new_n912));
  INV_X1    g487(.A(new_n911), .ZN(new_n913));
  NAND3_X1  g488(.A1(new_n913), .A2(new_n902), .A3(new_n900), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n912), .A2(new_n914), .ZN(new_n915));
  AOI21_X1  g490(.A(G37), .B1(new_n893), .B2(new_n915), .ZN(new_n916));
  INV_X1    g491(.A(KEYINPUT105), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n914), .A2(new_n917), .ZN(new_n918));
  NAND4_X1  g493(.A1(new_n913), .A2(KEYINPUT105), .A3(new_n902), .A4(new_n900), .ZN(new_n919));
  NAND4_X1  g494(.A1(new_n918), .A2(new_n919), .A3(new_n912), .A4(new_n892), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n916), .A2(new_n920), .ZN(new_n921));
  XNOR2_X1  g496(.A(new_n921), .B(KEYINPUT40), .ZN(G395));
  XNOR2_X1  g497(.A(new_n881), .B(new_n625), .ZN(new_n923));
  XNOR2_X1  g498(.A(new_n616), .B(new_n844), .ZN(new_n924));
  XOR2_X1   g499(.A(new_n924), .B(KEYINPUT41), .Z(new_n925));
  AND2_X1   g500(.A1(new_n923), .A2(new_n925), .ZN(new_n926));
  INV_X1    g501(.A(new_n924), .ZN(new_n927));
  NOR2_X1   g502(.A1(new_n923), .A2(new_n927), .ZN(new_n928));
  XNOR2_X1  g503(.A(KEYINPUT106), .B(KEYINPUT42), .ZN(new_n929));
  OR3_X1    g504(.A1(new_n926), .A2(new_n928), .A3(new_n929), .ZN(new_n930));
  XNOR2_X1  g505(.A(new_n729), .B(G305), .ZN(new_n931));
  INV_X1    g506(.A(new_n931), .ZN(new_n932));
  NAND3_X1  g507(.A1(new_n603), .A2(G303), .A3(new_n604), .ZN(new_n933));
  INV_X1    g508(.A(new_n933), .ZN(new_n934));
  AOI21_X1  g509(.A(G303), .B1(new_n603), .B2(new_n604), .ZN(new_n935));
  OAI21_X1  g510(.A(new_n932), .B1(new_n934), .B2(new_n935), .ZN(new_n936));
  INV_X1    g511(.A(new_n935), .ZN(new_n937));
  NAND3_X1  g512(.A1(new_n937), .A2(new_n933), .A3(new_n931), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n936), .A2(new_n938), .ZN(new_n939));
  INV_X1    g514(.A(new_n939), .ZN(new_n940));
  OAI21_X1  g515(.A(new_n929), .B1(new_n926), .B2(new_n928), .ZN(new_n941));
  AND3_X1   g516(.A1(new_n930), .A2(new_n940), .A3(new_n941), .ZN(new_n942));
  AOI21_X1  g517(.A(new_n940), .B1(new_n930), .B2(new_n941), .ZN(new_n943));
  OAI21_X1  g518(.A(G868), .B1(new_n942), .B2(new_n943), .ZN(new_n944));
  INV_X1    g519(.A(new_n887), .ZN(new_n945));
  OAI21_X1  g520(.A(new_n944), .B1(G868), .B2(new_n945), .ZN(G295));
  OAI21_X1  g521(.A(new_n944), .B1(G868), .B2(new_n945), .ZN(G331));
  XNOR2_X1  g522(.A(G168), .B(G171), .ZN(new_n948));
  INV_X1    g523(.A(new_n948), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n881), .A2(new_n949), .ZN(new_n950));
  NAND3_X1  g525(.A1(new_n878), .A2(new_n948), .A3(new_n880), .ZN(new_n951));
  NAND3_X1  g526(.A1(new_n950), .A2(new_n951), .A3(KEYINPUT107), .ZN(new_n952));
  OR3_X1    g527(.A1(new_n881), .A2(new_n949), .A3(KEYINPUT107), .ZN(new_n953));
  NAND3_X1  g528(.A1(new_n925), .A2(new_n952), .A3(new_n953), .ZN(new_n954));
  NAND3_X1  g529(.A1(new_n950), .A2(new_n951), .A3(new_n924), .ZN(new_n955));
  NAND3_X1  g530(.A1(new_n954), .A2(new_n939), .A3(new_n955), .ZN(new_n956));
  INV_X1    g531(.A(G37), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n956), .A2(new_n957), .ZN(new_n958));
  AOI21_X1  g533(.A(new_n939), .B1(new_n954), .B2(new_n955), .ZN(new_n959));
  OAI21_X1  g534(.A(KEYINPUT43), .B1(new_n958), .B2(new_n959), .ZN(new_n960));
  NAND2_X1  g535(.A1(new_n950), .A2(new_n951), .ZN(new_n961));
  AND2_X1   g536(.A1(new_n925), .A2(new_n961), .ZN(new_n962));
  AOI21_X1  g537(.A(new_n927), .B1(new_n952), .B2(new_n953), .ZN(new_n963));
  OAI21_X1  g538(.A(new_n940), .B1(new_n962), .B2(new_n963), .ZN(new_n964));
  INV_X1    g539(.A(KEYINPUT43), .ZN(new_n965));
  NAND4_X1  g540(.A1(new_n964), .A2(new_n965), .A3(new_n957), .A4(new_n956), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n960), .A2(new_n966), .ZN(new_n967));
  OAI21_X1  g542(.A(new_n965), .B1(new_n958), .B2(new_n959), .ZN(new_n968));
  NAND3_X1  g543(.A1(new_n964), .A2(new_n957), .A3(new_n956), .ZN(new_n969));
  OAI21_X1  g544(.A(new_n968), .B1(new_n965), .B2(new_n969), .ZN(new_n970));
  MUX2_X1   g545(.A(new_n967), .B(new_n970), .S(KEYINPUT44), .Z(G397));
  INV_X1    g546(.A(G1384), .ZN(new_n972));
  OAI21_X1  g547(.A(new_n972), .B1(new_n493), .B2(new_n503), .ZN(new_n973));
  INV_X1    g548(.A(KEYINPUT45), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n973), .A2(new_n974), .ZN(new_n975));
  NAND2_X1  g550(.A1(G160), .A2(G40), .ZN(new_n976));
  NOR2_X1   g551(.A1(new_n975), .A2(new_n976), .ZN(new_n977));
  XNOR2_X1  g552(.A(new_n790), .B(new_n796), .ZN(new_n978));
  INV_X1    g553(.A(new_n769), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n979), .A2(G1996), .ZN(new_n980));
  OAI211_X1 g555(.A(new_n978), .B(new_n980), .C1(new_n770), .C2(G1996), .ZN(new_n981));
  XNOR2_X1  g556(.A(new_n708), .B(new_n711), .ZN(new_n982));
  OAI21_X1  g557(.A(new_n977), .B1(new_n981), .B2(new_n982), .ZN(new_n983));
  INV_X1    g558(.A(new_n983), .ZN(new_n984));
  XNOR2_X1  g559(.A(G290), .B(G1986), .ZN(new_n985));
  AOI21_X1  g560(.A(new_n984), .B1(new_n985), .B2(new_n977), .ZN(new_n986));
  INV_X1    g561(.A(G8), .ZN(new_n987));
  AOI22_X1  g562(.A1(new_n470), .A2(KEYINPUT66), .B1(G113), .B2(G2104), .ZN(new_n988));
  AOI21_X1  g563(.A(new_n480), .B1(new_n988), .B2(new_n473), .ZN(new_n989));
  INV_X1    g564(.A(G40), .ZN(new_n990));
  NOR3_X1   g565(.A1(new_n989), .A2(new_n990), .A3(new_n468), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n489), .A2(new_n491), .ZN(new_n992));
  NOR2_X1   g567(.A1(new_n477), .A2(new_n492), .ZN(new_n993));
  NOR2_X1   g568(.A1(new_n992), .A2(new_n993), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n497), .A2(new_n502), .ZN(new_n995));
  INV_X1    g570(.A(new_n494), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n995), .A2(new_n996), .ZN(new_n997));
  AOI21_X1  g572(.A(G1384), .B1(new_n994), .B2(new_n997), .ZN(new_n998));
  AOI21_X1  g573(.A(new_n987), .B1(new_n991), .B2(new_n998), .ZN(new_n999));
  INV_X1    g574(.A(KEYINPUT49), .ZN(new_n1000));
  INV_X1    g575(.A(new_n737), .ZN(new_n1001));
  OAI211_X1 g576(.A(new_n1001), .B(new_n582), .C1(KEYINPUT109), .C2(new_n700), .ZN(new_n1002));
  AOI21_X1  g577(.A(new_n700), .B1(new_n582), .B2(KEYINPUT109), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n1003), .A2(G305), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n1002), .A2(new_n1004), .ZN(new_n1005));
  OAI21_X1  g580(.A(new_n999), .B1(new_n1000), .B2(new_n1005), .ZN(new_n1006));
  NAND3_X1  g581(.A1(new_n1002), .A2(new_n1004), .A3(KEYINPUT110), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n1007), .A2(new_n1000), .ZN(new_n1008));
  AOI21_X1  g583(.A(KEYINPUT110), .B1(new_n1002), .B2(new_n1004), .ZN(new_n1009));
  OAI21_X1  g584(.A(KEYINPUT111), .B1(new_n1008), .B2(new_n1009), .ZN(new_n1010));
  INV_X1    g585(.A(KEYINPUT110), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n1005), .A2(new_n1011), .ZN(new_n1012));
  INV_X1    g587(.A(KEYINPUT111), .ZN(new_n1013));
  NAND4_X1  g588(.A1(new_n1012), .A2(new_n1013), .A3(new_n1000), .A4(new_n1007), .ZN(new_n1014));
  AOI21_X1  g589(.A(new_n1006), .B1(new_n1010), .B2(new_n1014), .ZN(new_n1015));
  NAND2_X1  g590(.A1(new_n991), .A2(new_n998), .ZN(new_n1016));
  NAND3_X1  g591(.A1(new_n727), .A2(G1976), .A3(new_n728), .ZN(new_n1017));
  NAND3_X1  g592(.A1(new_n1016), .A2(G8), .A3(new_n1017), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n1018), .A2(KEYINPUT52), .ZN(new_n1019));
  XNOR2_X1  g594(.A(KEYINPUT108), .B(G1976), .ZN(new_n1020));
  AOI21_X1  g595(.A(KEYINPUT52), .B1(G288), .B2(new_n1020), .ZN(new_n1021));
  NAND3_X1  g596(.A1(new_n999), .A2(new_n1017), .A3(new_n1021), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n1019), .A2(new_n1022), .ZN(new_n1023));
  NOR3_X1   g598(.A1(new_n1015), .A2(new_n1023), .A3(KEYINPUT112), .ZN(new_n1024));
  INV_X1    g599(.A(KEYINPUT55), .ZN(new_n1025));
  AOI21_X1  g600(.A(new_n1025), .B1(G303), .B2(G8), .ZN(new_n1026));
  NOR3_X1   g601(.A1(G166), .A2(KEYINPUT55), .A3(new_n987), .ZN(new_n1027));
  NOR2_X1   g602(.A1(new_n1026), .A2(new_n1027), .ZN(new_n1028));
  INV_X1    g603(.A(new_n1028), .ZN(new_n1029));
  INV_X1    g604(.A(KEYINPUT50), .ZN(new_n1030));
  NAND2_X1  g605(.A1(new_n994), .A2(new_n997), .ZN(new_n1031));
  AOI21_X1  g606(.A(new_n1030), .B1(new_n1031), .B2(new_n972), .ZN(new_n1032));
  NOR2_X1   g607(.A1(KEYINPUT50), .A2(G1384), .ZN(new_n1033));
  OAI21_X1  g608(.A(new_n1033), .B1(new_n493), .B2(new_n503), .ZN(new_n1034));
  NAND3_X1  g609(.A1(new_n1034), .A2(G40), .A3(G160), .ZN(new_n1035));
  NOR2_X1   g610(.A1(new_n1032), .A2(new_n1035), .ZN(new_n1036));
  OAI211_X1 g611(.A(KEYINPUT45), .B(new_n972), .C1(new_n493), .C2(new_n503), .ZN(new_n1037));
  NAND3_X1  g612(.A1(new_n975), .A2(new_n991), .A3(new_n1037), .ZN(new_n1038));
  INV_X1    g613(.A(G1971), .ZN(new_n1039));
  AOI22_X1  g614(.A1(new_n1036), .A2(new_n779), .B1(new_n1038), .B2(new_n1039), .ZN(new_n1040));
  OAI21_X1  g615(.A(new_n1029), .B1(new_n1040), .B2(new_n987), .ZN(new_n1041));
  AOI21_X1  g616(.A(new_n976), .B1(new_n974), .B2(new_n973), .ZN(new_n1042));
  AOI21_X1  g617(.A(G1971), .B1(new_n1042), .B2(new_n1037), .ZN(new_n1043));
  OAI211_X1 g618(.A(new_n991), .B(new_n1034), .C1(new_n998), .C2(new_n1030), .ZN(new_n1044));
  NOR2_X1   g619(.A1(new_n1044), .A2(G2090), .ZN(new_n1045));
  OAI211_X1 g620(.A(G8), .B(new_n1028), .C1(new_n1043), .C2(new_n1045), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n1041), .A2(new_n1046), .ZN(new_n1047));
  NOR2_X1   g622(.A1(new_n1024), .A2(new_n1047), .ZN(new_n1048));
  OAI21_X1  g623(.A(KEYINPUT112), .B1(new_n1015), .B2(new_n1023), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n1048), .A2(new_n1049), .ZN(new_n1050));
  NAND2_X1  g625(.A1(new_n973), .A2(KEYINPUT50), .ZN(new_n1051));
  XOR2_X1   g626(.A(KEYINPUT113), .B(G2084), .Z(new_n1052));
  NAND4_X1  g627(.A1(new_n1051), .A2(new_n991), .A3(new_n1034), .A4(new_n1052), .ZN(new_n1053));
  INV_X1    g628(.A(KEYINPUT114), .ZN(new_n1054));
  NAND2_X1  g629(.A1(new_n1053), .A2(new_n1054), .ZN(new_n1055));
  AND3_X1   g630(.A1(new_n1034), .A2(G40), .A3(G160), .ZN(new_n1056));
  NAND4_X1  g631(.A1(new_n1056), .A2(KEYINPUT114), .A3(new_n1051), .A4(new_n1052), .ZN(new_n1057));
  NAND2_X1  g632(.A1(new_n1038), .A2(new_n805), .ZN(new_n1058));
  NAND3_X1  g633(.A1(new_n1055), .A2(new_n1057), .A3(new_n1058), .ZN(new_n1059));
  NAND3_X1  g634(.A1(new_n1059), .A2(G8), .A3(G168), .ZN(new_n1060));
  NOR3_X1   g635(.A1(new_n1050), .A2(KEYINPUT63), .A3(new_n1060), .ZN(new_n1061));
  NOR2_X1   g636(.A1(new_n1015), .A2(new_n1023), .ZN(new_n1062));
  AND3_X1   g637(.A1(new_n1059), .A2(G8), .A3(G168), .ZN(new_n1063));
  NAND3_X1  g638(.A1(new_n1062), .A2(new_n1063), .A3(new_n1041), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n1064), .A2(KEYINPUT63), .ZN(new_n1065));
  OR2_X1    g640(.A1(G288), .A2(G1976), .ZN(new_n1066));
  OAI22_X1  g641(.A1(new_n1015), .A2(new_n1066), .B1(G1981), .B2(G305), .ZN(new_n1067));
  INV_X1    g642(.A(new_n1046), .ZN(new_n1068));
  AOI22_X1  g643(.A1(new_n1067), .A2(new_n999), .B1(new_n1062), .B2(new_n1068), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n1065), .A2(new_n1069), .ZN(new_n1070));
  NOR2_X1   g645(.A1(new_n1061), .A2(new_n1070), .ZN(new_n1071));
  AOI21_X1  g646(.A(KEYINPUT119), .B1(new_n608), .B2(new_n615), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n1044), .A2(new_n802), .ZN(new_n1073));
  NAND3_X1  g648(.A1(new_n991), .A2(new_n998), .A3(new_n796), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n1073), .A2(new_n1074), .ZN(new_n1075));
  INV_X1    g650(.A(KEYINPUT60), .ZN(new_n1076));
  OAI21_X1  g651(.A(new_n1072), .B1(new_n1075), .B2(new_n1076), .ZN(new_n1077));
  AND3_X1   g652(.A1(new_n608), .A2(KEYINPUT119), .A3(new_n615), .ZN(new_n1078));
  NOR2_X1   g653(.A1(new_n1078), .A2(new_n1072), .ZN(new_n1079));
  NAND4_X1  g654(.A1(new_n1079), .A2(new_n1074), .A3(KEYINPUT60), .A4(new_n1073), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1075), .A2(new_n1076), .ZN(new_n1081));
  NAND3_X1  g656(.A1(new_n1077), .A2(new_n1080), .A3(new_n1081), .ZN(new_n1082));
  NAND2_X1  g657(.A1(KEYINPUT118), .A2(KEYINPUT59), .ZN(new_n1083));
  XOR2_X1   g658(.A(KEYINPUT58), .B(G1341), .Z(new_n1084));
  NAND2_X1  g659(.A1(new_n1016), .A2(new_n1084), .ZN(new_n1085));
  INV_X1    g660(.A(G1996), .ZN(new_n1086));
  NAND4_X1  g661(.A1(new_n975), .A2(new_n1086), .A3(new_n991), .A4(new_n1037), .ZN(new_n1087));
  AOI211_X1 g662(.A(new_n549), .B(new_n1083), .C1(new_n1085), .C2(new_n1087), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n1085), .A2(new_n1087), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n1089), .A2(new_n550), .ZN(new_n1090));
  XOR2_X1   g665(.A(KEYINPUT118), .B(KEYINPUT59), .Z(new_n1091));
  AOI21_X1  g666(.A(new_n1088), .B1(new_n1090), .B2(new_n1091), .ZN(new_n1092));
  NAND2_X1  g667(.A1(G299), .A2(KEYINPUT57), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n564), .A2(new_n565), .ZN(new_n1094));
  INV_X1    g669(.A(KEYINPUT116), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n1094), .A2(new_n1095), .ZN(new_n1096));
  NAND3_X1  g671(.A1(new_n564), .A2(KEYINPUT116), .A3(new_n565), .ZN(new_n1097));
  NAND4_X1  g672(.A1(new_n1096), .A2(new_n567), .A3(new_n559), .A4(new_n1097), .ZN(new_n1098));
  AOI21_X1  g673(.A(new_n1093), .B1(new_n1098), .B2(KEYINPUT115), .ZN(new_n1099));
  INV_X1    g674(.A(KEYINPUT115), .ZN(new_n1100));
  AOI21_X1  g675(.A(KEYINPUT57), .B1(new_n1098), .B2(new_n1100), .ZN(new_n1101));
  NOR2_X1   g676(.A1(new_n1099), .A2(new_n1101), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n1044), .A2(new_n846), .ZN(new_n1103));
  XNOR2_X1  g678(.A(KEYINPUT56), .B(G2072), .ZN(new_n1104));
  NAND3_X1  g679(.A1(new_n1042), .A2(new_n1037), .A3(new_n1104), .ZN(new_n1105));
  AOI21_X1  g680(.A(new_n1102), .B1(new_n1103), .B2(new_n1105), .ZN(new_n1106));
  NAND3_X1  g681(.A1(new_n1102), .A2(new_n1105), .A3(new_n1103), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n1107), .A2(KEYINPUT61), .ZN(new_n1108));
  OAI211_X1 g683(.A(new_n1082), .B(new_n1092), .C1(new_n1106), .C2(new_n1108), .ZN(new_n1109));
  AOI21_X1  g684(.A(new_n1106), .B1(new_n617), .B2(new_n1075), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n1109), .A2(new_n1110), .ZN(new_n1111));
  XOR2_X1   g686(.A(new_n1107), .B(KEYINPUT117), .Z(new_n1112));
  NAND2_X1  g687(.A1(new_n1111), .A2(new_n1112), .ZN(new_n1113));
  INV_X1    g688(.A(KEYINPUT61), .ZN(new_n1114));
  OR2_X1    g689(.A1(new_n1109), .A2(new_n1114), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n1113), .A2(new_n1115), .ZN(new_n1116));
  OAI21_X1  g691(.A(KEYINPUT54), .B1(G301), .B2(KEYINPUT122), .ZN(new_n1117));
  INV_X1    g692(.A(new_n1117), .ZN(new_n1118));
  NAND4_X1  g693(.A1(new_n1042), .A2(KEYINPUT53), .A3(new_n810), .A4(new_n1037), .ZN(new_n1119));
  NAND4_X1  g694(.A1(new_n975), .A2(new_n810), .A3(new_n991), .A4(new_n1037), .ZN(new_n1120));
  INV_X1    g695(.A(KEYINPUT53), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n1120), .A2(new_n1121), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n1044), .A2(new_n831), .ZN(new_n1123));
  AND4_X1   g698(.A1(G301), .A2(new_n1119), .A3(new_n1122), .A4(new_n1123), .ZN(new_n1124));
  AOI22_X1  g699(.A1(new_n1120), .A2(new_n1121), .B1(new_n1044), .B2(new_n831), .ZN(new_n1125));
  AOI21_X1  g700(.A(G301), .B1(new_n1125), .B2(new_n1119), .ZN(new_n1126));
  OAI21_X1  g701(.A(new_n1118), .B1(new_n1124), .B2(new_n1126), .ZN(new_n1127));
  NAND3_X1  g702(.A1(new_n1119), .A2(new_n1122), .A3(new_n1123), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n1128), .A2(G171), .ZN(new_n1129));
  NAND3_X1  g704(.A1(new_n1125), .A2(G301), .A3(new_n1119), .ZN(new_n1130));
  NAND3_X1  g705(.A1(new_n1129), .A2(new_n1117), .A3(new_n1130), .ZN(new_n1131));
  NAND2_X1  g706(.A1(new_n1127), .A2(new_n1131), .ZN(new_n1132));
  NAND3_X1  g707(.A1(new_n1132), .A2(new_n1048), .A3(new_n1049), .ZN(new_n1133));
  INV_X1    g708(.A(KEYINPUT121), .ZN(new_n1134));
  NOR2_X1   g709(.A1(G168), .A2(new_n987), .ZN(new_n1135));
  INV_X1    g710(.A(KEYINPUT51), .ZN(new_n1136));
  AOI21_X1  g711(.A(new_n1135), .B1(KEYINPUT120), .B2(new_n1136), .ZN(new_n1137));
  AOI21_X1  g712(.A(new_n1137), .B1(new_n1059), .B2(G8), .ZN(new_n1138));
  NOR2_X1   g713(.A1(new_n1063), .A2(new_n1138), .ZN(new_n1139));
  NAND3_X1  g714(.A1(new_n1059), .A2(KEYINPUT120), .A3(G8), .ZN(new_n1140));
  INV_X1    g715(.A(new_n1135), .ZN(new_n1141));
  AOI21_X1  g716(.A(KEYINPUT51), .B1(new_n1140), .B2(new_n1141), .ZN(new_n1142));
  OAI21_X1  g717(.A(new_n1134), .B1(new_n1139), .B2(new_n1142), .ZN(new_n1143));
  AOI22_X1  g718(.A1(new_n1054), .A2(new_n1053), .B1(new_n1038), .B2(new_n805), .ZN(new_n1144));
  AOI21_X1  g719(.A(new_n987), .B1(new_n1144), .B2(new_n1057), .ZN(new_n1145));
  OAI21_X1  g720(.A(new_n1060), .B1(new_n1145), .B2(new_n1137), .ZN(new_n1146));
  AOI21_X1  g721(.A(new_n1135), .B1(new_n1145), .B2(KEYINPUT120), .ZN(new_n1147));
  OAI211_X1 g722(.A(new_n1146), .B(KEYINPUT121), .C1(new_n1147), .C2(KEYINPUT51), .ZN(new_n1148));
  AOI21_X1  g723(.A(new_n1133), .B1(new_n1143), .B2(new_n1148), .ZN(new_n1149));
  OAI21_X1  g724(.A(new_n1116), .B1(new_n1149), .B2(KEYINPUT123), .ZN(new_n1150));
  INV_X1    g725(.A(KEYINPUT123), .ZN(new_n1151));
  AOI211_X1 g726(.A(new_n1151), .B(new_n1133), .C1(new_n1143), .C2(new_n1148), .ZN(new_n1152));
  OAI21_X1  g727(.A(new_n1071), .B1(new_n1150), .B2(new_n1152), .ZN(new_n1153));
  INV_X1    g728(.A(KEYINPUT62), .ZN(new_n1154));
  NAND3_X1  g729(.A1(new_n1143), .A2(new_n1154), .A3(new_n1148), .ZN(new_n1155));
  NOR2_X1   g730(.A1(new_n1050), .A2(new_n1129), .ZN(new_n1156));
  AND3_X1   g731(.A1(new_n1155), .A2(new_n1156), .A3(KEYINPUT124), .ZN(new_n1157));
  AOI21_X1  g732(.A(KEYINPUT124), .B1(new_n1155), .B2(new_n1156), .ZN(new_n1158));
  AOI21_X1  g733(.A(new_n1154), .B1(new_n1143), .B2(new_n1148), .ZN(new_n1159));
  NOR3_X1   g734(.A1(new_n1157), .A2(new_n1158), .A3(new_n1159), .ZN(new_n1160));
  OAI21_X1  g735(.A(new_n986), .B1(new_n1153), .B2(new_n1160), .ZN(new_n1161));
  INV_X1    g736(.A(new_n977), .ZN(new_n1162));
  AOI21_X1  g737(.A(new_n1162), .B1(new_n978), .B2(new_n769), .ZN(new_n1163));
  INV_X1    g738(.A(KEYINPUT46), .ZN(new_n1164));
  NOR3_X1   g739(.A1(new_n1162), .A2(new_n1164), .A3(G1996), .ZN(new_n1165));
  AOI21_X1  g740(.A(KEYINPUT46), .B1(new_n977), .B2(new_n1086), .ZN(new_n1166));
  NOR3_X1   g741(.A1(new_n1163), .A2(new_n1165), .A3(new_n1166), .ZN(new_n1167));
  XNOR2_X1  g742(.A(new_n1167), .B(KEYINPUT47), .ZN(new_n1168));
  INV_X1    g743(.A(KEYINPUT48), .ZN(new_n1169));
  NAND3_X1  g744(.A1(new_n716), .A2(new_n695), .A3(new_n977), .ZN(new_n1170));
  AOI21_X1  g745(.A(new_n984), .B1(new_n1169), .B2(new_n1170), .ZN(new_n1171));
  OAI21_X1  g746(.A(new_n1171), .B1(new_n1169), .B2(new_n1170), .ZN(new_n1172));
  NOR2_X1   g747(.A1(new_n790), .A2(G2067), .ZN(new_n1173));
  NAND2_X1  g748(.A1(new_n981), .A2(new_n977), .ZN(new_n1174));
  INV_X1    g749(.A(new_n711), .ZN(new_n1175));
  NOR2_X1   g750(.A1(new_n709), .A2(new_n1175), .ZN(new_n1176));
  AOI21_X1  g751(.A(new_n1173), .B1(new_n1174), .B2(new_n1176), .ZN(new_n1177));
  NOR2_X1   g752(.A1(new_n1177), .A2(new_n1162), .ZN(new_n1178));
  OAI21_X1  g753(.A(new_n1172), .B1(KEYINPUT125), .B2(new_n1178), .ZN(new_n1179));
  AOI211_X1 g754(.A(new_n1168), .B(new_n1179), .C1(KEYINPUT125), .C2(new_n1178), .ZN(new_n1180));
  NAND2_X1  g755(.A1(new_n1161), .A2(new_n1180), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g756(.A1(G227), .A2(new_n458), .ZN(new_n1183));
  INV_X1    g757(.A(new_n1183), .ZN(new_n1184));
  OAI21_X1  g758(.A(KEYINPUT126), .B1(G401), .B2(new_n1184), .ZN(new_n1185));
  AND2_X1   g759(.A1(new_n659), .A2(G14), .ZN(new_n1186));
  AOI21_X1  g760(.A(KEYINPUT81), .B1(new_n665), .B2(new_n656), .ZN(new_n1187));
  AOI211_X1 g761(.A(new_n661), .B(new_n657), .C1(new_n655), .C2(new_n658), .ZN(new_n1188));
  OAI21_X1  g762(.A(new_n1186), .B1(new_n1187), .B2(new_n1188), .ZN(new_n1189));
  INV_X1    g763(.A(KEYINPUT126), .ZN(new_n1190));
  NAND3_X1  g764(.A1(new_n1189), .A2(new_n1190), .A3(new_n1183), .ZN(new_n1191));
  NAND3_X1  g765(.A1(new_n1185), .A2(new_n1191), .A3(new_n702), .ZN(new_n1192));
  AOI21_X1  g766(.A(new_n1192), .B1(new_n916), .B2(new_n920), .ZN(new_n1193));
  INV_X1    g767(.A(KEYINPUT127), .ZN(new_n1194));
  AND3_X1   g768(.A1(new_n1193), .A2(new_n967), .A3(new_n1194), .ZN(new_n1195));
  AOI21_X1  g769(.A(new_n1194), .B1(new_n1193), .B2(new_n967), .ZN(new_n1196));
  NOR2_X1   g770(.A1(new_n1195), .A2(new_n1196), .ZN(G308));
  NAND2_X1  g771(.A1(new_n1193), .A2(new_n967), .ZN(new_n1198));
  NAND2_X1  g772(.A1(new_n1198), .A2(KEYINPUT127), .ZN(new_n1199));
  NAND3_X1  g773(.A1(new_n1193), .A2(new_n967), .A3(new_n1194), .ZN(new_n1200));
  NAND2_X1  g774(.A1(new_n1199), .A2(new_n1200), .ZN(G225));
endmodule


