//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 0 0 0 1 1 0 0 0 1 0 0 0 1 1 0 1 1 0 0 0 0 0 1 0 0 1 0 1 0 1 0 0 0 1 0 0 1 1 1 0 1 1 1 1 1 0 1 1 0 1 0 0 1 0 1 0 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:27:27 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n616, new_n617, new_n618, new_n619, new_n620, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n627, new_n628, new_n629, new_n630,
    new_n631, new_n632, new_n634, new_n635, new_n636, new_n637, new_n638,
    new_n639, new_n640, new_n641, new_n642, new_n643, new_n644, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n694, new_n696, new_n697, new_n698, new_n699,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n705, new_n707,
    new_n708, new_n709, new_n710, new_n711, new_n712, new_n713, new_n714,
    new_n715, new_n716, new_n717, new_n719, new_n720, new_n721, new_n722,
    new_n723, new_n724, new_n725, new_n726, new_n727, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n748, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n782,
    new_n783, new_n784, new_n785, new_n786, new_n787, new_n788, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n926, new_n927,
    new_n928, new_n929, new_n930, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n945, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n984, new_n985, new_n986, new_n987,
    new_n988, new_n989, new_n990, new_n991, new_n992, new_n993, new_n994,
    new_n995;
  INV_X1    g000(.A(G221), .ZN(new_n187));
  XOR2_X1   g001(.A(KEYINPUT9), .B(G234), .Z(new_n188));
  INV_X1    g002(.A(G902), .ZN(new_n189));
  AOI21_X1  g003(.A(new_n187), .B1(new_n188), .B2(new_n189), .ZN(new_n190));
  INV_X1    g004(.A(new_n190), .ZN(new_n191));
  OAI21_X1  g005(.A(G214), .B1(G237), .B2(G902), .ZN(new_n192));
  INV_X1    g006(.A(G113), .ZN(new_n193));
  XOR2_X1   g007(.A(KEYINPUT78), .B(KEYINPUT5), .Z(new_n194));
  INV_X1    g008(.A(G116), .ZN(new_n195));
  NOR2_X1   g009(.A1(new_n195), .A2(G119), .ZN(new_n196));
  AOI21_X1  g010(.A(new_n193), .B1(new_n194), .B2(new_n196), .ZN(new_n197));
  INV_X1    g011(.A(KEYINPUT65), .ZN(new_n198));
  INV_X1    g012(.A(G119), .ZN(new_n199));
  OAI21_X1  g013(.A(new_n198), .B1(new_n199), .B2(G116), .ZN(new_n200));
  NAND3_X1  g014(.A1(new_n195), .A2(KEYINPUT65), .A3(G119), .ZN(new_n201));
  AOI21_X1  g015(.A(new_n196), .B1(new_n200), .B2(new_n201), .ZN(new_n202));
  INV_X1    g016(.A(new_n202), .ZN(new_n203));
  OAI21_X1  g017(.A(new_n197), .B1(new_n203), .B2(new_n194), .ZN(new_n204));
  XOR2_X1   g018(.A(KEYINPUT2), .B(G113), .Z(new_n205));
  NAND2_X1  g019(.A1(new_n202), .A2(new_n205), .ZN(new_n206));
  INV_X1    g020(.A(G104), .ZN(new_n207));
  OAI21_X1  g021(.A(KEYINPUT3), .B1(new_n207), .B2(G107), .ZN(new_n208));
  INV_X1    g022(.A(KEYINPUT3), .ZN(new_n209));
  INV_X1    g023(.A(G107), .ZN(new_n210));
  NAND3_X1  g024(.A1(new_n209), .A2(new_n210), .A3(G104), .ZN(new_n211));
  INV_X1    g025(.A(G101), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n207), .A2(G107), .ZN(new_n213));
  NAND4_X1  g027(.A1(new_n208), .A2(new_n211), .A3(new_n212), .A4(new_n213), .ZN(new_n214));
  NOR2_X1   g028(.A1(new_n207), .A2(G107), .ZN(new_n215));
  NOR2_X1   g029(.A1(new_n210), .A2(G104), .ZN(new_n216));
  OAI21_X1  g030(.A(G101), .B1(new_n215), .B2(new_n216), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n214), .A2(new_n217), .ZN(new_n218));
  NAND3_X1  g032(.A1(new_n204), .A2(new_n206), .A3(new_n218), .ZN(new_n219));
  XNOR2_X1  g033(.A(G110), .B(G122), .ZN(new_n220));
  XNOR2_X1  g034(.A(new_n220), .B(KEYINPUT8), .ZN(new_n221));
  INV_X1    g035(.A(new_n206), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n202), .A2(KEYINPUT5), .ZN(new_n223));
  AOI21_X1  g037(.A(new_n222), .B1(new_n197), .B2(new_n223), .ZN(new_n224));
  OAI211_X1 g038(.A(new_n219), .B(new_n221), .C1(new_n224), .C2(new_n218), .ZN(new_n225));
  INV_X1    g039(.A(G146), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n226), .A2(G143), .ZN(new_n227));
  INV_X1    g041(.A(G143), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n228), .A2(G146), .ZN(new_n229));
  NAND4_X1  g043(.A1(new_n227), .A2(new_n229), .A3(KEYINPUT0), .A4(G128), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n227), .A2(new_n229), .ZN(new_n231));
  INV_X1    g045(.A(new_n231), .ZN(new_n232));
  XNOR2_X1  g046(.A(KEYINPUT0), .B(G128), .ZN(new_n233));
  OAI211_X1 g047(.A(new_n230), .B(G125), .C1(new_n232), .C2(new_n233), .ZN(new_n234));
  INV_X1    g048(.A(KEYINPUT1), .ZN(new_n235));
  NAND4_X1  g049(.A1(new_n227), .A2(new_n229), .A3(new_n235), .A4(G128), .ZN(new_n236));
  INV_X1    g050(.A(new_n236), .ZN(new_n237));
  OAI21_X1  g051(.A(KEYINPUT1), .B1(new_n228), .B2(G146), .ZN(new_n238));
  AOI22_X1  g052(.A1(new_n238), .A2(G128), .B1(new_n227), .B2(new_n229), .ZN(new_n239));
  NOR2_X1   g053(.A1(new_n237), .A2(new_n239), .ZN(new_n240));
  OAI21_X1  g054(.A(new_n234), .B1(new_n240), .B2(G125), .ZN(new_n241));
  INV_X1    g055(.A(KEYINPUT79), .ZN(new_n242));
  INV_X1    g056(.A(G224), .ZN(new_n243));
  NOR2_X1   g057(.A1(new_n243), .A2(G953), .ZN(new_n244));
  INV_X1    g058(.A(new_n244), .ZN(new_n245));
  NAND4_X1  g059(.A1(new_n241), .A2(new_n242), .A3(KEYINPUT7), .A4(new_n245), .ZN(new_n246));
  INV_X1    g060(.A(new_n234), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n238), .A2(G128), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n248), .A2(new_n231), .ZN(new_n249));
  AOI21_X1  g063(.A(G125), .B1(new_n249), .B2(new_n236), .ZN(new_n250));
  OAI211_X1 g064(.A(KEYINPUT7), .B(new_n245), .C1(new_n247), .C2(new_n250), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n251), .A2(KEYINPUT79), .ZN(new_n252));
  AND3_X1   g066(.A1(new_n225), .A2(new_n246), .A3(new_n252), .ZN(new_n253));
  INV_X1    g067(.A(new_n218), .ZN(new_n254));
  NAND3_X1  g068(.A1(new_n204), .A2(new_n206), .A3(new_n254), .ZN(new_n255));
  NAND3_X1  g069(.A1(new_n208), .A2(new_n211), .A3(new_n213), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n256), .A2(G101), .ZN(new_n257));
  NAND3_X1  g071(.A1(new_n257), .A2(KEYINPUT4), .A3(new_n214), .ZN(new_n258));
  INV_X1    g072(.A(new_n258), .ZN(new_n259));
  INV_X1    g073(.A(KEYINPUT4), .ZN(new_n260));
  NAND3_X1  g074(.A1(new_n256), .A2(new_n260), .A3(G101), .ZN(new_n261));
  NOR2_X1   g075(.A1(new_n202), .A2(new_n205), .ZN(new_n262));
  OAI21_X1  g076(.A(new_n261), .B1(new_n222), .B2(new_n262), .ZN(new_n263));
  OAI211_X1 g077(.A(new_n255), .B(new_n220), .C1(new_n259), .C2(new_n263), .ZN(new_n264));
  AND2_X1   g078(.A1(new_n245), .A2(KEYINPUT7), .ZN(new_n265));
  OR2_X1    g079(.A1(new_n241), .A2(new_n265), .ZN(new_n266));
  AND2_X1   g080(.A1(new_n264), .A2(new_n266), .ZN(new_n267));
  AOI21_X1  g081(.A(G902), .B1(new_n253), .B2(new_n267), .ZN(new_n268));
  OAI21_X1  g082(.A(new_n255), .B1(new_n259), .B2(new_n263), .ZN(new_n269));
  INV_X1    g083(.A(new_n220), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  NAND3_X1  g085(.A1(new_n271), .A2(KEYINPUT6), .A3(new_n264), .ZN(new_n272));
  XNOR2_X1  g086(.A(new_n241), .B(new_n245), .ZN(new_n273));
  INV_X1    g087(.A(KEYINPUT6), .ZN(new_n274));
  NAND3_X1  g088(.A1(new_n269), .A2(new_n274), .A3(new_n270), .ZN(new_n275));
  NAND3_X1  g089(.A1(new_n272), .A2(new_n273), .A3(new_n275), .ZN(new_n276));
  OAI21_X1  g090(.A(G210), .B1(G237), .B2(G902), .ZN(new_n277));
  XNOR2_X1  g091(.A(new_n277), .B(KEYINPUT80), .ZN(new_n278));
  INV_X1    g092(.A(new_n278), .ZN(new_n279));
  AND3_X1   g093(.A1(new_n268), .A2(new_n276), .A3(new_n279), .ZN(new_n280));
  AOI21_X1  g094(.A(new_n279), .B1(new_n268), .B2(new_n276), .ZN(new_n281));
  OAI21_X1  g095(.A(new_n192), .B1(new_n280), .B2(new_n281), .ZN(new_n282));
  INV_X1    g096(.A(KEYINPUT81), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n268), .A2(new_n276), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n285), .A2(new_n278), .ZN(new_n286));
  NAND3_X1  g100(.A1(new_n268), .A2(new_n276), .A3(new_n279), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  NAND3_X1  g102(.A1(new_n288), .A2(KEYINPUT81), .A3(new_n192), .ZN(new_n289));
  AND3_X1   g103(.A1(new_n249), .A2(KEYINPUT67), .A3(new_n236), .ZN(new_n290));
  AOI21_X1  g104(.A(KEYINPUT67), .B1(new_n249), .B2(new_n236), .ZN(new_n291));
  OAI211_X1 g105(.A(KEYINPUT10), .B(new_n254), .C1(new_n290), .C2(new_n291), .ZN(new_n292));
  INV_X1    g106(.A(KEYINPUT66), .ZN(new_n293));
  INV_X1    g107(.A(G131), .ZN(new_n294));
  INV_X1    g108(.A(G137), .ZN(new_n295));
  AOI21_X1  g109(.A(KEYINPUT11), .B1(new_n295), .B2(G134), .ZN(new_n296));
  NOR2_X1   g110(.A1(new_n295), .A2(G134), .ZN(new_n297));
  NOR2_X1   g111(.A1(new_n296), .A2(new_n297), .ZN(new_n298));
  NAND3_X1  g112(.A1(new_n295), .A2(KEYINPUT11), .A3(G134), .ZN(new_n299));
  AOI21_X1  g113(.A(new_n294), .B1(new_n298), .B2(new_n299), .ZN(new_n300));
  INV_X1    g114(.A(KEYINPUT11), .ZN(new_n301));
  INV_X1    g115(.A(G134), .ZN(new_n302));
  OAI21_X1  g116(.A(new_n301), .B1(new_n302), .B2(G137), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n302), .A2(G137), .ZN(new_n304));
  NAND4_X1  g118(.A1(new_n303), .A2(new_n299), .A3(new_n294), .A4(new_n304), .ZN(new_n305));
  INV_X1    g119(.A(new_n305), .ZN(new_n306));
  OAI21_X1  g120(.A(new_n293), .B1(new_n300), .B2(new_n306), .ZN(new_n307));
  NAND3_X1  g121(.A1(new_n303), .A2(new_n299), .A3(new_n304), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n308), .A2(G131), .ZN(new_n309));
  NAND3_X1  g123(.A1(new_n309), .A2(KEYINPUT66), .A3(new_n305), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n307), .A2(new_n310), .ZN(new_n311));
  OAI21_X1  g125(.A(new_n230), .B1(new_n232), .B2(new_n233), .ZN(new_n312));
  INV_X1    g126(.A(new_n312), .ZN(new_n313));
  NAND3_X1  g127(.A1(new_n313), .A2(new_n258), .A3(new_n261), .ZN(new_n314));
  OAI211_X1 g128(.A(new_n214), .B(new_n217), .C1(new_n237), .C2(new_n239), .ZN(new_n315));
  INV_X1    g129(.A(KEYINPUT10), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n315), .A2(new_n316), .ZN(new_n317));
  NAND4_X1  g131(.A1(new_n292), .A2(new_n311), .A3(new_n314), .A4(new_n317), .ZN(new_n318));
  XNOR2_X1  g132(.A(G110), .B(G140), .ZN(new_n319));
  INV_X1    g133(.A(G953), .ZN(new_n320));
  AND2_X1   g134(.A1(new_n320), .A2(G227), .ZN(new_n321));
  XNOR2_X1  g135(.A(new_n319), .B(new_n321), .ZN(new_n322));
  INV_X1    g136(.A(new_n322), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n318), .A2(new_n323), .ZN(new_n324));
  INV_X1    g138(.A(KEYINPUT77), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n324), .A2(new_n325), .ZN(new_n326));
  NAND3_X1  g140(.A1(new_n292), .A2(new_n317), .A3(new_n314), .ZN(new_n327));
  INV_X1    g141(.A(new_n310), .ZN(new_n328));
  AOI21_X1  g142(.A(KEYINPUT66), .B1(new_n309), .B2(new_n305), .ZN(new_n329));
  NOR2_X1   g143(.A1(new_n328), .A2(new_n329), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n327), .A2(new_n330), .ZN(new_n331));
  NAND3_X1  g145(.A1(new_n318), .A2(KEYINPUT77), .A3(new_n323), .ZN(new_n332));
  NAND3_X1  g146(.A1(new_n326), .A2(new_n331), .A3(new_n332), .ZN(new_n333));
  INV_X1    g147(.A(new_n318), .ZN(new_n334));
  INV_X1    g148(.A(KEYINPUT12), .ZN(new_n335));
  NAND3_X1  g149(.A1(new_n218), .A2(new_n236), .A3(new_n249), .ZN(new_n336));
  AND2_X1   g150(.A1(new_n336), .A2(new_n315), .ZN(new_n337));
  OAI21_X1  g151(.A(new_n335), .B1(new_n337), .B2(new_n311), .ZN(new_n338));
  INV_X1    g152(.A(KEYINPUT76), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n338), .A2(new_n339), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n336), .A2(new_n315), .ZN(new_n341));
  NAND3_X1  g155(.A1(new_n341), .A2(new_n310), .A3(new_n307), .ZN(new_n342));
  NAND3_X1  g156(.A1(new_n342), .A2(KEYINPUT76), .A3(new_n335), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n340), .A2(new_n343), .ZN(new_n344));
  OAI211_X1 g158(.A(new_n341), .B(KEYINPUT12), .C1(new_n300), .C2(new_n306), .ZN(new_n345));
  AOI21_X1  g159(.A(new_n334), .B1(new_n344), .B2(new_n345), .ZN(new_n346));
  XOR2_X1   g160(.A(new_n322), .B(KEYINPUT75), .Z(new_n347));
  INV_X1    g161(.A(new_n347), .ZN(new_n348));
  OAI211_X1 g162(.A(G469), .B(new_n333), .C1(new_n346), .C2(new_n348), .ZN(new_n349));
  INV_X1    g163(.A(G469), .ZN(new_n350));
  AOI21_X1  g164(.A(new_n324), .B1(new_n344), .B2(new_n345), .ZN(new_n351));
  AOI21_X1  g165(.A(new_n323), .B1(new_n331), .B2(new_n318), .ZN(new_n352));
  OAI211_X1 g166(.A(new_n350), .B(new_n189), .C1(new_n351), .C2(new_n352), .ZN(new_n353));
  NAND2_X1  g167(.A1(G469), .A2(G902), .ZN(new_n354));
  NAND3_X1  g168(.A1(new_n349), .A2(new_n353), .A3(new_n354), .ZN(new_n355));
  AND4_X1   g169(.A1(new_n191), .A2(new_n284), .A3(new_n289), .A4(new_n355), .ZN(new_n356));
  INV_X1    g170(.A(G475), .ZN(new_n357));
  XNOR2_X1  g171(.A(G125), .B(G140), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n358), .A2(KEYINPUT16), .ZN(new_n359));
  INV_X1    g173(.A(G140), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n360), .A2(G125), .ZN(new_n361));
  OR2_X1    g175(.A1(new_n361), .A2(KEYINPUT16), .ZN(new_n362));
  NAND3_X1  g176(.A1(new_n359), .A2(G146), .A3(new_n362), .ZN(new_n363));
  INV_X1    g177(.A(new_n363), .ZN(new_n364));
  AOI21_X1  g178(.A(G146), .B1(new_n359), .B2(new_n362), .ZN(new_n365));
  OR3_X1    g179(.A1(new_n364), .A2(new_n365), .A3(KEYINPUT85), .ZN(new_n366));
  NOR2_X1   g180(.A1(G237), .A2(G953), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n367), .A2(G214), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n368), .A2(new_n228), .ZN(new_n369));
  NAND3_X1  g183(.A1(new_n367), .A2(G143), .A3(G214), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n369), .A2(new_n370), .ZN(new_n371));
  NOR2_X1   g185(.A1(new_n371), .A2(G131), .ZN(new_n372));
  AOI21_X1  g186(.A(new_n294), .B1(new_n369), .B2(new_n370), .ZN(new_n373));
  OR3_X1    g187(.A1(new_n372), .A2(KEYINPUT17), .A3(new_n373), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n373), .A2(KEYINPUT17), .ZN(new_n375));
  OAI21_X1  g189(.A(KEYINPUT85), .B1(new_n364), .B2(new_n365), .ZN(new_n376));
  NAND4_X1  g190(.A1(new_n366), .A2(new_n374), .A3(new_n375), .A4(new_n376), .ZN(new_n377));
  NAND2_X1  g191(.A1(KEYINPUT18), .A2(G131), .ZN(new_n378));
  INV_X1    g192(.A(new_n378), .ZN(new_n379));
  AND3_X1   g193(.A1(new_n369), .A2(new_n370), .A3(new_n379), .ZN(new_n380));
  AOI22_X1  g194(.A1(new_n369), .A2(new_n370), .B1(KEYINPUT18), .B2(G131), .ZN(new_n381));
  NOR2_X1   g195(.A1(new_n380), .A2(new_n381), .ZN(new_n382));
  INV_X1    g196(.A(G125), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n383), .A2(G140), .ZN(new_n384));
  AND3_X1   g198(.A1(new_n361), .A2(new_n384), .A3(KEYINPUT72), .ZN(new_n385));
  AOI21_X1  g199(.A(KEYINPUT72), .B1(new_n361), .B2(new_n384), .ZN(new_n386));
  NOR3_X1   g200(.A1(new_n385), .A2(new_n386), .A3(G146), .ZN(new_n387));
  NOR2_X1   g201(.A1(new_n358), .A2(new_n226), .ZN(new_n388));
  OAI21_X1  g202(.A(KEYINPUT82), .B1(new_n387), .B2(new_n388), .ZN(new_n389));
  INV_X1    g203(.A(KEYINPUT72), .ZN(new_n390));
  NOR2_X1   g204(.A1(new_n383), .A2(G140), .ZN(new_n391));
  NOR2_X1   g205(.A1(new_n360), .A2(G125), .ZN(new_n392));
  OAI21_X1  g206(.A(new_n390), .B1(new_n391), .B2(new_n392), .ZN(new_n393));
  NAND3_X1  g207(.A1(new_n361), .A2(new_n384), .A3(KEYINPUT72), .ZN(new_n394));
  NAND3_X1  g208(.A1(new_n393), .A2(new_n226), .A3(new_n394), .ZN(new_n395));
  INV_X1    g209(.A(KEYINPUT82), .ZN(new_n396));
  OAI211_X1 g210(.A(new_n395), .B(new_n396), .C1(new_n226), .C2(new_n358), .ZN(new_n397));
  AOI21_X1  g211(.A(new_n382), .B1(new_n389), .B2(new_n397), .ZN(new_n398));
  INV_X1    g212(.A(new_n398), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n377), .A2(new_n399), .ZN(new_n400));
  XNOR2_X1  g214(.A(G113), .B(G122), .ZN(new_n401));
  XNOR2_X1  g215(.A(new_n401), .B(new_n207), .ZN(new_n402));
  INV_X1    g216(.A(new_n402), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n400), .A2(new_n403), .ZN(new_n404));
  NAND3_X1  g218(.A1(new_n377), .A2(new_n399), .A3(new_n402), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n404), .A2(new_n405), .ZN(new_n406));
  AOI21_X1  g220(.A(new_n357), .B1(new_n406), .B2(new_n189), .ZN(new_n407));
  INV_X1    g221(.A(new_n407), .ZN(new_n408));
  NOR2_X1   g222(.A1(new_n372), .A2(new_n373), .ZN(new_n409));
  INV_X1    g223(.A(KEYINPUT19), .ZN(new_n410));
  NAND3_X1  g224(.A1(new_n393), .A2(new_n410), .A3(new_n394), .ZN(new_n411));
  OAI21_X1  g225(.A(KEYINPUT19), .B1(new_n391), .B2(new_n392), .ZN(new_n412));
  NAND3_X1  g226(.A1(new_n411), .A2(new_n226), .A3(new_n412), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n413), .A2(new_n363), .ZN(new_n414));
  AOI21_X1  g228(.A(new_n409), .B1(new_n414), .B2(KEYINPUT83), .ZN(new_n415));
  INV_X1    g229(.A(KEYINPUT83), .ZN(new_n416));
  NAND3_X1  g230(.A1(new_n413), .A2(new_n416), .A3(new_n363), .ZN(new_n417));
  AOI21_X1  g231(.A(new_n398), .B1(new_n415), .B2(new_n417), .ZN(new_n418));
  OAI21_X1  g232(.A(KEYINPUT84), .B1(new_n418), .B2(new_n402), .ZN(new_n419));
  INV_X1    g233(.A(KEYINPUT84), .ZN(new_n420));
  AND3_X1   g234(.A1(new_n413), .A2(new_n416), .A3(new_n363), .ZN(new_n421));
  AOI21_X1  g235(.A(new_n416), .B1(new_n413), .B2(new_n363), .ZN(new_n422));
  NOR3_X1   g236(.A1(new_n421), .A2(new_n422), .A3(new_n409), .ZN(new_n423));
  OAI211_X1 g237(.A(new_n420), .B(new_n403), .C1(new_n423), .C2(new_n398), .ZN(new_n424));
  NAND3_X1  g238(.A1(new_n419), .A2(new_n424), .A3(new_n405), .ZN(new_n425));
  INV_X1    g239(.A(KEYINPUT20), .ZN(new_n426));
  NOR2_X1   g240(.A1(G475), .A2(G902), .ZN(new_n427));
  AND3_X1   g241(.A1(new_n425), .A2(new_n426), .A3(new_n427), .ZN(new_n428));
  AOI21_X1  g242(.A(new_n426), .B1(new_n425), .B2(new_n427), .ZN(new_n429));
  OAI21_X1  g243(.A(new_n408), .B1(new_n428), .B2(new_n429), .ZN(new_n430));
  INV_X1    g244(.A(KEYINPUT87), .ZN(new_n431));
  XNOR2_X1  g245(.A(G128), .B(G143), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n432), .A2(KEYINPUT13), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n228), .A2(G128), .ZN(new_n434));
  OAI211_X1 g248(.A(new_n433), .B(G134), .C1(KEYINPUT13), .C2(new_n434), .ZN(new_n435));
  XOR2_X1   g249(.A(G116), .B(G122), .Z(new_n436));
  NAND2_X1  g250(.A1(new_n436), .A2(G107), .ZN(new_n437));
  XNOR2_X1  g251(.A(G116), .B(G122), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n438), .A2(new_n210), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n437), .A2(new_n439), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n432), .A2(new_n302), .ZN(new_n441));
  NAND3_X1  g255(.A1(new_n435), .A2(new_n440), .A3(new_n441), .ZN(new_n442));
  XNOR2_X1  g256(.A(new_n432), .B(new_n302), .ZN(new_n443));
  NAND3_X1  g257(.A1(new_n195), .A2(KEYINPUT14), .A3(G122), .ZN(new_n444));
  OAI211_X1 g258(.A(G107), .B(new_n444), .C1(new_n436), .C2(KEYINPUT14), .ZN(new_n445));
  NAND3_X1  g259(.A1(new_n443), .A2(new_n439), .A3(new_n445), .ZN(new_n446));
  XOR2_X1   g260(.A(KEYINPUT70), .B(G217), .Z(new_n447));
  NAND3_X1  g261(.A1(new_n447), .A2(new_n188), .A3(new_n320), .ZN(new_n448));
  INV_X1    g262(.A(new_n448), .ZN(new_n449));
  NAND3_X1  g263(.A1(new_n442), .A2(new_n446), .A3(new_n449), .ZN(new_n450));
  AOI21_X1  g264(.A(new_n449), .B1(new_n442), .B2(new_n446), .ZN(new_n451));
  OAI21_X1  g265(.A(new_n450), .B1(new_n451), .B2(KEYINPUT86), .ZN(new_n452));
  INV_X1    g266(.A(KEYINPUT86), .ZN(new_n453));
  AOI211_X1 g267(.A(new_n453), .B(new_n449), .C1(new_n442), .C2(new_n446), .ZN(new_n454));
  OAI211_X1 g268(.A(new_n431), .B(new_n189), .C1(new_n452), .C2(new_n454), .ZN(new_n455));
  INV_X1    g269(.A(G478), .ZN(new_n456));
  NOR2_X1   g270(.A1(new_n456), .A2(KEYINPUT15), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n455), .A2(new_n457), .ZN(new_n458));
  AND2_X1   g272(.A1(new_n442), .A2(new_n446), .ZN(new_n459));
  OAI21_X1  g273(.A(new_n453), .B1(new_n459), .B2(new_n449), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n451), .A2(KEYINPUT86), .ZN(new_n461));
  NAND3_X1  g275(.A1(new_n460), .A2(new_n461), .A3(new_n450), .ZN(new_n462));
  INV_X1    g276(.A(new_n457), .ZN(new_n463));
  NAND4_X1  g277(.A1(new_n462), .A2(new_n431), .A3(new_n189), .A4(new_n463), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n458), .A2(new_n464), .ZN(new_n465));
  INV_X1    g279(.A(KEYINPUT88), .ZN(new_n466));
  XNOR2_X1  g280(.A(new_n465), .B(new_n466), .ZN(new_n467));
  AOI211_X1 g281(.A(new_n189), .B(new_n320), .C1(G234), .C2(G237), .ZN(new_n468));
  XNOR2_X1  g282(.A(KEYINPUT21), .B(G898), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  INV_X1    g284(.A(G952), .ZN(new_n471));
  AOI211_X1 g285(.A(G953), .B(new_n471), .C1(G234), .C2(G237), .ZN(new_n472));
  INV_X1    g286(.A(new_n472), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n470), .A2(new_n473), .ZN(new_n474));
  XOR2_X1   g288(.A(new_n474), .B(KEYINPUT89), .Z(new_n475));
  INV_X1    g289(.A(new_n475), .ZN(new_n476));
  NOR3_X1   g290(.A1(new_n430), .A2(new_n467), .A3(new_n476), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n356), .A2(new_n477), .ZN(new_n478));
  INV_X1    g292(.A(KEYINPUT68), .ZN(new_n479));
  NAND3_X1  g293(.A1(new_n307), .A2(new_n313), .A3(new_n310), .ZN(new_n480));
  OAI21_X1  g294(.A(KEYINPUT64), .B1(new_n302), .B2(G137), .ZN(new_n481));
  INV_X1    g295(.A(KEYINPUT64), .ZN(new_n482));
  NAND3_X1  g296(.A1(new_n482), .A2(new_n295), .A3(G134), .ZN(new_n483));
  NAND3_X1  g297(.A1(new_n481), .A2(new_n483), .A3(new_n304), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n484), .A2(G131), .ZN(new_n485));
  AND2_X1   g299(.A1(new_n485), .A2(new_n305), .ZN(new_n486));
  OAI21_X1  g300(.A(new_n486), .B1(new_n290), .B2(new_n291), .ZN(new_n487));
  NOR2_X1   g301(.A1(new_n222), .A2(new_n262), .ZN(new_n488));
  AND3_X1   g302(.A1(new_n480), .A2(new_n487), .A3(new_n488), .ZN(new_n489));
  AOI21_X1  g303(.A(new_n488), .B1(new_n480), .B2(new_n487), .ZN(new_n490));
  OAI211_X1 g304(.A(new_n479), .B(KEYINPUT28), .C1(new_n489), .C2(new_n490), .ZN(new_n491));
  INV_X1    g305(.A(KEYINPUT28), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n480), .A2(new_n487), .ZN(new_n493));
  INV_X1    g307(.A(new_n488), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  NAND3_X1  g309(.A1(new_n480), .A2(new_n487), .A3(new_n488), .ZN(new_n496));
  AOI21_X1  g310(.A(new_n492), .B1(new_n495), .B2(new_n496), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n496), .A2(new_n492), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n498), .A2(KEYINPUT68), .ZN(new_n499));
  OAI21_X1  g313(.A(new_n491), .B1(new_n497), .B2(new_n499), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n367), .A2(G210), .ZN(new_n501));
  XNOR2_X1  g315(.A(new_n501), .B(KEYINPUT27), .ZN(new_n502));
  XNOR2_X1  g316(.A(KEYINPUT26), .B(G101), .ZN(new_n503));
  XNOR2_X1  g317(.A(new_n502), .B(new_n503), .ZN(new_n504));
  INV_X1    g318(.A(new_n504), .ZN(new_n505));
  INV_X1    g319(.A(KEYINPUT29), .ZN(new_n506));
  NOR2_X1   g320(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n500), .A2(new_n507), .ZN(new_n508));
  NAND3_X1  g322(.A1(new_n480), .A2(new_n487), .A3(KEYINPUT30), .ZN(new_n509));
  INV_X1    g323(.A(KEYINPUT30), .ZN(new_n510));
  AOI21_X1  g324(.A(new_n312), .B1(new_n309), .B2(new_n305), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n485), .A2(new_n305), .ZN(new_n512));
  NOR2_X1   g326(.A1(new_n512), .A2(new_n240), .ZN(new_n513));
  OAI21_X1  g327(.A(new_n510), .B1(new_n511), .B2(new_n513), .ZN(new_n514));
  NAND3_X1  g328(.A1(new_n509), .A2(new_n494), .A3(new_n514), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n515), .A2(new_n496), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n516), .A2(new_n505), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n489), .A2(KEYINPUT28), .ZN(new_n518));
  OAI21_X1  g332(.A(new_n494), .B1(new_n513), .B2(new_n511), .ZN(new_n519));
  NAND4_X1  g333(.A1(new_n518), .A2(new_n504), .A3(new_n498), .A4(new_n519), .ZN(new_n520));
  NAND3_X1  g334(.A1(new_n517), .A2(new_n520), .A3(new_n506), .ZN(new_n521));
  NAND3_X1  g335(.A1(new_n508), .A2(new_n521), .A3(new_n189), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n522), .A2(G472), .ZN(new_n523));
  INV_X1    g337(.A(KEYINPUT32), .ZN(new_n524));
  NAND3_X1  g338(.A1(new_n515), .A2(new_n504), .A3(new_n496), .ZN(new_n525));
  INV_X1    g339(.A(KEYINPUT31), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  NAND4_X1  g341(.A1(new_n515), .A2(KEYINPUT31), .A3(new_n504), .A4(new_n496), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  NAND3_X1  g343(.A1(new_n518), .A2(new_n498), .A3(new_n519), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n530), .A2(new_n505), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n529), .A2(new_n531), .ZN(new_n532));
  NOR2_X1   g346(.A1(G472), .A2(G902), .ZN(new_n533));
  AOI21_X1  g347(.A(new_n524), .B1(new_n532), .B2(new_n533), .ZN(new_n534));
  AOI22_X1  g348(.A1(new_n527), .A2(new_n528), .B1(new_n505), .B2(new_n530), .ZN(new_n535));
  INV_X1    g349(.A(new_n533), .ZN(new_n536));
  NOR3_X1   g350(.A1(new_n535), .A2(KEYINPUT32), .A3(new_n536), .ZN(new_n537));
  OAI21_X1  g351(.A(new_n523), .B1(new_n534), .B2(new_n537), .ZN(new_n538));
  INV_X1    g352(.A(KEYINPUT69), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  NAND3_X1  g354(.A1(new_n532), .A2(new_n524), .A3(new_n533), .ZN(new_n541));
  OAI21_X1  g355(.A(KEYINPUT32), .B1(new_n535), .B2(new_n536), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  NAND3_X1  g357(.A1(new_n543), .A2(KEYINPUT69), .A3(new_n523), .ZN(new_n544));
  INV_X1    g358(.A(KEYINPUT25), .ZN(new_n545));
  XNOR2_X1  g359(.A(KEYINPUT22), .B(G137), .ZN(new_n546));
  INV_X1    g360(.A(G234), .ZN(new_n547));
  NOR3_X1   g361(.A1(new_n187), .A2(new_n547), .A3(G953), .ZN(new_n548));
  XOR2_X1   g362(.A(new_n546), .B(new_n548), .Z(new_n549));
  INV_X1    g363(.A(new_n549), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n199), .A2(G128), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n551), .A2(KEYINPUT23), .ZN(new_n552));
  INV_X1    g366(.A(G128), .ZN(new_n553));
  AOI21_X1  g367(.A(KEYINPUT71), .B1(new_n553), .B2(G119), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n552), .A2(new_n554), .ZN(new_n555));
  NOR2_X1   g369(.A1(new_n199), .A2(G128), .ZN(new_n556));
  OAI211_X1 g370(.A(KEYINPUT23), .B(new_n551), .C1(new_n556), .C2(KEYINPUT71), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n555), .A2(new_n557), .ZN(new_n558));
  XNOR2_X1  g372(.A(G119), .B(G128), .ZN(new_n559));
  XOR2_X1   g373(.A(KEYINPUT24), .B(G110), .Z(new_n560));
  OAI22_X1  g374(.A1(new_n558), .A2(G110), .B1(new_n559), .B2(new_n560), .ZN(new_n561));
  NAND3_X1  g375(.A1(new_n561), .A2(new_n363), .A3(new_n395), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n558), .A2(G110), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n560), .A2(new_n559), .ZN(new_n564));
  OAI211_X1 g378(.A(new_n563), .B(new_n564), .C1(new_n364), .C2(new_n365), .ZN(new_n565));
  AND3_X1   g379(.A1(new_n562), .A2(KEYINPUT73), .A3(new_n565), .ZN(new_n566));
  AOI21_X1  g380(.A(KEYINPUT73), .B1(new_n562), .B2(new_n565), .ZN(new_n567));
  OAI21_X1  g381(.A(new_n550), .B1(new_n566), .B2(new_n567), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n562), .A2(new_n565), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n569), .A2(new_n549), .ZN(new_n570));
  AOI21_X1  g384(.A(G902), .B1(new_n568), .B2(new_n570), .ZN(new_n571));
  INV_X1    g385(.A(KEYINPUT74), .ZN(new_n572));
  OAI21_X1  g386(.A(new_n545), .B1(new_n571), .B2(new_n572), .ZN(new_n573));
  INV_X1    g387(.A(new_n570), .ZN(new_n574));
  INV_X1    g388(.A(KEYINPUT73), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n569), .A2(new_n575), .ZN(new_n576));
  NAND3_X1  g390(.A1(new_n562), .A2(new_n565), .A3(KEYINPUT73), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  AOI21_X1  g392(.A(new_n574), .B1(new_n578), .B2(new_n550), .ZN(new_n579));
  OAI211_X1 g393(.A(KEYINPUT74), .B(KEYINPUT25), .C1(new_n579), .C2(G902), .ZN(new_n580));
  OAI21_X1  g394(.A(new_n447), .B1(new_n547), .B2(G902), .ZN(new_n581));
  INV_X1    g395(.A(new_n581), .ZN(new_n582));
  NAND3_X1  g396(.A1(new_n573), .A2(new_n580), .A3(new_n582), .ZN(new_n583));
  INV_X1    g397(.A(new_n579), .ZN(new_n584));
  NOR2_X1   g398(.A1(new_n582), .A2(G902), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n583), .A2(new_n586), .ZN(new_n587));
  INV_X1    g401(.A(new_n587), .ZN(new_n588));
  NAND3_X1  g402(.A1(new_n540), .A2(new_n544), .A3(new_n588), .ZN(new_n589));
  NOR2_X1   g403(.A1(new_n478), .A2(new_n589), .ZN(new_n590));
  XNOR2_X1  g404(.A(new_n590), .B(new_n212), .ZN(G3));
  INV_X1    g405(.A(KEYINPUT90), .ZN(new_n592));
  OAI211_X1 g406(.A(new_n592), .B(G472), .C1(new_n535), .C2(G902), .ZN(new_n593));
  INV_X1    g407(.A(new_n593), .ZN(new_n594));
  OAI21_X1  g408(.A(G472), .B1(new_n535), .B2(G902), .ZN(new_n595));
  OAI21_X1  g409(.A(new_n592), .B1(new_n535), .B2(new_n536), .ZN(new_n596));
  AOI21_X1  g410(.A(new_n594), .B1(new_n595), .B2(new_n596), .ZN(new_n597));
  INV_X1    g411(.A(new_n282), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n355), .A2(new_n191), .ZN(new_n599));
  NOR2_X1   g413(.A1(new_n599), .A2(new_n587), .ZN(new_n600));
  AND3_X1   g414(.A1(new_n597), .A2(new_n598), .A3(new_n600), .ZN(new_n601));
  INV_X1    g415(.A(KEYINPUT33), .ZN(new_n602));
  NOR2_X1   g416(.A1(new_n451), .A2(new_n602), .ZN(new_n603));
  AOI22_X1  g417(.A1(new_n462), .A2(new_n602), .B1(new_n450), .B2(new_n603), .ZN(new_n604));
  NAND3_X1  g418(.A1(new_n604), .A2(G478), .A3(new_n189), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n462), .A2(new_n189), .ZN(new_n606));
  XNOR2_X1  g420(.A(KEYINPUT91), .B(G478), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n605), .A2(new_n608), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n430), .A2(new_n609), .ZN(new_n610));
  NOR2_X1   g424(.A1(new_n610), .A2(new_n476), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n601), .A2(new_n611), .ZN(new_n612));
  XNOR2_X1  g426(.A(new_n612), .B(new_n207), .ZN(new_n613));
  XNOR2_X1  g427(.A(KEYINPUT92), .B(KEYINPUT34), .ZN(new_n614));
  XNOR2_X1  g428(.A(new_n613), .B(new_n614), .ZN(G6));
  NAND2_X1  g429(.A1(new_n425), .A2(new_n427), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n616), .A2(KEYINPUT20), .ZN(new_n617));
  INV_X1    g431(.A(KEYINPUT93), .ZN(new_n618));
  NAND3_X1  g432(.A1(new_n425), .A2(new_n426), .A3(new_n427), .ZN(new_n619));
  NAND3_X1  g433(.A1(new_n617), .A2(new_n618), .A3(new_n619), .ZN(new_n620));
  AOI21_X1  g434(.A(new_n407), .B1(new_n429), .B2(KEYINPUT93), .ZN(new_n621));
  NAND4_X1  g435(.A1(new_n467), .A2(new_n620), .A3(new_n475), .A4(new_n621), .ZN(new_n622));
  XNOR2_X1  g436(.A(new_n622), .B(KEYINPUT94), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n623), .A2(new_n601), .ZN(new_n624));
  XOR2_X1   g438(.A(KEYINPUT35), .B(G107), .Z(new_n625));
  XNOR2_X1  g439(.A(new_n624), .B(new_n625), .ZN(G9));
  NOR2_X1   g440(.A1(new_n550), .A2(KEYINPUT36), .ZN(new_n627));
  XOR2_X1   g441(.A(new_n578), .B(new_n627), .Z(new_n628));
  NAND2_X1  g442(.A1(new_n628), .A2(new_n585), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n583), .A2(new_n629), .ZN(new_n630));
  NAND4_X1  g444(.A1(new_n356), .A2(new_n597), .A3(new_n477), .A4(new_n630), .ZN(new_n631));
  XOR2_X1   g445(.A(KEYINPUT37), .B(G110), .Z(new_n632));
  XNOR2_X1  g446(.A(new_n631), .B(new_n632), .ZN(G12));
  NAND2_X1  g447(.A1(new_n620), .A2(new_n621), .ZN(new_n634));
  XNOR2_X1  g448(.A(new_n465), .B(KEYINPUT88), .ZN(new_n635));
  INV_X1    g449(.A(G900), .ZN(new_n636));
  AOI21_X1  g450(.A(new_n472), .B1(new_n468), .B2(new_n636), .ZN(new_n637));
  NOR3_X1   g451(.A1(new_n634), .A2(new_n635), .A3(new_n637), .ZN(new_n638));
  AND2_X1   g452(.A1(new_n583), .A2(new_n629), .ZN(new_n639));
  NOR2_X1   g453(.A1(new_n639), .A2(new_n282), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n638), .A2(new_n640), .ZN(new_n641));
  INV_X1    g455(.A(new_n599), .ZN(new_n642));
  NAND3_X1  g456(.A1(new_n540), .A2(new_n544), .A3(new_n642), .ZN(new_n643));
  NOR2_X1   g457(.A1(new_n641), .A2(new_n643), .ZN(new_n644));
  XNOR2_X1  g458(.A(new_n644), .B(new_n553), .ZN(G30));
  XOR2_X1   g459(.A(new_n288), .B(KEYINPUT38), .Z(new_n646));
  INV_X1    g460(.A(new_n192), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n430), .A2(new_n467), .ZN(new_n648));
  NOR4_X1   g462(.A1(new_n646), .A2(new_n647), .A3(new_n648), .A4(new_n630), .ZN(new_n649));
  XOR2_X1   g463(.A(new_n637), .B(KEYINPUT39), .Z(new_n650));
  INV_X1    g464(.A(new_n650), .ZN(new_n651));
  NOR2_X1   g465(.A1(new_n599), .A2(new_n651), .ZN(new_n652));
  INV_X1    g466(.A(new_n652), .ZN(new_n653));
  XNOR2_X1  g467(.A(KEYINPUT97), .B(KEYINPUT40), .ZN(new_n654));
  OR2_X1    g468(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  AOI21_X1  g469(.A(new_n505), .B1(new_n515), .B2(new_n496), .ZN(new_n656));
  NOR3_X1   g470(.A1(new_n489), .A2(new_n490), .A3(new_n504), .ZN(new_n657));
  OAI21_X1  g471(.A(KEYINPUT95), .B1(new_n656), .B2(new_n657), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n658), .A2(new_n189), .ZN(new_n659));
  NOR3_X1   g473(.A1(new_n656), .A2(new_n657), .A3(KEYINPUT95), .ZN(new_n660));
  OAI21_X1  g474(.A(G472), .B1(new_n659), .B2(new_n660), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n543), .A2(new_n661), .ZN(new_n662));
  INV_X1    g476(.A(KEYINPUT96), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  NAND3_X1  g478(.A1(new_n543), .A2(KEYINPUT96), .A3(new_n661), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  NAND2_X1  g480(.A1(new_n653), .A2(new_n654), .ZN(new_n667));
  NAND4_X1  g481(.A1(new_n649), .A2(new_n655), .A3(new_n666), .A4(new_n667), .ZN(new_n668));
  XNOR2_X1  g482(.A(new_n668), .B(G143), .ZN(G45));
  INV_X1    g483(.A(new_n637), .ZN(new_n670));
  NAND3_X1  g484(.A1(new_n430), .A2(new_n609), .A3(new_n670), .ZN(new_n671));
  INV_X1    g485(.A(KEYINPUT98), .ZN(new_n672));
  NAND2_X1  g486(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  NAND4_X1  g487(.A1(new_n430), .A2(KEYINPUT98), .A3(new_n609), .A4(new_n670), .ZN(new_n674));
  AND3_X1   g488(.A1(new_n673), .A2(new_n640), .A3(new_n674), .ZN(new_n675));
  AND3_X1   g489(.A1(new_n540), .A2(new_n544), .A3(new_n642), .ZN(new_n676));
  NAND2_X1  g490(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  XNOR2_X1  g491(.A(new_n677), .B(G146), .ZN(G48));
  AOI211_X1 g492(.A(new_n339), .B(KEYINPUT12), .C1(new_n330), .C2(new_n341), .ZN(new_n679));
  AOI21_X1  g493(.A(KEYINPUT76), .B1(new_n342), .B2(new_n335), .ZN(new_n680));
  OAI21_X1  g494(.A(new_n345), .B1(new_n679), .B2(new_n680), .ZN(new_n681));
  INV_X1    g495(.A(new_n324), .ZN(new_n682));
  AOI21_X1  g496(.A(new_n352), .B1(new_n681), .B2(new_n682), .ZN(new_n683));
  OAI21_X1  g497(.A(G469), .B1(new_n683), .B2(G902), .ZN(new_n684));
  NAND3_X1  g498(.A1(new_n684), .A2(new_n191), .A3(new_n353), .ZN(new_n685));
  NAND2_X1  g499(.A1(new_n685), .A2(KEYINPUT99), .ZN(new_n686));
  INV_X1    g500(.A(KEYINPUT99), .ZN(new_n687));
  NAND4_X1  g501(.A1(new_n684), .A2(new_n353), .A3(new_n687), .A4(new_n191), .ZN(new_n688));
  NAND3_X1  g502(.A1(new_n686), .A2(new_n598), .A3(new_n688), .ZN(new_n689));
  NOR2_X1   g503(.A1(new_n589), .A2(new_n689), .ZN(new_n690));
  NAND2_X1  g504(.A1(new_n690), .A2(new_n611), .ZN(new_n691));
  XNOR2_X1  g505(.A(KEYINPUT41), .B(G113), .ZN(new_n692));
  XNOR2_X1  g506(.A(new_n691), .B(new_n692), .ZN(G15));
  NAND2_X1  g507(.A1(new_n690), .A2(new_n623), .ZN(new_n694));
  XNOR2_X1  g508(.A(new_n694), .B(G116), .ZN(G18));
  AND3_X1   g509(.A1(new_n686), .A2(new_n598), .A3(new_n688), .ZN(new_n696));
  AOI21_X1  g510(.A(new_n407), .B1(new_n617), .B2(new_n619), .ZN(new_n697));
  AND4_X1   g511(.A1(new_n697), .A2(new_n630), .A3(new_n635), .A4(new_n475), .ZN(new_n698));
  NAND4_X1  g512(.A1(new_n696), .A2(new_n698), .A3(new_n540), .A4(new_n544), .ZN(new_n699));
  INV_X1    g513(.A(KEYINPUT100), .ZN(new_n700));
  NAND2_X1  g514(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  NAND4_X1  g515(.A1(new_n697), .A2(new_n630), .A3(new_n635), .A4(new_n475), .ZN(new_n702));
  NOR2_X1   g516(.A1(new_n689), .A2(new_n702), .ZN(new_n703));
  NAND4_X1  g517(.A1(new_n703), .A2(KEYINPUT100), .A3(new_n540), .A4(new_n544), .ZN(new_n704));
  NAND2_X1  g518(.A1(new_n701), .A2(new_n704), .ZN(new_n705));
  XNOR2_X1  g519(.A(new_n705), .B(G119), .ZN(G21));
  INV_X1    g520(.A(KEYINPUT102), .ZN(new_n707));
  OAI21_X1  g521(.A(new_n707), .B1(new_n697), .B2(new_n635), .ZN(new_n708));
  NAND3_X1  g522(.A1(new_n430), .A2(new_n467), .A3(KEYINPUT102), .ZN(new_n709));
  NAND2_X1  g523(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  NAND4_X1  g524(.A1(new_n686), .A2(new_n475), .A3(new_n598), .A4(new_n688), .ZN(new_n711));
  OAI21_X1  g525(.A(new_n529), .B1(new_n504), .B2(new_n500), .ZN(new_n712));
  NAND2_X1  g526(.A1(new_n712), .A2(new_n533), .ZN(new_n713));
  XOR2_X1   g527(.A(KEYINPUT101), .B(G472), .Z(new_n714));
  OAI21_X1  g528(.A(new_n714), .B1(new_n535), .B2(G902), .ZN(new_n715));
  NAND3_X1  g529(.A1(new_n588), .A2(new_n713), .A3(new_n715), .ZN(new_n716));
  NOR3_X1   g530(.A1(new_n710), .A2(new_n711), .A3(new_n716), .ZN(new_n717));
  XOR2_X1   g531(.A(new_n717), .B(G122), .Z(G24));
  NAND2_X1  g532(.A1(new_n673), .A2(new_n674), .ZN(new_n719));
  NAND2_X1  g533(.A1(new_n719), .A2(KEYINPUT103), .ZN(new_n720));
  NAND2_X1  g534(.A1(new_n713), .A2(new_n715), .ZN(new_n721));
  NOR2_X1   g535(.A1(new_n639), .A2(new_n721), .ZN(new_n722));
  INV_X1    g536(.A(new_n722), .ZN(new_n723));
  NOR2_X1   g537(.A1(new_n723), .A2(new_n689), .ZN(new_n724));
  INV_X1    g538(.A(KEYINPUT103), .ZN(new_n725));
  NAND3_X1  g539(.A1(new_n673), .A2(new_n725), .A3(new_n674), .ZN(new_n726));
  NAND3_X1  g540(.A1(new_n720), .A2(new_n724), .A3(new_n726), .ZN(new_n727));
  XNOR2_X1  g541(.A(new_n727), .B(G125), .ZN(G27));
  AND3_X1   g542(.A1(new_n540), .A2(new_n544), .A3(new_n588), .ZN(new_n729));
  INV_X1    g543(.A(KEYINPUT104), .ZN(new_n730));
  NAND2_X1  g544(.A1(new_n599), .A2(new_n730), .ZN(new_n731));
  NAND3_X1  g545(.A1(new_n355), .A2(KEYINPUT104), .A3(new_n191), .ZN(new_n732));
  NOR2_X1   g546(.A1(new_n288), .A2(new_n647), .ZN(new_n733));
  AND3_X1   g547(.A1(new_n731), .A2(new_n732), .A3(new_n733), .ZN(new_n734));
  NAND4_X1  g548(.A1(new_n720), .A2(new_n729), .A3(new_n726), .A4(new_n734), .ZN(new_n735));
  INV_X1    g549(.A(KEYINPUT42), .ZN(new_n736));
  AND3_X1   g550(.A1(new_n673), .A2(new_n725), .A3(new_n674), .ZN(new_n737));
  AOI21_X1  g551(.A(new_n725), .B1(new_n673), .B2(new_n674), .ZN(new_n738));
  NOR2_X1   g552(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  NAND4_X1  g553(.A1(new_n731), .A2(KEYINPUT42), .A3(new_n732), .A4(new_n733), .ZN(new_n740));
  NAND2_X1  g554(.A1(new_n538), .A2(new_n588), .ZN(new_n741));
  NAND2_X1  g555(.A1(new_n741), .A2(KEYINPUT105), .ZN(new_n742));
  INV_X1    g556(.A(KEYINPUT105), .ZN(new_n743));
  NAND3_X1  g557(.A1(new_n538), .A2(new_n743), .A3(new_n588), .ZN(new_n744));
  AOI21_X1  g558(.A(new_n740), .B1(new_n742), .B2(new_n744), .ZN(new_n745));
  AOI22_X1  g559(.A1(new_n735), .A2(new_n736), .B1(new_n739), .B2(new_n745), .ZN(new_n746));
  XNOR2_X1  g560(.A(new_n746), .B(new_n294), .ZN(G33));
  NAND3_X1  g561(.A1(new_n729), .A2(new_n638), .A3(new_n734), .ZN(new_n748));
  XNOR2_X1  g562(.A(new_n748), .B(G134), .ZN(G36));
  NOR2_X1   g563(.A1(new_n597), .A2(new_n639), .ZN(new_n750));
  NAND2_X1  g564(.A1(new_n697), .A2(new_n609), .ZN(new_n751));
  NAND2_X1  g565(.A1(new_n751), .A2(KEYINPUT107), .ZN(new_n752));
  INV_X1    g566(.A(KEYINPUT43), .ZN(new_n753));
  NAND2_X1  g567(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  NAND3_X1  g568(.A1(new_n751), .A2(KEYINPUT107), .A3(KEYINPUT43), .ZN(new_n755));
  NAND4_X1  g569(.A1(new_n750), .A2(new_n754), .A3(KEYINPUT44), .A4(new_n755), .ZN(new_n756));
  XOR2_X1   g570(.A(new_n756), .B(KEYINPUT108), .Z(new_n757));
  INV_X1    g571(.A(new_n681), .ZN(new_n758));
  OAI21_X1  g572(.A(new_n347), .B1(new_n758), .B2(new_n334), .ZN(new_n759));
  NAND2_X1  g573(.A1(new_n759), .A2(new_n333), .ZN(new_n760));
  INV_X1    g574(.A(KEYINPUT45), .ZN(new_n761));
  NAND2_X1  g575(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  NAND3_X1  g576(.A1(new_n759), .A2(KEYINPUT45), .A3(new_n333), .ZN(new_n763));
  NAND3_X1  g577(.A1(new_n762), .A2(G469), .A3(new_n763), .ZN(new_n764));
  NAND2_X1  g578(.A1(new_n764), .A2(new_n354), .ZN(new_n765));
  INV_X1    g579(.A(KEYINPUT46), .ZN(new_n766));
  NAND3_X1  g580(.A1(new_n765), .A2(KEYINPUT106), .A3(new_n766), .ZN(new_n767));
  NAND3_X1  g581(.A1(new_n764), .A2(KEYINPUT46), .A3(new_n354), .ZN(new_n768));
  NAND3_X1  g582(.A1(new_n767), .A2(new_n353), .A3(new_n768), .ZN(new_n769));
  INV_X1    g583(.A(new_n769), .ZN(new_n770));
  NAND2_X1  g584(.A1(new_n765), .A2(new_n766), .ZN(new_n771));
  INV_X1    g585(.A(KEYINPUT106), .ZN(new_n772));
  NAND2_X1  g586(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  AOI21_X1  g587(.A(new_n190), .B1(new_n770), .B2(new_n773), .ZN(new_n774));
  INV_X1    g588(.A(new_n733), .ZN(new_n775));
  NAND3_X1  g589(.A1(new_n750), .A2(new_n754), .A3(new_n755), .ZN(new_n776));
  INV_X1    g590(.A(KEYINPUT44), .ZN(new_n777));
  AOI21_X1  g591(.A(new_n775), .B1(new_n776), .B2(new_n777), .ZN(new_n778));
  NAND3_X1  g592(.A1(new_n774), .A2(new_n650), .A3(new_n778), .ZN(new_n779));
  OR2_X1    g593(.A1(new_n757), .A2(new_n779), .ZN(new_n780));
  XNOR2_X1  g594(.A(new_n780), .B(G137), .ZN(G39));
  INV_X1    g595(.A(KEYINPUT47), .ZN(new_n782));
  INV_X1    g596(.A(new_n773), .ZN(new_n783));
  OAI221_X1 g597(.A(new_n191), .B1(KEYINPUT109), .B2(new_n782), .C1(new_n783), .C2(new_n769), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n733), .A2(new_n587), .ZN(new_n785));
  AOI211_X1 g599(.A(new_n785), .B(new_n719), .C1(new_n540), .C2(new_n544), .ZN(new_n786));
  XNOR2_X1  g600(.A(KEYINPUT109), .B(KEYINPUT47), .ZN(new_n787));
  OAI211_X1 g601(.A(new_n784), .B(new_n786), .C1(new_n774), .C2(new_n787), .ZN(new_n788));
  XNOR2_X1  g602(.A(new_n788), .B(G140), .ZN(G42));
  NAND2_X1  g603(.A1(new_n696), .A2(new_n722), .ZN(new_n790));
  NOR3_X1   g604(.A1(new_n737), .A2(new_n738), .A3(new_n790), .ZN(new_n791));
  OAI21_X1  g605(.A(KEYINPUT110), .B1(new_n791), .B2(new_n644), .ZN(new_n792));
  NAND3_X1  g606(.A1(new_n642), .A2(new_n639), .A3(new_n670), .ZN(new_n793));
  AOI21_X1  g607(.A(new_n793), .B1(new_n664), .B2(new_n665), .ZN(new_n794));
  NOR2_X1   g608(.A1(new_n710), .A2(new_n282), .ZN(new_n795));
  NAND2_X1  g609(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  NAND3_X1  g610(.A1(new_n676), .A2(new_n640), .A3(new_n638), .ZN(new_n797));
  INV_X1    g611(.A(KEYINPUT110), .ZN(new_n798));
  NAND3_X1  g612(.A1(new_n727), .A2(new_n797), .A3(new_n798), .ZN(new_n799));
  NAND4_X1  g613(.A1(new_n792), .A2(new_n677), .A3(new_n796), .A4(new_n799), .ZN(new_n800));
  NAND2_X1  g614(.A1(new_n800), .A2(KEYINPUT52), .ZN(new_n801));
  AOI22_X1  g615(.A1(new_n795), .A2(new_n794), .B1(new_n675), .B2(new_n676), .ZN(new_n802));
  INV_X1    g616(.A(KEYINPUT52), .ZN(new_n803));
  NAND4_X1  g617(.A1(new_n802), .A2(new_n803), .A3(new_n797), .A4(new_n727), .ZN(new_n804));
  NAND2_X1  g618(.A1(new_n801), .A2(new_n804), .ZN(new_n805));
  NAND2_X1  g619(.A1(new_n735), .A2(new_n736), .ZN(new_n806));
  NAND2_X1  g620(.A1(new_n739), .A2(new_n745), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n806), .A2(new_n807), .ZN(new_n808));
  INV_X1    g622(.A(KEYINPUT111), .ZN(new_n809));
  AOI21_X1  g623(.A(new_n717), .B1(new_n690), .B2(new_n611), .ZN(new_n810));
  AOI22_X1  g624(.A1(new_n701), .A2(new_n704), .B1(new_n690), .B2(new_n623), .ZN(new_n811));
  NAND4_X1  g625(.A1(new_n808), .A2(new_n809), .A3(new_n810), .A4(new_n811), .ZN(new_n812));
  NAND3_X1  g626(.A1(new_n810), .A2(new_n705), .A3(new_n694), .ZN(new_n813));
  OAI21_X1  g627(.A(KEYINPUT111), .B1(new_n813), .B2(new_n746), .ZN(new_n814));
  INV_X1    g628(.A(new_n465), .ZN(new_n815));
  NAND3_X1  g629(.A1(new_n630), .A2(new_n815), .A3(new_n670), .ZN(new_n816));
  NOR3_X1   g630(.A1(new_n816), .A2(new_n775), .A3(new_n634), .ZN(new_n817));
  NAND2_X1  g631(.A1(new_n676), .A2(new_n817), .ZN(new_n818));
  NAND2_X1  g632(.A1(new_n748), .A2(new_n818), .ZN(new_n819));
  OAI21_X1  g633(.A(new_n610), .B1(new_n430), .B2(new_n815), .ZN(new_n820));
  AND3_X1   g634(.A1(new_n284), .A2(new_n289), .A3(new_n475), .ZN(new_n821));
  NAND4_X1  g635(.A1(new_n820), .A2(new_n821), .A3(new_n597), .A4(new_n600), .ZN(new_n822));
  OAI211_X1 g636(.A(new_n631), .B(new_n822), .C1(new_n589), .C2(new_n478), .ZN(new_n823));
  NAND4_X1  g637(.A1(new_n722), .A2(new_n731), .A3(new_n732), .A4(new_n733), .ZN(new_n824));
  NOR3_X1   g638(.A1(new_n737), .A2(new_n738), .A3(new_n824), .ZN(new_n825));
  INV_X1    g639(.A(KEYINPUT53), .ZN(new_n826));
  NOR4_X1   g640(.A1(new_n819), .A2(new_n823), .A3(new_n825), .A4(new_n826), .ZN(new_n827));
  NAND3_X1  g641(.A1(new_n812), .A2(new_n814), .A3(new_n827), .ZN(new_n828));
  OR2_X1    g642(.A1(new_n805), .A2(new_n828), .ZN(new_n829));
  INV_X1    g643(.A(KEYINPUT54), .ZN(new_n830));
  AND3_X1   g644(.A1(new_n810), .A2(new_n705), .A3(new_n694), .ZN(new_n831));
  NOR3_X1   g645(.A1(new_n819), .A2(new_n823), .A3(new_n825), .ZN(new_n832));
  NAND3_X1  g646(.A1(new_n831), .A2(new_n832), .A3(new_n808), .ZN(new_n833));
  NAND4_X1  g647(.A1(new_n727), .A2(new_n796), .A3(new_n797), .A4(new_n677), .ZN(new_n834));
  NAND2_X1  g648(.A1(new_n834), .A2(KEYINPUT52), .ZN(new_n835));
  NAND2_X1  g649(.A1(new_n835), .A2(new_n804), .ZN(new_n836));
  OAI21_X1  g650(.A(new_n826), .B1(new_n833), .B2(new_n836), .ZN(new_n837));
  NAND3_X1  g651(.A1(new_n829), .A2(new_n830), .A3(new_n837), .ZN(new_n838));
  INV_X1    g652(.A(KEYINPUT112), .ZN(new_n839));
  NAND2_X1  g653(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  NAND4_X1  g654(.A1(new_n829), .A2(KEYINPUT112), .A3(new_n830), .A4(new_n837), .ZN(new_n841));
  OR3_X1    g655(.A1(new_n805), .A2(KEYINPUT53), .A3(new_n833), .ZN(new_n842));
  OAI21_X1  g656(.A(KEYINPUT53), .B1(new_n833), .B2(new_n836), .ZN(new_n843));
  NAND3_X1  g657(.A1(new_n842), .A2(KEYINPUT54), .A3(new_n843), .ZN(new_n844));
  NAND3_X1  g658(.A1(new_n840), .A2(new_n841), .A3(new_n844), .ZN(new_n845));
  AND3_X1   g659(.A1(new_n754), .A2(new_n472), .A3(new_n755), .ZN(new_n846));
  AND3_X1   g660(.A1(new_n686), .A2(new_n688), .A3(new_n733), .ZN(new_n847));
  NAND2_X1  g661(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  INV_X1    g662(.A(new_n666), .ZN(new_n849));
  NAND4_X1  g663(.A1(new_n849), .A2(new_n588), .A3(new_n472), .A4(new_n847), .ZN(new_n850));
  NAND3_X1  g664(.A1(new_n697), .A2(new_n608), .A3(new_n605), .ZN(new_n851));
  OAI22_X1  g665(.A1(new_n848), .A2(new_n723), .B1(new_n850), .B2(new_n851), .ZN(new_n852));
  INV_X1    g666(.A(new_n716), .ZN(new_n853));
  NAND2_X1  g667(.A1(new_n846), .A2(new_n853), .ZN(new_n854));
  INV_X1    g668(.A(KEYINPUT50), .ZN(new_n855));
  AND4_X1   g669(.A1(new_n647), .A2(new_n646), .A3(new_n688), .A4(new_n686), .ZN(new_n856));
  INV_X1    g670(.A(new_n856), .ZN(new_n857));
  NOR3_X1   g671(.A1(new_n854), .A2(new_n855), .A3(new_n857), .ZN(new_n858));
  XOR2_X1   g672(.A(new_n858), .B(KEYINPUT114), .Z(new_n859));
  OAI21_X1  g673(.A(new_n855), .B1(new_n854), .B2(new_n857), .ZN(new_n860));
  XNOR2_X1  g674(.A(new_n860), .B(KEYINPUT113), .ZN(new_n861));
  AOI21_X1  g675(.A(new_n852), .B1(new_n859), .B2(new_n861), .ZN(new_n862));
  NAND2_X1  g676(.A1(new_n684), .A2(new_n353), .ZN(new_n863));
  NOR2_X1   g677(.A1(new_n863), .A2(new_n191), .ZN(new_n864));
  OR2_X1    g678(.A1(new_n774), .A2(new_n787), .ZN(new_n865));
  AOI21_X1  g679(.A(new_n864), .B1(new_n865), .B2(new_n784), .ZN(new_n866));
  INV_X1    g680(.A(KEYINPUT115), .ZN(new_n867));
  AND2_X1   g681(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  NOR2_X1   g682(.A1(new_n854), .A2(new_n775), .ZN(new_n869));
  OAI21_X1  g683(.A(new_n869), .B1(new_n866), .B2(new_n867), .ZN(new_n870));
  OAI211_X1 g684(.A(new_n862), .B(KEYINPUT51), .C1(new_n868), .C2(new_n870), .ZN(new_n871));
  AND2_X1   g685(.A1(new_n742), .A2(new_n744), .ZN(new_n872));
  NOR2_X1   g686(.A1(new_n848), .A2(new_n872), .ZN(new_n873));
  XNOR2_X1  g687(.A(new_n873), .B(KEYINPUT48), .ZN(new_n874));
  NOR2_X1   g688(.A1(new_n471), .A2(G953), .ZN(new_n875));
  OAI221_X1 g689(.A(new_n875), .B1(new_n850), .B2(new_n610), .C1(new_n854), .C2(new_n689), .ZN(new_n876));
  NOR2_X1   g690(.A1(new_n874), .A2(new_n876), .ZN(new_n877));
  OR3_X1    g691(.A1(new_n866), .A2(new_n775), .A3(new_n854), .ZN(new_n878));
  AND2_X1   g692(.A1(new_n862), .A2(new_n878), .ZN(new_n879));
  OAI211_X1 g693(.A(new_n871), .B(new_n877), .C1(new_n879), .C2(KEYINPUT51), .ZN(new_n880));
  OAI22_X1  g694(.A1(new_n845), .A2(new_n880), .B1(G952), .B2(G953), .ZN(new_n881));
  NAND4_X1  g695(.A1(new_n646), .A2(new_n588), .A3(new_n191), .A4(new_n192), .ZN(new_n882));
  XNOR2_X1  g696(.A(new_n863), .B(KEYINPUT49), .ZN(new_n883));
  OR4_X1    g697(.A1(new_n666), .A2(new_n882), .A3(new_n883), .A4(new_n751), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n881), .A2(new_n884), .ZN(G75));
  OAI21_X1  g699(.A(new_n837), .B1(new_n805), .B2(new_n828), .ZN(new_n886));
  NAND3_X1  g700(.A1(new_n886), .A2(G902), .A3(new_n278), .ZN(new_n887));
  INV_X1    g701(.A(KEYINPUT116), .ZN(new_n888));
  NOR2_X1   g702(.A1(new_n888), .A2(KEYINPUT56), .ZN(new_n889));
  NAND2_X1  g703(.A1(new_n887), .A2(new_n889), .ZN(new_n890));
  NAND2_X1  g704(.A1(new_n272), .A2(new_n275), .ZN(new_n891));
  XNOR2_X1  g705(.A(new_n891), .B(new_n273), .ZN(new_n892));
  XOR2_X1   g706(.A(new_n892), .B(KEYINPUT55), .Z(new_n893));
  NAND2_X1  g707(.A1(new_n890), .A2(new_n893), .ZN(new_n894));
  INV_X1    g708(.A(new_n893), .ZN(new_n895));
  NAND3_X1  g709(.A1(new_n887), .A2(new_n889), .A3(new_n895), .ZN(new_n896));
  NOR2_X1   g710(.A1(new_n320), .A2(G952), .ZN(new_n897));
  INV_X1    g711(.A(new_n897), .ZN(new_n898));
  NAND3_X1  g712(.A1(new_n894), .A2(new_n896), .A3(new_n898), .ZN(new_n899));
  INV_X1    g713(.A(KEYINPUT117), .ZN(new_n900));
  NAND2_X1  g714(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  NAND4_X1  g715(.A1(new_n894), .A2(KEYINPUT117), .A3(new_n896), .A4(new_n898), .ZN(new_n902));
  NAND2_X1  g716(.A1(new_n901), .A2(new_n902), .ZN(G51));
  XOR2_X1   g717(.A(new_n354), .B(KEYINPUT57), .Z(new_n904));
  INV_X1    g718(.A(new_n838), .ZN(new_n905));
  AND2_X1   g719(.A1(new_n886), .A2(KEYINPUT54), .ZN(new_n906));
  OAI21_X1  g720(.A(new_n904), .B1(new_n905), .B2(new_n906), .ZN(new_n907));
  XNOR2_X1  g721(.A(new_n683), .B(KEYINPUT118), .ZN(new_n908));
  NAND2_X1  g722(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  INV_X1    g723(.A(new_n764), .ZN(new_n910));
  NAND3_X1  g724(.A1(new_n886), .A2(G902), .A3(new_n910), .ZN(new_n911));
  AOI21_X1  g725(.A(new_n897), .B1(new_n909), .B2(new_n911), .ZN(G54));
  AND2_X1   g726(.A1(KEYINPUT58), .A2(G475), .ZN(new_n913));
  NAND4_X1  g727(.A1(new_n886), .A2(G902), .A3(new_n425), .A4(new_n913), .ZN(new_n914));
  AND2_X1   g728(.A1(new_n914), .A2(new_n898), .ZN(new_n915));
  NAND3_X1  g729(.A1(new_n886), .A2(G902), .A3(new_n913), .ZN(new_n916));
  INV_X1    g730(.A(KEYINPUT119), .ZN(new_n917));
  INV_X1    g731(.A(new_n425), .ZN(new_n918));
  AND3_X1   g732(.A1(new_n916), .A2(new_n917), .A3(new_n918), .ZN(new_n919));
  AOI21_X1  g733(.A(new_n917), .B1(new_n916), .B2(new_n918), .ZN(new_n920));
  OAI21_X1  g734(.A(new_n915), .B1(new_n919), .B2(new_n920), .ZN(new_n921));
  NAND2_X1  g735(.A1(new_n921), .A2(KEYINPUT120), .ZN(new_n922));
  INV_X1    g736(.A(KEYINPUT120), .ZN(new_n923));
  OAI211_X1 g737(.A(new_n923), .B(new_n915), .C1(new_n919), .C2(new_n920), .ZN(new_n924));
  NAND2_X1  g738(.A1(new_n922), .A2(new_n924), .ZN(G60));
  NAND2_X1  g739(.A1(G478), .A2(G902), .ZN(new_n926));
  XNOR2_X1  g740(.A(new_n926), .B(KEYINPUT59), .ZN(new_n927));
  AOI21_X1  g741(.A(new_n604), .B1(new_n845), .B2(new_n927), .ZN(new_n928));
  OAI211_X1 g742(.A(new_n604), .B(new_n927), .C1(new_n905), .C2(new_n906), .ZN(new_n929));
  NAND2_X1  g743(.A1(new_n929), .A2(new_n898), .ZN(new_n930));
  NOR2_X1   g744(.A1(new_n928), .A2(new_n930), .ZN(G63));
  NAND2_X1  g745(.A1(G217), .A2(G902), .ZN(new_n932));
  XOR2_X1   g746(.A(new_n932), .B(KEYINPUT60), .Z(new_n933));
  NAND2_X1  g747(.A1(new_n886), .A2(new_n933), .ZN(new_n934));
  AOI21_X1  g748(.A(new_n897), .B1(new_n934), .B2(new_n579), .ZN(new_n935));
  NAND3_X1  g749(.A1(new_n886), .A2(new_n628), .A3(new_n933), .ZN(new_n936));
  NAND2_X1  g750(.A1(new_n935), .A2(new_n936), .ZN(new_n937));
  NAND2_X1  g751(.A1(KEYINPUT121), .A2(KEYINPUT61), .ZN(new_n938));
  INV_X1    g752(.A(KEYINPUT121), .ZN(new_n939));
  INV_X1    g753(.A(KEYINPUT61), .ZN(new_n940));
  NAND2_X1  g754(.A1(new_n939), .A2(new_n940), .ZN(new_n941));
  AND3_X1   g755(.A1(new_n937), .A2(new_n938), .A3(new_n941), .ZN(new_n942));
  AOI21_X1  g756(.A(new_n941), .B1(new_n937), .B2(new_n938), .ZN(new_n943));
  NOR2_X1   g757(.A1(new_n942), .A2(new_n943), .ZN(G66));
  OR2_X1    g758(.A1(new_n813), .A2(new_n823), .ZN(new_n945));
  NAND2_X1  g759(.A1(new_n945), .A2(new_n320), .ZN(new_n946));
  OAI21_X1  g760(.A(G953), .B1(new_n469), .B2(new_n243), .ZN(new_n947));
  NAND2_X1  g761(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  OAI21_X1  g762(.A(new_n891), .B1(G898), .B2(new_n320), .ZN(new_n949));
  XNOR2_X1  g763(.A(new_n949), .B(KEYINPUT122), .ZN(new_n950));
  XNOR2_X1  g764(.A(new_n948), .B(new_n950), .ZN(G69));
  AOI21_X1  g765(.A(new_n320), .B1(G227), .B2(G900), .ZN(new_n952));
  NOR2_X1   g766(.A1(new_n952), .A2(KEYINPUT125), .ZN(new_n953));
  INV_X1    g767(.A(new_n952), .ZN(new_n954));
  INV_X1    g768(.A(KEYINPUT125), .ZN(new_n955));
  NOR2_X1   g769(.A1(new_n954), .A2(new_n955), .ZN(new_n956));
  NOR3_X1   g770(.A1(new_n872), .A2(new_n282), .A3(new_n710), .ZN(new_n957));
  NAND3_X1  g771(.A1(new_n774), .A2(new_n957), .A3(new_n650), .ZN(new_n958));
  OAI211_X1 g772(.A(new_n788), .B(new_n958), .C1(new_n779), .C2(new_n757), .ZN(new_n959));
  AND2_X1   g773(.A1(new_n792), .A2(new_n677), .ZN(new_n960));
  NAND2_X1  g774(.A1(new_n960), .A2(new_n799), .ZN(new_n961));
  NOR2_X1   g775(.A1(new_n959), .A2(new_n961), .ZN(new_n962));
  NAND2_X1  g776(.A1(new_n808), .A2(new_n748), .ZN(new_n963));
  INV_X1    g777(.A(KEYINPUT124), .ZN(new_n964));
  XNOR2_X1  g778(.A(new_n963), .B(new_n964), .ZN(new_n965));
  NAND2_X1  g779(.A1(new_n962), .A2(new_n965), .ZN(new_n966));
  NAND2_X1  g780(.A1(new_n509), .A2(new_n514), .ZN(new_n967));
  XOR2_X1   g781(.A(new_n967), .B(KEYINPUT123), .Z(new_n968));
  NAND2_X1  g782(.A1(new_n411), .A2(new_n412), .ZN(new_n969));
  XOR2_X1   g783(.A(new_n968), .B(new_n969), .Z(new_n970));
  INV_X1    g784(.A(new_n970), .ZN(new_n971));
  AOI21_X1  g785(.A(G953), .B1(new_n966), .B2(new_n971), .ZN(new_n972));
  NAND3_X1  g786(.A1(new_n960), .A2(new_n668), .A3(new_n799), .ZN(new_n973));
  INV_X1    g787(.A(KEYINPUT62), .ZN(new_n974));
  XNOR2_X1  g788(.A(new_n973), .B(new_n974), .ZN(new_n975));
  NAND4_X1  g789(.A1(new_n729), .A2(new_n652), .A3(new_n733), .A4(new_n820), .ZN(new_n976));
  AND3_X1   g790(.A1(new_n780), .A2(new_n788), .A3(new_n976), .ZN(new_n977));
  NAND3_X1  g791(.A1(new_n975), .A2(new_n970), .A3(new_n977), .ZN(new_n978));
  NAND2_X1  g792(.A1(new_n972), .A2(new_n978), .ZN(new_n979));
  NAND3_X1  g793(.A1(new_n971), .A2(G900), .A3(G953), .ZN(new_n980));
  AOI211_X1 g794(.A(new_n953), .B(new_n956), .C1(new_n979), .C2(new_n980), .ZN(new_n981));
  AND4_X1   g795(.A1(new_n955), .A2(new_n979), .A3(new_n954), .A4(new_n980), .ZN(new_n982));
  NOR2_X1   g796(.A1(new_n981), .A2(new_n982), .ZN(G72));
  OR3_X1    g797(.A1(new_n966), .A2(new_n504), .A3(new_n516), .ZN(new_n984));
  NAND3_X1  g798(.A1(new_n975), .A2(new_n656), .A3(new_n977), .ZN(new_n985));
  AOI21_X1  g799(.A(new_n945), .B1(new_n984), .B2(new_n985), .ZN(new_n986));
  AND2_X1   g800(.A1(new_n517), .A2(new_n525), .ZN(new_n987));
  XOR2_X1   g801(.A(KEYINPUT126), .B(KEYINPUT63), .Z(new_n988));
  NAND2_X1  g802(.A1(G472), .A2(G902), .ZN(new_n989));
  XNOR2_X1  g803(.A(new_n988), .B(new_n989), .ZN(new_n990));
  XOR2_X1   g804(.A(new_n990), .B(KEYINPUT127), .Z(new_n991));
  AOI21_X1  g805(.A(new_n897), .B1(new_n987), .B2(new_n991), .ZN(new_n992));
  NAND2_X1  g806(.A1(new_n842), .A2(new_n843), .ZN(new_n993));
  OR2_X1    g807(.A1(new_n987), .A2(new_n990), .ZN(new_n994));
  OAI21_X1  g808(.A(new_n992), .B1(new_n993), .B2(new_n994), .ZN(new_n995));
  NOR2_X1   g809(.A1(new_n986), .A2(new_n995), .ZN(G57));
endmodule


