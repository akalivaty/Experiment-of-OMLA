//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 0 1 1 1 0 0 0 0 0 1 0 0 1 0 0 1 0 1 0 1 0 0 0 1 1 1 1 1 0 1 0 1 1 1 0 1 0 1 1 0 0 0 1 1 0 1 0 1 0 0 1 1 1 0 0 1 0 0 1 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:19:32 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n689, new_n690, new_n691, new_n692,
    new_n693, new_n694, new_n695, new_n696, new_n697, new_n698, new_n699,
    new_n701, new_n702, new_n703, new_n704, new_n705, new_n706, new_n707,
    new_n709, new_n710, new_n711, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n739, new_n740, new_n741, new_n742, new_n743, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n781, new_n782, new_n783, new_n784, new_n786,
    new_n788, new_n789, new_n790, new_n791, new_n792, new_n793, new_n794,
    new_n795, new_n796, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n804, new_n805, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n857, new_n858, new_n859, new_n861, new_n862, new_n863,
    new_n865, new_n866, new_n867, new_n868, new_n869, new_n870, new_n871,
    new_n872, new_n873, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n925, new_n926, new_n928, new_n929, new_n930, new_n931,
    new_n932, new_n933, new_n934, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n944, new_n945, new_n946, new_n948,
    new_n949, new_n950, new_n951, new_n952, new_n953, new_n954, new_n955,
    new_n957, new_n958, new_n959, new_n960, new_n961, new_n962, new_n963,
    new_n964, new_n965, new_n967, new_n968, new_n969, new_n970, new_n971,
    new_n972, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n981, new_n982, new_n983, new_n984, new_n985, new_n986, new_n987,
    new_n988, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001;
  NAND2_X1  g000(.A1(G229gat), .A2(G233gat), .ZN(new_n202));
  INV_X1    g001(.A(KEYINPUT16), .ZN(new_n203));
  NOR2_X1   g002(.A1(new_n203), .A2(G1gat), .ZN(new_n204));
  OR2_X1    g003(.A1(G15gat), .A2(G22gat), .ZN(new_n205));
  NAND2_X1  g004(.A1(G15gat), .A2(G22gat), .ZN(new_n206));
  NAND3_X1  g005(.A1(new_n205), .A2(KEYINPUT88), .A3(new_n206), .ZN(new_n207));
  INV_X1    g006(.A(KEYINPUT88), .ZN(new_n208));
  AND2_X1   g007(.A1(G15gat), .A2(G22gat), .ZN(new_n209));
  NOR2_X1   g008(.A1(G15gat), .A2(G22gat), .ZN(new_n210));
  OAI21_X1  g009(.A(new_n208), .B1(new_n209), .B2(new_n210), .ZN(new_n211));
  AOI21_X1  g010(.A(new_n204), .B1(new_n207), .B2(new_n211), .ZN(new_n212));
  INV_X1    g011(.A(KEYINPUT89), .ZN(new_n213));
  XNOR2_X1  g012(.A(new_n212), .B(new_n213), .ZN(new_n214));
  INV_X1    g013(.A(G1gat), .ZN(new_n215));
  NAND3_X1  g014(.A1(new_n207), .A2(new_n211), .A3(new_n215), .ZN(new_n216));
  XOR2_X1   g015(.A(KEYINPUT90), .B(G8gat), .Z(new_n217));
  AND2_X1   g016(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n207), .A2(new_n211), .ZN(new_n219));
  INV_X1    g018(.A(new_n204), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n221), .A2(new_n216), .ZN(new_n222));
  AOI22_X1  g021(.A1(new_n214), .A2(new_n218), .B1(G8gat), .B2(new_n222), .ZN(new_n223));
  INV_X1    g022(.A(G29gat), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n224), .A2(KEYINPUT85), .ZN(new_n225));
  INV_X1    g024(.A(KEYINPUT85), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n226), .A2(G29gat), .ZN(new_n227));
  NAND3_X1  g026(.A1(new_n225), .A2(new_n227), .A3(G36gat), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n228), .A2(KEYINPUT86), .ZN(new_n229));
  XNOR2_X1  g028(.A(KEYINPUT85), .B(G29gat), .ZN(new_n230));
  INV_X1    g029(.A(KEYINPUT86), .ZN(new_n231));
  NAND3_X1  g030(.A1(new_n230), .A2(new_n231), .A3(G36gat), .ZN(new_n232));
  NOR2_X1   g031(.A1(G29gat), .A2(G36gat), .ZN(new_n233));
  INV_X1    g032(.A(KEYINPUT14), .ZN(new_n234));
  XNOR2_X1  g033(.A(new_n233), .B(new_n234), .ZN(new_n235));
  NAND3_X1  g034(.A1(new_n229), .A2(new_n232), .A3(new_n235), .ZN(new_n236));
  INV_X1    g035(.A(G43gat), .ZN(new_n237));
  OAI21_X1  g036(.A(KEYINPUT15), .B1(new_n237), .B2(G50gat), .ZN(new_n238));
  AOI21_X1  g037(.A(new_n238), .B1(new_n237), .B2(G50gat), .ZN(new_n239));
  INV_X1    g038(.A(new_n239), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n236), .A2(new_n240), .ZN(new_n241));
  OR2_X1    g040(.A1(new_n237), .A2(G50gat), .ZN(new_n242));
  XNOR2_X1  g041(.A(KEYINPUT87), .B(G50gat), .ZN(new_n243));
  OAI21_X1  g042(.A(new_n242), .B1(new_n243), .B2(G43gat), .ZN(new_n244));
  INV_X1    g043(.A(KEYINPUT15), .ZN(new_n245));
  AOI21_X1  g044(.A(new_n239), .B1(new_n244), .B2(new_n245), .ZN(new_n246));
  OAI21_X1  g045(.A(new_n241), .B1(new_n236), .B2(new_n246), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n247), .A2(KEYINPUT17), .ZN(new_n248));
  INV_X1    g047(.A(KEYINPUT17), .ZN(new_n249));
  OAI211_X1 g048(.A(new_n241), .B(new_n249), .C1(new_n236), .C2(new_n246), .ZN(new_n250));
  NAND3_X1  g049(.A1(new_n223), .A2(new_n248), .A3(new_n250), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n221), .A2(new_n213), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n212), .A2(KEYINPUT89), .ZN(new_n253));
  NAND3_X1  g052(.A1(new_n252), .A2(new_n218), .A3(new_n253), .ZN(new_n254));
  NAND2_X1  g053(.A1(new_n222), .A2(G8gat), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n254), .A2(new_n255), .ZN(new_n256));
  AND2_X1   g055(.A1(new_n236), .A2(new_n240), .ZN(new_n257));
  NOR2_X1   g056(.A1(new_n246), .A2(new_n236), .ZN(new_n258));
  NOR2_X1   g057(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  INV_X1    g058(.A(KEYINPUT91), .ZN(new_n260));
  AND3_X1   g059(.A1(new_n256), .A2(new_n259), .A3(new_n260), .ZN(new_n261));
  AOI21_X1  g060(.A(new_n260), .B1(new_n256), .B2(new_n259), .ZN(new_n262));
  OAI211_X1 g061(.A(new_n202), .B(new_n251), .C1(new_n261), .C2(new_n262), .ZN(new_n263));
  INV_X1    g062(.A(KEYINPUT18), .ZN(new_n264));
  NAND3_X1  g063(.A1(new_n263), .A2(KEYINPUT92), .A3(new_n264), .ZN(new_n265));
  XOR2_X1   g064(.A(new_n202), .B(KEYINPUT13), .Z(new_n266));
  NOR2_X1   g065(.A1(new_n261), .A2(new_n262), .ZN(new_n267));
  NAND3_X1  g066(.A1(new_n223), .A2(KEYINPUT93), .A3(new_n247), .ZN(new_n268));
  INV_X1    g067(.A(KEYINPUT93), .ZN(new_n269));
  OAI21_X1  g068(.A(new_n269), .B1(new_n256), .B2(new_n259), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n268), .A2(new_n270), .ZN(new_n271));
  OAI21_X1  g070(.A(new_n266), .B1(new_n267), .B2(new_n271), .ZN(new_n272));
  OAI21_X1  g071(.A(KEYINPUT91), .B1(new_n223), .B2(new_n247), .ZN(new_n273));
  NAND3_X1  g072(.A1(new_n256), .A2(new_n259), .A3(new_n260), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  NAND2_X1  g074(.A1(new_n264), .A2(KEYINPUT92), .ZN(new_n276));
  NAND4_X1  g075(.A1(new_n275), .A2(new_n202), .A3(new_n251), .A4(new_n276), .ZN(new_n277));
  NAND3_X1  g076(.A1(new_n265), .A2(new_n272), .A3(new_n277), .ZN(new_n278));
  XNOR2_X1  g077(.A(G113gat), .B(G141gat), .ZN(new_n279));
  XNOR2_X1  g078(.A(KEYINPUT84), .B(KEYINPUT11), .ZN(new_n280));
  XNOR2_X1  g079(.A(new_n279), .B(new_n280), .ZN(new_n281));
  XNOR2_X1  g080(.A(G169gat), .B(G197gat), .ZN(new_n282));
  XNOR2_X1  g081(.A(new_n281), .B(new_n282), .ZN(new_n283));
  XNOR2_X1  g082(.A(new_n283), .B(KEYINPUT12), .ZN(new_n284));
  INV_X1    g083(.A(new_n284), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n278), .A2(new_n285), .ZN(new_n286));
  NAND4_X1  g085(.A1(new_n265), .A2(new_n272), .A3(new_n277), .A4(new_n284), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  INV_X1    g087(.A(new_n288), .ZN(new_n289));
  NAND2_X1  g088(.A1(G211gat), .A2(G218gat), .ZN(new_n290));
  AND2_X1   g089(.A1(KEYINPUT73), .A2(KEYINPUT22), .ZN(new_n291));
  NOR2_X1   g090(.A1(KEYINPUT73), .A2(KEYINPUT22), .ZN(new_n292));
  OAI21_X1  g091(.A(new_n290), .B1(new_n291), .B2(new_n292), .ZN(new_n293));
  XNOR2_X1  g092(.A(G211gat), .B(G218gat), .ZN(new_n294));
  XNOR2_X1  g093(.A(G197gat), .B(G204gat), .ZN(new_n295));
  NAND3_X1  g094(.A1(new_n293), .A2(new_n294), .A3(new_n295), .ZN(new_n296));
  NAND2_X1  g095(.A1(new_n296), .A2(KEYINPUT74), .ZN(new_n297));
  INV_X1    g096(.A(new_n294), .ZN(new_n298));
  INV_X1    g097(.A(new_n295), .ZN(new_n299));
  OR2_X1    g098(.A1(new_n291), .A2(new_n292), .ZN(new_n300));
  OAI21_X1  g099(.A(new_n298), .B1(new_n299), .B2(new_n300), .ZN(new_n301));
  INV_X1    g100(.A(KEYINPUT74), .ZN(new_n302));
  NAND4_X1  g101(.A1(new_n293), .A2(new_n302), .A3(new_n294), .A4(new_n295), .ZN(new_n303));
  NAND3_X1  g102(.A1(new_n297), .A2(new_n301), .A3(new_n303), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n304), .A2(KEYINPUT75), .ZN(new_n305));
  INV_X1    g104(.A(KEYINPUT75), .ZN(new_n306));
  NAND4_X1  g105(.A1(new_n297), .A2(new_n306), .A3(new_n301), .A4(new_n303), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n305), .A2(new_n307), .ZN(new_n308));
  INV_X1    g107(.A(KEYINPUT76), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n308), .A2(new_n309), .ZN(new_n310));
  NAND3_X1  g109(.A1(new_n305), .A2(KEYINPUT76), .A3(new_n307), .ZN(new_n311));
  AND3_X1   g110(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n312));
  AOI21_X1  g111(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n313));
  NOR2_X1   g112(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  INV_X1    g113(.A(G190gat), .ZN(new_n315));
  AND2_X1   g114(.A1(KEYINPUT66), .A2(G183gat), .ZN(new_n316));
  NOR2_X1   g115(.A1(KEYINPUT66), .A2(G183gat), .ZN(new_n317));
  OAI21_X1  g116(.A(new_n315), .B1(new_n316), .B2(new_n317), .ZN(new_n318));
  AND2_X1   g117(.A1(new_n314), .A2(new_n318), .ZN(new_n319));
  OAI21_X1  g118(.A(KEYINPUT64), .B1(G169gat), .B2(G176gat), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n320), .A2(KEYINPUT23), .ZN(new_n321));
  NAND2_X1  g120(.A1(G169gat), .A2(G176gat), .ZN(new_n322));
  INV_X1    g121(.A(KEYINPUT23), .ZN(new_n323));
  OAI211_X1 g122(.A(new_n323), .B(KEYINPUT64), .C1(G169gat), .C2(G176gat), .ZN(new_n324));
  NAND3_X1  g123(.A1(new_n321), .A2(new_n322), .A3(new_n324), .ZN(new_n325));
  OAI21_X1  g124(.A(KEYINPUT25), .B1(new_n319), .B2(new_n325), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n325), .A2(KEYINPUT65), .ZN(new_n327));
  INV_X1    g126(.A(G183gat), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n328), .A2(new_n315), .ZN(new_n329));
  AOI21_X1  g128(.A(KEYINPUT25), .B1(new_n314), .B2(new_n329), .ZN(new_n330));
  INV_X1    g129(.A(KEYINPUT65), .ZN(new_n331));
  NAND4_X1  g130(.A1(new_n321), .A2(new_n331), .A3(new_n324), .A4(new_n322), .ZN(new_n332));
  NAND3_X1  g131(.A1(new_n327), .A2(new_n330), .A3(new_n332), .ZN(new_n333));
  AND2_X1   g132(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n334));
  NOR2_X1   g133(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n335));
  OAI211_X1 g134(.A(KEYINPUT28), .B(new_n315), .C1(new_n334), .C2(new_n335), .ZN(new_n336));
  INV_X1    g135(.A(new_n336), .ZN(new_n337));
  INV_X1    g136(.A(KEYINPUT27), .ZN(new_n338));
  NOR3_X1   g137(.A1(new_n316), .A2(new_n317), .A3(new_n338), .ZN(new_n339));
  OAI21_X1  g138(.A(new_n315), .B1(new_n339), .B2(new_n335), .ZN(new_n340));
  INV_X1    g139(.A(KEYINPUT28), .ZN(new_n341));
  AOI21_X1  g140(.A(new_n337), .B1(new_n340), .B2(new_n341), .ZN(new_n342));
  INV_X1    g141(.A(G169gat), .ZN(new_n343));
  INV_X1    g142(.A(G176gat), .ZN(new_n344));
  AOI21_X1  g143(.A(KEYINPUT26), .B1(new_n343), .B2(new_n344), .ZN(new_n345));
  AND2_X1   g144(.A1(new_n345), .A2(new_n322), .ZN(new_n346));
  NAND3_X1  g145(.A1(new_n343), .A2(new_n344), .A3(KEYINPUT26), .ZN(new_n347));
  OAI21_X1  g146(.A(new_n347), .B1(new_n328), .B2(new_n315), .ZN(new_n348));
  NOR2_X1   g147(.A1(new_n346), .A2(new_n348), .ZN(new_n349));
  INV_X1    g148(.A(new_n349), .ZN(new_n350));
  OAI211_X1 g149(.A(new_n326), .B(new_n333), .C1(new_n342), .C2(new_n350), .ZN(new_n351));
  INV_X1    g150(.A(G226gat), .ZN(new_n352));
  INV_X1    g151(.A(G233gat), .ZN(new_n353));
  NOR2_X1   g152(.A1(new_n352), .A2(new_n353), .ZN(new_n354));
  NOR2_X1   g153(.A1(new_n351), .A2(new_n354), .ZN(new_n355));
  NOR2_X1   g154(.A1(new_n354), .A2(KEYINPUT29), .ZN(new_n356));
  INV_X1    g155(.A(KEYINPUT66), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n357), .A2(new_n328), .ZN(new_n358));
  NAND2_X1  g157(.A1(KEYINPUT66), .A2(G183gat), .ZN(new_n359));
  NAND3_X1  g158(.A1(new_n358), .A2(KEYINPUT27), .A3(new_n359), .ZN(new_n360));
  INV_X1    g159(.A(new_n335), .ZN(new_n361));
  AOI21_X1  g160(.A(G190gat), .B1(new_n360), .B2(new_n361), .ZN(new_n362));
  OAI21_X1  g161(.A(new_n336), .B1(new_n362), .B2(KEYINPUT28), .ZN(new_n363));
  AND3_X1   g162(.A1(new_n321), .A2(new_n322), .A3(new_n324), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n314), .A2(new_n318), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  AOI22_X1  g165(.A1(new_n363), .A2(new_n349), .B1(KEYINPUT25), .B2(new_n366), .ZN(new_n367));
  AOI21_X1  g166(.A(new_n356), .B1(new_n367), .B2(new_n333), .ZN(new_n368));
  OAI211_X1 g167(.A(new_n310), .B(new_n311), .C1(new_n355), .C2(new_n368), .ZN(new_n369));
  XNOR2_X1  g168(.A(G8gat), .B(G36gat), .ZN(new_n370));
  INV_X1    g169(.A(G64gat), .ZN(new_n371));
  XNOR2_X1  g170(.A(new_n370), .B(new_n371), .ZN(new_n372));
  INV_X1    g171(.A(G92gat), .ZN(new_n373));
  XNOR2_X1  g172(.A(new_n372), .B(new_n373), .ZN(new_n374));
  INV_X1    g173(.A(new_n374), .ZN(new_n375));
  INV_X1    g174(.A(new_n356), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n351), .A2(new_n376), .ZN(new_n377));
  INV_X1    g176(.A(new_n354), .ZN(new_n378));
  NAND3_X1  g177(.A1(new_n367), .A2(new_n333), .A3(new_n378), .ZN(new_n379));
  NAND3_X1  g178(.A1(new_n377), .A2(new_n379), .A3(new_n308), .ZN(new_n380));
  AND3_X1   g179(.A1(new_n369), .A2(new_n375), .A3(new_n380), .ZN(new_n381));
  AOI21_X1  g180(.A(new_n375), .B1(new_n369), .B2(new_n380), .ZN(new_n382));
  INV_X1    g181(.A(KEYINPUT30), .ZN(new_n383));
  NOR3_X1   g182(.A1(new_n381), .A2(new_n382), .A3(new_n383), .ZN(new_n384));
  AND3_X1   g183(.A1(new_n377), .A2(new_n308), .A3(new_n379), .ZN(new_n385));
  AND2_X1   g184(.A1(new_n310), .A2(new_n311), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n377), .A2(new_n379), .ZN(new_n387));
  AOI21_X1  g186(.A(new_n385), .B1(new_n386), .B2(new_n387), .ZN(new_n388));
  AND3_X1   g187(.A1(new_n388), .A2(new_n383), .A3(new_n375), .ZN(new_n389));
  NOR2_X1   g188(.A1(new_n384), .A2(new_n389), .ZN(new_n390));
  INV_X1    g189(.A(KEYINPUT68), .ZN(new_n391));
  XNOR2_X1  g190(.A(G127gat), .B(G134gat), .ZN(new_n392));
  XNOR2_X1  g191(.A(G113gat), .B(G120gat), .ZN(new_n393));
  AOI21_X1  g192(.A(KEYINPUT1), .B1(new_n393), .B2(KEYINPUT67), .ZN(new_n394));
  INV_X1    g193(.A(KEYINPUT67), .ZN(new_n395));
  INV_X1    g194(.A(G113gat), .ZN(new_n396));
  NOR2_X1   g195(.A1(new_n396), .A2(G120gat), .ZN(new_n397));
  INV_X1    g196(.A(G120gat), .ZN(new_n398));
  NOR2_X1   g197(.A1(new_n398), .A2(G113gat), .ZN(new_n399));
  OAI21_X1  g198(.A(new_n395), .B1(new_n397), .B2(new_n399), .ZN(new_n400));
  AOI211_X1 g199(.A(new_n391), .B(new_n392), .C1(new_n394), .C2(new_n400), .ZN(new_n401));
  INV_X1    g200(.A(KEYINPUT1), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n398), .A2(G113gat), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n396), .A2(G120gat), .ZN(new_n404));
  NAND3_X1  g203(.A1(new_n403), .A2(new_n404), .A3(KEYINPUT67), .ZN(new_n405));
  NAND3_X1  g204(.A1(new_n400), .A2(new_n402), .A3(new_n405), .ZN(new_n406));
  XOR2_X1   g205(.A(G127gat), .B(G134gat), .Z(new_n407));
  AOI21_X1  g206(.A(KEYINPUT68), .B1(new_n406), .B2(new_n407), .ZN(new_n408));
  NOR2_X1   g207(.A1(new_n401), .A2(new_n408), .ZN(new_n409));
  INV_X1    g208(.A(KEYINPUT79), .ZN(new_n410));
  AOI21_X1  g209(.A(KEYINPUT1), .B1(new_n407), .B2(KEYINPUT69), .ZN(new_n411));
  INV_X1    g210(.A(new_n393), .ZN(new_n412));
  OAI211_X1 g211(.A(new_n411), .B(new_n412), .C1(KEYINPUT69), .C2(new_n407), .ZN(new_n413));
  INV_X1    g212(.A(G141gat), .ZN(new_n414));
  NOR2_X1   g213(.A1(new_n414), .A2(G148gat), .ZN(new_n415));
  INV_X1    g214(.A(new_n415), .ZN(new_n416));
  XNOR2_X1  g215(.A(KEYINPUT78), .B(G141gat), .ZN(new_n417));
  INV_X1    g216(.A(G148gat), .ZN(new_n418));
  OAI21_X1  g217(.A(new_n416), .B1(new_n417), .B2(new_n418), .ZN(new_n419));
  NAND2_X1  g218(.A1(G155gat), .A2(G162gat), .ZN(new_n420));
  OR2_X1    g219(.A1(G155gat), .A2(G162gat), .ZN(new_n421));
  OAI21_X1  g220(.A(new_n420), .B1(new_n421), .B2(KEYINPUT2), .ZN(new_n422));
  NOR2_X1   g221(.A1(new_n418), .A2(G141gat), .ZN(new_n423));
  AND2_X1   g222(.A1(KEYINPUT77), .A2(KEYINPUT2), .ZN(new_n424));
  NOR2_X1   g223(.A1(KEYINPUT77), .A2(KEYINPUT2), .ZN(new_n425));
  OAI22_X1  g224(.A1(new_n415), .A2(new_n423), .B1(new_n424), .B2(new_n425), .ZN(new_n426));
  AND2_X1   g225(.A1(new_n421), .A2(new_n420), .ZN(new_n427));
  AOI22_X1  g226(.A1(new_n419), .A2(new_n422), .B1(new_n426), .B2(new_n427), .ZN(new_n428));
  NAND4_X1  g227(.A1(new_n409), .A2(new_n410), .A3(new_n413), .A4(new_n428), .ZN(new_n429));
  NAND2_X1  g228(.A1(new_n405), .A2(new_n402), .ZN(new_n430));
  NOR2_X1   g229(.A1(new_n393), .A2(KEYINPUT67), .ZN(new_n431));
  OAI21_X1  g230(.A(new_n407), .B1(new_n430), .B2(new_n431), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n432), .A2(new_n391), .ZN(new_n433));
  NAND3_X1  g232(.A1(new_n406), .A2(KEYINPUT68), .A3(new_n407), .ZN(new_n434));
  NAND4_X1  g233(.A1(new_n433), .A2(new_n413), .A3(new_n434), .A4(new_n428), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n435), .A2(KEYINPUT79), .ZN(new_n436));
  NAND2_X1  g235(.A1(G225gat), .A2(G233gat), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n437), .A2(KEYINPUT4), .ZN(new_n438));
  NAND3_X1  g237(.A1(new_n429), .A2(new_n436), .A3(new_n438), .ZN(new_n439));
  INV_X1    g238(.A(new_n435), .ZN(new_n440));
  XNOR2_X1  g239(.A(new_n428), .B(KEYINPUT3), .ZN(new_n441));
  NAND3_X1  g240(.A1(new_n433), .A2(new_n413), .A3(new_n434), .ZN(new_n442));
  AOI22_X1  g241(.A1(new_n440), .A2(KEYINPUT4), .B1(new_n441), .B2(new_n442), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n439), .A2(new_n443), .ZN(new_n444));
  INV_X1    g243(.A(new_n428), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n442), .A2(new_n445), .ZN(new_n446));
  NAND3_X1  g245(.A1(new_n429), .A2(new_n436), .A3(new_n446), .ZN(new_n447));
  INV_X1    g246(.A(new_n437), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n447), .A2(new_n448), .ZN(new_n449));
  NAND3_X1  g248(.A1(new_n444), .A2(new_n449), .A3(KEYINPUT5), .ZN(new_n450));
  INV_X1    g249(.A(KEYINPUT3), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n428), .A2(new_n451), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n445), .A2(KEYINPUT3), .ZN(new_n453));
  AND3_X1   g252(.A1(new_n442), .A2(new_n452), .A3(new_n453), .ZN(new_n454));
  INV_X1    g253(.A(KEYINPUT4), .ZN(new_n455));
  OAI21_X1  g254(.A(new_n435), .B1(new_n454), .B2(new_n455), .ZN(new_n456));
  NOR2_X1   g255(.A1(new_n448), .A2(KEYINPUT5), .ZN(new_n457));
  AND2_X1   g256(.A1(new_n429), .A2(new_n436), .ZN(new_n458));
  OAI211_X1 g257(.A(new_n456), .B(new_n457), .C1(new_n455), .C2(new_n458), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n450), .A2(new_n459), .ZN(new_n460));
  XNOR2_X1  g259(.A(KEYINPUT0), .B(G57gat), .ZN(new_n461));
  XNOR2_X1  g260(.A(new_n461), .B(G85gat), .ZN(new_n462));
  XNOR2_X1  g261(.A(G1gat), .B(G29gat), .ZN(new_n463));
  XOR2_X1   g262(.A(new_n462), .B(new_n463), .Z(new_n464));
  INV_X1    g263(.A(new_n464), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n460), .A2(new_n465), .ZN(new_n466));
  NAND3_X1  g265(.A1(new_n450), .A2(new_n459), .A3(new_n464), .ZN(new_n467));
  XNOR2_X1  g266(.A(KEYINPUT80), .B(KEYINPUT6), .ZN(new_n468));
  NAND3_X1  g267(.A1(new_n466), .A2(new_n467), .A3(new_n468), .ZN(new_n469));
  INV_X1    g268(.A(new_n468), .ZN(new_n470));
  NAND3_X1  g269(.A1(new_n460), .A2(new_n465), .A3(new_n470), .ZN(new_n471));
  AOI21_X1  g270(.A(new_n390), .B1(new_n469), .B2(new_n471), .ZN(new_n472));
  INV_X1    g271(.A(G227gat), .ZN(new_n473));
  NOR2_X1   g272(.A1(new_n473), .A2(new_n353), .ZN(new_n474));
  AND2_X1   g273(.A1(new_n351), .A2(new_n442), .ZN(new_n475));
  NOR2_X1   g274(.A1(new_n351), .A2(new_n442), .ZN(new_n476));
  OAI21_X1  g275(.A(new_n474), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  INV_X1    g276(.A(KEYINPUT70), .ZN(new_n478));
  INV_X1    g277(.A(KEYINPUT33), .ZN(new_n479));
  NAND3_X1  g278(.A1(new_n477), .A2(new_n478), .A3(new_n479), .ZN(new_n480));
  INV_X1    g279(.A(new_n474), .ZN(new_n481));
  NAND4_X1  g280(.A1(new_n409), .A2(new_n367), .A3(new_n413), .A4(new_n333), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n351), .A2(new_n442), .ZN(new_n483));
  AOI21_X1  g282(.A(new_n481), .B1(new_n482), .B2(new_n483), .ZN(new_n484));
  OAI21_X1  g283(.A(KEYINPUT70), .B1(new_n484), .B2(KEYINPUT33), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n477), .A2(KEYINPUT32), .ZN(new_n486));
  XNOR2_X1  g285(.A(G15gat), .B(G43gat), .ZN(new_n487));
  XNOR2_X1  g286(.A(new_n487), .B(G71gat), .ZN(new_n488));
  INV_X1    g287(.A(G99gat), .ZN(new_n489));
  XNOR2_X1  g288(.A(new_n488), .B(new_n489), .ZN(new_n490));
  NAND4_X1  g289(.A1(new_n480), .A2(new_n485), .A3(new_n486), .A4(new_n490), .ZN(new_n491));
  OR2_X1    g290(.A1(new_n490), .A2(KEYINPUT71), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n490), .A2(KEYINPUT71), .ZN(new_n493));
  NAND3_X1  g292(.A1(new_n492), .A2(KEYINPUT33), .A3(new_n493), .ZN(new_n494));
  NAND3_X1  g293(.A1(new_n477), .A2(KEYINPUT32), .A3(new_n494), .ZN(new_n495));
  NAND3_X1  g294(.A1(new_n482), .A2(new_n481), .A3(new_n483), .ZN(new_n496));
  XOR2_X1   g295(.A(new_n496), .B(KEYINPUT34), .Z(new_n497));
  AND3_X1   g296(.A1(new_n491), .A2(new_n495), .A3(new_n497), .ZN(new_n498));
  AOI21_X1  g297(.A(new_n497), .B1(new_n491), .B2(new_n495), .ZN(new_n499));
  NOR2_X1   g298(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  INV_X1    g299(.A(KEYINPUT29), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n452), .A2(new_n501), .ZN(new_n502));
  NAND3_X1  g301(.A1(new_n310), .A2(new_n502), .A3(new_n311), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n304), .A2(new_n501), .ZN(new_n504));
  AOI21_X1  g303(.A(new_n428), .B1(new_n504), .B2(new_n451), .ZN(new_n505));
  INV_X1    g304(.A(new_n505), .ZN(new_n506));
  NAND4_X1  g305(.A1(new_n503), .A2(G228gat), .A3(G233gat), .A4(new_n506), .ZN(new_n507));
  NAND2_X1  g306(.A1(G228gat), .A2(G233gat), .ZN(new_n508));
  AOI21_X1  g307(.A(new_n308), .B1(new_n501), .B2(new_n452), .ZN(new_n509));
  OAI21_X1  g308(.A(new_n508), .B1(new_n509), .B2(new_n505), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n507), .A2(new_n510), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n511), .A2(G22gat), .ZN(new_n512));
  INV_X1    g311(.A(G22gat), .ZN(new_n513));
  NAND3_X1  g312(.A1(new_n507), .A2(new_n510), .A3(new_n513), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n512), .A2(new_n514), .ZN(new_n515));
  XNOR2_X1  g314(.A(G78gat), .B(G106gat), .ZN(new_n516));
  XNOR2_X1  g315(.A(KEYINPUT31), .B(G50gat), .ZN(new_n517));
  XNOR2_X1  g316(.A(new_n516), .B(new_n517), .ZN(new_n518));
  AOI21_X1  g317(.A(new_n513), .B1(new_n507), .B2(new_n510), .ZN(new_n519));
  OAI21_X1  g318(.A(new_n518), .B1(new_n519), .B2(KEYINPUT81), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n515), .A2(new_n520), .ZN(new_n521));
  NAND4_X1  g320(.A1(new_n512), .A2(KEYINPUT81), .A3(new_n514), .A4(new_n518), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  INV_X1    g322(.A(KEYINPUT83), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n524), .A2(KEYINPUT35), .ZN(new_n525));
  NAND4_X1  g324(.A1(new_n472), .A2(new_n500), .A3(new_n523), .A4(new_n525), .ZN(new_n526));
  NOR2_X1   g325(.A1(new_n524), .A2(KEYINPUT35), .ZN(new_n527));
  INV_X1    g326(.A(new_n527), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n526), .A2(new_n528), .ZN(new_n529));
  NAND4_X1  g328(.A1(new_n472), .A2(new_n500), .A3(new_n523), .A4(new_n527), .ZN(new_n530));
  NAND2_X1  g329(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n441), .A2(new_n442), .ZN(new_n532));
  AOI21_X1  g331(.A(new_n440), .B1(new_n532), .B2(KEYINPUT4), .ZN(new_n533));
  AOI21_X1  g332(.A(new_n455), .B1(new_n429), .B2(new_n436), .ZN(new_n534));
  OAI21_X1  g333(.A(new_n448), .B1(new_n533), .B2(new_n534), .ZN(new_n535));
  NAND3_X1  g334(.A1(new_n458), .A2(new_n437), .A3(new_n446), .ZN(new_n536));
  AND3_X1   g335(.A1(new_n535), .A2(KEYINPUT39), .A3(new_n536), .ZN(new_n537));
  OAI21_X1  g336(.A(new_n464), .B1(new_n535), .B2(KEYINPUT39), .ZN(new_n538));
  INV_X1    g337(.A(KEYINPUT40), .ZN(new_n539));
  OR3_X1    g338(.A1(new_n537), .A2(new_n538), .A3(new_n539), .ZN(new_n540));
  OAI21_X1  g339(.A(new_n539), .B1(new_n537), .B2(new_n538), .ZN(new_n541));
  NAND4_X1  g340(.A1(new_n540), .A2(new_n466), .A3(new_n390), .A4(new_n541), .ZN(new_n542));
  INV_X1    g341(.A(KEYINPUT37), .ZN(new_n543));
  OAI211_X1 g342(.A(KEYINPUT82), .B(new_n374), .C1(new_n388), .C2(new_n543), .ZN(new_n544));
  INV_X1    g343(.A(KEYINPUT82), .ZN(new_n545));
  AOI21_X1  g344(.A(new_n543), .B1(new_n369), .B2(new_n380), .ZN(new_n546));
  OAI21_X1  g345(.A(new_n545), .B1(new_n546), .B2(new_n375), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n388), .A2(new_n543), .ZN(new_n548));
  NAND3_X1  g347(.A1(new_n544), .A2(new_n547), .A3(new_n548), .ZN(new_n549));
  NAND2_X1  g348(.A1(new_n549), .A2(KEYINPUT38), .ZN(new_n550));
  INV_X1    g349(.A(new_n381), .ZN(new_n551));
  NAND4_X1  g350(.A1(new_n550), .A2(new_n471), .A3(new_n469), .A4(new_n551), .ZN(new_n552));
  INV_X1    g351(.A(KEYINPUT38), .ZN(new_n553));
  AOI21_X1  g352(.A(new_n543), .B1(new_n387), .B2(new_n308), .ZN(new_n554));
  INV_X1    g353(.A(new_n386), .ZN(new_n555));
  OAI21_X1  g354(.A(new_n554), .B1(new_n555), .B2(new_n387), .ZN(new_n556));
  AND4_X1   g355(.A1(new_n553), .A2(new_n548), .A3(new_n374), .A4(new_n556), .ZN(new_n557));
  OAI211_X1 g356(.A(new_n523), .B(new_n542), .C1(new_n552), .C2(new_n557), .ZN(new_n558));
  NAND2_X1  g357(.A1(new_n491), .A2(new_n495), .ZN(new_n559));
  INV_X1    g358(.A(new_n497), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  NAND3_X1  g360(.A1(new_n491), .A2(new_n495), .A3(new_n497), .ZN(new_n562));
  NAND2_X1  g361(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  INV_X1    g362(.A(KEYINPUT72), .ZN(new_n564));
  AOI21_X1  g363(.A(KEYINPUT36), .B1(new_n563), .B2(new_n564), .ZN(new_n565));
  OAI211_X1 g364(.A(new_n564), .B(KEYINPUT36), .C1(new_n498), .C2(new_n499), .ZN(new_n566));
  INV_X1    g365(.A(new_n566), .ZN(new_n567));
  NOR2_X1   g366(.A1(new_n565), .A2(new_n567), .ZN(new_n568));
  OR2_X1    g367(.A1(new_n472), .A2(new_n523), .ZN(new_n569));
  NAND3_X1  g368(.A1(new_n558), .A2(new_n568), .A3(new_n569), .ZN(new_n570));
  AOI21_X1  g369(.A(new_n289), .B1(new_n531), .B2(new_n570), .ZN(new_n571));
  XNOR2_X1  g370(.A(G127gat), .B(G155gat), .ZN(new_n572));
  XOR2_X1   g371(.A(new_n572), .B(G211gat), .Z(new_n573));
  INV_X1    g372(.A(new_n573), .ZN(new_n574));
  INV_X1    g373(.A(KEYINPUT21), .ZN(new_n575));
  INV_X1    g374(.A(G57gat), .ZN(new_n576));
  OAI21_X1  g375(.A(KEYINPUT94), .B1(new_n576), .B2(G64gat), .ZN(new_n577));
  INV_X1    g376(.A(KEYINPUT94), .ZN(new_n578));
  NAND3_X1  g377(.A1(new_n578), .A2(new_n371), .A3(G57gat), .ZN(new_n579));
  NAND2_X1  g378(.A1(new_n576), .A2(G64gat), .ZN(new_n580));
  NAND3_X1  g379(.A1(new_n577), .A2(new_n579), .A3(new_n580), .ZN(new_n581));
  INV_X1    g380(.A(G71gat), .ZN(new_n582));
  INV_X1    g381(.A(G78gat), .ZN(new_n583));
  NAND2_X1  g382(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  NAND2_X1  g383(.A1(G71gat), .A2(G78gat), .ZN(new_n585));
  NAND2_X1  g384(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  INV_X1    g385(.A(KEYINPUT9), .ZN(new_n587));
  NAND2_X1  g386(.A1(new_n585), .A2(new_n587), .ZN(new_n588));
  INV_X1    g387(.A(KEYINPUT95), .ZN(new_n589));
  NAND2_X1  g388(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  NAND3_X1  g389(.A1(new_n585), .A2(KEYINPUT95), .A3(new_n587), .ZN(new_n591));
  NAND4_X1  g390(.A1(new_n581), .A2(new_n586), .A3(new_n590), .A4(new_n591), .ZN(new_n592));
  XNOR2_X1  g391(.A(G57gat), .B(G64gat), .ZN(new_n593));
  OAI211_X1 g392(.A(new_n585), .B(new_n584), .C1(new_n593), .C2(new_n587), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n592), .A2(new_n594), .ZN(new_n595));
  OAI211_X1 g394(.A(new_n254), .B(new_n255), .C1(new_n575), .C2(new_n595), .ZN(new_n596));
  NAND2_X1  g395(.A1(new_n596), .A2(G183gat), .ZN(new_n597));
  INV_X1    g396(.A(new_n597), .ZN(new_n598));
  NOR2_X1   g397(.A1(new_n596), .A2(G183gat), .ZN(new_n599));
  INV_X1    g398(.A(G231gat), .ZN(new_n600));
  OAI22_X1  g399(.A1(new_n598), .A2(new_n599), .B1(new_n600), .B2(new_n353), .ZN(new_n601));
  INV_X1    g400(.A(new_n599), .ZN(new_n602));
  NOR2_X1   g401(.A1(new_n600), .A2(new_n353), .ZN(new_n603));
  NAND3_X1  g402(.A1(new_n602), .A2(new_n597), .A3(new_n603), .ZN(new_n604));
  AOI21_X1  g403(.A(new_n574), .B1(new_n601), .B2(new_n604), .ZN(new_n605));
  INV_X1    g404(.A(new_n605), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n595), .A2(new_n575), .ZN(new_n607));
  XNOR2_X1  g406(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n608));
  XOR2_X1   g407(.A(new_n607), .B(new_n608), .Z(new_n609));
  NAND3_X1  g408(.A1(new_n601), .A2(new_n604), .A3(new_n574), .ZN(new_n610));
  NAND3_X1  g409(.A1(new_n606), .A2(new_n609), .A3(new_n610), .ZN(new_n611));
  INV_X1    g410(.A(new_n609), .ZN(new_n612));
  INV_X1    g411(.A(new_n610), .ZN(new_n613));
  OAI21_X1  g412(.A(new_n612), .B1(new_n613), .B2(new_n605), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n611), .A2(new_n614), .ZN(new_n615));
  XOR2_X1   g414(.A(G190gat), .B(G218gat), .Z(new_n616));
  INV_X1    g415(.A(new_n616), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n617), .A2(KEYINPUT97), .ZN(new_n618));
  XOR2_X1   g417(.A(G134gat), .B(G162gat), .Z(new_n619));
  XNOR2_X1  g418(.A(new_n618), .B(new_n619), .ZN(new_n620));
  INV_X1    g419(.A(new_n620), .ZN(new_n621));
  INV_X1    g420(.A(KEYINPUT96), .ZN(new_n622));
  NAND2_X1  g421(.A1(G99gat), .A2(G106gat), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n623), .A2(KEYINPUT8), .ZN(new_n624));
  NAND2_X1  g423(.A1(G85gat), .A2(G92gat), .ZN(new_n625));
  INV_X1    g424(.A(KEYINPUT7), .ZN(new_n626));
  NAND2_X1  g425(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  INV_X1    g426(.A(G85gat), .ZN(new_n628));
  NAND2_X1  g427(.A1(new_n628), .A2(new_n373), .ZN(new_n629));
  NAND3_X1  g428(.A1(KEYINPUT7), .A2(G85gat), .A3(G92gat), .ZN(new_n630));
  NAND4_X1  g429(.A1(new_n624), .A2(new_n627), .A3(new_n629), .A4(new_n630), .ZN(new_n631));
  XNOR2_X1  g430(.A(G99gat), .B(G106gat), .ZN(new_n632));
  INV_X1    g431(.A(new_n632), .ZN(new_n633));
  NOR2_X1   g432(.A1(new_n631), .A2(new_n633), .ZN(new_n634));
  INV_X1    g433(.A(new_n630), .ZN(new_n635));
  AOI21_X1  g434(.A(KEYINPUT7), .B1(G85gat), .B2(G92gat), .ZN(new_n636));
  NOR2_X1   g435(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  AOI22_X1  g436(.A1(KEYINPUT8), .A2(new_n623), .B1(new_n628), .B2(new_n373), .ZN(new_n638));
  AOI21_X1  g437(.A(new_n632), .B1(new_n637), .B2(new_n638), .ZN(new_n639));
  OAI21_X1  g438(.A(new_n622), .B1(new_n634), .B2(new_n639), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n631), .A2(new_n633), .ZN(new_n641));
  NAND3_X1  g440(.A1(new_n637), .A2(new_n632), .A3(new_n638), .ZN(new_n642));
  NAND3_X1  g441(.A1(new_n641), .A2(new_n642), .A3(KEYINPUT96), .ZN(new_n643));
  NAND2_X1  g442(.A1(new_n640), .A2(new_n643), .ZN(new_n644));
  NAND3_X1  g443(.A1(new_n248), .A2(new_n250), .A3(new_n644), .ZN(new_n645));
  NAND3_X1  g444(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n646));
  OAI211_X1 g445(.A(new_n645), .B(new_n646), .C1(new_n247), .C2(new_n644), .ZN(new_n647));
  OR2_X1    g446(.A1(new_n617), .A2(KEYINPUT97), .ZN(new_n648));
  AOI21_X1  g447(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n649));
  INV_X1    g448(.A(new_n649), .ZN(new_n650));
  NAND3_X1  g449(.A1(new_n647), .A2(new_n648), .A3(new_n650), .ZN(new_n651));
  INV_X1    g450(.A(new_n651), .ZN(new_n652));
  AOI21_X1  g451(.A(new_n650), .B1(new_n647), .B2(new_n648), .ZN(new_n653));
  OAI21_X1  g452(.A(new_n621), .B1(new_n652), .B2(new_n653), .ZN(new_n654));
  INV_X1    g453(.A(new_n653), .ZN(new_n655));
  NAND3_X1  g454(.A1(new_n655), .A2(new_n651), .A3(new_n620), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n654), .A2(new_n656), .ZN(new_n657));
  NAND2_X1  g456(.A1(G230gat), .A2(G233gat), .ZN(new_n658));
  INV_X1    g457(.A(new_n658), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n641), .A2(new_n642), .ZN(new_n660));
  NAND2_X1  g459(.A1(new_n595), .A2(new_n660), .ZN(new_n661));
  XOR2_X1   g460(.A(KEYINPUT98), .B(KEYINPUT10), .Z(new_n662));
  NAND4_X1  g461(.A1(new_n592), .A2(new_n641), .A3(new_n642), .A4(new_n594), .ZN(new_n663));
  NAND3_X1  g462(.A1(new_n661), .A2(new_n662), .A3(new_n663), .ZN(new_n664));
  AND3_X1   g463(.A1(new_n592), .A2(KEYINPUT10), .A3(new_n594), .ZN(new_n665));
  NAND3_X1  g464(.A1(new_n665), .A2(new_n640), .A3(new_n643), .ZN(new_n666));
  AOI21_X1  g465(.A(new_n659), .B1(new_n664), .B2(new_n666), .ZN(new_n667));
  AOI21_X1  g466(.A(new_n658), .B1(new_n661), .B2(new_n663), .ZN(new_n668));
  OR2_X1    g467(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  XNOR2_X1  g468(.A(G120gat), .B(G148gat), .ZN(new_n670));
  INV_X1    g469(.A(G204gat), .ZN(new_n671));
  XNOR2_X1  g470(.A(new_n670), .B(new_n671), .ZN(new_n672));
  OR2_X1    g471(.A1(new_n672), .A2(KEYINPUT99), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n672), .A2(KEYINPUT99), .ZN(new_n674));
  AND3_X1   g473(.A1(new_n673), .A2(G176gat), .A3(new_n674), .ZN(new_n675));
  AOI21_X1  g474(.A(G176gat), .B1(new_n673), .B2(new_n674), .ZN(new_n676));
  NOR2_X1   g475(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  INV_X1    g476(.A(new_n677), .ZN(new_n678));
  XNOR2_X1  g477(.A(new_n669), .B(new_n678), .ZN(new_n679));
  INV_X1    g478(.A(new_n679), .ZN(new_n680));
  NAND3_X1  g479(.A1(new_n615), .A2(new_n657), .A3(new_n680), .ZN(new_n681));
  INV_X1    g480(.A(KEYINPUT100), .ZN(new_n682));
  XNOR2_X1  g481(.A(new_n681), .B(new_n682), .ZN(new_n683));
  INV_X1    g482(.A(new_n683), .ZN(new_n684));
  NAND2_X1  g483(.A1(new_n571), .A2(new_n684), .ZN(new_n685));
  NAND2_X1  g484(.A1(new_n469), .A2(new_n471), .ZN(new_n686));
  NOR2_X1   g485(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  XNOR2_X1  g486(.A(new_n687), .B(new_n215), .ZN(G1324gat));
  INV_X1    g487(.A(new_n685), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n689), .A2(new_n390), .ZN(new_n690));
  AND2_X1   g489(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n691));
  NOR2_X1   g490(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n692));
  NOR3_X1   g491(.A1(new_n690), .A2(new_n691), .A3(new_n692), .ZN(new_n693));
  INV_X1    g492(.A(new_n693), .ZN(new_n694));
  INV_X1    g493(.A(KEYINPUT42), .ZN(new_n695));
  AOI22_X1  g494(.A1(new_n694), .A2(new_n695), .B1(G8gat), .B2(new_n690), .ZN(new_n696));
  INV_X1    g495(.A(KEYINPUT101), .ZN(new_n697));
  OAI21_X1  g496(.A(new_n697), .B1(new_n694), .B2(new_n695), .ZN(new_n698));
  NAND3_X1  g497(.A1(new_n693), .A2(KEYINPUT101), .A3(KEYINPUT42), .ZN(new_n699));
  NAND3_X1  g498(.A1(new_n696), .A2(new_n698), .A3(new_n699), .ZN(G1325gat));
  AOI21_X1  g499(.A(G15gat), .B1(new_n689), .B2(new_n500), .ZN(new_n701));
  NAND2_X1  g500(.A1(new_n568), .A2(KEYINPUT102), .ZN(new_n702));
  INV_X1    g501(.A(KEYINPUT102), .ZN(new_n703));
  OAI21_X1  g502(.A(new_n703), .B1(new_n565), .B2(new_n567), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n702), .A2(new_n704), .ZN(new_n705));
  NAND2_X1  g504(.A1(new_n705), .A2(G15gat), .ZN(new_n706));
  XOR2_X1   g505(.A(new_n706), .B(KEYINPUT103), .Z(new_n707));
  AOI21_X1  g506(.A(new_n701), .B1(new_n707), .B2(new_n689), .ZN(G1326gat));
  NOR2_X1   g507(.A1(new_n685), .A2(new_n523), .ZN(new_n709));
  XOR2_X1   g508(.A(KEYINPUT43), .B(G22gat), .Z(new_n710));
  XNOR2_X1  g509(.A(new_n710), .B(KEYINPUT104), .ZN(new_n711));
  XNOR2_X1  g510(.A(new_n709), .B(new_n711), .ZN(G1327gat));
  AOI21_X1  g511(.A(new_n657), .B1(new_n531), .B2(new_n570), .ZN(new_n713));
  INV_X1    g512(.A(new_n615), .ZN(new_n714));
  NAND2_X1  g513(.A1(new_n714), .A2(new_n680), .ZN(new_n715));
  NOR2_X1   g514(.A1(new_n715), .A2(new_n289), .ZN(new_n716));
  AND2_X1   g515(.A1(new_n713), .A2(new_n716), .ZN(new_n717));
  INV_X1    g516(.A(new_n686), .ZN(new_n718));
  INV_X1    g517(.A(new_n230), .ZN(new_n719));
  NAND3_X1  g518(.A1(new_n717), .A2(new_n718), .A3(new_n719), .ZN(new_n720));
  XNOR2_X1  g519(.A(new_n720), .B(KEYINPUT45), .ZN(new_n721));
  NAND2_X1  g520(.A1(new_n531), .A2(new_n570), .ZN(new_n722));
  INV_X1    g521(.A(new_n657), .ZN(new_n723));
  INV_X1    g522(.A(KEYINPUT44), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n724), .A2(KEYINPUT106), .ZN(new_n725));
  NOR2_X1   g524(.A1(new_n724), .A2(KEYINPUT106), .ZN(new_n726));
  INV_X1    g525(.A(new_n726), .ZN(new_n727));
  AOI22_X1  g526(.A1(new_n722), .A2(new_n723), .B1(new_n725), .B2(new_n727), .ZN(new_n728));
  AOI211_X1 g527(.A(new_n657), .B(new_n726), .C1(new_n531), .C2(new_n570), .ZN(new_n729));
  OR2_X1    g528(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  NAND3_X1  g529(.A1(new_n286), .A2(KEYINPUT105), .A3(new_n287), .ZN(new_n731));
  INV_X1    g530(.A(new_n731), .ZN(new_n732));
  AOI21_X1  g531(.A(KEYINPUT105), .B1(new_n286), .B2(new_n287), .ZN(new_n733));
  NOR2_X1   g532(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  NOR2_X1   g533(.A1(new_n715), .A2(new_n734), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n730), .A2(new_n735), .ZN(new_n736));
  OAI21_X1  g535(.A(new_n230), .B1(new_n736), .B2(new_n686), .ZN(new_n737));
  NAND2_X1  g536(.A1(new_n721), .A2(new_n737), .ZN(G1328gat));
  NAND2_X1  g537(.A1(new_n717), .A2(new_n390), .ZN(new_n739));
  NOR2_X1   g538(.A1(new_n739), .A2(G36gat), .ZN(new_n740));
  XNOR2_X1  g539(.A(new_n740), .B(KEYINPUT46), .ZN(new_n741));
  INV_X1    g540(.A(new_n390), .ZN(new_n742));
  OAI21_X1  g541(.A(G36gat), .B1(new_n736), .B2(new_n742), .ZN(new_n743));
  NAND2_X1  g542(.A1(new_n741), .A2(new_n743), .ZN(G1329gat));
  OAI21_X1  g543(.A(G43gat), .B1(new_n736), .B2(new_n568), .ZN(new_n745));
  NAND3_X1  g544(.A1(new_n717), .A2(new_n237), .A3(new_n500), .ZN(new_n746));
  NAND2_X1  g545(.A1(new_n746), .A2(KEYINPUT108), .ZN(new_n747));
  INV_X1    g546(.A(KEYINPUT108), .ZN(new_n748));
  NAND4_X1  g547(.A1(new_n717), .A2(new_n748), .A3(new_n237), .A4(new_n500), .ZN(new_n749));
  NAND2_X1  g548(.A1(new_n747), .A2(new_n749), .ZN(new_n750));
  NAND3_X1  g549(.A1(new_n745), .A2(KEYINPUT47), .A3(new_n750), .ZN(new_n751));
  NAND3_X1  g550(.A1(new_n730), .A2(new_n705), .A3(new_n735), .ZN(new_n752));
  AOI22_X1  g551(.A1(new_n752), .A2(G43gat), .B1(new_n747), .B2(new_n749), .ZN(new_n753));
  XOR2_X1   g552(.A(KEYINPUT107), .B(KEYINPUT47), .Z(new_n754));
  OAI21_X1  g553(.A(new_n751), .B1(new_n753), .B2(new_n754), .ZN(G1330gat));
  INV_X1    g554(.A(new_n523), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n717), .A2(new_n756), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n757), .A2(new_n243), .ZN(new_n758));
  INV_X1    g557(.A(new_n243), .ZN(new_n759));
  NAND3_X1  g558(.A1(new_n730), .A2(new_n759), .A3(new_n735), .ZN(new_n760));
  OAI21_X1  g559(.A(new_n758), .B1(new_n760), .B2(new_n523), .ZN(new_n761));
  XNOR2_X1  g560(.A(new_n761), .B(KEYINPUT48), .ZN(G1331gat));
  AOI211_X1 g561(.A(new_n714), .B(new_n723), .C1(new_n531), .C2(new_n570), .ZN(new_n763));
  INV_X1    g562(.A(new_n734), .ZN(new_n764));
  NOR2_X1   g563(.A1(new_n764), .A2(new_n680), .ZN(new_n765));
  NAND2_X1  g564(.A1(new_n763), .A2(new_n765), .ZN(new_n766));
  XNOR2_X1  g565(.A(new_n686), .B(KEYINPUT109), .ZN(new_n767));
  NOR2_X1   g566(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  XNOR2_X1  g567(.A(new_n768), .B(new_n576), .ZN(G1332gat));
  INV_X1    g568(.A(new_n766), .ZN(new_n770));
  AND2_X1   g569(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n771));
  INV_X1    g570(.A(new_n771), .ZN(new_n772));
  NAND3_X1  g571(.A1(new_n770), .A2(new_n390), .A3(new_n772), .ZN(new_n773));
  NAND2_X1  g572(.A1(new_n773), .A2(KEYINPUT110), .ZN(new_n774));
  NOR2_X1   g573(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n775));
  INV_X1    g574(.A(KEYINPUT110), .ZN(new_n776));
  NAND4_X1  g575(.A1(new_n770), .A2(new_n776), .A3(new_n390), .A4(new_n772), .ZN(new_n777));
  AND3_X1   g576(.A1(new_n774), .A2(new_n775), .A3(new_n777), .ZN(new_n778));
  AOI21_X1  g577(.A(new_n775), .B1(new_n774), .B2(new_n777), .ZN(new_n779));
  NOR2_X1   g578(.A1(new_n778), .A2(new_n779), .ZN(G1333gat));
  NAND3_X1  g579(.A1(new_n770), .A2(new_n582), .A3(new_n500), .ZN(new_n781));
  INV_X1    g580(.A(new_n705), .ZN(new_n782));
  OAI21_X1  g581(.A(G71gat), .B1(new_n766), .B2(new_n782), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n781), .A2(new_n783), .ZN(new_n784));
  XOR2_X1   g583(.A(new_n784), .B(KEYINPUT50), .Z(G1334gat));
  NOR2_X1   g584(.A1(new_n766), .A2(new_n523), .ZN(new_n786));
  XNOR2_X1  g585(.A(new_n786), .B(new_n583), .ZN(G1335gat));
  NOR3_X1   g586(.A1(new_n764), .A2(new_n615), .A3(new_n680), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n730), .A2(new_n788), .ZN(new_n789));
  NOR3_X1   g588(.A1(new_n789), .A2(new_n628), .A3(new_n686), .ZN(new_n790));
  NAND4_X1  g589(.A1(new_n722), .A2(new_n714), .A3(new_n723), .A4(new_n734), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n791), .A2(KEYINPUT51), .ZN(new_n792));
  INV_X1    g591(.A(KEYINPUT51), .ZN(new_n793));
  NAND4_X1  g592(.A1(new_n713), .A2(new_n793), .A3(new_n714), .A4(new_n734), .ZN(new_n794));
  AND2_X1   g593(.A1(new_n792), .A2(new_n794), .ZN(new_n795));
  NAND3_X1  g594(.A1(new_n795), .A2(new_n718), .A3(new_n679), .ZN(new_n796));
  AOI21_X1  g595(.A(new_n790), .B1(new_n628), .B2(new_n796), .ZN(G1336gat));
  NAND4_X1  g596(.A1(new_n792), .A2(new_n390), .A3(new_n679), .A4(new_n794), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n798), .A2(new_n373), .ZN(new_n799));
  NAND4_X1  g598(.A1(new_n730), .A2(G92gat), .A3(new_n390), .A4(new_n788), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  INV_X1    g600(.A(KEYINPUT52), .ZN(new_n802));
  XNOR2_X1  g601(.A(new_n801), .B(new_n802), .ZN(G1337gat));
  OAI21_X1  g602(.A(G99gat), .B1(new_n789), .B2(new_n782), .ZN(new_n804));
  NAND3_X1  g603(.A1(new_n795), .A2(new_n489), .A3(new_n679), .ZN(new_n805));
  OAI21_X1  g604(.A(new_n804), .B1(new_n563), .B2(new_n805), .ZN(G1338gat));
  OAI211_X1 g605(.A(new_n756), .B(new_n788), .C1(new_n728), .C2(new_n729), .ZN(new_n807));
  INV_X1    g606(.A(KEYINPUT53), .ZN(new_n808));
  NAND3_X1  g607(.A1(new_n807), .A2(new_n808), .A3(G106gat), .ZN(new_n809));
  NOR2_X1   g608(.A1(new_n523), .A2(G106gat), .ZN(new_n810));
  NAND4_X1  g609(.A1(new_n792), .A2(new_n679), .A3(new_n794), .A4(new_n810), .ZN(new_n811));
  OAI211_X1 g610(.A(new_n809), .B(new_n811), .C1(KEYINPUT112), .C2(new_n808), .ZN(new_n812));
  AND3_X1   g611(.A1(new_n807), .A2(KEYINPUT111), .A3(G106gat), .ZN(new_n813));
  NOR2_X1   g612(.A1(new_n811), .A2(KEYINPUT112), .ZN(new_n814));
  AOI21_X1  g613(.A(KEYINPUT111), .B1(new_n807), .B2(G106gat), .ZN(new_n815));
  NOR3_X1   g614(.A1(new_n813), .A2(new_n814), .A3(new_n815), .ZN(new_n816));
  OAI21_X1  g615(.A(new_n812), .B1(new_n816), .B2(new_n808), .ZN(G1339gat));
  NAND2_X1  g616(.A1(new_n523), .A2(new_n500), .ZN(new_n818));
  NAND3_X1  g617(.A1(new_n664), .A2(new_n666), .A3(new_n659), .ZN(new_n819));
  INV_X1    g618(.A(KEYINPUT113), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n664), .A2(new_n666), .ZN(new_n822));
  NAND2_X1  g621(.A1(new_n822), .A2(new_n658), .ZN(new_n823));
  NAND4_X1  g622(.A1(new_n664), .A2(new_n666), .A3(KEYINPUT113), .A4(new_n659), .ZN(new_n824));
  NAND4_X1  g623(.A1(new_n821), .A2(new_n823), .A3(KEYINPUT54), .A4(new_n824), .ZN(new_n825));
  INV_X1    g624(.A(KEYINPUT54), .ZN(new_n826));
  AOI21_X1  g625(.A(new_n677), .B1(new_n826), .B2(new_n667), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n825), .A2(new_n827), .ZN(new_n828));
  INV_X1    g627(.A(KEYINPUT55), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n828), .A2(new_n829), .ZN(new_n830));
  OR2_X1    g629(.A1(new_n669), .A2(new_n678), .ZN(new_n831));
  NAND3_X1  g630(.A1(new_n825), .A2(new_n827), .A3(KEYINPUT55), .ZN(new_n832));
  NAND3_X1  g631(.A1(new_n830), .A2(new_n831), .A3(new_n832), .ZN(new_n833));
  INV_X1    g632(.A(new_n833), .ZN(new_n834));
  OAI21_X1  g633(.A(new_n834), .B1(new_n732), .B2(new_n733), .ZN(new_n835));
  NOR3_X1   g634(.A1(new_n267), .A2(new_n271), .A3(new_n266), .ZN(new_n836));
  AOI21_X1  g635(.A(new_n202), .B1(new_n275), .B2(new_n251), .ZN(new_n837));
  OAI21_X1  g636(.A(new_n283), .B1(new_n836), .B2(new_n837), .ZN(new_n838));
  AND3_X1   g637(.A1(new_n287), .A2(new_n838), .A3(new_n679), .ZN(new_n839));
  INV_X1    g638(.A(new_n839), .ZN(new_n840));
  AOI21_X1  g639(.A(new_n723), .B1(new_n835), .B2(new_n840), .ZN(new_n841));
  AND2_X1   g640(.A1(new_n287), .A2(new_n838), .ZN(new_n842));
  NAND3_X1  g641(.A1(new_n723), .A2(new_n834), .A3(new_n842), .ZN(new_n843));
  INV_X1    g642(.A(new_n843), .ZN(new_n844));
  OAI21_X1  g643(.A(new_n714), .B1(new_n841), .B2(new_n844), .ZN(new_n845));
  INV_X1    g644(.A(new_n681), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n846), .A2(new_n734), .ZN(new_n847));
  AOI21_X1  g646(.A(new_n818), .B1(new_n845), .B2(new_n847), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n718), .A2(new_n742), .ZN(new_n849));
  INV_X1    g648(.A(new_n849), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n848), .A2(new_n850), .ZN(new_n851));
  OAI21_X1  g650(.A(G113gat), .B1(new_n851), .B2(new_n289), .ZN(new_n852));
  INV_X1    g651(.A(new_n767), .ZN(new_n853));
  NAND3_X1  g652(.A1(new_n848), .A2(new_n742), .A3(new_n853), .ZN(new_n854));
  NAND2_X1  g653(.A1(new_n764), .A2(new_n396), .ZN(new_n855));
  OAI21_X1  g654(.A(new_n852), .B1(new_n854), .B2(new_n855), .ZN(G1340gat));
  INV_X1    g655(.A(new_n854), .ZN(new_n857));
  NAND3_X1  g656(.A1(new_n857), .A2(new_n398), .A3(new_n679), .ZN(new_n858));
  OAI21_X1  g657(.A(G120gat), .B1(new_n851), .B2(new_n680), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n858), .A2(new_n859), .ZN(G1341gat));
  INV_X1    g659(.A(G127gat), .ZN(new_n861));
  NOR3_X1   g660(.A1(new_n851), .A2(new_n861), .A3(new_n714), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n857), .A2(new_n615), .ZN(new_n863));
  AOI21_X1  g662(.A(new_n862), .B1(new_n863), .B2(new_n861), .ZN(G1342gat));
  NAND4_X1  g663(.A1(new_n848), .A2(new_n742), .A3(new_n723), .A4(new_n853), .ZN(new_n865));
  OAI21_X1  g664(.A(KEYINPUT56), .B1(new_n865), .B2(G134gat), .ZN(new_n866));
  INV_X1    g665(.A(KEYINPUT115), .ZN(new_n867));
  XNOR2_X1  g666(.A(new_n866), .B(new_n867), .ZN(new_n868));
  OAI21_X1  g667(.A(G134gat), .B1(new_n851), .B2(new_n657), .ZN(new_n869));
  NOR2_X1   g668(.A1(new_n865), .A2(G134gat), .ZN(new_n870));
  INV_X1    g669(.A(KEYINPUT56), .ZN(new_n871));
  AOI21_X1  g670(.A(KEYINPUT114), .B1(new_n870), .B2(new_n871), .ZN(new_n872));
  AND3_X1   g671(.A1(new_n870), .A2(KEYINPUT114), .A3(new_n871), .ZN(new_n873));
  OAI211_X1 g672(.A(new_n868), .B(new_n869), .C1(new_n872), .C2(new_n873), .ZN(G1343gat));
  INV_X1    g673(.A(KEYINPUT105), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n288), .A2(new_n875), .ZN(new_n876));
  AOI21_X1  g675(.A(new_n833), .B1(new_n876), .B2(new_n731), .ZN(new_n877));
  OAI21_X1  g676(.A(new_n657), .B1(new_n877), .B2(new_n839), .ZN(new_n878));
  AOI21_X1  g677(.A(new_n615), .B1(new_n878), .B2(new_n843), .ZN(new_n879));
  INV_X1    g678(.A(new_n847), .ZN(new_n880));
  OAI21_X1  g679(.A(new_n756), .B1(new_n879), .B2(new_n880), .ZN(new_n881));
  NOR2_X1   g680(.A1(new_n881), .A2(new_n767), .ZN(new_n882));
  NOR2_X1   g681(.A1(new_n705), .A2(new_n390), .ZN(new_n883));
  AND4_X1   g682(.A1(new_n414), .A2(new_n882), .A3(new_n288), .A4(new_n883), .ZN(new_n884));
  NOR2_X1   g683(.A1(new_n884), .A2(KEYINPUT58), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n850), .A2(new_n568), .ZN(new_n886));
  AOI21_X1  g685(.A(new_n833), .B1(new_n286), .B2(new_n287), .ZN(new_n887));
  OAI21_X1  g686(.A(new_n657), .B1(new_n887), .B2(new_n839), .ZN(new_n888));
  AOI21_X1  g687(.A(new_n615), .B1(new_n888), .B2(new_n843), .ZN(new_n889));
  OAI21_X1  g688(.A(new_n847), .B1(new_n889), .B2(KEYINPUT116), .ZN(new_n890));
  INV_X1    g689(.A(KEYINPUT116), .ZN(new_n891));
  AOI211_X1 g690(.A(new_n891), .B(new_n615), .C1(new_n888), .C2(new_n843), .ZN(new_n892));
  OAI21_X1  g691(.A(new_n756), .B1(new_n890), .B2(new_n892), .ZN(new_n893));
  AOI21_X1  g692(.A(new_n886), .B1(new_n893), .B2(KEYINPUT57), .ZN(new_n894));
  INV_X1    g693(.A(KEYINPUT57), .ZN(new_n895));
  OAI211_X1 g694(.A(new_n895), .B(new_n756), .C1(new_n879), .C2(new_n880), .ZN(new_n896));
  NAND2_X1  g695(.A1(new_n894), .A2(new_n896), .ZN(new_n897));
  OAI21_X1  g696(.A(new_n417), .B1(new_n897), .B2(new_n289), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n885), .A2(new_n898), .ZN(new_n899));
  NAND2_X1  g698(.A1(new_n893), .A2(KEYINPUT57), .ZN(new_n900));
  INV_X1    g699(.A(new_n886), .ZN(new_n901));
  AND4_X1   g700(.A1(KEYINPUT117), .A2(new_n900), .A3(new_n896), .A4(new_n901), .ZN(new_n902));
  AOI21_X1  g701(.A(KEYINPUT117), .B1(new_n894), .B2(new_n896), .ZN(new_n903));
  OAI21_X1  g702(.A(new_n764), .B1(new_n902), .B2(new_n903), .ZN(new_n904));
  AOI21_X1  g703(.A(new_n884), .B1(new_n904), .B2(new_n417), .ZN(new_n905));
  INV_X1    g704(.A(KEYINPUT58), .ZN(new_n906));
  OAI21_X1  g705(.A(new_n899), .B1(new_n905), .B2(new_n906), .ZN(G1344gat));
  INV_X1    g706(.A(KEYINPUT59), .ZN(new_n908));
  AND2_X1   g707(.A1(new_n882), .A2(new_n883), .ZN(new_n909));
  AOI211_X1 g708(.A(new_n908), .B(G148gat), .C1(new_n909), .C2(new_n679), .ZN(new_n910));
  NAND2_X1  g709(.A1(new_n881), .A2(KEYINPUT57), .ZN(new_n911));
  NOR2_X1   g710(.A1(new_n683), .A2(new_n288), .ZN(new_n912));
  AND3_X1   g711(.A1(new_n888), .A2(KEYINPUT118), .A3(new_n843), .ZN(new_n913));
  AOI21_X1  g712(.A(KEYINPUT118), .B1(new_n888), .B2(new_n843), .ZN(new_n914));
  NOR3_X1   g713(.A1(new_n913), .A2(new_n914), .A3(new_n615), .ZN(new_n915));
  OAI211_X1 g714(.A(new_n895), .B(new_n756), .C1(new_n912), .C2(new_n915), .ZN(new_n916));
  NAND3_X1  g715(.A1(new_n911), .A2(new_n679), .A3(new_n916), .ZN(new_n917));
  OR3_X1    g716(.A1(new_n917), .A2(new_n908), .A3(new_n886), .ZN(new_n918));
  INV_X1    g717(.A(KEYINPUT117), .ZN(new_n919));
  NAND2_X1  g718(.A1(new_n897), .A2(new_n919), .ZN(new_n920));
  NAND3_X1  g719(.A1(new_n894), .A2(KEYINPUT117), .A3(new_n896), .ZN(new_n921));
  AOI21_X1  g720(.A(new_n680), .B1(new_n920), .B2(new_n921), .ZN(new_n922));
  OAI21_X1  g721(.A(new_n918), .B1(new_n922), .B2(KEYINPUT59), .ZN(new_n923));
  AOI21_X1  g722(.A(new_n910), .B1(new_n923), .B2(G148gat), .ZN(G1345gat));
  AOI21_X1  g723(.A(G155gat), .B1(new_n909), .B2(new_n615), .ZN(new_n925));
  AOI21_X1  g724(.A(new_n714), .B1(new_n920), .B2(new_n921), .ZN(new_n926));
  AOI21_X1  g725(.A(new_n925), .B1(new_n926), .B2(G155gat), .ZN(G1346gat));
  OAI21_X1  g726(.A(new_n723), .B1(new_n902), .B2(new_n903), .ZN(new_n928));
  NAND2_X1  g727(.A1(new_n928), .A2(KEYINPUT119), .ZN(new_n929));
  INV_X1    g728(.A(KEYINPUT119), .ZN(new_n930));
  OAI211_X1 g729(.A(new_n930), .B(new_n723), .C1(new_n902), .C2(new_n903), .ZN(new_n931));
  NAND3_X1  g730(.A1(new_n929), .A2(G162gat), .A3(new_n931), .ZN(new_n932));
  INV_X1    g731(.A(G162gat), .ZN(new_n933));
  NAND3_X1  g732(.A1(new_n909), .A2(new_n933), .A3(new_n723), .ZN(new_n934));
  NAND2_X1  g733(.A1(new_n932), .A2(new_n934), .ZN(G1347gat));
  NAND2_X1  g734(.A1(new_n848), .A2(new_n390), .ZN(new_n936));
  NOR2_X1   g735(.A1(new_n936), .A2(new_n718), .ZN(new_n937));
  NAND3_X1  g736(.A1(new_n937), .A2(new_n343), .A3(new_n764), .ZN(new_n938));
  NOR2_X1   g737(.A1(new_n936), .A2(new_n853), .ZN(new_n939));
  NAND2_X1  g738(.A1(new_n939), .A2(new_n288), .ZN(new_n940));
  AND3_X1   g739(.A1(new_n940), .A2(KEYINPUT120), .A3(G169gat), .ZN(new_n941));
  AOI21_X1  g740(.A(KEYINPUT120), .B1(new_n940), .B2(G169gat), .ZN(new_n942));
  OAI21_X1  g741(.A(new_n938), .B1(new_n941), .B2(new_n942), .ZN(G1348gat));
  AOI21_X1  g742(.A(G176gat), .B1(new_n937), .B2(new_n679), .ZN(new_n944));
  INV_X1    g743(.A(new_n939), .ZN(new_n945));
  NOR2_X1   g744(.A1(new_n945), .A2(new_n680), .ZN(new_n946));
  AOI21_X1  g745(.A(new_n944), .B1(G176gat), .B2(new_n946), .ZN(G1349gat));
  OAI211_X1 g746(.A(new_n937), .B(new_n615), .C1(new_n335), .C2(new_n334), .ZN(new_n948));
  NAND2_X1  g747(.A1(new_n948), .A2(KEYINPUT121), .ZN(new_n949));
  AOI211_X1 g748(.A(new_n317), .B(new_n316), .C1(new_n939), .C2(new_n615), .ZN(new_n950));
  OAI21_X1  g749(.A(KEYINPUT60), .B1(new_n949), .B2(new_n950), .ZN(new_n951));
  NOR2_X1   g750(.A1(new_n316), .A2(new_n317), .ZN(new_n952));
  OAI21_X1  g751(.A(new_n952), .B1(new_n945), .B2(new_n714), .ZN(new_n953));
  INV_X1    g752(.A(KEYINPUT60), .ZN(new_n954));
  NAND4_X1  g753(.A1(new_n953), .A2(KEYINPUT121), .A3(new_n954), .A4(new_n948), .ZN(new_n955));
  NAND2_X1  g754(.A1(new_n951), .A2(new_n955), .ZN(G1350gat));
  INV_X1    g755(.A(KEYINPUT123), .ZN(new_n957));
  INV_X1    g756(.A(KEYINPUT61), .ZN(new_n958));
  NOR2_X1   g757(.A1(new_n957), .A2(new_n958), .ZN(new_n959));
  AOI211_X1 g758(.A(new_n315), .B(new_n959), .C1(new_n939), .C2(new_n723), .ZN(new_n960));
  OAI21_X1  g759(.A(new_n960), .B1(KEYINPUT123), .B2(KEYINPUT61), .ZN(new_n961));
  OAI21_X1  g760(.A(G190gat), .B1(new_n945), .B2(new_n657), .ZN(new_n962));
  NAND3_X1  g761(.A1(new_n962), .A2(new_n957), .A3(new_n958), .ZN(new_n963));
  NOR4_X1   g762(.A1(new_n936), .A2(G190gat), .A3(new_n718), .A4(new_n657), .ZN(new_n964));
  XNOR2_X1  g763(.A(new_n964), .B(KEYINPUT122), .ZN(new_n965));
  NAND3_X1  g764(.A1(new_n961), .A2(new_n963), .A3(new_n965), .ZN(G1351gat));
  NOR3_X1   g765(.A1(new_n705), .A2(new_n742), .A3(new_n853), .ZN(new_n967));
  AOI21_X1  g766(.A(new_n523), .B1(new_n845), .B2(new_n847), .ZN(new_n968));
  OAI211_X1 g767(.A(new_n916), .B(new_n967), .C1(new_n968), .C2(new_n895), .ZN(new_n969));
  OAI21_X1  g768(.A(G197gat), .B1(new_n969), .B2(new_n289), .ZN(new_n970));
  NAND4_X1  g769(.A1(new_n968), .A2(new_n686), .A3(new_n390), .A4(new_n782), .ZN(new_n971));
  OR2_X1    g770(.A1(new_n734), .A2(G197gat), .ZN(new_n972));
  OAI21_X1  g771(.A(new_n970), .B1(new_n971), .B2(new_n972), .ZN(G1352gat));
  NOR3_X1   g772(.A1(new_n971), .A2(G204gat), .A3(new_n680), .ZN(new_n974));
  INV_X1    g773(.A(KEYINPUT62), .ZN(new_n975));
  OR2_X1    g774(.A1(new_n974), .A2(new_n975), .ZN(new_n976));
  INV_X1    g775(.A(new_n967), .ZN(new_n977));
  OAI21_X1  g776(.A(G204gat), .B1(new_n917), .B2(new_n977), .ZN(new_n978));
  NAND2_X1  g777(.A1(new_n974), .A2(new_n975), .ZN(new_n979));
  NAND3_X1  g778(.A1(new_n976), .A2(new_n978), .A3(new_n979), .ZN(G1353gat));
  OAI21_X1  g779(.A(G211gat), .B1(new_n969), .B2(new_n714), .ZN(new_n981));
  INV_X1    g780(.A(KEYINPUT63), .ZN(new_n982));
  NAND2_X1  g781(.A1(new_n981), .A2(new_n982), .ZN(new_n983));
  OAI211_X1 g782(.A(KEYINPUT63), .B(G211gat), .C1(new_n969), .C2(new_n714), .ZN(new_n984));
  NAND3_X1  g783(.A1(new_n983), .A2(KEYINPUT124), .A3(new_n984), .ZN(new_n985));
  OR3_X1    g784(.A1(new_n971), .A2(G211gat), .A3(new_n714), .ZN(new_n986));
  INV_X1    g785(.A(KEYINPUT124), .ZN(new_n987));
  NAND3_X1  g786(.A1(new_n981), .A2(new_n987), .A3(new_n982), .ZN(new_n988));
  NAND3_X1  g787(.A1(new_n985), .A2(new_n986), .A3(new_n988), .ZN(G1354gat));
  NAND2_X1  g788(.A1(new_n969), .A2(KEYINPUT125), .ZN(new_n990));
  NAND2_X1  g789(.A1(new_n723), .A2(G218gat), .ZN(new_n991));
  XNOR2_X1  g790(.A(new_n991), .B(KEYINPUT126), .ZN(new_n992));
  INV_X1    g791(.A(KEYINPUT125), .ZN(new_n993));
  NAND4_X1  g792(.A1(new_n911), .A2(new_n993), .A3(new_n916), .A4(new_n967), .ZN(new_n994));
  NAND3_X1  g793(.A1(new_n990), .A2(new_n992), .A3(new_n994), .ZN(new_n995));
  INV_X1    g794(.A(G218gat), .ZN(new_n996));
  OAI21_X1  g795(.A(new_n996), .B1(new_n971), .B2(new_n657), .ZN(new_n997));
  NAND2_X1  g796(.A1(new_n995), .A2(new_n997), .ZN(new_n998));
  INV_X1    g797(.A(KEYINPUT127), .ZN(new_n999));
  NAND2_X1  g798(.A1(new_n998), .A2(new_n999), .ZN(new_n1000));
  NAND3_X1  g799(.A1(new_n995), .A2(KEYINPUT127), .A3(new_n997), .ZN(new_n1001));
  NAND2_X1  g800(.A1(new_n1000), .A2(new_n1001), .ZN(G1355gat));
endmodule


