

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n339, n340, n341, n342, n343, n344, n345, n346, n347, n348, n349,
         n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360,
         n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371,
         n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382,
         n383, n384, n385, n386, n387, n388, n389, n390, n392, n393, n394,
         n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405,
         n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416,
         n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427,
         n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438,
         n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449,
         n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460,
         n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471,
         n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482,
         n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493,
         n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504,
         n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515,
         n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526,
         n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537,
         n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
         n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559,
         n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570,
         n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581,
         n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592,
         n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603,
         n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614,
         n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625,
         n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636,
         n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647,
         n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658,
         n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669,
         n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680,
         n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691,
         n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702,
         n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713,
         n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724,
         n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735,
         n736, n737;

  OR2_X1 U361 ( .A1(n737), .A2(n685), .ZN(n575) );
  BUF_X1 U362 ( .A(n501), .Z(n518) );
  NOR2_X1 U363 ( .A1(G953), .A2(G237), .ZN(n472) );
  XNOR2_X1 U364 ( .A(n421), .B(KEYINPUT67), .ZN(n626) );
  INV_X1 U365 ( .A(G953), .ZN(n727) );
  NOR2_X1 U366 ( .A1(n547), .A2(n632), .ZN(n540) );
  XNOR2_X2 U367 ( .A(n411), .B(n725), .ZN(n431) );
  INV_X1 U368 ( .A(n611), .ZN(n589) );
  AND2_X1 U369 ( .A1(n526), .A2(n525), .ZN(n359) );
  XNOR2_X1 U370 ( .A(n417), .B(n416), .ZN(n622) );
  BUF_X1 U371 ( .A(n551), .Z(n339) );
  BUF_X1 U372 ( .A(n688), .Z(n716) );
  XNOR2_X2 U373 ( .A(n487), .B(n399), .ZN(n725) );
  XNOR2_X1 U374 ( .A(G119), .B(G113), .ZN(n422) );
  XNOR2_X1 U375 ( .A(KEYINPUT15), .B(G902), .ZN(n590) );
  XNOR2_X1 U376 ( .A(n443), .B(KEYINPUT10), .ZN(n462) );
  INV_X1 U377 ( .A(G146), .ZN(n411) );
  INV_X1 U378 ( .A(G237), .ZN(n447) );
  XOR2_X1 U379 ( .A(KEYINPUT11), .B(G143), .Z(n471) );
  XNOR2_X1 U380 ( .A(n372), .B(G146), .ZN(n443) );
  INV_X1 U381 ( .A(G125), .ZN(n372) );
  XNOR2_X1 U382 ( .A(n363), .B(KEYINPUT17), .ZN(n362) );
  XNOR2_X1 U383 ( .A(KEYINPUT85), .B(KEYINPUT18), .ZN(n363) );
  XNOR2_X1 U384 ( .A(KEYINPUT74), .B(KEYINPUT4), .ZN(n361) );
  NAND2_X1 U385 ( .A1(n369), .A2(n340), .ZN(n364) );
  XNOR2_X1 U386 ( .A(n355), .B(n519), .ZN(n354) );
  NAND2_X1 U387 ( .A1(n518), .A2(n652), .ZN(n355) );
  XNOR2_X1 U388 ( .A(n491), .B(n490), .ZN(n520) );
  XNOR2_X1 U389 ( .A(n374), .B(n437), .ZN(n373) );
  NAND2_X1 U390 ( .A1(G234), .A2(G237), .ZN(n450) );
  XOR2_X1 U391 ( .A(G137), .B(G140), .Z(n412) );
  XNOR2_X1 U392 ( .A(G101), .B(G104), .ZN(n392) );
  NAND2_X1 U393 ( .A1(n611), .A2(n349), .ZN(n386) );
  XNOR2_X1 U394 ( .A(n517), .B(n516), .ZN(n652) );
  NAND2_X1 U395 ( .A1(n627), .A2(n626), .ZN(n515) );
  INV_X1 U396 ( .A(G902), .ZN(n489) );
  AND2_X2 U397 ( .A1(n356), .A2(n587), .ZN(n726) );
  XNOR2_X1 U398 ( .A(n357), .B(n578), .ZN(n356) );
  XNOR2_X1 U399 ( .A(KEYINPUT71), .B(KEYINPUT16), .ZN(n374) );
  INV_X1 U400 ( .A(G110), .ZN(n437) );
  XNOR2_X1 U401 ( .A(n352), .B(KEYINPUT83), .ZN(n551) );
  INV_X1 U402 ( .A(n560), .ZN(n371) );
  NOR2_X1 U403 ( .A1(n717), .A2(G902), .ZN(n417) );
  OR2_X1 U404 ( .A1(n689), .A2(G902), .ZN(n433) );
  AND2_X1 U405 ( .A1(n626), .A2(n542), .ZN(n557) );
  XNOR2_X1 U406 ( .A(n484), .B(n483), .ZN(n485) );
  XNOR2_X1 U407 ( .A(n476), .B(n475), .ZN(n602) );
  XNOR2_X1 U408 ( .A(n474), .B(n473), .ZN(n475) );
  XNOR2_X1 U409 ( .A(n362), .B(n361), .ZN(n445) );
  NOR2_X1 U410 ( .A1(n727), .A2(G952), .ZN(n722) );
  NOR2_X1 U411 ( .A1(n570), .A2(n654), .ZN(n571) );
  NAND2_X1 U412 ( .A1(n341), .A2(n365), .ZN(n574) );
  NAND2_X1 U413 ( .A1(n354), .A2(n522), .ZN(n353) );
  XNOR2_X1 U414 ( .A(n460), .B(n459), .ZN(n709) );
  XNOR2_X1 U415 ( .A(n493), .B(KEYINPUT102), .ZN(n707) );
  XOR2_X1 U416 ( .A(n559), .B(KEYINPUT30), .Z(n340) );
  AND2_X1 U417 ( .A1(n364), .A2(n368), .ZN(n341) );
  AND2_X1 U418 ( .A1(G217), .A2(n418), .ZN(n342) );
  AND2_X1 U419 ( .A1(G227), .A2(n727), .ZN(n343) );
  XOR2_X1 U420 ( .A(KEYINPUT24), .B(KEYINPUT93), .Z(n344) );
  XNOR2_X1 U421 ( .A(n551), .B(KEYINPUT19), .ZN(n544) );
  AND2_X1 U422 ( .A1(n340), .A2(n371), .ZN(n345) );
  AND2_X1 U423 ( .A1(n371), .A2(n638), .ZN(n346) );
  AND2_X1 U424 ( .A1(n449), .A2(G210), .ZN(n347) );
  AND2_X1 U425 ( .A1(n557), .A2(n632), .ZN(n348) );
  INV_X1 U426 ( .A(KEYINPUT39), .ZN(n370) );
  INV_X1 U427 ( .A(n707), .ZN(n368) );
  AND2_X1 U428 ( .A1(n591), .A2(KEYINPUT2), .ZN(n349) );
  AND2_X1 U429 ( .A1(n387), .A2(KEYINPUT64), .ZN(n350) );
  INV_X1 U430 ( .A(n388), .ZN(n387) );
  XNOR2_X1 U431 ( .A(KEYINPUT59), .B(KEYINPUT87), .ZN(n351) );
  NAND2_X1 U432 ( .A1(n561), .A2(n390), .ZN(n352) );
  XNOR2_X2 U433 ( .A(n448), .B(n347), .ZN(n561) );
  XNOR2_X2 U434 ( .A(n353), .B(n523), .ZN(n687) );
  NAND2_X2 U435 ( .A1(n617), .A2(n726), .ZN(n611) );
  AND2_X1 U436 ( .A1(n576), .A2(n577), .ZN(n357) );
  XNOR2_X2 U437 ( .A(n358), .B(KEYINPUT45), .ZN(n617) );
  NAND2_X1 U438 ( .A1(n360), .A2(n359), .ZN(n358) );
  NAND2_X1 U439 ( .A1(n531), .A2(n532), .ZN(n360) );
  NAND2_X1 U440 ( .A1(n380), .A2(n378), .ZN(n377) );
  XNOR2_X2 U441 ( .A(n441), .B(n398), .ZN(n487) );
  INV_X2 U442 ( .A(G104), .ZN(n376) );
  XNOR2_X2 U443 ( .A(n461), .B(KEYINPUT96), .ZN(n697) );
  NOR2_X1 U444 ( .A1(n589), .A2(KEYINPUT64), .ZN(n385) );
  XNOR2_X1 U445 ( .A(n599), .B(n598), .ZN(n601) );
  XOR2_X2 U446 ( .A(G116), .B(G107), .Z(n482) );
  NAND2_X1 U447 ( .A1(n365), .A2(n364), .ZN(n579) );
  NAND2_X1 U448 ( .A1(n366), .A2(n370), .ZN(n365) );
  NAND2_X1 U449 ( .A1(n346), .A2(n340), .ZN(n366) );
  NOR2_X1 U450 ( .A1(n560), .A2(n367), .ZN(n369) );
  NAND2_X1 U451 ( .A1(n638), .A2(KEYINPUT39), .ZN(n367) );
  XNOR2_X1 U452 ( .A(n375), .B(n373), .ZN(n439) );
  XNOR2_X1 U453 ( .A(n482), .B(n463), .ZN(n375) );
  XNOR2_X2 U454 ( .A(n376), .B(G122), .ZN(n463) );
  NAND2_X2 U455 ( .A1(n382), .A2(n377), .ZN(n688) );
  NAND2_X1 U456 ( .A1(n386), .A2(n379), .ZN(n378) );
  NAND2_X1 U457 ( .A1(n388), .A2(n592), .ZN(n379) );
  NAND2_X1 U458 ( .A1(n381), .A2(n592), .ZN(n380) );
  INV_X1 U459 ( .A(n386), .ZN(n381) );
  AND2_X2 U460 ( .A1(n384), .A2(n383), .ZN(n382) );
  NAND2_X1 U461 ( .A1(n589), .A2(n350), .ZN(n383) );
  NAND2_X1 U462 ( .A1(n385), .A2(n386), .ZN(n384) );
  NAND2_X1 U463 ( .A1(n589), .A2(n588), .ZN(n615) );
  NAND2_X1 U464 ( .A1(n591), .A2(n588), .ZN(n388) );
  OR2_X1 U465 ( .A1(n645), .A2(n644), .ZN(n389) );
  NAND2_X1 U466 ( .A1(n449), .A2(G214), .ZN(n390) );
  AND2_X1 U467 ( .A1(n601), .A2(n600), .ZN(G54) );
  INV_X1 U468 ( .A(KEYINPUT23), .ZN(n405) );
  XNOR2_X1 U469 ( .A(n406), .B(n405), .ZN(n407) );
  INV_X1 U470 ( .A(KEYINPUT2), .ZN(n588) );
  INV_X1 U471 ( .A(KEYINPUT7), .ZN(n483) );
  XNOR2_X1 U472 ( .A(KEYINPUT108), .B(KEYINPUT28), .ZN(n539) );
  NOR2_X1 U473 ( .A1(n547), .A2(n707), .ZN(n550) );
  XNOR2_X1 U474 ( .A(n540), .B(n539), .ZN(n541) );
  XNOR2_X1 U475 ( .A(n486), .B(n485), .ZN(n488) );
  XNOR2_X1 U476 ( .A(n717), .B(n718), .ZN(n719) );
  INV_X1 U477 ( .A(n607), .ZN(n608) );
  XNOR2_X1 U478 ( .A(n720), .B(n719), .ZN(n721) );
  NOR2_X1 U479 ( .A1(n610), .A2(n722), .ZN(G63) );
  XNOR2_X1 U480 ( .A(KEYINPUT73), .B(KEYINPUT92), .ZN(n397) );
  XOR2_X1 U481 ( .A(G107), .B(G110), .Z(n393) );
  XNOR2_X1 U482 ( .A(n393), .B(n392), .ZN(n395) );
  XNOR2_X1 U483 ( .A(n412), .B(n343), .ZN(n394) );
  XNOR2_X1 U484 ( .A(n395), .B(n394), .ZN(n396) );
  XNOR2_X1 U485 ( .A(n397), .B(n396), .ZN(n400) );
  XNOR2_X2 U486 ( .A(G143), .B(G128), .ZN(n441) );
  INV_X1 U487 ( .A(G134), .ZN(n398) );
  XNOR2_X1 U488 ( .A(KEYINPUT4), .B(G131), .ZN(n399) );
  XNOR2_X1 U489 ( .A(n400), .B(n431), .ZN(n593) );
  NAND2_X1 U490 ( .A1(n593), .A2(n489), .ZN(n402) );
  XOR2_X1 U491 ( .A(KEYINPUT69), .B(G469), .Z(n401) );
  XNOR2_X2 U492 ( .A(n402), .B(n401), .ZN(n542) );
  XNOR2_X2 U493 ( .A(n542), .B(KEYINPUT1), .ZN(n627) );
  NAND2_X1 U494 ( .A1(G234), .A2(n727), .ZN(n403) );
  XOR2_X1 U495 ( .A(n403), .B(KEYINPUT8), .Z(n479) );
  NAND2_X1 U496 ( .A1(n479), .A2(G221), .ZN(n410) );
  XNOR2_X1 U497 ( .A(G128), .B(KEYINPUT77), .ZN(n404) );
  XNOR2_X1 U498 ( .A(n344), .B(n404), .ZN(n408) );
  XNOR2_X1 U499 ( .A(G119), .B(G110), .ZN(n406) );
  XNOR2_X1 U500 ( .A(n408), .B(n407), .ZN(n409) );
  XNOR2_X1 U501 ( .A(n410), .B(n409), .ZN(n413) );
  XNOR2_X1 U502 ( .A(n412), .B(n462), .ZN(n723) );
  XNOR2_X1 U503 ( .A(n413), .B(n723), .ZN(n717) );
  XOR2_X1 U504 ( .A(KEYINPUT25), .B(KEYINPUT72), .Z(n415) );
  NAND2_X1 U505 ( .A1(G234), .A2(n590), .ZN(n414) );
  XNOR2_X1 U506 ( .A(KEYINPUT20), .B(n414), .ZN(n418) );
  XNOR2_X1 U507 ( .A(n415), .B(n342), .ZN(n416) );
  AND2_X1 U508 ( .A1(n418), .A2(G221), .ZN(n420) );
  XNOR2_X1 U509 ( .A(KEYINPUT94), .B(KEYINPUT21), .ZN(n419) );
  XNOR2_X1 U510 ( .A(n420), .B(n419), .ZN(n623) );
  NAND2_X1 U511 ( .A1(n622), .A2(n623), .ZN(n421) );
  INV_X1 U512 ( .A(n515), .ZN(n434) );
  XNOR2_X1 U513 ( .A(n422), .B(KEYINPUT3), .ZN(n424) );
  XNOR2_X1 U514 ( .A(G101), .B(KEYINPUT89), .ZN(n423) );
  XNOR2_X1 U515 ( .A(n424), .B(n423), .ZN(n438) );
  NAND2_X1 U516 ( .A1(n472), .A2(G210), .ZN(n426) );
  XNOR2_X1 U517 ( .A(G137), .B(G116), .ZN(n425) );
  XNOR2_X1 U518 ( .A(n426), .B(n425), .ZN(n428) );
  XNOR2_X1 U519 ( .A(KEYINPUT95), .B(KEYINPUT5), .ZN(n427) );
  XNOR2_X1 U520 ( .A(n428), .B(n427), .ZN(n429) );
  XNOR2_X1 U521 ( .A(n438), .B(n429), .ZN(n430) );
  XNOR2_X1 U522 ( .A(n431), .B(n430), .ZN(n689) );
  XNOR2_X1 U523 ( .A(G472), .B(KEYINPUT70), .ZN(n432) );
  XNOR2_X2 U524 ( .A(n433), .B(n432), .ZN(n558) );
  NAND2_X1 U525 ( .A1(n434), .A2(n558), .ZN(n436) );
  INV_X1 U526 ( .A(KEYINPUT97), .ZN(n435) );
  XNOR2_X1 U527 ( .A(n436), .B(n435), .ZN(n635) );
  INV_X1 U528 ( .A(n635), .ZN(n458) );
  XNOR2_X1 U529 ( .A(n439), .B(n438), .ZN(n679) );
  NAND2_X1 U530 ( .A1(G224), .A2(n727), .ZN(n440) );
  XNOR2_X1 U531 ( .A(n441), .B(n440), .ZN(n442) );
  XNOR2_X1 U532 ( .A(n443), .B(n442), .ZN(n444) );
  XNOR2_X1 U533 ( .A(n445), .B(n444), .ZN(n446) );
  XNOR2_X1 U534 ( .A(n679), .B(n446), .ZN(n666) );
  NAND2_X1 U535 ( .A1(n666), .A2(n590), .ZN(n448) );
  NAND2_X1 U536 ( .A1(n489), .A2(n447), .ZN(n449) );
  XNOR2_X1 U537 ( .A(n450), .B(KEYINPUT14), .ZN(n453) );
  NAND2_X1 U538 ( .A1(G952), .A2(n453), .ZN(n651) );
  NOR2_X1 U539 ( .A1(G953), .A2(n651), .ZN(n452) );
  INV_X1 U540 ( .A(KEYINPUT90), .ZN(n451) );
  XNOR2_X1 U541 ( .A(n452), .B(n451), .ZN(n536) );
  NAND2_X1 U542 ( .A1(G902), .A2(n453), .ZN(n533) );
  XNOR2_X1 U543 ( .A(G898), .B(KEYINPUT91), .ZN(n675) );
  NAND2_X1 U544 ( .A1(G953), .A2(n675), .ZN(n680) );
  OR2_X1 U545 ( .A1(n533), .A2(n680), .ZN(n454) );
  AND2_X1 U546 ( .A1(n536), .A2(n454), .ZN(n455) );
  OR2_X2 U547 ( .A1(n544), .A2(n455), .ZN(n457) );
  XNOR2_X1 U548 ( .A(KEYINPUT65), .B(KEYINPUT0), .ZN(n456) );
  XNOR2_X2 U549 ( .A(n457), .B(n456), .ZN(n501) );
  NAND2_X1 U550 ( .A1(n458), .A2(n501), .ZN(n460) );
  INV_X1 U551 ( .A(KEYINPUT31), .ZN(n459) );
  NAND2_X1 U552 ( .A1(n518), .A2(n348), .ZN(n461) );
  NAND2_X1 U553 ( .A1(n709), .A2(n697), .ZN(n494) );
  INV_X1 U554 ( .A(n462), .ZN(n469) );
  XNOR2_X1 U555 ( .A(n463), .B(KEYINPUT100), .ZN(n467) );
  XOR2_X1 U556 ( .A(KEYINPUT12), .B(KEYINPUT98), .Z(n465) );
  XNOR2_X1 U557 ( .A(G140), .B(KEYINPUT99), .ZN(n464) );
  XNOR2_X1 U558 ( .A(n465), .B(n464), .ZN(n466) );
  XNOR2_X1 U559 ( .A(n467), .B(n466), .ZN(n468) );
  XOR2_X1 U560 ( .A(n469), .B(n468), .Z(n476) );
  XNOR2_X1 U561 ( .A(G113), .B(G131), .ZN(n470) );
  XNOR2_X1 U562 ( .A(n471), .B(n470), .ZN(n474) );
  NAND2_X1 U563 ( .A1(G214), .A2(n472), .ZN(n473) );
  NOR2_X1 U564 ( .A1(G902), .A2(n602), .ZN(n478) );
  XNOR2_X1 U565 ( .A(KEYINPUT13), .B(G475), .ZN(n477) );
  XNOR2_X1 U566 ( .A(n478), .B(n477), .ZN(n496) );
  NAND2_X1 U567 ( .A1(G217), .A2(n479), .ZN(n481) );
  XOR2_X1 U568 ( .A(KEYINPUT9), .B(KEYINPUT101), .Z(n480) );
  XNOR2_X1 U569 ( .A(n481), .B(n480), .ZN(n486) );
  XNOR2_X1 U570 ( .A(G122), .B(n482), .ZN(n484) );
  XNOR2_X1 U571 ( .A(n488), .B(n487), .ZN(n607) );
  NAND2_X1 U572 ( .A1(n607), .A2(n489), .ZN(n491) );
  INV_X1 U573 ( .A(G478), .ZN(n490) );
  NOR2_X1 U574 ( .A1(n496), .A2(n520), .ZN(n492) );
  XOR2_X1 U575 ( .A(KEYINPUT103), .B(n492), .Z(n702) );
  INV_X1 U576 ( .A(n702), .ZN(n710) );
  NAND2_X1 U577 ( .A1(n520), .A2(n496), .ZN(n493) );
  NAND2_X1 U578 ( .A1(n710), .A2(n707), .ZN(n641) );
  NAND2_X1 U579 ( .A1(n494), .A2(n641), .ZN(n495) );
  XNOR2_X1 U580 ( .A(n495), .B(KEYINPUT104), .ZN(n507) );
  INV_X1 U581 ( .A(n496), .ZN(n521) );
  NAND2_X1 U582 ( .A1(n521), .A2(n520), .ZN(n498) );
  INV_X1 U583 ( .A(KEYINPUT105), .ZN(n497) );
  XNOR2_X1 U584 ( .A(n498), .B(n497), .ZN(n640) );
  INV_X1 U585 ( .A(n623), .ZN(n499) );
  NOR2_X1 U586 ( .A1(n640), .A2(n499), .ZN(n500) );
  NAND2_X1 U587 ( .A1(n501), .A2(n500), .ZN(n503) );
  INV_X1 U588 ( .A(KEYINPUT22), .ZN(n502) );
  XNOR2_X2 U589 ( .A(n503), .B(n502), .ZN(n510) );
  XNOR2_X1 U590 ( .A(n558), .B(KEYINPUT6), .ZN(n548) );
  NAND2_X1 U591 ( .A1(n510), .A2(n548), .ZN(n504) );
  XNOR2_X1 U592 ( .A(n504), .B(KEYINPUT81), .ZN(n506) );
  INV_X1 U593 ( .A(n622), .ZN(n538) );
  NOR2_X1 U594 ( .A1(n627), .A2(n538), .ZN(n505) );
  NAND2_X1 U595 ( .A1(n506), .A2(n505), .ZN(n695) );
  AND2_X1 U596 ( .A1(n507), .A2(n695), .ZN(n526) );
  XNOR2_X1 U597 ( .A(n627), .B(KEYINPUT86), .ZN(n554) );
  AND2_X1 U598 ( .A1(n554), .A2(n538), .ZN(n508) );
  AND2_X1 U599 ( .A1(n548), .A2(n508), .ZN(n509) );
  NAND2_X1 U600 ( .A1(n510), .A2(n509), .ZN(n511) );
  XNOR2_X2 U601 ( .A(n511), .B(KEYINPUT32), .ZN(n686) );
  OR2_X1 U602 ( .A1(n622), .A2(n558), .ZN(n512) );
  NOR2_X1 U603 ( .A1(n627), .A2(n512), .ZN(n513) );
  AND2_X1 U604 ( .A1(n510), .A2(n513), .ZN(n701) );
  INV_X1 U605 ( .A(n701), .ZN(n514) );
  AND2_X2 U606 ( .A1(n686), .A2(n514), .ZN(n527) );
  OR2_X1 U607 ( .A1(n515), .A2(n548), .ZN(n517) );
  XNOR2_X1 U608 ( .A(KEYINPUT106), .B(KEYINPUT33), .ZN(n516) );
  INV_X1 U609 ( .A(KEYINPUT34), .ZN(n519) );
  OR2_X1 U610 ( .A1(n521), .A2(n520), .ZN(n562) );
  INV_X1 U611 ( .A(n562), .ZN(n522) );
  XNOR2_X1 U612 ( .A(KEYINPUT79), .B(KEYINPUT35), .ZN(n523) );
  NAND2_X1 U613 ( .A1(n527), .A2(n687), .ZN(n524) );
  NAND2_X1 U614 ( .A1(n524), .A2(KEYINPUT44), .ZN(n525) );
  XNOR2_X1 U615 ( .A(n527), .B(KEYINPUT82), .ZN(n532) );
  INV_X1 U616 ( .A(KEYINPUT44), .ZN(n528) );
  NAND2_X1 U617 ( .A1(n687), .A2(n528), .ZN(n530) );
  INV_X1 U618 ( .A(KEYINPUT66), .ZN(n529) );
  XNOR2_X1 U619 ( .A(n530), .B(n529), .ZN(n531) );
  NOR2_X1 U620 ( .A1(G900), .A2(n533), .ZN(n534) );
  NAND2_X1 U621 ( .A1(n534), .A2(G953), .ZN(n535) );
  NAND2_X1 U622 ( .A1(n536), .A2(n535), .ZN(n556) );
  AND2_X1 U623 ( .A1(n623), .A2(n556), .ZN(n537) );
  NAND2_X1 U624 ( .A1(n538), .A2(n537), .ZN(n547) );
  INV_X1 U625 ( .A(n558), .ZN(n632) );
  NAND2_X1 U626 ( .A1(n542), .A2(n541), .ZN(n543) );
  XOR2_X1 U627 ( .A(KEYINPUT109), .B(n543), .Z(n570) );
  NOR2_X1 U628 ( .A1(n570), .A2(n544), .ZN(n705) );
  NAND2_X1 U629 ( .A1(n705), .A2(n641), .ZN(n546) );
  INV_X1 U630 ( .A(KEYINPUT47), .ZN(n545) );
  XNOR2_X1 U631 ( .A(n546), .B(n545), .ZN(n567) );
  INV_X1 U632 ( .A(n548), .ZN(n549) );
  NAND2_X1 U633 ( .A1(n550), .A2(n549), .ZN(n581) );
  INV_X1 U634 ( .A(n339), .ZN(n552) );
  NOR2_X1 U635 ( .A1(n581), .A2(n552), .ZN(n553) );
  XNOR2_X1 U636 ( .A(n553), .B(KEYINPUT36), .ZN(n555) );
  NAND2_X1 U637 ( .A1(n555), .A2(n554), .ZN(n713) );
  XNOR2_X1 U638 ( .A(n713), .B(KEYINPUT80), .ZN(n565) );
  NAND2_X1 U639 ( .A1(n557), .A2(n556), .ZN(n560) );
  NAND2_X1 U640 ( .A1(n558), .A2(n390), .ZN(n559) );
  INV_X1 U641 ( .A(n561), .ZN(n586) );
  NOR2_X1 U642 ( .A1(n562), .A2(n586), .ZN(n563) );
  NAND2_X1 U643 ( .A1(n345), .A2(n563), .ZN(n671) );
  XNOR2_X1 U644 ( .A(n671), .B(KEYINPUT76), .ZN(n564) );
  AND2_X1 U645 ( .A1(n565), .A2(n564), .ZN(n566) );
  AND2_X1 U646 ( .A1(n567), .A2(n566), .ZN(n577) );
  INV_X1 U647 ( .A(KEYINPUT38), .ZN(n568) );
  XNOR2_X1 U648 ( .A(n586), .B(n568), .ZN(n572) );
  INV_X1 U649 ( .A(n572), .ZN(n638) );
  NAND2_X1 U650 ( .A1(n638), .A2(n390), .ZN(n642) );
  NOR2_X1 U651 ( .A1(n642), .A2(n640), .ZN(n569) );
  XNOR2_X1 U652 ( .A(n569), .B(KEYINPUT41), .ZN(n654) );
  XNOR2_X1 U653 ( .A(n571), .B(KEYINPUT42), .ZN(n737) );
  INV_X1 U654 ( .A(KEYINPUT40), .ZN(n573) );
  XNOR2_X1 U655 ( .A(n574), .B(n573), .ZN(n685) );
  XOR2_X1 U656 ( .A(n575), .B(KEYINPUT46), .Z(n576) );
  XNOR2_X1 U657 ( .A(KEYINPUT68), .B(KEYINPUT48), .ZN(n578) );
  OR2_X1 U658 ( .A1(n579), .A2(n710), .ZN(n580) );
  XNOR2_X1 U659 ( .A(n580), .B(KEYINPUT110), .ZN(n735) );
  XOR2_X1 U660 ( .A(KEYINPUT43), .B(KEYINPUT107), .Z(n584) );
  NOR2_X1 U661 ( .A1(n627), .A2(n581), .ZN(n582) );
  NAND2_X1 U662 ( .A1(n390), .A2(n582), .ZN(n583) );
  XNOR2_X1 U663 ( .A(n584), .B(n583), .ZN(n585) );
  NAND2_X1 U664 ( .A1(n586), .A2(n585), .ZN(n714) );
  AND2_X1 U665 ( .A1(n735), .A2(n714), .ZN(n587) );
  INV_X1 U666 ( .A(n590), .ZN(n591) );
  INV_X1 U667 ( .A(KEYINPUT64), .ZN(n592) );
  NAND2_X1 U668 ( .A1(n716), .A2(G469), .ZN(n599) );
  XNOR2_X1 U669 ( .A(KEYINPUT58), .B(KEYINPUT118), .ZN(n595) );
  XOR2_X1 U670 ( .A(KEYINPUT119), .B(n593), .Z(n594) );
  XNOR2_X1 U671 ( .A(n595), .B(n594), .ZN(n597) );
  XOR2_X1 U672 ( .A(KEYINPUT120), .B(KEYINPUT57), .Z(n596) );
  XNOR2_X1 U673 ( .A(n597), .B(n596), .ZN(n598) );
  INV_X1 U674 ( .A(n722), .ZN(n600) );
  NAND2_X1 U675 ( .A1(n688), .A2(G475), .ZN(n604) );
  XNOR2_X1 U676 ( .A(n602), .B(n351), .ZN(n603) );
  XNOR2_X1 U677 ( .A(n604), .B(n603), .ZN(n605) );
  NOR2_X2 U678 ( .A1(n605), .A2(n722), .ZN(n606) );
  XNOR2_X1 U679 ( .A(n606), .B(KEYINPUT60), .ZN(G60) );
  NAND2_X1 U680 ( .A1(n716), .A2(G478), .ZN(n609) );
  XNOR2_X1 U681 ( .A(n609), .B(n608), .ZN(n610) );
  NAND2_X1 U682 ( .A1(n611), .A2(KEYINPUT78), .ZN(n612) );
  NAND2_X1 U683 ( .A1(n612), .A2(KEYINPUT2), .ZN(n614) );
  INV_X1 U684 ( .A(KEYINPUT78), .ZN(n618) );
  OR2_X1 U685 ( .A1(n618), .A2(KEYINPUT2), .ZN(n613) );
  NAND2_X1 U686 ( .A1(n614), .A2(n613), .ZN(n616) );
  NAND2_X1 U687 ( .A1(n616), .A2(n615), .ZN(n621) );
  INV_X1 U688 ( .A(n617), .ZN(n672) );
  NAND2_X1 U689 ( .A1(n672), .A2(n726), .ZN(n619) );
  NAND2_X1 U690 ( .A1(n619), .A2(n618), .ZN(n620) );
  NAND2_X1 U691 ( .A1(n621), .A2(n620), .ZN(n658) );
  XNOR2_X1 U692 ( .A(KEYINPUT113), .B(KEYINPUT49), .ZN(n625) );
  NOR2_X1 U693 ( .A1(n623), .A2(n622), .ZN(n624) );
  XNOR2_X1 U694 ( .A(n625), .B(n624), .ZN(n631) );
  XOR2_X1 U695 ( .A(KEYINPUT50), .B(KEYINPUT114), .Z(n629) );
  OR2_X1 U696 ( .A1(n627), .A2(n626), .ZN(n628) );
  XNOR2_X1 U697 ( .A(n629), .B(n628), .ZN(n630) );
  NOR2_X1 U698 ( .A1(n631), .A2(n630), .ZN(n633) );
  NAND2_X1 U699 ( .A1(n633), .A2(n632), .ZN(n634) );
  NAND2_X1 U700 ( .A1(n635), .A2(n634), .ZN(n636) );
  XNOR2_X1 U701 ( .A(KEYINPUT51), .B(n636), .ZN(n637) );
  NOR2_X1 U702 ( .A1(n637), .A2(n654), .ZN(n647) );
  NOR2_X1 U703 ( .A1(n638), .A2(n390), .ZN(n639) );
  NOR2_X1 U704 ( .A1(n640), .A2(n639), .ZN(n645) );
  INV_X1 U705 ( .A(n641), .ZN(n643) );
  NOR2_X1 U706 ( .A1(n643), .A2(n642), .ZN(n644) );
  AND2_X1 U707 ( .A1(n652), .A2(n389), .ZN(n646) );
  NOR2_X1 U708 ( .A1(n647), .A2(n646), .ZN(n648) );
  XOR2_X1 U709 ( .A(n648), .B(KEYINPUT52), .Z(n649) );
  XNOR2_X1 U710 ( .A(KEYINPUT115), .B(n649), .ZN(n650) );
  NOR2_X1 U711 ( .A1(n651), .A2(n650), .ZN(n656) );
  INV_X1 U712 ( .A(n652), .ZN(n653) );
  NOR2_X1 U713 ( .A1(n654), .A2(n653), .ZN(n655) );
  NOR2_X1 U714 ( .A1(n656), .A2(n655), .ZN(n657) );
  NAND2_X1 U715 ( .A1(n658), .A2(n657), .ZN(n659) );
  XOR2_X1 U716 ( .A(KEYINPUT116), .B(n659), .Z(n660) );
  NAND2_X1 U717 ( .A1(n727), .A2(n660), .ZN(n662) );
  XNOR2_X1 U718 ( .A(KEYINPUT53), .B(KEYINPUT117), .ZN(n661) );
  XNOR2_X1 U719 ( .A(n662), .B(n661), .ZN(G75) );
  NAND2_X1 U720 ( .A1(n688), .A2(G210), .ZN(n668) );
  XOR2_X1 U721 ( .A(KEYINPUT84), .B(KEYINPUT75), .Z(n664) );
  XNOR2_X1 U722 ( .A(KEYINPUT55), .B(KEYINPUT54), .ZN(n663) );
  XNOR2_X1 U723 ( .A(n664), .B(n663), .ZN(n665) );
  XNOR2_X1 U724 ( .A(n666), .B(n665), .ZN(n667) );
  XNOR2_X1 U725 ( .A(n668), .B(n667), .ZN(n669) );
  NOR2_X2 U726 ( .A1(n669), .A2(n722), .ZN(n670) );
  XNOR2_X1 U727 ( .A(n670), .B(KEYINPUT56), .ZN(G51) );
  XNOR2_X1 U728 ( .A(n671), .B(G143), .ZN(G45) );
  NOR2_X1 U729 ( .A1(n672), .A2(G953), .ZN(n678) );
  XOR2_X1 U730 ( .A(KEYINPUT61), .B(KEYINPUT122), .Z(n674) );
  NAND2_X1 U731 ( .A1(G224), .A2(G953), .ZN(n673) );
  XNOR2_X1 U732 ( .A(n674), .B(n673), .ZN(n676) );
  NOR2_X1 U733 ( .A1(n676), .A2(n675), .ZN(n677) );
  NOR2_X1 U734 ( .A1(n678), .A2(n677), .ZN(n683) );
  NAND2_X1 U735 ( .A1(n679), .A2(n680), .ZN(n681) );
  XOR2_X1 U736 ( .A(n681), .B(KEYINPUT123), .Z(n682) );
  XNOR2_X1 U737 ( .A(n683), .B(n682), .ZN(G69) );
  XOR2_X1 U738 ( .A(G131), .B(KEYINPUT126), .Z(n684) );
  XNOR2_X1 U739 ( .A(n685), .B(n684), .ZN(G33) );
  XNOR2_X1 U740 ( .A(n686), .B(G119), .ZN(G21) );
  XNOR2_X1 U741 ( .A(n687), .B(G122), .ZN(G24) );
  NAND2_X1 U742 ( .A1(n688), .A2(G472), .ZN(n691) );
  XNOR2_X1 U743 ( .A(n689), .B(KEYINPUT62), .ZN(n690) );
  XNOR2_X1 U744 ( .A(n691), .B(n690), .ZN(n692) );
  NOR2_X2 U745 ( .A1(n692), .A2(n722), .ZN(n694) );
  XOR2_X1 U746 ( .A(KEYINPUT88), .B(KEYINPUT63), .Z(n693) );
  XNOR2_X1 U747 ( .A(n694), .B(n693), .ZN(G57) );
  XNOR2_X1 U748 ( .A(G101), .B(n695), .ZN(G3) );
  NOR2_X1 U749 ( .A1(n707), .A2(n697), .ZN(n696) );
  XOR2_X1 U750 ( .A(G104), .B(n696), .Z(G6) );
  NOR2_X1 U751 ( .A1(n697), .A2(n710), .ZN(n699) );
  XNOR2_X1 U752 ( .A(KEYINPUT27), .B(KEYINPUT26), .ZN(n698) );
  XNOR2_X1 U753 ( .A(n699), .B(n698), .ZN(n700) );
  XNOR2_X1 U754 ( .A(G107), .B(n700), .ZN(G9) );
  XOR2_X1 U755 ( .A(G110), .B(n701), .Z(G12) );
  XOR2_X1 U756 ( .A(G128), .B(KEYINPUT29), .Z(n704) );
  NAND2_X1 U757 ( .A1(n705), .A2(n702), .ZN(n703) );
  XNOR2_X1 U758 ( .A(n704), .B(n703), .ZN(G30) );
  NAND2_X1 U759 ( .A1(n705), .A2(n368), .ZN(n706) );
  XNOR2_X1 U760 ( .A(G146), .B(n706), .ZN(G48) );
  NOR2_X1 U761 ( .A1(n707), .A2(n709), .ZN(n708) );
  XOR2_X1 U762 ( .A(G113), .B(n708), .Z(G15) );
  NOR2_X1 U763 ( .A1(n710), .A2(n709), .ZN(n711) );
  XOR2_X1 U764 ( .A(G116), .B(n711), .Z(G18) );
  XOR2_X1 U765 ( .A(G125), .B(KEYINPUT37), .Z(n712) );
  XNOR2_X1 U766 ( .A(n713), .B(n712), .ZN(G27) );
  XNOR2_X1 U767 ( .A(n714), .B(G140), .ZN(n715) );
  XNOR2_X1 U768 ( .A(KEYINPUT112), .B(n715), .ZN(G42) );
  NAND2_X1 U769 ( .A1(n716), .A2(G217), .ZN(n720) );
  INV_X1 U770 ( .A(KEYINPUT121), .ZN(n718) );
  NOR2_X1 U771 ( .A1(n722), .A2(n721), .ZN(G66) );
  XNOR2_X1 U772 ( .A(n723), .B(KEYINPUT124), .ZN(n724) );
  XOR2_X1 U773 ( .A(n725), .B(n724), .Z(n729) );
  XNOR2_X1 U774 ( .A(n726), .B(n729), .ZN(n728) );
  NAND2_X1 U775 ( .A1(n728), .A2(n727), .ZN(n734) );
  XOR2_X1 U776 ( .A(n729), .B(G227), .Z(n730) );
  NAND2_X1 U777 ( .A1(n730), .A2(G900), .ZN(n731) );
  XOR2_X1 U778 ( .A(KEYINPUT125), .B(n731), .Z(n732) );
  NAND2_X1 U779 ( .A1(G953), .A2(n732), .ZN(n733) );
  NAND2_X1 U780 ( .A1(n734), .A2(n733), .ZN(G72) );
  XOR2_X1 U781 ( .A(G134), .B(n735), .Z(n736) );
  XNOR2_X1 U782 ( .A(KEYINPUT111), .B(n736), .ZN(G36) );
  XOR2_X1 U783 ( .A(G137), .B(n737), .Z(G39) );
endmodule

