//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 0 0 0 0 1 0 1 1 1 1 1 1 1 0 1 0 0 0 0 1 0 1 1 1 1 0 1 1 1 0 0 0 1 1 0 1 1 1 1 0 1 0 0 1 0 1 1 1 1 1 0 1 0 1 0 1 1 1 0 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:18:07 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n675, new_n676, new_n677, new_n678, new_n680,
    new_n681, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n714, new_n715, new_n716, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n751, new_n752, new_n753, new_n754, new_n755, new_n756,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n763, new_n764,
    new_n765, new_n766, new_n767, new_n768, new_n770, new_n771, new_n773,
    new_n774, new_n775, new_n776, new_n777, new_n778, new_n779, new_n780,
    new_n781, new_n782, new_n783, new_n784, new_n785, new_n786, new_n787,
    new_n788, new_n789, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n804, new_n805, new_n806, new_n807, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n864, new_n865, new_n867, new_n868, new_n869, new_n870, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n911, new_n912, new_n913, new_n914, new_n916, new_n917,
    new_n918, new_n919, new_n920, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n928, new_n929, new_n930, new_n932, new_n933, new_n934,
    new_n935, new_n936, new_n938, new_n939, new_n940, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n961, new_n962, new_n963, new_n965, new_n966, new_n967,
    new_n968;
  INV_X1    g000(.A(KEYINPUT35), .ZN(new_n202));
  XNOR2_X1  g001(.A(G1gat), .B(G29gat), .ZN(new_n203));
  XNOR2_X1  g002(.A(new_n203), .B(G85gat), .ZN(new_n204));
  XNOR2_X1  g003(.A(KEYINPUT0), .B(G57gat), .ZN(new_n205));
  XOR2_X1   g004(.A(new_n204), .B(new_n205), .Z(new_n206));
  INV_X1    g005(.A(KEYINPUT72), .ZN(new_n207));
  INV_X1    g006(.A(G148gat), .ZN(new_n208));
  NOR2_X1   g007(.A1(new_n208), .A2(G141gat), .ZN(new_n209));
  INV_X1    g008(.A(G141gat), .ZN(new_n210));
  NOR2_X1   g009(.A1(new_n210), .A2(G148gat), .ZN(new_n211));
  OAI21_X1  g010(.A(new_n207), .B1(new_n209), .B2(new_n211), .ZN(new_n212));
  NAND2_X1  g011(.A1(G155gat), .A2(G162gat), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n213), .A2(KEYINPUT2), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n210), .A2(G148gat), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n208), .A2(G141gat), .ZN(new_n216));
  NAND3_X1  g015(.A1(new_n215), .A2(new_n216), .A3(KEYINPUT72), .ZN(new_n217));
  NAND3_X1  g016(.A1(new_n212), .A2(new_n214), .A3(new_n217), .ZN(new_n218));
  INV_X1    g017(.A(KEYINPUT71), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n213), .A2(new_n219), .ZN(new_n220));
  NAND3_X1  g019(.A1(KEYINPUT71), .A2(G155gat), .A3(G162gat), .ZN(new_n221));
  INV_X1    g020(.A(G155gat), .ZN(new_n222));
  INV_X1    g021(.A(G162gat), .ZN(new_n223));
  AOI22_X1  g022(.A1(new_n220), .A2(new_n221), .B1(new_n222), .B2(new_n223), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n218), .A2(new_n224), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n222), .A2(KEYINPUT74), .ZN(new_n226));
  INV_X1    g025(.A(KEYINPUT74), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n227), .A2(G155gat), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n226), .A2(new_n228), .ZN(new_n229));
  OAI21_X1  g028(.A(KEYINPUT2), .B1(new_n229), .B2(new_n223), .ZN(new_n230));
  XNOR2_X1  g029(.A(KEYINPUT73), .B(G148gat), .ZN(new_n231));
  OAI21_X1  g030(.A(new_n215), .B1(new_n231), .B2(new_n210), .ZN(new_n232));
  XNOR2_X1  g031(.A(G155gat), .B(G162gat), .ZN(new_n233));
  NAND3_X1  g032(.A1(new_n230), .A2(new_n232), .A3(new_n233), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n225), .A2(new_n234), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n235), .A2(KEYINPUT3), .ZN(new_n236));
  INV_X1    g035(.A(G134gat), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n237), .A2(G127gat), .ZN(new_n238));
  INV_X1    g037(.A(G127gat), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n239), .A2(G134gat), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n238), .A2(new_n240), .ZN(new_n241));
  XNOR2_X1  g040(.A(G113gat), .B(G120gat), .ZN(new_n242));
  OAI21_X1  g041(.A(new_n241), .B1(new_n242), .B2(KEYINPUT1), .ZN(new_n243));
  INV_X1    g042(.A(G120gat), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n244), .A2(G113gat), .ZN(new_n245));
  INV_X1    g044(.A(G113gat), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n246), .A2(G120gat), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n245), .A2(new_n247), .ZN(new_n248));
  XNOR2_X1  g047(.A(G127gat), .B(G134gat), .ZN(new_n249));
  INV_X1    g048(.A(KEYINPUT1), .ZN(new_n250));
  NAND3_X1  g049(.A1(new_n248), .A2(new_n249), .A3(new_n250), .ZN(new_n251));
  AND2_X1   g050(.A1(new_n243), .A2(new_n251), .ZN(new_n252));
  INV_X1    g051(.A(new_n252), .ZN(new_n253));
  INV_X1    g052(.A(KEYINPUT3), .ZN(new_n254));
  NAND3_X1  g053(.A1(new_n225), .A2(new_n254), .A3(new_n234), .ZN(new_n255));
  NAND3_X1  g054(.A1(new_n236), .A2(new_n253), .A3(new_n255), .ZN(new_n256));
  NAND2_X1  g055(.A1(G225gat), .A2(G233gat), .ZN(new_n257));
  NAND3_X1  g056(.A1(new_n225), .A2(new_n252), .A3(new_n234), .ZN(new_n258));
  XNOR2_X1  g057(.A(KEYINPUT75), .B(KEYINPUT4), .ZN(new_n259));
  INV_X1    g058(.A(new_n259), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n258), .A2(new_n260), .ZN(new_n261));
  AND3_X1   g060(.A1(new_n225), .A2(new_n252), .A3(new_n234), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n262), .A2(KEYINPUT4), .ZN(new_n263));
  NAND4_X1  g062(.A1(new_n256), .A2(new_n257), .A3(new_n261), .A4(new_n263), .ZN(new_n264));
  INV_X1    g063(.A(new_n257), .ZN(new_n265));
  AOI21_X1  g064(.A(new_n252), .B1(new_n225), .B2(new_n234), .ZN(new_n266));
  OAI21_X1  g065(.A(new_n265), .B1(new_n262), .B2(new_n266), .ZN(new_n267));
  INV_X1    g066(.A(KEYINPUT76), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  OAI211_X1 g068(.A(KEYINPUT76), .B(new_n265), .C1(new_n262), .C2(new_n266), .ZN(new_n270));
  NAND4_X1  g069(.A1(new_n264), .A2(KEYINPUT5), .A3(new_n269), .A4(new_n270), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n258), .A2(KEYINPUT4), .ZN(new_n272));
  OAI211_X1 g071(.A(new_n272), .B(KEYINPUT77), .C1(new_n258), .C2(new_n259), .ZN(new_n273));
  NOR2_X1   g072(.A1(new_n265), .A2(KEYINPUT5), .ZN(new_n274));
  INV_X1    g073(.A(KEYINPUT77), .ZN(new_n275));
  NAND3_X1  g074(.A1(new_n258), .A2(new_n275), .A3(KEYINPUT4), .ZN(new_n276));
  NAND4_X1  g075(.A1(new_n273), .A2(new_n274), .A3(new_n256), .A4(new_n276), .ZN(new_n277));
  AOI21_X1  g076(.A(new_n206), .B1(new_n271), .B2(new_n277), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n278), .A2(KEYINPUT6), .ZN(new_n279));
  NAND3_X1  g078(.A1(new_n271), .A2(new_n206), .A3(new_n277), .ZN(new_n280));
  INV_X1    g079(.A(KEYINPUT6), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  XOR2_X1   g081(.A(new_n206), .B(KEYINPUT82), .Z(new_n283));
  AOI21_X1  g082(.A(new_n283), .B1(new_n271), .B2(new_n277), .ZN(new_n284));
  OAI21_X1  g083(.A(new_n279), .B1(new_n282), .B2(new_n284), .ZN(new_n285));
  XNOR2_X1  g084(.A(G8gat), .B(G36gat), .ZN(new_n286));
  XNOR2_X1  g085(.A(G64gat), .B(G92gat), .ZN(new_n287));
  XNOR2_X1  g086(.A(new_n286), .B(new_n287), .ZN(new_n288));
  INV_X1    g087(.A(new_n288), .ZN(new_n289));
  NAND2_X1  g088(.A1(G226gat), .A2(G233gat), .ZN(new_n290));
  INV_X1    g089(.A(new_n290), .ZN(new_n291));
  AOI21_X1  g090(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n292));
  OAI21_X1  g091(.A(new_n292), .B1(G169gat), .B2(G176gat), .ZN(new_n293));
  NOR2_X1   g092(.A1(G169gat), .A2(G176gat), .ZN(new_n294));
  AOI22_X1  g093(.A1(new_n294), .A2(KEYINPUT26), .B1(G183gat), .B2(G190gat), .ZN(new_n295));
  INV_X1    g094(.A(KEYINPUT65), .ZN(new_n296));
  AND3_X1   g095(.A1(new_n293), .A2(new_n295), .A3(new_n296), .ZN(new_n297));
  AOI21_X1  g096(.A(new_n296), .B1(new_n293), .B2(new_n295), .ZN(new_n298));
  NOR2_X1   g097(.A1(new_n297), .A2(new_n298), .ZN(new_n299));
  INV_X1    g098(.A(G190gat), .ZN(new_n300));
  INV_X1    g099(.A(KEYINPUT27), .ZN(new_n301));
  OAI21_X1  g100(.A(KEYINPUT64), .B1(new_n301), .B2(G183gat), .ZN(new_n302));
  XNOR2_X1  g101(.A(KEYINPUT27), .B(G183gat), .ZN(new_n303));
  OAI211_X1 g102(.A(new_n300), .B(new_n302), .C1(new_n303), .C2(KEYINPUT64), .ZN(new_n304));
  INV_X1    g103(.A(KEYINPUT28), .ZN(new_n305));
  NOR2_X1   g104(.A1(new_n305), .A2(G190gat), .ZN(new_n306));
  AOI22_X1  g105(.A1(new_n304), .A2(new_n305), .B1(new_n303), .B2(new_n306), .ZN(new_n307));
  OAI21_X1  g106(.A(KEYINPUT66), .B1(new_n299), .B2(new_n307), .ZN(new_n308));
  INV_X1    g107(.A(KEYINPUT23), .ZN(new_n309));
  INV_X1    g108(.A(G169gat), .ZN(new_n310));
  INV_X1    g109(.A(G176gat), .ZN(new_n311));
  NAND3_X1  g110(.A1(new_n309), .A2(new_n310), .A3(new_n311), .ZN(new_n312));
  OAI21_X1  g111(.A(KEYINPUT23), .B1(G169gat), .B2(G176gat), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  INV_X1    g113(.A(G183gat), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n315), .A2(new_n300), .ZN(new_n316));
  NAND2_X1  g115(.A1(G183gat), .A2(G190gat), .ZN(new_n317));
  NAND3_X1  g116(.A1(new_n316), .A2(KEYINPUT24), .A3(new_n317), .ZN(new_n318));
  OR2_X1    g117(.A1(new_n317), .A2(KEYINPUT24), .ZN(new_n319));
  NAND2_X1  g118(.A1(G169gat), .A2(G176gat), .ZN(new_n320));
  NAND4_X1  g119(.A1(new_n314), .A2(new_n318), .A3(new_n319), .A4(new_n320), .ZN(new_n321));
  INV_X1    g120(.A(KEYINPUT25), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  AOI22_X1  g122(.A1(new_n312), .A2(new_n313), .B1(G169gat), .B2(G176gat), .ZN(new_n324));
  NAND4_X1  g123(.A1(new_n324), .A2(KEYINPUT25), .A3(new_n319), .A4(new_n318), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n323), .A2(new_n325), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n293), .A2(new_n295), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n327), .A2(KEYINPUT65), .ZN(new_n328));
  NAND3_X1  g127(.A1(new_n293), .A2(new_n295), .A3(new_n296), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n328), .A2(new_n329), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n315), .A2(KEYINPUT27), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n301), .A2(G183gat), .ZN(new_n332));
  AOI21_X1  g131(.A(KEYINPUT64), .B1(new_n331), .B2(new_n332), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n302), .A2(new_n300), .ZN(new_n334));
  OAI21_X1  g133(.A(new_n305), .B1(new_n333), .B2(new_n334), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n303), .A2(new_n306), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n335), .A2(new_n336), .ZN(new_n337));
  INV_X1    g136(.A(KEYINPUT66), .ZN(new_n338));
  NAND3_X1  g137(.A1(new_n330), .A2(new_n337), .A3(new_n338), .ZN(new_n339));
  NAND3_X1  g138(.A1(new_n308), .A2(new_n326), .A3(new_n339), .ZN(new_n340));
  INV_X1    g139(.A(KEYINPUT29), .ZN(new_n341));
  AOI21_X1  g140(.A(new_n291), .B1(new_n340), .B2(new_n341), .ZN(new_n342));
  AOI22_X1  g141(.A1(new_n330), .A2(new_n337), .B1(new_n323), .B2(new_n325), .ZN(new_n343));
  OAI21_X1  g142(.A(KEYINPUT69), .B1(new_n343), .B2(new_n290), .ZN(new_n344));
  INV_X1    g143(.A(KEYINPUT69), .ZN(new_n345));
  AND2_X1   g144(.A1(new_n323), .A2(new_n325), .ZN(new_n346));
  AOI22_X1  g145(.A1(new_n329), .A2(new_n328), .B1(new_n335), .B2(new_n336), .ZN(new_n347));
  OAI211_X1 g146(.A(new_n345), .B(new_n291), .C1(new_n346), .C2(new_n347), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n344), .A2(new_n348), .ZN(new_n349));
  XNOR2_X1  g148(.A(G197gat), .B(G204gat), .ZN(new_n350));
  INV_X1    g149(.A(G211gat), .ZN(new_n351));
  INV_X1    g150(.A(G218gat), .ZN(new_n352));
  NOR2_X1   g151(.A1(new_n351), .A2(new_n352), .ZN(new_n353));
  OAI21_X1  g152(.A(new_n350), .B1(KEYINPUT22), .B2(new_n353), .ZN(new_n354));
  XNOR2_X1  g153(.A(G211gat), .B(G218gat), .ZN(new_n355));
  XNOR2_X1  g154(.A(new_n354), .B(new_n355), .ZN(new_n356));
  INV_X1    g155(.A(new_n356), .ZN(new_n357));
  NOR3_X1   g156(.A1(new_n342), .A2(new_n349), .A3(new_n357), .ZN(new_n358));
  OAI211_X1 g157(.A(new_n341), .B(new_n290), .C1(new_n346), .C2(new_n347), .ZN(new_n359));
  OAI21_X1  g158(.A(new_n359), .B1(new_n340), .B2(new_n290), .ZN(new_n360));
  NOR2_X1   g159(.A1(new_n360), .A2(new_n356), .ZN(new_n361));
  OAI211_X1 g160(.A(KEYINPUT30), .B(new_n289), .C1(new_n358), .C2(new_n361), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n340), .A2(new_n341), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n363), .A2(new_n290), .ZN(new_n364));
  AND2_X1   g163(.A1(new_n344), .A2(new_n348), .ZN(new_n365));
  NAND3_X1  g164(.A1(new_n364), .A2(new_n356), .A3(new_n365), .ZN(new_n366));
  OR2_X1    g165(.A1(new_n360), .A2(new_n356), .ZN(new_n367));
  NAND3_X1  g166(.A1(new_n366), .A2(new_n367), .A3(new_n288), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n362), .A2(new_n368), .ZN(new_n369));
  INV_X1    g168(.A(new_n369), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n366), .A2(new_n367), .ZN(new_n371));
  AOI21_X1  g170(.A(KEYINPUT30), .B1(new_n371), .B2(new_n289), .ZN(new_n372));
  INV_X1    g171(.A(new_n372), .ZN(new_n373));
  AND4_X1   g172(.A1(new_n202), .A2(new_n285), .A3(new_n370), .A4(new_n373), .ZN(new_n374));
  XNOR2_X1  g173(.A(G15gat), .B(G43gat), .ZN(new_n375));
  INV_X1    g174(.A(G71gat), .ZN(new_n376));
  XNOR2_X1  g175(.A(new_n375), .B(new_n376), .ZN(new_n377));
  XNOR2_X1  g176(.A(new_n377), .B(G99gat), .ZN(new_n378));
  INV_X1    g177(.A(G227gat), .ZN(new_n379));
  INV_X1    g178(.A(G233gat), .ZN(new_n380));
  NOR2_X1   g179(.A1(new_n379), .A2(new_n380), .ZN(new_n381));
  INV_X1    g180(.A(new_n381), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n340), .A2(new_n253), .ZN(new_n383));
  NAND4_X1  g182(.A1(new_n308), .A2(new_n252), .A3(new_n326), .A4(new_n339), .ZN(new_n384));
  AOI21_X1  g183(.A(new_n382), .B1(new_n383), .B2(new_n384), .ZN(new_n385));
  OAI21_X1  g184(.A(new_n378), .B1(new_n385), .B2(KEYINPUT33), .ZN(new_n386));
  INV_X1    g185(.A(KEYINPUT32), .ZN(new_n387));
  NOR2_X1   g186(.A1(new_n385), .A2(new_n387), .ZN(new_n388));
  NOR2_X1   g187(.A1(new_n386), .A2(new_n388), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n383), .A2(new_n384), .ZN(new_n390));
  AOI221_X4 g189(.A(new_n387), .B1(KEYINPUT33), .B2(new_n378), .C1(new_n390), .C2(new_n381), .ZN(new_n391));
  OAI21_X1  g190(.A(KEYINPUT68), .B1(new_n389), .B2(new_n391), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n390), .A2(new_n381), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n393), .A2(KEYINPUT32), .ZN(new_n394));
  INV_X1    g193(.A(KEYINPUT33), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n393), .A2(new_n395), .ZN(new_n396));
  NAND3_X1  g195(.A1(new_n394), .A2(new_n396), .A3(new_n378), .ZN(new_n397));
  INV_X1    g196(.A(KEYINPUT68), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n386), .A2(new_n388), .ZN(new_n399));
  NAND3_X1  g198(.A1(new_n397), .A2(new_n398), .A3(new_n399), .ZN(new_n400));
  NAND3_X1  g199(.A1(new_n383), .A2(new_n382), .A3(new_n384), .ZN(new_n401));
  XNOR2_X1  g200(.A(new_n401), .B(KEYINPUT34), .ZN(new_n402));
  INV_X1    g201(.A(new_n402), .ZN(new_n403));
  NAND3_X1  g202(.A1(new_n392), .A2(new_n400), .A3(new_n403), .ZN(new_n404));
  NAND4_X1  g203(.A1(new_n397), .A2(new_n402), .A3(new_n398), .A4(new_n399), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n404), .A2(new_n405), .ZN(new_n406));
  XNOR2_X1  g205(.A(G78gat), .B(G106gat), .ZN(new_n407));
  XNOR2_X1  g206(.A(new_n407), .B(G22gat), .ZN(new_n408));
  INV_X1    g207(.A(new_n408), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n255), .A2(new_n341), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n410), .A2(new_n356), .ZN(new_n411));
  XNOR2_X1  g210(.A(new_n411), .B(KEYINPUT80), .ZN(new_n412));
  OAI21_X1  g211(.A(new_n254), .B1(new_n356), .B2(KEYINPUT29), .ZN(new_n413));
  NAND2_X1  g212(.A1(new_n413), .A2(new_n235), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n412), .A2(new_n414), .ZN(new_n415));
  NAND2_X1  g214(.A1(G228gat), .A2(G233gat), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n415), .A2(new_n416), .ZN(new_n417));
  NAND4_X1  g216(.A1(new_n411), .A2(new_n414), .A3(G228gat), .A4(G233gat), .ZN(new_n418));
  INV_X1    g217(.A(KEYINPUT81), .ZN(new_n419));
  XNOR2_X1  g218(.A(new_n418), .B(new_n419), .ZN(new_n420));
  XNOR2_X1  g219(.A(KEYINPUT31), .B(G50gat), .ZN(new_n421));
  INV_X1    g220(.A(new_n421), .ZN(new_n422));
  AND3_X1   g221(.A1(new_n417), .A2(new_n420), .A3(new_n422), .ZN(new_n423));
  AOI21_X1  g222(.A(new_n422), .B1(new_n417), .B2(new_n420), .ZN(new_n424));
  OAI21_X1  g223(.A(new_n409), .B1(new_n423), .B2(new_n424), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n417), .A2(new_n420), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n426), .A2(new_n421), .ZN(new_n427));
  NAND3_X1  g226(.A1(new_n417), .A2(new_n420), .A3(new_n422), .ZN(new_n428));
  NAND3_X1  g227(.A1(new_n427), .A2(new_n408), .A3(new_n428), .ZN(new_n429));
  NAND2_X1  g228(.A1(new_n425), .A2(new_n429), .ZN(new_n430));
  AND3_X1   g229(.A1(new_n374), .A2(new_n406), .A3(new_n430), .ZN(new_n431));
  INV_X1    g230(.A(KEYINPUT79), .ZN(new_n432));
  AOI21_X1  g231(.A(new_n278), .B1(new_n282), .B2(KEYINPUT78), .ZN(new_n433));
  INV_X1    g232(.A(KEYINPUT78), .ZN(new_n434));
  NAND3_X1  g233(.A1(new_n280), .A2(new_n434), .A3(new_n281), .ZN(new_n435));
  AOI22_X1  g234(.A1(new_n433), .A2(new_n435), .B1(KEYINPUT6), .B2(new_n278), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n369), .A2(KEYINPUT70), .ZN(new_n437));
  INV_X1    g236(.A(KEYINPUT70), .ZN(new_n438));
  NAND3_X1  g237(.A1(new_n362), .A2(new_n438), .A3(new_n368), .ZN(new_n439));
  NAND3_X1  g238(.A1(new_n437), .A2(new_n439), .A3(new_n373), .ZN(new_n440));
  OAI21_X1  g239(.A(new_n432), .B1(new_n436), .B2(new_n440), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n282), .A2(KEYINPUT78), .ZN(new_n442));
  INV_X1    g241(.A(new_n278), .ZN(new_n443));
  NAND3_X1  g242(.A1(new_n442), .A2(new_n443), .A3(new_n435), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n444), .A2(new_n279), .ZN(new_n445));
  AND3_X1   g244(.A1(new_n362), .A2(new_n438), .A3(new_n368), .ZN(new_n446));
  AOI21_X1  g245(.A(new_n438), .B1(new_n362), .B2(new_n368), .ZN(new_n447));
  NOR3_X1   g246(.A1(new_n446), .A2(new_n447), .A3(new_n372), .ZN(new_n448));
  NAND3_X1  g247(.A1(new_n445), .A2(new_n448), .A3(KEYINPUT79), .ZN(new_n449));
  OAI22_X1  g248(.A1(new_n389), .A2(new_n391), .B1(new_n403), .B2(KEYINPUT67), .ZN(new_n450));
  INV_X1    g249(.A(KEYINPUT67), .ZN(new_n451));
  NAND4_X1  g250(.A1(new_n397), .A2(new_n451), .A3(new_n402), .A4(new_n399), .ZN(new_n452));
  AOI22_X1  g251(.A1(new_n425), .A2(new_n429), .B1(new_n450), .B2(new_n452), .ZN(new_n453));
  NAND3_X1  g252(.A1(new_n441), .A2(new_n449), .A3(new_n453), .ZN(new_n454));
  AOI21_X1  g253(.A(new_n431), .B1(new_n454), .B2(KEYINPUT35), .ZN(new_n455));
  AOI21_X1  g254(.A(new_n430), .B1(new_n441), .B2(new_n449), .ZN(new_n456));
  INV_X1    g255(.A(KEYINPUT36), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n406), .A2(new_n457), .ZN(new_n458));
  NAND3_X1  g257(.A1(new_n450), .A2(KEYINPUT36), .A3(new_n452), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  NOR2_X1   g259(.A1(new_n456), .A2(new_n460), .ZN(new_n461));
  INV_X1    g260(.A(new_n284), .ZN(new_n462));
  INV_X1    g261(.A(new_n272), .ZN(new_n463));
  OAI21_X1  g262(.A(KEYINPUT77), .B1(new_n258), .B2(new_n259), .ZN(new_n464));
  OAI211_X1 g263(.A(new_n256), .B(new_n276), .C1(new_n463), .C2(new_n464), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n465), .A2(new_n265), .ZN(new_n466));
  OR3_X1    g265(.A1(new_n262), .A2(new_n266), .A3(new_n265), .ZN(new_n467));
  NAND3_X1  g266(.A1(new_n466), .A2(KEYINPUT39), .A3(new_n467), .ZN(new_n468));
  INV_X1    g267(.A(new_n468), .ZN(new_n469));
  INV_X1    g268(.A(KEYINPUT83), .ZN(new_n470));
  INV_X1    g269(.A(KEYINPUT39), .ZN(new_n471));
  NAND3_X1  g270(.A1(new_n465), .A2(new_n471), .A3(new_n265), .ZN(new_n472));
  AOI21_X1  g271(.A(new_n470), .B1(new_n472), .B2(new_n283), .ZN(new_n473));
  INV_X1    g272(.A(new_n473), .ZN(new_n474));
  NAND3_X1  g273(.A1(new_n472), .A2(new_n470), .A3(new_n283), .ZN(new_n475));
  AOI21_X1  g274(.A(new_n469), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  OAI21_X1  g275(.A(new_n462), .B1(new_n476), .B2(KEYINPUT40), .ZN(new_n477));
  AND3_X1   g276(.A1(new_n472), .A2(new_n470), .A3(new_n283), .ZN(new_n478));
  OAI211_X1 g277(.A(KEYINPUT40), .B(new_n468), .C1(new_n478), .C2(new_n473), .ZN(new_n479));
  OAI21_X1  g278(.A(new_n479), .B1(new_n369), .B2(new_n372), .ZN(new_n480));
  OAI21_X1  g279(.A(KEYINPUT84), .B1(new_n477), .B2(new_n480), .ZN(new_n481));
  INV_X1    g280(.A(KEYINPUT37), .ZN(new_n482));
  OAI21_X1  g281(.A(new_n482), .B1(new_n358), .B2(new_n361), .ZN(new_n483));
  NAND3_X1  g282(.A1(new_n366), .A2(new_n367), .A3(KEYINPUT37), .ZN(new_n484));
  NAND3_X1  g283(.A1(new_n483), .A2(new_n484), .A3(new_n288), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n485), .A2(KEYINPUT38), .ZN(new_n486));
  INV_X1    g285(.A(KEYINPUT87), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n486), .A2(new_n487), .ZN(new_n488));
  NAND2_X1  g287(.A1(new_n371), .A2(new_n289), .ZN(new_n489));
  OAI211_X1 g288(.A(new_n279), .B(new_n489), .C1(new_n282), .C2(new_n284), .ZN(new_n490));
  INV_X1    g289(.A(new_n490), .ZN(new_n491));
  NAND3_X1  g290(.A1(new_n364), .A2(new_n357), .A3(new_n365), .ZN(new_n492));
  INV_X1    g291(.A(KEYINPUT85), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  OAI211_X1 g293(.A(new_n359), .B(new_n356), .C1(new_n340), .C2(new_n290), .ZN(new_n495));
  OR2_X1    g294(.A1(new_n495), .A2(KEYINPUT86), .ZN(new_n496));
  NAND4_X1  g295(.A1(new_n364), .A2(new_n365), .A3(KEYINPUT85), .A4(new_n357), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n495), .A2(KEYINPUT86), .ZN(new_n498));
  NAND4_X1  g297(.A1(new_n494), .A2(new_n496), .A3(new_n497), .A4(new_n498), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n499), .A2(KEYINPUT37), .ZN(new_n500));
  AOI211_X1 g299(.A(KEYINPUT38), .B(new_n289), .C1(new_n371), .C2(new_n482), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  NAND3_X1  g301(.A1(new_n485), .A2(KEYINPUT87), .A3(KEYINPUT38), .ZN(new_n503));
  NAND4_X1  g302(.A1(new_n488), .A2(new_n491), .A3(new_n502), .A4(new_n503), .ZN(new_n504));
  OAI21_X1  g303(.A(new_n468), .B1(new_n478), .B2(new_n473), .ZN(new_n505));
  INV_X1    g304(.A(KEYINPUT40), .ZN(new_n506));
  AOI21_X1  g305(.A(new_n284), .B1(new_n505), .B2(new_n506), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n370), .A2(new_n373), .ZN(new_n508));
  INV_X1    g307(.A(KEYINPUT84), .ZN(new_n509));
  NAND4_X1  g308(.A1(new_n507), .A2(new_n508), .A3(new_n509), .A4(new_n479), .ZN(new_n510));
  NAND4_X1  g309(.A1(new_n481), .A2(new_n504), .A3(new_n510), .A4(new_n430), .ZN(new_n511));
  AOI21_X1  g310(.A(new_n455), .B1(new_n461), .B2(new_n511), .ZN(new_n512));
  XNOR2_X1  g311(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n513));
  INV_X1    g312(.A(new_n513), .ZN(new_n514));
  XNOR2_X1  g313(.A(G57gat), .B(G64gat), .ZN(new_n515));
  AOI21_X1  g314(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n516));
  OR2_X1    g315(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  XNOR2_X1  g316(.A(G71gat), .B(G78gat), .ZN(new_n518));
  XNOR2_X1  g317(.A(new_n517), .B(new_n518), .ZN(new_n519));
  XNOR2_X1  g318(.A(KEYINPUT94), .B(KEYINPUT21), .ZN(new_n520));
  NOR2_X1   g319(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  INV_X1    g320(.A(new_n521), .ZN(new_n522));
  XNOR2_X1  g321(.A(G15gat), .B(G22gat), .ZN(new_n523));
  OR2_X1    g322(.A1(new_n523), .A2(G1gat), .ZN(new_n524));
  INV_X1    g323(.A(KEYINPUT16), .ZN(new_n525));
  OAI21_X1  g324(.A(new_n523), .B1(new_n525), .B2(G1gat), .ZN(new_n526));
  INV_X1    g325(.A(G8gat), .ZN(new_n527));
  NAND3_X1  g326(.A1(new_n524), .A2(new_n526), .A3(new_n527), .ZN(new_n528));
  XNOR2_X1  g327(.A(new_n528), .B(KEYINPUT92), .ZN(new_n529));
  NAND2_X1  g328(.A1(new_n524), .A2(KEYINPUT91), .ZN(new_n530));
  OR3_X1    g329(.A1(new_n523), .A2(KEYINPUT91), .A3(G1gat), .ZN(new_n531));
  NAND3_X1  g330(.A1(new_n530), .A2(new_n526), .A3(new_n531), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n532), .A2(G8gat), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n529), .A2(new_n533), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n534), .A2(KEYINPUT93), .ZN(new_n535));
  INV_X1    g334(.A(KEYINPUT93), .ZN(new_n536));
  NAND3_X1  g335(.A1(new_n529), .A2(new_n536), .A3(new_n533), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n519), .A2(KEYINPUT21), .ZN(new_n538));
  NAND3_X1  g337(.A1(new_n535), .A2(new_n537), .A3(new_n538), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n539), .A2(G183gat), .ZN(new_n540));
  NAND4_X1  g339(.A1(new_n535), .A2(new_n315), .A3(new_n537), .A4(new_n538), .ZN(new_n541));
  INV_X1    g340(.A(G231gat), .ZN(new_n542));
  NOR2_X1   g341(.A1(new_n542), .A2(new_n380), .ZN(new_n543));
  INV_X1    g342(.A(new_n543), .ZN(new_n544));
  AND3_X1   g343(.A1(new_n540), .A2(new_n541), .A3(new_n544), .ZN(new_n545));
  AOI21_X1  g344(.A(new_n544), .B1(new_n540), .B2(new_n541), .ZN(new_n546));
  OAI21_X1  g345(.A(new_n522), .B1(new_n545), .B2(new_n546), .ZN(new_n547));
  XNOR2_X1  g346(.A(G127gat), .B(G155gat), .ZN(new_n548));
  XNOR2_X1  g347(.A(new_n548), .B(G211gat), .ZN(new_n549));
  INV_X1    g348(.A(new_n549), .ZN(new_n550));
  AND3_X1   g349(.A1(new_n529), .A2(new_n536), .A3(new_n533), .ZN(new_n551));
  AOI21_X1  g350(.A(new_n536), .B1(new_n529), .B2(new_n533), .ZN(new_n552));
  NOR2_X1   g351(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  AOI21_X1  g352(.A(new_n315), .B1(new_n553), .B2(new_n538), .ZN(new_n554));
  INV_X1    g353(.A(new_n541), .ZN(new_n555));
  OAI21_X1  g354(.A(new_n543), .B1(new_n554), .B2(new_n555), .ZN(new_n556));
  NAND3_X1  g355(.A1(new_n540), .A2(new_n541), .A3(new_n544), .ZN(new_n557));
  NAND3_X1  g356(.A1(new_n556), .A2(new_n557), .A3(new_n521), .ZN(new_n558));
  AND3_X1   g357(.A1(new_n547), .A2(new_n550), .A3(new_n558), .ZN(new_n559));
  AOI21_X1  g358(.A(new_n550), .B1(new_n547), .B2(new_n558), .ZN(new_n560));
  OAI21_X1  g359(.A(new_n514), .B1(new_n559), .B2(new_n560), .ZN(new_n561));
  INV_X1    g360(.A(new_n558), .ZN(new_n562));
  AOI21_X1  g361(.A(new_n521), .B1(new_n556), .B2(new_n557), .ZN(new_n563));
  OAI21_X1  g362(.A(new_n549), .B1(new_n562), .B2(new_n563), .ZN(new_n564));
  NAND3_X1  g363(.A1(new_n547), .A2(new_n550), .A3(new_n558), .ZN(new_n565));
  NAND3_X1  g364(.A1(new_n564), .A2(new_n513), .A3(new_n565), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n561), .A2(new_n566), .ZN(new_n567));
  INV_X1    g366(.A(new_n567), .ZN(new_n568));
  XOR2_X1   g367(.A(G43gat), .B(G50gat), .Z(new_n569));
  INV_X1    g368(.A(KEYINPUT15), .ZN(new_n570));
  AOI22_X1  g369(.A1(new_n569), .A2(new_n570), .B1(G29gat), .B2(G36gat), .ZN(new_n571));
  XNOR2_X1  g370(.A(G43gat), .B(G50gat), .ZN(new_n572));
  NAND2_X1  g371(.A1(new_n572), .A2(KEYINPUT15), .ZN(new_n573));
  NOR3_X1   g372(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n574));
  XNOR2_X1  g373(.A(new_n574), .B(KEYINPUT89), .ZN(new_n575));
  OAI21_X1  g374(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n576));
  INV_X1    g375(.A(new_n576), .ZN(new_n577));
  OAI211_X1 g376(.A(new_n571), .B(new_n573), .C1(new_n575), .C2(new_n577), .ZN(new_n578));
  INV_X1    g377(.A(G29gat), .ZN(new_n579));
  INV_X1    g378(.A(G36gat), .ZN(new_n580));
  OAI22_X1  g379(.A1(new_n577), .A2(new_n574), .B1(new_n579), .B2(new_n580), .ZN(new_n581));
  NAND3_X1  g380(.A1(new_n581), .A2(KEYINPUT15), .A3(new_n572), .ZN(new_n582));
  NAND2_X1  g381(.A1(new_n578), .A2(new_n582), .ZN(new_n583));
  XNOR2_X1  g382(.A(new_n583), .B(KEYINPUT90), .ZN(new_n584));
  INV_X1    g383(.A(KEYINPUT17), .ZN(new_n585));
  NAND2_X1  g384(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  NAND3_X1  g385(.A1(new_n578), .A2(KEYINPUT17), .A3(new_n582), .ZN(new_n587));
  XOR2_X1   g386(.A(G99gat), .B(G106gat), .Z(new_n588));
  NAND2_X1  g387(.A1(G99gat), .A2(G106gat), .ZN(new_n589));
  AOI22_X1  g388(.A1(new_n588), .A2(KEYINPUT96), .B1(KEYINPUT8), .B2(new_n589), .ZN(new_n590));
  NAND2_X1  g389(.A1(G85gat), .A2(G92gat), .ZN(new_n591));
  XNOR2_X1  g390(.A(new_n591), .B(KEYINPUT7), .ZN(new_n592));
  OAI211_X1 g391(.A(new_n590), .B(new_n592), .C1(G85gat), .C2(G92gat), .ZN(new_n593));
  NOR2_X1   g392(.A1(new_n588), .A2(KEYINPUT96), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  OR2_X1    g394(.A1(new_n593), .A2(new_n594), .ZN(new_n596));
  NAND4_X1  g395(.A1(new_n586), .A2(new_n587), .A3(new_n595), .A4(new_n596), .ZN(new_n597));
  XNOR2_X1  g396(.A(new_n593), .B(new_n594), .ZN(new_n598));
  NAND2_X1  g397(.A1(new_n584), .A2(new_n598), .ZN(new_n599));
  NAND3_X1  g398(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n600));
  NAND3_X1  g399(.A1(new_n597), .A2(new_n599), .A3(new_n600), .ZN(new_n601));
  XNOR2_X1  g400(.A(G190gat), .B(G218gat), .ZN(new_n602));
  XOR2_X1   g401(.A(new_n602), .B(KEYINPUT97), .Z(new_n603));
  INV_X1    g402(.A(new_n603), .ZN(new_n604));
  NAND2_X1  g403(.A1(new_n601), .A2(new_n604), .ZN(new_n605));
  NAND4_X1  g404(.A1(new_n597), .A2(new_n599), .A3(new_n600), .A4(new_n603), .ZN(new_n606));
  NAND3_X1  g405(.A1(new_n605), .A2(KEYINPUT98), .A3(new_n606), .ZN(new_n607));
  AOI21_X1  g406(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n608));
  XNOR2_X1  g407(.A(new_n608), .B(KEYINPUT95), .ZN(new_n609));
  XNOR2_X1  g408(.A(G134gat), .B(G162gat), .ZN(new_n610));
  XNOR2_X1  g409(.A(new_n609), .B(new_n610), .ZN(new_n611));
  NOR2_X1   g410(.A1(new_n607), .A2(new_n611), .ZN(new_n612));
  NAND2_X1  g411(.A1(new_n605), .A2(new_n606), .ZN(new_n613));
  XNOR2_X1  g412(.A(new_n613), .B(KEYINPUT98), .ZN(new_n614));
  AOI21_X1  g413(.A(new_n612), .B1(new_n614), .B2(new_n611), .ZN(new_n615));
  INV_X1    g414(.A(new_n615), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n568), .A2(new_n616), .ZN(new_n617));
  NOR2_X1   g416(.A1(new_n512), .A2(new_n617), .ZN(new_n618));
  NAND4_X1  g417(.A1(new_n586), .A2(new_n533), .A3(new_n529), .A4(new_n587), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n535), .A2(new_n537), .ZN(new_n620));
  NAND2_X1  g419(.A1(new_n620), .A2(new_n584), .ZN(new_n621));
  AND2_X1   g420(.A1(new_n619), .A2(new_n621), .ZN(new_n622));
  NAND2_X1  g421(.A1(G229gat), .A2(G233gat), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  INV_X1    g423(.A(KEYINPUT18), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  XNOR2_X1  g425(.A(new_n620), .B(new_n584), .ZN(new_n627));
  XOR2_X1   g426(.A(new_n623), .B(KEYINPUT13), .Z(new_n628));
  NAND2_X1  g427(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  NAND3_X1  g428(.A1(new_n622), .A2(KEYINPUT18), .A3(new_n623), .ZN(new_n630));
  NAND3_X1  g429(.A1(new_n626), .A2(new_n629), .A3(new_n630), .ZN(new_n631));
  XOR2_X1   g430(.A(KEYINPUT88), .B(KEYINPUT11), .Z(new_n632));
  XNOR2_X1  g431(.A(G169gat), .B(G197gat), .ZN(new_n633));
  XNOR2_X1  g432(.A(new_n632), .B(new_n633), .ZN(new_n634));
  XNOR2_X1  g433(.A(G113gat), .B(G141gat), .ZN(new_n635));
  XNOR2_X1  g434(.A(new_n634), .B(new_n635), .ZN(new_n636));
  XOR2_X1   g435(.A(new_n636), .B(KEYINPUT12), .Z(new_n637));
  NAND2_X1  g436(.A1(new_n631), .A2(new_n637), .ZN(new_n638));
  INV_X1    g437(.A(new_n637), .ZN(new_n639));
  NAND4_X1  g438(.A1(new_n626), .A2(new_n639), .A3(new_n629), .A4(new_n630), .ZN(new_n640));
  AND2_X1   g439(.A1(new_n638), .A2(new_n640), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n598), .A2(new_n519), .ZN(new_n642));
  INV_X1    g441(.A(KEYINPUT10), .ZN(new_n643));
  INV_X1    g442(.A(new_n519), .ZN(new_n644));
  NAND3_X1  g443(.A1(new_n596), .A2(new_n644), .A3(new_n595), .ZN(new_n645));
  NAND3_X1  g444(.A1(new_n642), .A2(new_n643), .A3(new_n645), .ZN(new_n646));
  NAND3_X1  g445(.A1(new_n598), .A2(KEYINPUT10), .A3(new_n519), .ZN(new_n647));
  INV_X1    g446(.A(KEYINPUT99), .ZN(new_n648));
  NAND2_X1  g447(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  NAND4_X1  g448(.A1(new_n598), .A2(KEYINPUT99), .A3(KEYINPUT10), .A4(new_n519), .ZN(new_n650));
  NAND3_X1  g449(.A1(new_n646), .A2(new_n649), .A3(new_n650), .ZN(new_n651));
  NAND2_X1  g450(.A1(G230gat), .A2(G233gat), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  AND2_X1   g452(.A1(new_n642), .A2(new_n645), .ZN(new_n654));
  OAI21_X1  g453(.A(new_n653), .B1(new_n652), .B2(new_n654), .ZN(new_n655));
  XNOR2_X1  g454(.A(G120gat), .B(G148gat), .ZN(new_n656));
  XNOR2_X1  g455(.A(G176gat), .B(G204gat), .ZN(new_n657));
  XNOR2_X1  g456(.A(new_n656), .B(new_n657), .ZN(new_n658));
  OR2_X1    g457(.A1(new_n655), .A2(new_n658), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n655), .A2(new_n658), .ZN(new_n660));
  NAND2_X1  g459(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  NOR2_X1   g460(.A1(new_n641), .A2(new_n661), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n618), .A2(new_n662), .ZN(new_n663));
  INV_X1    g462(.A(new_n663), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n664), .A2(new_n436), .ZN(new_n665));
  XNOR2_X1  g464(.A(new_n665), .B(G1gat), .ZN(G1324gat));
  INV_X1    g465(.A(new_n508), .ZN(new_n667));
  NOR2_X1   g466(.A1(new_n663), .A2(new_n667), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n525), .A2(new_n527), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  AOI21_X1  g469(.A(new_n670), .B1(KEYINPUT16), .B2(G8gat), .ZN(new_n671));
  OR2_X1    g470(.A1(new_n671), .A2(KEYINPUT42), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n671), .A2(KEYINPUT42), .ZN(new_n673));
  OAI211_X1 g472(.A(new_n672), .B(new_n673), .C1(new_n527), .C2(new_n668), .ZN(G1325gat));
  INV_X1    g473(.A(G15gat), .ZN(new_n675));
  AND2_X1   g474(.A1(new_n458), .A2(new_n459), .ZN(new_n676));
  NOR3_X1   g475(.A1(new_n663), .A2(new_n675), .A3(new_n676), .ZN(new_n677));
  NAND2_X1  g476(.A1(new_n664), .A2(new_n406), .ZN(new_n678));
  AOI21_X1  g477(.A(new_n677), .B1(new_n675), .B2(new_n678), .ZN(G1326gat));
  NOR2_X1   g478(.A1(new_n663), .A2(new_n430), .ZN(new_n680));
  XOR2_X1   g479(.A(KEYINPUT43), .B(G22gat), .Z(new_n681));
  XNOR2_X1  g480(.A(new_n680), .B(new_n681), .ZN(G1327gat));
  NAND2_X1  g481(.A1(new_n454), .A2(KEYINPUT35), .ZN(new_n683));
  INV_X1    g482(.A(new_n431), .ZN(new_n684));
  NAND2_X1  g483(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  INV_X1    g484(.A(new_n430), .ZN(new_n686));
  NOR3_X1   g485(.A1(new_n436), .A2(new_n440), .A3(new_n432), .ZN(new_n687));
  AOI21_X1  g486(.A(KEYINPUT79), .B1(new_n445), .B2(new_n448), .ZN(new_n688));
  OAI21_X1  g487(.A(new_n686), .B1(new_n687), .B2(new_n688), .ZN(new_n689));
  NAND3_X1  g488(.A1(new_n689), .A2(new_n676), .A3(new_n511), .ZN(new_n690));
  AOI21_X1  g489(.A(new_n616), .B1(new_n685), .B2(new_n690), .ZN(new_n691));
  NAND2_X1  g490(.A1(new_n662), .A2(new_n567), .ZN(new_n692));
  INV_X1    g491(.A(new_n692), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n691), .A2(new_n693), .ZN(new_n694));
  INV_X1    g493(.A(new_n694), .ZN(new_n695));
  NAND3_X1  g494(.A1(new_n695), .A2(new_n579), .A3(new_n436), .ZN(new_n696));
  XNOR2_X1  g495(.A(new_n696), .B(KEYINPUT45), .ZN(new_n697));
  NOR2_X1   g496(.A1(KEYINPUT100), .A2(KEYINPUT44), .ZN(new_n698));
  NAND2_X1  g497(.A1(new_n685), .A2(new_n690), .ZN(new_n699));
  AOI21_X1  g498(.A(new_n698), .B1(new_n699), .B2(new_n615), .ZN(new_n700));
  XOR2_X1   g499(.A(KEYINPUT100), .B(KEYINPUT44), .Z(new_n701));
  AOI211_X1 g500(.A(new_n616), .B(new_n701), .C1(new_n685), .C2(new_n690), .ZN(new_n702));
  OAI21_X1  g501(.A(new_n693), .B1(new_n700), .B2(new_n702), .ZN(new_n703));
  INV_X1    g502(.A(KEYINPUT101), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  INV_X1    g504(.A(new_n701), .ZN(new_n706));
  AND4_X1   g505(.A1(new_n430), .A2(new_n481), .A3(new_n504), .A4(new_n510), .ZN(new_n707));
  NOR3_X1   g506(.A1(new_n707), .A2(new_n456), .A3(new_n460), .ZN(new_n708));
  OAI211_X1 g507(.A(new_n615), .B(new_n706), .C1(new_n708), .C2(new_n455), .ZN(new_n709));
  OAI21_X1  g508(.A(new_n709), .B1(new_n691), .B2(new_n698), .ZN(new_n710));
  NAND3_X1  g509(.A1(new_n710), .A2(KEYINPUT101), .A3(new_n693), .ZN(new_n711));
  AOI21_X1  g510(.A(new_n445), .B1(new_n705), .B2(new_n711), .ZN(new_n712));
  OAI21_X1  g511(.A(new_n697), .B1(new_n712), .B2(new_n579), .ZN(G1328gat));
  NOR3_X1   g512(.A1(new_n694), .A2(G36gat), .A3(new_n667), .ZN(new_n714));
  XNOR2_X1  g513(.A(new_n714), .B(KEYINPUT46), .ZN(new_n715));
  AOI21_X1  g514(.A(new_n667), .B1(new_n705), .B2(new_n711), .ZN(new_n716));
  OAI21_X1  g515(.A(new_n715), .B1(new_n716), .B2(new_n580), .ZN(G1329gat));
  OAI21_X1  g516(.A(G43gat), .B1(new_n703), .B2(new_n676), .ZN(new_n718));
  INV_X1    g517(.A(new_n406), .ZN(new_n719));
  NOR3_X1   g518(.A1(new_n694), .A2(G43gat), .A3(new_n719), .ZN(new_n720));
  INV_X1    g519(.A(new_n720), .ZN(new_n721));
  NAND3_X1  g520(.A1(new_n718), .A2(KEYINPUT47), .A3(new_n721), .ZN(new_n722));
  INV_X1    g521(.A(new_n698), .ZN(new_n723));
  OAI21_X1  g522(.A(new_n723), .B1(new_n512), .B2(new_n616), .ZN(new_n724));
  AOI211_X1 g523(.A(new_n704), .B(new_n692), .C1(new_n724), .C2(new_n709), .ZN(new_n725));
  AOI21_X1  g524(.A(KEYINPUT101), .B1(new_n710), .B2(new_n693), .ZN(new_n726));
  OAI21_X1  g525(.A(new_n460), .B1(new_n725), .B2(new_n726), .ZN(new_n727));
  AOI21_X1  g526(.A(new_n720), .B1(new_n727), .B2(G43gat), .ZN(new_n728));
  OAI21_X1  g527(.A(new_n722), .B1(new_n728), .B2(KEYINPUT47), .ZN(G1330gat));
  INV_X1    g528(.A(KEYINPUT102), .ZN(new_n730));
  AOI21_X1  g529(.A(new_n430), .B1(new_n705), .B2(new_n711), .ZN(new_n731));
  INV_X1    g530(.A(G50gat), .ZN(new_n732));
  OAI21_X1  g531(.A(new_n730), .B1(new_n731), .B2(new_n732), .ZN(new_n733));
  NAND3_X1  g532(.A1(new_n695), .A2(new_n732), .A3(new_n686), .ZN(new_n734));
  OAI21_X1  g533(.A(new_n686), .B1(new_n725), .B2(new_n726), .ZN(new_n735));
  NAND3_X1  g534(.A1(new_n735), .A2(KEYINPUT102), .A3(G50gat), .ZN(new_n736));
  NAND3_X1  g535(.A1(new_n733), .A2(new_n734), .A3(new_n736), .ZN(new_n737));
  INV_X1    g536(.A(KEYINPUT48), .ZN(new_n738));
  NAND2_X1  g537(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  OAI21_X1  g538(.A(G50gat), .B1(new_n703), .B2(new_n430), .ZN(new_n740));
  NAND3_X1  g539(.A1(new_n740), .A2(KEYINPUT48), .A3(new_n734), .ZN(new_n741));
  XNOR2_X1  g540(.A(new_n741), .B(KEYINPUT103), .ZN(new_n742));
  NAND2_X1  g541(.A1(new_n739), .A2(new_n742), .ZN(G1331gat));
  NAND3_X1  g542(.A1(new_n618), .A2(new_n641), .A3(new_n661), .ZN(new_n744));
  OR2_X1    g543(.A1(new_n744), .A2(KEYINPUT104), .ZN(new_n745));
  NAND2_X1  g544(.A1(new_n744), .A2(KEYINPUT104), .ZN(new_n746));
  NAND2_X1  g545(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  NOR2_X1   g546(.A1(new_n747), .A2(new_n445), .ZN(new_n748));
  XNOR2_X1  g547(.A(KEYINPUT105), .B(G57gat), .ZN(new_n749));
  XNOR2_X1  g548(.A(new_n748), .B(new_n749), .ZN(G1332gat));
  NOR2_X1   g549(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n751));
  XNOR2_X1  g550(.A(new_n751), .B(KEYINPUT107), .ZN(new_n752));
  NAND2_X1  g551(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n753));
  NAND4_X1  g552(.A1(new_n745), .A2(new_n508), .A3(new_n746), .A4(new_n753), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n754), .A2(KEYINPUT106), .ZN(new_n755));
  INV_X1    g554(.A(new_n755), .ZN(new_n756));
  NOR2_X1   g555(.A1(new_n754), .A2(KEYINPUT106), .ZN(new_n757));
  OAI21_X1  g556(.A(new_n752), .B1(new_n756), .B2(new_n757), .ZN(new_n758));
  INV_X1    g557(.A(new_n757), .ZN(new_n759));
  INV_X1    g558(.A(new_n752), .ZN(new_n760));
  NAND3_X1  g559(.A1(new_n759), .A2(new_n755), .A3(new_n760), .ZN(new_n761));
  NAND2_X1  g560(.A1(new_n758), .A2(new_n761), .ZN(G1333gat));
  OAI21_X1  g561(.A(new_n376), .B1(new_n747), .B2(new_n719), .ZN(new_n763));
  NAND4_X1  g562(.A1(new_n745), .A2(G71gat), .A3(new_n460), .A4(new_n746), .ZN(new_n764));
  NAND2_X1  g563(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  NAND2_X1  g564(.A1(new_n765), .A2(KEYINPUT50), .ZN(new_n766));
  INV_X1    g565(.A(KEYINPUT50), .ZN(new_n767));
  NAND3_X1  g566(.A1(new_n763), .A2(new_n767), .A3(new_n764), .ZN(new_n768));
  NAND2_X1  g567(.A1(new_n766), .A2(new_n768), .ZN(G1334gat));
  NOR2_X1   g568(.A1(new_n747), .A2(new_n430), .ZN(new_n770));
  XNOR2_X1  g569(.A(KEYINPUT108), .B(G78gat), .ZN(new_n771));
  XNOR2_X1  g570(.A(new_n770), .B(new_n771), .ZN(G1335gat));
  NAND2_X1  g571(.A1(new_n567), .A2(new_n641), .ZN(new_n773));
  INV_X1    g572(.A(KEYINPUT109), .ZN(new_n774));
  XNOR2_X1  g573(.A(new_n773), .B(new_n774), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n691), .A2(new_n775), .ZN(new_n776));
  INV_X1    g575(.A(KEYINPUT51), .ZN(new_n777));
  NAND2_X1  g576(.A1(new_n776), .A2(new_n777), .ZN(new_n778));
  NAND2_X1  g577(.A1(new_n778), .A2(KEYINPUT110), .ZN(new_n779));
  NAND3_X1  g578(.A1(new_n691), .A2(new_n775), .A3(KEYINPUT51), .ZN(new_n780));
  INV_X1    g579(.A(KEYINPUT110), .ZN(new_n781));
  NAND3_X1  g580(.A1(new_n776), .A2(new_n781), .A3(new_n777), .ZN(new_n782));
  NAND3_X1  g581(.A1(new_n779), .A2(new_n780), .A3(new_n782), .ZN(new_n783));
  INV_X1    g582(.A(new_n783), .ZN(new_n784));
  INV_X1    g583(.A(new_n661), .ZN(new_n785));
  OR4_X1    g584(.A1(G85gat), .A2(new_n784), .A3(new_n445), .A4(new_n785), .ZN(new_n786));
  AOI21_X1  g585(.A(new_n785), .B1(new_n724), .B2(new_n709), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n787), .A2(new_n775), .ZN(new_n788));
  OAI21_X1  g587(.A(G85gat), .B1(new_n788), .B2(new_n445), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n786), .A2(new_n789), .ZN(G1336gat));
  INV_X1    g589(.A(KEYINPUT52), .ZN(new_n791));
  AND3_X1   g590(.A1(new_n776), .A2(KEYINPUT112), .A3(new_n777), .ZN(new_n792));
  AOI21_X1  g591(.A(new_n776), .B1(KEYINPUT112), .B2(new_n777), .ZN(new_n793));
  OR2_X1    g592(.A1(new_n792), .A2(new_n793), .ZN(new_n794));
  OR3_X1    g593(.A1(new_n785), .A2(G92gat), .A3(new_n667), .ZN(new_n795));
  XNOR2_X1  g594(.A(new_n795), .B(KEYINPUT111), .ZN(new_n796));
  INV_X1    g595(.A(new_n796), .ZN(new_n797));
  NAND3_X1  g596(.A1(new_n787), .A2(new_n508), .A3(new_n775), .ZN(new_n798));
  AOI22_X1  g597(.A1(new_n794), .A2(new_n797), .B1(new_n798), .B2(G92gat), .ZN(new_n799));
  NOR2_X1   g598(.A1(new_n784), .A2(new_n796), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n798), .A2(G92gat), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n801), .A2(new_n791), .ZN(new_n802));
  OAI22_X1  g601(.A1(new_n791), .A2(new_n799), .B1(new_n800), .B2(new_n802), .ZN(G1337gat));
  XNOR2_X1  g602(.A(KEYINPUT113), .B(G99gat), .ZN(new_n804));
  OAI21_X1  g603(.A(new_n804), .B1(new_n788), .B2(new_n676), .ZN(new_n805));
  NOR3_X1   g604(.A1(new_n719), .A2(new_n785), .A3(new_n804), .ZN(new_n806));
  XOR2_X1   g605(.A(new_n806), .B(KEYINPUT114), .Z(new_n807));
  OAI21_X1  g606(.A(new_n805), .B1(new_n784), .B2(new_n807), .ZN(G1338gat));
  NOR2_X1   g607(.A1(new_n430), .A2(G106gat), .ZN(new_n809));
  NAND3_X1  g608(.A1(new_n783), .A2(new_n661), .A3(new_n809), .ZN(new_n810));
  INV_X1    g609(.A(KEYINPUT53), .ZN(new_n811));
  OAI21_X1  g610(.A(G106gat), .B1(new_n788), .B2(new_n430), .ZN(new_n812));
  AND3_X1   g611(.A1(new_n810), .A2(new_n811), .A3(new_n812), .ZN(new_n813));
  OAI211_X1 g612(.A(new_n661), .B(new_n809), .C1(new_n792), .C2(new_n793), .ZN(new_n814));
  AOI21_X1  g613(.A(new_n811), .B1(new_n812), .B2(new_n814), .ZN(new_n815));
  OAI21_X1  g614(.A(KEYINPUT115), .B1(new_n813), .B2(new_n815), .ZN(new_n816));
  NAND3_X1  g615(.A1(new_n810), .A2(new_n811), .A3(new_n812), .ZN(new_n817));
  INV_X1    g616(.A(KEYINPUT115), .ZN(new_n818));
  AND2_X1   g617(.A1(new_n812), .A2(new_n814), .ZN(new_n819));
  OAI211_X1 g618(.A(new_n817), .B(new_n818), .C1(new_n819), .C2(new_n811), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n816), .A2(new_n820), .ZN(G1339gat));
  INV_X1    g620(.A(new_n652), .ZN(new_n822));
  NAND4_X1  g621(.A1(new_n649), .A2(new_n646), .A3(new_n822), .A4(new_n650), .ZN(new_n823));
  NAND3_X1  g622(.A1(new_n653), .A2(KEYINPUT54), .A3(new_n823), .ZN(new_n824));
  INV_X1    g623(.A(KEYINPUT54), .ZN(new_n825));
  NAND3_X1  g624(.A1(new_n651), .A2(new_n825), .A3(new_n652), .ZN(new_n826));
  NAND3_X1  g625(.A1(new_n824), .A2(new_n658), .A3(new_n826), .ZN(new_n827));
  INV_X1    g626(.A(KEYINPUT55), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n827), .A2(new_n828), .ZN(new_n829));
  NAND4_X1  g628(.A1(new_n824), .A2(KEYINPUT55), .A3(new_n658), .A4(new_n826), .ZN(new_n830));
  NAND3_X1  g629(.A1(new_n829), .A2(new_n659), .A3(new_n830), .ZN(new_n831));
  INV_X1    g630(.A(KEYINPUT116), .ZN(new_n832));
  NAND2_X1  g631(.A1(new_n831), .A2(new_n832), .ZN(new_n833));
  NAND2_X1  g632(.A1(new_n638), .A2(new_n640), .ZN(new_n834));
  NAND4_X1  g633(.A1(new_n829), .A2(new_n830), .A3(new_n659), .A4(KEYINPUT116), .ZN(new_n835));
  NAND3_X1  g634(.A1(new_n833), .A2(new_n834), .A3(new_n835), .ZN(new_n836));
  NOR2_X1   g635(.A1(new_n622), .A2(new_n623), .ZN(new_n837));
  NOR2_X1   g636(.A1(new_n627), .A2(new_n628), .ZN(new_n838));
  OAI21_X1  g637(.A(new_n636), .B1(new_n837), .B2(new_n838), .ZN(new_n839));
  AND2_X1   g638(.A1(new_n640), .A2(new_n839), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n840), .A2(new_n661), .ZN(new_n841));
  AOI21_X1  g640(.A(new_n615), .B1(new_n836), .B2(new_n841), .ZN(new_n842));
  AND4_X1   g641(.A1(new_n615), .A2(new_n833), .A3(new_n835), .A4(new_n840), .ZN(new_n843));
  OAI21_X1  g642(.A(new_n567), .B1(new_n842), .B2(new_n843), .ZN(new_n844));
  NAND4_X1  g643(.A1(new_n568), .A2(new_n616), .A3(new_n641), .A4(new_n785), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  AND2_X1   g645(.A1(new_n846), .A2(new_n453), .ZN(new_n847));
  NOR2_X1   g646(.A1(new_n445), .A2(new_n508), .ZN(new_n848));
  AND2_X1   g647(.A1(new_n847), .A2(new_n848), .ZN(new_n849));
  NAND3_X1  g648(.A1(new_n849), .A2(new_n246), .A3(new_n834), .ZN(new_n850));
  NOR2_X1   g649(.A1(new_n719), .A2(new_n686), .ZN(new_n851));
  AND3_X1   g650(.A1(new_n846), .A2(new_n851), .A3(new_n848), .ZN(new_n852));
  INV_X1    g651(.A(new_n852), .ZN(new_n853));
  OAI21_X1  g652(.A(G113gat), .B1(new_n853), .B2(new_n641), .ZN(new_n854));
  NAND2_X1  g653(.A1(new_n850), .A2(new_n854), .ZN(G1340gat));
  NAND3_X1  g654(.A1(new_n849), .A2(new_n244), .A3(new_n661), .ZN(new_n856));
  INV_X1    g655(.A(KEYINPUT117), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n852), .A2(new_n661), .ZN(new_n858));
  AOI21_X1  g657(.A(new_n857), .B1(new_n858), .B2(G120gat), .ZN(new_n859));
  AOI211_X1 g658(.A(KEYINPUT117), .B(new_n244), .C1(new_n852), .C2(new_n661), .ZN(new_n860));
  OAI21_X1  g659(.A(new_n856), .B1(new_n859), .B2(new_n860), .ZN(new_n861));
  INV_X1    g660(.A(KEYINPUT118), .ZN(new_n862));
  XNOR2_X1  g661(.A(new_n861), .B(new_n862), .ZN(G1341gat));
  AOI21_X1  g662(.A(G127gat), .B1(new_n849), .B2(new_n568), .ZN(new_n864));
  NOR2_X1   g663(.A1(new_n567), .A2(new_n239), .ZN(new_n865));
  AOI21_X1  g664(.A(new_n864), .B1(new_n852), .B2(new_n865), .ZN(G1342gat));
  NAND3_X1  g665(.A1(new_n849), .A2(new_n237), .A3(new_n615), .ZN(new_n867));
  XOR2_X1   g666(.A(new_n867), .B(KEYINPUT56), .Z(new_n868));
  AOI21_X1  g667(.A(new_n237), .B1(new_n852), .B2(new_n615), .ZN(new_n869));
  XOR2_X1   g668(.A(new_n869), .B(KEYINPUT119), .Z(new_n870));
  NAND2_X1  g669(.A1(new_n868), .A2(new_n870), .ZN(G1343gat));
  NAND2_X1  g670(.A1(new_n846), .A2(new_n686), .ZN(new_n872));
  INV_X1    g671(.A(KEYINPUT120), .ZN(new_n873));
  INV_X1    g672(.A(KEYINPUT57), .ZN(new_n874));
  NAND3_X1  g673(.A1(new_n872), .A2(new_n873), .A3(new_n874), .ZN(new_n875));
  OAI21_X1  g674(.A(new_n841), .B1(new_n641), .B2(new_n831), .ZN(new_n876));
  AOI21_X1  g675(.A(new_n843), .B1(new_n616), .B2(new_n876), .ZN(new_n877));
  OAI21_X1  g676(.A(new_n845), .B1(new_n877), .B2(new_n568), .ZN(new_n878));
  NAND3_X1  g677(.A1(new_n878), .A2(KEYINPUT57), .A3(new_n686), .ZN(new_n879));
  AOI21_X1  g678(.A(new_n430), .B1(new_n844), .B2(new_n845), .ZN(new_n880));
  OAI21_X1  g679(.A(KEYINPUT120), .B1(new_n880), .B2(KEYINPUT57), .ZN(new_n881));
  NAND3_X1  g680(.A1(new_n875), .A2(new_n879), .A3(new_n881), .ZN(new_n882));
  NAND2_X1  g681(.A1(new_n676), .A2(new_n848), .ZN(new_n883));
  INV_X1    g682(.A(new_n883), .ZN(new_n884));
  NAND3_X1  g683(.A1(new_n882), .A2(new_n834), .A3(new_n884), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n885), .A2(G141gat), .ZN(new_n886));
  NOR2_X1   g685(.A1(new_n872), .A2(new_n883), .ZN(new_n887));
  NAND3_X1  g686(.A1(new_n887), .A2(new_n210), .A3(new_n834), .ZN(new_n888));
  NAND2_X1  g687(.A1(new_n886), .A2(new_n888), .ZN(new_n889));
  NAND2_X1  g688(.A1(new_n889), .A2(KEYINPUT58), .ZN(new_n890));
  INV_X1    g689(.A(KEYINPUT58), .ZN(new_n891));
  NAND3_X1  g690(.A1(new_n886), .A2(new_n891), .A3(new_n888), .ZN(new_n892));
  NAND2_X1  g691(.A1(new_n890), .A2(new_n892), .ZN(G1344gat));
  INV_X1    g692(.A(KEYINPUT59), .ZN(new_n894));
  NAND2_X1  g693(.A1(new_n882), .A2(new_n884), .ZN(new_n895));
  OAI211_X1 g694(.A(new_n894), .B(new_n231), .C1(new_n895), .C2(new_n785), .ZN(new_n896));
  NAND2_X1  g695(.A1(new_n872), .A2(KEYINPUT57), .ZN(new_n897));
  NAND2_X1  g696(.A1(new_n876), .A2(new_n616), .ZN(new_n898));
  INV_X1    g697(.A(new_n831), .ZN(new_n899));
  NAND3_X1  g698(.A1(new_n615), .A2(new_n899), .A3(new_n840), .ZN(new_n900));
  AOI21_X1  g699(.A(new_n568), .B1(new_n898), .B2(new_n900), .ZN(new_n901));
  INV_X1    g700(.A(new_n845), .ZN(new_n902));
  OAI211_X1 g701(.A(new_n874), .B(new_n686), .C1(new_n901), .C2(new_n902), .ZN(new_n903));
  NAND3_X1  g702(.A1(new_n897), .A2(new_n661), .A3(new_n903), .ZN(new_n904));
  INV_X1    g703(.A(new_n904), .ZN(new_n905));
  AOI21_X1  g704(.A(new_n208), .B1(new_n905), .B2(new_n884), .ZN(new_n906));
  OAI21_X1  g705(.A(new_n896), .B1(new_n894), .B2(new_n906), .ZN(new_n907));
  INV_X1    g706(.A(new_n231), .ZN(new_n908));
  NAND3_X1  g707(.A1(new_n887), .A2(new_n908), .A3(new_n661), .ZN(new_n909));
  NAND2_X1  g708(.A1(new_n907), .A2(new_n909), .ZN(G1345gat));
  INV_X1    g709(.A(new_n895), .ZN(new_n911));
  NOR2_X1   g710(.A1(new_n567), .A2(new_n229), .ZN(new_n912));
  XNOR2_X1  g711(.A(new_n912), .B(KEYINPUT121), .ZN(new_n913));
  NAND2_X1  g712(.A1(new_n887), .A2(new_n568), .ZN(new_n914));
  AOI22_X1  g713(.A1(new_n911), .A2(new_n913), .B1(new_n229), .B2(new_n914), .ZN(G1346gat));
  NAND3_X1  g714(.A1(new_n911), .A2(KEYINPUT122), .A3(new_n615), .ZN(new_n916));
  INV_X1    g715(.A(KEYINPUT122), .ZN(new_n917));
  OAI21_X1  g716(.A(new_n917), .B1(new_n895), .B2(new_n616), .ZN(new_n918));
  NAND3_X1  g717(.A1(new_n916), .A2(G162gat), .A3(new_n918), .ZN(new_n919));
  NAND3_X1  g718(.A1(new_n887), .A2(new_n223), .A3(new_n615), .ZN(new_n920));
  NAND2_X1  g719(.A1(new_n919), .A2(new_n920), .ZN(G1347gat));
  NOR2_X1   g720(.A1(new_n667), .A2(new_n436), .ZN(new_n922));
  AND2_X1   g721(.A1(new_n847), .A2(new_n922), .ZN(new_n923));
  NAND3_X1  g722(.A1(new_n923), .A2(new_n310), .A3(new_n834), .ZN(new_n924));
  NAND3_X1  g723(.A1(new_n846), .A2(new_n851), .A3(new_n922), .ZN(new_n925));
  OAI21_X1  g724(.A(G169gat), .B1(new_n925), .B2(new_n641), .ZN(new_n926));
  NAND2_X1  g725(.A1(new_n924), .A2(new_n926), .ZN(G1348gat));
  NAND3_X1  g726(.A1(new_n923), .A2(new_n311), .A3(new_n661), .ZN(new_n928));
  OAI21_X1  g727(.A(G176gat), .B1(new_n925), .B2(new_n785), .ZN(new_n929));
  NAND2_X1  g728(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  XNOR2_X1  g729(.A(new_n930), .B(KEYINPUT123), .ZN(G1349gat));
  NAND3_X1  g730(.A1(new_n923), .A2(new_n303), .A3(new_n568), .ZN(new_n932));
  NAND2_X1  g731(.A1(KEYINPUT124), .A2(KEYINPUT60), .ZN(new_n933));
  OAI21_X1  g732(.A(G183gat), .B1(new_n925), .B2(new_n567), .ZN(new_n934));
  NAND3_X1  g733(.A1(new_n932), .A2(new_n933), .A3(new_n934), .ZN(new_n935));
  NOR2_X1   g734(.A1(KEYINPUT124), .A2(KEYINPUT60), .ZN(new_n936));
  XOR2_X1   g735(.A(new_n935), .B(new_n936), .Z(G1350gat));
  OAI21_X1  g736(.A(G190gat), .B1(new_n925), .B2(new_n616), .ZN(new_n938));
  XNOR2_X1  g737(.A(new_n938), .B(KEYINPUT61), .ZN(new_n939));
  NAND3_X1  g738(.A1(new_n923), .A2(new_n300), .A3(new_n615), .ZN(new_n940));
  NAND2_X1  g739(.A1(new_n939), .A2(new_n940), .ZN(G1351gat));
  NAND2_X1  g740(.A1(new_n676), .A2(new_n922), .ZN(new_n942));
  INV_X1    g741(.A(new_n942), .ZN(new_n943));
  NAND3_X1  g742(.A1(new_n897), .A2(new_n903), .A3(new_n943), .ZN(new_n944));
  OAI21_X1  g743(.A(G197gat), .B1(new_n944), .B2(new_n641), .ZN(new_n945));
  NAND2_X1  g744(.A1(new_n880), .A2(new_n943), .ZN(new_n946));
  OR2_X1    g745(.A1(new_n641), .A2(G197gat), .ZN(new_n947));
  OAI21_X1  g746(.A(new_n945), .B1(new_n946), .B2(new_n947), .ZN(G1352gat));
  NAND3_X1  g747(.A1(new_n905), .A2(KEYINPUT126), .A3(new_n943), .ZN(new_n949));
  INV_X1    g748(.A(KEYINPUT126), .ZN(new_n950));
  OAI21_X1  g749(.A(new_n950), .B1(new_n904), .B2(new_n942), .ZN(new_n951));
  NAND3_X1  g750(.A1(new_n949), .A2(G204gat), .A3(new_n951), .ZN(new_n952));
  INV_X1    g751(.A(KEYINPUT62), .ZN(new_n953));
  NAND2_X1  g752(.A1(new_n953), .A2(KEYINPUT125), .ZN(new_n954));
  NOR2_X1   g753(.A1(new_n946), .A2(G204gat), .ZN(new_n955));
  NAND2_X1  g754(.A1(new_n955), .A2(new_n661), .ZN(new_n956));
  NOR2_X1   g755(.A1(new_n953), .A2(KEYINPUT125), .ZN(new_n957));
  OAI21_X1  g756(.A(new_n954), .B1(new_n956), .B2(new_n957), .ZN(new_n958));
  NAND4_X1  g757(.A1(new_n955), .A2(KEYINPUT125), .A3(new_n953), .A4(new_n661), .ZN(new_n959));
  NAND3_X1  g758(.A1(new_n952), .A2(new_n958), .A3(new_n959), .ZN(G1353gat));
  OAI21_X1  g759(.A(G211gat), .B1(new_n944), .B2(new_n567), .ZN(new_n961));
  XOR2_X1   g760(.A(new_n961), .B(KEYINPUT63), .Z(new_n962));
  NAND4_X1  g761(.A1(new_n880), .A2(new_n351), .A3(new_n568), .A4(new_n943), .ZN(new_n963));
  NAND2_X1  g762(.A1(new_n962), .A2(new_n963), .ZN(G1354gat));
  OAI21_X1  g763(.A(G218gat), .B1(new_n944), .B2(new_n616), .ZN(new_n965));
  NAND2_X1  g764(.A1(new_n615), .A2(new_n352), .ZN(new_n966));
  OAI21_X1  g765(.A(new_n965), .B1(new_n946), .B2(new_n966), .ZN(new_n967));
  INV_X1    g766(.A(KEYINPUT127), .ZN(new_n968));
  XNOR2_X1  g767(.A(new_n967), .B(new_n968), .ZN(G1355gat));
endmodule


