//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 0 0 1 1 0 0 1 1 1 1 0 0 0 1 1 1 1 0 0 1 0 1 1 0 1 0 0 0 1 1 1 0 1 0 1 1 0 0 1 0 0 0 0 1 1 1 1 1 1 1 1 1 0 1 0 1 0 0 0 0 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:36:23 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n236, new_n237,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n244, new_n245,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n252, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n601, new_n602, new_n603, new_n604, new_n605,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1183, new_n1184, new_n1185, new_n1186, new_n1187,
    new_n1188, new_n1189, new_n1190, new_n1191, new_n1192, new_n1193,
    new_n1194, new_n1195, new_n1196, new_n1197, new_n1198, new_n1199,
    new_n1200, new_n1201, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1213,
    new_n1214, new_n1216, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1267, new_n1268, new_n1269,
    new_n1270, new_n1271, new_n1272, new_n1273, new_n1274, new_n1275;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(new_n201), .ZN(new_n202));
  NOR3_X1   g0002(.A1(new_n202), .A2(G50), .A3(G77), .ZN(G353));
  OAI21_X1  g0003(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0004(.A(G1), .ZN(new_n205));
  INV_X1    g0005(.A(G20), .ZN(new_n206));
  NOR2_X1   g0006(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  INV_X1    g0007(.A(new_n207), .ZN(new_n208));
  AOI22_X1  g0008(.A1(G77), .A2(G244), .B1(G97), .B2(G257), .ZN(new_n209));
  INV_X1    g0009(.A(G50), .ZN(new_n210));
  INV_X1    g0010(.A(G226), .ZN(new_n211));
  INV_X1    g0011(.A(G87), .ZN(new_n212));
  INV_X1    g0012(.A(G250), .ZN(new_n213));
  OAI221_X1 g0013(.A(new_n209), .B1(new_n210), .B2(new_n211), .C1(new_n212), .C2(new_n213), .ZN(new_n214));
  AOI22_X1  g0014(.A1(G107), .A2(G264), .B1(G116), .B2(G270), .ZN(new_n215));
  INV_X1    g0015(.A(G58), .ZN(new_n216));
  INV_X1    g0016(.A(G232), .ZN(new_n217));
  INV_X1    g0017(.A(G68), .ZN(new_n218));
  INV_X1    g0018(.A(G238), .ZN(new_n219));
  OAI221_X1 g0019(.A(new_n215), .B1(new_n216), .B2(new_n217), .C1(new_n218), .C2(new_n219), .ZN(new_n220));
  OAI21_X1  g0020(.A(new_n208), .B1(new_n214), .B2(new_n220), .ZN(new_n221));
  XNOR2_X1  g0021(.A(new_n221), .B(KEYINPUT67), .ZN(new_n222));
  INV_X1    g0022(.A(KEYINPUT1), .ZN(new_n223));
  NOR2_X1   g0023(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  XNOR2_X1  g0024(.A(new_n224), .B(KEYINPUT68), .ZN(new_n225));
  NOR2_X1   g0025(.A1(new_n208), .A2(G13), .ZN(new_n226));
  OAI211_X1 g0026(.A(new_n226), .B(G250), .C1(G257), .C2(G264), .ZN(new_n227));
  XNOR2_X1  g0027(.A(new_n227), .B(KEYINPUT0), .ZN(new_n228));
  XNOR2_X1  g0028(.A(KEYINPUT64), .B(G20), .ZN(new_n229));
  NAND2_X1  g0029(.A1(G1), .A2(G13), .ZN(new_n230));
  NOR2_X1   g0030(.A1(new_n229), .A2(new_n230), .ZN(new_n231));
  INV_X1    g0031(.A(new_n231), .ZN(new_n232));
  OR2_X1    g0032(.A1(new_n201), .A2(KEYINPUT65), .ZN(new_n233));
  NAND2_X1  g0033(.A1(new_n201), .A2(KEYINPUT65), .ZN(new_n234));
  NAND3_X1  g0034(.A1(new_n233), .A2(G50), .A3(new_n234), .ZN(new_n235));
  OAI21_X1  g0035(.A(new_n228), .B1(new_n232), .B2(new_n235), .ZN(new_n236));
  XOR2_X1   g0036(.A(new_n236), .B(KEYINPUT66), .Z(new_n237));
  AOI211_X1 g0037(.A(new_n225), .B(new_n237), .C1(new_n223), .C2(new_n222), .ZN(G361));
  XNOR2_X1  g0038(.A(G238), .B(G244), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n239), .B(G232), .ZN(new_n240));
  XOR2_X1   g0040(.A(KEYINPUT2), .B(G226), .Z(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XOR2_X1   g0042(.A(G250), .B(G257), .Z(new_n243));
  XNOR2_X1  g0043(.A(G264), .B(G270), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XOR2_X1   g0045(.A(new_n242), .B(new_n245), .Z(G358));
  XNOR2_X1  g0046(.A(G50), .B(G68), .ZN(new_n247));
  XNOR2_X1  g0047(.A(G58), .B(G77), .ZN(new_n248));
  XOR2_X1   g0048(.A(new_n247), .B(new_n248), .Z(new_n249));
  XOR2_X1   g0049(.A(G87), .B(G116), .Z(new_n250));
  XNOR2_X1  g0050(.A(G97), .B(G107), .ZN(new_n251));
  XNOR2_X1  g0051(.A(new_n250), .B(new_n251), .ZN(new_n252));
  XNOR2_X1  g0052(.A(new_n249), .B(new_n252), .ZN(G351));
  INV_X1    g0053(.A(KEYINPUT13), .ZN(new_n254));
  INV_X1    g0054(.A(G1698), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n255), .A2(KEYINPUT69), .ZN(new_n256));
  INV_X1    g0056(.A(KEYINPUT69), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n257), .A2(G1698), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n256), .A2(new_n258), .ZN(new_n259));
  XNOR2_X1  g0059(.A(KEYINPUT3), .B(G33), .ZN(new_n260));
  AND2_X1   g0060(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n261), .A2(G226), .ZN(new_n262));
  INV_X1    g0062(.A(G33), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n263), .A2(KEYINPUT3), .ZN(new_n264));
  INV_X1    g0064(.A(KEYINPUT3), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n265), .A2(G33), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n264), .A2(new_n266), .ZN(new_n267));
  NOR2_X1   g0067(.A1(new_n267), .A2(new_n255), .ZN(new_n268));
  INV_X1    g0068(.A(KEYINPUT71), .ZN(new_n269));
  NAND3_X1  g0069(.A1(new_n268), .A2(new_n269), .A3(G232), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n260), .A2(G1698), .ZN(new_n271));
  OAI21_X1  g0071(.A(KEYINPUT71), .B1(new_n271), .B2(new_n217), .ZN(new_n272));
  NAND2_X1  g0072(.A1(G33), .A2(G97), .ZN(new_n273));
  NAND4_X1  g0073(.A1(new_n262), .A2(new_n270), .A3(new_n272), .A4(new_n273), .ZN(new_n274));
  AOI21_X1  g0074(.A(new_n230), .B1(G33), .B2(G41), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  OAI21_X1  g0076(.A(new_n205), .B1(G41), .B2(G45), .ZN(new_n277));
  INV_X1    g0077(.A(G274), .ZN(new_n278));
  NOR2_X1   g0078(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  INV_X1    g0079(.A(new_n279), .ZN(new_n280));
  INV_X1    g0080(.A(new_n275), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n281), .A2(new_n277), .ZN(new_n282));
  OAI21_X1  g0082(.A(new_n280), .B1(new_n282), .B2(new_n219), .ZN(new_n283));
  INV_X1    g0083(.A(new_n283), .ZN(new_n284));
  AOI21_X1  g0084(.A(new_n254), .B1(new_n276), .B2(new_n284), .ZN(new_n285));
  AOI211_X1 g0085(.A(KEYINPUT13), .B(new_n283), .C1(new_n274), .C2(new_n275), .ZN(new_n286));
  OAI21_X1  g0086(.A(G169), .B1(new_n285), .B2(new_n286), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n287), .A2(KEYINPUT14), .ZN(new_n288));
  INV_X1    g0088(.A(KEYINPUT14), .ZN(new_n289));
  OAI211_X1 g0089(.A(new_n289), .B(G169), .C1(new_n285), .C2(new_n286), .ZN(new_n290));
  INV_X1    g0090(.A(G179), .ZN(new_n291));
  OR2_X1    g0091(.A1(new_n285), .A2(new_n286), .ZN(new_n292));
  OAI211_X1 g0092(.A(new_n288), .B(new_n290), .C1(new_n291), .C2(new_n292), .ZN(new_n293));
  NAND3_X1  g0093(.A1(new_n205), .A2(G13), .A3(G20), .ZN(new_n294));
  INV_X1    g0094(.A(new_n294), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n295), .A2(new_n218), .ZN(new_n296));
  AND2_X1   g0096(.A1(new_n296), .A2(KEYINPUT12), .ZN(new_n297));
  OR2_X1    g0097(.A1(new_n297), .A2(KEYINPUT72), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n297), .A2(KEYINPUT72), .ZN(new_n299));
  OAI211_X1 g0099(.A(new_n298), .B(new_n299), .C1(KEYINPUT12), .C2(new_n296), .ZN(new_n300));
  NAND3_X1  g0100(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n301), .A2(new_n230), .ZN(new_n302));
  INV_X1    g0102(.A(new_n302), .ZN(new_n303));
  OAI21_X1  g0103(.A(new_n303), .B1(G1), .B2(new_n206), .ZN(new_n304));
  OAI21_X1  g0104(.A(new_n300), .B1(new_n218), .B2(new_n304), .ZN(new_n305));
  NOR2_X1   g0105(.A1(G20), .A2(G33), .ZN(new_n306));
  AOI22_X1  g0106(.A1(new_n306), .A2(G50), .B1(G20), .B2(new_n218), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n229), .A2(G33), .ZN(new_n308));
  INV_X1    g0108(.A(G77), .ZN(new_n309));
  OAI21_X1  g0109(.A(new_n307), .B1(new_n308), .B2(new_n309), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n310), .A2(new_n302), .ZN(new_n311));
  XOR2_X1   g0111(.A(new_n311), .B(KEYINPUT11), .Z(new_n312));
  NOR2_X1   g0112(.A1(new_n305), .A2(new_n312), .ZN(new_n313));
  INV_X1    g0113(.A(new_n313), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n293), .A2(new_n314), .ZN(new_n315));
  INV_X1    g0115(.A(new_n315), .ZN(new_n316));
  OAI211_X1 g0116(.A(new_n303), .B(G77), .C1(G1), .C2(new_n206), .ZN(new_n317));
  OAI21_X1  g0117(.A(new_n317), .B1(G77), .B2(new_n294), .ZN(new_n318));
  XNOR2_X1  g0118(.A(KEYINPUT8), .B(G58), .ZN(new_n319));
  INV_X1    g0119(.A(new_n319), .ZN(new_n320));
  AND2_X1   g0120(.A1(KEYINPUT64), .A2(G20), .ZN(new_n321));
  NOR2_X1   g0121(.A1(KEYINPUT64), .A2(G20), .ZN(new_n322));
  NOR2_X1   g0122(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  AOI22_X1  g0123(.A1(new_n320), .A2(new_n306), .B1(new_n323), .B2(G77), .ZN(new_n324));
  XOR2_X1   g0124(.A(KEYINPUT15), .B(G87), .Z(new_n325));
  INV_X1    g0125(.A(new_n325), .ZN(new_n326));
  OAI21_X1  g0126(.A(new_n324), .B1(new_n308), .B2(new_n326), .ZN(new_n327));
  AOI21_X1  g0127(.A(new_n318), .B1(new_n327), .B2(new_n302), .ZN(new_n328));
  INV_X1    g0128(.A(new_n328), .ZN(new_n329));
  INV_X1    g0129(.A(G107), .ZN(new_n330));
  OAI22_X1  g0130(.A1(new_n271), .A2(new_n219), .B1(new_n330), .B2(new_n260), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n259), .A2(new_n260), .ZN(new_n332));
  NOR2_X1   g0132(.A1(new_n332), .A2(new_n217), .ZN(new_n333));
  OAI21_X1  g0133(.A(new_n275), .B1(new_n331), .B2(new_n333), .ZN(new_n334));
  INV_X1    g0134(.A(new_n282), .ZN(new_n335));
  AOI21_X1  g0135(.A(new_n279), .B1(new_n335), .B2(G244), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n334), .A2(new_n336), .ZN(new_n337));
  INV_X1    g0137(.A(new_n337), .ZN(new_n338));
  OAI21_X1  g0138(.A(new_n329), .B1(new_n338), .B2(G169), .ZN(new_n339));
  NOR2_X1   g0139(.A1(new_n337), .A2(G179), .ZN(new_n340));
  NOR2_X1   g0140(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  NOR2_X1   g0141(.A1(new_n316), .A2(new_n341), .ZN(new_n342));
  OAI21_X1  g0142(.A(G200), .B1(new_n285), .B2(new_n286), .ZN(new_n343));
  INV_X1    g0143(.A(G190), .ZN(new_n344));
  OAI211_X1 g0144(.A(new_n313), .B(new_n343), .C1(new_n292), .C2(new_n344), .ZN(new_n345));
  OAI21_X1  g0145(.A(new_n328), .B1(new_n337), .B2(new_n344), .ZN(new_n346));
  AOI21_X1  g0146(.A(new_n346), .B1(G200), .B2(new_n337), .ZN(new_n347));
  OAI21_X1  g0147(.A(G20), .B1(new_n202), .B2(G50), .ZN(new_n348));
  INV_X1    g0148(.A(G150), .ZN(new_n349));
  INV_X1    g0149(.A(new_n306), .ZN(new_n350));
  OAI221_X1 g0150(.A(new_n348), .B1(new_n349), .B2(new_n350), .C1(new_n308), .C2(new_n319), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n351), .A2(new_n302), .ZN(new_n352));
  MUX2_X1   g0152(.A(new_n294), .B(new_n304), .S(G50), .Z(new_n353));
  NAND2_X1  g0153(.A1(new_n352), .A2(new_n353), .ZN(new_n354));
  XNOR2_X1  g0154(.A(new_n354), .B(KEYINPUT9), .ZN(new_n355));
  INV_X1    g0155(.A(G200), .ZN(new_n356));
  OAI21_X1  g0156(.A(new_n280), .B1(new_n282), .B2(new_n211), .ZN(new_n357));
  AOI22_X1  g0157(.A1(new_n268), .A2(G223), .B1(G77), .B2(new_n267), .ZN(new_n358));
  INV_X1    g0158(.A(G222), .ZN(new_n359));
  OAI21_X1  g0159(.A(new_n358), .B1(new_n359), .B2(new_n332), .ZN(new_n360));
  AOI21_X1  g0160(.A(new_n357), .B1(new_n360), .B2(new_n275), .ZN(new_n361));
  OAI21_X1  g0161(.A(new_n355), .B1(new_n356), .B2(new_n361), .ZN(new_n362));
  AND2_X1   g0162(.A1(new_n361), .A2(G190), .ZN(new_n363));
  OR3_X1    g0163(.A1(new_n362), .A2(KEYINPUT10), .A3(new_n363), .ZN(new_n364));
  OAI21_X1  g0164(.A(KEYINPUT10), .B1(new_n362), .B2(new_n363), .ZN(new_n365));
  AOI21_X1  g0165(.A(new_n347), .B1(new_n364), .B2(new_n365), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n361), .A2(new_n291), .ZN(new_n367));
  OAI211_X1 g0167(.A(new_n367), .B(new_n354), .C1(G169), .C2(new_n361), .ZN(new_n368));
  XOR2_X1   g0168(.A(new_n368), .B(KEYINPUT70), .Z(new_n369));
  NAND4_X1  g0169(.A1(new_n342), .A2(new_n345), .A3(new_n366), .A4(new_n369), .ZN(new_n370));
  NOR2_X1   g0170(.A1(new_n320), .A2(new_n295), .ZN(new_n371));
  AOI21_X1  g0171(.A(new_n371), .B1(new_n304), .B2(new_n320), .ZN(new_n372));
  INV_X1    g0172(.A(new_n372), .ZN(new_n373));
  NOR2_X1   g0173(.A1(new_n216), .A2(new_n218), .ZN(new_n374));
  OAI21_X1  g0174(.A(G20), .B1(new_n374), .B2(new_n201), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n306), .A2(G159), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n375), .A2(new_n376), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n267), .A2(new_n206), .ZN(new_n378));
  AOI21_X1  g0178(.A(new_n218), .B1(new_n378), .B2(KEYINPUT7), .ZN(new_n379));
  INV_X1    g0179(.A(KEYINPUT7), .ZN(new_n380));
  NAND3_X1  g0180(.A1(new_n267), .A2(new_n229), .A3(new_n380), .ZN(new_n381));
  AOI21_X1  g0181(.A(new_n377), .B1(new_n379), .B2(new_n381), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n382), .A2(KEYINPUT16), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n383), .A2(new_n302), .ZN(new_n384));
  NOR2_X1   g0184(.A1(new_n323), .A2(new_n380), .ZN(new_n385));
  INV_X1    g0185(.A(KEYINPUT73), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n264), .A2(new_n386), .ZN(new_n387));
  NAND3_X1  g0187(.A1(new_n263), .A2(KEYINPUT73), .A3(KEYINPUT3), .ZN(new_n388));
  NAND3_X1  g0188(.A1(new_n387), .A2(new_n266), .A3(new_n388), .ZN(new_n389));
  AND2_X1   g0189(.A1(new_n385), .A2(new_n389), .ZN(new_n390));
  AOI21_X1  g0190(.A(KEYINPUT7), .B1(new_n267), .B2(new_n206), .ZN(new_n391));
  OAI21_X1  g0191(.A(G68), .B1(new_n390), .B2(new_n391), .ZN(new_n392));
  INV_X1    g0192(.A(new_n377), .ZN(new_n393));
  AOI21_X1  g0193(.A(KEYINPUT16), .B1(new_n392), .B2(new_n393), .ZN(new_n394));
  OAI21_X1  g0194(.A(new_n373), .B1(new_n384), .B2(new_n394), .ZN(new_n395));
  INV_X1    g0195(.A(KEYINPUT76), .ZN(new_n396));
  OAI21_X1  g0196(.A(new_n280), .B1(new_n282), .B2(new_n217), .ZN(new_n397));
  NAND3_X1  g0197(.A1(new_n259), .A2(new_n260), .A3(G223), .ZN(new_n398));
  NAND3_X1  g0198(.A1(new_n260), .A2(G226), .A3(G1698), .ZN(new_n399));
  NAND2_X1  g0199(.A1(G33), .A2(G87), .ZN(new_n400));
  NAND3_X1  g0200(.A1(new_n398), .A2(new_n399), .A3(new_n400), .ZN(new_n401));
  INV_X1    g0201(.A(KEYINPUT74), .ZN(new_n402));
  AOI21_X1  g0202(.A(new_n281), .B1(new_n401), .B2(new_n402), .ZN(new_n403));
  NAND4_X1  g0203(.A1(new_n398), .A2(new_n399), .A3(KEYINPUT74), .A4(new_n400), .ZN(new_n404));
  AOI211_X1 g0204(.A(G190), .B(new_n397), .C1(new_n403), .C2(new_n404), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n401), .A2(new_n402), .ZN(new_n406));
  NAND3_X1  g0206(.A1(new_n406), .A2(new_n404), .A3(new_n275), .ZN(new_n407));
  INV_X1    g0207(.A(new_n397), .ZN(new_n408));
  AOI21_X1  g0208(.A(G200), .B1(new_n407), .B2(new_n408), .ZN(new_n409));
  OAI21_X1  g0209(.A(new_n396), .B1(new_n405), .B2(new_n409), .ZN(new_n410));
  NAND3_X1  g0210(.A1(new_n407), .A2(new_n344), .A3(new_n408), .ZN(new_n411));
  AOI21_X1  g0211(.A(new_n397), .B1(new_n403), .B2(new_n404), .ZN(new_n412));
  OAI211_X1 g0212(.A(new_n411), .B(KEYINPUT76), .C1(G200), .C2(new_n412), .ZN(new_n413));
  AOI21_X1  g0213(.A(new_n395), .B1(new_n410), .B2(new_n413), .ZN(new_n414));
  INV_X1    g0214(.A(KEYINPUT17), .ZN(new_n415));
  XNOR2_X1  g0215(.A(new_n414), .B(new_n415), .ZN(new_n416));
  AOI211_X1 g0216(.A(G179), .B(new_n397), .C1(new_n403), .C2(new_n404), .ZN(new_n417));
  AOI21_X1  g0217(.A(G169), .B1(new_n407), .B2(new_n408), .ZN(new_n418));
  OAI21_X1  g0218(.A(KEYINPUT75), .B1(new_n417), .B2(new_n418), .ZN(new_n419));
  NAND3_X1  g0219(.A1(new_n407), .A2(new_n291), .A3(new_n408), .ZN(new_n420));
  INV_X1    g0220(.A(KEYINPUT75), .ZN(new_n421));
  OAI211_X1 g0221(.A(new_n420), .B(new_n421), .C1(G169), .C2(new_n412), .ZN(new_n422));
  NAND3_X1  g0222(.A1(new_n419), .A2(new_n395), .A3(new_n422), .ZN(new_n423));
  INV_X1    g0223(.A(KEYINPUT18), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n423), .A2(new_n424), .ZN(new_n425));
  NAND4_X1  g0225(.A1(new_n419), .A2(KEYINPUT18), .A3(new_n422), .A4(new_n395), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n425), .A2(new_n426), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n416), .A2(new_n427), .ZN(new_n428));
  INV_X1    g0228(.A(G45), .ZN(new_n429));
  NOR2_X1   g0229(.A1(new_n429), .A2(G1), .ZN(new_n430));
  INV_X1    g0230(.A(new_n430), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n431), .A2(G250), .ZN(new_n432));
  OAI22_X1  g0232(.A1(new_n432), .A2(new_n275), .B1(new_n278), .B2(new_n431), .ZN(new_n433));
  INV_X1    g0233(.A(KEYINPUT79), .ZN(new_n434));
  OAI21_X1  g0234(.A(new_n434), .B1(new_n332), .B2(new_n219), .ZN(new_n435));
  NAND4_X1  g0235(.A1(new_n259), .A2(new_n260), .A3(KEYINPUT79), .A4(G238), .ZN(new_n436));
  NAND4_X1  g0236(.A1(new_n264), .A2(new_n266), .A3(G244), .A4(G1698), .ZN(new_n437));
  NAND2_X1  g0237(.A1(G33), .A2(G116), .ZN(new_n438));
  AND2_X1   g0238(.A1(new_n437), .A2(new_n438), .ZN(new_n439));
  NAND3_X1  g0239(.A1(new_n435), .A2(new_n436), .A3(new_n439), .ZN(new_n440));
  AOI21_X1  g0240(.A(new_n433), .B1(new_n440), .B2(new_n275), .ZN(new_n441));
  INV_X1    g0241(.A(new_n441), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n442), .A2(G200), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n440), .A2(new_n275), .ZN(new_n444));
  INV_X1    g0244(.A(new_n433), .ZN(new_n445));
  NAND3_X1  g0245(.A1(new_n444), .A2(G190), .A3(new_n445), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n446), .A2(KEYINPUT83), .ZN(new_n447));
  NOR2_X1   g0247(.A1(new_n325), .A2(new_n294), .ZN(new_n448));
  OAI211_X1 g0248(.A(new_n303), .B(new_n294), .C1(G1), .C2(new_n263), .ZN(new_n449));
  NOR2_X1   g0249(.A1(new_n449), .A2(new_n212), .ZN(new_n450));
  OAI211_X1 g0250(.A(G33), .B(G97), .C1(new_n321), .C2(new_n322), .ZN(new_n451));
  INV_X1    g0251(.A(KEYINPUT19), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n451), .A2(new_n452), .ZN(new_n453));
  INV_X1    g0253(.A(G97), .ZN(new_n454));
  NAND3_X1  g0254(.A1(new_n212), .A2(new_n454), .A3(new_n330), .ZN(new_n455));
  NOR2_X1   g0255(.A1(new_n273), .A2(new_n452), .ZN(new_n456));
  OAI21_X1  g0256(.A(new_n455), .B1(new_n323), .B2(new_n456), .ZN(new_n457));
  NAND3_X1  g0257(.A1(new_n229), .A2(new_n260), .A3(G68), .ZN(new_n458));
  NAND3_X1  g0258(.A1(new_n453), .A2(new_n457), .A3(new_n458), .ZN(new_n459));
  INV_X1    g0259(.A(KEYINPUT82), .ZN(new_n460));
  AOI21_X1  g0260(.A(new_n303), .B1(new_n459), .B2(new_n460), .ZN(new_n461));
  NAND4_X1  g0261(.A1(new_n453), .A2(new_n457), .A3(new_n458), .A4(KEYINPUT82), .ZN(new_n462));
  AOI211_X1 g0262(.A(new_n448), .B(new_n450), .C1(new_n461), .C2(new_n462), .ZN(new_n463));
  INV_X1    g0263(.A(KEYINPUT83), .ZN(new_n464));
  NAND3_X1  g0264(.A1(new_n441), .A2(new_n464), .A3(G190), .ZN(new_n465));
  AND4_X1   g0265(.A1(new_n443), .A2(new_n447), .A3(new_n463), .A4(new_n465), .ZN(new_n466));
  AOI21_X1  g0266(.A(new_n448), .B1(new_n461), .B2(new_n462), .ZN(new_n467));
  INV_X1    g0267(.A(new_n449), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n468), .A2(new_n325), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n467), .A2(new_n469), .ZN(new_n470));
  INV_X1    g0270(.A(new_n470), .ZN(new_n471));
  INV_X1    g0271(.A(KEYINPUT80), .ZN(new_n472));
  NAND3_X1  g0272(.A1(new_n441), .A2(new_n472), .A3(new_n291), .ZN(new_n473));
  OAI21_X1  g0273(.A(KEYINPUT80), .B1(new_n441), .B2(G169), .ZN(new_n474));
  AOI211_X1 g0274(.A(G179), .B(new_n433), .C1(new_n440), .C2(new_n275), .ZN(new_n475));
  OAI21_X1  g0275(.A(new_n473), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  INV_X1    g0276(.A(KEYINPUT81), .ZN(new_n477));
  AOI21_X1  g0277(.A(new_n471), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  OAI211_X1 g0278(.A(KEYINPUT81), .B(new_n473), .C1(new_n474), .C2(new_n475), .ZN(new_n479));
  AOI21_X1  g0279(.A(new_n466), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n263), .A2(G97), .ZN(new_n481));
  INV_X1    g0281(.A(G283), .ZN(new_n482));
  OAI221_X1 g0282(.A(new_n481), .B1(new_n263), .B2(new_n482), .C1(new_n321), .C2(new_n322), .ZN(new_n483));
  INV_X1    g0283(.A(G116), .ZN(new_n484));
  AOI22_X1  g0284(.A1(new_n301), .A2(new_n230), .B1(G20), .B2(new_n484), .ZN(new_n485));
  NAND3_X1  g0285(.A1(new_n483), .A2(KEYINPUT20), .A3(new_n485), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n486), .A2(KEYINPUT84), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n483), .A2(new_n485), .ZN(new_n488));
  INV_X1    g0288(.A(KEYINPUT20), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  INV_X1    g0290(.A(KEYINPUT84), .ZN(new_n491));
  NAND4_X1  g0291(.A1(new_n483), .A2(new_n491), .A3(KEYINPUT20), .A4(new_n485), .ZN(new_n492));
  NAND3_X1  g0292(.A1(new_n487), .A2(new_n490), .A3(new_n492), .ZN(new_n493));
  NOR2_X1   g0293(.A1(new_n294), .A2(G116), .ZN(new_n494));
  AOI21_X1  g0294(.A(new_n494), .B1(new_n468), .B2(G116), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n493), .A2(new_n495), .ZN(new_n496));
  INV_X1    g0296(.A(G264), .ZN(new_n497));
  INV_X1    g0297(.A(G303), .ZN(new_n498));
  OAI22_X1  g0298(.A1(new_n271), .A2(new_n497), .B1(new_n498), .B2(new_n260), .ZN(new_n499));
  INV_X1    g0299(.A(G257), .ZN(new_n500));
  NOR2_X1   g0300(.A1(new_n332), .A2(new_n500), .ZN(new_n501));
  OAI21_X1  g0301(.A(new_n275), .B1(new_n499), .B2(new_n501), .ZN(new_n502));
  INV_X1    g0302(.A(G41), .ZN(new_n503));
  OAI211_X1 g0303(.A(new_n205), .B(G45), .C1(new_n503), .C2(KEYINPUT5), .ZN(new_n504));
  INV_X1    g0304(.A(KEYINPUT78), .ZN(new_n505));
  AOI22_X1  g0305(.A1(new_n504), .A2(new_n505), .B1(KEYINPUT5), .B2(new_n503), .ZN(new_n506));
  OAI211_X1 g0306(.A(new_n430), .B(KEYINPUT78), .C1(KEYINPUT5), .C2(new_n503), .ZN(new_n507));
  NAND4_X1  g0307(.A1(new_n506), .A2(G274), .A3(new_n281), .A4(new_n507), .ZN(new_n508));
  AOI21_X1  g0308(.A(new_n275), .B1(new_n506), .B2(new_n507), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n509), .A2(G270), .ZN(new_n510));
  NAND3_X1  g0310(.A1(new_n502), .A2(new_n508), .A3(new_n510), .ZN(new_n511));
  NAND3_X1  g0311(.A1(new_n496), .A2(G169), .A3(new_n511), .ZN(new_n512));
  INV_X1    g0312(.A(KEYINPUT21), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  NAND4_X1  g0314(.A1(new_n496), .A2(KEYINPUT21), .A3(new_n511), .A4(G169), .ZN(new_n515));
  INV_X1    g0315(.A(new_n511), .ZN(new_n516));
  NAND3_X1  g0316(.A1(new_n516), .A2(new_n496), .A3(G179), .ZN(new_n517));
  NAND3_X1  g0317(.A1(new_n514), .A2(new_n515), .A3(new_n517), .ZN(new_n518));
  NOR2_X1   g0318(.A1(new_n294), .A2(G107), .ZN(new_n519));
  INV_X1    g0319(.A(KEYINPUT25), .ZN(new_n520));
  XNOR2_X1  g0320(.A(new_n519), .B(new_n520), .ZN(new_n521));
  AOI21_X1  g0321(.A(new_n521), .B1(new_n468), .B2(G107), .ZN(new_n522));
  NAND3_X1  g0322(.A1(new_n229), .A2(new_n260), .A3(G87), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n523), .A2(KEYINPUT22), .ZN(new_n524));
  INV_X1    g0324(.A(KEYINPUT22), .ZN(new_n525));
  NAND4_X1  g0325(.A1(new_n229), .A2(new_n260), .A3(new_n525), .A4(G87), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n524), .A2(new_n526), .ZN(new_n527));
  INV_X1    g0327(.A(KEYINPUT23), .ZN(new_n528));
  NAND3_X1  g0328(.A1(new_n323), .A2(new_n528), .A3(new_n330), .ZN(new_n529));
  AOI21_X1  g0329(.A(new_n528), .B1(G20), .B2(new_n330), .ZN(new_n530));
  NOR2_X1   g0330(.A1(new_n438), .A2(G20), .ZN(new_n531));
  NOR2_X1   g0331(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  NAND3_X1  g0332(.A1(new_n527), .A2(new_n529), .A3(new_n532), .ZN(new_n533));
  INV_X1    g0333(.A(KEYINPUT24), .ZN(new_n534));
  NOR2_X1   g0334(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n529), .A2(new_n532), .ZN(new_n536));
  AOI21_X1  g0336(.A(new_n536), .B1(new_n524), .B2(new_n526), .ZN(new_n537));
  OAI21_X1  g0337(.A(new_n302), .B1(new_n537), .B2(KEYINPUT24), .ZN(new_n538));
  OAI21_X1  g0338(.A(new_n522), .B1(new_n535), .B2(new_n538), .ZN(new_n539));
  INV_X1    g0339(.A(G294), .ZN(new_n540));
  OAI22_X1  g0340(.A1(new_n271), .A2(new_n500), .B1(new_n263), .B2(new_n540), .ZN(new_n541));
  NOR2_X1   g0341(.A1(new_n332), .A2(new_n213), .ZN(new_n542));
  OAI21_X1  g0342(.A(new_n275), .B1(new_n541), .B2(new_n542), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n509), .A2(G264), .ZN(new_n544));
  NAND3_X1  g0344(.A1(new_n543), .A2(new_n508), .A3(new_n544), .ZN(new_n545));
  INV_X1    g0345(.A(G169), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  AND2_X1   g0347(.A1(new_n543), .A2(new_n544), .ZN(new_n548));
  NAND3_X1  g0348(.A1(new_n548), .A2(new_n291), .A3(new_n508), .ZN(new_n549));
  AND3_X1   g0349(.A1(new_n539), .A2(new_n547), .A3(new_n549), .ZN(new_n550));
  NOR2_X1   g0350(.A1(new_n518), .A2(new_n550), .ZN(new_n551));
  AOI21_X1  g0351(.A(new_n496), .B1(new_n516), .B2(G190), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n511), .A2(G200), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  NAND3_X1  g0354(.A1(new_n330), .A2(KEYINPUT6), .A3(G97), .ZN(new_n555));
  INV_X1    g0355(.A(new_n251), .ZN(new_n556));
  OAI21_X1  g0356(.A(new_n555), .B1(new_n556), .B2(KEYINPUT6), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n557), .A2(new_n323), .ZN(new_n558));
  OAI21_X1  g0358(.A(new_n558), .B1(new_n309), .B2(new_n350), .ZN(new_n559));
  AOI22_X1  g0359(.A1(new_n389), .A2(new_n385), .B1(new_n378), .B2(new_n380), .ZN(new_n560));
  NOR2_X1   g0360(.A1(new_n560), .A2(new_n330), .ZN(new_n561));
  OAI21_X1  g0361(.A(new_n302), .B1(new_n559), .B2(new_n561), .ZN(new_n562));
  NOR2_X1   g0362(.A1(new_n294), .A2(G97), .ZN(new_n563));
  AOI21_X1  g0363(.A(new_n563), .B1(new_n468), .B2(G97), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n562), .A2(new_n564), .ZN(new_n565));
  NAND3_X1  g0365(.A1(new_n260), .A2(G250), .A3(G1698), .ZN(new_n566));
  INV_X1    g0366(.A(KEYINPUT4), .ZN(new_n567));
  AOI22_X1  g0367(.A1(new_n567), .A2(KEYINPUT77), .B1(G33), .B2(G283), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n566), .A2(new_n568), .ZN(new_n569));
  NOR2_X1   g0369(.A1(new_n567), .A2(KEYINPUT77), .ZN(new_n570));
  INV_X1    g0370(.A(G244), .ZN(new_n571));
  NOR2_X1   g0371(.A1(new_n332), .A2(new_n571), .ZN(new_n572));
  AOI21_X1  g0372(.A(new_n569), .B1(new_n570), .B2(new_n572), .ZN(new_n573));
  OAI22_X1  g0373(.A1(new_n332), .A2(new_n571), .B1(KEYINPUT77), .B2(new_n567), .ZN(new_n574));
  AOI21_X1  g0374(.A(new_n281), .B1(new_n573), .B2(new_n574), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n509), .A2(G257), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n576), .A2(new_n508), .ZN(new_n577));
  OAI21_X1  g0377(.A(new_n546), .B1(new_n575), .B2(new_n577), .ZN(new_n578));
  NAND3_X1  g0378(.A1(new_n261), .A2(G244), .A3(new_n570), .ZN(new_n579));
  NAND3_X1  g0379(.A1(new_n579), .A2(new_n566), .A3(new_n568), .ZN(new_n580));
  INV_X1    g0380(.A(new_n574), .ZN(new_n581));
  OAI21_X1  g0381(.A(new_n275), .B1(new_n580), .B2(new_n581), .ZN(new_n582));
  INV_X1    g0382(.A(new_n577), .ZN(new_n583));
  NAND3_X1  g0383(.A1(new_n582), .A2(new_n583), .A3(new_n291), .ZN(new_n584));
  NAND3_X1  g0384(.A1(new_n565), .A2(new_n578), .A3(new_n584), .ZN(new_n585));
  OAI21_X1  g0385(.A(G200), .B1(new_n575), .B2(new_n577), .ZN(new_n586));
  NAND3_X1  g0386(.A1(new_n582), .A2(new_n583), .A3(G190), .ZN(new_n587));
  INV_X1    g0387(.A(new_n564), .ZN(new_n588));
  OAI221_X1 g0388(.A(new_n558), .B1(new_n309), .B2(new_n350), .C1(new_n560), .C2(new_n330), .ZN(new_n589));
  AOI21_X1  g0389(.A(new_n588), .B1(new_n589), .B2(new_n302), .ZN(new_n590));
  NAND3_X1  g0390(.A1(new_n586), .A2(new_n587), .A3(new_n590), .ZN(new_n591));
  NAND3_X1  g0391(.A1(new_n554), .A2(new_n585), .A3(new_n591), .ZN(new_n592));
  INV_X1    g0392(.A(KEYINPUT85), .ZN(new_n593));
  NAND4_X1  g0393(.A1(new_n543), .A2(new_n544), .A3(new_n344), .A4(new_n508), .ZN(new_n594));
  AOI22_X1  g0394(.A1(new_n593), .A2(new_n594), .B1(new_n545), .B2(new_n356), .ZN(new_n595));
  OR2_X1    g0395(.A1(new_n594), .A2(new_n593), .ZN(new_n596));
  AOI21_X1  g0396(.A(new_n539), .B1(new_n595), .B2(new_n596), .ZN(new_n597));
  NOR2_X1   g0397(.A1(new_n592), .A2(new_n597), .ZN(new_n598));
  NAND3_X1  g0398(.A1(new_n480), .A2(new_n551), .A3(new_n598), .ZN(new_n599));
  NOR3_X1   g0399(.A1(new_n370), .A2(new_n428), .A3(new_n599), .ZN(G372));
  NOR2_X1   g0400(.A1(new_n370), .A2(new_n428), .ZN(new_n601));
  INV_X1    g0401(.A(KEYINPUT26), .ZN(new_n602));
  INV_X1    g0402(.A(new_n585), .ZN(new_n603));
  AOI21_X1  g0403(.A(new_n602), .B1(new_n480), .B2(new_n603), .ZN(new_n604));
  OAI21_X1  g0404(.A(KEYINPUT86), .B1(new_n518), .B2(new_n550), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n442), .A2(new_n546), .ZN(new_n606));
  INV_X1    g0406(.A(new_n475), .ZN(new_n607));
  NAND3_X1  g0407(.A1(new_n606), .A2(new_n607), .A3(new_n470), .ZN(new_n608));
  NAND3_X1  g0408(.A1(new_n443), .A2(new_n463), .A3(new_n446), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  NOR2_X1   g0410(.A1(new_n610), .A2(new_n597), .ZN(new_n611));
  AND2_X1   g0411(.A1(new_n517), .A2(new_n515), .ZN(new_n612));
  NAND3_X1  g0412(.A1(new_n539), .A2(new_n547), .A3(new_n549), .ZN(new_n613));
  INV_X1    g0413(.A(KEYINPUT86), .ZN(new_n614));
  NAND4_X1  g0414(.A1(new_n612), .A2(new_n613), .A3(new_n614), .A4(new_n514), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n585), .A2(new_n591), .ZN(new_n616));
  INV_X1    g0416(.A(new_n616), .ZN(new_n617));
  NAND4_X1  g0417(.A1(new_n605), .A2(new_n611), .A3(new_n615), .A4(new_n617), .ZN(new_n618));
  INV_X1    g0418(.A(new_n608), .ZN(new_n619));
  NOR2_X1   g0419(.A1(new_n610), .A2(new_n585), .ZN(new_n620));
  AOI21_X1  g0420(.A(new_n619), .B1(new_n620), .B2(new_n602), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n618), .A2(new_n621), .ZN(new_n622));
  OAI21_X1  g0422(.A(new_n601), .B1(new_n604), .B2(new_n622), .ZN(new_n623));
  INV_X1    g0423(.A(new_n369), .ZN(new_n624));
  AND3_X1   g0424(.A1(new_n425), .A2(KEYINPUT87), .A3(new_n426), .ZN(new_n625));
  AOI21_X1  g0425(.A(KEYINPUT87), .B1(new_n425), .B2(new_n426), .ZN(new_n626));
  NOR2_X1   g0426(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n416), .A2(new_n345), .ZN(new_n628));
  OAI21_X1  g0428(.A(new_n627), .B1(new_n342), .B2(new_n628), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n364), .A2(new_n365), .ZN(new_n630));
  AOI21_X1  g0430(.A(new_n624), .B1(new_n629), .B2(new_n630), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n623), .A2(new_n631), .ZN(G369));
  NAND3_X1  g0432(.A1(new_n229), .A2(new_n205), .A3(G13), .ZN(new_n633));
  AND2_X1   g0433(.A1(new_n633), .A2(KEYINPUT27), .ZN(new_n634));
  NOR2_X1   g0434(.A1(new_n633), .A2(KEYINPUT27), .ZN(new_n635));
  INV_X1    g0435(.A(G213), .ZN(new_n636));
  NOR3_X1   g0436(.A1(new_n634), .A2(new_n635), .A3(new_n636), .ZN(new_n637));
  XNOR2_X1  g0437(.A(KEYINPUT88), .B(G343), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  INV_X1    g0439(.A(new_n639), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n640), .A2(new_n496), .ZN(new_n641));
  OR2_X1    g0441(.A1(new_n518), .A2(new_n641), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n518), .A2(new_n641), .ZN(new_n643));
  NAND3_X1  g0443(.A1(new_n642), .A2(new_n554), .A3(new_n643), .ZN(new_n644));
  INV_X1    g0444(.A(KEYINPUT89), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  NAND4_X1  g0446(.A1(new_n642), .A2(KEYINPUT89), .A3(new_n554), .A4(new_n643), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n595), .A2(new_n596), .ZN(new_n648));
  OR2_X1    g0448(.A1(new_n535), .A2(new_n538), .ZN(new_n649));
  NAND3_X1  g0449(.A1(new_n648), .A2(new_n649), .A3(new_n522), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n539), .A2(new_n640), .ZN(new_n651));
  AOI21_X1  g0451(.A(new_n550), .B1(new_n650), .B2(new_n651), .ZN(new_n652));
  NOR2_X1   g0452(.A1(new_n613), .A2(new_n640), .ZN(new_n653));
  NOR2_X1   g0453(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  NAND4_X1  g0454(.A1(new_n646), .A2(G330), .A3(new_n647), .A4(new_n654), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n518), .A2(new_n639), .ZN(new_n656));
  INV_X1    g0456(.A(new_n656), .ZN(new_n657));
  INV_X1    g0457(.A(new_n651), .ZN(new_n658));
  OAI21_X1  g0458(.A(new_n613), .B1(new_n597), .B2(new_n658), .ZN(new_n659));
  AOI21_X1  g0459(.A(new_n653), .B1(new_n657), .B2(new_n659), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n655), .A2(new_n660), .ZN(G399));
  INV_X1    g0461(.A(new_n226), .ZN(new_n662));
  NOR2_X1   g0462(.A1(new_n662), .A2(G41), .ZN(new_n663));
  INV_X1    g0463(.A(new_n663), .ZN(new_n664));
  NOR2_X1   g0464(.A1(new_n455), .A2(G116), .ZN(new_n665));
  NAND3_X1  g0465(.A1(new_n664), .A2(G1), .A3(new_n665), .ZN(new_n666));
  OAI21_X1  g0466(.A(new_n666), .B1(new_n235), .B2(new_n664), .ZN(new_n667));
  XNOR2_X1  g0467(.A(new_n667), .B(KEYINPUT28), .ZN(new_n668));
  INV_X1    g0468(.A(KEYINPUT31), .ZN(new_n669));
  NAND4_X1  g0469(.A1(new_n548), .A2(new_n582), .A3(new_n583), .A4(new_n441), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n516), .A2(G179), .ZN(new_n671));
  OAI21_X1  g0471(.A(KEYINPUT90), .B1(new_n670), .B2(new_n671), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n672), .A2(KEYINPUT30), .ZN(new_n673));
  INV_X1    g0473(.A(KEYINPUT30), .ZN(new_n674));
  OAI211_X1 g0474(.A(KEYINPUT90), .B(new_n674), .C1(new_n670), .C2(new_n671), .ZN(new_n675));
  NOR2_X1   g0475(.A1(new_n516), .A2(G179), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n582), .A2(new_n583), .ZN(new_n677));
  NAND4_X1  g0477(.A1(new_n676), .A2(new_n442), .A3(new_n545), .A4(new_n677), .ZN(new_n678));
  NAND3_X1  g0478(.A1(new_n673), .A2(new_n675), .A3(new_n678), .ZN(new_n679));
  AOI21_X1  g0479(.A(new_n669), .B1(new_n679), .B2(new_n640), .ZN(new_n680));
  OAI21_X1  g0480(.A(new_n680), .B1(new_n599), .B2(new_n640), .ZN(new_n681));
  NAND3_X1  g0481(.A1(new_n679), .A2(new_n669), .A3(new_n640), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  INV_X1    g0483(.A(new_n683), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n684), .A2(G330), .ZN(new_n685));
  INV_X1    g0485(.A(new_n685), .ZN(new_n686));
  NOR3_X1   g0486(.A1(new_n551), .A2(new_n597), .A3(new_n610), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n616), .A2(KEYINPUT92), .ZN(new_n688));
  INV_X1    g0488(.A(KEYINPUT92), .ZN(new_n689));
  NAND3_X1  g0489(.A1(new_n585), .A2(new_n591), .A3(new_n689), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n688), .A2(new_n690), .ZN(new_n691));
  AOI21_X1  g0491(.A(new_n619), .B1(new_n687), .B2(new_n691), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n620), .A2(KEYINPUT26), .ZN(new_n693));
  AOI21_X1  g0493(.A(KEYINPUT26), .B1(new_n480), .B2(new_n603), .ZN(new_n694));
  INV_X1    g0494(.A(KEYINPUT91), .ZN(new_n695));
  OAI21_X1  g0495(.A(new_n693), .B1(new_n694), .B2(new_n695), .ZN(new_n696));
  AOI211_X1 g0496(.A(new_n585), .B(new_n466), .C1(new_n478), .C2(new_n479), .ZN(new_n697));
  NOR3_X1   g0497(.A1(new_n697), .A2(KEYINPUT91), .A3(KEYINPUT26), .ZN(new_n698));
  OAI21_X1  g0498(.A(new_n692), .B1(new_n696), .B2(new_n698), .ZN(new_n699));
  NAND3_X1  g0499(.A1(new_n699), .A2(KEYINPUT29), .A3(new_n639), .ZN(new_n700));
  OAI21_X1  g0500(.A(new_n639), .B1(new_n622), .B2(new_n604), .ZN(new_n701));
  INV_X1    g0501(.A(KEYINPUT29), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  INV_X1    g0503(.A(KEYINPUT93), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n700), .A2(new_n705), .ZN(new_n706));
  NAND4_X1  g0506(.A1(new_n699), .A2(new_n704), .A3(KEYINPUT29), .A4(new_n639), .ZN(new_n707));
  AOI21_X1  g0507(.A(new_n686), .B1(new_n706), .B2(new_n707), .ZN(new_n708));
  OAI21_X1  g0508(.A(new_n668), .B1(new_n708), .B2(G1), .ZN(G364));
  NOR2_X1   g0509(.A1(G13), .A2(G33), .ZN(new_n710));
  INV_X1    g0510(.A(new_n710), .ZN(new_n711));
  NOR2_X1   g0511(.A1(new_n711), .A2(G20), .ZN(new_n712));
  XNOR2_X1  g0512(.A(new_n712), .B(KEYINPUT100), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n644), .A2(new_n713), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n229), .A2(G13), .ZN(new_n715));
  XOR2_X1   g0515(.A(new_n715), .B(KEYINPUT94), .Z(new_n716));
  NAND2_X1  g0516(.A1(new_n716), .A2(G45), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n717), .A2(G1), .ZN(new_n718));
  NOR2_X1   g0518(.A1(new_n718), .A2(new_n663), .ZN(new_n719));
  INV_X1    g0519(.A(new_n719), .ZN(new_n720));
  NAND3_X1  g0520(.A1(new_n226), .A2(G355), .A3(new_n260), .ZN(new_n721));
  NOR2_X1   g0521(.A1(new_n662), .A2(new_n260), .ZN(new_n722));
  NOR2_X1   g0522(.A1(new_n249), .A2(new_n429), .ZN(new_n723));
  OAI221_X1 g0523(.A(new_n722), .B1(G45), .B2(new_n235), .C1(new_n723), .C2(KEYINPUT95), .ZN(new_n724));
  AND2_X1   g0524(.A1(new_n723), .A2(KEYINPUT95), .ZN(new_n725));
  OAI221_X1 g0525(.A(new_n721), .B1(G116), .B2(new_n226), .C1(new_n724), .C2(new_n725), .ZN(new_n726));
  AOI21_X1  g0526(.A(new_n230), .B1(G20), .B2(new_n546), .ZN(new_n727));
  NOR2_X1   g0527(.A1(new_n712), .A2(new_n727), .ZN(new_n728));
  AOI21_X1  g0528(.A(new_n720), .B1(new_n726), .B2(new_n728), .ZN(new_n729));
  NOR2_X1   g0529(.A1(new_n229), .A2(new_n291), .ZN(new_n730));
  INV_X1    g0530(.A(new_n730), .ZN(new_n731));
  NOR3_X1   g0531(.A1(new_n731), .A2(G190), .A3(new_n356), .ZN(new_n732));
  INV_X1    g0532(.A(new_n732), .ZN(new_n733));
  NOR2_X1   g0533(.A1(new_n344), .A2(new_n356), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n730), .A2(new_n734), .ZN(new_n735));
  OAI22_X1  g0535(.A1(new_n733), .A2(new_n218), .B1(new_n210), .B2(new_n735), .ZN(new_n736));
  NOR2_X1   g0536(.A1(new_n344), .A2(G200), .ZN(new_n737));
  NAND2_X1  g0537(.A1(new_n737), .A2(new_n291), .ZN(new_n738));
  NAND2_X1  g0538(.A1(new_n738), .A2(new_n323), .ZN(new_n739));
  OR2_X1    g0539(.A1(new_n739), .A2(KEYINPUT99), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n739), .A2(KEYINPUT99), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  INV_X1    g0542(.A(new_n742), .ZN(new_n743));
  AOI21_X1  g0543(.A(new_n736), .B1(G97), .B2(new_n743), .ZN(new_n744));
  OR2_X1    g0544(.A1(new_n731), .A2(KEYINPUT96), .ZN(new_n745));
  NAND2_X1  g0545(.A1(new_n731), .A2(KEYINPUT96), .ZN(new_n746));
  NAND3_X1  g0546(.A1(new_n745), .A2(new_n746), .A3(new_n737), .ZN(new_n747));
  NOR2_X1   g0547(.A1(G190), .A2(G200), .ZN(new_n748));
  NAND3_X1  g0548(.A1(new_n745), .A2(new_n746), .A3(new_n748), .ZN(new_n749));
  OAI221_X1 g0549(.A(new_n744), .B1(new_n216), .B2(new_n747), .C1(new_n309), .C2(new_n749), .ZN(new_n750));
  AOI21_X1  g0550(.A(KEYINPUT97), .B1(new_n323), .B2(new_n344), .ZN(new_n751));
  NOR2_X1   g0551(.A1(new_n751), .A2(G179), .ZN(new_n752));
  NAND3_X1  g0552(.A1(new_n323), .A2(KEYINPUT97), .A3(new_n344), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  NOR2_X1   g0554(.A1(new_n754), .A2(new_n356), .ZN(new_n755));
  NAND2_X1  g0555(.A1(new_n755), .A2(G107), .ZN(new_n756));
  NAND3_X1  g0556(.A1(new_n734), .A2(G20), .A3(new_n291), .ZN(new_n757));
  OAI211_X1 g0557(.A(new_n756), .B(new_n260), .C1(new_n212), .C2(new_n757), .ZN(new_n758));
  AOI21_X1  g0558(.A(new_n750), .B1(KEYINPUT98), .B2(new_n758), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n754), .A2(G200), .ZN(new_n760));
  NAND2_X1  g0560(.A1(new_n760), .A2(G159), .ZN(new_n761));
  XOR2_X1   g0561(.A(new_n761), .B(KEYINPUT32), .Z(new_n762));
  OAI211_X1 g0562(.A(new_n759), .B(new_n762), .C1(KEYINPUT98), .C2(new_n758), .ZN(new_n763));
  OAI21_X1  g0563(.A(new_n267), .B1(new_n757), .B2(new_n498), .ZN(new_n764));
  AOI21_X1  g0564(.A(new_n764), .B1(G294), .B2(new_n739), .ZN(new_n765));
  INV_X1    g0565(.A(G326), .ZN(new_n766));
  XOR2_X1   g0566(.A(KEYINPUT33), .B(G317), .Z(new_n767));
  OAI221_X1 g0567(.A(new_n765), .B1(new_n766), .B2(new_n735), .C1(new_n733), .C2(new_n767), .ZN(new_n768));
  INV_X1    g0568(.A(new_n749), .ZN(new_n769));
  AOI21_X1  g0569(.A(new_n768), .B1(G311), .B2(new_n769), .ZN(new_n770));
  INV_X1    g0570(.A(new_n747), .ZN(new_n771));
  NAND2_X1  g0571(.A1(new_n771), .A2(G322), .ZN(new_n772));
  AOI22_X1  g0572(.A1(G283), .A2(new_n755), .B1(new_n760), .B2(G329), .ZN(new_n773));
  NAND3_X1  g0573(.A1(new_n770), .A2(new_n772), .A3(new_n773), .ZN(new_n774));
  AND2_X1   g0574(.A1(new_n763), .A2(new_n774), .ZN(new_n775));
  INV_X1    g0575(.A(new_n727), .ZN(new_n776));
  OAI211_X1 g0576(.A(new_n714), .B(new_n729), .C1(new_n775), .C2(new_n776), .ZN(new_n777));
  AND2_X1   g0577(.A1(new_n646), .A2(new_n647), .ZN(new_n778));
  NAND2_X1  g0578(.A1(new_n778), .A2(G330), .ZN(new_n779));
  NAND2_X1  g0579(.A1(new_n779), .A2(new_n720), .ZN(new_n780));
  NOR2_X1   g0580(.A1(new_n778), .A2(G330), .ZN(new_n781));
  OAI21_X1  g0581(.A(new_n777), .B1(new_n780), .B2(new_n781), .ZN(G396));
  NAND2_X1  g0582(.A1(new_n640), .A2(new_n329), .ZN(new_n783));
  XNOR2_X1  g0583(.A(new_n783), .B(KEYINPUT102), .ZN(new_n784));
  OAI22_X1  g0584(.A1(new_n784), .A2(new_n347), .B1(new_n340), .B2(new_n339), .ZN(new_n785));
  NAND2_X1  g0585(.A1(new_n341), .A2(new_n639), .ZN(new_n786));
  NAND2_X1  g0586(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  NAND2_X1  g0587(.A1(new_n701), .A2(new_n787), .ZN(new_n788));
  INV_X1    g0588(.A(new_n787), .ZN(new_n789));
  OAI211_X1 g0589(.A(new_n639), .B(new_n789), .C1(new_n622), .C2(new_n604), .ZN(new_n790));
  NAND2_X1  g0590(.A1(new_n788), .A2(new_n790), .ZN(new_n791));
  OR2_X1    g0591(.A1(new_n791), .A2(new_n685), .ZN(new_n792));
  OR2_X1    g0592(.A1(new_n792), .A2(KEYINPUT103), .ZN(new_n793));
  INV_X1    g0593(.A(KEYINPUT104), .ZN(new_n794));
  AOI21_X1  g0594(.A(new_n719), .B1(new_n792), .B2(KEYINPUT103), .ZN(new_n795));
  NAND3_X1  g0595(.A1(new_n793), .A2(new_n794), .A3(new_n795), .ZN(new_n796));
  NAND2_X1  g0596(.A1(new_n791), .A2(new_n685), .ZN(new_n797));
  NAND2_X1  g0597(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  AOI21_X1  g0598(.A(new_n794), .B1(new_n793), .B2(new_n795), .ZN(new_n799));
  INV_X1    g0599(.A(new_n739), .ZN(new_n800));
  OAI221_X1 g0600(.A(new_n260), .B1(new_n210), .B2(new_n757), .C1(new_n800), .C2(new_n216), .ZN(new_n801));
  INV_X1    g0601(.A(new_n755), .ZN(new_n802));
  NOR2_X1   g0602(.A1(new_n802), .A2(new_n218), .ZN(new_n803));
  AOI211_X1 g0603(.A(new_n801), .B(new_n803), .C1(G132), .C2(new_n760), .ZN(new_n804));
  INV_X1    g0604(.A(new_n735), .ZN(new_n805));
  AOI22_X1  g0605(.A1(new_n732), .A2(G150), .B1(G137), .B2(new_n805), .ZN(new_n806));
  INV_X1    g0606(.A(G159), .ZN(new_n807));
  INV_X1    g0607(.A(G143), .ZN(new_n808));
  OAI221_X1 g0608(.A(new_n806), .B1(new_n749), .B2(new_n807), .C1(new_n808), .C2(new_n747), .ZN(new_n809));
  INV_X1    g0609(.A(KEYINPUT34), .ZN(new_n810));
  NAND2_X1  g0610(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  OR2_X1    g0611(.A1(new_n809), .A2(new_n810), .ZN(new_n812));
  NAND3_X1  g0612(.A1(new_n804), .A2(new_n811), .A3(new_n812), .ZN(new_n813));
  INV_X1    g0613(.A(new_n757), .ZN(new_n814));
  AOI21_X1  g0614(.A(new_n260), .B1(new_n814), .B2(G107), .ZN(new_n815));
  OAI221_X1 g0615(.A(new_n815), .B1(new_n498), .B2(new_n735), .C1(new_n733), .C2(new_n482), .ZN(new_n816));
  AOI21_X1  g0616(.A(new_n816), .B1(G97), .B2(new_n743), .ZN(new_n817));
  AOI22_X1  g0617(.A1(G116), .A2(new_n769), .B1(new_n771), .B2(G294), .ZN(new_n818));
  NAND2_X1  g0618(.A1(new_n760), .A2(G311), .ZN(new_n819));
  NAND2_X1  g0619(.A1(new_n755), .A2(G87), .ZN(new_n820));
  NAND4_X1  g0620(.A1(new_n817), .A2(new_n818), .A3(new_n819), .A4(new_n820), .ZN(new_n821));
  AND3_X1   g0621(.A1(new_n813), .A2(KEYINPUT101), .A3(new_n821), .ZN(new_n822));
  AOI21_X1  g0622(.A(KEYINPUT101), .B1(new_n813), .B2(new_n821), .ZN(new_n823));
  NOR3_X1   g0623(.A1(new_n822), .A2(new_n823), .A3(new_n776), .ZN(new_n824));
  NAND2_X1  g0624(.A1(new_n776), .A2(new_n711), .ZN(new_n825));
  OAI221_X1 g0625(.A(new_n719), .B1(G77), .B2(new_n825), .C1(new_n789), .C2(new_n711), .ZN(new_n826));
  OAI22_X1  g0626(.A1(new_n798), .A2(new_n799), .B1(new_n824), .B2(new_n826), .ZN(G384));
  OAI211_X1 g0627(.A(G116), .B(new_n231), .C1(new_n557), .C2(KEYINPUT35), .ZN(new_n828));
  AOI21_X1  g0628(.A(new_n828), .B1(KEYINPUT35), .B2(new_n557), .ZN(new_n829));
  XNOR2_X1  g0629(.A(new_n829), .B(KEYINPUT36), .ZN(new_n830));
  OR3_X1    g0630(.A1(new_n235), .A2(new_n309), .A3(new_n374), .ZN(new_n831));
  NAND2_X1  g0631(.A1(new_n210), .A2(G68), .ZN(new_n832));
  AOI211_X1 g0632(.A(new_n205), .B(G13), .C1(new_n831), .C2(new_n832), .ZN(new_n833));
  NOR2_X1   g0633(.A1(new_n830), .A2(new_n833), .ZN(new_n834));
  NOR2_X1   g0634(.A1(new_n382), .A2(KEYINPUT16), .ZN(new_n835));
  OAI21_X1  g0635(.A(new_n373), .B1(new_n384), .B2(new_n835), .ZN(new_n836));
  NAND2_X1  g0636(.A1(new_n836), .A2(new_n637), .ZN(new_n837));
  INV_X1    g0637(.A(new_n837), .ZN(new_n838));
  NAND2_X1  g0638(.A1(new_n428), .A2(new_n838), .ZN(new_n839));
  INV_X1    g0639(.A(KEYINPUT37), .ZN(new_n840));
  NAND2_X1  g0640(.A1(new_n410), .A2(new_n413), .ZN(new_n841));
  INV_X1    g0641(.A(new_n395), .ZN(new_n842));
  NAND2_X1  g0642(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  NAND3_X1  g0643(.A1(new_n419), .A2(new_n422), .A3(new_n836), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  INV_X1    g0645(.A(KEYINPUT105), .ZN(new_n846));
  AOI21_X1  g0646(.A(new_n838), .B1(new_n845), .B2(new_n846), .ZN(new_n847));
  NAND3_X1  g0647(.A1(new_n843), .A2(KEYINPUT105), .A3(new_n844), .ZN(new_n848));
  AOI21_X1  g0648(.A(new_n840), .B1(new_n847), .B2(new_n848), .ZN(new_n849));
  NAND2_X1  g0649(.A1(new_n395), .A2(new_n637), .ZN(new_n850));
  NAND4_X1  g0650(.A1(new_n843), .A2(new_n840), .A3(new_n423), .A4(new_n850), .ZN(new_n851));
  INV_X1    g0651(.A(new_n851), .ZN(new_n852));
  OAI211_X1 g0652(.A(new_n839), .B(KEYINPUT38), .C1(new_n849), .C2(new_n852), .ZN(new_n853));
  INV_X1    g0653(.A(KEYINPUT38), .ZN(new_n854));
  AND3_X1   g0654(.A1(new_n419), .A2(new_n422), .A3(new_n836), .ZN(new_n855));
  OAI21_X1  g0655(.A(new_n846), .B1(new_n855), .B2(new_n414), .ZN(new_n856));
  NAND3_X1  g0656(.A1(new_n856), .A2(new_n848), .A3(new_n837), .ZN(new_n857));
  AOI21_X1  g0657(.A(new_n852), .B1(new_n857), .B2(KEYINPUT37), .ZN(new_n858));
  AOI21_X1  g0658(.A(new_n837), .B1(new_n416), .B2(new_n427), .ZN(new_n859));
  OAI21_X1  g0659(.A(new_n854), .B1(new_n858), .B2(new_n859), .ZN(new_n860));
  INV_X1    g0660(.A(KEYINPUT106), .ZN(new_n861));
  NAND3_X1  g0661(.A1(new_n853), .A2(new_n860), .A3(new_n861), .ZN(new_n862));
  OAI211_X1 g0662(.A(KEYINPUT106), .B(new_n854), .C1(new_n858), .C2(new_n859), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n316), .A2(new_n639), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n314), .A2(new_n640), .ZN(new_n865));
  AOI22_X1  g0665(.A1(new_n293), .A2(new_n314), .B1(new_n345), .B2(new_n865), .ZN(new_n866));
  INV_X1    g0666(.A(new_n866), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n864), .A2(new_n867), .ZN(new_n868));
  NOR3_X1   g0668(.A1(new_n683), .A2(new_n868), .A3(new_n787), .ZN(new_n869));
  NAND3_X1  g0669(.A1(new_n862), .A2(new_n863), .A3(new_n869), .ZN(new_n870));
  INV_X1    g0670(.A(KEYINPUT40), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  NOR2_X1   g0672(.A1(new_n315), .A2(new_n640), .ZN(new_n873));
  NOR3_X1   g0673(.A1(new_n873), .A2(new_n866), .A3(new_n787), .ZN(new_n874));
  NAND4_X1  g0674(.A1(new_n874), .A2(KEYINPUT40), .A3(new_n681), .A4(new_n682), .ZN(new_n875));
  AOI21_X1  g0675(.A(new_n850), .B1(new_n627), .B2(new_n416), .ZN(new_n876));
  INV_X1    g0676(.A(KEYINPUT107), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n423), .A2(new_n850), .ZN(new_n878));
  OR4_X1    g0678(.A1(new_n877), .A2(new_n878), .A3(KEYINPUT37), .A4(new_n414), .ZN(new_n879));
  OAI21_X1  g0679(.A(KEYINPUT37), .B1(new_n878), .B2(new_n414), .ZN(new_n880));
  NAND3_X1  g0680(.A1(new_n880), .A2(new_n877), .A3(new_n851), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n879), .A2(new_n881), .ZN(new_n882));
  OAI21_X1  g0682(.A(new_n854), .B1(new_n876), .B2(new_n882), .ZN(new_n883));
  AOI21_X1  g0683(.A(new_n875), .B1(new_n883), .B2(new_n853), .ZN(new_n884));
  INV_X1    g0684(.A(new_n884), .ZN(new_n885));
  NAND3_X1  g0685(.A1(new_n872), .A2(G330), .A3(new_n885), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n686), .A2(new_n601), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  AOI21_X1  g0688(.A(new_n884), .B1(new_n870), .B2(new_n871), .ZN(new_n889));
  NAND3_X1  g0689(.A1(new_n889), .A2(new_n601), .A3(new_n684), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n888), .A2(new_n890), .ZN(new_n891));
  OAI21_X1  g0691(.A(KEYINPUT91), .B1(new_n697), .B2(KEYINPUT26), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n480), .A2(new_n603), .ZN(new_n893));
  NAND3_X1  g0693(.A1(new_n893), .A2(new_n695), .A3(new_n602), .ZN(new_n894));
  NAND3_X1  g0694(.A1(new_n892), .A2(new_n894), .A3(new_n693), .ZN(new_n895));
  AOI211_X1 g0695(.A(new_n702), .B(new_n640), .C1(new_n895), .C2(new_n692), .ZN(new_n896));
  AOI21_X1  g0696(.A(KEYINPUT93), .B1(new_n701), .B2(new_n702), .ZN(new_n897));
  OAI211_X1 g0697(.A(new_n601), .B(new_n707), .C1(new_n896), .C2(new_n897), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n898), .A2(new_n631), .ZN(new_n899));
  XOR2_X1   g0699(.A(new_n891), .B(new_n899), .Z(new_n900));
  NAND2_X1  g0700(.A1(new_n790), .A2(new_n786), .ZN(new_n901));
  INV_X1    g0701(.A(new_n868), .ZN(new_n902));
  NAND4_X1  g0702(.A1(new_n862), .A2(new_n863), .A3(new_n901), .A4(new_n902), .ZN(new_n903));
  OR2_X1    g0703(.A1(new_n627), .A2(new_n637), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  NAND3_X1  g0705(.A1(new_n862), .A2(KEYINPUT39), .A3(new_n863), .ZN(new_n906));
  INV_X1    g0706(.A(KEYINPUT39), .ZN(new_n907));
  NAND3_X1  g0707(.A1(new_n883), .A2(new_n907), .A3(new_n853), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n906), .A2(new_n908), .ZN(new_n909));
  AOI21_X1  g0709(.A(new_n905), .B1(new_n873), .B2(new_n909), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n900), .A2(new_n910), .ZN(new_n911));
  OAI21_X1  g0711(.A(new_n911), .B1(new_n205), .B2(new_n716), .ZN(new_n912));
  NOR2_X1   g0712(.A1(new_n900), .A2(new_n910), .ZN(new_n913));
  OAI21_X1  g0713(.A(new_n834), .B1(new_n912), .B2(new_n913), .ZN(G367));
  INV_X1    g0714(.A(KEYINPUT45), .ZN(new_n915));
  NOR2_X1   g0715(.A1(new_n585), .A2(new_n639), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n565), .A2(new_n640), .ZN(new_n917));
  AOI21_X1  g0717(.A(new_n916), .B1(new_n691), .B2(new_n917), .ZN(new_n918));
  OAI22_X1  g0718(.A1(new_n652), .A2(new_n656), .B1(new_n613), .B2(new_n640), .ZN(new_n919));
  OAI21_X1  g0719(.A(new_n915), .B1(new_n918), .B2(new_n919), .ZN(new_n920));
  AND3_X1   g0720(.A1(new_n585), .A2(new_n591), .A3(new_n689), .ZN(new_n921));
  AOI21_X1  g0721(.A(new_n689), .B1(new_n585), .B2(new_n591), .ZN(new_n922));
  OAI21_X1  g0722(.A(new_n917), .B1(new_n921), .B2(new_n922), .ZN(new_n923));
  INV_X1    g0723(.A(new_n916), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  NAND3_X1  g0725(.A1(new_n925), .A2(KEYINPUT45), .A3(new_n660), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n920), .A2(new_n926), .ZN(new_n927));
  INV_X1    g0727(.A(KEYINPUT44), .ZN(new_n928));
  OAI21_X1  g0728(.A(new_n928), .B1(new_n925), .B2(new_n660), .ZN(new_n929));
  NAND3_X1  g0729(.A1(new_n918), .A2(new_n919), .A3(KEYINPUT44), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  AND3_X1   g0731(.A1(new_n927), .A2(new_n931), .A3(new_n655), .ZN(new_n932));
  AOI21_X1  g0732(.A(new_n655), .B1(new_n927), .B2(new_n931), .ZN(new_n933));
  OR2_X1    g0733(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  NOR2_X1   g0734(.A1(new_n654), .A2(new_n657), .ZN(new_n935));
  NOR3_X1   g0735(.A1(new_n652), .A2(new_n653), .A3(new_n656), .ZN(new_n936));
  NOR2_X1   g0736(.A1(new_n935), .A2(new_n936), .ZN(new_n937));
  XNOR2_X1  g0737(.A(new_n779), .B(new_n937), .ZN(new_n938));
  INV_X1    g0738(.A(new_n938), .ZN(new_n939));
  OAI21_X1  g0739(.A(new_n708), .B1(new_n934), .B2(new_n939), .ZN(new_n940));
  XNOR2_X1  g0740(.A(new_n663), .B(KEYINPUT41), .ZN(new_n941));
  AOI21_X1  g0741(.A(new_n718), .B1(new_n940), .B2(new_n941), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n936), .A2(new_n925), .ZN(new_n943));
  AND2_X1   g0743(.A1(new_n943), .A2(KEYINPUT42), .ZN(new_n944));
  NAND3_X1  g0744(.A1(new_n691), .A2(new_n550), .A3(new_n917), .ZN(new_n945));
  AOI21_X1  g0745(.A(new_n640), .B1(new_n945), .B2(new_n585), .ZN(new_n946));
  NOR2_X1   g0746(.A1(new_n944), .A2(new_n946), .ZN(new_n947));
  OAI21_X1  g0747(.A(new_n947), .B1(KEYINPUT42), .B2(new_n943), .ZN(new_n948));
  OR2_X1    g0748(.A1(new_n463), .A2(new_n639), .ZN(new_n949));
  OR2_X1    g0749(.A1(new_n949), .A2(new_n608), .ZN(new_n950));
  NAND3_X1  g0750(.A1(new_n949), .A2(new_n608), .A3(new_n609), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n950), .A2(new_n951), .ZN(new_n952));
  INV_X1    g0752(.A(KEYINPUT108), .ZN(new_n953));
  AOI21_X1  g0753(.A(KEYINPUT43), .B1(new_n952), .B2(new_n953), .ZN(new_n954));
  NAND3_X1  g0754(.A1(new_n950), .A2(KEYINPUT108), .A3(new_n951), .ZN(new_n955));
  AND2_X1   g0755(.A1(new_n954), .A2(new_n955), .ZN(new_n956));
  AOI21_X1  g0756(.A(new_n956), .B1(KEYINPUT43), .B2(new_n952), .ZN(new_n957));
  AND2_X1   g0757(.A1(new_n948), .A2(new_n957), .ZN(new_n958));
  INV_X1    g0758(.A(new_n956), .ZN(new_n959));
  NOR2_X1   g0759(.A1(new_n948), .A2(new_n959), .ZN(new_n960));
  OAI22_X1  g0760(.A1(new_n958), .A2(new_n960), .B1(new_n655), .B2(new_n918), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n948), .A2(new_n957), .ZN(new_n962));
  NOR2_X1   g0762(.A1(new_n655), .A2(new_n918), .ZN(new_n963));
  OAI211_X1 g0763(.A(new_n962), .B(new_n963), .C1(new_n948), .C2(new_n959), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n961), .A2(new_n964), .ZN(new_n965));
  INV_X1    g0765(.A(new_n713), .ZN(new_n966));
  NOR2_X1   g0766(.A1(new_n952), .A2(new_n966), .ZN(new_n967));
  INV_X1    g0767(.A(G311), .ZN(new_n968));
  OAI22_X1  g0768(.A1(new_n733), .A2(new_n540), .B1(new_n968), .B2(new_n735), .ZN(new_n969));
  INV_X1    g0769(.A(KEYINPUT46), .ZN(new_n970));
  OAI21_X1  g0770(.A(new_n970), .B1(new_n757), .B2(new_n484), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n971), .A2(new_n267), .ZN(new_n972));
  NOR3_X1   g0772(.A1(new_n757), .A2(new_n970), .A3(new_n484), .ZN(new_n973));
  NOR2_X1   g0773(.A1(new_n800), .A2(new_n330), .ZN(new_n974));
  NOR4_X1   g0774(.A1(new_n969), .A2(new_n972), .A3(new_n973), .A4(new_n974), .ZN(new_n975));
  OAI221_X1 g0775(.A(new_n975), .B1(new_n482), .B2(new_n749), .C1(new_n498), .C2(new_n747), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n755), .A2(G97), .ZN(new_n977));
  INV_X1    g0777(.A(new_n760), .ZN(new_n978));
  INV_X1    g0778(.A(G317), .ZN(new_n979));
  OAI21_X1  g0779(.A(new_n977), .B1(new_n978), .B2(new_n979), .ZN(new_n980));
  AOI22_X1  g0780(.A1(G50), .A2(new_n769), .B1(new_n771), .B2(G150), .ZN(new_n981));
  OAI221_X1 g0781(.A(new_n260), .B1(new_n216), .B2(new_n757), .C1(new_n735), .C2(new_n808), .ZN(new_n982));
  AOI21_X1  g0782(.A(new_n982), .B1(G159), .B2(new_n732), .ZN(new_n983));
  OAI211_X1 g0783(.A(new_n981), .B(new_n983), .C1(new_n218), .C2(new_n742), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n755), .A2(G77), .ZN(new_n985));
  XOR2_X1   g0785(.A(KEYINPUT109), .B(G137), .Z(new_n986));
  OAI21_X1  g0786(.A(new_n985), .B1(new_n978), .B2(new_n986), .ZN(new_n987));
  OAI22_X1  g0787(.A1(new_n976), .A2(new_n980), .B1(new_n984), .B2(new_n987), .ZN(new_n988));
  INV_X1    g0788(.A(KEYINPUT47), .ZN(new_n989));
  AOI21_X1  g0789(.A(new_n776), .B1(new_n988), .B2(new_n989), .ZN(new_n990));
  OAI21_X1  g0790(.A(new_n990), .B1(new_n989), .B2(new_n988), .ZN(new_n991));
  INV_X1    g0791(.A(new_n722), .ZN(new_n992));
  OAI221_X1 g0792(.A(new_n728), .B1(new_n226), .B2(new_n326), .C1(new_n992), .C2(new_n245), .ZN(new_n993));
  NAND3_X1  g0793(.A1(new_n991), .A2(new_n719), .A3(new_n993), .ZN(new_n994));
  XNOR2_X1  g0794(.A(new_n994), .B(KEYINPUT110), .ZN(new_n995));
  OAI22_X1  g0795(.A1(new_n942), .A2(new_n965), .B1(new_n967), .B2(new_n995), .ZN(G387));
  NAND2_X1  g0796(.A1(new_n938), .A2(new_n718), .ZN(new_n997));
  XOR2_X1   g0797(.A(KEYINPUT112), .B(G150), .Z(new_n998));
  OAI21_X1  g0798(.A(new_n977), .B1(new_n978), .B2(new_n998), .ZN(new_n999));
  OAI22_X1  g0799(.A1(new_n210), .A2(new_n747), .B1(new_n749), .B2(new_n218), .ZN(new_n1000));
  AOI21_X1  g0800(.A(new_n267), .B1(new_n814), .B2(G77), .ZN(new_n1001));
  OAI221_X1 g0801(.A(new_n1001), .B1(new_n807), .B2(new_n735), .C1(new_n733), .C2(new_n319), .ZN(new_n1002));
  NOR2_X1   g0802(.A1(new_n742), .A2(new_n326), .ZN(new_n1003));
  NOR4_X1   g0803(.A1(new_n999), .A2(new_n1000), .A3(new_n1002), .A4(new_n1003), .ZN(new_n1004));
  AOI22_X1  g0804(.A1(new_n732), .A2(G311), .B1(G322), .B2(new_n805), .ZN(new_n1005));
  OAI221_X1 g0805(.A(new_n1005), .B1(new_n749), .B2(new_n498), .C1(new_n979), .C2(new_n747), .ZN(new_n1006));
  XNOR2_X1  g0806(.A(new_n1006), .B(KEYINPUT113), .ZN(new_n1007));
  INV_X1    g0807(.A(KEYINPUT48), .ZN(new_n1008));
  OR2_X1    g0808(.A1(new_n1007), .A2(new_n1008), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n1007), .A2(new_n1008), .ZN(new_n1010));
  AOI22_X1  g0810(.A1(G294), .A2(new_n814), .B1(new_n739), .B2(G283), .ZN(new_n1011));
  NAND3_X1  g0811(.A1(new_n1009), .A2(new_n1010), .A3(new_n1011), .ZN(new_n1012));
  INV_X1    g0812(.A(KEYINPUT49), .ZN(new_n1013));
  OR2_X1    g0813(.A1(new_n1012), .A2(new_n1013), .ZN(new_n1014));
  OAI221_X1 g0814(.A(new_n267), .B1(new_n802), .B2(new_n484), .C1(new_n766), .C2(new_n978), .ZN(new_n1015));
  AOI21_X1  g0815(.A(new_n1015), .B1(new_n1012), .B2(new_n1013), .ZN(new_n1016));
  AOI21_X1  g0816(.A(new_n1004), .B1(new_n1014), .B2(new_n1016), .ZN(new_n1017));
  NOR2_X1   g0817(.A1(new_n1017), .A2(new_n776), .ZN(new_n1018));
  INV_X1    g0818(.A(new_n728), .ZN(new_n1019));
  INV_X1    g0819(.A(new_n665), .ZN(new_n1020));
  NAND3_X1  g0820(.A1(new_n1020), .A2(new_n226), .A3(new_n260), .ZN(new_n1021));
  OAI21_X1  g0821(.A(new_n1021), .B1(G107), .B2(new_n226), .ZN(new_n1022));
  AOI21_X1  g0822(.A(KEYINPUT111), .B1(new_n242), .B2(G45), .ZN(new_n1023));
  NAND2_X1  g0823(.A1(new_n320), .A2(new_n210), .ZN(new_n1024));
  OR2_X1    g0824(.A1(new_n1024), .A2(KEYINPUT50), .ZN(new_n1025));
  OAI21_X1  g0825(.A(new_n429), .B1(new_n218), .B2(new_n309), .ZN(new_n1026));
  AOI211_X1 g0826(.A(new_n1026), .B(new_n1020), .C1(KEYINPUT50), .C2(new_n1024), .ZN(new_n1027));
  AOI211_X1 g0827(.A(new_n992), .B(new_n1023), .C1(new_n1025), .C2(new_n1027), .ZN(new_n1028));
  NAND3_X1  g0828(.A1(new_n242), .A2(KEYINPUT111), .A3(G45), .ZN(new_n1029));
  AOI21_X1  g0829(.A(new_n1022), .B1(new_n1028), .B2(new_n1029), .ZN(new_n1030));
  OAI221_X1 g0830(.A(new_n719), .B1(new_n1019), .B2(new_n1030), .C1(new_n654), .C2(new_n966), .ZN(new_n1031));
  OAI21_X1  g0831(.A(new_n707), .B1(new_n896), .B2(new_n897), .ZN(new_n1032));
  NAND3_X1  g0832(.A1(new_n1032), .A2(new_n685), .A3(new_n938), .ZN(new_n1033));
  NAND2_X1  g0833(.A1(new_n1033), .A2(new_n663), .ZN(new_n1034));
  NOR2_X1   g0834(.A1(new_n708), .A2(new_n938), .ZN(new_n1035));
  OAI221_X1 g0835(.A(new_n997), .B1(new_n1018), .B2(new_n1031), .C1(new_n1034), .C2(new_n1035), .ZN(G393));
  NOR2_X1   g0836(.A1(new_n932), .A2(new_n933), .ZN(new_n1037));
  NAND4_X1  g0837(.A1(new_n1032), .A2(new_n685), .A3(new_n1037), .A4(new_n938), .ZN(new_n1038));
  NAND2_X1  g0838(.A1(new_n1038), .A2(new_n663), .ZN(new_n1039));
  AOI21_X1  g0839(.A(new_n1037), .B1(new_n708), .B2(new_n938), .ZN(new_n1040));
  OAI21_X1  g0840(.A(KEYINPUT117), .B1(new_n1039), .B2(new_n1040), .ZN(new_n1041));
  NAND2_X1  g0841(.A1(new_n1033), .A2(new_n934), .ZN(new_n1042));
  INV_X1    g0842(.A(KEYINPUT117), .ZN(new_n1043));
  NAND4_X1  g0843(.A1(new_n1042), .A2(new_n1043), .A3(new_n663), .A4(new_n1038), .ZN(new_n1044));
  NAND2_X1  g0844(.A1(new_n1041), .A2(new_n1044), .ZN(new_n1045));
  NAND2_X1  g0845(.A1(new_n934), .A2(KEYINPUT114), .ZN(new_n1046));
  INV_X1    g0846(.A(KEYINPUT114), .ZN(new_n1047));
  NAND2_X1  g0847(.A1(new_n1037), .A2(new_n1047), .ZN(new_n1048));
  NAND3_X1  g0848(.A1(new_n1046), .A2(new_n718), .A3(new_n1048), .ZN(new_n1049));
  OAI22_X1  g0849(.A1(new_n747), .A2(new_n807), .B1(new_n349), .B2(new_n735), .ZN(new_n1050));
  XOR2_X1   g0850(.A(new_n1050), .B(KEYINPUT51), .Z(new_n1051));
  OAI221_X1 g0851(.A(new_n260), .B1(new_n218), .B2(new_n757), .C1(new_n733), .C2(new_n210), .ZN(new_n1052));
  AOI21_X1  g0852(.A(new_n1052), .B1(G77), .B2(new_n743), .ZN(new_n1053));
  OAI211_X1 g0853(.A(new_n1053), .B(new_n820), .C1(new_n319), .C2(new_n749), .ZN(new_n1054));
  AOI211_X1 g0854(.A(new_n1051), .B(new_n1054), .C1(G143), .C2(new_n760), .ZN(new_n1055));
  XNOR2_X1  g0855(.A(new_n1055), .B(KEYINPUT115), .ZN(new_n1056));
  OAI221_X1 g0856(.A(new_n267), .B1(new_n482), .B2(new_n757), .C1(new_n800), .C2(new_n484), .ZN(new_n1057));
  AOI21_X1  g0857(.A(new_n1057), .B1(G303), .B2(new_n732), .ZN(new_n1058));
  OAI211_X1 g0858(.A(new_n1058), .B(new_n756), .C1(new_n540), .C2(new_n749), .ZN(new_n1059));
  OAI22_X1  g0859(.A1(new_n747), .A2(new_n968), .B1(new_n979), .B2(new_n735), .ZN(new_n1060));
  XOR2_X1   g0860(.A(new_n1060), .B(KEYINPUT52), .Z(new_n1061));
  AOI211_X1 g0861(.A(new_n1059), .B(new_n1061), .C1(G322), .C2(new_n760), .ZN(new_n1062));
  XNOR2_X1  g0862(.A(new_n1062), .B(KEYINPUT116), .ZN(new_n1063));
  OAI21_X1  g0863(.A(new_n727), .B1(new_n1056), .B2(new_n1063), .ZN(new_n1064));
  NAND2_X1  g0864(.A1(new_n918), .A2(new_n712), .ZN(new_n1065));
  OAI221_X1 g0865(.A(new_n728), .B1(new_n454), .B2(new_n226), .C1(new_n992), .C2(new_n252), .ZN(new_n1066));
  NAND4_X1  g0866(.A1(new_n1064), .A2(new_n719), .A3(new_n1065), .A4(new_n1066), .ZN(new_n1067));
  NAND2_X1  g0867(.A1(new_n1049), .A2(new_n1067), .ZN(new_n1068));
  INV_X1    g0868(.A(new_n1068), .ZN(new_n1069));
  NAND2_X1  g0869(.A1(new_n1045), .A2(new_n1069), .ZN(G390));
  NAND4_X1  g0870(.A1(new_n874), .A2(G330), .A3(new_n681), .A4(new_n682), .ZN(new_n1071));
  INV_X1    g0871(.A(new_n1071), .ZN(new_n1072));
  NAND2_X1  g0872(.A1(new_n901), .A2(new_n902), .ZN(new_n1073));
  NAND2_X1  g0873(.A1(new_n1073), .A2(new_n864), .ZN(new_n1074));
  AND3_X1   g0874(.A1(new_n906), .A2(new_n908), .A3(new_n1074), .ZN(new_n1075));
  NAND3_X1  g0875(.A1(new_n699), .A2(new_n639), .A3(new_n785), .ZN(new_n1076));
  NAND3_X1  g0876(.A1(new_n1076), .A2(new_n786), .A3(new_n864), .ZN(new_n1077));
  AOI22_X1  g0877(.A1(new_n1077), .A2(new_n867), .B1(new_n853), .B2(new_n883), .ZN(new_n1078));
  OAI21_X1  g0878(.A(new_n1072), .B1(new_n1075), .B2(new_n1078), .ZN(new_n1079));
  NAND3_X1  g0879(.A1(new_n906), .A2(new_n908), .A3(new_n1074), .ZN(new_n1080));
  AND2_X1   g0880(.A1(new_n1077), .A2(new_n867), .ZN(new_n1081));
  AND2_X1   g0881(.A1(new_n883), .A2(new_n853), .ZN(new_n1082));
  OAI211_X1 g0882(.A(new_n1080), .B(new_n1071), .C1(new_n1081), .C2(new_n1082), .ZN(new_n1083));
  NAND2_X1  g0883(.A1(new_n1079), .A2(new_n1083), .ZN(new_n1084));
  NAND3_X1  g0884(.A1(new_n898), .A2(new_n631), .A3(new_n887), .ZN(new_n1085));
  NAND4_X1  g0885(.A1(new_n681), .A2(G330), .A3(new_n682), .A4(new_n789), .ZN(new_n1086));
  NAND2_X1  g0886(.A1(new_n1086), .A2(new_n868), .ZN(new_n1087));
  AOI22_X1  g0887(.A1(new_n1087), .A2(new_n1071), .B1(new_n786), .B2(new_n790), .ZN(new_n1088));
  AND2_X1   g0888(.A1(new_n1076), .A2(new_n786), .ZN(new_n1089));
  AND2_X1   g0889(.A1(new_n1087), .A2(new_n1071), .ZN(new_n1090));
  AOI21_X1  g0890(.A(new_n1088), .B1(new_n1089), .B2(new_n1090), .ZN(new_n1091));
  NOR2_X1   g0891(.A1(new_n1085), .A2(new_n1091), .ZN(new_n1092));
  INV_X1    g0892(.A(new_n1092), .ZN(new_n1093));
  NAND2_X1  g0893(.A1(new_n1084), .A2(new_n1093), .ZN(new_n1094));
  NAND3_X1  g0894(.A1(new_n1079), .A2(new_n1083), .A3(new_n1092), .ZN(new_n1095));
  NAND3_X1  g0895(.A1(new_n1094), .A2(new_n663), .A3(new_n1095), .ZN(new_n1096));
  NAND3_X1  g0896(.A1(new_n1079), .A2(new_n1083), .A3(new_n718), .ZN(new_n1097));
  OAI21_X1  g0897(.A(new_n719), .B1(new_n320), .B2(new_n825), .ZN(new_n1098));
  NOR2_X1   g0898(.A1(new_n757), .A2(new_n998), .ZN(new_n1099));
  INV_X1    g0899(.A(KEYINPUT53), .ZN(new_n1100));
  OAI21_X1  g0900(.A(new_n260), .B1(new_n1099), .B2(new_n1100), .ZN(new_n1101));
  NAND2_X1  g0901(.A1(new_n805), .A2(G128), .ZN(new_n1102));
  OAI21_X1  g0902(.A(new_n1102), .B1(new_n733), .B2(new_n986), .ZN(new_n1103));
  AOI211_X1 g0903(.A(new_n1101), .B(new_n1103), .C1(new_n1100), .C2(new_n1099), .ZN(new_n1104));
  XOR2_X1   g0904(.A(KEYINPUT54), .B(G143), .Z(new_n1105));
  AOI22_X1  g0905(.A1(G132), .A2(new_n771), .B1(new_n769), .B2(new_n1105), .ZN(new_n1106));
  OAI211_X1 g0906(.A(new_n1104), .B(new_n1106), .C1(new_n807), .C2(new_n742), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n760), .A2(G125), .ZN(new_n1108));
  OAI21_X1  g0908(.A(new_n1108), .B1(new_n802), .B2(new_n210), .ZN(new_n1109));
  INV_X1    g0909(.A(new_n803), .ZN(new_n1110));
  NAND2_X1  g0910(.A1(new_n760), .A2(G294), .ZN(new_n1111));
  NAND2_X1  g0911(.A1(new_n769), .A2(G97), .ZN(new_n1112));
  OAI221_X1 g0912(.A(new_n267), .B1(new_n212), .B2(new_n757), .C1(new_n735), .C2(new_n482), .ZN(new_n1113));
  AOI21_X1  g0913(.A(new_n1113), .B1(G107), .B2(new_n732), .ZN(new_n1114));
  NAND4_X1  g0914(.A1(new_n1110), .A2(new_n1111), .A3(new_n1112), .A4(new_n1114), .ZN(new_n1115));
  OAI22_X1  g0915(.A1(new_n747), .A2(new_n484), .B1(new_n742), .B2(new_n309), .ZN(new_n1116));
  XOR2_X1   g0916(.A(new_n1116), .B(KEYINPUT118), .Z(new_n1117));
  OAI22_X1  g0917(.A1(new_n1107), .A2(new_n1109), .B1(new_n1115), .B2(new_n1117), .ZN(new_n1118));
  AOI21_X1  g0918(.A(new_n1098), .B1(new_n1118), .B2(new_n727), .ZN(new_n1119));
  OAI21_X1  g0919(.A(new_n1119), .B1(new_n909), .B2(new_n711), .ZN(new_n1120));
  AND2_X1   g0920(.A1(new_n1097), .A2(new_n1120), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n1096), .A2(new_n1121), .ZN(G378));
  NAND2_X1  g0922(.A1(new_n909), .A2(new_n873), .ZN(new_n1123));
  NAND3_X1  g0923(.A1(new_n1123), .A2(new_n904), .A3(new_n903), .ZN(new_n1124));
  NAND2_X1  g0924(.A1(new_n630), .A2(new_n368), .ZN(new_n1125));
  AND3_X1   g0925(.A1(new_n1125), .A2(new_n354), .A3(new_n637), .ZN(new_n1126));
  AOI21_X1  g0926(.A(new_n1125), .B1(new_n354), .B2(new_n637), .ZN(new_n1127));
  XNOR2_X1  g0927(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1128));
  INV_X1    g0928(.A(new_n1128), .ZN(new_n1129));
  OR3_X1    g0929(.A1(new_n1126), .A2(new_n1127), .A3(new_n1129), .ZN(new_n1130));
  OAI21_X1  g0930(.A(new_n1129), .B1(new_n1126), .B2(new_n1127), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n1130), .A2(new_n1131), .ZN(new_n1132));
  AND4_X1   g0932(.A1(G330), .A2(new_n872), .A3(new_n885), .A4(new_n1132), .ZN(new_n1133));
  AOI21_X1  g0933(.A(new_n1132), .B1(new_n889), .B2(G330), .ZN(new_n1134));
  OAI21_X1  g0934(.A(new_n1124), .B1(new_n1133), .B2(new_n1134), .ZN(new_n1135));
  INV_X1    g0935(.A(new_n1132), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n886), .A2(new_n1136), .ZN(new_n1137));
  NAND3_X1  g0937(.A1(new_n889), .A2(G330), .A3(new_n1132), .ZN(new_n1138));
  NAND3_X1  g0938(.A1(new_n1137), .A2(new_n910), .A3(new_n1138), .ZN(new_n1139));
  INV_X1    g0939(.A(KEYINPUT120), .ZN(new_n1140));
  NAND3_X1  g0940(.A1(new_n1135), .A2(new_n1139), .A3(new_n1140), .ZN(new_n1141));
  AOI21_X1  g0941(.A(new_n910), .B1(new_n1137), .B2(new_n1138), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n1142), .A2(KEYINPUT120), .ZN(new_n1143));
  INV_X1    g0943(.A(KEYINPUT121), .ZN(new_n1144));
  XNOR2_X1  g0944(.A(new_n1085), .B(new_n1144), .ZN(new_n1145));
  NAND2_X1  g0945(.A1(new_n1095), .A2(new_n1145), .ZN(new_n1146));
  NAND3_X1  g0946(.A1(new_n1141), .A2(new_n1143), .A3(new_n1146), .ZN(new_n1147));
  INV_X1    g0947(.A(KEYINPUT57), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n1147), .A2(new_n1148), .ZN(new_n1149));
  AOI21_X1  g0949(.A(new_n1148), .B1(new_n1135), .B2(new_n1139), .ZN(new_n1150));
  AOI21_X1  g0950(.A(new_n664), .B1(new_n1150), .B2(new_n1146), .ZN(new_n1151));
  NAND2_X1  g0951(.A1(new_n1149), .A2(new_n1151), .ZN(new_n1152));
  NAND3_X1  g0952(.A1(new_n1141), .A2(new_n718), .A3(new_n1143), .ZN(new_n1153));
  OAI21_X1  g0953(.A(new_n719), .B1(G50), .B2(new_n825), .ZN(new_n1154));
  NOR2_X1   g0954(.A1(new_n260), .A2(G41), .ZN(new_n1155));
  AOI211_X1 g0955(.A(G50), .B(new_n1155), .C1(new_n263), .C2(new_n503), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n755), .A2(G58), .ZN(new_n1157));
  OAI21_X1  g0957(.A(new_n1157), .B1(new_n978), .B2(new_n482), .ZN(new_n1158));
  OAI21_X1  g0958(.A(new_n1155), .B1(new_n309), .B2(new_n757), .ZN(new_n1159));
  AOI21_X1  g0959(.A(new_n1159), .B1(new_n732), .B2(G97), .ZN(new_n1160));
  OAI221_X1 g0960(.A(new_n1160), .B1(new_n484), .B2(new_n735), .C1(new_n218), .C2(new_n742), .ZN(new_n1161));
  OAI22_X1  g0961(.A1(new_n330), .A2(new_n747), .B1(new_n749), .B2(new_n326), .ZN(new_n1162));
  NOR3_X1   g0962(.A1(new_n1158), .A2(new_n1161), .A3(new_n1162), .ZN(new_n1163));
  AOI21_X1  g0963(.A(new_n1156), .B1(new_n1163), .B2(KEYINPUT58), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n760), .A2(G124), .ZN(new_n1165));
  AOI211_X1 g0965(.A(G33), .B(G41), .C1(new_n755), .C2(G159), .ZN(new_n1166));
  AOI22_X1  g0966(.A1(new_n732), .A2(G132), .B1(G125), .B2(new_n805), .ZN(new_n1167));
  INV_X1    g0967(.A(G137), .ZN(new_n1168));
  OAI221_X1 g0968(.A(new_n1167), .B1(new_n349), .B2(new_n742), .C1(new_n749), .C2(new_n1168), .ZN(new_n1169));
  AOI22_X1  g0969(.A1(new_n771), .A2(G128), .B1(new_n814), .B2(new_n1105), .ZN(new_n1170));
  OR2_X1    g0970(.A1(new_n1170), .A2(KEYINPUT119), .ZN(new_n1171));
  NAND2_X1  g0971(.A1(new_n1170), .A2(KEYINPUT119), .ZN(new_n1172));
  AOI21_X1  g0972(.A(new_n1169), .B1(new_n1171), .B2(new_n1172), .ZN(new_n1173));
  INV_X1    g0973(.A(KEYINPUT59), .ZN(new_n1174));
  OAI211_X1 g0974(.A(new_n1165), .B(new_n1166), .C1(new_n1173), .C2(new_n1174), .ZN(new_n1175));
  AND2_X1   g0975(.A1(new_n1173), .A2(new_n1174), .ZN(new_n1176));
  OAI221_X1 g0976(.A(new_n1164), .B1(KEYINPUT58), .B2(new_n1163), .C1(new_n1175), .C2(new_n1176), .ZN(new_n1177));
  AOI21_X1  g0977(.A(new_n1154), .B1(new_n1177), .B2(new_n727), .ZN(new_n1178));
  OAI21_X1  g0978(.A(new_n1178), .B1(new_n1132), .B2(new_n711), .ZN(new_n1179));
  NAND2_X1  g0979(.A1(new_n1153), .A2(new_n1179), .ZN(new_n1180));
  INV_X1    g0980(.A(new_n1180), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n1152), .A2(new_n1181), .ZN(G375));
  NAND2_X1  g0982(.A1(new_n1085), .A2(new_n1091), .ZN(new_n1183));
  NAND3_X1  g0983(.A1(new_n1093), .A2(new_n941), .A3(new_n1183), .ZN(new_n1184));
  OAI21_X1  g0984(.A(new_n719), .B1(G68), .B2(new_n825), .ZN(new_n1185));
  OAI221_X1 g0985(.A(new_n267), .B1(new_n454), .B2(new_n757), .C1(new_n733), .C2(new_n484), .ZN(new_n1186));
  AOI211_X1 g0986(.A(new_n1003), .B(new_n1186), .C1(G294), .C2(new_n805), .ZN(new_n1187));
  AOI22_X1  g0987(.A1(G107), .A2(new_n769), .B1(new_n771), .B2(G283), .ZN(new_n1188));
  NAND2_X1  g0988(.A1(new_n760), .A2(G303), .ZN(new_n1189));
  NAND4_X1  g0989(.A1(new_n1187), .A2(new_n985), .A3(new_n1188), .A4(new_n1189), .ZN(new_n1190));
  AOI21_X1  g0990(.A(new_n267), .B1(new_n732), .B2(new_n1105), .ZN(new_n1191));
  INV_X1    g0991(.A(G132), .ZN(new_n1192));
  OAI21_X1  g0992(.A(new_n1191), .B1(new_n1192), .B2(new_n735), .ZN(new_n1193));
  OAI22_X1  g0993(.A1(new_n349), .A2(new_n749), .B1(new_n747), .B2(new_n986), .ZN(new_n1194));
  AOI211_X1 g0994(.A(new_n1193), .B(new_n1194), .C1(G50), .C2(new_n743), .ZN(new_n1195));
  AOI22_X1  g0995(.A1(new_n760), .A2(G128), .B1(G159), .B2(new_n814), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(new_n1196), .A2(KEYINPUT122), .ZN(new_n1197));
  NAND3_X1  g0997(.A1(new_n1195), .A2(new_n1157), .A3(new_n1197), .ZN(new_n1198));
  NOR2_X1   g0998(.A1(new_n1196), .A2(KEYINPUT122), .ZN(new_n1199));
  OAI21_X1  g0999(.A(new_n1190), .B1(new_n1198), .B2(new_n1199), .ZN(new_n1200));
  AOI21_X1  g1000(.A(new_n1185), .B1(new_n1200), .B2(new_n727), .ZN(new_n1201));
  XNOR2_X1  g1001(.A(new_n1201), .B(KEYINPUT123), .ZN(new_n1202));
  AOI21_X1  g1002(.A(new_n1202), .B1(new_n710), .B2(new_n868), .ZN(new_n1203));
  INV_X1    g1003(.A(new_n1091), .ZN(new_n1204));
  AOI21_X1  g1004(.A(new_n1203), .B1(new_n1204), .B2(new_n718), .ZN(new_n1205));
  NAND2_X1  g1005(.A1(new_n1184), .A2(new_n1205), .ZN(G381));
  INV_X1    g1006(.A(G378), .ZN(new_n1207));
  AND3_X1   g1007(.A1(new_n1152), .A2(new_n1207), .A3(new_n1181), .ZN(new_n1208));
  AOI21_X1  g1008(.A(new_n1068), .B1(new_n1041), .B2(new_n1044), .ZN(new_n1209));
  OR2_X1    g1009(.A1(G393), .A2(G396), .ZN(new_n1210));
  NOR4_X1   g1010(.A1(new_n1210), .A2(G381), .A3(G384), .A4(G387), .ZN(new_n1211));
  NAND3_X1  g1011(.A1(new_n1208), .A2(new_n1209), .A3(new_n1211), .ZN(G407));
  AOI21_X1  g1012(.A(new_n1180), .B1(new_n1149), .B2(new_n1151), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(new_n1213), .A2(new_n1207), .ZN(new_n1214));
  OAI211_X1 g1014(.A(G407), .B(G213), .C1(new_n638), .C2(new_n1214), .ZN(G409));
  NOR2_X1   g1015(.A1(new_n638), .A2(new_n636), .ZN(new_n1216));
  NAND2_X1  g1016(.A1(new_n1135), .A2(new_n1139), .ZN(new_n1217));
  NAND2_X1  g1017(.A1(new_n1217), .A2(new_n718), .ZN(new_n1218));
  AND4_X1   g1018(.A1(new_n1096), .A2(new_n1218), .A3(new_n1121), .A4(new_n1179), .ZN(new_n1219));
  NAND4_X1  g1019(.A1(new_n1141), .A2(new_n1143), .A3(new_n1146), .A4(new_n941), .ZN(new_n1220));
  AOI21_X1  g1020(.A(new_n1216), .B1(new_n1219), .B2(new_n1220), .ZN(new_n1221));
  INV_X1    g1021(.A(G384), .ZN(new_n1222));
  INV_X1    g1022(.A(KEYINPUT60), .ZN(new_n1223));
  NAND2_X1  g1023(.A1(new_n1183), .A2(new_n1223), .ZN(new_n1224));
  NAND3_X1  g1024(.A1(new_n1085), .A2(new_n1091), .A3(KEYINPUT60), .ZN(new_n1225));
  NAND4_X1  g1025(.A1(new_n1224), .A2(new_n1093), .A3(new_n663), .A4(new_n1225), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n1226), .A2(new_n1205), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(new_n1222), .A2(new_n1227), .ZN(new_n1228));
  NAND3_X1  g1028(.A1(G384), .A2(new_n1205), .A3(new_n1226), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n1228), .A2(new_n1229), .ZN(new_n1230));
  INV_X1    g1030(.A(new_n1230), .ZN(new_n1231));
  OAI211_X1 g1031(.A(new_n1221), .B(new_n1231), .C1(new_n1213), .C2(new_n1207), .ZN(new_n1232));
  INV_X1    g1032(.A(KEYINPUT63), .ZN(new_n1233));
  OR2_X1    g1033(.A1(new_n1232), .A2(new_n1233), .ZN(new_n1234));
  XOR2_X1   g1034(.A(G393), .B(G396), .Z(new_n1235));
  NOR2_X1   g1035(.A1(new_n1209), .A2(G387), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n1209), .A2(G387), .ZN(new_n1237));
  INV_X1    g1037(.A(new_n1237), .ZN(new_n1238));
  NOR3_X1   g1038(.A1(new_n1235), .A2(new_n1236), .A3(new_n1238), .ZN(new_n1239));
  INV_X1    g1039(.A(KEYINPUT124), .ZN(new_n1240));
  NOR2_X1   g1040(.A1(new_n995), .A2(new_n967), .ZN(new_n1241));
  INV_X1    g1041(.A(new_n942), .ZN(new_n1242));
  AND2_X1   g1042(.A1(new_n961), .A2(new_n964), .ZN(new_n1243));
  AOI21_X1  g1043(.A(new_n1241), .B1(new_n1242), .B2(new_n1243), .ZN(new_n1244));
  NAND3_X1  g1044(.A1(G390), .A2(new_n1240), .A3(new_n1244), .ZN(new_n1245));
  OAI21_X1  g1045(.A(KEYINPUT124), .B1(new_n1209), .B2(G387), .ZN(new_n1246));
  NAND3_X1  g1046(.A1(new_n1245), .A2(new_n1246), .A3(new_n1237), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n1247), .A2(new_n1235), .ZN(new_n1248));
  INV_X1    g1048(.A(KEYINPUT125), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n1248), .A2(new_n1249), .ZN(new_n1250));
  NAND3_X1  g1050(.A1(new_n1247), .A2(KEYINPUT125), .A3(new_n1235), .ZN(new_n1251));
  AOI21_X1  g1051(.A(new_n1239), .B1(new_n1250), .B2(new_n1251), .ZN(new_n1252));
  INV_X1    g1052(.A(new_n1252), .ZN(new_n1253));
  OAI21_X1  g1053(.A(new_n1221), .B1(new_n1213), .B2(new_n1207), .ZN(new_n1254));
  NAND2_X1  g1054(.A1(new_n1216), .A2(G2897), .ZN(new_n1255));
  XNOR2_X1  g1055(.A(new_n1230), .B(new_n1255), .ZN(new_n1256));
  AOI21_X1  g1056(.A(KEYINPUT61), .B1(new_n1254), .B2(new_n1256), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(new_n1232), .A2(new_n1233), .ZN(new_n1258));
  NAND4_X1  g1058(.A1(new_n1234), .A2(new_n1253), .A3(new_n1257), .A4(new_n1258), .ZN(new_n1259));
  INV_X1    g1059(.A(KEYINPUT126), .ZN(new_n1260));
  NAND3_X1  g1060(.A1(new_n1232), .A2(new_n1260), .A3(KEYINPUT62), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(G375), .A2(G378), .ZN(new_n1262));
  XNOR2_X1  g1062(.A(KEYINPUT126), .B(KEYINPUT62), .ZN(new_n1263));
  NAND4_X1  g1063(.A1(new_n1262), .A2(new_n1221), .A3(new_n1231), .A4(new_n1263), .ZN(new_n1264));
  AND3_X1   g1064(.A1(new_n1261), .A2(new_n1257), .A3(new_n1264), .ZN(new_n1265));
  OAI21_X1  g1065(.A(new_n1259), .B1(new_n1265), .B2(new_n1253), .ZN(G405));
  AOI21_X1  g1066(.A(new_n1207), .B1(new_n1152), .B2(new_n1181), .ZN(new_n1267));
  OAI21_X1  g1067(.A(new_n1230), .B1(new_n1208), .B2(new_n1267), .ZN(new_n1268));
  NAND3_X1  g1068(.A1(new_n1262), .A2(new_n1214), .A3(new_n1231), .ZN(new_n1269));
  NAND3_X1  g1069(.A1(new_n1268), .A2(new_n1269), .A3(new_n1252), .ZN(new_n1270));
  NAND2_X1  g1070(.A1(new_n1270), .A2(KEYINPUT127), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(new_n1268), .A2(new_n1269), .ZN(new_n1272));
  NAND2_X1  g1072(.A1(new_n1272), .A2(new_n1253), .ZN(new_n1273));
  INV_X1    g1073(.A(KEYINPUT127), .ZN(new_n1274));
  NAND4_X1  g1074(.A1(new_n1268), .A2(new_n1269), .A3(new_n1252), .A4(new_n1274), .ZN(new_n1275));
  AND3_X1   g1075(.A1(new_n1271), .A2(new_n1273), .A3(new_n1275), .ZN(G402));
endmodule


