//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 1 1 1 1 0 0 1 0 1 1 1 1 1 0 1 1 1 1 0 1 1 1 0 1 1 1 1 0 0 1 1 1 0 0 0 0 1 0 0 0 1 1 1 0 1 1 1 1 1 1 0 0 1 0 0 0 1 0 1 0 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:21:40 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n711, new_n712, new_n713,
    new_n714, new_n716, new_n717, new_n718, new_n719, new_n720, new_n721,
    new_n722, new_n723, new_n724, new_n725, new_n726, new_n727, new_n728,
    new_n729, new_n730, new_n732, new_n733, new_n734, new_n735, new_n736,
    new_n737, new_n738, new_n739, new_n740, new_n741, new_n742, new_n743,
    new_n744, new_n745, new_n746, new_n747, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n777, new_n778, new_n779, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n800, new_n801, new_n802, new_n803,
    new_n804, new_n805, new_n806, new_n807, new_n808, new_n809, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n928, new_n929, new_n930, new_n931,
    new_n932, new_n933, new_n934, new_n935, new_n936, new_n937, new_n938,
    new_n939, new_n940, new_n941, new_n942, new_n943, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n957, new_n958, new_n959, new_n960, new_n962,
    new_n963, new_n964, new_n965, new_n966, new_n967, new_n969, new_n970,
    new_n971, new_n972, new_n973, new_n974, new_n975, new_n976, new_n977,
    new_n978, new_n979, new_n980, new_n981, new_n982, new_n984, new_n985,
    new_n986, new_n987, new_n988, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1021, new_n1022, new_n1023, new_n1024;
  NOR2_X1   g000(.A1(G237), .A2(G953), .ZN(new_n187));
  NAND2_X1  g001(.A1(new_n187), .A2(G210), .ZN(new_n188));
  INV_X1    g002(.A(G101), .ZN(new_n189));
  XNOR2_X1  g003(.A(new_n188), .B(new_n189), .ZN(new_n190));
  XNOR2_X1  g004(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n191));
  XOR2_X1   g005(.A(new_n190), .B(new_n191), .Z(new_n192));
  INV_X1    g006(.A(new_n192), .ZN(new_n193));
  INV_X1    g007(.A(G137), .ZN(new_n194));
  OAI21_X1  g008(.A(KEYINPUT65), .B1(new_n194), .B2(G134), .ZN(new_n195));
  INV_X1    g009(.A(KEYINPUT65), .ZN(new_n196));
  INV_X1    g010(.A(G134), .ZN(new_n197));
  NAND3_X1  g011(.A1(new_n196), .A2(new_n197), .A3(G137), .ZN(new_n198));
  AND2_X1   g012(.A1(new_n195), .A2(new_n198), .ZN(new_n199));
  INV_X1    g013(.A(KEYINPUT11), .ZN(new_n200));
  OAI21_X1  g014(.A(new_n200), .B1(new_n197), .B2(G137), .ZN(new_n201));
  NAND3_X1  g015(.A1(new_n194), .A2(KEYINPUT11), .A3(G134), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  OAI21_X1  g017(.A(G131), .B1(new_n199), .B2(new_n203), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n195), .A2(new_n198), .ZN(new_n205));
  INV_X1    g019(.A(G131), .ZN(new_n206));
  NAND4_X1  g020(.A1(new_n205), .A2(new_n206), .A3(new_n201), .A4(new_n202), .ZN(new_n207));
  NAND3_X1  g021(.A1(new_n204), .A2(KEYINPUT66), .A3(new_n207), .ZN(new_n208));
  XNOR2_X1  g022(.A(G143), .B(G146), .ZN(new_n209));
  NAND3_X1  g023(.A1(new_n209), .A2(KEYINPUT0), .A3(G128), .ZN(new_n210));
  NOR3_X1   g024(.A1(KEYINPUT64), .A2(KEYINPUT0), .A3(G128), .ZN(new_n211));
  OAI21_X1  g025(.A(KEYINPUT64), .B1(KEYINPUT0), .B2(G128), .ZN(new_n212));
  INV_X1    g026(.A(new_n212), .ZN(new_n213));
  NAND2_X1  g027(.A1(KEYINPUT0), .A2(G128), .ZN(new_n214));
  AOI21_X1  g028(.A(new_n211), .B1(new_n213), .B2(new_n214), .ZN(new_n215));
  OAI21_X1  g029(.A(new_n210), .B1(new_n215), .B2(new_n209), .ZN(new_n216));
  INV_X1    g030(.A(new_n216), .ZN(new_n217));
  INV_X1    g031(.A(KEYINPUT66), .ZN(new_n218));
  OAI211_X1 g032(.A(new_n218), .B(G131), .C1(new_n199), .C2(new_n203), .ZN(new_n219));
  NAND3_X1  g033(.A1(new_n208), .A2(new_n217), .A3(new_n219), .ZN(new_n220));
  INV_X1    g034(.A(G146), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n221), .A2(G143), .ZN(new_n222));
  INV_X1    g036(.A(G143), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n223), .A2(G146), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n222), .A2(new_n224), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n222), .A2(KEYINPUT1), .ZN(new_n226));
  NAND3_X1  g040(.A1(new_n225), .A2(new_n226), .A3(G128), .ZN(new_n227));
  INV_X1    g041(.A(G128), .ZN(new_n228));
  OAI211_X1 g042(.A(new_n222), .B(new_n224), .C1(KEYINPUT1), .C2(new_n228), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n227), .A2(new_n229), .ZN(new_n230));
  INV_X1    g044(.A(new_n230), .ZN(new_n231));
  NOR2_X1   g045(.A1(new_n194), .A2(G134), .ZN(new_n232));
  NOR2_X1   g046(.A1(new_n197), .A2(G137), .ZN(new_n233));
  OAI21_X1  g047(.A(G131), .B1(new_n232), .B2(new_n233), .ZN(new_n234));
  NAND3_X1  g048(.A1(new_n231), .A2(new_n207), .A3(new_n234), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n220), .A2(new_n235), .ZN(new_n236));
  INV_X1    g050(.A(KEYINPUT30), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n236), .A2(new_n237), .ZN(new_n238));
  OR2_X1    g052(.A1(KEYINPUT2), .A2(G113), .ZN(new_n239));
  NAND2_X1  g053(.A1(KEYINPUT2), .A2(G113), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n239), .A2(new_n240), .ZN(new_n241));
  INV_X1    g055(.A(G119), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n242), .A2(G116), .ZN(new_n243));
  INV_X1    g057(.A(G116), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n244), .A2(G119), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n243), .A2(new_n245), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n241), .A2(new_n246), .ZN(new_n247));
  NAND4_X1  g061(.A1(new_n239), .A2(new_n243), .A3(new_n245), .A4(new_n240), .ZN(new_n248));
  NAND3_X1  g062(.A1(new_n247), .A2(KEYINPUT67), .A3(new_n248), .ZN(new_n249));
  INV_X1    g063(.A(KEYINPUT67), .ZN(new_n250));
  NAND3_X1  g064(.A1(new_n241), .A2(new_n246), .A3(new_n250), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n249), .A2(new_n251), .ZN(new_n252));
  INV_X1    g066(.A(new_n252), .ZN(new_n253));
  NAND3_X1  g067(.A1(new_n220), .A2(KEYINPUT30), .A3(new_n235), .ZN(new_n254));
  AND3_X1   g068(.A1(new_n238), .A2(new_n253), .A3(new_n254), .ZN(new_n255));
  NAND3_X1  g069(.A1(new_n220), .A2(new_n252), .A3(new_n235), .ZN(new_n256));
  INV_X1    g070(.A(new_n256), .ZN(new_n257));
  OAI21_X1  g071(.A(new_n193), .B1(new_n255), .B2(new_n257), .ZN(new_n258));
  INV_X1    g072(.A(KEYINPUT28), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n256), .A2(new_n259), .ZN(new_n260));
  AOI21_X1  g074(.A(new_n252), .B1(new_n220), .B2(new_n235), .ZN(new_n261));
  NOR2_X1   g075(.A1(new_n257), .A2(new_n261), .ZN(new_n262));
  XNOR2_X1  g076(.A(KEYINPUT68), .B(KEYINPUT28), .ZN(new_n263));
  INV_X1    g077(.A(new_n263), .ZN(new_n264));
  OAI211_X1 g078(.A(new_n192), .B(new_n260), .C1(new_n262), .C2(new_n264), .ZN(new_n265));
  INV_X1    g079(.A(KEYINPUT29), .ZN(new_n266));
  NAND3_X1  g080(.A1(new_n258), .A2(new_n265), .A3(new_n266), .ZN(new_n267));
  INV_X1    g081(.A(new_n260), .ZN(new_n268));
  OAI21_X1  g082(.A(KEYINPUT28), .B1(new_n257), .B2(new_n261), .ZN(new_n269));
  AOI21_X1  g083(.A(new_n268), .B1(new_n269), .B2(KEYINPUT70), .ZN(new_n270));
  INV_X1    g084(.A(KEYINPUT70), .ZN(new_n271));
  OAI211_X1 g085(.A(new_n271), .B(KEYINPUT28), .C1(new_n257), .C2(new_n261), .ZN(new_n272));
  NAND4_X1  g086(.A1(new_n270), .A2(KEYINPUT29), .A3(new_n192), .A4(new_n272), .ZN(new_n273));
  INV_X1    g087(.A(G902), .ZN(new_n274));
  NAND3_X1  g088(.A1(new_n267), .A2(new_n273), .A3(new_n274), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n275), .A2(G472), .ZN(new_n276));
  NAND3_X1  g090(.A1(new_n238), .A2(new_n253), .A3(new_n254), .ZN(new_n277));
  NAND3_X1  g091(.A1(new_n277), .A2(new_n192), .A3(new_n256), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n278), .A2(KEYINPUT31), .ZN(new_n279));
  INV_X1    g093(.A(new_n261), .ZN(new_n280));
  AOI21_X1  g094(.A(new_n264), .B1(new_n280), .B2(new_n256), .ZN(new_n281));
  OAI21_X1  g095(.A(new_n193), .B1(new_n281), .B2(new_n268), .ZN(new_n282));
  INV_X1    g096(.A(KEYINPUT31), .ZN(new_n283));
  NAND4_X1  g097(.A1(new_n277), .A2(new_n283), .A3(new_n192), .A4(new_n256), .ZN(new_n284));
  NAND3_X1  g098(.A1(new_n279), .A2(new_n282), .A3(new_n284), .ZN(new_n285));
  NOR2_X1   g099(.A1(G472), .A2(G902), .ZN(new_n286));
  XNOR2_X1  g100(.A(new_n286), .B(KEYINPUT69), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n285), .A2(new_n287), .ZN(new_n288));
  INV_X1    g102(.A(KEYINPUT32), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  NAND3_X1  g104(.A1(new_n285), .A2(KEYINPUT32), .A3(new_n287), .ZN(new_n291));
  NAND3_X1  g105(.A1(new_n276), .A2(new_n290), .A3(new_n291), .ZN(new_n292));
  XNOR2_X1  g106(.A(KEYINPUT22), .B(G137), .ZN(new_n293));
  INV_X1    g107(.A(G221), .ZN(new_n294));
  INV_X1    g108(.A(G234), .ZN(new_n295));
  NOR3_X1   g109(.A1(new_n294), .A2(new_n295), .A3(G953), .ZN(new_n296));
  XOR2_X1   g110(.A(new_n293), .B(new_n296), .Z(new_n297));
  INV_X1    g111(.A(new_n297), .ZN(new_n298));
  INV_X1    g112(.A(G140), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n299), .A2(G125), .ZN(new_n300));
  INV_X1    g114(.A(G125), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n301), .A2(G140), .ZN(new_n302));
  NAND3_X1  g116(.A1(new_n300), .A2(new_n302), .A3(new_n221), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n303), .A2(KEYINPUT75), .ZN(new_n304));
  XNOR2_X1  g118(.A(G125), .B(G140), .ZN(new_n305));
  INV_X1    g119(.A(KEYINPUT75), .ZN(new_n306));
  NAND3_X1  g120(.A1(new_n305), .A2(new_n306), .A3(new_n221), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n304), .A2(new_n307), .ZN(new_n308));
  NAND3_X1  g122(.A1(new_n300), .A2(new_n302), .A3(KEYINPUT16), .ZN(new_n309));
  OR3_X1    g123(.A1(new_n301), .A2(KEYINPUT16), .A3(G140), .ZN(new_n310));
  NAND3_X1  g124(.A1(new_n309), .A2(new_n310), .A3(G146), .ZN(new_n311));
  AND2_X1   g125(.A1(new_n308), .A2(new_n311), .ZN(new_n312));
  XOR2_X1   g126(.A(KEYINPUT73), .B(G110), .Z(new_n313));
  OAI21_X1  g127(.A(KEYINPUT23), .B1(new_n228), .B2(G119), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n314), .A2(KEYINPUT71), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n242), .A2(G128), .ZN(new_n316));
  INV_X1    g130(.A(KEYINPUT71), .ZN(new_n317));
  NAND3_X1  g131(.A1(new_n316), .A2(new_n317), .A3(KEYINPUT23), .ZN(new_n318));
  NAND3_X1  g132(.A1(new_n315), .A2(KEYINPUT72), .A3(new_n318), .ZN(new_n319));
  NOR2_X1   g133(.A1(new_n242), .A2(G128), .ZN(new_n320));
  INV_X1    g134(.A(new_n320), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n319), .A2(new_n321), .ZN(new_n322));
  INV_X1    g136(.A(KEYINPUT23), .ZN(new_n323));
  OAI211_X1 g137(.A(new_n320), .B(new_n323), .C1(KEYINPUT71), .C2(KEYINPUT72), .ZN(new_n324));
  AOI21_X1  g138(.A(new_n313), .B1(new_n322), .B2(new_n324), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n321), .A2(new_n316), .ZN(new_n326));
  XNOR2_X1  g140(.A(KEYINPUT24), .B(G110), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n326), .A2(new_n327), .ZN(new_n328));
  INV_X1    g142(.A(KEYINPUT74), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n328), .A2(new_n329), .ZN(new_n330));
  NAND3_X1  g144(.A1(new_n326), .A2(new_n327), .A3(KEYINPUT74), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n330), .A2(new_n331), .ZN(new_n332));
  OAI21_X1  g146(.A(new_n312), .B1(new_n325), .B2(new_n332), .ZN(new_n333));
  INV_X1    g147(.A(KEYINPUT76), .ZN(new_n334));
  NAND3_X1  g148(.A1(new_n322), .A2(G110), .A3(new_n324), .ZN(new_n335));
  NOR2_X1   g149(.A1(new_n326), .A2(new_n327), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n309), .A2(new_n310), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n337), .A2(new_n221), .ZN(new_n338));
  AOI21_X1  g152(.A(new_n336), .B1(new_n338), .B2(new_n311), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n335), .A2(new_n339), .ZN(new_n340));
  AND3_X1   g154(.A1(new_n333), .A2(new_n334), .A3(new_n340), .ZN(new_n341));
  AOI21_X1  g155(.A(new_n334), .B1(new_n333), .B2(new_n340), .ZN(new_n342));
  OAI21_X1  g156(.A(new_n298), .B1(new_n341), .B2(new_n342), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n333), .A2(new_n340), .ZN(new_n344));
  NOR2_X1   g158(.A1(new_n344), .A2(new_n298), .ZN(new_n345));
  INV_X1    g159(.A(new_n345), .ZN(new_n346));
  NAND3_X1  g160(.A1(new_n343), .A2(new_n274), .A3(new_n346), .ZN(new_n347));
  INV_X1    g161(.A(KEYINPUT25), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n347), .A2(new_n348), .ZN(new_n349));
  NAND4_X1  g163(.A1(new_n343), .A2(KEYINPUT25), .A3(new_n346), .A4(new_n274), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n349), .A2(new_n350), .ZN(new_n351));
  INV_X1    g165(.A(G217), .ZN(new_n352));
  AOI21_X1  g166(.A(new_n352), .B1(G234), .B2(new_n274), .ZN(new_n353));
  NOR2_X1   g167(.A1(new_n353), .A2(G902), .ZN(new_n354));
  XNOR2_X1  g168(.A(new_n354), .B(KEYINPUT77), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n344), .A2(KEYINPUT76), .ZN(new_n356));
  NAND3_X1  g170(.A1(new_n333), .A2(new_n334), .A3(new_n340), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  AOI21_X1  g172(.A(new_n345), .B1(new_n358), .B2(new_n298), .ZN(new_n359));
  AOI22_X1  g173(.A1(new_n351), .A2(new_n353), .B1(new_n355), .B2(new_n359), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n292), .A2(new_n360), .ZN(new_n361));
  NOR2_X1   g175(.A1(new_n361), .A2(KEYINPUT78), .ZN(new_n362));
  INV_X1    g176(.A(KEYINPUT78), .ZN(new_n363));
  AOI21_X1  g177(.A(new_n363), .B1(new_n292), .B2(new_n360), .ZN(new_n364));
  NOR2_X1   g178(.A1(new_n362), .A2(new_n364), .ZN(new_n365));
  INV_X1    g179(.A(KEYINPUT3), .ZN(new_n366));
  INV_X1    g180(.A(G107), .ZN(new_n367));
  NAND3_X1  g181(.A1(new_n366), .A2(new_n367), .A3(G104), .ZN(new_n368));
  INV_X1    g182(.A(G104), .ZN(new_n369));
  AOI21_X1  g183(.A(KEYINPUT3), .B1(new_n369), .B2(G107), .ZN(new_n370));
  NOR2_X1   g184(.A1(new_n369), .A2(G107), .ZN(new_n371));
  OAI211_X1 g185(.A(new_n189), .B(new_n368), .C1(new_n370), .C2(new_n371), .ZN(new_n372));
  NOR2_X1   g186(.A1(new_n367), .A2(G104), .ZN(new_n373));
  OAI21_X1  g187(.A(G101), .B1(new_n371), .B2(new_n373), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n372), .A2(new_n374), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n230), .A2(new_n375), .ZN(new_n376));
  NAND4_X1  g190(.A1(new_n227), .A2(new_n372), .A3(new_n229), .A4(new_n374), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n376), .A2(new_n377), .ZN(new_n378));
  NAND3_X1  g192(.A1(new_n378), .A2(new_n219), .A3(new_n208), .ZN(new_n379));
  INV_X1    g193(.A(KEYINPUT12), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n379), .A2(new_n380), .ZN(new_n381));
  AND2_X1   g195(.A1(new_n208), .A2(new_n219), .ZN(new_n382));
  NAND3_X1  g196(.A1(new_n382), .A2(KEYINPUT12), .A3(new_n378), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n381), .A2(new_n383), .ZN(new_n384));
  INV_X1    g198(.A(KEYINPUT81), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n384), .A2(new_n385), .ZN(new_n386));
  XNOR2_X1  g200(.A(G110), .B(G140), .ZN(new_n387));
  INV_X1    g201(.A(G227), .ZN(new_n388));
  NOR2_X1   g202(.A1(new_n388), .A2(G953), .ZN(new_n389));
  XOR2_X1   g203(.A(new_n387), .B(new_n389), .Z(new_n390));
  INV_X1    g204(.A(new_n390), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n208), .A2(new_n219), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n392), .A2(KEYINPUT80), .ZN(new_n393));
  INV_X1    g207(.A(KEYINPUT80), .ZN(new_n394));
  NAND3_X1  g208(.A1(new_n208), .A2(new_n394), .A3(new_n219), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n393), .A2(new_n395), .ZN(new_n396));
  INV_X1    g210(.A(new_n375), .ZN(new_n397));
  NAND3_X1  g211(.A1(new_n231), .A2(new_n397), .A3(KEYINPUT10), .ZN(new_n398));
  INV_X1    g212(.A(KEYINPUT10), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n377), .A2(new_n399), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n398), .A2(new_n400), .ZN(new_n401));
  INV_X1    g215(.A(KEYINPUT79), .ZN(new_n402));
  NAND3_X1  g216(.A1(new_n372), .A2(new_n402), .A3(KEYINPUT4), .ZN(new_n403));
  OAI21_X1  g217(.A(new_n368), .B1(new_n370), .B2(new_n371), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n404), .A2(G101), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n403), .A2(new_n405), .ZN(new_n406));
  NAND4_X1  g220(.A1(new_n404), .A2(new_n402), .A3(KEYINPUT4), .A4(G101), .ZN(new_n407));
  AOI21_X1  g221(.A(new_n216), .B1(new_n406), .B2(new_n407), .ZN(new_n408));
  NOR2_X1   g222(.A1(new_n401), .A2(new_n408), .ZN(new_n409));
  AOI21_X1  g223(.A(new_n391), .B1(new_n396), .B2(new_n409), .ZN(new_n410));
  NAND3_X1  g224(.A1(new_n381), .A2(new_n383), .A3(KEYINPUT81), .ZN(new_n411));
  NAND3_X1  g225(.A1(new_n386), .A2(new_n410), .A3(new_n411), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n396), .A2(new_n409), .ZN(new_n413));
  OAI21_X1  g227(.A(new_n382), .B1(new_n401), .B2(new_n408), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n413), .A2(new_n414), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n415), .A2(new_n391), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n412), .A2(new_n416), .ZN(new_n417));
  INV_X1    g231(.A(G469), .ZN(new_n418));
  NAND3_X1  g232(.A1(new_n417), .A2(new_n418), .A3(new_n274), .ZN(new_n419));
  NAND2_X1  g233(.A1(G469), .A2(G902), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n413), .A2(new_n384), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n421), .A2(new_n391), .ZN(new_n422));
  NAND3_X1  g236(.A1(new_n413), .A2(new_n414), .A3(new_n390), .ZN(new_n423));
  NAND3_X1  g237(.A1(new_n422), .A2(G469), .A3(new_n423), .ZN(new_n424));
  NAND3_X1  g238(.A1(new_n419), .A2(new_n420), .A3(new_n424), .ZN(new_n425));
  XOR2_X1   g239(.A(KEYINPUT9), .B(G234), .Z(new_n426));
  AOI21_X1  g240(.A(new_n294), .B1(new_n426), .B2(new_n274), .ZN(new_n427));
  INV_X1    g241(.A(new_n427), .ZN(new_n428));
  AND2_X1   g242(.A1(new_n425), .A2(new_n428), .ZN(new_n429));
  OAI21_X1  g243(.A(G214), .B1(G237), .B2(G902), .ZN(new_n430));
  AOI21_X1  g244(.A(new_n252), .B1(new_n406), .B2(new_n407), .ZN(new_n431));
  NAND3_X1  g245(.A1(new_n243), .A2(new_n245), .A3(KEYINPUT5), .ZN(new_n432));
  OAI211_X1 g246(.A(new_n432), .B(G113), .C1(KEYINPUT5), .C2(new_n243), .ZN(new_n433));
  AND4_X1   g247(.A1(new_n248), .A2(new_n433), .A3(new_n372), .A4(new_n374), .ZN(new_n434));
  XNOR2_X1  g248(.A(G110), .B(G122), .ZN(new_n435));
  INV_X1    g249(.A(new_n435), .ZN(new_n436));
  NOR3_X1   g250(.A1(new_n431), .A2(new_n434), .A3(new_n436), .ZN(new_n437));
  XNOR2_X1  g251(.A(new_n435), .B(KEYINPUT8), .ZN(new_n438));
  AOI22_X1  g252(.A1(new_n433), .A2(new_n248), .B1(new_n372), .B2(new_n374), .ZN(new_n439));
  OAI21_X1  g253(.A(new_n438), .B1(new_n434), .B2(new_n439), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n216), .A2(G125), .ZN(new_n441));
  AOI21_X1  g255(.A(G125), .B1(new_n227), .B2(new_n229), .ZN(new_n442));
  INV_X1    g256(.A(new_n442), .ZN(new_n443));
  INV_X1    g257(.A(G224), .ZN(new_n444));
  NOR2_X1   g258(.A1(new_n444), .A2(G953), .ZN(new_n445));
  INV_X1    g259(.A(new_n445), .ZN(new_n446));
  NAND4_X1  g260(.A1(new_n441), .A2(new_n443), .A3(KEYINPUT7), .A4(new_n446), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n440), .A2(new_n447), .ZN(new_n448));
  NOR2_X1   g262(.A1(new_n437), .A2(new_n448), .ZN(new_n449));
  INV_X1    g263(.A(KEYINPUT84), .ZN(new_n450));
  INV_X1    g264(.A(KEYINPUT7), .ZN(new_n451));
  AOI21_X1  g265(.A(new_n445), .B1(new_n450), .B2(new_n451), .ZN(new_n452));
  OAI21_X1  g266(.A(new_n452), .B1(new_n450), .B2(new_n451), .ZN(new_n453));
  INV_X1    g267(.A(KEYINPUT83), .ZN(new_n454));
  AOI21_X1  g268(.A(new_n454), .B1(new_n441), .B2(new_n443), .ZN(new_n455));
  NOR2_X1   g269(.A1(new_n442), .A2(KEYINPUT83), .ZN(new_n456));
  OAI21_X1  g270(.A(new_n453), .B1(new_n455), .B2(new_n456), .ZN(new_n457));
  AOI21_X1  g271(.A(G902), .B1(new_n449), .B2(new_n457), .ZN(new_n458));
  AOI21_X1  g272(.A(new_n212), .B1(KEYINPUT0), .B2(G128), .ZN(new_n459));
  OAI21_X1  g273(.A(new_n225), .B1(new_n459), .B2(new_n211), .ZN(new_n460));
  AOI21_X1  g274(.A(new_n301), .B1(new_n460), .B2(new_n210), .ZN(new_n461));
  OAI21_X1  g275(.A(new_n445), .B1(new_n461), .B2(new_n442), .ZN(new_n462));
  NAND3_X1  g276(.A1(new_n441), .A2(new_n443), .A3(new_n446), .ZN(new_n463));
  AND3_X1   g277(.A1(new_n462), .A2(new_n463), .A3(KEYINPUT82), .ZN(new_n464));
  AOI21_X1  g278(.A(KEYINPUT82), .B1(new_n462), .B2(new_n463), .ZN(new_n465));
  NOR2_X1   g279(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  INV_X1    g280(.A(new_n434), .ZN(new_n467));
  AND2_X1   g281(.A1(new_n406), .A2(new_n407), .ZN(new_n468));
  OAI211_X1 g282(.A(new_n467), .B(new_n435), .C1(new_n468), .C2(new_n252), .ZN(new_n469));
  OAI21_X1  g283(.A(new_n436), .B1(new_n431), .B2(new_n434), .ZN(new_n470));
  NAND3_X1  g284(.A1(new_n469), .A2(new_n470), .A3(KEYINPUT6), .ZN(new_n471));
  INV_X1    g285(.A(KEYINPUT6), .ZN(new_n472));
  OAI211_X1 g286(.A(new_n472), .B(new_n436), .C1(new_n431), .C2(new_n434), .ZN(new_n473));
  NAND3_X1  g287(.A1(new_n466), .A2(new_n471), .A3(new_n473), .ZN(new_n474));
  OAI21_X1  g288(.A(G210), .B1(G237), .B2(G902), .ZN(new_n475));
  AND3_X1   g289(.A1(new_n458), .A2(new_n474), .A3(new_n475), .ZN(new_n476));
  AOI21_X1  g290(.A(new_n475), .B1(new_n458), .B2(new_n474), .ZN(new_n477));
  OAI21_X1  g291(.A(new_n430), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  INV_X1    g292(.A(KEYINPUT85), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  OAI211_X1 g294(.A(KEYINPUT85), .B(new_n430), .C1(new_n476), .C2(new_n477), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  INV_X1    g296(.A(KEYINPUT89), .ZN(new_n483));
  NOR2_X1   g297(.A1(G475), .A2(G902), .ZN(new_n484));
  INV_X1    g298(.A(new_n484), .ZN(new_n485));
  INV_X1    g299(.A(KEYINPUT87), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n300), .A2(new_n302), .ZN(new_n487));
  XNOR2_X1  g301(.A(new_n487), .B(KEYINPUT19), .ZN(new_n488));
  OAI21_X1  g302(.A(new_n486), .B1(new_n488), .B2(G146), .ZN(new_n489));
  INV_X1    g303(.A(new_n311), .ZN(new_n490));
  NAND3_X1  g304(.A1(new_n187), .A2(G143), .A3(G214), .ZN(new_n491));
  INV_X1    g305(.A(new_n491), .ZN(new_n492));
  AOI21_X1  g306(.A(G143), .B1(new_n187), .B2(G214), .ZN(new_n493));
  OAI21_X1  g307(.A(G131), .B1(new_n492), .B2(new_n493), .ZN(new_n494));
  INV_X1    g308(.A(new_n493), .ZN(new_n495));
  NAND3_X1  g309(.A1(new_n495), .A2(new_n206), .A3(new_n491), .ZN(new_n496));
  AOI21_X1  g310(.A(new_n490), .B1(new_n494), .B2(new_n496), .ZN(new_n497));
  XNOR2_X1  g311(.A(new_n305), .B(KEYINPUT19), .ZN(new_n498));
  NAND3_X1  g312(.A1(new_n498), .A2(KEYINPUT87), .A3(new_n221), .ZN(new_n499));
  NAND3_X1  g313(.A1(new_n489), .A2(new_n497), .A3(new_n499), .ZN(new_n500));
  INV_X1    g314(.A(KEYINPUT86), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n487), .A2(G146), .ZN(new_n502));
  NOR2_X1   g316(.A1(new_n492), .A2(new_n493), .ZN(new_n503));
  NAND2_X1  g317(.A1(KEYINPUT18), .A2(G131), .ZN(new_n504));
  AOI22_X1  g318(.A1(new_n308), .A2(new_n502), .B1(new_n503), .B2(new_n504), .ZN(new_n505));
  OAI211_X1 g319(.A(KEYINPUT18), .B(G131), .C1(new_n492), .C2(new_n493), .ZN(new_n506));
  AOI21_X1  g320(.A(new_n501), .B1(new_n505), .B2(new_n506), .ZN(new_n507));
  AOI21_X1  g321(.A(new_n306), .B1(new_n305), .B2(new_n221), .ZN(new_n508));
  AND4_X1   g322(.A1(new_n306), .A2(new_n300), .A3(new_n302), .A4(new_n221), .ZN(new_n509));
  OAI21_X1  g323(.A(new_n502), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n503), .A2(new_n504), .ZN(new_n511));
  AND4_X1   g325(.A1(new_n501), .A2(new_n510), .A3(new_n511), .A4(new_n506), .ZN(new_n512));
  OAI21_X1  g326(.A(new_n500), .B1(new_n507), .B2(new_n512), .ZN(new_n513));
  XNOR2_X1  g327(.A(G113), .B(G122), .ZN(new_n514));
  XNOR2_X1  g328(.A(new_n514), .B(new_n369), .ZN(new_n515));
  INV_X1    g329(.A(new_n515), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n513), .A2(new_n516), .ZN(new_n517));
  INV_X1    g331(.A(KEYINPUT17), .ZN(new_n518));
  OR2_X1    g332(.A1(new_n494), .A2(new_n518), .ZN(new_n519));
  INV_X1    g333(.A(KEYINPUT88), .ZN(new_n520));
  AOI21_X1  g334(.A(G146), .B1(new_n309), .B2(new_n310), .ZN(new_n521));
  OAI21_X1  g335(.A(new_n520), .B1(new_n490), .B2(new_n521), .ZN(new_n522));
  NAND3_X1  g336(.A1(new_n338), .A2(KEYINPUT88), .A3(new_n311), .ZN(new_n523));
  NAND3_X1  g337(.A1(new_n494), .A2(new_n496), .A3(new_n518), .ZN(new_n524));
  NAND4_X1  g338(.A1(new_n519), .A2(new_n522), .A3(new_n523), .A4(new_n524), .ZN(new_n525));
  OAI211_X1 g339(.A(new_n525), .B(new_n515), .C1(new_n507), .C2(new_n512), .ZN(new_n526));
  AOI21_X1  g340(.A(new_n485), .B1(new_n517), .B2(new_n526), .ZN(new_n527));
  INV_X1    g341(.A(KEYINPUT20), .ZN(new_n528));
  OAI21_X1  g342(.A(new_n483), .B1(new_n527), .B2(new_n528), .ZN(new_n529));
  INV_X1    g343(.A(new_n526), .ZN(new_n530));
  NAND3_X1  g344(.A1(new_n510), .A2(new_n511), .A3(new_n506), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n531), .A2(KEYINPUT86), .ZN(new_n532));
  NAND4_X1  g346(.A1(new_n510), .A2(new_n511), .A3(new_n501), .A4(new_n506), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  AOI21_X1  g348(.A(new_n515), .B1(new_n534), .B2(new_n500), .ZN(new_n535));
  OAI21_X1  g349(.A(new_n484), .B1(new_n530), .B2(new_n535), .ZN(new_n536));
  NAND3_X1  g350(.A1(new_n536), .A2(KEYINPUT89), .A3(KEYINPUT20), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n517), .A2(new_n526), .ZN(new_n538));
  XNOR2_X1  g352(.A(new_n484), .B(KEYINPUT90), .ZN(new_n539));
  NAND3_X1  g353(.A1(new_n538), .A2(new_n528), .A3(new_n539), .ZN(new_n540));
  NAND3_X1  g354(.A1(new_n529), .A2(new_n537), .A3(new_n540), .ZN(new_n541));
  AOI21_X1  g355(.A(new_n515), .B1(new_n534), .B2(new_n525), .ZN(new_n542));
  OAI21_X1  g356(.A(new_n274), .B1(new_n530), .B2(new_n542), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n543), .A2(G475), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n541), .A2(new_n544), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n228), .A2(G143), .ZN(new_n546));
  INV_X1    g360(.A(KEYINPUT93), .ZN(new_n547));
  XNOR2_X1  g361(.A(new_n546), .B(new_n547), .ZN(new_n548));
  OAI21_X1  g362(.A(KEYINPUT91), .B1(new_n228), .B2(G143), .ZN(new_n549));
  INV_X1    g363(.A(KEYINPUT91), .ZN(new_n550));
  NAND3_X1  g364(.A1(new_n550), .A2(new_n223), .A3(G128), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n549), .A2(new_n551), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n548), .A2(new_n552), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n553), .A2(G134), .ZN(new_n554));
  NAND3_X1  g368(.A1(new_n548), .A2(new_n197), .A3(new_n552), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  INV_X1    g370(.A(G122), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n557), .A2(G116), .ZN(new_n558));
  AOI21_X1  g372(.A(new_n367), .B1(new_n558), .B2(KEYINPUT14), .ZN(new_n559));
  XNOR2_X1  g373(.A(G116), .B(G122), .ZN(new_n560));
  XOR2_X1   g374(.A(new_n559), .B(new_n560), .Z(new_n561));
  INV_X1    g375(.A(new_n561), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n556), .A2(new_n562), .ZN(new_n563));
  INV_X1    g377(.A(G953), .ZN(new_n564));
  NAND3_X1  g378(.A1(new_n426), .A2(G217), .A3(new_n564), .ZN(new_n565));
  INV_X1    g379(.A(new_n565), .ZN(new_n566));
  INV_X1    g380(.A(new_n548), .ZN(new_n567));
  INV_X1    g381(.A(KEYINPUT92), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n552), .A2(new_n568), .ZN(new_n569));
  NAND3_X1  g383(.A1(new_n549), .A2(new_n551), .A3(KEYINPUT92), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  AOI21_X1  g385(.A(new_n567), .B1(new_n571), .B2(KEYINPUT13), .ZN(new_n572));
  INV_X1    g386(.A(KEYINPUT13), .ZN(new_n573));
  NAND3_X1  g387(.A1(new_n569), .A2(new_n573), .A3(new_n570), .ZN(new_n574));
  AOI21_X1  g388(.A(new_n197), .B1(new_n572), .B2(new_n574), .ZN(new_n575));
  XNOR2_X1  g389(.A(new_n560), .B(new_n367), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n555), .A2(new_n576), .ZN(new_n577));
  OAI211_X1 g391(.A(new_n563), .B(new_n566), .C1(new_n575), .C2(new_n577), .ZN(new_n578));
  AND3_X1   g392(.A1(new_n549), .A2(new_n551), .A3(KEYINPUT92), .ZN(new_n579));
  AOI21_X1  g393(.A(KEYINPUT92), .B1(new_n549), .B2(new_n551), .ZN(new_n580));
  OAI21_X1  g394(.A(KEYINPUT13), .B1(new_n579), .B2(new_n580), .ZN(new_n581));
  NAND3_X1  g395(.A1(new_n581), .A2(new_n574), .A3(new_n548), .ZN(new_n582));
  AOI21_X1  g396(.A(new_n577), .B1(new_n582), .B2(G134), .ZN(new_n583));
  AOI21_X1  g397(.A(new_n561), .B1(new_n554), .B2(new_n555), .ZN(new_n584));
  OAI21_X1  g398(.A(new_n565), .B1(new_n583), .B2(new_n584), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n578), .A2(new_n585), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n586), .A2(new_n274), .ZN(new_n587));
  INV_X1    g401(.A(G478), .ZN(new_n588));
  NOR2_X1   g402(.A1(KEYINPUT94), .A2(KEYINPUT15), .ZN(new_n589));
  INV_X1    g403(.A(new_n589), .ZN(new_n590));
  NAND2_X1  g404(.A1(KEYINPUT94), .A2(KEYINPUT15), .ZN(new_n591));
  AOI21_X1  g405(.A(new_n588), .B1(new_n590), .B2(new_n591), .ZN(new_n592));
  INV_X1    g406(.A(new_n592), .ZN(new_n593));
  NAND3_X1  g407(.A1(new_n587), .A2(KEYINPUT95), .A3(new_n593), .ZN(new_n594));
  AOI21_X1  g408(.A(G902), .B1(new_n578), .B2(new_n585), .ZN(new_n595));
  INV_X1    g409(.A(KEYINPUT95), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  INV_X1    g411(.A(new_n597), .ZN(new_n598));
  OAI21_X1  g412(.A(new_n592), .B1(new_n595), .B2(new_n596), .ZN(new_n599));
  OAI21_X1  g413(.A(new_n594), .B1(new_n598), .B2(new_n599), .ZN(new_n600));
  INV_X1    g414(.A(new_n600), .ZN(new_n601));
  INV_X1    g415(.A(G952), .ZN(new_n602));
  NOR2_X1   g416(.A1(new_n602), .A2(G953), .ZN(new_n603));
  INV_X1    g417(.A(G237), .ZN(new_n604));
  OAI21_X1  g418(.A(new_n603), .B1(new_n295), .B2(new_n604), .ZN(new_n605));
  INV_X1    g419(.A(new_n605), .ZN(new_n606));
  OAI211_X1 g420(.A(G902), .B(G953), .C1(new_n295), .C2(new_n604), .ZN(new_n607));
  XOR2_X1   g421(.A(new_n607), .B(KEYINPUT96), .Z(new_n608));
  XNOR2_X1  g422(.A(KEYINPUT21), .B(G898), .ZN(new_n609));
  AOI21_X1  g423(.A(new_n606), .B1(new_n608), .B2(new_n609), .ZN(new_n610));
  NOR3_X1   g424(.A1(new_n545), .A2(new_n601), .A3(new_n610), .ZN(new_n611));
  AND3_X1   g425(.A1(new_n429), .A2(new_n482), .A3(new_n611), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n365), .A2(new_n612), .ZN(new_n613));
  XNOR2_X1  g427(.A(new_n613), .B(G101), .ZN(G3));
  AND3_X1   g428(.A1(new_n360), .A2(new_n428), .A3(new_n425), .ZN(new_n615));
  AND3_X1   g429(.A1(new_n578), .A2(new_n585), .A3(KEYINPUT33), .ZN(new_n616));
  AOI21_X1  g430(.A(KEYINPUT33), .B1(new_n578), .B2(new_n585), .ZN(new_n617));
  NOR2_X1   g431(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  NOR2_X1   g432(.A1(new_n588), .A2(G902), .ZN(new_n619));
  AOI22_X1  g433(.A1(new_n618), .A2(new_n619), .B1(new_n588), .B2(new_n587), .ZN(new_n620));
  INV_X1    g434(.A(new_n620), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n545), .A2(new_n621), .ZN(new_n622));
  INV_X1    g436(.A(new_n430), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n458), .A2(new_n474), .ZN(new_n624));
  INV_X1    g438(.A(new_n475), .ZN(new_n625));
  NAND2_X1  g439(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  NAND3_X1  g440(.A1(new_n458), .A2(new_n474), .A3(new_n475), .ZN(new_n627));
  AOI21_X1  g441(.A(new_n623), .B1(new_n626), .B2(new_n627), .ZN(new_n628));
  INV_X1    g442(.A(new_n610), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  NOR2_X1   g444(.A1(new_n622), .A2(new_n630), .ZN(new_n631));
  INV_X1    g445(.A(G472), .ZN(new_n632));
  AOI21_X1  g446(.A(new_n632), .B1(new_n285), .B2(new_n274), .ZN(new_n633));
  AOI21_X1  g447(.A(new_n633), .B1(new_n285), .B2(new_n287), .ZN(new_n634));
  NAND3_X1  g448(.A1(new_n615), .A2(new_n631), .A3(new_n634), .ZN(new_n635));
  XOR2_X1   g449(.A(KEYINPUT34), .B(G104), .Z(new_n636));
  XNOR2_X1  g450(.A(new_n635), .B(new_n636), .ZN(G6));
  NAND2_X1  g451(.A1(new_n615), .A2(new_n634), .ZN(new_n638));
  NAND3_X1  g452(.A1(new_n538), .A2(new_n528), .A3(new_n484), .ZN(new_n639));
  NAND3_X1  g453(.A1(new_n529), .A2(new_n537), .A3(new_n639), .ZN(new_n640));
  AND2_X1   g454(.A1(new_n640), .A2(new_n544), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n641), .A2(new_n601), .ZN(new_n642));
  NOR3_X1   g456(.A1(new_n638), .A2(new_n630), .A3(new_n642), .ZN(new_n643));
  XNOR2_X1  g457(.A(KEYINPUT35), .B(G107), .ZN(new_n644));
  XNOR2_X1  g458(.A(new_n643), .B(new_n644), .ZN(G9));
  NAND2_X1  g459(.A1(new_n351), .A2(new_n353), .ZN(new_n646));
  NOR2_X1   g460(.A1(new_n298), .A2(KEYINPUT36), .ZN(new_n647));
  XNOR2_X1  g461(.A(new_n358), .B(new_n647), .ZN(new_n648));
  NAND2_X1  g462(.A1(new_n648), .A2(new_n355), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n646), .A2(new_n649), .ZN(new_n650));
  INV_X1    g464(.A(new_n633), .ZN(new_n651));
  AND3_X1   g465(.A1(new_n650), .A2(new_n288), .A3(new_n651), .ZN(new_n652));
  NAND2_X1  g466(.A1(new_n612), .A2(new_n652), .ZN(new_n653));
  XOR2_X1   g467(.A(KEYINPUT37), .B(G110), .Z(new_n654));
  XNOR2_X1  g468(.A(new_n653), .B(new_n654), .ZN(G12));
  NAND3_X1  g469(.A1(new_n292), .A2(new_n429), .A3(new_n650), .ZN(new_n656));
  INV_X1    g470(.A(G900), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n608), .A2(new_n657), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n658), .A2(new_n605), .ZN(new_n659));
  NAND4_X1  g473(.A1(new_n641), .A2(new_n628), .A3(new_n601), .A4(new_n659), .ZN(new_n660));
  NOR2_X1   g474(.A1(new_n656), .A2(new_n660), .ZN(new_n661));
  XNOR2_X1  g475(.A(new_n661), .B(new_n228), .ZN(G30));
  XOR2_X1   g476(.A(new_n659), .B(KEYINPUT39), .Z(new_n663));
  INV_X1    g477(.A(new_n663), .ZN(new_n664));
  NAND2_X1  g478(.A1(new_n429), .A2(new_n664), .ZN(new_n665));
  XOR2_X1   g479(.A(new_n665), .B(KEYINPUT40), .Z(new_n666));
  NAND2_X1  g480(.A1(new_n290), .A2(new_n291), .ZN(new_n667));
  OAI21_X1  g481(.A(new_n278), .B1(new_n262), .B2(new_n192), .ZN(new_n668));
  AOI21_X1  g482(.A(new_n632), .B1(new_n668), .B2(new_n274), .ZN(new_n669));
  NOR2_X1   g483(.A1(new_n667), .A2(new_n669), .ZN(new_n670));
  INV_X1    g484(.A(new_n670), .ZN(new_n671));
  NOR2_X1   g485(.A1(new_n476), .A2(new_n477), .ZN(new_n672));
  XNOR2_X1  g486(.A(KEYINPUT97), .B(KEYINPUT38), .ZN(new_n673));
  XOR2_X1   g487(.A(new_n672), .B(new_n673), .Z(new_n674));
  AOI22_X1  g488(.A1(new_n351), .A2(new_n353), .B1(new_n355), .B2(new_n648), .ZN(new_n675));
  AOI21_X1  g489(.A(new_n600), .B1(new_n541), .B2(new_n544), .ZN(new_n676));
  AND4_X1   g490(.A1(new_n430), .A2(new_n674), .A3(new_n675), .A4(new_n676), .ZN(new_n677));
  NAND3_X1  g491(.A1(new_n666), .A2(new_n671), .A3(new_n677), .ZN(new_n678));
  XNOR2_X1  g492(.A(new_n678), .B(G143), .ZN(G45));
  NAND4_X1  g493(.A1(new_n545), .A2(new_n628), .A3(new_n621), .A4(new_n659), .ZN(new_n680));
  INV_X1    g494(.A(KEYINPUT98), .ZN(new_n681));
  NAND2_X1  g495(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  AOI21_X1  g496(.A(new_n620), .B1(new_n541), .B2(new_n544), .ZN(new_n683));
  NAND4_X1  g497(.A1(new_n683), .A2(KEYINPUT98), .A3(new_n628), .A4(new_n659), .ZN(new_n684));
  NAND2_X1  g498(.A1(new_n682), .A2(new_n684), .ZN(new_n685));
  NOR2_X1   g499(.A1(new_n685), .A2(new_n656), .ZN(new_n686));
  XNOR2_X1  g500(.A(new_n686), .B(new_n221), .ZN(G48));
  AOI21_X1  g501(.A(G902), .B1(new_n412), .B2(new_n416), .ZN(new_n688));
  AOI21_X1  g502(.A(KEYINPUT99), .B1(new_n688), .B2(new_n418), .ZN(new_n689));
  INV_X1    g503(.A(new_n395), .ZN(new_n690));
  AOI21_X1  g504(.A(new_n394), .B1(new_n208), .B2(new_n219), .ZN(new_n691));
  NOR2_X1   g505(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  OAI211_X1 g506(.A(new_n400), .B(new_n398), .C1(new_n468), .C2(new_n216), .ZN(new_n693));
  OAI21_X1  g507(.A(new_n390), .B1(new_n692), .B2(new_n693), .ZN(new_n694));
  AOI21_X1  g508(.A(KEYINPUT81), .B1(new_n381), .B2(new_n383), .ZN(new_n695));
  NOR2_X1   g509(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  AOI22_X1  g510(.A1(new_n696), .A2(new_n411), .B1(new_n415), .B2(new_n391), .ZN(new_n697));
  OAI21_X1  g511(.A(G469), .B1(new_n697), .B2(G902), .ZN(new_n698));
  NAND2_X1  g512(.A1(new_n689), .A2(new_n698), .ZN(new_n699));
  OAI211_X1 g513(.A(KEYINPUT99), .B(G469), .C1(new_n697), .C2(G902), .ZN(new_n700));
  AOI21_X1  g514(.A(new_n427), .B1(new_n699), .B2(new_n700), .ZN(new_n701));
  NAND4_X1  g515(.A1(new_n631), .A2(new_n701), .A3(new_n292), .A4(new_n360), .ZN(new_n702));
  XNOR2_X1  g516(.A(KEYINPUT41), .B(G113), .ZN(new_n703));
  XNOR2_X1  g517(.A(new_n702), .B(new_n703), .ZN(G15));
  INV_X1    g518(.A(new_n361), .ZN(new_n705));
  AOI211_X1 g519(.A(new_n478), .B(new_n427), .C1(new_n699), .C2(new_n700), .ZN(new_n706));
  AND4_X1   g520(.A1(new_n544), .A2(new_n601), .A3(new_n640), .A4(new_n629), .ZN(new_n707));
  NAND3_X1  g521(.A1(new_n705), .A2(new_n706), .A3(new_n707), .ZN(new_n708));
  XOR2_X1   g522(.A(KEYINPUT100), .B(G116), .Z(new_n709));
  XNOR2_X1  g523(.A(new_n708), .B(new_n709), .ZN(G18));
  NAND3_X1  g524(.A1(new_n292), .A2(new_n611), .A3(new_n650), .ZN(new_n711));
  NAND2_X1  g525(.A1(new_n699), .A2(new_n700), .ZN(new_n712));
  NAND3_X1  g526(.A1(new_n712), .A2(new_n628), .A3(new_n428), .ZN(new_n713));
  OR2_X1    g527(.A1(new_n711), .A2(new_n713), .ZN(new_n714));
  XNOR2_X1  g528(.A(new_n714), .B(G119), .ZN(G21));
  XOR2_X1   g529(.A(new_n287), .B(KEYINPUT101), .Z(new_n716));
  INV_X1    g530(.A(new_n716), .ZN(new_n717));
  AND2_X1   g531(.A1(new_n279), .A2(new_n284), .ZN(new_n718));
  AOI21_X1  g532(.A(new_n259), .B1(new_n280), .B2(new_n256), .ZN(new_n719));
  OAI21_X1  g533(.A(new_n260), .B1(new_n719), .B2(new_n271), .ZN(new_n720));
  INV_X1    g534(.A(new_n272), .ZN(new_n721));
  OAI21_X1  g535(.A(new_n193), .B1(new_n720), .B2(new_n721), .ZN(new_n722));
  AOI21_X1  g536(.A(new_n717), .B1(new_n718), .B2(new_n722), .ZN(new_n723));
  NOR2_X1   g537(.A1(new_n723), .A2(new_n633), .ZN(new_n724));
  NAND4_X1  g538(.A1(new_n701), .A2(new_n360), .A3(new_n629), .A4(new_n724), .ZN(new_n725));
  AND3_X1   g539(.A1(new_n676), .A2(KEYINPUT102), .A3(new_n628), .ZN(new_n726));
  AOI21_X1  g540(.A(KEYINPUT102), .B1(new_n676), .B2(new_n628), .ZN(new_n727));
  NOR2_X1   g541(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  OR2_X1    g542(.A1(new_n725), .A2(new_n728), .ZN(new_n729));
  XOR2_X1   g543(.A(KEYINPUT103), .B(G122), .Z(new_n730));
  XNOR2_X1  g544(.A(new_n729), .B(new_n730), .ZN(G24));
  NAND2_X1  g545(.A1(new_n718), .A2(new_n722), .ZN(new_n732));
  NAND2_X1  g546(.A1(new_n732), .A2(new_n716), .ZN(new_n733));
  NAND3_X1  g547(.A1(new_n650), .A2(new_n733), .A3(new_n651), .ZN(new_n734));
  NAND2_X1  g548(.A1(new_n683), .A2(new_n659), .ZN(new_n735));
  NAND2_X1  g549(.A1(new_n735), .A2(KEYINPUT104), .ZN(new_n736));
  INV_X1    g550(.A(KEYINPUT104), .ZN(new_n737));
  NAND3_X1  g551(.A1(new_n683), .A2(new_n737), .A3(new_n659), .ZN(new_n738));
  AOI21_X1  g552(.A(new_n734), .B1(new_n736), .B2(new_n738), .ZN(new_n739));
  AOI21_X1  g553(.A(KEYINPUT105), .B1(new_n739), .B2(new_n706), .ZN(new_n740));
  NOR3_X1   g554(.A1(new_n675), .A2(new_n723), .A3(new_n633), .ZN(new_n741));
  AND4_X1   g555(.A1(new_n737), .A2(new_n545), .A3(new_n621), .A4(new_n659), .ZN(new_n742));
  AOI21_X1  g556(.A(new_n737), .B1(new_n683), .B2(new_n659), .ZN(new_n743));
  OAI21_X1  g557(.A(new_n741), .B1(new_n742), .B2(new_n743), .ZN(new_n744));
  INV_X1    g558(.A(KEYINPUT105), .ZN(new_n745));
  NOR3_X1   g559(.A1(new_n744), .A2(new_n745), .A3(new_n713), .ZN(new_n746));
  NOR2_X1   g560(.A1(new_n740), .A2(new_n746), .ZN(new_n747));
  XNOR2_X1  g561(.A(new_n747), .B(new_n301), .ZN(G27));
  INV_X1    g562(.A(new_n291), .ZN(new_n749));
  AOI21_X1  g563(.A(KEYINPUT32), .B1(new_n285), .B2(new_n287), .ZN(new_n750));
  OAI21_X1  g564(.A(KEYINPUT107), .B1(new_n749), .B2(new_n750), .ZN(new_n751));
  INV_X1    g565(.A(KEYINPUT108), .ZN(new_n752));
  OAI211_X1 g566(.A(new_n751), .B(new_n752), .C1(KEYINPUT107), .C2(new_n750), .ZN(new_n753));
  INV_X1    g567(.A(KEYINPUT107), .ZN(new_n754));
  AOI21_X1  g568(.A(new_n754), .B1(new_n290), .B2(new_n291), .ZN(new_n755));
  NOR2_X1   g569(.A1(new_n750), .A2(KEYINPUT107), .ZN(new_n756));
  OAI21_X1  g570(.A(KEYINPUT108), .B1(new_n755), .B2(new_n756), .ZN(new_n757));
  NAND3_X1  g571(.A1(new_n753), .A2(new_n757), .A3(new_n276), .ZN(new_n758));
  INV_X1    g572(.A(KEYINPUT106), .ZN(new_n759));
  NAND2_X1  g573(.A1(new_n422), .A2(new_n759), .ZN(new_n760));
  NAND3_X1  g574(.A1(new_n421), .A2(KEYINPUT106), .A3(new_n391), .ZN(new_n761));
  NAND4_X1  g575(.A1(new_n760), .A2(G469), .A3(new_n423), .A4(new_n761), .ZN(new_n762));
  NAND3_X1  g576(.A1(new_n762), .A2(new_n419), .A3(new_n420), .ZN(new_n763));
  NOR3_X1   g577(.A1(new_n476), .A2(new_n477), .A3(new_n623), .ZN(new_n764));
  NAND4_X1  g578(.A1(new_n763), .A2(KEYINPUT42), .A3(new_n428), .A4(new_n764), .ZN(new_n765));
  AOI21_X1  g579(.A(new_n765), .B1(new_n736), .B2(new_n738), .ZN(new_n766));
  NAND3_X1  g580(.A1(new_n758), .A2(new_n360), .A3(new_n766), .ZN(new_n767));
  NAND2_X1  g581(.A1(new_n736), .A2(new_n738), .ZN(new_n768));
  NAND2_X1  g582(.A1(new_n763), .A2(new_n428), .ZN(new_n769));
  INV_X1    g583(.A(new_n764), .ZN(new_n770));
  NOR2_X1   g584(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  NAND3_X1  g585(.A1(new_n705), .A2(new_n768), .A3(new_n771), .ZN(new_n772));
  INV_X1    g586(.A(KEYINPUT42), .ZN(new_n773));
  NAND2_X1  g587(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  NAND2_X1  g588(.A1(new_n767), .A2(new_n774), .ZN(new_n775));
  XNOR2_X1  g589(.A(new_n775), .B(G131), .ZN(G33));
  INV_X1    g590(.A(new_n659), .ZN(new_n777));
  NOR2_X1   g591(.A1(new_n642), .A2(new_n777), .ZN(new_n778));
  NAND3_X1  g592(.A1(new_n705), .A2(new_n778), .A3(new_n771), .ZN(new_n779));
  XNOR2_X1  g593(.A(new_n779), .B(G134), .ZN(G36));
  NAND4_X1  g594(.A1(new_n760), .A2(KEYINPUT45), .A3(new_n423), .A4(new_n761), .ZN(new_n781));
  AND2_X1   g595(.A1(new_n422), .A2(new_n423), .ZN(new_n782));
  OAI211_X1 g596(.A(new_n781), .B(G469), .C1(KEYINPUT45), .C2(new_n782), .ZN(new_n783));
  NAND3_X1  g597(.A1(new_n783), .A2(KEYINPUT46), .A3(new_n420), .ZN(new_n784));
  AND2_X1   g598(.A1(new_n784), .A2(new_n419), .ZN(new_n785));
  NAND2_X1  g599(.A1(new_n783), .A2(new_n420), .ZN(new_n786));
  INV_X1    g600(.A(KEYINPUT46), .ZN(new_n787));
  NAND2_X1  g601(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  NAND2_X1  g602(.A1(new_n785), .A2(new_n788), .ZN(new_n789));
  NAND2_X1  g603(.A1(new_n789), .A2(new_n428), .ZN(new_n790));
  NOR2_X1   g604(.A1(new_n790), .A2(new_n663), .ZN(new_n791));
  NOR2_X1   g605(.A1(new_n545), .A2(new_n620), .ZN(new_n792));
  XNOR2_X1  g606(.A(new_n792), .B(KEYINPUT43), .ZN(new_n793));
  INV_X1    g607(.A(new_n634), .ZN(new_n794));
  NAND3_X1  g608(.A1(new_n793), .A2(new_n794), .A3(new_n650), .ZN(new_n795));
  INV_X1    g609(.A(KEYINPUT44), .ZN(new_n796));
  AOI21_X1  g610(.A(new_n770), .B1(new_n795), .B2(new_n796), .ZN(new_n797));
  OAI211_X1 g611(.A(new_n791), .B(new_n797), .C1(new_n796), .C2(new_n795), .ZN(new_n798));
  XNOR2_X1  g612(.A(new_n798), .B(G137), .ZN(G39));
  INV_X1    g613(.A(KEYINPUT47), .ZN(new_n800));
  NOR2_X1   g614(.A1(new_n800), .A2(KEYINPUT109), .ZN(new_n801));
  NAND2_X1  g615(.A1(new_n790), .A2(new_n801), .ZN(new_n802));
  INV_X1    g616(.A(new_n801), .ZN(new_n803));
  AOI21_X1  g617(.A(new_n427), .B1(new_n785), .B2(new_n788), .ZN(new_n804));
  NAND2_X1  g618(.A1(new_n800), .A2(KEYINPUT109), .ZN(new_n805));
  INV_X1    g619(.A(new_n805), .ZN(new_n806));
  OAI21_X1  g620(.A(new_n803), .B1(new_n804), .B2(new_n806), .ZN(new_n807));
  NOR4_X1   g621(.A1(new_n292), .A2(new_n735), .A3(new_n360), .A4(new_n770), .ZN(new_n808));
  NAND3_X1  g622(.A1(new_n802), .A2(new_n807), .A3(new_n808), .ZN(new_n809));
  XNOR2_X1  g623(.A(new_n809), .B(G140), .ZN(G42));
  NOR2_X1   g624(.A1(G952), .A2(G953), .ZN(new_n811));
  INV_X1    g625(.A(KEYINPUT53), .ZN(new_n812));
  INV_X1    g626(.A(new_n656), .ZN(new_n813));
  AND2_X1   g627(.A1(new_n682), .A2(new_n684), .ZN(new_n814));
  INV_X1    g628(.A(new_n660), .ZN(new_n815));
  OAI21_X1  g629(.A(new_n813), .B1(new_n814), .B2(new_n815), .ZN(new_n816));
  INV_X1    g630(.A(new_n728), .ZN(new_n817));
  XOR2_X1   g631(.A(new_n659), .B(KEYINPUT112), .Z(new_n818));
  NOR3_X1   g632(.A1(new_n769), .A2(new_n650), .A3(new_n818), .ZN(new_n819));
  NAND3_X1  g633(.A1(new_n817), .A2(new_n671), .A3(new_n819), .ZN(new_n820));
  OAI211_X1 g634(.A(new_n816), .B(new_n820), .C1(new_n740), .C2(new_n746), .ZN(new_n821));
  NAND2_X1  g635(.A1(new_n821), .A2(KEYINPUT113), .ZN(new_n822));
  INV_X1    g636(.A(KEYINPUT52), .ZN(new_n823));
  AOI21_X1  g637(.A(new_n656), .B1(new_n685), .B2(new_n660), .ZN(new_n824));
  OAI21_X1  g638(.A(new_n745), .B1(new_n744), .B2(new_n713), .ZN(new_n825));
  NAND4_X1  g639(.A1(new_n768), .A2(new_n706), .A3(KEYINPUT105), .A4(new_n741), .ZN(new_n826));
  AOI21_X1  g640(.A(new_n824), .B1(new_n825), .B2(new_n826), .ZN(new_n827));
  INV_X1    g641(.A(KEYINPUT113), .ZN(new_n828));
  NAND3_X1  g642(.A1(new_n827), .A2(new_n828), .A3(new_n820), .ZN(new_n829));
  NAND3_X1  g643(.A1(new_n822), .A2(new_n823), .A3(new_n829), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n775), .A2(new_n779), .ZN(new_n831));
  OAI21_X1  g645(.A(new_n622), .B1(new_n545), .B2(new_n600), .ZN(new_n832));
  AOI21_X1  g646(.A(new_n610), .B1(new_n480), .B2(new_n481), .ZN(new_n833));
  NAND4_X1  g647(.A1(new_n615), .A2(new_n832), .A3(new_n833), .A4(new_n634), .ZN(new_n834));
  OAI21_X1  g648(.A(new_n834), .B1(new_n725), .B2(new_n728), .ZN(new_n835));
  NAND3_X1  g649(.A1(new_n701), .A2(new_n628), .A3(new_n707), .ZN(new_n836));
  OAI22_X1  g650(.A1(new_n836), .A2(new_n361), .B1(new_n711), .B2(new_n713), .ZN(new_n837));
  NOR2_X1   g651(.A1(new_n835), .A2(new_n837), .ZN(new_n838));
  AND2_X1   g652(.A1(new_n653), .A2(new_n702), .ZN(new_n839));
  AND2_X1   g653(.A1(new_n292), .A2(new_n429), .ZN(new_n840));
  NOR2_X1   g654(.A1(new_n601), .A2(new_n777), .ZN(new_n841));
  AND4_X1   g655(.A1(new_n641), .A2(new_n650), .A3(new_n764), .A4(new_n841), .ZN(new_n842));
  AOI22_X1  g656(.A1(new_n739), .A2(new_n771), .B1(new_n840), .B2(new_n842), .ZN(new_n843));
  NAND4_X1  g657(.A1(new_n838), .A2(new_n613), .A3(new_n839), .A4(new_n843), .ZN(new_n844));
  NOR2_X1   g658(.A1(new_n831), .A2(new_n844), .ZN(new_n845));
  NAND2_X1  g659(.A1(new_n830), .A2(new_n845), .ZN(new_n846));
  AOI21_X1  g660(.A(new_n823), .B1(new_n822), .B2(new_n829), .ZN(new_n847));
  OAI21_X1  g661(.A(new_n812), .B1(new_n846), .B2(new_n847), .ZN(new_n848));
  INV_X1    g662(.A(KEYINPUT54), .ZN(new_n849));
  NAND2_X1  g663(.A1(new_n821), .A2(KEYINPUT52), .ZN(new_n850));
  NAND4_X1  g664(.A1(new_n830), .A2(new_n845), .A3(KEYINPUT53), .A4(new_n850), .ZN(new_n851));
  AND3_X1   g665(.A1(new_n848), .A2(new_n849), .A3(new_n851), .ZN(new_n852));
  AND2_X1   g666(.A1(new_n830), .A2(new_n845), .ZN(new_n853));
  NOR2_X1   g667(.A1(new_n821), .A2(KEYINPUT113), .ZN(new_n854));
  AOI21_X1  g668(.A(new_n828), .B1(new_n827), .B2(new_n820), .ZN(new_n855));
  OAI21_X1  g669(.A(KEYINPUT52), .B1(new_n854), .B2(new_n855), .ZN(new_n856));
  NAND4_X1  g670(.A1(new_n853), .A2(KEYINPUT114), .A3(KEYINPUT53), .A4(new_n856), .ZN(new_n857));
  NAND4_X1  g671(.A1(new_n856), .A2(KEYINPUT53), .A3(new_n830), .A4(new_n845), .ZN(new_n858));
  INV_X1    g672(.A(KEYINPUT114), .ZN(new_n859));
  NAND2_X1  g673(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  AND3_X1   g674(.A1(new_n838), .A2(new_n613), .A3(new_n839), .ZN(new_n861));
  INV_X1    g675(.A(KEYINPUT111), .ZN(new_n862));
  INV_X1    g676(.A(new_n779), .ZN(new_n863));
  AOI21_X1  g677(.A(new_n863), .B1(new_n767), .B2(new_n774), .ZN(new_n864));
  NAND4_X1  g678(.A1(new_n861), .A2(new_n862), .A3(new_n864), .A4(new_n843), .ZN(new_n865));
  OAI21_X1  g679(.A(KEYINPUT111), .B1(new_n831), .B2(new_n844), .ZN(new_n866));
  NAND4_X1  g680(.A1(new_n865), .A2(new_n866), .A3(new_n830), .A4(new_n850), .ZN(new_n867));
  NAND2_X1  g681(.A1(new_n867), .A2(new_n812), .ZN(new_n868));
  NAND3_X1  g682(.A1(new_n857), .A2(new_n860), .A3(new_n868), .ZN(new_n869));
  AOI21_X1  g683(.A(new_n852), .B1(KEYINPUT54), .B2(new_n869), .ZN(new_n870));
  NAND2_X1  g684(.A1(new_n802), .A2(new_n807), .ZN(new_n871));
  NAND2_X1  g685(.A1(new_n712), .A2(new_n427), .ZN(new_n872));
  NAND2_X1  g686(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  NAND2_X1  g687(.A1(new_n793), .A2(new_n606), .ZN(new_n874));
  INV_X1    g688(.A(new_n874), .ZN(new_n875));
  INV_X1    g689(.A(new_n360), .ZN(new_n876));
  NOR3_X1   g690(.A1(new_n876), .A2(new_n633), .A3(new_n723), .ZN(new_n877));
  NAND3_X1  g691(.A1(new_n875), .A2(new_n877), .A3(new_n764), .ZN(new_n878));
  OR2_X1    g692(.A1(new_n878), .A2(KEYINPUT115), .ZN(new_n879));
  NAND2_X1  g693(.A1(new_n878), .A2(KEYINPUT115), .ZN(new_n880));
  NAND3_X1  g694(.A1(new_n873), .A2(new_n879), .A3(new_n880), .ZN(new_n881));
  NAND2_X1  g695(.A1(new_n701), .A2(new_n764), .ZN(new_n882));
  NOR2_X1   g696(.A1(new_n874), .A2(new_n882), .ZN(new_n883));
  NAND2_X1  g697(.A1(new_n883), .A2(new_n741), .ZN(new_n884));
  NOR2_X1   g698(.A1(new_n876), .A2(new_n605), .ZN(new_n885));
  NAND4_X1  g699(.A1(new_n670), .A2(new_n885), .A3(new_n701), .A4(new_n764), .ZN(new_n886));
  OR3_X1    g700(.A1(new_n886), .A2(new_n545), .A3(new_n621), .ZN(new_n887));
  NAND2_X1  g701(.A1(new_n884), .A2(new_n887), .ZN(new_n888));
  NAND2_X1  g702(.A1(new_n712), .A2(new_n428), .ZN(new_n889));
  NOR3_X1   g703(.A1(new_n889), .A2(new_n674), .A3(new_n430), .ZN(new_n890));
  NAND4_X1  g704(.A1(new_n875), .A2(KEYINPUT50), .A3(new_n877), .A4(new_n890), .ZN(new_n891));
  INV_X1    g705(.A(KEYINPUT50), .ZN(new_n892));
  NAND2_X1  g706(.A1(new_n875), .A2(new_n877), .ZN(new_n893));
  INV_X1    g707(.A(new_n890), .ZN(new_n894));
  OAI21_X1  g708(.A(new_n892), .B1(new_n893), .B2(new_n894), .ZN(new_n895));
  AOI21_X1  g709(.A(new_n888), .B1(new_n891), .B2(new_n895), .ZN(new_n896));
  NAND3_X1  g710(.A1(new_n881), .A2(new_n896), .A3(KEYINPUT51), .ZN(new_n897));
  INV_X1    g711(.A(KEYINPUT117), .ZN(new_n898));
  NAND2_X1  g712(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  NAND4_X1  g713(.A1(new_n881), .A2(new_n896), .A3(KEYINPUT117), .A4(KEYINPUT51), .ZN(new_n900));
  NAND2_X1  g714(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  XOR2_X1   g715(.A(new_n872), .B(KEYINPUT116), .Z(new_n902));
  NAND2_X1  g716(.A1(new_n871), .A2(new_n902), .ZN(new_n903));
  NAND3_X1  g717(.A1(new_n903), .A2(new_n879), .A3(new_n880), .ZN(new_n904));
  AOI21_X1  g718(.A(KEYINPUT51), .B1(new_n904), .B2(new_n896), .ZN(new_n905));
  AND2_X1   g719(.A1(new_n758), .A2(new_n360), .ZN(new_n906));
  NAND2_X1  g720(.A1(new_n906), .A2(new_n883), .ZN(new_n907));
  XOR2_X1   g721(.A(new_n907), .B(KEYINPUT48), .Z(new_n908));
  OAI221_X1 g722(.A(new_n603), .B1(new_n622), .B2(new_n886), .C1(new_n893), .C2(new_n713), .ZN(new_n909));
  NOR3_X1   g723(.A1(new_n905), .A2(new_n908), .A3(new_n909), .ZN(new_n910));
  AND2_X1   g724(.A1(new_n901), .A2(new_n910), .ZN(new_n911));
  AOI21_X1  g725(.A(new_n811), .B1(new_n870), .B2(new_n911), .ZN(new_n912));
  INV_X1    g726(.A(KEYINPUT49), .ZN(new_n913));
  AOI211_X1 g727(.A(new_n674), .B(new_n671), .C1(new_n913), .C2(new_n712), .ZN(new_n914));
  NOR3_X1   g728(.A1(new_n876), .A2(new_n623), .A3(new_n427), .ZN(new_n915));
  OAI211_X1 g729(.A(new_n915), .B(new_n792), .C1(new_n913), .C2(new_n712), .ZN(new_n916));
  OR2_X1    g730(.A1(new_n916), .A2(KEYINPUT110), .ZN(new_n917));
  NAND2_X1  g731(.A1(new_n916), .A2(KEYINPUT110), .ZN(new_n918));
  NAND3_X1  g732(.A1(new_n914), .A2(new_n917), .A3(new_n918), .ZN(new_n919));
  INV_X1    g733(.A(new_n919), .ZN(new_n920));
  OAI21_X1  g734(.A(KEYINPUT118), .B1(new_n912), .B2(new_n920), .ZN(new_n921));
  INV_X1    g735(.A(KEYINPUT118), .ZN(new_n922));
  NAND2_X1  g736(.A1(new_n869), .A2(KEYINPUT54), .ZN(new_n923));
  INV_X1    g737(.A(new_n852), .ZN(new_n924));
  AND3_X1   g738(.A1(new_n923), .A2(new_n924), .A3(new_n911), .ZN(new_n925));
  OAI211_X1 g739(.A(new_n922), .B(new_n919), .C1(new_n925), .C2(new_n811), .ZN(new_n926));
  NAND2_X1  g740(.A1(new_n921), .A2(new_n926), .ZN(G75));
  NAND2_X1  g741(.A1(new_n471), .A2(new_n473), .ZN(new_n928));
  XOR2_X1   g742(.A(new_n928), .B(new_n466), .Z(new_n929));
  XNOR2_X1  g743(.A(new_n929), .B(KEYINPUT55), .ZN(new_n930));
  INV_X1    g744(.A(KEYINPUT56), .ZN(new_n931));
  NAND2_X1  g745(.A1(new_n848), .A2(new_n851), .ZN(new_n932));
  NAND2_X1  g746(.A1(new_n932), .A2(G902), .ZN(new_n933));
  INV_X1    g747(.A(G210), .ZN(new_n934));
  OAI21_X1  g748(.A(new_n931), .B1(new_n933), .B2(new_n934), .ZN(new_n935));
  NAND2_X1  g749(.A1(new_n935), .A2(KEYINPUT119), .ZN(new_n936));
  INV_X1    g750(.A(KEYINPUT119), .ZN(new_n937));
  OAI211_X1 g751(.A(new_n937), .B(new_n931), .C1(new_n933), .C2(new_n934), .ZN(new_n938));
  AOI21_X1  g752(.A(new_n930), .B1(new_n936), .B2(new_n938), .ZN(new_n939));
  NAND2_X1  g753(.A1(new_n938), .A2(new_n930), .ZN(new_n940));
  NAND2_X1  g754(.A1(new_n602), .A2(G953), .ZN(new_n941));
  XOR2_X1   g755(.A(new_n941), .B(KEYINPUT120), .Z(new_n942));
  NAND2_X1  g756(.A1(new_n940), .A2(new_n942), .ZN(new_n943));
  NOR2_X1   g757(.A1(new_n939), .A2(new_n943), .ZN(G51));
  INV_X1    g758(.A(new_n942), .ZN(new_n945));
  NOR2_X1   g759(.A1(new_n933), .A2(new_n783), .ZN(new_n946));
  AOI21_X1  g760(.A(new_n849), .B1(new_n848), .B2(new_n851), .ZN(new_n947));
  NOR2_X1   g761(.A1(new_n852), .A2(new_n947), .ZN(new_n948));
  XNOR2_X1  g762(.A(new_n420), .B(KEYINPUT121), .ZN(new_n949));
  XNOR2_X1  g763(.A(new_n949), .B(KEYINPUT57), .ZN(new_n950));
  INV_X1    g764(.A(new_n950), .ZN(new_n951));
  OAI21_X1  g765(.A(new_n417), .B1(new_n948), .B2(new_n951), .ZN(new_n952));
  INV_X1    g766(.A(KEYINPUT122), .ZN(new_n953));
  AOI21_X1  g767(.A(new_n946), .B1(new_n952), .B2(new_n953), .ZN(new_n954));
  OAI211_X1 g768(.A(KEYINPUT122), .B(new_n417), .C1(new_n948), .C2(new_n951), .ZN(new_n955));
  AOI21_X1  g769(.A(new_n945), .B1(new_n954), .B2(new_n955), .ZN(G54));
  AND4_X1   g770(.A1(KEYINPUT58), .A2(new_n932), .A3(G475), .A4(G902), .ZN(new_n957));
  INV_X1    g771(.A(new_n538), .ZN(new_n958));
  OR2_X1    g772(.A1(new_n957), .A2(new_n958), .ZN(new_n959));
  NAND2_X1  g773(.A1(new_n957), .A2(new_n958), .ZN(new_n960));
  AOI21_X1  g774(.A(new_n945), .B1(new_n959), .B2(new_n960), .ZN(G60));
  INV_X1    g775(.A(new_n618), .ZN(new_n962));
  NAND2_X1  g776(.A1(G478), .A2(G902), .ZN(new_n963));
  XOR2_X1   g777(.A(new_n963), .B(KEYINPUT59), .Z(new_n964));
  OR2_X1    g778(.A1(new_n962), .A2(new_n964), .ZN(new_n965));
  OAI21_X1  g779(.A(new_n942), .B1(new_n948), .B2(new_n965), .ZN(new_n966));
  OR2_X1    g780(.A1(new_n870), .A2(new_n964), .ZN(new_n967));
  AOI21_X1  g781(.A(new_n966), .B1(new_n967), .B2(new_n962), .ZN(G63));
  AND2_X1   g782(.A1(new_n848), .A2(new_n851), .ZN(new_n969));
  NAND2_X1  g783(.A1(G217), .A2(G902), .ZN(new_n970));
  XNOR2_X1  g784(.A(new_n970), .B(KEYINPUT60), .ZN(new_n971));
  NOR2_X1   g785(.A1(new_n969), .A2(new_n971), .ZN(new_n972));
  AOI21_X1  g786(.A(new_n945), .B1(new_n972), .B2(new_n648), .ZN(new_n973));
  XNOR2_X1  g787(.A(new_n359), .B(KEYINPUT123), .ZN(new_n974));
  OAI21_X1  g788(.A(new_n974), .B1(new_n969), .B2(new_n971), .ZN(new_n975));
  NAND2_X1  g789(.A1(new_n973), .A2(new_n975), .ZN(new_n976));
  NAND2_X1  g790(.A1(new_n972), .A2(new_n648), .ZN(new_n977));
  INV_X1    g791(.A(KEYINPUT124), .ZN(new_n978));
  AOI21_X1  g792(.A(KEYINPUT61), .B1(new_n977), .B2(new_n978), .ZN(new_n979));
  NAND2_X1  g793(.A1(new_n976), .A2(new_n979), .ZN(new_n980));
  AOI21_X1  g794(.A(KEYINPUT124), .B1(new_n972), .B2(new_n648), .ZN(new_n981));
  OAI211_X1 g795(.A(new_n975), .B(new_n973), .C1(new_n981), .C2(KEYINPUT61), .ZN(new_n982));
  NAND2_X1  g796(.A1(new_n980), .A2(new_n982), .ZN(G66));
  NOR2_X1   g797(.A1(new_n861), .A2(G953), .ZN(new_n984));
  XNOR2_X1  g798(.A(new_n984), .B(KEYINPUT125), .ZN(new_n985));
  OAI21_X1  g799(.A(G953), .B1(new_n609), .B2(new_n444), .ZN(new_n986));
  NAND2_X1  g800(.A1(new_n985), .A2(new_n986), .ZN(new_n987));
  OAI21_X1  g801(.A(new_n928), .B1(G898), .B2(new_n564), .ZN(new_n988));
  XNOR2_X1  g802(.A(new_n987), .B(new_n988), .ZN(G69));
  NAND2_X1  g803(.A1(new_n238), .A2(new_n254), .ZN(new_n990));
  XNOR2_X1  g804(.A(new_n990), .B(new_n498), .ZN(new_n991));
  NAND2_X1  g805(.A1(new_n798), .A2(new_n809), .ZN(new_n992));
  NOR3_X1   g806(.A1(new_n992), .A2(new_n747), .A3(new_n824), .ZN(new_n993));
  NAND3_X1  g807(.A1(new_n791), .A2(new_n817), .A3(new_n906), .ZN(new_n994));
  NAND3_X1  g808(.A1(new_n993), .A2(new_n864), .A3(new_n994), .ZN(new_n995));
  NAND2_X1  g809(.A1(new_n995), .A2(new_n564), .ZN(new_n996));
  NAND3_X1  g810(.A1(new_n388), .A2(G900), .A3(G953), .ZN(new_n997));
  AOI21_X1  g811(.A(new_n991), .B1(new_n996), .B2(new_n997), .ZN(new_n998));
  NOR2_X1   g812(.A1(new_n665), .A2(new_n770), .ZN(new_n999));
  NAND3_X1  g813(.A1(new_n365), .A2(new_n832), .A3(new_n999), .ZN(new_n1000));
  INV_X1    g814(.A(KEYINPUT126), .ZN(new_n1001));
  AND2_X1   g815(.A1(new_n1000), .A2(new_n1001), .ZN(new_n1002));
  NAND2_X1  g816(.A1(new_n678), .A2(new_n827), .ZN(new_n1003));
  INV_X1    g817(.A(new_n1003), .ZN(new_n1004));
  OR2_X1    g818(.A1(new_n1004), .A2(KEYINPUT62), .ZN(new_n1005));
  NAND2_X1  g819(.A1(new_n1004), .A2(KEYINPUT62), .ZN(new_n1006));
  AOI211_X1 g820(.A(new_n1002), .B(new_n992), .C1(new_n1005), .C2(new_n1006), .ZN(new_n1007));
  OAI211_X1 g821(.A(new_n1007), .B(new_n564), .C1(new_n1001), .C2(new_n1000), .ZN(new_n1008));
  NAND3_X1  g822(.A1(G227), .A2(G900), .A3(G953), .ZN(new_n1009));
  NAND2_X1  g823(.A1(new_n1008), .A2(new_n1009), .ZN(new_n1010));
  AOI21_X1  g824(.A(new_n998), .B1(new_n1010), .B2(new_n991), .ZN(G72));
  NAND2_X1  g825(.A1(G472), .A2(G902), .ZN(new_n1012));
  XOR2_X1   g826(.A(new_n1012), .B(KEYINPUT63), .Z(new_n1013));
  INV_X1    g827(.A(new_n861), .ZN(new_n1014));
  OAI21_X1  g828(.A(new_n1013), .B1(new_n995), .B2(new_n1014), .ZN(new_n1015));
  NAND4_X1  g829(.A1(new_n1015), .A2(new_n193), .A3(new_n256), .A4(new_n277), .ZN(new_n1016));
  INV_X1    g830(.A(new_n1013), .ZN(new_n1017));
  NOR2_X1   g831(.A1(new_n1000), .A2(new_n1001), .ZN(new_n1018));
  NOR2_X1   g832(.A1(new_n1014), .A2(new_n1018), .ZN(new_n1019));
  AOI21_X1  g833(.A(new_n1017), .B1(new_n1007), .B2(new_n1019), .ZN(new_n1020));
  OAI21_X1  g834(.A(new_n192), .B1(new_n255), .B2(new_n257), .ZN(new_n1021));
  OAI211_X1 g835(.A(new_n1016), .B(new_n942), .C1(new_n1020), .C2(new_n1021), .ZN(new_n1022));
  AOI21_X1  g836(.A(new_n1017), .B1(new_n258), .B2(new_n278), .ZN(new_n1023));
  XOR2_X1   g837(.A(new_n1023), .B(KEYINPUT127), .Z(new_n1024));
  AOI21_X1  g838(.A(new_n1022), .B1(new_n869), .B2(new_n1024), .ZN(G57));
endmodule


