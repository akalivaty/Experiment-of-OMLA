

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
         n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597,
         n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608,
         n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619,
         n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630,
         n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641,
         n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652,
         n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663,
         n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674,
         n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685,
         n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696,
         n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707,
         n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718,
         n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729,
         n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740,
         n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751,
         n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762,
         n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773,
         n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784,
         n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, n795,
         n796, n797, n798, n799, n800, n801, n802, n803, n804, n805, n806,
         n807, n808, n809, n810, n811, n812, n813, n814, n815, n816, n817,
         n818, n819, n820, n821, n822, n823, n824, n825, n826, n827, n828,
         n829, n830, n831, n832, n833, n834, n835, n836, n837, n838, n839,
         n840, n841, n842, n843, n844, n845, n846, n847, n848, n849, n850,
         n851, n852, n853, n854, n855, n856, n857, n858, n859, n860, n861,
         n862, n863, n864, n865, n866, n867, n868, n869, n870, n871, n872,
         n873, n874, n875, n876, n877, n878, n879, n880, n881, n882, n883,
         n884, n885, n886, n887, n888, n889, n890, n891, n892, n893, n894,
         n895, n896, n897, n898, n899, n900, n901, n902, n903, n904, n905,
         n906, n907, n908, n909, n910, n911, n912, n913, n914, n915, n916,
         n917, n918, n919, n920, n921, n922, n923, n924, n925, n926, n927,
         n928, n929, n930, n931, n932, n933, n934, n935, n936, n937, n938,
         n939, n940, n941, n942, n943, n944, n945, n946, n947, n948, n949,
         n950, n951, n952, n953, n954, n955, n956, n957, n958, n959, n960,
         n961, n962, n963, n964, n965, n966, n967, n968, n969, n970, n971,
         n972, n973, n974, n975, n976, n977, n978, n979, n980, n981, n982,
         n983, n984, n985, n986, n987, n988, n989, n990, n991, n992, n993,
         n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NAND2_X1 U547 ( .A1(n765), .A2(n688), .ZN(n736) );
  OR2_X1 U548 ( .A1(n758), .A2(n751), .ZN(n517) );
  OR2_X1 U549 ( .A1(n763), .A2(n762), .ZN(n518) );
  AND2_X1 U550 ( .A1(n812), .A2(n988), .ZN(n519) );
  INV_X1 U551 ( .A(KEYINPUT26), .ZN(n693) );
  XNOR2_X1 U552 ( .A(n694), .B(n693), .ZN(n696) );
  NOR2_X1 U553 ( .A1(n713), .A2(n712), .ZN(n714) );
  NAND2_X1 U554 ( .A1(n901), .A2(n517), .ZN(n752) );
  NOR2_X1 U555 ( .A1(G164), .A2(G1384), .ZN(n765) );
  NOR2_X1 U556 ( .A1(n799), .A2(n519), .ZN(n800) );
  NOR2_X1 U557 ( .A1(G651), .A2(n640), .ZN(n655) );
  INV_X1 U558 ( .A(G2104), .ZN(n524) );
  AND2_X1 U559 ( .A1(n524), .A2(G2105), .ZN(n876) );
  NAND2_X1 U560 ( .A1(G126), .A2(n876), .ZN(n522) );
  NAND2_X1 U561 ( .A1(G2104), .A2(G2105), .ZN(n520) );
  XOR2_X2 U562 ( .A(KEYINPUT66), .B(n520), .Z(n877) );
  NAND2_X1 U563 ( .A1(G114), .A2(n877), .ZN(n521) );
  NAND2_X1 U564 ( .A1(n522), .A2(n521), .ZN(n523) );
  XNOR2_X1 U565 ( .A(KEYINPUT90), .B(n523), .ZN(n531) );
  NOR2_X4 U566 ( .A1(G2105), .A2(n524), .ZN(n880) );
  NAND2_X1 U567 ( .A1(G102), .A2(n880), .ZN(n529) );
  XNOR2_X1 U568 ( .A(KEYINPUT68), .B(KEYINPUT17), .ZN(n526) );
  NOR2_X1 U569 ( .A1(G2105), .A2(G2104), .ZN(n525) );
  XNOR2_X1 U570 ( .A(n526), .B(n525), .ZN(n527) );
  XNOR2_X2 U571 ( .A(KEYINPUT67), .B(n527), .ZN(n881) );
  NAND2_X1 U572 ( .A1(G138), .A2(n881), .ZN(n528) );
  NAND2_X1 U573 ( .A1(n529), .A2(n528), .ZN(n530) );
  NOR2_X1 U574 ( .A1(n531), .A2(n530), .ZN(G164) );
  NAND2_X1 U575 ( .A1(G101), .A2(n880), .ZN(n532) );
  XNOR2_X1 U576 ( .A(n532), .B(KEYINPUT23), .ZN(n533) );
  XNOR2_X1 U577 ( .A(n533), .B(KEYINPUT65), .ZN(n535) );
  NAND2_X1 U578 ( .A1(G113), .A2(n877), .ZN(n534) );
  NAND2_X1 U579 ( .A1(n535), .A2(n534), .ZN(n539) );
  NAND2_X1 U580 ( .A1(G125), .A2(n876), .ZN(n537) );
  NAND2_X1 U581 ( .A1(G137), .A2(n881), .ZN(n536) );
  NAND2_X1 U582 ( .A1(n537), .A2(n536), .ZN(n538) );
  NOR2_X1 U583 ( .A1(n539), .A2(n538), .ZN(G160) );
  INV_X1 U584 ( .A(G651), .ZN(n544) );
  NOR2_X1 U585 ( .A1(G543), .A2(n544), .ZN(n540) );
  XOR2_X1 U586 ( .A(KEYINPUT1), .B(n540), .Z(n650) );
  NAND2_X1 U587 ( .A1(G65), .A2(n650), .ZN(n543) );
  NOR2_X1 U588 ( .A1(G543), .A2(G651), .ZN(n541) );
  XNOR2_X1 U589 ( .A(n541), .B(KEYINPUT64), .ZN(n651) );
  NAND2_X1 U590 ( .A1(G91), .A2(n651), .ZN(n542) );
  NAND2_X1 U591 ( .A1(n543), .A2(n542), .ZN(n548) );
  XOR2_X1 U592 ( .A(KEYINPUT0), .B(G543), .Z(n640) );
  NOR2_X1 U593 ( .A1(n640), .A2(n544), .ZN(n654) );
  NAND2_X1 U594 ( .A1(G78), .A2(n654), .ZN(n546) );
  NAND2_X1 U595 ( .A1(G53), .A2(n655), .ZN(n545) );
  NAND2_X1 U596 ( .A1(n546), .A2(n545), .ZN(n547) );
  OR2_X1 U597 ( .A1(n548), .A2(n547), .ZN(G299) );
  XOR2_X1 U598 ( .A(G2438), .B(G2454), .Z(n550) );
  XNOR2_X1 U599 ( .A(G2435), .B(G2430), .ZN(n549) );
  XNOR2_X1 U600 ( .A(n550), .B(n549), .ZN(n551) );
  XOR2_X1 U601 ( .A(n551), .B(KEYINPUT106), .Z(n553) );
  XNOR2_X1 U602 ( .A(G1341), .B(G1348), .ZN(n552) );
  XNOR2_X1 U603 ( .A(n553), .B(n552), .ZN(n557) );
  XOR2_X1 U604 ( .A(G2446), .B(G2451), .Z(n555) );
  XNOR2_X1 U605 ( .A(G2443), .B(G2427), .ZN(n554) );
  XNOR2_X1 U606 ( .A(n555), .B(n554), .ZN(n556) );
  XOR2_X1 U607 ( .A(n557), .B(n556), .Z(n558) );
  AND2_X1 U608 ( .A1(G14), .A2(n558), .ZN(G401) );
  NAND2_X1 U609 ( .A1(G64), .A2(n650), .ZN(n560) );
  NAND2_X1 U610 ( .A1(G52), .A2(n655), .ZN(n559) );
  NAND2_X1 U611 ( .A1(n560), .A2(n559), .ZN(n566) );
  NAND2_X1 U612 ( .A1(n654), .A2(G77), .ZN(n562) );
  NAND2_X1 U613 ( .A1(G90), .A2(n651), .ZN(n561) );
  NAND2_X1 U614 ( .A1(n562), .A2(n561), .ZN(n563) );
  XOR2_X1 U615 ( .A(KEYINPUT9), .B(n563), .Z(n564) );
  XNOR2_X1 U616 ( .A(KEYINPUT70), .B(n564), .ZN(n565) );
  NOR2_X1 U617 ( .A1(n566), .A2(n565), .ZN(G171) );
  AND2_X1 U618 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U619 ( .A(G132), .ZN(G219) );
  INV_X1 U620 ( .A(G82), .ZN(G220) );
  INV_X1 U621 ( .A(G120), .ZN(G236) );
  NAND2_X1 U622 ( .A1(n654), .A2(G75), .ZN(n567) );
  XOR2_X1 U623 ( .A(KEYINPUT83), .B(n567), .Z(n569) );
  NAND2_X1 U624 ( .A1(G88), .A2(n651), .ZN(n568) );
  NAND2_X1 U625 ( .A1(n569), .A2(n568), .ZN(n570) );
  XOR2_X1 U626 ( .A(KEYINPUT84), .B(n570), .Z(n574) );
  NAND2_X1 U627 ( .A1(G62), .A2(n650), .ZN(n572) );
  NAND2_X1 U628 ( .A1(G50), .A2(n655), .ZN(n571) );
  AND2_X1 U629 ( .A1(n572), .A2(n571), .ZN(n573) );
  NAND2_X1 U630 ( .A1(n574), .A2(n573), .ZN(G303) );
  NAND2_X1 U631 ( .A1(G7), .A2(G661), .ZN(n575) );
  XNOR2_X1 U632 ( .A(n575), .B(KEYINPUT10), .ZN(G223) );
  XOR2_X1 U633 ( .A(G223), .B(KEYINPUT72), .Z(n816) );
  NAND2_X1 U634 ( .A1(n816), .A2(G567), .ZN(n576) );
  XOR2_X1 U635 ( .A(KEYINPUT11), .B(n576), .Z(G234) );
  NAND2_X1 U636 ( .A1(G56), .A2(n650), .ZN(n577) );
  XOR2_X1 U637 ( .A(KEYINPUT14), .B(n577), .Z(n583) );
  NAND2_X1 U638 ( .A1(G81), .A2(n651), .ZN(n578) );
  XNOR2_X1 U639 ( .A(n578), .B(KEYINPUT12), .ZN(n580) );
  NAND2_X1 U640 ( .A1(G68), .A2(n654), .ZN(n579) );
  NAND2_X1 U641 ( .A1(n580), .A2(n579), .ZN(n581) );
  XOR2_X1 U642 ( .A(KEYINPUT13), .B(n581), .Z(n582) );
  NOR2_X1 U643 ( .A1(n583), .A2(n582), .ZN(n585) );
  NAND2_X1 U644 ( .A1(n655), .A2(G43), .ZN(n584) );
  NAND2_X1 U645 ( .A1(n585), .A2(n584), .ZN(n904) );
  INV_X1 U646 ( .A(G860), .ZN(n610) );
  OR2_X1 U647 ( .A1(n904), .A2(n610), .ZN(n586) );
  XOR2_X1 U648 ( .A(KEYINPUT73), .B(n586), .Z(G153) );
  INV_X1 U649 ( .A(G171), .ZN(G301) );
  NAND2_X1 U650 ( .A1(G868), .A2(G301), .ZN(n597) );
  NAND2_X1 U651 ( .A1(G54), .A2(n655), .ZN(n593) );
  NAND2_X1 U652 ( .A1(G66), .A2(n650), .ZN(n588) );
  NAND2_X1 U653 ( .A1(G92), .A2(n651), .ZN(n587) );
  NAND2_X1 U654 ( .A1(n588), .A2(n587), .ZN(n591) );
  NAND2_X1 U655 ( .A1(n654), .A2(G79), .ZN(n589) );
  XOR2_X1 U656 ( .A(KEYINPUT74), .B(n589), .Z(n590) );
  NOR2_X1 U657 ( .A1(n591), .A2(n590), .ZN(n592) );
  NAND2_X1 U658 ( .A1(n593), .A2(n592), .ZN(n594) );
  XNOR2_X1 U659 ( .A(n594), .B(KEYINPUT15), .ZN(n595) );
  XNOR2_X1 U660 ( .A(KEYINPUT75), .B(n595), .ZN(n905) );
  INV_X1 U661 ( .A(G868), .ZN(n670) );
  NAND2_X1 U662 ( .A1(n905), .A2(n670), .ZN(n596) );
  NAND2_X1 U663 ( .A1(n597), .A2(n596), .ZN(G284) );
  NAND2_X1 U664 ( .A1(G89), .A2(n651), .ZN(n598) );
  XNOR2_X1 U665 ( .A(n598), .B(KEYINPUT4), .ZN(n600) );
  NAND2_X1 U666 ( .A1(G76), .A2(n654), .ZN(n599) );
  NAND2_X1 U667 ( .A1(n600), .A2(n599), .ZN(n601) );
  XNOR2_X1 U668 ( .A(n601), .B(KEYINPUT5), .ZN(n606) );
  NAND2_X1 U669 ( .A1(G63), .A2(n650), .ZN(n603) );
  NAND2_X1 U670 ( .A1(G51), .A2(n655), .ZN(n602) );
  NAND2_X1 U671 ( .A1(n603), .A2(n602), .ZN(n604) );
  XOR2_X1 U672 ( .A(KEYINPUT6), .B(n604), .Z(n605) );
  NAND2_X1 U673 ( .A1(n606), .A2(n605), .ZN(n607) );
  XNOR2_X1 U674 ( .A(n607), .B(KEYINPUT7), .ZN(G168) );
  XOR2_X1 U675 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NOR2_X1 U676 ( .A1(G286), .A2(n670), .ZN(n609) );
  NOR2_X1 U677 ( .A1(G868), .A2(G299), .ZN(n608) );
  NOR2_X1 U678 ( .A1(n609), .A2(n608), .ZN(G297) );
  NAND2_X1 U679 ( .A1(n610), .A2(G559), .ZN(n611) );
  INV_X1 U680 ( .A(n905), .ZN(n826) );
  NAND2_X1 U681 ( .A1(n611), .A2(n826), .ZN(n612) );
  XNOR2_X1 U682 ( .A(n612), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U683 ( .A1(G868), .A2(n904), .ZN(n615) );
  NAND2_X1 U684 ( .A1(G868), .A2(n826), .ZN(n613) );
  NOR2_X1 U685 ( .A1(G559), .A2(n613), .ZN(n614) );
  NOR2_X1 U686 ( .A1(n615), .A2(n614), .ZN(n616) );
  XNOR2_X1 U687 ( .A(KEYINPUT76), .B(n616), .ZN(G282) );
  NAND2_X1 U688 ( .A1(G123), .A2(n876), .ZN(n617) );
  XNOR2_X1 U689 ( .A(n617), .B(KEYINPUT18), .ZN(n620) );
  NAND2_X1 U690 ( .A1(n881), .A2(G135), .ZN(n618) );
  XOR2_X1 U691 ( .A(KEYINPUT77), .B(n618), .Z(n619) );
  NAND2_X1 U692 ( .A1(n620), .A2(n619), .ZN(n624) );
  NAND2_X1 U693 ( .A1(n880), .A2(G99), .ZN(n622) );
  NAND2_X1 U694 ( .A1(G111), .A2(n877), .ZN(n621) );
  NAND2_X1 U695 ( .A1(n622), .A2(n621), .ZN(n623) );
  NOR2_X1 U696 ( .A1(n624), .A2(n623), .ZN(n986) );
  XOR2_X1 U697 ( .A(G2096), .B(n986), .Z(n625) );
  NOR2_X1 U698 ( .A1(G2100), .A2(n625), .ZN(n626) );
  XOR2_X1 U699 ( .A(KEYINPUT78), .B(n626), .Z(G156) );
  NAND2_X1 U700 ( .A1(n651), .A2(G86), .ZN(n635) );
  NAND2_X1 U701 ( .A1(G73), .A2(n654), .ZN(n627) );
  XNOR2_X1 U702 ( .A(n627), .B(KEYINPUT2), .ZN(n630) );
  NAND2_X1 U703 ( .A1(G61), .A2(n650), .ZN(n628) );
  XNOR2_X1 U704 ( .A(n628), .B(KEYINPUT80), .ZN(n629) );
  NAND2_X1 U705 ( .A1(n630), .A2(n629), .ZN(n633) );
  NAND2_X1 U706 ( .A1(G48), .A2(n655), .ZN(n631) );
  XNOR2_X1 U707 ( .A(KEYINPUT81), .B(n631), .ZN(n632) );
  NOR2_X1 U708 ( .A1(n633), .A2(n632), .ZN(n634) );
  NAND2_X1 U709 ( .A1(n635), .A2(n634), .ZN(n636) );
  XNOR2_X1 U710 ( .A(n636), .B(KEYINPUT82), .ZN(G305) );
  NAND2_X1 U711 ( .A1(G49), .A2(n655), .ZN(n638) );
  NAND2_X1 U712 ( .A1(G74), .A2(G651), .ZN(n637) );
  NAND2_X1 U713 ( .A1(n638), .A2(n637), .ZN(n639) );
  NOR2_X1 U714 ( .A1(n650), .A2(n639), .ZN(n642) );
  NAND2_X1 U715 ( .A1(n640), .A2(G87), .ZN(n641) );
  NAND2_X1 U716 ( .A1(n642), .A2(n641), .ZN(G288) );
  NAND2_X1 U717 ( .A1(n654), .A2(G72), .ZN(n644) );
  NAND2_X1 U718 ( .A1(G85), .A2(n651), .ZN(n643) );
  NAND2_X1 U719 ( .A1(n644), .A2(n643), .ZN(n648) );
  NAND2_X1 U720 ( .A1(G60), .A2(n650), .ZN(n646) );
  NAND2_X1 U721 ( .A1(G47), .A2(n655), .ZN(n645) );
  NAND2_X1 U722 ( .A1(n646), .A2(n645), .ZN(n647) );
  NOR2_X1 U723 ( .A1(n648), .A2(n647), .ZN(n649) );
  XNOR2_X1 U724 ( .A(KEYINPUT69), .B(n649), .ZN(G290) );
  XNOR2_X1 U725 ( .A(G305), .B(G303), .ZN(n666) );
  XNOR2_X1 U726 ( .A(KEYINPUT85), .B(KEYINPUT19), .ZN(n662) );
  NAND2_X1 U727 ( .A1(G67), .A2(n650), .ZN(n653) );
  NAND2_X1 U728 ( .A1(G93), .A2(n651), .ZN(n652) );
  NAND2_X1 U729 ( .A1(n653), .A2(n652), .ZN(n659) );
  NAND2_X1 U730 ( .A1(G80), .A2(n654), .ZN(n657) );
  NAND2_X1 U731 ( .A1(G55), .A2(n655), .ZN(n656) );
  NAND2_X1 U732 ( .A1(n657), .A2(n656), .ZN(n658) );
  NOR2_X1 U733 ( .A1(n659), .A2(n658), .ZN(n660) );
  XNOR2_X1 U734 ( .A(KEYINPUT79), .B(n660), .ZN(n823) );
  XOR2_X1 U735 ( .A(G288), .B(n823), .Z(n661) );
  XNOR2_X1 U736 ( .A(n662), .B(n661), .ZN(n663) );
  XOR2_X1 U737 ( .A(n663), .B(G290), .Z(n664) );
  XNOR2_X1 U738 ( .A(G299), .B(n664), .ZN(n665) );
  XNOR2_X1 U739 ( .A(n666), .B(n665), .ZN(n825) );
  NAND2_X1 U740 ( .A1(G559), .A2(n826), .ZN(n667) );
  XNOR2_X1 U741 ( .A(n667), .B(n904), .ZN(n822) );
  XNOR2_X1 U742 ( .A(n825), .B(n822), .ZN(n668) );
  NAND2_X1 U743 ( .A1(n668), .A2(G868), .ZN(n669) );
  XNOR2_X1 U744 ( .A(n669), .B(KEYINPUT86), .ZN(n672) );
  NAND2_X1 U745 ( .A1(n670), .A2(n823), .ZN(n671) );
  NAND2_X1 U746 ( .A1(n672), .A2(n671), .ZN(G295) );
  NAND2_X1 U747 ( .A1(G2078), .A2(G2084), .ZN(n673) );
  XOR2_X1 U748 ( .A(KEYINPUT20), .B(n673), .Z(n674) );
  NAND2_X1 U749 ( .A1(G2090), .A2(n674), .ZN(n675) );
  XNOR2_X1 U750 ( .A(KEYINPUT21), .B(n675), .ZN(n676) );
  NAND2_X1 U751 ( .A1(n676), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U752 ( .A(KEYINPUT71), .B(G57), .ZN(G237) );
  XOR2_X1 U753 ( .A(KEYINPUT87), .B(G44), .Z(n677) );
  XNOR2_X1 U754 ( .A(KEYINPUT3), .B(n677), .ZN(G218) );
  NOR2_X1 U755 ( .A1(G237), .A2(G236), .ZN(n678) );
  NAND2_X1 U756 ( .A1(G69), .A2(n678), .ZN(n679) );
  XNOR2_X1 U757 ( .A(KEYINPUT89), .B(n679), .ZN(n680) );
  NAND2_X1 U758 ( .A1(n680), .A2(G108), .ZN(n820) );
  NAND2_X1 U759 ( .A1(n820), .A2(G567), .ZN(n686) );
  NOR2_X1 U760 ( .A1(G220), .A2(G219), .ZN(n681) );
  XNOR2_X1 U761 ( .A(KEYINPUT22), .B(n681), .ZN(n682) );
  NAND2_X1 U762 ( .A1(n682), .A2(G96), .ZN(n683) );
  NOR2_X1 U763 ( .A1(G218), .A2(n683), .ZN(n684) );
  XOR2_X1 U764 ( .A(KEYINPUT88), .B(n684), .Z(n821) );
  NAND2_X1 U765 ( .A1(n821), .A2(G2106), .ZN(n685) );
  NAND2_X1 U766 ( .A1(n686), .A2(n685), .ZN(n899) );
  NAND2_X1 U767 ( .A1(G483), .A2(G661), .ZN(n687) );
  NOR2_X1 U768 ( .A1(n899), .A2(n687), .ZN(n819) );
  NAND2_X1 U769 ( .A1(n819), .A2(G36), .ZN(G176) );
  NAND2_X1 U770 ( .A1(G160), .A2(G40), .ZN(n764) );
  INV_X1 U771 ( .A(n764), .ZN(n688) );
  NAND2_X1 U772 ( .A1(G8), .A2(n736), .ZN(n758) );
  NOR2_X1 U773 ( .A1(G1981), .A2(G305), .ZN(n689) );
  XOR2_X1 U774 ( .A(n689), .B(KEYINPUT24), .Z(n690) );
  NOR2_X1 U775 ( .A1(n758), .A2(n690), .ZN(n763) );
  NOR2_X1 U776 ( .A1(G2084), .A2(n736), .ZN(n720) );
  NAND2_X1 U777 ( .A1(G8), .A2(n720), .ZN(n734) );
  NOR2_X1 U778 ( .A1(G1966), .A2(n758), .ZN(n732) );
  NAND2_X1 U779 ( .A1(G1348), .A2(n736), .ZN(n692) );
  INV_X1 U780 ( .A(n736), .ZN(n715) );
  NAND2_X1 U781 ( .A1(G2067), .A2(n715), .ZN(n691) );
  NAND2_X1 U782 ( .A1(n692), .A2(n691), .ZN(n700) );
  NOR2_X1 U783 ( .A1(n905), .A2(n700), .ZN(n699) );
  AND2_X1 U784 ( .A1(n715), .A2(G1996), .ZN(n694) );
  NAND2_X1 U785 ( .A1(n736), .A2(G1341), .ZN(n695) );
  NAND2_X1 U786 ( .A1(n696), .A2(n695), .ZN(n697) );
  NOR2_X1 U787 ( .A1(n697), .A2(n904), .ZN(n698) );
  NOR2_X1 U788 ( .A1(n699), .A2(n698), .ZN(n702) );
  AND2_X1 U789 ( .A1(n905), .A2(n700), .ZN(n701) );
  NOR2_X1 U790 ( .A1(n702), .A2(n701), .ZN(n709) );
  INV_X1 U791 ( .A(G2072), .ZN(n981) );
  NOR2_X1 U792 ( .A1(n736), .A2(n981), .ZN(n704) );
  XNOR2_X1 U793 ( .A(KEYINPUT27), .B(KEYINPUT100), .ZN(n703) );
  XNOR2_X1 U794 ( .A(n704), .B(n703), .ZN(n706) );
  NAND2_X1 U795 ( .A1(n736), .A2(G1956), .ZN(n705) );
  NAND2_X1 U796 ( .A1(n706), .A2(n705), .ZN(n710) );
  NOR2_X1 U797 ( .A1(G299), .A2(n710), .ZN(n707) );
  XOR2_X1 U798 ( .A(KEYINPUT101), .B(n707), .Z(n708) );
  NOR2_X1 U799 ( .A1(n709), .A2(n708), .ZN(n713) );
  NAND2_X1 U800 ( .A1(G299), .A2(n710), .ZN(n711) );
  XOR2_X1 U801 ( .A(KEYINPUT28), .B(n711), .Z(n712) );
  XNOR2_X1 U802 ( .A(n714), .B(KEYINPUT29), .ZN(n719) );
  XNOR2_X1 U803 ( .A(G1961), .B(KEYINPUT99), .ZN(n926) );
  NAND2_X1 U804 ( .A1(n736), .A2(n926), .ZN(n717) );
  XNOR2_X1 U805 ( .A(G2078), .B(KEYINPUT25), .ZN(n957) );
  NAND2_X1 U806 ( .A1(n715), .A2(n957), .ZN(n716) );
  NAND2_X1 U807 ( .A1(n717), .A2(n716), .ZN(n724) );
  NAND2_X1 U808 ( .A1(G171), .A2(n724), .ZN(n718) );
  NAND2_X1 U809 ( .A1(n719), .A2(n718), .ZN(n729) );
  NOR2_X1 U810 ( .A1(n732), .A2(n720), .ZN(n721) );
  NAND2_X1 U811 ( .A1(G8), .A2(n721), .ZN(n722) );
  XNOR2_X1 U812 ( .A(KEYINPUT30), .B(n722), .ZN(n723) );
  NOR2_X1 U813 ( .A1(G168), .A2(n723), .ZN(n726) );
  NOR2_X1 U814 ( .A1(G171), .A2(n724), .ZN(n725) );
  NOR2_X1 U815 ( .A1(n726), .A2(n725), .ZN(n727) );
  XOR2_X1 U816 ( .A(KEYINPUT31), .B(n727), .Z(n728) );
  NAND2_X1 U817 ( .A1(n729), .A2(n728), .ZN(n730) );
  XNOR2_X1 U818 ( .A(n730), .B(KEYINPUT102), .ZN(n735) );
  INV_X1 U819 ( .A(n735), .ZN(n731) );
  NOR2_X1 U820 ( .A1(n732), .A2(n731), .ZN(n733) );
  NAND2_X1 U821 ( .A1(n734), .A2(n733), .ZN(n745) );
  NAND2_X1 U822 ( .A1(n735), .A2(G286), .ZN(n741) );
  NOR2_X1 U823 ( .A1(G1971), .A2(n758), .ZN(n738) );
  NOR2_X1 U824 ( .A1(G2090), .A2(n736), .ZN(n737) );
  NOR2_X1 U825 ( .A1(n738), .A2(n737), .ZN(n739) );
  NAND2_X1 U826 ( .A1(n739), .A2(G303), .ZN(n740) );
  NAND2_X1 U827 ( .A1(n741), .A2(n740), .ZN(n742) );
  NAND2_X1 U828 ( .A1(n742), .A2(G8), .ZN(n743) );
  XNOR2_X1 U829 ( .A(n743), .B(KEYINPUT32), .ZN(n744) );
  NAND2_X1 U830 ( .A1(n745), .A2(n744), .ZN(n756) );
  NOR2_X1 U831 ( .A1(G1976), .A2(G288), .ZN(n750) );
  NOR2_X1 U832 ( .A1(G1971), .A2(G303), .ZN(n746) );
  NOR2_X1 U833 ( .A1(n750), .A2(n746), .ZN(n916) );
  NAND2_X1 U834 ( .A1(n756), .A2(n916), .ZN(n747) );
  NAND2_X1 U835 ( .A1(G1976), .A2(G288), .ZN(n909) );
  NAND2_X1 U836 ( .A1(n747), .A2(n909), .ZN(n748) );
  NOR2_X1 U837 ( .A1(n748), .A2(n758), .ZN(n749) );
  NOR2_X1 U838 ( .A1(KEYINPUT33), .A2(n749), .ZN(n753) );
  XOR2_X1 U839 ( .A(G1981), .B(G305), .Z(n901) );
  NAND2_X1 U840 ( .A1(n750), .A2(KEYINPUT33), .ZN(n751) );
  OR2_X1 U841 ( .A1(n753), .A2(n752), .ZN(n761) );
  NOR2_X1 U842 ( .A1(G2090), .A2(G303), .ZN(n754) );
  NAND2_X1 U843 ( .A1(G8), .A2(n754), .ZN(n755) );
  NAND2_X1 U844 ( .A1(n756), .A2(n755), .ZN(n757) );
  XOR2_X1 U845 ( .A(KEYINPUT103), .B(n757), .Z(n759) );
  NAND2_X1 U846 ( .A1(n759), .A2(n758), .ZN(n760) );
  NAND2_X1 U847 ( .A1(n761), .A2(n760), .ZN(n762) );
  XNOR2_X1 U848 ( .A(G1986), .B(G290), .ZN(n908) );
  NOR2_X1 U849 ( .A1(n765), .A2(n764), .ZN(n766) );
  XOR2_X1 U850 ( .A(KEYINPUT91), .B(n766), .Z(n812) );
  NAND2_X1 U851 ( .A1(n908), .A2(n812), .ZN(n767) );
  XNOR2_X1 U852 ( .A(n767), .B(KEYINPUT92), .ZN(n780) );
  NAND2_X1 U853 ( .A1(G104), .A2(n880), .ZN(n769) );
  NAND2_X1 U854 ( .A1(G140), .A2(n881), .ZN(n768) );
  NAND2_X1 U855 ( .A1(n769), .A2(n768), .ZN(n770) );
  XNOR2_X1 U856 ( .A(KEYINPUT34), .B(n770), .ZN(n777) );
  XNOR2_X1 U857 ( .A(KEYINPUT94), .B(KEYINPUT35), .ZN(n775) );
  NAND2_X1 U858 ( .A1(n876), .A2(G128), .ZN(n773) );
  NAND2_X1 U859 ( .A1(G116), .A2(n877), .ZN(n771) );
  XOR2_X1 U860 ( .A(KEYINPUT93), .B(n771), .Z(n772) );
  NAND2_X1 U861 ( .A1(n773), .A2(n772), .ZN(n774) );
  XOR2_X1 U862 ( .A(n775), .B(n774), .Z(n776) );
  NOR2_X1 U863 ( .A1(n777), .A2(n776), .ZN(n778) );
  XNOR2_X1 U864 ( .A(KEYINPUT36), .B(n778), .ZN(n866) );
  XNOR2_X1 U865 ( .A(KEYINPUT37), .B(G2067), .ZN(n808) );
  NOR2_X1 U866 ( .A1(n866), .A2(n808), .ZN(n779) );
  XOR2_X1 U867 ( .A(KEYINPUT95), .B(n779), .Z(n999) );
  NAND2_X1 U868 ( .A1(n812), .A2(n999), .ZN(n806) );
  NAND2_X1 U869 ( .A1(n780), .A2(n806), .ZN(n799) );
  NAND2_X1 U870 ( .A1(G119), .A2(n876), .ZN(n782) );
  NAND2_X1 U871 ( .A1(G107), .A2(n877), .ZN(n781) );
  NAND2_X1 U872 ( .A1(n782), .A2(n781), .ZN(n785) );
  NAND2_X1 U873 ( .A1(n880), .A2(G95), .ZN(n783) );
  XOR2_X1 U874 ( .A(KEYINPUT96), .B(n783), .Z(n784) );
  NOR2_X1 U875 ( .A1(n785), .A2(n784), .ZN(n787) );
  NAND2_X1 U876 ( .A1(G131), .A2(n881), .ZN(n786) );
  NAND2_X1 U877 ( .A1(n787), .A2(n786), .ZN(n868) );
  NAND2_X1 U878 ( .A1(G1991), .A2(n868), .ZN(n798) );
  XOR2_X1 U879 ( .A(KEYINPUT98), .B(KEYINPUT38), .Z(n789) );
  NAND2_X1 U880 ( .A1(G105), .A2(n880), .ZN(n788) );
  XNOR2_X1 U881 ( .A(n789), .B(n788), .ZN(n794) );
  NAND2_X1 U882 ( .A1(G129), .A2(n876), .ZN(n791) );
  NAND2_X1 U883 ( .A1(G117), .A2(n877), .ZN(n790) );
  NAND2_X1 U884 ( .A1(n791), .A2(n790), .ZN(n792) );
  XOR2_X1 U885 ( .A(KEYINPUT97), .B(n792), .Z(n793) );
  NOR2_X1 U886 ( .A1(n794), .A2(n793), .ZN(n796) );
  NAND2_X1 U887 ( .A1(G141), .A2(n881), .ZN(n795) );
  NAND2_X1 U888 ( .A1(n796), .A2(n795), .ZN(n887) );
  NAND2_X1 U889 ( .A1(G1996), .A2(n887), .ZN(n797) );
  NAND2_X1 U890 ( .A1(n798), .A2(n797), .ZN(n988) );
  NAND2_X1 U891 ( .A1(n518), .A2(n800), .ZN(n814) );
  NOR2_X1 U892 ( .A1(G1996), .A2(n887), .ZN(n992) );
  NOR2_X1 U893 ( .A1(n868), .A2(G1991), .ZN(n801) );
  XNOR2_X1 U894 ( .A(n801), .B(KEYINPUT104), .ZN(n987) );
  NOR2_X1 U895 ( .A1(G1986), .A2(G290), .ZN(n802) );
  NOR2_X1 U896 ( .A1(n987), .A2(n802), .ZN(n803) );
  NOR2_X1 U897 ( .A1(n519), .A2(n803), .ZN(n804) );
  NOR2_X1 U898 ( .A1(n992), .A2(n804), .ZN(n805) );
  XNOR2_X1 U899 ( .A(n805), .B(KEYINPUT39), .ZN(n807) );
  NAND2_X1 U900 ( .A1(n807), .A2(n806), .ZN(n810) );
  NAND2_X1 U901 ( .A1(n866), .A2(n808), .ZN(n809) );
  XOR2_X1 U902 ( .A(KEYINPUT105), .B(n809), .Z(n996) );
  NAND2_X1 U903 ( .A1(n810), .A2(n996), .ZN(n811) );
  NAND2_X1 U904 ( .A1(n812), .A2(n811), .ZN(n813) );
  NAND2_X1 U905 ( .A1(n814), .A2(n813), .ZN(n815) );
  XNOR2_X1 U906 ( .A(KEYINPUT40), .B(n815), .ZN(G329) );
  NAND2_X1 U907 ( .A1(G2106), .A2(n816), .ZN(G217) );
  AND2_X1 U908 ( .A1(G15), .A2(G2), .ZN(n817) );
  NAND2_X1 U909 ( .A1(G661), .A2(n817), .ZN(G259) );
  NAND2_X1 U910 ( .A1(G3), .A2(G1), .ZN(n818) );
  NAND2_X1 U911 ( .A1(n819), .A2(n818), .ZN(G188) );
  INV_X1 U913 ( .A(G108), .ZN(G238) );
  INV_X1 U914 ( .A(G96), .ZN(G221) );
  NOR2_X1 U915 ( .A1(n821), .A2(n820), .ZN(G325) );
  INV_X1 U916 ( .A(G325), .ZN(G261) );
  NOR2_X1 U917 ( .A1(n822), .A2(G860), .ZN(n824) );
  XOR2_X1 U918 ( .A(n824), .B(n823), .Z(G145) );
  XOR2_X1 U919 ( .A(n825), .B(G286), .Z(n828) );
  XNOR2_X1 U920 ( .A(G171), .B(n826), .ZN(n827) );
  XNOR2_X1 U921 ( .A(n828), .B(n827), .ZN(n829) );
  XNOR2_X1 U922 ( .A(n829), .B(n904), .ZN(n830) );
  NOR2_X1 U923 ( .A1(G37), .A2(n830), .ZN(G397) );
  XOR2_X1 U924 ( .A(KEYINPUT108), .B(G2678), .Z(n832) );
  XNOR2_X1 U925 ( .A(KEYINPUT107), .B(KEYINPUT43), .ZN(n831) );
  XNOR2_X1 U926 ( .A(n832), .B(n831), .ZN(n836) );
  XOR2_X1 U927 ( .A(KEYINPUT42), .B(G2090), .Z(n834) );
  XNOR2_X1 U928 ( .A(G2067), .B(G2072), .ZN(n833) );
  XNOR2_X1 U929 ( .A(n834), .B(n833), .ZN(n835) );
  XOR2_X1 U930 ( .A(n836), .B(n835), .Z(n838) );
  XNOR2_X1 U931 ( .A(G2096), .B(G2100), .ZN(n837) );
  XNOR2_X1 U932 ( .A(n838), .B(n837), .ZN(n840) );
  XOR2_X1 U933 ( .A(G2078), .B(G2084), .Z(n839) );
  XNOR2_X1 U934 ( .A(n840), .B(n839), .ZN(G227) );
  XOR2_X1 U935 ( .A(G1981), .B(G1961), .Z(n842) );
  XNOR2_X1 U936 ( .A(G1996), .B(G1966), .ZN(n841) );
  XNOR2_X1 U937 ( .A(n842), .B(n841), .ZN(n846) );
  XOR2_X1 U938 ( .A(G1976), .B(G1971), .Z(n844) );
  XNOR2_X1 U939 ( .A(G1986), .B(G1956), .ZN(n843) );
  XNOR2_X1 U940 ( .A(n844), .B(n843), .ZN(n845) );
  XOR2_X1 U941 ( .A(n846), .B(n845), .Z(n848) );
  XNOR2_X1 U942 ( .A(KEYINPUT109), .B(G2474), .ZN(n847) );
  XNOR2_X1 U943 ( .A(n848), .B(n847), .ZN(n850) );
  XOR2_X1 U944 ( .A(G1991), .B(KEYINPUT41), .Z(n849) );
  XNOR2_X1 U945 ( .A(n850), .B(n849), .ZN(G229) );
  NAND2_X1 U946 ( .A1(n876), .A2(G124), .ZN(n851) );
  XNOR2_X1 U947 ( .A(n851), .B(KEYINPUT44), .ZN(n853) );
  NAND2_X1 U948 ( .A1(G100), .A2(n880), .ZN(n852) );
  NAND2_X1 U949 ( .A1(n853), .A2(n852), .ZN(n857) );
  NAND2_X1 U950 ( .A1(G112), .A2(n877), .ZN(n855) );
  NAND2_X1 U951 ( .A1(G136), .A2(n881), .ZN(n854) );
  NAND2_X1 U952 ( .A1(n855), .A2(n854), .ZN(n856) );
  NOR2_X1 U953 ( .A1(n857), .A2(n856), .ZN(G162) );
  NAND2_X1 U954 ( .A1(G103), .A2(n880), .ZN(n859) );
  NAND2_X1 U955 ( .A1(G139), .A2(n881), .ZN(n858) );
  NAND2_X1 U956 ( .A1(n859), .A2(n858), .ZN(n864) );
  NAND2_X1 U957 ( .A1(G127), .A2(n876), .ZN(n861) );
  NAND2_X1 U958 ( .A1(G115), .A2(n877), .ZN(n860) );
  NAND2_X1 U959 ( .A1(n861), .A2(n860), .ZN(n862) );
  XOR2_X1 U960 ( .A(KEYINPUT47), .B(n862), .Z(n863) );
  NOR2_X1 U961 ( .A1(n864), .A2(n863), .ZN(n980) );
  XOR2_X1 U962 ( .A(n986), .B(n980), .Z(n865) );
  XNOR2_X1 U963 ( .A(n866), .B(n865), .ZN(n870) );
  XOR2_X1 U964 ( .A(G160), .B(G162), .Z(n867) );
  XNOR2_X1 U965 ( .A(n868), .B(n867), .ZN(n869) );
  XOR2_X1 U966 ( .A(n870), .B(n869), .Z(n875) );
  XOR2_X1 U967 ( .A(KEYINPUT111), .B(KEYINPUT110), .Z(n872) );
  XNOR2_X1 U968 ( .A(KEYINPUT112), .B(KEYINPUT48), .ZN(n871) );
  XNOR2_X1 U969 ( .A(n872), .B(n871), .ZN(n873) );
  XNOR2_X1 U970 ( .A(KEYINPUT46), .B(n873), .ZN(n874) );
  XNOR2_X1 U971 ( .A(n875), .B(n874), .ZN(n891) );
  NAND2_X1 U972 ( .A1(G130), .A2(n876), .ZN(n879) );
  NAND2_X1 U973 ( .A1(G118), .A2(n877), .ZN(n878) );
  NAND2_X1 U974 ( .A1(n879), .A2(n878), .ZN(n886) );
  NAND2_X1 U975 ( .A1(G106), .A2(n880), .ZN(n883) );
  NAND2_X1 U976 ( .A1(G142), .A2(n881), .ZN(n882) );
  NAND2_X1 U977 ( .A1(n883), .A2(n882), .ZN(n884) );
  XOR2_X1 U978 ( .A(n884), .B(KEYINPUT45), .Z(n885) );
  NOR2_X1 U979 ( .A1(n886), .A2(n885), .ZN(n888) );
  XNOR2_X1 U980 ( .A(n888), .B(n887), .ZN(n889) );
  XOR2_X1 U981 ( .A(G164), .B(n889), .Z(n890) );
  XNOR2_X1 U982 ( .A(n891), .B(n890), .ZN(n892) );
  NOR2_X1 U983 ( .A1(G37), .A2(n892), .ZN(G395) );
  NOR2_X1 U984 ( .A1(G401), .A2(n899), .ZN(n896) );
  NOR2_X1 U985 ( .A1(G227), .A2(G229), .ZN(n893) );
  XNOR2_X1 U986 ( .A(KEYINPUT49), .B(n893), .ZN(n894) );
  NOR2_X1 U987 ( .A1(G397), .A2(n894), .ZN(n895) );
  NAND2_X1 U988 ( .A1(n896), .A2(n895), .ZN(n897) );
  NOR2_X1 U989 ( .A1(n897), .A2(G395), .ZN(n898) );
  XNOR2_X1 U990 ( .A(n898), .B(KEYINPUT113), .ZN(G225) );
  INV_X1 U991 ( .A(G225), .ZN(G308) );
  INV_X1 U992 ( .A(G303), .ZN(G166) );
  INV_X1 U993 ( .A(n899), .ZN(G319) );
  INV_X1 U994 ( .A(G69), .ZN(G235) );
  XNOR2_X1 U995 ( .A(G16), .B(KEYINPUT56), .ZN(n925) );
  XOR2_X1 U996 ( .A(G1966), .B(G168), .Z(n900) );
  XNOR2_X1 U997 ( .A(KEYINPUT121), .B(n900), .ZN(n902) );
  NAND2_X1 U998 ( .A1(n902), .A2(n901), .ZN(n903) );
  XNOR2_X1 U999 ( .A(n903), .B(KEYINPUT57), .ZN(n923) );
  XNOR2_X1 U1000 ( .A(n904), .B(G1341), .ZN(n921) );
  XNOR2_X1 U1001 ( .A(G1348), .B(KEYINPUT122), .ZN(n906) );
  XNOR2_X1 U1002 ( .A(n906), .B(n905), .ZN(n907) );
  NOR2_X1 U1003 ( .A1(n908), .A2(n907), .ZN(n914) );
  XNOR2_X1 U1004 ( .A(G171), .B(G1961), .ZN(n910) );
  NAND2_X1 U1005 ( .A1(n910), .A2(n909), .ZN(n912) );
  XNOR2_X1 U1006 ( .A(G1956), .B(G299), .ZN(n911) );
  NOR2_X1 U1007 ( .A1(n912), .A2(n911), .ZN(n913) );
  NAND2_X1 U1008 ( .A1(n914), .A2(n913), .ZN(n918) );
  NAND2_X1 U1009 ( .A1(G1971), .A2(G303), .ZN(n915) );
  NAND2_X1 U1010 ( .A1(n916), .A2(n915), .ZN(n917) );
  NOR2_X1 U1011 ( .A1(n918), .A2(n917), .ZN(n919) );
  XNOR2_X1 U1012 ( .A(KEYINPUT123), .B(n919), .ZN(n920) );
  NOR2_X1 U1013 ( .A1(n921), .A2(n920), .ZN(n922) );
  NAND2_X1 U1014 ( .A1(n923), .A2(n922), .ZN(n924) );
  NAND2_X1 U1015 ( .A1(n925), .A2(n924), .ZN(n952) );
  INV_X1 U1016 ( .A(G16), .ZN(n950) );
  XNOR2_X1 U1017 ( .A(G5), .B(n926), .ZN(n945) );
  XNOR2_X1 U1018 ( .A(G1341), .B(G19), .ZN(n928) );
  XNOR2_X1 U1019 ( .A(G1981), .B(G6), .ZN(n927) );
  NOR2_X1 U1020 ( .A1(n928), .A2(n927), .ZN(n929) );
  XOR2_X1 U1021 ( .A(KEYINPUT124), .B(n929), .Z(n931) );
  XNOR2_X1 U1022 ( .A(G1956), .B(G20), .ZN(n930) );
  NOR2_X1 U1023 ( .A1(n931), .A2(n930), .ZN(n935) );
  XOR2_X1 U1024 ( .A(G4), .B(KEYINPUT125), .Z(n933) );
  XNOR2_X1 U1025 ( .A(G1348), .B(KEYINPUT59), .ZN(n932) );
  XNOR2_X1 U1026 ( .A(n933), .B(n932), .ZN(n934) );
  NAND2_X1 U1027 ( .A1(n935), .A2(n934), .ZN(n936) );
  XNOR2_X1 U1028 ( .A(n936), .B(KEYINPUT60), .ZN(n943) );
  XNOR2_X1 U1029 ( .A(G1986), .B(G24), .ZN(n938) );
  XNOR2_X1 U1030 ( .A(G1971), .B(G22), .ZN(n937) );
  NOR2_X1 U1031 ( .A1(n938), .A2(n937), .ZN(n940) );
  XOR2_X1 U1032 ( .A(G1976), .B(G23), .Z(n939) );
  NAND2_X1 U1033 ( .A1(n940), .A2(n939), .ZN(n941) );
  XNOR2_X1 U1034 ( .A(KEYINPUT58), .B(n941), .ZN(n942) );
  NOR2_X1 U1035 ( .A1(n943), .A2(n942), .ZN(n944) );
  NAND2_X1 U1036 ( .A1(n945), .A2(n944), .ZN(n947) );
  XNOR2_X1 U1037 ( .A(G21), .B(G1966), .ZN(n946) );
  NOR2_X1 U1038 ( .A1(n947), .A2(n946), .ZN(n948) );
  XNOR2_X1 U1039 ( .A(KEYINPUT61), .B(n948), .ZN(n949) );
  NAND2_X1 U1040 ( .A1(n950), .A2(n949), .ZN(n951) );
  NAND2_X1 U1041 ( .A1(n952), .A2(n951), .ZN(n979) );
  XNOR2_X1 U1042 ( .A(G29), .B(KEYINPUT119), .ZN(n975) );
  XOR2_X1 U1043 ( .A(G2090), .B(G35), .Z(n956) );
  XOR2_X1 U1044 ( .A(G2084), .B(G34), .Z(n953) );
  XNOR2_X1 U1045 ( .A(KEYINPUT118), .B(n953), .ZN(n954) );
  XNOR2_X1 U1046 ( .A(n954), .B(KEYINPUT54), .ZN(n955) );
  NAND2_X1 U1047 ( .A1(n956), .A2(n955), .ZN(n972) );
  XNOR2_X1 U1048 ( .A(n957), .B(G27), .ZN(n968) );
  XOR2_X1 U1049 ( .A(G1991), .B(G25), .Z(n958) );
  NAND2_X1 U1050 ( .A1(G28), .A2(n958), .ZN(n959) );
  XNOR2_X1 U1051 ( .A(n959), .B(KEYINPUT115), .ZN(n963) );
  XNOR2_X1 U1052 ( .A(G2067), .B(G26), .ZN(n961) );
  XNOR2_X1 U1053 ( .A(G1996), .B(G32), .ZN(n960) );
  NOR2_X1 U1054 ( .A1(n961), .A2(n960), .ZN(n962) );
  NAND2_X1 U1055 ( .A1(n963), .A2(n962), .ZN(n966) );
  XOR2_X1 U1056 ( .A(KEYINPUT116), .B(n981), .Z(n964) );
  XNOR2_X1 U1057 ( .A(G33), .B(n964), .ZN(n965) );
  NOR2_X1 U1058 ( .A1(n966), .A2(n965), .ZN(n967) );
  NAND2_X1 U1059 ( .A1(n968), .A2(n967), .ZN(n969) );
  XNOR2_X1 U1060 ( .A(n969), .B(KEYINPUT117), .ZN(n970) );
  XNOR2_X1 U1061 ( .A(n970), .B(KEYINPUT53), .ZN(n971) );
  NOR2_X1 U1062 ( .A1(n972), .A2(n971), .ZN(n973) );
  XNOR2_X1 U1063 ( .A(KEYINPUT55), .B(n973), .ZN(n974) );
  NAND2_X1 U1064 ( .A1(n975), .A2(n974), .ZN(n976) );
  NAND2_X1 U1065 ( .A1(G11), .A2(n976), .ZN(n977) );
  XNOR2_X1 U1066 ( .A(KEYINPUT120), .B(n977), .ZN(n978) );
  NOR2_X1 U1067 ( .A1(n979), .A2(n978), .ZN(n1008) );
  XOR2_X1 U1068 ( .A(G164), .B(G2078), .Z(n983) );
  XNOR2_X1 U1069 ( .A(n981), .B(n980), .ZN(n982) );
  NOR2_X1 U1070 ( .A1(n983), .A2(n982), .ZN(n984) );
  XOR2_X1 U1071 ( .A(KEYINPUT50), .B(n984), .Z(n1002) );
  XOR2_X1 U1072 ( .A(G2084), .B(G160), .Z(n985) );
  NOR2_X1 U1073 ( .A1(n986), .A2(n985), .ZN(n990) );
  NOR2_X1 U1074 ( .A1(n988), .A2(n987), .ZN(n989) );
  NAND2_X1 U1075 ( .A1(n990), .A2(n989), .ZN(n995) );
  XOR2_X1 U1076 ( .A(G2090), .B(G162), .Z(n991) );
  NOR2_X1 U1077 ( .A1(n992), .A2(n991), .ZN(n993) );
  XNOR2_X1 U1078 ( .A(n993), .B(KEYINPUT51), .ZN(n994) );
  NOR2_X1 U1079 ( .A1(n995), .A2(n994), .ZN(n997) );
  NAND2_X1 U1080 ( .A1(n997), .A2(n996), .ZN(n998) );
  NOR2_X1 U1081 ( .A1(n999), .A2(n998), .ZN(n1000) );
  XOR2_X1 U1082 ( .A(KEYINPUT114), .B(n1000), .Z(n1001) );
  NOR2_X1 U1083 ( .A1(n1002), .A2(n1001), .ZN(n1003) );
  XNOR2_X1 U1084 ( .A(KEYINPUT52), .B(n1003), .ZN(n1005) );
  INV_X1 U1085 ( .A(KEYINPUT55), .ZN(n1004) );
  NAND2_X1 U1086 ( .A1(n1005), .A2(n1004), .ZN(n1006) );
  NAND2_X1 U1087 ( .A1(n1006), .A2(G29), .ZN(n1007) );
  NAND2_X1 U1088 ( .A1(n1008), .A2(n1007), .ZN(n1009) );
  XOR2_X1 U1089 ( .A(KEYINPUT62), .B(n1009), .Z(G311) );
  XOR2_X1 U1090 ( .A(KEYINPUT126), .B(G311), .Z(G150) );
endmodule

