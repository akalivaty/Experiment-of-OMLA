//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 1 0 0 1 0 1 1 0 0 1 0 0 0 1 0 1 1 0 1 1 0 1 0 1 1 0 0 0 1 1 0 1 0 0 0 0 1 1 0 0 1 1 0 1 1 0 1 1 1 1 0 1 1 1 1 0 1 0 1 0 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:42:45 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n205, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n597, new_n598,
    new_n599, new_n600, new_n601, new_n602, new_n603, new_n604, new_n605,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1184, new_n1185, new_n1186, new_n1187,
    new_n1188, new_n1189, new_n1190, new_n1191, new_n1192, new_n1193,
    new_n1194, new_n1195, new_n1196, new_n1197, new_n1198, new_n1199,
    new_n1200, new_n1201, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1217, new_n1219,
    new_n1220, new_n1221, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1307, new_n1308, new_n1309, new_n1310;
  INV_X1    g0000(.A(G50), .ZN(new_n201));
  INV_X1    g0001(.A(G58), .ZN(new_n202));
  INV_X1    g0002(.A(G68), .ZN(new_n203));
  INV_X1    g0003(.A(G77), .ZN(new_n204));
  NAND4_X1  g0004(.A1(new_n201), .A2(new_n202), .A3(new_n203), .A4(new_n204), .ZN(new_n205));
  XNOR2_X1  g0005(.A(new_n205), .B(KEYINPUT64), .ZN(G353));
  OAI21_X1  g0006(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0007(.A1(G1), .A2(G20), .ZN(new_n208));
  NOR2_X1   g0008(.A1(new_n208), .A2(G13), .ZN(new_n209));
  OAI211_X1 g0009(.A(new_n209), .B(G250), .C1(G257), .C2(G264), .ZN(new_n210));
  XNOR2_X1  g0010(.A(new_n210), .B(KEYINPUT0), .ZN(new_n211));
  NAND2_X1  g0011(.A1(G1), .A2(G13), .ZN(new_n212));
  INV_X1    g0012(.A(G20), .ZN(new_n213));
  NOR2_X1   g0013(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  XOR2_X1   g0014(.A(new_n214), .B(KEYINPUT65), .Z(new_n215));
  OAI21_X1  g0015(.A(G50), .B1(G58), .B2(G68), .ZN(new_n216));
  AOI22_X1  g0016(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n217));
  INV_X1    g0017(.A(G238), .ZN(new_n218));
  INV_X1    g0018(.A(G244), .ZN(new_n219));
  OAI221_X1 g0019(.A(new_n217), .B1(new_n203), .B2(new_n218), .C1(new_n204), .C2(new_n219), .ZN(new_n220));
  NAND2_X1  g0020(.A1(new_n220), .A2(KEYINPUT66), .ZN(new_n221));
  AOI22_X1  g0021(.A1(G87), .A2(G250), .B1(G107), .B2(G264), .ZN(new_n222));
  AOI22_X1  g0022(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n223));
  NAND3_X1  g0023(.A1(new_n221), .A2(new_n222), .A3(new_n223), .ZN(new_n224));
  NOR2_X1   g0024(.A1(new_n220), .A2(KEYINPUT66), .ZN(new_n225));
  OAI21_X1  g0025(.A(new_n208), .B1(new_n224), .B2(new_n225), .ZN(new_n226));
  OAI221_X1 g0026(.A(new_n211), .B1(new_n215), .B2(new_n216), .C1(new_n226), .C2(KEYINPUT1), .ZN(new_n227));
  AOI21_X1  g0027(.A(new_n227), .B1(KEYINPUT1), .B2(new_n226), .ZN(G361));
  XOR2_X1   g0028(.A(G238), .B(G244), .Z(new_n229));
  XNOR2_X1  g0029(.A(G226), .B(G232), .ZN(new_n230));
  XNOR2_X1  g0030(.A(new_n229), .B(new_n230), .ZN(new_n231));
  XNOR2_X1  g0031(.A(KEYINPUT67), .B(KEYINPUT2), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n231), .B(new_n232), .ZN(new_n233));
  XOR2_X1   g0033(.A(G264), .B(G270), .Z(new_n234));
  XNOR2_X1  g0034(.A(G250), .B(G257), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n233), .B(new_n236), .ZN(G358));
  XOR2_X1   g0037(.A(G87), .B(G97), .Z(new_n238));
  XOR2_X1   g0038(.A(G107), .B(G116), .Z(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n240), .B(KEYINPUT68), .ZN(new_n241));
  XOR2_X1   g0041(.A(G68), .B(G77), .Z(new_n242));
  XOR2_X1   g0042(.A(G50), .B(G58), .Z(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XOR2_X1   g0044(.A(new_n241), .B(new_n244), .Z(G351));
  NOR2_X1   g0045(.A1(new_n202), .A2(new_n203), .ZN(new_n246));
  NOR2_X1   g0046(.A1(G58), .A2(G68), .ZN(new_n247));
  OAI21_X1  g0047(.A(G20), .B1(new_n246), .B2(new_n247), .ZN(new_n248));
  NOR2_X1   g0048(.A1(G20), .A2(G33), .ZN(new_n249));
  NAND2_X1  g0049(.A1(new_n249), .A2(G159), .ZN(new_n250));
  NAND2_X1  g0050(.A1(new_n248), .A2(new_n250), .ZN(new_n251));
  INV_X1    g0051(.A(new_n251), .ZN(new_n252));
  INV_X1    g0052(.A(KEYINPUT3), .ZN(new_n253));
  INV_X1    g0053(.A(G33), .ZN(new_n254));
  NAND2_X1  g0054(.A1(new_n253), .A2(new_n254), .ZN(new_n255));
  NAND2_X1  g0055(.A1(KEYINPUT3), .A2(G33), .ZN(new_n256));
  NAND3_X1  g0056(.A1(new_n255), .A2(new_n213), .A3(new_n256), .ZN(new_n257));
  INV_X1    g0057(.A(KEYINPUT7), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  INV_X1    g0059(.A(KEYINPUT74), .ZN(new_n260));
  NAND4_X1  g0060(.A1(new_n255), .A2(KEYINPUT7), .A3(new_n213), .A4(new_n256), .ZN(new_n261));
  AND3_X1   g0061(.A1(new_n259), .A2(new_n260), .A3(new_n261), .ZN(new_n262));
  OAI21_X1  g0062(.A(G68), .B1(new_n261), .B2(new_n260), .ZN(new_n263));
  OAI211_X1 g0063(.A(KEYINPUT16), .B(new_n252), .C1(new_n262), .C2(new_n263), .ZN(new_n264));
  NAND3_X1  g0064(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n265), .A2(new_n212), .ZN(new_n266));
  INV_X1    g0066(.A(KEYINPUT16), .ZN(new_n267));
  AOI21_X1  g0067(.A(new_n203), .B1(new_n259), .B2(new_n261), .ZN(new_n268));
  OAI21_X1  g0068(.A(new_n267), .B1(new_n268), .B2(new_n251), .ZN(new_n269));
  NAND3_X1  g0069(.A1(new_n264), .A2(new_n266), .A3(new_n269), .ZN(new_n270));
  INV_X1    g0070(.A(KEYINPUT17), .ZN(new_n271));
  XNOR2_X1  g0071(.A(KEYINPUT8), .B(G58), .ZN(new_n272));
  INV_X1    g0072(.A(KEYINPUT70), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  OR3_X1    g0074(.A1(new_n273), .A2(new_n202), .A3(KEYINPUT8), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  INV_X1    g0076(.A(G1), .ZN(new_n277));
  NAND3_X1  g0077(.A1(new_n277), .A2(G13), .A3(G20), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n276), .A2(new_n278), .ZN(new_n279));
  AOI21_X1  g0079(.A(new_n266), .B1(new_n277), .B2(G20), .ZN(new_n280));
  OAI21_X1  g0080(.A(new_n279), .B1(new_n276), .B2(new_n280), .ZN(new_n281));
  INV_X1    g0081(.A(G226), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n282), .A2(G1698), .ZN(new_n283));
  AND2_X1   g0083(.A1(KEYINPUT3), .A2(G33), .ZN(new_n284));
  NOR2_X1   g0084(.A1(KEYINPUT3), .A2(G33), .ZN(new_n285));
  OAI221_X1 g0085(.A(new_n283), .B1(G223), .B2(G1698), .C1(new_n284), .C2(new_n285), .ZN(new_n286));
  NAND2_X1  g0086(.A1(G33), .A2(G87), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  AOI21_X1  g0088(.A(new_n212), .B1(G33), .B2(G41), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  INV_X1    g0090(.A(G190), .ZN(new_n291));
  OR2_X1    g0091(.A1(KEYINPUT69), .A2(G41), .ZN(new_n292));
  INV_X1    g0092(.A(G45), .ZN(new_n293));
  NAND2_X1  g0093(.A1(KEYINPUT69), .A2(G41), .ZN(new_n294));
  NAND3_X1  g0094(.A1(new_n292), .A2(new_n293), .A3(new_n294), .ZN(new_n295));
  INV_X1    g0095(.A(G274), .ZN(new_n296));
  NOR2_X1   g0096(.A1(new_n296), .A2(G1), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n295), .A2(new_n297), .ZN(new_n298));
  INV_X1    g0098(.A(G41), .ZN(new_n299));
  OAI211_X1 g0099(.A(G1), .B(G13), .C1(new_n254), .C2(new_n299), .ZN(new_n300));
  OAI21_X1  g0100(.A(new_n277), .B1(G41), .B2(G45), .ZN(new_n301));
  NAND3_X1  g0101(.A1(new_n300), .A2(G232), .A3(new_n301), .ZN(new_n302));
  AND2_X1   g0102(.A1(new_n298), .A2(new_n302), .ZN(new_n303));
  NAND3_X1  g0103(.A1(new_n290), .A2(new_n291), .A3(new_n303), .ZN(new_n304));
  INV_X1    g0104(.A(G200), .ZN(new_n305));
  AOI21_X1  g0105(.A(new_n300), .B1(new_n286), .B2(new_n287), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n298), .A2(new_n302), .ZN(new_n307));
  OAI21_X1  g0107(.A(new_n305), .B1(new_n306), .B2(new_n307), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n304), .A2(new_n308), .ZN(new_n309));
  NAND4_X1  g0109(.A1(new_n270), .A2(new_n271), .A3(new_n281), .A4(new_n309), .ZN(new_n310));
  INV_X1    g0110(.A(KEYINPUT76), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  INV_X1    g0112(.A(new_n281), .ZN(new_n313));
  INV_X1    g0113(.A(new_n266), .ZN(new_n314));
  NOR2_X1   g0114(.A1(new_n284), .A2(new_n285), .ZN(new_n315));
  AOI21_X1  g0115(.A(KEYINPUT7), .B1(new_n315), .B2(new_n213), .ZN(new_n316));
  INV_X1    g0116(.A(new_n261), .ZN(new_n317));
  OAI21_X1  g0117(.A(G68), .B1(new_n316), .B2(new_n317), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n318), .A2(new_n252), .ZN(new_n319));
  AOI21_X1  g0119(.A(new_n314), .B1(new_n319), .B2(new_n267), .ZN(new_n320));
  AOI21_X1  g0120(.A(new_n313), .B1(new_n320), .B2(new_n264), .ZN(new_n321));
  NAND4_X1  g0121(.A1(new_n321), .A2(KEYINPUT76), .A3(new_n271), .A4(new_n309), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n312), .A2(new_n322), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n269), .A2(new_n266), .ZN(new_n324));
  INV_X1    g0124(.A(new_n263), .ZN(new_n325));
  NAND3_X1  g0125(.A1(new_n259), .A2(new_n260), .A3(new_n261), .ZN(new_n326));
  AOI211_X1 g0126(.A(new_n267), .B(new_n251), .C1(new_n325), .C2(new_n326), .ZN(new_n327));
  OAI211_X1 g0127(.A(new_n281), .B(new_n309), .C1(new_n324), .C2(new_n327), .ZN(new_n328));
  INV_X1    g0128(.A(KEYINPUT75), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n328), .A2(new_n329), .ZN(new_n330));
  NAND4_X1  g0130(.A1(new_n270), .A2(KEYINPUT75), .A3(new_n281), .A4(new_n309), .ZN(new_n331));
  NAND3_X1  g0131(.A1(new_n330), .A2(KEYINPUT17), .A3(new_n331), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n323), .A2(new_n332), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n270), .A2(new_n281), .ZN(new_n334));
  INV_X1    g0134(.A(KEYINPUT18), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n290), .A2(new_n303), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n336), .A2(G169), .ZN(new_n337));
  INV_X1    g0137(.A(G179), .ZN(new_n338));
  OAI21_X1  g0138(.A(new_n337), .B1(new_n336), .B2(new_n338), .ZN(new_n339));
  AND3_X1   g0139(.A1(new_n334), .A2(new_n335), .A3(new_n339), .ZN(new_n340));
  AOI21_X1  g0140(.A(new_n335), .B1(new_n334), .B2(new_n339), .ZN(new_n341));
  NOR2_X1   g0141(.A1(new_n340), .A2(new_n341), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n333), .A2(new_n342), .ZN(new_n343));
  INV_X1    g0143(.A(new_n343), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n280), .A2(G50), .ZN(new_n345));
  OAI21_X1  g0145(.A(new_n345), .B1(G50), .B2(new_n278), .ZN(new_n346));
  INV_X1    g0146(.A(new_n276), .ZN(new_n347));
  NOR2_X1   g0147(.A1(new_n254), .A2(G20), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n347), .A2(new_n348), .ZN(new_n349));
  NAND3_X1  g0149(.A1(new_n201), .A2(new_n202), .A3(new_n203), .ZN(new_n350));
  AOI22_X1  g0150(.A1(new_n350), .A2(G20), .B1(G150), .B2(new_n249), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n349), .A2(new_n351), .ZN(new_n352));
  AOI21_X1  g0152(.A(new_n346), .B1(new_n266), .B2(new_n352), .ZN(new_n353));
  INV_X1    g0153(.A(KEYINPUT9), .ZN(new_n354));
  XNOR2_X1  g0154(.A(new_n353), .B(new_n354), .ZN(new_n355));
  INV_X1    g0155(.A(G1698), .ZN(new_n356));
  NOR2_X1   g0156(.A1(new_n315), .A2(new_n356), .ZN(new_n357));
  AOI22_X1  g0157(.A1(new_n357), .A2(G223), .B1(G77), .B2(new_n315), .ZN(new_n358));
  INV_X1    g0158(.A(G222), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n255), .A2(new_n256), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n360), .A2(new_n356), .ZN(new_n361));
  OAI21_X1  g0161(.A(new_n358), .B1(new_n359), .B2(new_n361), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n362), .A2(new_n289), .ZN(new_n363));
  AND2_X1   g0163(.A1(new_n300), .A2(new_n301), .ZN(new_n364));
  AOI22_X1  g0164(.A1(new_n364), .A2(G226), .B1(new_n295), .B2(new_n297), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n363), .A2(new_n365), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n366), .A2(G200), .ZN(new_n367));
  INV_X1    g0167(.A(KEYINPUT10), .ZN(new_n368));
  NOR2_X1   g0168(.A1(new_n368), .A2(KEYINPUT72), .ZN(new_n369));
  INV_X1    g0169(.A(new_n366), .ZN(new_n370));
  AOI21_X1  g0170(.A(new_n369), .B1(new_n370), .B2(G190), .ZN(new_n371));
  NAND3_X1  g0171(.A1(new_n355), .A2(new_n367), .A3(new_n371), .ZN(new_n372));
  NAND3_X1  g0172(.A1(new_n372), .A2(KEYINPUT72), .A3(new_n368), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n368), .A2(KEYINPUT72), .ZN(new_n374));
  NAND4_X1  g0174(.A1(new_n355), .A2(new_n374), .A3(new_n367), .A4(new_n371), .ZN(new_n375));
  INV_X1    g0175(.A(G169), .ZN(new_n376));
  AOI21_X1  g0176(.A(new_n353), .B1(new_n376), .B2(new_n366), .ZN(new_n377));
  OAI21_X1  g0177(.A(new_n377), .B1(G179), .B2(new_n366), .ZN(new_n378));
  AND3_X1   g0178(.A1(new_n373), .A2(new_n375), .A3(new_n378), .ZN(new_n379));
  NAND3_X1  g0179(.A1(new_n360), .A2(G232), .A3(G1698), .ZN(new_n380));
  NAND2_X1  g0180(.A1(G33), .A2(G97), .ZN(new_n381));
  OAI211_X1 g0181(.A(new_n380), .B(new_n381), .C1(new_n361), .C2(new_n282), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n382), .A2(new_n289), .ZN(new_n383));
  INV_X1    g0183(.A(KEYINPUT13), .ZN(new_n384));
  AOI22_X1  g0184(.A1(new_n364), .A2(G238), .B1(new_n295), .B2(new_n297), .ZN(new_n385));
  NAND3_X1  g0185(.A1(new_n383), .A2(new_n384), .A3(new_n385), .ZN(new_n386));
  INV_X1    g0186(.A(new_n386), .ZN(new_n387));
  AOI21_X1  g0187(.A(new_n384), .B1(new_n383), .B2(new_n385), .ZN(new_n388));
  OAI21_X1  g0188(.A(G169), .B1(new_n387), .B2(new_n388), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n389), .A2(KEYINPUT14), .ZN(new_n390));
  INV_X1    g0190(.A(KEYINPUT14), .ZN(new_n391));
  OAI211_X1 g0191(.A(new_n391), .B(G169), .C1(new_n387), .C2(new_n388), .ZN(new_n392));
  NOR2_X1   g0192(.A1(new_n387), .A2(new_n388), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n393), .A2(G179), .ZN(new_n394));
  NAND3_X1  g0194(.A1(new_n390), .A2(new_n392), .A3(new_n394), .ZN(new_n395));
  AOI22_X1  g0195(.A1(new_n348), .A2(G77), .B1(G20), .B2(new_n203), .ZN(new_n396));
  INV_X1    g0196(.A(new_n249), .ZN(new_n397));
  OAI21_X1  g0197(.A(new_n396), .B1(new_n201), .B2(new_n397), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n398), .A2(new_n266), .ZN(new_n399));
  INV_X1    g0199(.A(KEYINPUT11), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n399), .A2(new_n400), .ZN(new_n401));
  NAND3_X1  g0201(.A1(new_n398), .A2(KEYINPUT11), .A3(new_n266), .ZN(new_n402));
  INV_X1    g0202(.A(new_n278), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n403), .A2(new_n203), .ZN(new_n404));
  XNOR2_X1  g0204(.A(new_n404), .B(KEYINPUT12), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n280), .A2(G68), .ZN(new_n406));
  NAND4_X1  g0206(.A1(new_n401), .A2(new_n402), .A3(new_n405), .A4(new_n406), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n395), .A2(new_n407), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n364), .A2(G244), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n409), .A2(new_n298), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n315), .A2(G107), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n360), .A2(G1698), .ZN(new_n412));
  INV_X1    g0212(.A(G232), .ZN(new_n413));
  OAI221_X1 g0213(.A(new_n411), .B1(new_n412), .B2(new_n218), .C1(new_n413), .C2(new_n361), .ZN(new_n414));
  AOI21_X1  g0214(.A(new_n410), .B1(new_n414), .B2(new_n289), .ZN(new_n415));
  INV_X1    g0215(.A(new_n415), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n416), .A2(new_n376), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n415), .A2(new_n338), .ZN(new_n418));
  XNOR2_X1  g0218(.A(KEYINPUT15), .B(G87), .ZN(new_n419));
  INV_X1    g0219(.A(new_n419), .ZN(new_n420));
  AOI22_X1  g0220(.A1(new_n420), .A2(new_n348), .B1(G20), .B2(G77), .ZN(new_n421));
  OAI21_X1  g0221(.A(new_n421), .B1(new_n397), .B2(new_n272), .ZN(new_n422));
  AOI22_X1  g0222(.A1(new_n422), .A2(new_n266), .B1(new_n204), .B2(new_n403), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n280), .A2(G77), .ZN(new_n424));
  XNOR2_X1  g0224(.A(new_n424), .B(KEYINPUT71), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n423), .A2(new_n425), .ZN(new_n426));
  NAND3_X1  g0226(.A1(new_n417), .A2(new_n418), .A3(new_n426), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n416), .A2(G200), .ZN(new_n428));
  INV_X1    g0228(.A(new_n426), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n415), .A2(G190), .ZN(new_n430));
  NAND3_X1  g0230(.A1(new_n428), .A2(new_n429), .A3(new_n430), .ZN(new_n431));
  AND3_X1   g0231(.A1(new_n408), .A2(new_n427), .A3(new_n431), .ZN(new_n432));
  AOI21_X1  g0232(.A(new_n407), .B1(new_n393), .B2(G190), .ZN(new_n433));
  OAI21_X1  g0233(.A(G200), .B1(new_n387), .B2(new_n388), .ZN(new_n434));
  NAND3_X1  g0234(.A1(new_n433), .A2(KEYINPUT73), .A3(new_n434), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n383), .A2(new_n385), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n436), .A2(KEYINPUT13), .ZN(new_n437));
  NAND3_X1  g0237(.A1(new_n437), .A2(G190), .A3(new_n386), .ZN(new_n438));
  INV_X1    g0238(.A(new_n407), .ZN(new_n439));
  NAND3_X1  g0239(.A1(new_n434), .A2(new_n438), .A3(new_n439), .ZN(new_n440));
  INV_X1    g0240(.A(KEYINPUT73), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n440), .A2(new_n441), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n435), .A2(new_n442), .ZN(new_n443));
  AND4_X1   g0243(.A1(new_n344), .A2(new_n379), .A3(new_n432), .A4(new_n443), .ZN(new_n444));
  NAND3_X1  g0244(.A1(new_n277), .A2(new_n296), .A3(G45), .ZN(new_n445));
  INV_X1    g0245(.A(G250), .ZN(new_n446));
  OAI21_X1  g0246(.A(new_n446), .B1(new_n293), .B2(G1), .ZN(new_n447));
  NAND3_X1  g0247(.A1(new_n300), .A2(new_n445), .A3(new_n447), .ZN(new_n448));
  INV_X1    g0248(.A(new_n448), .ZN(new_n449));
  NAND3_X1  g0249(.A1(new_n360), .A2(G244), .A3(G1698), .ZN(new_n450));
  NAND2_X1  g0250(.A1(G33), .A2(G116), .ZN(new_n451));
  OAI211_X1 g0251(.A(new_n450), .B(new_n451), .C1(new_n361), .C2(new_n218), .ZN(new_n452));
  AOI21_X1  g0252(.A(new_n449), .B1(new_n452), .B2(new_n289), .ZN(new_n453));
  NOR2_X1   g0253(.A1(new_n453), .A2(new_n305), .ZN(new_n454));
  AOI21_X1  g0254(.A(new_n454), .B1(G190), .B2(new_n453), .ZN(new_n455));
  NAND3_X1  g0255(.A1(new_n360), .A2(new_n213), .A3(G68), .ZN(new_n456));
  INV_X1    g0256(.A(KEYINPUT79), .ZN(new_n457));
  NOR3_X1   g0257(.A1(G87), .A2(G97), .A3(G107), .ZN(new_n458));
  AOI21_X1  g0258(.A(G20), .B1(G33), .B2(G97), .ZN(new_n459));
  OAI21_X1  g0259(.A(KEYINPUT19), .B1(new_n458), .B2(new_n459), .ZN(new_n460));
  INV_X1    g0260(.A(KEYINPUT19), .ZN(new_n461));
  NAND3_X1  g0261(.A1(new_n348), .A2(new_n461), .A3(G97), .ZN(new_n462));
  AOI22_X1  g0262(.A1(new_n456), .A2(new_n457), .B1(new_n460), .B2(new_n462), .ZN(new_n463));
  NOR2_X1   g0263(.A1(new_n315), .A2(G20), .ZN(new_n464));
  NAND3_X1  g0264(.A1(new_n464), .A2(KEYINPUT79), .A3(G68), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n463), .A2(new_n465), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n466), .A2(new_n266), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n419), .A2(new_n403), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n277), .A2(G33), .ZN(new_n469));
  NAND4_X1  g0269(.A1(new_n314), .A2(G87), .A3(new_n278), .A4(new_n469), .ZN(new_n470));
  NAND3_X1  g0270(.A1(new_n467), .A2(new_n468), .A3(new_n470), .ZN(new_n471));
  INV_X1    g0271(.A(new_n471), .ZN(new_n472));
  AOI22_X1  g0272(.A1(new_n466), .A2(new_n266), .B1(new_n403), .B2(new_n419), .ZN(new_n473));
  NAND3_X1  g0273(.A1(new_n314), .A2(new_n278), .A3(new_n469), .ZN(new_n474));
  OAI21_X1  g0274(.A(new_n473), .B1(new_n419), .B2(new_n474), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n453), .A2(G179), .ZN(new_n476));
  OAI21_X1  g0276(.A(new_n476), .B1(new_n376), .B2(new_n453), .ZN(new_n477));
  AOI22_X1  g0277(.A1(new_n455), .A2(new_n472), .B1(new_n475), .B2(new_n477), .ZN(new_n478));
  NOR2_X1   g0278(.A1(new_n451), .A2(G20), .ZN(new_n479));
  INV_X1    g0279(.A(KEYINPUT23), .ZN(new_n480));
  OAI21_X1  g0280(.A(new_n480), .B1(new_n213), .B2(G107), .ZN(new_n481));
  INV_X1    g0281(.A(G107), .ZN(new_n482));
  NAND3_X1  g0282(.A1(new_n482), .A2(KEYINPUT23), .A3(G20), .ZN(new_n483));
  AOI21_X1  g0283(.A(new_n479), .B1(new_n481), .B2(new_n483), .ZN(new_n484));
  INV_X1    g0284(.A(KEYINPUT22), .ZN(new_n485));
  AOI21_X1  g0285(.A(new_n485), .B1(new_n464), .B2(G87), .ZN(new_n486));
  NAND3_X1  g0286(.A1(new_n360), .A2(new_n213), .A3(G87), .ZN(new_n487));
  NOR2_X1   g0287(.A1(new_n487), .A2(KEYINPUT22), .ZN(new_n488));
  OAI21_X1  g0288(.A(new_n484), .B1(new_n486), .B2(new_n488), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n489), .A2(KEYINPUT24), .ZN(new_n490));
  INV_X1    g0290(.A(KEYINPUT24), .ZN(new_n491));
  OAI211_X1 g0291(.A(new_n491), .B(new_n484), .C1(new_n486), .C2(new_n488), .ZN(new_n492));
  AOI21_X1  g0292(.A(new_n314), .B1(new_n490), .B2(new_n492), .ZN(new_n493));
  INV_X1    g0293(.A(new_n493), .ZN(new_n494));
  INV_X1    g0294(.A(KEYINPUT5), .ZN(new_n495));
  OAI211_X1 g0295(.A(new_n277), .B(G45), .C1(new_n495), .C2(G41), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n292), .A2(new_n294), .ZN(new_n497));
  AOI21_X1  g0297(.A(new_n496), .B1(new_n497), .B2(new_n495), .ZN(new_n498));
  NOR2_X1   g0298(.A1(new_n289), .A2(new_n296), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  AOI21_X1  g0300(.A(KEYINPUT5), .B1(new_n292), .B2(new_n294), .ZN(new_n501));
  OAI21_X1  g0301(.A(new_n300), .B1(new_n501), .B2(new_n496), .ZN(new_n502));
  INV_X1    g0302(.A(G264), .ZN(new_n503));
  OAI21_X1  g0303(.A(new_n500), .B1(new_n502), .B2(new_n503), .ZN(new_n504));
  INV_X1    g0304(.A(new_n504), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n360), .A2(G257), .ZN(new_n506));
  INV_X1    g0306(.A(G294), .ZN(new_n507));
  OAI22_X1  g0307(.A1(new_n506), .A2(new_n356), .B1(new_n254), .B2(new_n507), .ZN(new_n508));
  INV_X1    g0308(.A(KEYINPUT80), .ZN(new_n509));
  OAI21_X1  g0309(.A(new_n509), .B1(new_n361), .B2(new_n446), .ZN(new_n510));
  NOR2_X1   g0310(.A1(new_n315), .A2(G1698), .ZN(new_n511));
  NAND3_X1  g0311(.A1(new_n511), .A2(KEYINPUT80), .A3(G250), .ZN(new_n512));
  AOI21_X1  g0312(.A(new_n508), .B1(new_n510), .B2(new_n512), .ZN(new_n513));
  OAI211_X1 g0313(.A(new_n505), .B(G190), .C1(new_n513), .C2(new_n300), .ZN(new_n514));
  OAI21_X1  g0314(.A(new_n505), .B1(new_n513), .B2(new_n300), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n515), .A2(G200), .ZN(new_n516));
  NAND3_X1  g0316(.A1(new_n403), .A2(KEYINPUT25), .A3(new_n482), .ZN(new_n517));
  INV_X1    g0317(.A(new_n517), .ZN(new_n518));
  AOI21_X1  g0318(.A(KEYINPUT25), .B1(new_n403), .B2(new_n482), .ZN(new_n519));
  OAI22_X1  g0319(.A1(new_n518), .A2(new_n519), .B1(new_n474), .B2(new_n482), .ZN(new_n520));
  INV_X1    g0320(.A(new_n520), .ZN(new_n521));
  NAND4_X1  g0321(.A1(new_n494), .A2(new_n514), .A3(new_n516), .A4(new_n521), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n510), .A2(new_n512), .ZN(new_n523));
  INV_X1    g0323(.A(new_n508), .ZN(new_n524));
  AOI21_X1  g0324(.A(new_n300), .B1(new_n523), .B2(new_n524), .ZN(new_n525));
  OAI21_X1  g0325(.A(new_n376), .B1(new_n525), .B2(new_n504), .ZN(new_n526));
  OAI211_X1 g0326(.A(new_n505), .B(new_n338), .C1(new_n513), .C2(new_n300), .ZN(new_n527));
  OAI211_X1 g0327(.A(new_n526), .B(new_n527), .C1(new_n493), .C2(new_n520), .ZN(new_n528));
  NAND3_X1  g0328(.A1(new_n478), .A2(new_n522), .A3(new_n528), .ZN(new_n529));
  AOI21_X1  g0329(.A(G20), .B1(new_n254), .B2(G97), .ZN(new_n530));
  NAND2_X1  g0330(.A1(G33), .A2(G283), .ZN(new_n531));
  INV_X1    g0331(.A(KEYINPUT78), .ZN(new_n532));
  NOR2_X1   g0332(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  AOI21_X1  g0333(.A(KEYINPUT78), .B1(G33), .B2(G283), .ZN(new_n534));
  OAI21_X1  g0334(.A(new_n530), .B1(new_n533), .B2(new_n534), .ZN(new_n535));
  INV_X1    g0335(.A(G116), .ZN(new_n536));
  AOI22_X1  g0336(.A1(new_n265), .A2(new_n212), .B1(G20), .B2(new_n536), .ZN(new_n537));
  AND3_X1   g0337(.A1(new_n535), .A2(KEYINPUT20), .A3(new_n537), .ZN(new_n538));
  AOI21_X1  g0338(.A(KEYINPUT20), .B1(new_n535), .B2(new_n537), .ZN(new_n539));
  NOR2_X1   g0339(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n403), .A2(new_n536), .ZN(new_n541));
  OAI21_X1  g0341(.A(new_n541), .B1(new_n474), .B2(new_n536), .ZN(new_n542));
  NOR2_X1   g0342(.A1(new_n540), .A2(new_n542), .ZN(new_n543));
  NAND3_X1  g0343(.A1(new_n360), .A2(G257), .A3(new_n356), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n315), .A2(G303), .ZN(new_n545));
  OAI211_X1 g0345(.A(new_n544), .B(new_n545), .C1(new_n412), .C2(new_n503), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n546), .A2(new_n289), .ZN(new_n547));
  INV_X1    g0347(.A(new_n502), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n548), .A2(G270), .ZN(new_n549));
  NAND3_X1  g0349(.A1(new_n547), .A2(new_n549), .A3(new_n500), .ZN(new_n550));
  NOR3_X1   g0350(.A1(new_n543), .A2(new_n550), .A3(new_n338), .ZN(new_n551));
  OAI221_X1 g0351(.A(new_n541), .B1(new_n536), .B2(new_n474), .C1(new_n538), .C2(new_n539), .ZN(new_n552));
  NAND3_X1  g0352(.A1(new_n550), .A2(new_n552), .A3(G169), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n553), .A2(KEYINPUT21), .ZN(new_n554));
  INV_X1    g0354(.A(KEYINPUT21), .ZN(new_n555));
  NAND4_X1  g0355(.A1(new_n550), .A2(new_n552), .A3(new_n555), .A4(G169), .ZN(new_n556));
  AOI21_X1  g0356(.A(new_n551), .B1(new_n554), .B2(new_n556), .ZN(new_n557));
  AOI21_X1  g0357(.A(new_n552), .B1(new_n550), .B2(G200), .ZN(new_n558));
  OAI21_X1  g0358(.A(new_n558), .B1(new_n291), .B2(new_n550), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n557), .A2(new_n559), .ZN(new_n560));
  INV_X1    g0360(.A(KEYINPUT4), .ZN(new_n561));
  OAI21_X1  g0361(.A(new_n561), .B1(new_n361), .B2(new_n219), .ZN(new_n562));
  NAND3_X1  g0362(.A1(new_n511), .A2(KEYINPUT4), .A3(G244), .ZN(new_n563));
  OR2_X1    g0363(.A1(new_n533), .A2(new_n534), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n357), .A2(G250), .ZN(new_n565));
  NAND4_X1  g0365(.A1(new_n562), .A2(new_n563), .A3(new_n564), .A4(new_n565), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n566), .A2(new_n289), .ZN(new_n567));
  INV_X1    g0367(.A(G257), .ZN(new_n568));
  OAI21_X1  g0368(.A(new_n500), .B1(new_n568), .B2(new_n502), .ZN(new_n569));
  INV_X1    g0369(.A(new_n569), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n567), .A2(new_n570), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n571), .A2(new_n376), .ZN(new_n572));
  NAND3_X1  g0372(.A1(new_n482), .A2(KEYINPUT6), .A3(G97), .ZN(new_n573));
  OR2_X1    g0373(.A1(new_n573), .A2(KEYINPUT77), .ZN(new_n574));
  INV_X1    g0374(.A(KEYINPUT6), .ZN(new_n575));
  INV_X1    g0375(.A(G97), .ZN(new_n576));
  NOR2_X1   g0376(.A1(new_n576), .A2(new_n482), .ZN(new_n577));
  NOR2_X1   g0377(.A1(G97), .A2(G107), .ZN(new_n578));
  OAI21_X1  g0378(.A(new_n575), .B1(new_n577), .B2(new_n578), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n573), .A2(KEYINPUT77), .ZN(new_n580));
  NAND3_X1  g0380(.A1(new_n574), .A2(new_n579), .A3(new_n580), .ZN(new_n581));
  AOI22_X1  g0381(.A1(new_n581), .A2(G20), .B1(G77), .B2(new_n249), .ZN(new_n582));
  OAI21_X1  g0382(.A(G107), .B1(new_n316), .B2(new_n317), .ZN(new_n583));
  AOI21_X1  g0383(.A(new_n314), .B1(new_n582), .B2(new_n583), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n403), .A2(new_n576), .ZN(new_n585));
  OAI21_X1  g0385(.A(new_n585), .B1(new_n474), .B2(new_n576), .ZN(new_n586));
  OR2_X1    g0386(.A1(new_n584), .A2(new_n586), .ZN(new_n587));
  AOI21_X1  g0387(.A(new_n569), .B1(new_n566), .B2(new_n289), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n588), .A2(new_n338), .ZN(new_n589));
  NAND3_X1  g0389(.A1(new_n572), .A2(new_n587), .A3(new_n589), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n588), .A2(G190), .ZN(new_n591));
  NOR2_X1   g0391(.A1(new_n584), .A2(new_n586), .ZN(new_n592));
  OAI211_X1 g0392(.A(new_n591), .B(new_n592), .C1(new_n305), .C2(new_n588), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n590), .A2(new_n593), .ZN(new_n594));
  NOR3_X1   g0394(.A1(new_n529), .A2(new_n560), .A3(new_n594), .ZN(new_n595));
  AND2_X1   g0395(.A1(new_n444), .A2(new_n595), .ZN(G372));
  INV_X1    g0396(.A(KEYINPUT81), .ZN(new_n597));
  NOR2_X1   g0397(.A1(new_n471), .A2(new_n597), .ZN(new_n598));
  AOI21_X1  g0398(.A(KEYINPUT81), .B1(new_n473), .B2(new_n470), .ZN(new_n599));
  OAI21_X1  g0399(.A(new_n455), .B1(new_n598), .B2(new_n599), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n475), .A2(new_n477), .ZN(new_n601));
  AND3_X1   g0401(.A1(new_n522), .A2(new_n600), .A3(new_n601), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n557), .A2(new_n528), .ZN(new_n603));
  NAND4_X1  g0403(.A1(new_n602), .A2(new_n590), .A3(new_n593), .A4(new_n603), .ZN(new_n604));
  INV_X1    g0404(.A(new_n601), .ZN(new_n605));
  NAND4_X1  g0405(.A1(new_n478), .A2(new_n589), .A3(new_n587), .A4(new_n572), .ZN(new_n606));
  AOI21_X1  g0406(.A(new_n605), .B1(new_n606), .B2(KEYINPUT26), .ZN(new_n607));
  INV_X1    g0407(.A(new_n589), .ZN(new_n608));
  OAI22_X1  g0408(.A1(new_n588), .A2(G169), .B1(new_n584), .B2(new_n586), .ZN(new_n609));
  OAI21_X1  g0409(.A(KEYINPUT82), .B1(new_n608), .B2(new_n609), .ZN(new_n610));
  INV_X1    g0410(.A(KEYINPUT82), .ZN(new_n611));
  NAND4_X1  g0411(.A1(new_n572), .A2(new_n587), .A3(new_n611), .A4(new_n589), .ZN(new_n612));
  AND2_X1   g0412(.A1(new_n610), .A2(new_n612), .ZN(new_n613));
  AND2_X1   g0413(.A1(new_n600), .A2(new_n601), .ZN(new_n614));
  INV_X1    g0414(.A(KEYINPUT26), .ZN(new_n615));
  NAND3_X1  g0415(.A1(new_n613), .A2(new_n614), .A3(new_n615), .ZN(new_n616));
  NAND3_X1  g0416(.A1(new_n604), .A2(new_n607), .A3(new_n616), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n444), .A2(new_n617), .ZN(new_n618));
  XOR2_X1   g0418(.A(new_n618), .B(KEYINPUT83), .Z(new_n619));
  INV_X1    g0419(.A(new_n378), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n427), .A2(KEYINPUT84), .ZN(new_n621));
  INV_X1    g0421(.A(KEYINPUT84), .ZN(new_n622));
  NAND4_X1  g0422(.A1(new_n417), .A2(new_n622), .A3(new_n418), .A4(new_n426), .ZN(new_n623));
  NAND3_X1  g0423(.A1(new_n621), .A2(new_n440), .A3(new_n623), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n408), .A2(new_n624), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n625), .A2(new_n333), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n626), .A2(new_n342), .ZN(new_n627));
  AND2_X1   g0427(.A1(new_n373), .A2(new_n375), .ZN(new_n628));
  AOI21_X1  g0428(.A(new_n620), .B1(new_n627), .B2(new_n628), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n619), .A2(new_n629), .ZN(G369));
  INV_X1    g0430(.A(new_n557), .ZN(new_n631));
  NAND3_X1  g0431(.A1(new_n277), .A2(new_n213), .A3(G13), .ZN(new_n632));
  OR2_X1    g0432(.A1(new_n632), .A2(KEYINPUT27), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n632), .A2(KEYINPUT27), .ZN(new_n634));
  NAND3_X1  g0434(.A1(new_n633), .A2(G213), .A3(new_n634), .ZN(new_n635));
  INV_X1    g0435(.A(G343), .ZN(new_n636));
  NOR2_X1   g0436(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  INV_X1    g0437(.A(new_n637), .ZN(new_n638));
  NOR2_X1   g0438(.A1(new_n543), .A2(new_n638), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n631), .A2(new_n639), .ZN(new_n640));
  OAI21_X1  g0440(.A(new_n640), .B1(new_n560), .B2(new_n639), .ZN(new_n641));
  AND2_X1   g0441(.A1(new_n641), .A2(G330), .ZN(new_n642));
  NOR2_X1   g0442(.A1(new_n528), .A2(new_n637), .ZN(new_n643));
  OAI21_X1  g0443(.A(new_n637), .B1(new_n493), .B2(new_n520), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n522), .A2(new_n644), .ZN(new_n645));
  AOI21_X1  g0445(.A(new_n643), .B1(new_n645), .B2(new_n528), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n642), .A2(new_n646), .ZN(new_n647));
  NOR2_X1   g0447(.A1(new_n557), .A2(new_n637), .ZN(new_n648));
  AND2_X1   g0448(.A1(new_n646), .A2(new_n648), .ZN(new_n649));
  NOR2_X1   g0449(.A1(new_n649), .A2(new_n643), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n647), .A2(new_n650), .ZN(G399));
  NAND2_X1  g0451(.A1(new_n458), .A2(new_n536), .ZN(new_n652));
  XNOR2_X1  g0452(.A(new_n652), .B(KEYINPUT85), .ZN(new_n653));
  INV_X1    g0453(.A(new_n653), .ZN(new_n654));
  INV_X1    g0454(.A(new_n209), .ZN(new_n655));
  NOR2_X1   g0455(.A1(new_n655), .A2(new_n497), .ZN(new_n656));
  INV_X1    g0456(.A(new_n656), .ZN(new_n657));
  NAND3_X1  g0457(.A1(new_n654), .A2(G1), .A3(new_n657), .ZN(new_n658));
  OAI21_X1  g0458(.A(new_n658), .B1(new_n216), .B2(new_n657), .ZN(new_n659));
  XNOR2_X1  g0459(.A(new_n659), .B(KEYINPUT28), .ZN(new_n660));
  XNOR2_X1  g0460(.A(new_n603), .B(KEYINPUT88), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n594), .A2(KEYINPUT89), .ZN(new_n662));
  INV_X1    g0462(.A(KEYINPUT89), .ZN(new_n663));
  NAND3_X1  g0463(.A1(new_n590), .A2(new_n593), .A3(new_n663), .ZN(new_n664));
  NAND3_X1  g0464(.A1(new_n602), .A2(new_n662), .A3(new_n664), .ZN(new_n665));
  OAI21_X1  g0465(.A(new_n601), .B1(new_n661), .B2(new_n665), .ZN(new_n666));
  NAND4_X1  g0466(.A1(new_n613), .A2(new_n614), .A3(KEYINPUT87), .A4(KEYINPUT26), .ZN(new_n667));
  INV_X1    g0467(.A(KEYINPUT87), .ZN(new_n668));
  NAND4_X1  g0468(.A1(new_n610), .A2(new_n600), .A3(new_n612), .A4(new_n601), .ZN(new_n669));
  OAI21_X1  g0469(.A(new_n668), .B1(new_n669), .B2(new_n615), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n606), .A2(new_n615), .ZN(new_n671));
  AND3_X1   g0471(.A1(new_n667), .A2(new_n670), .A3(new_n671), .ZN(new_n672));
  OAI211_X1 g0472(.A(KEYINPUT29), .B(new_n638), .C1(new_n666), .C2(new_n672), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n617), .A2(new_n638), .ZN(new_n674));
  INV_X1    g0474(.A(KEYINPUT29), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  AND2_X1   g0476(.A1(new_n673), .A2(new_n676), .ZN(new_n677));
  NOR4_X1   g0477(.A1(new_n529), .A2(new_n560), .A3(new_n594), .A4(new_n637), .ZN(new_n678));
  INV_X1    g0478(.A(new_n678), .ZN(new_n679));
  INV_X1    g0479(.A(KEYINPUT86), .ZN(new_n680));
  AOI22_X1  g0480(.A1(new_n289), .A2(new_n546), .B1(new_n548), .B2(G270), .ZN(new_n681));
  OAI211_X1 g0481(.A(new_n681), .B(new_n505), .C1(new_n300), .C2(new_n513), .ZN(new_n682));
  INV_X1    g0482(.A(new_n682), .ZN(new_n683));
  AND2_X1   g0483(.A1(new_n453), .A2(G179), .ZN(new_n684));
  NAND4_X1  g0484(.A1(new_n683), .A2(KEYINPUT30), .A3(new_n588), .A4(new_n684), .ZN(new_n685));
  INV_X1    g0485(.A(KEYINPUT30), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n684), .A2(new_n588), .ZN(new_n687));
  OAI21_X1  g0487(.A(new_n686), .B1(new_n687), .B2(new_n682), .ZN(new_n688));
  NOR2_X1   g0488(.A1(new_n453), .A2(G179), .ZN(new_n689));
  NAND4_X1  g0489(.A1(new_n571), .A2(new_n515), .A3(new_n550), .A4(new_n689), .ZN(new_n690));
  NAND3_X1  g0490(.A1(new_n685), .A2(new_n688), .A3(new_n690), .ZN(new_n691));
  AND3_X1   g0491(.A1(new_n691), .A2(KEYINPUT31), .A3(new_n637), .ZN(new_n692));
  AOI21_X1  g0492(.A(KEYINPUT31), .B1(new_n691), .B2(new_n637), .ZN(new_n693));
  OAI21_X1  g0493(.A(new_n680), .B1(new_n692), .B2(new_n693), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n691), .A2(new_n637), .ZN(new_n695));
  INV_X1    g0495(.A(KEYINPUT31), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  NAND3_X1  g0497(.A1(new_n691), .A2(KEYINPUT31), .A3(new_n637), .ZN(new_n698));
  NAND3_X1  g0498(.A1(new_n697), .A2(KEYINPUT86), .A3(new_n698), .ZN(new_n699));
  NAND3_X1  g0499(.A1(new_n679), .A2(new_n694), .A3(new_n699), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n700), .A2(G330), .ZN(new_n701));
  INV_X1    g0501(.A(new_n701), .ZN(new_n702));
  NOR2_X1   g0502(.A1(new_n677), .A2(new_n702), .ZN(new_n703));
  OAI21_X1  g0503(.A(new_n660), .B1(new_n703), .B2(G1), .ZN(G364));
  AND2_X1   g0504(.A1(new_n213), .A2(G13), .ZN(new_n705));
  AOI21_X1  g0505(.A(new_n277), .B1(new_n705), .B2(G45), .ZN(new_n706));
  INV_X1    g0506(.A(new_n706), .ZN(new_n707));
  OR3_X1    g0507(.A1(new_n707), .A2(new_n656), .A3(KEYINPUT90), .ZN(new_n708));
  OAI21_X1  g0508(.A(KEYINPUT90), .B1(new_n707), .B2(new_n656), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  INV_X1    g0510(.A(new_n710), .ZN(new_n711));
  NOR2_X1   g0511(.A1(new_n642), .A2(new_n711), .ZN(new_n712));
  OAI21_X1  g0512(.A(new_n712), .B1(G330), .B2(new_n641), .ZN(new_n713));
  NAND3_X1  g0513(.A1(new_n360), .A2(G355), .A3(new_n209), .ZN(new_n714));
  OAI21_X1  g0514(.A(new_n714), .B1(G116), .B2(new_n209), .ZN(new_n715));
  NOR2_X1   g0515(.A1(new_n655), .A2(new_n360), .ZN(new_n716));
  XOR2_X1   g0516(.A(new_n716), .B(KEYINPUT91), .Z(new_n717));
  INV_X1    g0517(.A(new_n717), .ZN(new_n718));
  INV_X1    g0518(.A(new_n216), .ZN(new_n719));
  AOI21_X1  g0519(.A(new_n718), .B1(new_n293), .B2(new_n719), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n244), .A2(G45), .ZN(new_n721));
  AOI21_X1  g0521(.A(new_n715), .B1(new_n720), .B2(new_n721), .ZN(new_n722));
  NOR2_X1   g0522(.A1(G13), .A2(G33), .ZN(new_n723));
  INV_X1    g0523(.A(new_n723), .ZN(new_n724));
  NOR2_X1   g0524(.A1(new_n724), .A2(G20), .ZN(new_n725));
  AOI21_X1  g0525(.A(new_n212), .B1(G20), .B2(new_n376), .ZN(new_n726));
  NOR2_X1   g0526(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  INV_X1    g0527(.A(new_n727), .ZN(new_n728));
  OAI21_X1  g0528(.A(new_n711), .B1(new_n722), .B2(new_n728), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n291), .A2(G20), .ZN(new_n730));
  INV_X1    g0530(.A(KEYINPUT92), .ZN(new_n731));
  XNOR2_X1  g0531(.A(new_n730), .B(new_n731), .ZN(new_n732));
  NOR3_X1   g0532(.A1(new_n732), .A2(G179), .A3(G200), .ZN(new_n733));
  INV_X1    g0533(.A(new_n733), .ZN(new_n734));
  OR2_X1    g0534(.A1(new_n734), .A2(KEYINPUT94), .ZN(new_n735));
  NAND2_X1  g0535(.A1(new_n734), .A2(KEYINPUT94), .ZN(new_n736));
  NAND2_X1  g0536(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  INV_X1    g0537(.A(new_n737), .ZN(new_n738));
  NAND2_X1  g0538(.A1(new_n738), .A2(G329), .ZN(new_n739));
  NOR3_X1   g0539(.A1(new_n732), .A2(G179), .A3(new_n305), .ZN(new_n740));
  OR2_X1    g0540(.A1(new_n740), .A2(KEYINPUT93), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n740), .A2(KEYINPUT93), .ZN(new_n742));
  NAND2_X1  g0542(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  INV_X1    g0543(.A(new_n743), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n744), .A2(G283), .ZN(new_n745));
  NOR2_X1   g0545(.A1(new_n213), .A2(new_n338), .ZN(new_n746));
  NAND3_X1  g0546(.A1(new_n746), .A2(new_n291), .A3(G200), .ZN(new_n747));
  XOR2_X1   g0547(.A(KEYINPUT33), .B(G317), .Z(new_n748));
  NOR2_X1   g0548(.A1(G190), .A2(G200), .ZN(new_n749));
  NAND2_X1  g0549(.A1(new_n746), .A2(new_n749), .ZN(new_n750));
  INV_X1    g0550(.A(G311), .ZN(new_n751));
  OAI22_X1  g0551(.A1(new_n747), .A2(new_n748), .B1(new_n750), .B2(new_n751), .ZN(new_n752));
  NOR4_X1   g0552(.A1(new_n213), .A2(new_n291), .A3(new_n305), .A4(G179), .ZN(new_n753));
  AOI211_X1 g0553(.A(new_n360), .B(new_n752), .C1(G303), .C2(new_n753), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n746), .A2(G190), .ZN(new_n755));
  NOR2_X1   g0555(.A1(new_n755), .A2(new_n305), .ZN(new_n756));
  NAND2_X1  g0556(.A1(new_n756), .A2(G326), .ZN(new_n757));
  NOR2_X1   g0557(.A1(new_n755), .A2(G200), .ZN(new_n758));
  INV_X1    g0558(.A(new_n758), .ZN(new_n759));
  INV_X1    g0559(.A(G322), .ZN(new_n760));
  OAI21_X1  g0560(.A(new_n757), .B1(new_n759), .B2(new_n760), .ZN(new_n761));
  NOR2_X1   g0561(.A1(G179), .A2(G200), .ZN(new_n762));
  AOI21_X1  g0562(.A(new_n213), .B1(new_n762), .B2(G190), .ZN(new_n763));
  INV_X1    g0563(.A(new_n763), .ZN(new_n764));
  AOI21_X1  g0564(.A(new_n761), .B1(G294), .B2(new_n764), .ZN(new_n765));
  NAND4_X1  g0565(.A1(new_n739), .A2(new_n745), .A3(new_n754), .A4(new_n765), .ZN(new_n766));
  NAND2_X1  g0566(.A1(new_n744), .A2(G107), .ZN(new_n767));
  NAND2_X1  g0567(.A1(new_n733), .A2(G159), .ZN(new_n768));
  XOR2_X1   g0568(.A(new_n768), .B(KEYINPUT32), .Z(new_n769));
  AOI22_X1  g0569(.A1(G50), .A2(new_n756), .B1(new_n758), .B2(G58), .ZN(new_n770));
  OAI21_X1  g0570(.A(new_n770), .B1(new_n576), .B2(new_n763), .ZN(new_n771));
  AND2_X1   g0571(.A1(new_n753), .A2(G87), .ZN(new_n772));
  OAI22_X1  g0572(.A1(new_n747), .A2(new_n203), .B1(new_n750), .B2(new_n204), .ZN(new_n773));
  NOR4_X1   g0573(.A1(new_n771), .A2(new_n315), .A3(new_n772), .A4(new_n773), .ZN(new_n774));
  NAND3_X1  g0574(.A1(new_n767), .A2(new_n769), .A3(new_n774), .ZN(new_n775));
  NAND2_X1  g0575(.A1(new_n766), .A2(new_n775), .ZN(new_n776));
  AOI21_X1  g0576(.A(new_n729), .B1(new_n726), .B2(new_n776), .ZN(new_n777));
  INV_X1    g0577(.A(new_n725), .ZN(new_n778));
  OAI21_X1  g0578(.A(new_n777), .B1(new_n641), .B2(new_n778), .ZN(new_n779));
  AND2_X1   g0579(.A1(new_n713), .A2(new_n779), .ZN(new_n780));
  INV_X1    g0580(.A(new_n780), .ZN(G396));
  NAND2_X1  g0581(.A1(new_n426), .A2(new_n637), .ZN(new_n782));
  NAND3_X1  g0582(.A1(new_n431), .A2(new_n427), .A3(new_n782), .ZN(new_n783));
  INV_X1    g0583(.A(KEYINPUT99), .ZN(new_n784));
  NAND2_X1  g0584(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  NAND4_X1  g0585(.A1(new_n431), .A2(new_n427), .A3(KEYINPUT99), .A4(new_n782), .ZN(new_n786));
  NAND2_X1  g0586(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  INV_X1    g0587(.A(new_n782), .ZN(new_n788));
  NAND3_X1  g0588(.A1(new_n621), .A2(new_n623), .A3(new_n788), .ZN(new_n789));
  NAND2_X1  g0589(.A1(new_n789), .A2(KEYINPUT100), .ZN(new_n790));
  INV_X1    g0590(.A(KEYINPUT100), .ZN(new_n791));
  NAND4_X1  g0591(.A1(new_n621), .A2(new_n791), .A3(new_n623), .A4(new_n788), .ZN(new_n792));
  NAND3_X1  g0592(.A1(new_n787), .A2(new_n790), .A3(new_n792), .ZN(new_n793));
  XOR2_X1   g0593(.A(new_n674), .B(new_n793), .Z(new_n794));
  AOI21_X1  g0594(.A(new_n711), .B1(new_n794), .B2(new_n701), .ZN(new_n795));
  OAI21_X1  g0595(.A(new_n795), .B1(new_n701), .B2(new_n794), .ZN(new_n796));
  NOR2_X1   g0596(.A1(new_n726), .A2(new_n723), .ZN(new_n797));
  INV_X1    g0597(.A(new_n797), .ZN(new_n798));
  OAI21_X1  g0598(.A(new_n711), .B1(G77), .B2(new_n798), .ZN(new_n799));
  NAND2_X1  g0599(.A1(new_n738), .A2(G311), .ZN(new_n800));
  INV_X1    g0600(.A(G283), .ZN(new_n801));
  OAI22_X1  g0601(.A1(new_n747), .A2(new_n801), .B1(new_n750), .B2(new_n536), .ZN(new_n802));
  INV_X1    g0602(.A(new_n756), .ZN(new_n803));
  INV_X1    g0603(.A(G303), .ZN(new_n804));
  OAI22_X1  g0604(.A1(new_n507), .A2(new_n759), .B1(new_n803), .B2(new_n804), .ZN(new_n805));
  AOI211_X1 g0605(.A(new_n802), .B(new_n805), .C1(G97), .C2(new_n764), .ZN(new_n806));
  NAND2_X1  g0606(.A1(new_n744), .A2(G87), .ZN(new_n807));
  AOI21_X1  g0607(.A(new_n360), .B1(new_n753), .B2(G107), .ZN(new_n808));
  XNOR2_X1  g0608(.A(new_n808), .B(KEYINPUT95), .ZN(new_n809));
  NAND4_X1  g0609(.A1(new_n800), .A2(new_n806), .A3(new_n807), .A4(new_n809), .ZN(new_n810));
  NAND2_X1  g0610(.A1(new_n744), .A2(G68), .ZN(new_n811));
  INV_X1    g0611(.A(new_n753), .ZN(new_n812));
  OAI21_X1  g0612(.A(new_n811), .B1(new_n201), .B2(new_n812), .ZN(new_n813));
  XNOR2_X1  g0613(.A(new_n813), .B(KEYINPUT97), .ZN(new_n814));
  INV_X1    g0614(.A(new_n747), .ZN(new_n815));
  INV_X1    g0615(.A(new_n750), .ZN(new_n816));
  AOI22_X1  g0616(.A1(new_n815), .A2(G150), .B1(new_n816), .B2(G159), .ZN(new_n817));
  INV_X1    g0617(.A(G137), .ZN(new_n818));
  XNOR2_X1  g0618(.A(KEYINPUT96), .B(G143), .ZN(new_n819));
  OAI221_X1 g0619(.A(new_n817), .B1(new_n803), .B2(new_n818), .C1(new_n759), .C2(new_n819), .ZN(new_n820));
  XNOR2_X1  g0620(.A(new_n820), .B(KEYINPUT34), .ZN(new_n821));
  AOI21_X1  g0621(.A(new_n315), .B1(new_n764), .B2(G58), .ZN(new_n822));
  INV_X1    g0622(.A(G132), .ZN(new_n823));
  OAI211_X1 g0623(.A(new_n821), .B(new_n822), .C1(new_n823), .C2(new_n737), .ZN(new_n824));
  OAI21_X1  g0624(.A(new_n810), .B1(new_n814), .B2(new_n824), .ZN(new_n825));
  AOI21_X1  g0625(.A(new_n799), .B1(new_n825), .B2(new_n726), .ZN(new_n826));
  XOR2_X1   g0626(.A(new_n826), .B(KEYINPUT98), .Z(new_n827));
  OAI21_X1  g0627(.A(new_n827), .B1(new_n724), .B2(new_n793), .ZN(new_n828));
  NAND2_X1  g0628(.A1(new_n796), .A2(new_n828), .ZN(G384));
  NAND2_X1  g0629(.A1(new_n407), .A2(new_n637), .ZN(new_n830));
  NAND3_X1  g0630(.A1(new_n408), .A2(new_n440), .A3(new_n830), .ZN(new_n831));
  INV_X1    g0631(.A(KEYINPUT102), .ZN(new_n832));
  AND3_X1   g0632(.A1(new_n390), .A2(new_n392), .A3(new_n394), .ZN(new_n833));
  AOI21_X1  g0633(.A(KEYINPUT73), .B1(new_n433), .B2(new_n434), .ZN(new_n834));
  NOR2_X1   g0634(.A1(new_n440), .A2(new_n441), .ZN(new_n835));
  OAI21_X1  g0635(.A(new_n833), .B1(new_n834), .B2(new_n835), .ZN(new_n836));
  INV_X1    g0636(.A(new_n830), .ZN(new_n837));
  AOI21_X1  g0637(.A(new_n832), .B1(new_n836), .B2(new_n837), .ZN(new_n838));
  AOI21_X1  g0638(.A(new_n395), .B1(new_n435), .B2(new_n442), .ZN(new_n839));
  NOR3_X1   g0639(.A1(new_n839), .A2(KEYINPUT102), .A3(new_n830), .ZN(new_n840));
  OAI21_X1  g0640(.A(new_n831), .B1(new_n838), .B2(new_n840), .ZN(new_n841));
  NAND3_X1  g0641(.A1(new_n679), .A2(new_n697), .A3(new_n698), .ZN(new_n842));
  NAND3_X1  g0642(.A1(new_n841), .A2(new_n842), .A3(new_n793), .ZN(new_n843));
  AOI21_X1  g0643(.A(new_n251), .B1(new_n325), .B2(new_n326), .ZN(new_n844));
  OAI21_X1  g0644(.A(new_n266), .B1(new_n844), .B2(KEYINPUT16), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n845), .A2(KEYINPUT103), .ZN(new_n846));
  INV_X1    g0646(.A(KEYINPUT103), .ZN(new_n847));
  OAI211_X1 g0647(.A(new_n847), .B(new_n266), .C1(new_n844), .C2(KEYINPUT16), .ZN(new_n848));
  NAND3_X1  g0648(.A1(new_n846), .A2(new_n264), .A3(new_n848), .ZN(new_n849));
  AOI21_X1  g0649(.A(new_n635), .B1(new_n849), .B2(new_n281), .ZN(new_n850));
  INV_X1    g0650(.A(new_n635), .ZN(new_n851));
  NOR2_X1   g0651(.A1(new_n339), .A2(new_n851), .ZN(new_n852));
  AOI21_X1  g0652(.A(new_n852), .B1(new_n849), .B2(new_n281), .ZN(new_n853));
  NAND2_X1  g0653(.A1(new_n330), .A2(new_n331), .ZN(new_n854));
  OAI21_X1  g0654(.A(KEYINPUT37), .B1(new_n853), .B2(new_n854), .ZN(new_n855));
  XNOR2_X1  g0655(.A(new_n635), .B(KEYINPUT104), .ZN(new_n856));
  OAI21_X1  g0656(.A(new_n334), .B1(new_n339), .B2(new_n856), .ZN(new_n857));
  INV_X1    g0657(.A(KEYINPUT37), .ZN(new_n858));
  NAND4_X1  g0658(.A1(new_n857), .A2(new_n858), .A3(new_n330), .A4(new_n331), .ZN(new_n859));
  AOI22_X1  g0659(.A1(new_n343), .A2(new_n850), .B1(new_n855), .B2(new_n859), .ZN(new_n860));
  OAI21_X1  g0660(.A(KEYINPUT105), .B1(new_n860), .B2(KEYINPUT38), .ZN(new_n861));
  INV_X1    g0661(.A(KEYINPUT105), .ZN(new_n862));
  INV_X1    g0662(.A(KEYINPUT38), .ZN(new_n863));
  AND2_X1   g0663(.A1(new_n855), .A2(new_n859), .ZN(new_n864));
  INV_X1    g0664(.A(new_n850), .ZN(new_n865));
  AOI21_X1  g0665(.A(new_n865), .B1(new_n333), .B2(new_n342), .ZN(new_n866));
  OAI211_X1 g0666(.A(new_n862), .B(new_n863), .C1(new_n864), .C2(new_n866), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n860), .A2(KEYINPUT38), .ZN(new_n868));
  NAND3_X1  g0668(.A1(new_n861), .A2(new_n867), .A3(new_n868), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n869), .A2(KEYINPUT106), .ZN(new_n870));
  INV_X1    g0670(.A(KEYINPUT106), .ZN(new_n871));
  NAND4_X1  g0671(.A1(new_n861), .A2(new_n871), .A3(new_n867), .A4(new_n868), .ZN(new_n872));
  AOI21_X1  g0672(.A(new_n843), .B1(new_n870), .B2(new_n872), .ZN(new_n873));
  OR2_X1    g0673(.A1(new_n873), .A2(KEYINPUT40), .ZN(new_n874));
  NAND3_X1  g0674(.A1(new_n321), .A2(KEYINPUT107), .A3(new_n309), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n857), .A2(new_n875), .ZN(new_n876));
  AOI21_X1  g0676(.A(KEYINPUT107), .B1(new_n321), .B2(new_n309), .ZN(new_n877));
  OAI21_X1  g0677(.A(KEYINPUT37), .B1(new_n876), .B2(new_n877), .ZN(new_n878));
  AND2_X1   g0678(.A1(new_n878), .A2(new_n859), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n334), .A2(new_n856), .ZN(new_n880));
  AOI21_X1  g0680(.A(new_n880), .B1(new_n333), .B2(new_n342), .ZN(new_n881));
  OAI21_X1  g0681(.A(new_n863), .B1(new_n879), .B2(new_n881), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n868), .A2(new_n882), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n883), .A2(KEYINPUT40), .ZN(new_n884));
  OR2_X1    g0684(.A1(new_n884), .A2(new_n843), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n874), .A2(new_n885), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n444), .A2(new_n842), .ZN(new_n887));
  OAI21_X1  g0687(.A(G330), .B1(new_n886), .B2(new_n887), .ZN(new_n888));
  AOI21_X1  g0688(.A(new_n888), .B1(new_n887), .B2(new_n886), .ZN(new_n889));
  OR2_X1    g0689(.A1(new_n342), .A2(new_n856), .ZN(new_n890));
  NOR2_X1   g0690(.A1(new_n883), .A2(KEYINPUT39), .ZN(new_n891));
  AOI21_X1  g0691(.A(new_n891), .B1(KEYINPUT39), .B2(new_n869), .ZN(new_n892));
  NAND3_X1  g0692(.A1(new_n395), .A2(new_n407), .A3(new_n638), .ZN(new_n893));
  OAI21_X1  g0693(.A(new_n890), .B1(new_n892), .B2(new_n893), .ZN(new_n894));
  NAND3_X1  g0694(.A1(new_n617), .A2(new_n638), .A3(new_n793), .ZN(new_n895));
  NOR2_X1   g0695(.A1(new_n427), .A2(new_n637), .ZN(new_n896));
  INV_X1    g0696(.A(new_n896), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n895), .A2(new_n897), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n898), .A2(new_n841), .ZN(new_n899));
  AOI21_X1  g0699(.A(new_n899), .B1(new_n870), .B2(new_n872), .ZN(new_n900));
  NOR2_X1   g0700(.A1(new_n894), .A2(new_n900), .ZN(new_n901));
  NAND3_X1  g0701(.A1(new_n673), .A2(new_n444), .A3(new_n676), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n902), .A2(new_n629), .ZN(new_n903));
  XNOR2_X1  g0703(.A(new_n901), .B(new_n903), .ZN(new_n904));
  OAI22_X1  g0704(.A1(new_n889), .A2(new_n904), .B1(new_n277), .B2(new_n705), .ZN(new_n905));
  AOI21_X1  g0705(.A(new_n905), .B1(new_n904), .B2(new_n889), .ZN(new_n906));
  AND2_X1   g0706(.A1(new_n581), .A2(KEYINPUT35), .ZN(new_n907));
  NOR2_X1   g0707(.A1(new_n581), .A2(KEYINPUT35), .ZN(new_n908));
  NOR4_X1   g0708(.A1(new_n907), .A2(new_n908), .A3(new_n536), .A4(new_n215), .ZN(new_n909));
  XNOR2_X1  g0709(.A(new_n909), .B(KEYINPUT36), .ZN(new_n910));
  NOR3_X1   g0710(.A1(new_n246), .A2(new_n216), .A3(new_n204), .ZN(new_n911));
  INV_X1    g0711(.A(new_n911), .ZN(new_n912));
  OR2_X1    g0712(.A1(new_n912), .A2(KEYINPUT101), .ZN(new_n913));
  AOI22_X1  g0713(.A1(new_n912), .A2(KEYINPUT101), .B1(new_n201), .B2(G68), .ZN(new_n914));
  AOI211_X1 g0714(.A(new_n277), .B(G13), .C1(new_n913), .C2(new_n914), .ZN(new_n915));
  OR3_X1    g0715(.A1(new_n906), .A2(new_n910), .A3(new_n915), .ZN(G367));
  INV_X1    g0716(.A(new_n703), .ZN(new_n917));
  AND2_X1   g0717(.A1(new_n662), .A2(new_n664), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n587), .A2(new_n637), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  NOR2_X1   g0720(.A1(new_n590), .A2(new_n638), .ZN(new_n921));
  INV_X1    g0721(.A(new_n921), .ZN(new_n922));
  OAI211_X1 g0722(.A(new_n920), .B(new_n922), .C1(new_n649), .C2(new_n643), .ZN(new_n923));
  XNOR2_X1  g0723(.A(new_n923), .B(KEYINPUT44), .ZN(new_n924));
  INV_X1    g0724(.A(new_n924), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n920), .A2(new_n922), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n650), .A2(new_n926), .ZN(new_n927));
  INV_X1    g0727(.A(KEYINPUT45), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  NAND3_X1  g0729(.A1(new_n650), .A2(new_n926), .A3(KEYINPUT45), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n647), .A2(KEYINPUT110), .ZN(new_n932));
  OR2_X1    g0732(.A1(new_n647), .A2(KEYINPUT110), .ZN(new_n933));
  NAND4_X1  g0733(.A1(new_n925), .A2(new_n931), .A3(new_n932), .A4(new_n933), .ZN(new_n934));
  AND2_X1   g0734(.A1(new_n929), .A2(new_n930), .ZN(new_n935));
  OAI211_X1 g0735(.A(KEYINPUT110), .B(new_n647), .C1(new_n935), .C2(new_n924), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n934), .A2(new_n936), .ZN(new_n937));
  NOR2_X1   g0737(.A1(new_n646), .A2(new_n648), .ZN(new_n938));
  NOR2_X1   g0738(.A1(new_n649), .A2(new_n938), .ZN(new_n939));
  XNOR2_X1  g0739(.A(new_n939), .B(new_n642), .ZN(new_n940));
  INV_X1    g0740(.A(new_n940), .ZN(new_n941));
  AOI21_X1  g0741(.A(new_n917), .B1(new_n937), .B2(new_n941), .ZN(new_n942));
  XOR2_X1   g0742(.A(new_n656), .B(KEYINPUT41), .Z(new_n943));
  OAI21_X1  g0743(.A(new_n706), .B1(new_n942), .B2(new_n943), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n926), .A2(new_n649), .ZN(new_n945));
  INV_X1    g0745(.A(KEYINPUT42), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n945), .A2(new_n946), .ZN(new_n947));
  NAND3_X1  g0747(.A1(new_n926), .A2(KEYINPUT42), .A3(new_n649), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  OR2_X1    g0749(.A1(new_n920), .A2(new_n528), .ZN(new_n950));
  AND2_X1   g0750(.A1(new_n950), .A2(new_n590), .ZN(new_n951));
  OAI21_X1  g0751(.A(new_n949), .B1(new_n637), .B2(new_n951), .ZN(new_n952));
  NAND3_X1  g0752(.A1(new_n952), .A2(KEYINPUT109), .A3(KEYINPUT43), .ZN(new_n953));
  INV_X1    g0753(.A(KEYINPUT43), .ZN(new_n954));
  AOI21_X1  g0754(.A(new_n637), .B1(new_n950), .B2(new_n590), .ZN(new_n955));
  AOI21_X1  g0755(.A(new_n955), .B1(new_n948), .B2(new_n947), .ZN(new_n956));
  INV_X1    g0756(.A(KEYINPUT109), .ZN(new_n957));
  OAI21_X1  g0757(.A(new_n954), .B1(new_n956), .B2(new_n957), .ZN(new_n958));
  OR2_X1    g0758(.A1(new_n598), .A2(new_n599), .ZN(new_n959));
  NOR2_X1   g0759(.A1(new_n959), .A2(new_n638), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n960), .A2(new_n601), .ZN(new_n961));
  OAI21_X1  g0761(.A(new_n961), .B1(new_n614), .B2(new_n960), .ZN(new_n962));
  XNOR2_X1  g0762(.A(new_n962), .B(KEYINPUT108), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n952), .A2(new_n963), .ZN(new_n964));
  NAND3_X1  g0764(.A1(new_n953), .A2(new_n958), .A3(new_n964), .ZN(new_n965));
  INV_X1    g0765(.A(new_n926), .ZN(new_n966));
  AND2_X1   g0766(.A1(new_n953), .A2(new_n958), .ZN(new_n967));
  INV_X1    g0767(.A(new_n963), .ZN(new_n968));
  OAI221_X1 g0768(.A(new_n965), .B1(new_n647), .B2(new_n966), .C1(new_n967), .C2(new_n968), .ZN(new_n969));
  NOR2_X1   g0769(.A1(new_n966), .A2(new_n647), .ZN(new_n970));
  INV_X1    g0770(.A(new_n965), .ZN(new_n971));
  AOI21_X1  g0771(.A(new_n968), .B1(new_n953), .B2(new_n958), .ZN(new_n972));
  OAI21_X1  g0772(.A(new_n970), .B1(new_n971), .B2(new_n972), .ZN(new_n973));
  NAND3_X1  g0773(.A1(new_n944), .A2(new_n969), .A3(new_n973), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n968), .A2(new_n725), .ZN(new_n975));
  OAI221_X1 g0775(.A(new_n727), .B1(new_n209), .B2(new_n419), .C1(new_n718), .C2(new_n236), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n976), .A2(new_n711), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n744), .A2(G97), .ZN(new_n978));
  OAI221_X1 g0778(.A(new_n315), .B1(new_n750), .B2(new_n801), .C1(new_n507), .C2(new_n747), .ZN(new_n979));
  NOR2_X1   g0779(.A1(new_n803), .A2(new_n751), .ZN(new_n980));
  NOR2_X1   g0780(.A1(new_n812), .A2(new_n536), .ZN(new_n981));
  AOI211_X1 g0781(.A(new_n979), .B(new_n980), .C1(KEYINPUT46), .C2(new_n981), .ZN(new_n982));
  OAI22_X1  g0782(.A1(new_n981), .A2(KEYINPUT46), .B1(new_n804), .B2(new_n759), .ZN(new_n983));
  AOI21_X1  g0783(.A(new_n983), .B1(G107), .B2(new_n764), .ZN(new_n984));
  XNOR2_X1  g0784(.A(KEYINPUT111), .B(G317), .ZN(new_n985));
  OR2_X1    g0785(.A1(new_n734), .A2(new_n985), .ZN(new_n986));
  NAND4_X1  g0786(.A1(new_n978), .A2(new_n982), .A3(new_n984), .A4(new_n986), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n744), .A2(G77), .ZN(new_n988));
  NAND2_X1  g0788(.A1(new_n988), .A2(new_n360), .ZN(new_n989));
  AND2_X1   g0789(.A1(new_n989), .A2(KEYINPUT112), .ZN(new_n990));
  AOI22_X1  g0790(.A1(new_n815), .A2(G159), .B1(new_n816), .B2(G50), .ZN(new_n991));
  OAI21_X1  g0791(.A(new_n991), .B1(new_n202), .B2(new_n812), .ZN(new_n992));
  AOI22_X1  g0792(.A1(new_n758), .A2(G150), .B1(G68), .B2(new_n764), .ZN(new_n993));
  OAI21_X1  g0793(.A(new_n993), .B1(new_n803), .B2(new_n819), .ZN(new_n994));
  AOI211_X1 g0794(.A(new_n992), .B(new_n994), .C1(G137), .C2(new_n733), .ZN(new_n995));
  OAI21_X1  g0795(.A(new_n995), .B1(new_n989), .B2(KEYINPUT112), .ZN(new_n996));
  OAI21_X1  g0796(.A(new_n987), .B1(new_n990), .B2(new_n996), .ZN(new_n997));
  XNOR2_X1  g0797(.A(new_n997), .B(KEYINPUT47), .ZN(new_n998));
  AOI21_X1  g0798(.A(new_n977), .B1(new_n998), .B2(new_n726), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n975), .A2(new_n999), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n974), .A2(new_n1000), .ZN(G387));
  NAND2_X1  g0801(.A1(new_n917), .A2(new_n940), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n703), .A2(new_n941), .ZN(new_n1003));
  NAND3_X1  g0803(.A1(new_n1002), .A2(new_n656), .A3(new_n1003), .ZN(new_n1004));
  NOR2_X1   g0804(.A1(new_n646), .A2(new_n778), .ZN(new_n1005));
  NAND3_X1  g0805(.A1(new_n653), .A2(new_n209), .A3(new_n360), .ZN(new_n1006));
  OAI21_X1  g0806(.A(new_n1006), .B1(G107), .B2(new_n209), .ZN(new_n1007));
  XNOR2_X1  g0807(.A(new_n1007), .B(KEYINPUT113), .ZN(new_n1008));
  NOR2_X1   g0808(.A1(new_n233), .A2(new_n293), .ZN(new_n1009));
  NOR2_X1   g0809(.A1(new_n272), .A2(G50), .ZN(new_n1010));
  XNOR2_X1  g0810(.A(KEYINPUT114), .B(KEYINPUT50), .ZN(new_n1011));
  XNOR2_X1  g0811(.A(new_n1010), .B(new_n1011), .ZN(new_n1012));
  AOI21_X1  g0812(.A(G45), .B1(G68), .B2(G77), .ZN(new_n1013));
  NAND3_X1  g0813(.A1(new_n1012), .A2(new_n654), .A3(new_n1013), .ZN(new_n1014));
  NAND2_X1  g0814(.A1(new_n1014), .A2(new_n717), .ZN(new_n1015));
  NOR2_X1   g0815(.A1(new_n1009), .A2(new_n1015), .ZN(new_n1016));
  OAI21_X1  g0816(.A(new_n727), .B1(new_n1008), .B2(new_n1016), .ZN(new_n1017));
  NAND2_X1  g0817(.A1(new_n1017), .A2(new_n711), .ZN(new_n1018));
  NAND2_X1  g0818(.A1(new_n764), .A2(new_n420), .ZN(new_n1019));
  INV_X1    g0819(.A(G159), .ZN(new_n1020));
  OAI21_X1  g0820(.A(new_n1019), .B1(new_n803), .B2(new_n1020), .ZN(new_n1021));
  OAI221_X1 g0821(.A(new_n360), .B1(new_n203), .B2(new_n750), .C1(new_n759), .C2(new_n201), .ZN(new_n1022));
  AOI211_X1 g0822(.A(new_n1021), .B(new_n1022), .C1(new_n347), .C2(new_n815), .ZN(new_n1023));
  AOI22_X1  g0823(.A1(new_n733), .A2(G150), .B1(G77), .B2(new_n753), .ZN(new_n1024));
  XNOR2_X1  g0824(.A(new_n1024), .B(KEYINPUT115), .ZN(new_n1025));
  NAND3_X1  g0825(.A1(new_n978), .A2(new_n1023), .A3(new_n1025), .ZN(new_n1026));
  AOI22_X1  g0826(.A1(new_n815), .A2(G311), .B1(new_n816), .B2(G303), .ZN(new_n1027));
  OAI221_X1 g0827(.A(new_n1027), .B1(new_n803), .B2(new_n760), .C1(new_n759), .C2(new_n985), .ZN(new_n1028));
  INV_X1    g0828(.A(KEYINPUT48), .ZN(new_n1029));
  OR2_X1    g0829(.A1(new_n1028), .A2(new_n1029), .ZN(new_n1030));
  NAND2_X1  g0830(.A1(new_n1028), .A2(new_n1029), .ZN(new_n1031));
  AOI22_X1  g0831(.A1(new_n753), .A2(G294), .B1(new_n764), .B2(G283), .ZN(new_n1032));
  NAND3_X1  g0832(.A1(new_n1030), .A2(new_n1031), .A3(new_n1032), .ZN(new_n1033));
  XNOR2_X1  g0833(.A(KEYINPUT116), .B(KEYINPUT49), .ZN(new_n1034));
  XNOR2_X1  g0834(.A(new_n1033), .B(new_n1034), .ZN(new_n1035));
  NAND2_X1  g0835(.A1(new_n1035), .A2(KEYINPUT117), .ZN(new_n1036));
  AOI21_X1  g0836(.A(new_n360), .B1(new_n733), .B2(G326), .ZN(new_n1037));
  OAI211_X1 g0837(.A(new_n1036), .B(new_n1037), .C1(new_n536), .C2(new_n743), .ZN(new_n1038));
  NOR2_X1   g0838(.A1(new_n1035), .A2(KEYINPUT117), .ZN(new_n1039));
  OAI21_X1  g0839(.A(new_n1026), .B1(new_n1038), .B2(new_n1039), .ZN(new_n1040));
  AOI211_X1 g0840(.A(new_n1005), .B(new_n1018), .C1(new_n1040), .C2(new_n726), .ZN(new_n1041));
  AOI21_X1  g0841(.A(new_n1041), .B1(new_n941), .B2(new_n707), .ZN(new_n1042));
  NAND2_X1  g0842(.A1(new_n1004), .A2(new_n1042), .ZN(G393));
  AOI21_X1  g0843(.A(new_n706), .B1(new_n934), .B2(new_n936), .ZN(new_n1044));
  INV_X1    g0844(.A(KEYINPUT118), .ZN(new_n1045));
  AOI22_X1  g0845(.A1(G150), .A2(new_n756), .B1(new_n758), .B2(G159), .ZN(new_n1046));
  XOR2_X1   g0846(.A(new_n1046), .B(KEYINPUT51), .Z(new_n1047));
  OR2_X1    g0847(.A1(new_n734), .A2(new_n819), .ZN(new_n1048));
  OAI21_X1  g0848(.A(new_n360), .B1(new_n750), .B2(new_n272), .ZN(new_n1049));
  OAI22_X1  g0849(.A1(new_n812), .A2(new_n203), .B1(new_n201), .B2(new_n747), .ZN(new_n1050));
  AOI211_X1 g0850(.A(new_n1049), .B(new_n1050), .C1(G77), .C2(new_n764), .ZN(new_n1051));
  NAND4_X1  g0851(.A1(new_n807), .A2(new_n1047), .A3(new_n1048), .A4(new_n1051), .ZN(new_n1052));
  OAI22_X1  g0852(.A1(new_n747), .A2(new_n804), .B1(new_n750), .B2(new_n507), .ZN(new_n1053));
  OAI21_X1  g0853(.A(new_n315), .B1(new_n812), .B2(new_n801), .ZN(new_n1054));
  AOI211_X1 g0854(.A(new_n1053), .B(new_n1054), .C1(G116), .C2(new_n764), .ZN(new_n1055));
  OAI211_X1 g0855(.A(new_n767), .B(new_n1055), .C1(new_n760), .C2(new_n734), .ZN(new_n1056));
  AOI22_X1  g0856(.A1(G311), .A2(new_n758), .B1(new_n756), .B2(G317), .ZN(new_n1057));
  XNOR2_X1  g0857(.A(new_n1057), .B(KEYINPUT52), .ZN(new_n1058));
  OAI21_X1  g0858(.A(new_n1052), .B1(new_n1056), .B2(new_n1058), .ZN(new_n1059));
  NAND2_X1  g0859(.A1(new_n1059), .A2(new_n726), .ZN(new_n1060));
  NAND2_X1  g0860(.A1(new_n717), .A2(new_n240), .ZN(new_n1061));
  AOI21_X1  g0861(.A(new_n728), .B1(G97), .B2(new_n655), .ZN(new_n1062));
  AOI21_X1  g0862(.A(new_n710), .B1(new_n1061), .B2(new_n1062), .ZN(new_n1063));
  OAI211_X1 g0863(.A(new_n1060), .B(new_n1063), .C1(new_n926), .C2(new_n778), .ZN(new_n1064));
  INV_X1    g0864(.A(new_n1064), .ZN(new_n1065));
  OR3_X1    g0865(.A1(new_n1044), .A2(new_n1045), .A3(new_n1065), .ZN(new_n1066));
  OAI21_X1  g0866(.A(new_n1045), .B1(new_n1044), .B2(new_n1065), .ZN(new_n1067));
  NAND2_X1  g0867(.A1(new_n1066), .A2(new_n1067), .ZN(new_n1068));
  INV_X1    g0868(.A(new_n1003), .ZN(new_n1069));
  AOI21_X1  g0869(.A(new_n657), .B1(new_n937), .B2(new_n1069), .ZN(new_n1070));
  OAI21_X1  g0870(.A(new_n1070), .B1(new_n1069), .B2(new_n937), .ZN(new_n1071));
  NAND2_X1  g0871(.A1(new_n1068), .A2(new_n1071), .ZN(G390));
  NAND2_X1  g0872(.A1(new_n697), .A2(new_n698), .ZN(new_n1073));
  OAI211_X1 g0873(.A(G330), .B(new_n793), .C1(new_n1073), .C2(new_n678), .ZN(new_n1074));
  INV_X1    g0874(.A(new_n831), .ZN(new_n1075));
  OAI21_X1  g0875(.A(KEYINPUT102), .B1(new_n839), .B2(new_n830), .ZN(new_n1076));
  NAND3_X1  g0876(.A1(new_n836), .A2(new_n832), .A3(new_n837), .ZN(new_n1077));
  AOI21_X1  g0877(.A(new_n1075), .B1(new_n1076), .B2(new_n1077), .ZN(new_n1078));
  NOR2_X1   g0878(.A1(new_n1074), .A2(new_n1078), .ZN(new_n1079));
  NAND2_X1  g0879(.A1(new_n899), .A2(new_n893), .ZN(new_n1080));
  NAND2_X1  g0880(.A1(new_n869), .A2(KEYINPUT39), .ZN(new_n1081));
  INV_X1    g0881(.A(new_n891), .ZN(new_n1082));
  AND3_X1   g0882(.A1(new_n1080), .A2(new_n1081), .A3(new_n1082), .ZN(new_n1083));
  NAND2_X1  g0883(.A1(new_n883), .A2(new_n893), .ZN(new_n1084));
  OAI211_X1 g0884(.A(new_n638), .B(new_n793), .C1(new_n666), .C2(new_n672), .ZN(new_n1085));
  NAND2_X1  g0885(.A1(new_n1085), .A2(new_n897), .ZN(new_n1086));
  AOI21_X1  g0886(.A(new_n1084), .B1(new_n1086), .B2(new_n841), .ZN(new_n1087));
  OAI21_X1  g0887(.A(new_n1079), .B1(new_n1083), .B2(new_n1087), .ZN(new_n1088));
  INV_X1    g0888(.A(new_n1087), .ZN(new_n1089));
  NAND2_X1  g0889(.A1(new_n892), .A2(new_n1080), .ZN(new_n1090));
  NAND4_X1  g0890(.A1(new_n841), .A2(new_n700), .A3(G330), .A4(new_n793), .ZN(new_n1091));
  NAND3_X1  g0891(.A1(new_n1089), .A2(new_n1090), .A3(new_n1091), .ZN(new_n1092));
  NAND2_X1  g0892(.A1(new_n1088), .A2(new_n1092), .ZN(new_n1093));
  NOR2_X1   g0893(.A1(new_n1093), .A2(new_n706), .ZN(new_n1094));
  NAND2_X1  g0894(.A1(new_n892), .A2(new_n723), .ZN(new_n1095));
  OAI21_X1  g0895(.A(new_n711), .B1(new_n347), .B2(new_n798), .ZN(new_n1096));
  AOI22_X1  g0896(.A1(new_n758), .A2(G116), .B1(G77), .B2(new_n764), .ZN(new_n1097));
  OAI21_X1  g0897(.A(new_n1097), .B1(new_n801), .B2(new_n803), .ZN(new_n1098));
  OAI22_X1  g0898(.A1(new_n747), .A2(new_n482), .B1(new_n750), .B2(new_n576), .ZN(new_n1099));
  NOR4_X1   g0899(.A1(new_n1098), .A2(new_n360), .A3(new_n772), .A4(new_n1099), .ZN(new_n1100));
  OAI211_X1 g0900(.A(new_n811), .B(new_n1100), .C1(new_n507), .C2(new_n737), .ZN(new_n1101));
  INV_X1    g0901(.A(KEYINPUT120), .ZN(new_n1102));
  OR2_X1    g0902(.A1(new_n1101), .A2(new_n1102), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n756), .A2(G128), .ZN(new_n1104));
  OAI21_X1  g0904(.A(new_n1104), .B1(new_n759), .B2(new_n823), .ZN(new_n1105));
  NAND2_X1  g0905(.A1(new_n753), .A2(G150), .ZN(new_n1106));
  OAI22_X1  g0906(.A1(new_n1106), .A2(KEYINPUT53), .B1(new_n1020), .B2(new_n763), .ZN(new_n1107));
  AND2_X1   g0907(.A1(new_n1106), .A2(KEYINPUT53), .ZN(new_n1108));
  XNOR2_X1  g0908(.A(KEYINPUT54), .B(G143), .ZN(new_n1109));
  OAI221_X1 g0909(.A(new_n360), .B1(new_n750), .B2(new_n1109), .C1(new_n818), .C2(new_n747), .ZN(new_n1110));
  NOR4_X1   g0910(.A1(new_n1105), .A2(new_n1107), .A3(new_n1108), .A4(new_n1110), .ZN(new_n1111));
  INV_X1    g0911(.A(G125), .ZN(new_n1112));
  OAI221_X1 g0912(.A(new_n1111), .B1(new_n743), .B2(new_n201), .C1(new_n737), .C2(new_n1112), .ZN(new_n1113));
  NAND2_X1  g0913(.A1(new_n1101), .A2(new_n1102), .ZN(new_n1114));
  NAND3_X1  g0914(.A1(new_n1103), .A2(new_n1113), .A3(new_n1114), .ZN(new_n1115));
  AOI21_X1  g0915(.A(new_n1096), .B1(new_n1115), .B2(new_n726), .ZN(new_n1116));
  AOI21_X1  g0916(.A(new_n1094), .B1(new_n1095), .B2(new_n1116), .ZN(new_n1117));
  NAND2_X1  g0917(.A1(new_n1074), .A2(new_n1078), .ZN(new_n1118));
  NAND4_X1  g0918(.A1(new_n1091), .A2(new_n1085), .A3(new_n897), .A4(new_n1118), .ZN(new_n1119));
  NAND3_X1  g0919(.A1(new_n700), .A2(G330), .A3(new_n793), .ZN(new_n1120));
  AOI21_X1  g0920(.A(new_n1079), .B1(new_n1078), .B2(new_n1120), .ZN(new_n1121));
  INV_X1    g0921(.A(new_n898), .ZN(new_n1122));
  OAI21_X1  g0922(.A(new_n1119), .B1(new_n1121), .B2(new_n1122), .ZN(new_n1123));
  NAND3_X1  g0923(.A1(new_n444), .A2(G330), .A3(new_n842), .ZN(new_n1124));
  AND3_X1   g0924(.A1(new_n902), .A2(new_n629), .A3(new_n1124), .ZN(new_n1125));
  AND3_X1   g0925(.A1(new_n1123), .A2(new_n1125), .A3(KEYINPUT119), .ZN(new_n1126));
  AOI21_X1  g0926(.A(KEYINPUT119), .B1(new_n1123), .B2(new_n1125), .ZN(new_n1127));
  NOR2_X1   g0927(.A1(new_n1126), .A2(new_n1127), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n1128), .A2(new_n1093), .ZN(new_n1129));
  OAI211_X1 g0929(.A(new_n1092), .B(new_n1088), .C1(new_n1126), .C2(new_n1127), .ZN(new_n1130));
  NAND3_X1  g0930(.A1(new_n1129), .A2(new_n656), .A3(new_n1130), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n1117), .A2(new_n1131), .ZN(G378));
  NAND2_X1  g0932(.A1(new_n744), .A2(G58), .ZN(new_n1133));
  AOI211_X1 g0933(.A(new_n360), .B(new_n497), .C1(new_n753), .C2(G77), .ZN(new_n1134));
  OAI211_X1 g0934(.A(new_n1133), .B(new_n1134), .C1(new_n801), .C2(new_n737), .ZN(new_n1135));
  XNOR2_X1  g0935(.A(new_n1135), .B(KEYINPUT121), .ZN(new_n1136));
  OAI22_X1  g0936(.A1(new_n747), .A2(new_n576), .B1(new_n750), .B2(new_n419), .ZN(new_n1137));
  OAI22_X1  g0937(.A1(new_n482), .A2(new_n759), .B1(new_n803), .B2(new_n536), .ZN(new_n1138));
  AOI211_X1 g0938(.A(new_n1137), .B(new_n1138), .C1(G68), .C2(new_n764), .ZN(new_n1139));
  NAND3_X1  g0939(.A1(new_n1136), .A2(KEYINPUT58), .A3(new_n1139), .ZN(new_n1140));
  OAI221_X1 g0940(.A(new_n201), .B1(G33), .B2(G41), .C1(new_n497), .C2(new_n360), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n758), .A2(G128), .ZN(new_n1142));
  OAI21_X1  g0942(.A(new_n1142), .B1(new_n803), .B2(new_n1112), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n816), .A2(G137), .ZN(new_n1144));
  OAI221_X1 g0944(.A(new_n1144), .B1(new_n823), .B2(new_n747), .C1(new_n812), .C2(new_n1109), .ZN(new_n1145));
  AOI211_X1 g0945(.A(new_n1143), .B(new_n1145), .C1(G150), .C2(new_n764), .ZN(new_n1146));
  INV_X1    g0946(.A(KEYINPUT59), .ZN(new_n1147));
  NOR2_X1   g0947(.A1(new_n1146), .A2(new_n1147), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n1146), .A2(new_n1147), .ZN(new_n1149));
  AOI211_X1 g0949(.A(G33), .B(G41), .C1(new_n733), .C2(G124), .ZN(new_n1150));
  OAI211_X1 g0950(.A(new_n1149), .B(new_n1150), .C1(new_n1020), .C2(new_n743), .ZN(new_n1151));
  OAI211_X1 g0951(.A(new_n1140), .B(new_n1141), .C1(new_n1148), .C2(new_n1151), .ZN(new_n1152));
  AOI21_X1  g0952(.A(KEYINPUT58), .B1(new_n1136), .B2(new_n1139), .ZN(new_n1153));
  OAI21_X1  g0953(.A(new_n726), .B1(new_n1152), .B2(new_n1153), .ZN(new_n1154));
  OAI211_X1 g0954(.A(new_n1154), .B(new_n711), .C1(G50), .C2(new_n798), .ZN(new_n1155));
  NOR2_X1   g0955(.A1(new_n353), .A2(new_n635), .ZN(new_n1156));
  XOR2_X1   g0956(.A(new_n379), .B(new_n1156), .Z(new_n1157));
  XNOR2_X1  g0957(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1158));
  XNOR2_X1  g0958(.A(new_n1157), .B(new_n1158), .ZN(new_n1159));
  AOI21_X1  g0959(.A(new_n1155), .B1(new_n1159), .B2(new_n723), .ZN(new_n1160));
  OAI211_X1 g0960(.A(G330), .B(new_n885), .C1(new_n873), .C2(KEYINPUT40), .ZN(new_n1161));
  AND2_X1   g0961(.A1(new_n1161), .A2(new_n1159), .ZN(new_n1162));
  NOR2_X1   g0962(.A1(new_n1161), .A2(new_n1159), .ZN(new_n1163));
  OAI21_X1  g0963(.A(KEYINPUT122), .B1(new_n1162), .B2(new_n1163), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n1164), .A2(new_n901), .ZN(new_n1165));
  INV_X1    g0965(.A(new_n1159), .ZN(new_n1166));
  NAND4_X1  g0966(.A1(new_n874), .A2(new_n1166), .A3(G330), .A4(new_n885), .ZN(new_n1167));
  NAND2_X1  g0967(.A1(new_n1161), .A2(new_n1159), .ZN(new_n1168));
  NAND2_X1  g0968(.A1(new_n1167), .A2(new_n1168), .ZN(new_n1169));
  INV_X1    g0969(.A(new_n901), .ZN(new_n1170));
  NAND3_X1  g0970(.A1(new_n1169), .A2(KEYINPUT122), .A3(new_n1170), .ZN(new_n1171));
  NAND2_X1  g0971(.A1(new_n1165), .A2(new_n1171), .ZN(new_n1172));
  AOI21_X1  g0972(.A(new_n1160), .B1(new_n1172), .B2(new_n707), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n1130), .A2(new_n1125), .ZN(new_n1174));
  AOI21_X1  g0974(.A(KEYINPUT57), .B1(new_n1172), .B2(new_n1174), .ZN(new_n1175));
  INV_X1    g0975(.A(KEYINPUT57), .ZN(new_n1176));
  AOI21_X1  g0976(.A(new_n1176), .B1(new_n1130), .B2(new_n1125), .ZN(new_n1177));
  OAI21_X1  g0977(.A(new_n1170), .B1(new_n1162), .B2(new_n1163), .ZN(new_n1178));
  NAND3_X1  g0978(.A1(new_n1167), .A2(new_n901), .A3(new_n1168), .ZN(new_n1179));
  NAND2_X1  g0979(.A1(new_n1178), .A2(new_n1179), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n1177), .A2(new_n1180), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n1181), .A2(new_n656), .ZN(new_n1182));
  OAI21_X1  g0982(.A(new_n1173), .B1(new_n1175), .B2(new_n1182), .ZN(G375));
  NAND2_X1  g0983(.A1(new_n1123), .A2(new_n707), .ZN(new_n1184));
  INV_X1    g0984(.A(KEYINPUT123), .ZN(new_n1185));
  AOI21_X1  g0985(.A(new_n710), .B1(new_n203), .B2(new_n797), .ZN(new_n1186));
  INV_X1    g0986(.A(new_n726), .ZN(new_n1187));
  NAND2_X1  g0987(.A1(new_n738), .A2(G303), .ZN(new_n1188));
  OAI22_X1  g0988(.A1(new_n747), .A2(new_n536), .B1(new_n750), .B2(new_n482), .ZN(new_n1189));
  AOI211_X1 g0989(.A(new_n360), .B(new_n1189), .C1(G97), .C2(new_n753), .ZN(new_n1190));
  OAI221_X1 g0990(.A(new_n1019), .B1(new_n803), .B2(new_n507), .C1(new_n801), .C2(new_n759), .ZN(new_n1191));
  INV_X1    g0991(.A(new_n1191), .ZN(new_n1192));
  NAND4_X1  g0992(.A1(new_n1188), .A2(new_n988), .A3(new_n1190), .A4(new_n1192), .ZN(new_n1193));
  NAND2_X1  g0993(.A1(new_n738), .A2(G128), .ZN(new_n1194));
  INV_X1    g0994(.A(G150), .ZN(new_n1195));
  OAI22_X1  g0995(.A1(new_n747), .A2(new_n1109), .B1(new_n750), .B2(new_n1195), .ZN(new_n1196));
  AOI211_X1 g0996(.A(new_n315), .B(new_n1196), .C1(G159), .C2(new_n753), .ZN(new_n1197));
  OAI22_X1  g0997(.A1(new_n759), .A2(new_n818), .B1(new_n763), .B2(new_n201), .ZN(new_n1198));
  AOI21_X1  g0998(.A(new_n1198), .B1(G132), .B2(new_n756), .ZN(new_n1199));
  NAND4_X1  g0999(.A1(new_n1194), .A2(new_n1133), .A3(new_n1197), .A4(new_n1199), .ZN(new_n1200));
  AND2_X1   g1000(.A1(new_n1193), .A2(new_n1200), .ZN(new_n1201));
  OAI221_X1 g1001(.A(new_n1186), .B1(new_n1187), .B2(new_n1201), .C1(new_n841), .C2(new_n724), .ZN(new_n1202));
  AND3_X1   g1002(.A1(new_n1184), .A2(new_n1185), .A3(new_n1202), .ZN(new_n1203));
  AOI21_X1  g1003(.A(new_n1185), .B1(new_n1184), .B2(new_n1202), .ZN(new_n1204));
  NOR2_X1   g1004(.A1(new_n1203), .A2(new_n1204), .ZN(new_n1205));
  INV_X1    g1005(.A(new_n1205), .ZN(new_n1206));
  INV_X1    g1006(.A(new_n943), .ZN(new_n1207));
  OR2_X1    g1007(.A1(new_n1123), .A2(new_n1125), .ZN(new_n1208));
  NAND3_X1  g1008(.A1(new_n1128), .A2(new_n1207), .A3(new_n1208), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(new_n1206), .A2(new_n1209), .ZN(G381));
  INV_X1    g1010(.A(G390), .ZN(new_n1211));
  INV_X1    g1011(.A(G384), .ZN(new_n1212));
  NOR2_X1   g1012(.A1(G393), .A2(G396), .ZN(new_n1213));
  NAND3_X1  g1013(.A1(new_n1211), .A2(new_n1212), .A3(new_n1213), .ZN(new_n1214));
  NOR3_X1   g1014(.A1(new_n1214), .A2(G387), .A3(G381), .ZN(new_n1215));
  INV_X1    g1015(.A(G375), .ZN(new_n1216));
  INV_X1    g1016(.A(G378), .ZN(new_n1217));
  NAND3_X1  g1017(.A1(new_n1215), .A2(new_n1216), .A3(new_n1217), .ZN(G407));
  NAND2_X1  g1018(.A1(new_n636), .A2(G213), .ZN(new_n1219));
  INV_X1    g1019(.A(new_n1219), .ZN(new_n1220));
  NAND3_X1  g1020(.A1(new_n1216), .A2(new_n1217), .A3(new_n1220), .ZN(new_n1221));
  NAND3_X1  g1021(.A1(G407), .A2(new_n1221), .A3(G213), .ZN(G409));
  INV_X1    g1022(.A(KEYINPUT127), .ZN(new_n1223));
  INV_X1    g1023(.A(KEYINPUT126), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(new_n1211), .A2(G387), .ZN(new_n1225));
  NAND3_X1  g1025(.A1(G390), .A2(new_n974), .A3(new_n1000), .ZN(new_n1226));
  AOI21_X1  g1026(.A(new_n780), .B1(new_n1004), .B2(new_n1042), .ZN(new_n1227));
  NOR2_X1   g1027(.A1(new_n1213), .A2(new_n1227), .ZN(new_n1228));
  AND4_X1   g1028(.A1(new_n1224), .A2(new_n1225), .A3(new_n1226), .A4(new_n1228), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n1226), .A2(KEYINPUT126), .ZN(new_n1230));
  AOI22_X1  g1030(.A1(new_n1230), .A2(new_n1228), .B1(new_n1225), .B2(new_n1226), .ZN(new_n1231));
  NOR2_X1   g1031(.A1(new_n1229), .A2(new_n1231), .ZN(new_n1232));
  INV_X1    g1032(.A(KEYINPUT61), .ZN(new_n1233));
  OAI211_X1 g1033(.A(G378), .B(new_n1173), .C1(new_n1175), .C2(new_n1182), .ZN(new_n1234));
  AOI21_X1  g1034(.A(new_n1160), .B1(new_n1180), .B2(new_n707), .ZN(new_n1235));
  AOI21_X1  g1035(.A(new_n1170), .B1(new_n1169), .B2(KEYINPUT122), .ZN(new_n1236));
  INV_X1    g1036(.A(KEYINPUT122), .ZN(new_n1237));
  AOI211_X1 g1037(.A(new_n1237), .B(new_n901), .C1(new_n1167), .C2(new_n1168), .ZN(new_n1238));
  OAI21_X1  g1038(.A(new_n1174), .B1(new_n1236), .B2(new_n1238), .ZN(new_n1239));
  OAI21_X1  g1039(.A(new_n1235), .B1(new_n1239), .B2(new_n943), .ZN(new_n1240));
  NAND2_X1  g1040(.A1(new_n1240), .A2(new_n1217), .ZN(new_n1241));
  AOI21_X1  g1041(.A(new_n1220), .B1(new_n1234), .B2(new_n1241), .ZN(new_n1242));
  NAND2_X1  g1042(.A1(new_n1220), .A2(G2897), .ZN(new_n1243));
  NOR2_X1   g1043(.A1(new_n1123), .A2(new_n1125), .ZN(new_n1244));
  OAI21_X1  g1044(.A(new_n656), .B1(new_n1244), .B2(KEYINPUT60), .ZN(new_n1245));
  INV_X1    g1045(.A(new_n1245), .ZN(new_n1246));
  NOR3_X1   g1046(.A1(new_n1126), .A2(new_n1127), .A3(new_n1244), .ZN(new_n1247));
  INV_X1    g1047(.A(KEYINPUT60), .ZN(new_n1248));
  OAI21_X1  g1048(.A(new_n1246), .B1(new_n1247), .B2(new_n1248), .ZN(new_n1249));
  NAND3_X1  g1049(.A1(new_n1249), .A2(new_n1206), .A3(G384), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(new_n1123), .A2(new_n1125), .ZN(new_n1251));
  INV_X1    g1051(.A(KEYINPUT119), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(new_n1251), .A2(new_n1252), .ZN(new_n1253));
  NAND3_X1  g1053(.A1(new_n1123), .A2(new_n1125), .A3(KEYINPUT119), .ZN(new_n1254));
  NAND3_X1  g1054(.A1(new_n1253), .A2(new_n1208), .A3(new_n1254), .ZN(new_n1255));
  AOI21_X1  g1055(.A(new_n1245), .B1(new_n1255), .B2(KEYINPUT60), .ZN(new_n1256));
  OAI21_X1  g1056(.A(new_n1212), .B1(new_n1256), .B2(new_n1205), .ZN(new_n1257));
  INV_X1    g1057(.A(KEYINPUT125), .ZN(new_n1258));
  AND3_X1   g1058(.A1(new_n1250), .A2(new_n1257), .A3(new_n1258), .ZN(new_n1259));
  AOI21_X1  g1059(.A(new_n1258), .B1(new_n1250), .B2(new_n1257), .ZN(new_n1260));
  OAI21_X1  g1060(.A(new_n1243), .B1(new_n1259), .B2(new_n1260), .ZN(new_n1261));
  NAND3_X1  g1061(.A1(new_n1250), .A2(new_n1257), .A3(new_n1258), .ZN(new_n1262));
  INV_X1    g1062(.A(new_n1243), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n1262), .A2(new_n1263), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(new_n1261), .A2(new_n1264), .ZN(new_n1265));
  OAI21_X1  g1065(.A(new_n1233), .B1(new_n1242), .B2(new_n1265), .ZN(new_n1266));
  INV_X1    g1066(.A(KEYINPUT62), .ZN(new_n1267));
  AOI21_X1  g1067(.A(G384), .B1(new_n1249), .B2(new_n1206), .ZN(new_n1268));
  NOR3_X1   g1068(.A1(new_n1256), .A2(new_n1205), .A3(new_n1212), .ZN(new_n1269));
  NOR2_X1   g1069(.A1(new_n1268), .A2(new_n1269), .ZN(new_n1270));
  AOI21_X1  g1070(.A(new_n1267), .B1(new_n1242), .B2(new_n1270), .ZN(new_n1271));
  NOR2_X1   g1071(.A1(new_n1266), .A2(new_n1271), .ZN(new_n1272));
  NAND2_X1  g1072(.A1(new_n1234), .A2(new_n1241), .ZN(new_n1273));
  NAND3_X1  g1073(.A1(new_n1273), .A2(new_n1219), .A3(new_n1270), .ZN(new_n1274));
  NOR2_X1   g1074(.A1(new_n1274), .A2(KEYINPUT62), .ZN(new_n1275));
  INV_X1    g1075(.A(new_n1275), .ZN(new_n1276));
  AOI21_X1  g1076(.A(new_n1232), .B1(new_n1272), .B2(new_n1276), .ZN(new_n1277));
  INV_X1    g1077(.A(KEYINPUT63), .ZN(new_n1278));
  NAND2_X1  g1078(.A1(new_n1274), .A2(new_n1278), .ZN(new_n1279));
  NAND3_X1  g1079(.A1(new_n1242), .A2(KEYINPUT63), .A3(new_n1270), .ZN(new_n1280));
  NOR3_X1   g1080(.A1(new_n1229), .A2(new_n1231), .A3(KEYINPUT61), .ZN(new_n1281));
  NAND3_X1  g1081(.A1(new_n1279), .A2(new_n1280), .A3(new_n1281), .ZN(new_n1282));
  OAI21_X1  g1082(.A(KEYINPUT125), .B1(new_n1268), .B2(new_n1269), .ZN(new_n1283));
  AOI21_X1  g1083(.A(new_n1263), .B1(new_n1283), .B2(new_n1262), .ZN(new_n1284));
  INV_X1    g1084(.A(new_n1264), .ZN(new_n1285));
  NOR2_X1   g1085(.A1(new_n1284), .A2(new_n1285), .ZN(new_n1286));
  OAI21_X1  g1086(.A(new_n1286), .B1(new_n1242), .B2(KEYINPUT124), .ZN(new_n1287));
  INV_X1    g1087(.A(KEYINPUT124), .ZN(new_n1288));
  AOI211_X1 g1088(.A(new_n1288), .B(new_n1220), .C1(new_n1234), .C2(new_n1241), .ZN(new_n1289));
  NOR2_X1   g1089(.A1(new_n1287), .A2(new_n1289), .ZN(new_n1290));
  NOR2_X1   g1090(.A1(new_n1282), .A2(new_n1290), .ZN(new_n1291));
  OAI21_X1  g1091(.A(new_n1223), .B1(new_n1277), .B2(new_n1291), .ZN(new_n1292));
  NAND2_X1  g1092(.A1(new_n1273), .A2(new_n1219), .ZN(new_n1293));
  NAND2_X1  g1093(.A1(new_n1293), .A2(new_n1288), .ZN(new_n1294));
  NAND2_X1  g1094(.A1(new_n1242), .A2(KEYINPUT124), .ZN(new_n1295));
  NAND3_X1  g1095(.A1(new_n1294), .A2(new_n1295), .A3(new_n1286), .ZN(new_n1296));
  NAND2_X1  g1096(.A1(new_n1230), .A2(new_n1228), .ZN(new_n1297));
  NAND2_X1  g1097(.A1(new_n1225), .A2(new_n1226), .ZN(new_n1298));
  NAND2_X1  g1098(.A1(new_n1297), .A2(new_n1298), .ZN(new_n1299));
  NAND4_X1  g1099(.A1(new_n1230), .A2(new_n1226), .A3(new_n1225), .A4(new_n1228), .ZN(new_n1300));
  NAND3_X1  g1100(.A1(new_n1299), .A2(new_n1233), .A3(new_n1300), .ZN(new_n1301));
  AOI21_X1  g1101(.A(new_n1301), .B1(new_n1278), .B2(new_n1274), .ZN(new_n1302));
  NAND3_X1  g1102(.A1(new_n1296), .A2(new_n1302), .A3(new_n1280), .ZN(new_n1303));
  NOR3_X1   g1103(.A1(new_n1275), .A2(new_n1266), .A3(new_n1271), .ZN(new_n1304));
  OAI211_X1 g1104(.A(new_n1303), .B(KEYINPUT127), .C1(new_n1232), .C2(new_n1304), .ZN(new_n1305));
  NAND2_X1  g1105(.A1(new_n1292), .A2(new_n1305), .ZN(G405));
  NAND2_X1  g1106(.A1(G375), .A2(new_n1217), .ZN(new_n1307));
  NAND2_X1  g1107(.A1(new_n1307), .A2(new_n1234), .ZN(new_n1308));
  INV_X1    g1108(.A(new_n1270), .ZN(new_n1309));
  XNOR2_X1  g1109(.A(new_n1308), .B(new_n1309), .ZN(new_n1310));
  XNOR2_X1  g1110(.A(new_n1310), .B(new_n1232), .ZN(G402));
endmodule


