//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 0 0 0 0 0 1 0 0 1 0 1 1 1 1 0 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 1 1 1 0 1 1 1 1 1 1 1 1 0 0 1 1 0 1 0 1 1 1 1 0 0 1 0 0' ..
//Module:
 module locked_locked_c1355( 
    KEYINPUT0, KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5,
    KEYINPUT6, KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11,
    KEYINPUT12, KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
    KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23,
    KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29,
    KEYINPUT30, KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35,
    KEYINPUT36, KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41,
    KEYINPUT42, KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
    KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53,
    KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59,
    KEYINPUT60, KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat,
    G22gat, G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat,
    G85gat, G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat,
    G141gat, G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat,
    G197gat, G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat,
    G229gat, G230gat, G231gat, G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  , KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64);
input KEYINPUT64;
input KEYINPUT65;
input KEYINPUT66;
input KEYINPUT67;
input KEYINPUT68;
input KEYINPUT69;
input KEYINPUT70;
input KEYINPUT71;
input KEYINPUT72;
input KEYINPUT73;
input KEYINPUT74;
input KEYINPUT75;
input KEYINPUT76;
input KEYINPUT77;
input KEYINPUT78;
input KEYINPUT79;
input KEYINPUT80;
input KEYINPUT81;
input KEYINPUT82;
input KEYINPUT83;
input KEYINPUT84;
input KEYINPUT85;
input KEYINPUT86;
input KEYINPUT87;
input KEYINPUT88;
input KEYINPUT89;
input KEYINPUT90;
input KEYINPUT91;
input KEYINPUT92;
input KEYINPUT93;
input KEYINPUT94;
input KEYINPUT95;
input KEYINPUT96;
input KEYINPUT97;
input KEYINPUT98;
input KEYINPUT99;
input KEYINPUT100;
input KEYINPUT101;
input KEYINPUT102;
input KEYINPUT103;
input KEYINPUT104;
input KEYINPUT105;
input KEYINPUT106;
input KEYINPUT107;
input KEYINPUT108;
input KEYINPUT109;
input KEYINPUT110;
input KEYINPUT111;
input KEYINPUT112;
input KEYINPUT113;
input KEYINPUT114;
input KEYINPUT115;
input KEYINPUT116;
input KEYINPUT117;
input KEYINPUT118;
input KEYINPUT119;
input KEYINPUT120;
input KEYINPUT121;
input KEYINPUT122;
input KEYINPUT123;
input KEYINPUT124;
input KEYINPUT125;
input KEYINPUT126;
input KEYINPUT127;
//Header:
   input  KEYINPUT0, KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4,
    KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10,
    KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16,
    KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
    KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28,
    KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34,
    KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40,
    KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46,
    KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
    KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58,
    KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat,
    G8gat, G15gat, G22gat, G29gat, G36gat, G43gat, G50gat, G57gat, G64gat,
    G71gat, G78gat, G85gat, G92gat, G99gat, G106gat, G113gat, G120gat,
    G127gat, G134gat, G141gat, G148gat, G155gat, G162gat, G169gat, G176gat,
    G183gat, G190gat, G197gat, G204gat, G211gat, G218gat, G225gat, G226gat,
    G227gat, G228gat, G229gat, G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n138, new_n139, new_n140, new_n141, new_n142, new_n143, new_n144,
    new_n145, new_n146, new_n147, new_n148, new_n149, new_n150, new_n151,
    new_n152, new_n153, new_n154, new_n155, new_n156, new_n157, new_n158,
    new_n159, new_n160, new_n161, new_n162, new_n163, new_n164, new_n165,
    new_n166, new_n167, new_n168, new_n169, new_n170, new_n171, new_n172,
    new_n173, new_n174, new_n175, new_n176, new_n177, new_n178, new_n179,
    new_n180, new_n181, new_n182, new_n183, new_n184, new_n185, new_n186,
    new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n521, new_n522, new_n523, new_n524,
    new_n526, new_n527, new_n529, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n536, new_n537, new_n538, new_n539, new_n540,
    new_n541, new_n542, new_n543, new_n544, new_n545, new_n547, new_n548,
    new_n549, new_n550, new_n552, new_n553, new_n554, new_n555, new_n556,
    new_n557, new_n558, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n570, new_n571, new_n572,
    new_n573, new_n575, new_n576, new_n577, new_n578, new_n579, new_n581,
    new_n582, new_n583, new_n584, new_n586, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n599, new_n600, new_n601, new_n602, new_n603, new_n604, new_n605,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n612, new_n613,
    new_n614, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n652, new_n653, new_n655, new_n656, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n702, new_n703, new_n705, new_n706,
    new_n708, new_n709, new_n710, new_n711, new_n712, new_n713, new_n714,
    new_n715, new_n717, new_n718, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n727, new_n728, new_n729, new_n730, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n747, new_n748,
    new_n749, new_n750, new_n752, new_n753, new_n754;
wire RLL_wire_A_64;
wire RLL_wire_A_65;
wire RLL_wire_A_66;
wire RLL_wire_A_67;
wire RLL_wire_A_68;
wire RLL_wire_A_69;
wire RLL_wire_A_70;
wire RLL_wire_A_71;
wire RLL_wire_A_72;
wire RLL_wire_A_73;
wire RLL_wire_A_74;
wire RLL_wire_A_75;
wire RLL_wire_A_76;
wire RLL_wire_A_77;
wire RLL_wire_A_78;
wire RLL_wire_A_79;
wire RLL_wire_A_80;
wire RLL_wire_A_81;
wire RLL_wire_A_82;
wire RLL_wire_A_83;
wire RLL_wire_A_84;
wire RLL_wire_A_85;
wire RLL_wire_A_86;
wire RLL_wire_A_87;
wire RLL_wire_A_88;
wire RLL_wire_A_89;
wire RLL_wire_A_90;
wire RLL_wire_A_91;
wire RLL_wire_A_92;
wire RLL_wire_A_93;
wire RLL_wire_A_94;
wire RLL_wire_A_95;
wire RLL_wire_A_96;
wire RLL_wire_A_97;
wire RLL_wire_A_98;
wire RLL_wire_A_99;
wire RLL_wire_A_100;
wire RLL_wire_A_101;
wire RLL_wire_A_102;
wire RLL_wire_A_103;
wire RLL_wire_A_104;
wire RLL_wire_A_105;
wire RLL_wire_A_106;
wire RLL_wire_A_107;
wire RLL_wire_A_108;
wire RLL_wire_A_109;
wire RLL_wire_A_110;
wire RLL_wire_A_111;
wire RLL_wire_A_112;
wire RLL_wire_A_113;
wire RLL_wire_A_114;
wire RLL_wire_A_115;
wire RLL_wire_A_116;
wire RLL_wire_A_117;
wire RLL_wire_A_118;
wire RLL_wire_A_119;
wire RLL_wire_A_120;
wire RLL_wire_A_121;
wire RLL_wire_A_122;
wire RLL_wire_A_123;
wire RLL_wire_A_124;
wire RLL_wire_A_125;
wire RLL_wire_A_126;
wire RLL_wire_A_127;

//Body:
  NAND2_X1  g000(.A1(G227gat), .A2(G233gat), .ZN(new_n138));
  INV_X1    g001(.A(new_n138), .ZN(RLL_wire_A_64));
  XOR2_X1 RLL_XOR_64 (.A(RLL_wire_A_64), .B(KEYINPUT64), .Z(new_n139) );
  INV_X1    g002(.A(KEYINPUT25), .ZN(new_n140));
  AND3_X1   g003(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n141));
  AOI21_X1  g004(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n142));
  NOR2_X1   g005(.A1(G183gat), .A2(G190gat), .ZN(new_n143));
  NOR3_X1   g006(.A1(new_n141), .A2(new_n142), .A3(new_n143), .ZN(RLL_wire_A_65));
  XNOR2_X1 RLL_XNOR_65 (.A(RLL_wire_A_65), .B(KEYINPUT65), .ZN(new_n144) );
  INV_X1    g007(.A(G169gat), .ZN(RLL_wire_A_66));
  XNOR2_X1 RLL_XNOR_66 (.A(RLL_wire_A_66), .B(KEYINPUT66), .ZN(new_n145) );
  INV_X1    g008(.A(G176gat), .ZN(new_n146));
  NAND3_X1  g009(.A1(new_n145), .A2(new_n146), .A3(KEYINPUT23), .ZN(new_n147));
  INV_X1    g010(.A(KEYINPUT23), .ZN(new_n148));
  OAI21_X1  g011(.A(new_n148), .B1(G169gat), .B2(G176gat), .ZN(new_n149));
  NAND2_X1  g012(.A1(G169gat), .A2(G176gat), .ZN(RLL_wire_A_67));
  XOR2_X1 RLL_XOR_67 (.A(RLL_wire_A_67), .B(KEYINPUT67), .Z(new_n150) );
  NAND3_X1  g013(.A1(new_n147), .A2(new_n149), .A3(new_n150), .ZN(new_n151));
  OAI21_X1  g014(.A(new_n140), .B1(new_n144), .B2(new_n151), .ZN(new_n152));
  INV_X1    g015(.A(new_n150), .ZN(new_n153));
  NOR2_X1   g016(.A1(G169gat), .A2(G176gat), .ZN(new_n154));
  AOI21_X1  g017(.A(new_n153), .B1(KEYINPUT23), .B2(new_n154), .ZN(new_n155));
  NAND2_X1  g018(.A1(G183gat), .A2(G190gat), .ZN(new_n156));
  INV_X1    g019(.A(KEYINPUT24), .ZN(new_n157));
  NAND2_X1  g020(.A1(new_n156), .A2(new_n157), .ZN(RLL_wire_A_68));
  XNOR2_X1 RLL_XNOR_68 (.A(RLL_wire_A_68), .B(KEYINPUT68), .ZN(new_n158) );
  NAND3_X1  g021(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n159));
  INV_X1    g022(.A(G183gat), .ZN(new_n160));
  INV_X1    g023(.A(G190gat), .ZN(RLL_wire_A_69));
  XNOR2_X1 RLL_XNOR_69 (.A(RLL_wire_A_69), .B(KEYINPUT69), .ZN(new_n161) );
  NAND2_X1  g024(.A1(new_n160), .A2(new_n161), .ZN(new_n162));
  NAND3_X1  g025(.A1(new_n158), .A2(new_n159), .A3(new_n162), .ZN(new_n163));
  NAND4_X1  g026(.A1(new_n155), .A2(new_n163), .A3(KEYINPUT25), .A4(new_n149), .ZN(new_n164));
  NAND2_X1  g027(.A1(new_n152), .A2(new_n164), .ZN(RLL_wire_A_70));
  XOR2_X1 RLL_XOR_70 (.A(RLL_wire_A_70), .B(KEYINPUT70), .Z(new_n165) );
  NAND2_X1  g028(.A1(new_n160), .A2(KEYINPUT27), .ZN(new_n166));
  INV_X1    g029(.A(KEYINPUT27), .ZN(new_n167));
  NAND2_X1  g030(.A1(new_n167), .A2(G183gat), .ZN(new_n168));
  NAND3_X1  g031(.A1(new_n166), .A2(new_n168), .A3(new_n161), .ZN(new_n169));
  INV_X1    g032(.A(KEYINPUT28), .ZN(new_n170));
  NAND2_X1  g033(.A1(new_n169), .A2(new_n170), .ZN(new_n171));
  XNOR2_X1  g034(.A(KEYINPUT27), .B(G183gat), .ZN(new_n172));
  NAND3_X1  g035(.A1(new_n172), .A2(KEYINPUT28), .A3(new_n161), .ZN(new_n173));
  NAND2_X1  g036(.A1(new_n171), .A2(new_n173), .ZN(RLL_wire_A_71));
  XOR2_X1 RLL_XOR_71 (.A(RLL_wire_A_71), .B(KEYINPUT71), .Z(new_n174) );
  OAI21_X1  g037(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n175));
  AND2_X1   g038(.A1(new_n175), .A2(new_n150), .ZN(new_n176));
  INV_X1    g039(.A(KEYINPUT26), .ZN(new_n177));
  NAND2_X1  g040(.A1(new_n154), .A2(new_n177), .ZN(new_n178));
  AOI22_X1  g041(.A1(new_n176), .A2(new_n178), .B1(G183gat), .B2(G190gat), .ZN(new_n179));
  NAND2_X1  g042(.A1(new_n174), .A2(new_n179), .ZN(new_n180));
  INV_X1    g043(.A(G134gat), .ZN(new_n181));
  NAND2_X1  g044(.A1(new_n181), .A2(G127gat), .ZN(new_n182));
  INV_X1    g045(.A(G127gat), .ZN(new_n183));
  NAND2_X1  g046(.A1(new_n183), .A2(G134gat), .ZN(new_n184));
  NAND2_X1  g047(.A1(new_n182), .A2(new_n184), .ZN(new_n185));
  XNOR2_X1  g048(.A(G113gat), .B(G120gat), .ZN(new_n186));
  OAI21_X1  g049(.A(new_n185), .B1(new_n186), .B2(KEYINPUT1), .ZN(new_n187));
  INV_X1    g050(.A(G120gat), .ZN(new_n188));
  NAND2_X1  g051(.A1(new_n188), .A2(G113gat), .ZN(new_n189));
  INV_X1    g052(.A(G113gat), .ZN(new_n190));
  NAND2_X1  g053(.A1(new_n190), .A2(G120gat), .ZN(new_n191));
  NAND2_X1  g054(.A1(new_n189), .A2(new_n191), .ZN(new_n192));
  XNOR2_X1  g055(.A(G127gat), .B(G134gat), .ZN(new_n193));
  INV_X1    g056(.A(KEYINPUT1), .ZN(new_n194));
  NAND3_X1  g057(.A1(new_n192), .A2(new_n193), .A3(new_n194), .ZN(new_n195));
  AND2_X1   g058(.A1(new_n187), .A2(new_n195), .ZN(new_n196));
  AND3_X1   g059(.A1(new_n165), .A2(new_n180), .A3(new_n196), .ZN(new_n197));
  AOI21_X1  g060(.A(new_n196), .B1(new_n165), .B2(new_n180), .ZN(new_n198));
  OAI21_X1  g061(.A(new_n139), .B1(new_n197), .B2(new_n198), .ZN(new_n199));
  INV_X1    g062(.A(KEYINPUT33), .ZN(RLL_wire_A_72));
  XOR2_X1 RLL_XOR_72 (.A(RLL_wire_A_72), .B(KEYINPUT72), .Z(new_n200) );
  NAND2_X1  g063(.A1(new_n199), .A2(new_n200), .ZN(new_n201));
  NAND2_X1  g064(.A1(new_n199), .A2(KEYINPUT32), .ZN(new_n202));
  XOR2_X1   g065(.A(G15gat), .B(G43gat), .Z(new_n203));
  XNOR2_X1  g066(.A(G71gat), .B(G99gat), .ZN(new_n204));
  XNOR2_X1  g067(.A(new_n203), .B(new_n204), .ZN(new_n205));
  NAND3_X1  g068(.A1(new_n201), .A2(new_n202), .A3(new_n205), .ZN(new_n206));
  INV_X1    g069(.A(new_n205), .ZN(new_n207));
  OAI211_X1 g070(.A(new_n199), .B(KEYINPUT32), .C1(new_n200), .C2(new_n207), .ZN(new_n208));
  NAND2_X1  g071(.A1(new_n206), .A2(new_n208), .ZN(new_n209));
  INV_X1    g072(.A(KEYINPUT34), .ZN(new_n210));
  NOR2_X1   g073(.A1(new_n197), .A2(new_n198), .ZN(new_n211));
  AOI21_X1  g074(.A(new_n210), .B1(new_n211), .B2(new_n138), .ZN(new_n212));
  NOR4_X1   g075(.A1(new_n197), .A2(new_n198), .A3(KEYINPUT34), .A4(new_n139), .ZN(new_n213));
  NOR2_X1   g076(.A1(new_n212), .A2(new_n213), .ZN(RLL_wire_A_73));
  XOR2_X1 RLL_XOR_73 (.A(RLL_wire_A_73), .B(KEYINPUT73), .Z(new_n214) );
  INV_X1    g077(.A(new_n214), .ZN(new_n215));
  NAND2_X1  g078(.A1(new_n209), .A2(new_n215), .ZN(new_n216));
  NAND3_X1  g079(.A1(new_n214), .A2(new_n206), .A3(new_n208), .ZN(new_n217));
  NAND3_X1  g080(.A1(new_n216), .A2(KEYINPUT36), .A3(new_n217), .ZN(new_n218));
  INV_X1    g081(.A(KEYINPUT36), .ZN(new_n219));
  INV_X1    g082(.A(new_n217), .ZN(new_n220));
  AOI21_X1  g083(.A(new_n214), .B1(new_n206), .B2(new_n208), .ZN(new_n221));
  OAI21_X1  g084(.A(new_n219), .B1(new_n220), .B2(new_n221), .ZN(new_n222));
  XNOR2_X1  g085(.A(G197gat), .B(G204gat), .ZN(new_n223));
  INV_X1    g086(.A(KEYINPUT22), .ZN(new_n224));
  INV_X1    g087(.A(G211gat), .ZN(new_n225));
  INV_X1    g088(.A(G218gat), .ZN(new_n226));
  OAI21_X1  g089(.A(new_n224), .B1(new_n225), .B2(new_n226), .ZN(new_n227));
  NAND2_X1  g090(.A1(new_n223), .A2(new_n227), .ZN(new_n228));
  XNOR2_X1  g091(.A(G211gat), .B(G218gat), .ZN(new_n229));
  INV_X1    g092(.A(new_n229), .ZN(new_n230));
  NAND2_X1  g093(.A1(new_n228), .A2(new_n230), .ZN(new_n231));
  NAND3_X1  g094(.A1(new_n229), .A2(new_n223), .A3(new_n227), .ZN(new_n232));
  NAND2_X1  g095(.A1(new_n231), .A2(new_n232), .ZN(new_n233));
  INV_X1    g096(.A(new_n233), .ZN(new_n234));
  NAND2_X1  g097(.A1(G226gat), .A2(G233gat), .ZN(new_n235));
  INV_X1    g098(.A(new_n235), .ZN(new_n236));
  NAND2_X1  g099(.A1(new_n165), .A2(new_n180), .ZN(RLL_wire_A_74));
  XOR2_X1 RLL_XOR_74 (.A(RLL_wire_A_74), .B(KEYINPUT74), .Z(new_n237) );
  INV_X1    g100(.A(KEYINPUT29), .ZN(new_n238));
  AOI21_X1  g101(.A(new_n236), .B1(new_n237), .B2(new_n238), .ZN(new_n239));
  AOI22_X1  g102(.A1(new_n152), .A2(new_n164), .B1(new_n174), .B2(new_n179), .ZN(new_n240));
  NOR2_X1   g103(.A1(new_n240), .A2(new_n235), .ZN(new_n241));
  OAI21_X1  g104(.A(new_n234), .B1(new_n239), .B2(new_n241), .ZN(new_n242));
  OAI21_X1  g105(.A(new_n235), .B1(new_n240), .B2(KEYINPUT29), .ZN(new_n243));
  NAND2_X1  g106(.A1(new_n237), .A2(new_n236), .ZN(RLL_wire_A_75));
  XNOR2_X1 RLL_XNOR_75 (.A(RLL_wire_A_75), .B(KEYINPUT75), .ZN(new_n244) );
  NAND3_X1  g107(.A1(new_n243), .A2(new_n233), .A3(new_n244), .ZN(new_n245));
  NAND2_X1  g108(.A1(new_n242), .A2(new_n245), .ZN(new_n246));
  XNOR2_X1  g109(.A(G8gat), .B(G36gat), .ZN(new_n247));
  XNOR2_X1  g110(.A(G64gat), .B(G92gat), .ZN(new_n248));
  XOR2_X1   g111(.A(new_n247), .B(new_n248), .Z(new_n249));
  INV_X1    g112(.A(new_n249), .ZN(new_n250));
  NAND2_X1  g113(.A1(new_n246), .A2(new_n250), .ZN(new_n251));
  NAND4_X1  g114(.A1(new_n242), .A2(new_n245), .A3(KEYINPUT30), .A4(new_n249), .ZN(new_n252));
  AND2_X1   g115(.A1(new_n251), .A2(new_n252), .ZN(new_n253));
  NAND3_X1  g116(.A1(new_n242), .A2(new_n245), .A3(new_n249), .ZN(new_n254));
  INV_X1    g117(.A(KEYINPUT30), .ZN(RLL_wire_A_76));
  XOR2_X1 RLL_XOR_76 (.A(RLL_wire_A_76), .B(KEYINPUT76), .Z(new_n255) );
  NAND2_X1  g118(.A1(new_n254), .A2(new_n255), .ZN(new_n256));
  AND2_X1   g119(.A1(G155gat), .A2(G162gat), .ZN(new_n257));
  NOR2_X1   g120(.A1(G155gat), .A2(G162gat), .ZN(new_n258));
  NOR2_X1   g121(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  XNOR2_X1  g122(.A(G141gat), .B(G148gat), .ZN(new_n260));
  INV_X1    g123(.A(KEYINPUT2), .ZN(new_n261));
  AOI21_X1  g124(.A(new_n261), .B1(G155gat), .B2(G162gat), .ZN(new_n262));
  OAI21_X1  g125(.A(new_n259), .B1(new_n260), .B2(new_n262), .ZN(new_n263));
  INV_X1    g126(.A(G141gat), .ZN(new_n264));
  NAND2_X1  g127(.A1(new_n264), .A2(G148gat), .ZN(new_n265));
  INV_X1    g128(.A(G148gat), .ZN(new_n266));
  NAND2_X1  g129(.A1(new_n266), .A2(G141gat), .ZN(new_n267));
  NAND2_X1  g130(.A1(new_n265), .A2(new_n267), .ZN(RLL_wire_A_77));
  XOR2_X1 RLL_XOR_77 (.A(RLL_wire_A_77), .B(KEYINPUT77), .Z(new_n268) );
  XNOR2_X1  g131(.A(G155gat), .B(G162gat), .ZN(new_n269));
  INV_X1    g132(.A(G155gat), .ZN(RLL_wire_A_78));
  XNOR2_X1 RLL_XNOR_78 (.A(RLL_wire_A_78), .B(KEYINPUT78), .ZN(new_n270) );
  INV_X1    g133(.A(G162gat), .ZN(new_n271));
  OAI21_X1  g134(.A(KEYINPUT2), .B1(new_n270), .B2(new_n271), .ZN(new_n272));
  NAND3_X1  g135(.A1(new_n268), .A2(new_n269), .A3(new_n272), .ZN(new_n273));
  NAND2_X1  g136(.A1(new_n263), .A2(new_n273), .ZN(new_n274));
  NAND2_X1  g137(.A1(new_n274), .A2(KEYINPUT3), .ZN(new_n275));
  NAND2_X1  g138(.A1(new_n187), .A2(new_n195), .ZN(new_n276));
  INV_X1    g139(.A(KEYINPUT3), .ZN(new_n277));
  NAND3_X1  g140(.A1(new_n263), .A2(new_n273), .A3(new_n277), .ZN(new_n278));
  NAND3_X1  g141(.A1(new_n275), .A2(new_n276), .A3(new_n278), .ZN(new_n279));
  NAND2_X1  g142(.A1(G225gat), .A2(G233gat), .ZN(new_n280));
  INV_X1    g143(.A(KEYINPUT4), .ZN(new_n281));
  AND2_X1   g144(.A1(new_n263), .A2(new_n273), .ZN(new_n282));
  AOI21_X1  g145(.A(new_n281), .B1(new_n282), .B2(new_n196), .ZN(new_n283));
  NAND4_X1  g146(.A1(new_n263), .A2(new_n187), .A3(new_n273), .A4(new_n195), .ZN(new_n284));
  NOR2_X1   g147(.A1(new_n284), .A2(KEYINPUT4), .ZN(new_n285));
  OAI211_X1 g148(.A(new_n279), .B(new_n280), .C1(new_n283), .C2(new_n285), .ZN(new_n286));
  NAND2_X1  g149(.A1(new_n274), .A2(new_n276), .ZN(new_n287));
  AOI21_X1  g150(.A(new_n280), .B1(new_n287), .B2(new_n284), .ZN(new_n288));
  INV_X1    g151(.A(KEYINPUT5), .ZN(new_n289));
  NOR2_X1   g152(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  NAND2_X1  g153(.A1(new_n286), .A2(new_n290), .ZN(new_n291));
  XOR2_X1   g154(.A(G1gat), .B(G29gat), .Z(RLL_wire_A_79));
  XOR2_X1 RLL_XOR_79 (.A(RLL_wire_A_79), .B(KEYINPUT79), .Z(new_n292) );
  XNOR2_X1  g155(.A(new_n292), .B(KEYINPUT0), .ZN(new_n293));
  XNOR2_X1  g156(.A(G57gat), .B(G85gat), .ZN(new_n294));
  XNOR2_X1  g157(.A(new_n293), .B(new_n294), .ZN(new_n295));
  NAND3_X1  g158(.A1(new_n282), .A2(new_n196), .A3(new_n281), .ZN(new_n296));
  NAND2_X1  g159(.A1(new_n284), .A2(KEYINPUT4), .ZN(new_n297));
  NAND2_X1  g160(.A1(new_n296), .A2(new_n297), .ZN(new_n298));
  NAND4_X1  g161(.A1(new_n298), .A2(new_n289), .A3(new_n280), .A4(new_n279), .ZN(new_n299));
  NAND3_X1  g162(.A1(new_n291), .A2(new_n295), .A3(new_n299), .ZN(new_n300));
  INV_X1    g163(.A(KEYINPUT6), .ZN(new_n301));
  NAND2_X1  g164(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  AOI21_X1  g165(.A(new_n295), .B1(new_n291), .B2(new_n299), .ZN(new_n303));
  NOR2_X1   g166(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  AOI211_X1 g167(.A(new_n301), .B(new_n295), .C1(new_n291), .C2(new_n299), .ZN(new_n305));
  OAI211_X1 g168(.A(new_n253), .B(new_n256), .C1(new_n304), .C2(new_n305), .ZN(new_n306));
  XNOR2_X1  g169(.A(G78gat), .B(G106gat), .ZN(new_n307));
  XNOR2_X1  g170(.A(new_n307), .B(KEYINPUT31), .ZN(new_n308));
  XNOR2_X1  g171(.A(new_n308), .B(G50gat), .ZN(new_n309));
  INV_X1    g172(.A(new_n309), .ZN(new_n310));
  NAND2_X1  g173(.A1(G228gat), .A2(G233gat), .ZN(new_n311));
  INV_X1    g174(.A(new_n232), .ZN(RLL_wire_A_80));
  XNOR2_X1 RLL_XNOR_80 (.A(RLL_wire_A_80), .B(KEYINPUT80), .ZN(new_n312) );
  AOI21_X1  g175(.A(new_n229), .B1(new_n227), .B2(new_n223), .ZN(new_n313));
  OAI21_X1  g176(.A(new_n238), .B1(new_n312), .B2(new_n313), .ZN(new_n314));
  AOI21_X1  g177(.A(new_n282), .B1(new_n314), .B2(new_n277), .ZN(new_n315));
  AOI21_X1  g178(.A(new_n233), .B1(new_n238), .B2(new_n278), .ZN(new_n316));
  OAI21_X1  g179(.A(new_n311), .B1(new_n315), .B2(new_n316), .ZN(new_n317));
  AOI21_X1  g180(.A(KEYINPUT29), .B1(new_n231), .B2(new_n232), .ZN(new_n318));
  OAI21_X1  g181(.A(new_n274), .B1(new_n318), .B2(KEYINPUT3), .ZN(new_n319));
  NAND2_X1  g182(.A1(new_n278), .A2(new_n238), .ZN(new_n320));
  NAND2_X1  g183(.A1(new_n320), .A2(new_n234), .ZN(RLL_wire_A_81));
  XNOR2_X1 RLL_XNOR_81 (.A(RLL_wire_A_81), .B(KEYINPUT81), .ZN(new_n321) );
  NAND4_X1  g184(.A1(new_n319), .A2(new_n321), .A3(G228gat), .A4(G233gat), .ZN(new_n322));
  INV_X1    g185(.A(G22gat), .ZN(new_n323));
  AND3_X1   g186(.A1(new_n317), .A2(new_n322), .A3(new_n323), .ZN(new_n324));
  AOI21_X1  g187(.A(new_n323), .B1(new_n317), .B2(new_n322), .ZN(RLL_wire_A_82));
  XNOR2_X1 RLL_XNOR_82 (.A(RLL_wire_A_82), .B(KEYINPUT82), .ZN(new_n325) );
  OAI21_X1  g188(.A(new_n310), .B1(new_n324), .B2(new_n325), .ZN(new_n326));
  NAND2_X1  g189(.A1(new_n317), .A2(new_n322), .ZN(new_n327));
  NAND2_X1  g190(.A1(new_n327), .A2(G22gat), .ZN(new_n328));
  NAND3_X1  g191(.A1(new_n317), .A2(new_n322), .A3(new_n323), .ZN(new_n329));
  NAND3_X1  g192(.A1(new_n328), .A2(new_n329), .A3(new_n309), .ZN(RLL_wire_A_83));
  XNOR2_X1 RLL_XNOR_83 (.A(RLL_wire_A_83), .B(KEYINPUT83), .ZN(new_n330) );
  NAND2_X1  g193(.A1(new_n326), .A2(new_n330), .ZN(new_n331));
  INV_X1    g194(.A(new_n331), .ZN(new_n332));
  AOI22_X1  g195(.A1(new_n218), .A2(new_n222), .B1(new_n306), .B2(new_n332), .ZN(new_n333));
  NAND3_X1  g196(.A1(new_n256), .A2(new_n251), .A3(new_n252), .ZN(new_n334));
  INV_X1    g197(.A(new_n295), .ZN(new_n335));
  AOI21_X1  g198(.A(new_n280), .B1(new_n298), .B2(new_n279), .ZN(new_n336));
  INV_X1    g199(.A(KEYINPUT39), .ZN(new_n337));
  AOI21_X1  g200(.A(new_n335), .B1(new_n336), .B2(new_n337), .ZN(RLL_wire_A_84));
  XOR2_X1 RLL_XOR_84 (.A(RLL_wire_A_84), .B(KEYINPUT84), .Z(new_n338) );
  NAND3_X1  g201(.A1(new_n287), .A2(new_n280), .A3(new_n284), .ZN(new_n339));
  NAND2_X1  g202(.A1(new_n339), .A2(KEYINPUT39), .ZN(new_n340));
  OAI21_X1  g203(.A(new_n338), .B1(new_n336), .B2(new_n340), .ZN(new_n341));
  INV_X1    g204(.A(KEYINPUT40), .ZN(new_n342));
  NAND2_X1  g205(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  NAND2_X1  g206(.A1(new_n291), .A2(new_n299), .ZN(RLL_wire_A_85));
  XNOR2_X1 RLL_XNOR_85 (.A(RLL_wire_A_85), .B(KEYINPUT85), .ZN(new_n344) );
  NAND2_X1  g207(.A1(new_n344), .A2(new_n335), .ZN(new_n345));
  OAI211_X1 g208(.A(new_n338), .B(KEYINPUT40), .C1(new_n336), .C2(new_n340), .ZN(new_n346));
  NAND4_X1  g209(.A1(new_n334), .A2(new_n343), .A3(new_n345), .A4(new_n346), .ZN(new_n347));
  NAND3_X1  g210(.A1(new_n345), .A2(new_n301), .A3(new_n300), .ZN(RLL_wire_A_86));
  XOR2_X1 RLL_XOR_86 (.A(RLL_wire_A_86), .B(KEYINPUT86), .Z(new_n348) );
  NOR3_X1   g211(.A1(new_n239), .A2(new_n241), .A3(new_n234), .ZN(new_n349));
  AOI21_X1  g212(.A(new_n233), .B1(new_n243), .B2(new_n244), .ZN(new_n350));
  OAI21_X1  g213(.A(KEYINPUT37), .B1(new_n349), .B2(new_n350), .ZN(new_n351));
  INV_X1    g214(.A(KEYINPUT38), .ZN(new_n352));
  INV_X1    g215(.A(KEYINPUT37), .ZN(new_n353));
  NAND3_X1  g216(.A1(new_n242), .A2(new_n353), .A3(new_n245), .ZN(new_n354));
  NAND4_X1  g217(.A1(new_n351), .A2(new_n352), .A3(new_n354), .A4(new_n250), .ZN(new_n355));
  INV_X1    g218(.A(new_n305), .ZN(new_n356));
  NAND4_X1  g219(.A1(new_n348), .A2(new_n355), .A3(new_n356), .A4(new_n254), .ZN(new_n357));
  AOI21_X1  g220(.A(new_n249), .B1(new_n246), .B2(KEYINPUT37), .ZN(new_n358));
  AOI21_X1  g221(.A(new_n352), .B1(new_n358), .B2(new_n354), .ZN(new_n359));
  OAI211_X1 g222(.A(new_n347), .B(new_n331), .C1(new_n357), .C2(new_n359), .ZN(new_n360));
  AOI21_X1  g223(.A(new_n334), .B1(new_n356), .B2(new_n348), .ZN(new_n361));
  NOR2_X1   g224(.A1(new_n220), .A2(new_n221), .ZN(new_n362));
  INV_X1    g225(.A(KEYINPUT35), .ZN(new_n363));
  NAND4_X1  g226(.A1(new_n361), .A2(new_n362), .A3(new_n363), .A4(new_n331), .ZN(new_n364));
  NAND3_X1  g227(.A1(new_n216), .A2(new_n331), .A3(new_n217), .ZN(new_n365));
  OAI21_X1  g228(.A(KEYINPUT35), .B1(new_n306), .B2(new_n365), .ZN(new_n366));
  AOI22_X1  g229(.A1(new_n333), .A2(new_n360), .B1(new_n364), .B2(new_n366), .ZN(new_n367));
  XNOR2_X1  g230(.A(G113gat), .B(G141gat), .ZN(new_n368));
  XNOR2_X1  g231(.A(new_n368), .B(KEYINPUT11), .ZN(new_n369));
  XOR2_X1   g232(.A(G169gat), .B(G197gat), .Z(new_n370));
  XNOR2_X1  g233(.A(new_n369), .B(new_n370), .ZN(new_n371));
  XNOR2_X1  g234(.A(new_n371), .B(KEYINPUT12), .ZN(new_n372));
  INV_X1    g235(.A(new_n372), .ZN(new_n373));
  XNOR2_X1  g236(.A(G43gat), .B(G50gat), .ZN(new_n374));
  OAI21_X1  g237(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n375));
  INV_X1    g238(.A(new_n375), .ZN(new_n376));
  NOR3_X1   g239(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n377));
  NOR2_X1   g240(.A1(new_n376), .A2(new_n377), .ZN(new_n378));
  INV_X1    g241(.A(G29gat), .ZN(new_n379));
  INV_X1    g242(.A(G36gat), .ZN(new_n380));
  NOR2_X1   g243(.A1(new_n379), .A2(new_n380), .ZN(new_n381));
  OAI211_X1 g244(.A(KEYINPUT15), .B(new_n374), .C1(new_n378), .C2(new_n381), .ZN(new_n382));
  NAND2_X1  g245(.A1(new_n374), .A2(KEYINPUT15), .ZN(new_n383));
  INV_X1    g246(.A(KEYINPUT15), .ZN(new_n384));
  INV_X1    g247(.A(G43gat), .ZN(RLL_wire_A_87));
  XNOR2_X1 RLL_XNOR_87 (.A(RLL_wire_A_87), .B(KEYINPUT87), .ZN(new_n385) );
  NOR2_X1   g248(.A1(new_n385), .A2(G50gat), .ZN(new_n386));
  INV_X1    g249(.A(G50gat), .ZN(new_n387));
  NOR2_X1   g250(.A1(new_n387), .A2(G43gat), .ZN(new_n388));
  OAI21_X1  g251(.A(new_n384), .B1(new_n386), .B2(new_n388), .ZN(new_n389));
  OR3_X1    g252(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(RLL_wire_A_88));
  XOR2_X1 RLL_XOR_88 (.A(RLL_wire_A_88), .B(KEYINPUT88), .Z(new_n390) );
  NAND2_X1  g253(.A1(new_n390), .A2(new_n375), .ZN(new_n391));
  INV_X1    g254(.A(new_n381), .ZN(new_n392));
  NAND4_X1  g255(.A1(new_n383), .A2(new_n389), .A3(new_n391), .A4(new_n392), .ZN(new_n393));
  NAND2_X1  g256(.A1(new_n382), .A2(new_n393), .ZN(new_n394));
  INV_X1    g257(.A(KEYINPUT17), .ZN(new_n395));
  NAND2_X1  g258(.A1(new_n394), .A2(new_n395), .ZN(new_n396));
  XNOR2_X1  g259(.A(G15gat), .B(G22gat), .ZN(new_n397));
  INV_X1    g260(.A(G1gat), .ZN(new_n398));
  NAND2_X1  g261(.A1(new_n398), .A2(KEYINPUT16), .ZN(new_n399));
  AND2_X1   g262(.A1(new_n397), .A2(new_n399), .ZN(new_n400));
  NOR2_X1   g263(.A1(new_n397), .A2(G1gat), .ZN(new_n401));
  OAI21_X1  g264(.A(G8gat), .B1(new_n400), .B2(new_n401), .ZN(new_n402));
  NAND2_X1  g265(.A1(new_n397), .A2(new_n399), .ZN(new_n403));
  INV_X1    g266(.A(G8gat), .ZN(new_n404));
  OAI211_X1 g267(.A(new_n403), .B(new_n404), .C1(G1gat), .C2(new_n397), .ZN(new_n405));
  AND2_X1   g268(.A1(new_n402), .A2(new_n405), .ZN(new_n406));
  NAND3_X1  g269(.A1(new_n382), .A2(new_n393), .A3(KEYINPUT17), .ZN(RLL_wire_A_89));
  XOR2_X1 RLL_XOR_89 (.A(RLL_wire_A_89), .B(KEYINPUT89), .Z(new_n407) );
  NAND3_X1  g270(.A1(new_n396), .A2(new_n406), .A3(new_n407), .ZN(new_n408));
  NAND2_X1  g271(.A1(G229gat), .A2(G233gat), .ZN(new_n409));
  NAND2_X1  g272(.A1(new_n402), .A2(new_n405), .ZN(new_n410));
  NAND2_X1  g273(.A1(new_n410), .A2(new_n394), .ZN(new_n411));
  NAND3_X1  g274(.A1(new_n408), .A2(new_n409), .A3(new_n411), .ZN(new_n412));
  INV_X1    g275(.A(KEYINPUT18), .ZN(new_n413));
  AND2_X1   g276(.A1(new_n412), .A2(new_n413), .ZN(new_n414));
  NAND4_X1  g277(.A1(new_n408), .A2(KEYINPUT18), .A3(new_n409), .A4(new_n411), .ZN(new_n415));
  XOR2_X1   g278(.A(new_n409), .B(KEYINPUT13), .Z(new_n416));
  INV_X1    g279(.A(new_n411), .ZN(RLL_wire_A_90));
  XOR2_X1 RLL_XOR_90 (.A(RLL_wire_A_90), .B(KEYINPUT90), .Z(new_n417) );
  NOR2_X1   g280(.A1(new_n410), .A2(new_n394), .ZN(new_n418));
  OAI21_X1  g281(.A(new_n416), .B1(new_n417), .B2(new_n418), .ZN(new_n419));
  NAND2_X1  g282(.A1(new_n415), .A2(new_n419), .ZN(new_n420));
  OAI21_X1  g283(.A(new_n373), .B1(new_n414), .B2(new_n420), .ZN(new_n421));
  NAND2_X1  g284(.A1(new_n412), .A2(new_n413), .ZN(new_n422));
  NAND4_X1  g285(.A1(new_n422), .A2(new_n419), .A3(new_n415), .A4(new_n372), .ZN(new_n423));
  AND2_X1   g286(.A1(new_n421), .A2(new_n423), .ZN(new_n424));
  NOR2_X1   g287(.A1(new_n367), .A2(new_n424), .ZN(new_n425));
  AND2_X1   g288(.A1(G71gat), .A2(G78gat), .ZN(new_n426));
  NOR2_X1   g289(.A1(G71gat), .A2(G78gat), .ZN(new_n427));
  NOR2_X1   g290(.A1(new_n426), .A2(new_n427), .ZN(new_n428));
  XNOR2_X1  g291(.A(G57gat), .B(G64gat), .ZN(new_n429));
  AOI21_X1  g292(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n430));
  OAI21_X1  g293(.A(new_n428), .B1(new_n429), .B2(new_n430), .ZN(new_n431));
  INV_X1    g294(.A(G57gat), .ZN(new_n432));
  NAND2_X1  g295(.A1(new_n432), .A2(G64gat), .ZN(new_n433));
  INV_X1    g296(.A(G64gat), .ZN(new_n434));
  NAND2_X1  g297(.A1(new_n434), .A2(G57gat), .ZN(new_n435));
  NAND2_X1  g298(.A1(new_n433), .A2(new_n435), .ZN(new_n436));
  XNOR2_X1  g299(.A(G71gat), .B(G78gat), .ZN(RLL_wire_A_91));
  XNOR2_X1 RLL_XNOR_91 (.A(RLL_wire_A_91), .B(KEYINPUT91), .ZN(new_n437) );
  INV_X1    g300(.A(new_n430), .ZN(new_n438));
  NAND3_X1  g301(.A1(new_n436), .A2(new_n437), .A3(new_n438), .ZN(new_n439));
  NAND2_X1  g302(.A1(new_n431), .A2(new_n439), .ZN(new_n440));
  INV_X1    g303(.A(KEYINPUT21), .ZN(new_n441));
  NAND2_X1  g304(.A1(new_n440), .A2(new_n441), .ZN(new_n442));
  NAND2_X1  g305(.A1(G231gat), .A2(G233gat), .ZN(new_n443));
  XNOR2_X1  g306(.A(new_n442), .B(new_n443), .ZN(new_n444));
  XNOR2_X1  g307(.A(G127gat), .B(G155gat), .ZN(new_n445));
  XNOR2_X1  g308(.A(new_n445), .B(KEYINPUT19), .ZN(new_n446));
  XOR2_X1   g309(.A(new_n446), .B(KEYINPUT20), .Z(new_n447));
  XNOR2_X1  g310(.A(new_n444), .B(new_n447), .ZN(new_n448));
  INV_X1    g311(.A(new_n440), .ZN(new_n449));
  AOI21_X1  g312(.A(new_n410), .B1(KEYINPUT21), .B2(new_n449), .ZN(new_n450));
  XNOR2_X1  g313(.A(G183gat), .B(G211gat), .ZN(new_n451));
  XNOR2_X1  g314(.A(new_n450), .B(new_n451), .ZN(new_n452));
  XOR2_X1   g315(.A(new_n448), .B(new_n452), .Z(new_n453));
  AND2_X1   g316(.A1(G232gat), .A2(G233gat), .ZN(RLL_wire_A_92));
  XNOR2_X1 RLL_XNOR_92 (.A(RLL_wire_A_92), .B(KEYINPUT92), .ZN(new_n454) );
  NOR2_X1   g317(.A1(new_n454), .A2(KEYINPUT41), .ZN(new_n455));
  XNOR2_X1  g318(.A(G134gat), .B(G162gat), .ZN(new_n456));
  XNOR2_X1  g319(.A(new_n455), .B(new_n456), .ZN(new_n457));
  INV_X1    g320(.A(new_n457), .ZN(new_n458));
  NAND2_X1  g321(.A1(G85gat), .A2(G92gat), .ZN(RLL_wire_A_93));
  XNOR2_X1 RLL_XNOR_93 (.A(RLL_wire_A_93), .B(KEYINPUT93), .ZN(new_n459) );
  NAND2_X1  g322(.A1(new_n459), .A2(KEYINPUT7), .ZN(new_n460));
  INV_X1    g323(.A(KEYINPUT7), .ZN(new_n461));
  NAND3_X1  g324(.A1(new_n461), .A2(G85gat), .A3(G92gat), .ZN(new_n462));
  NAND2_X1  g325(.A1(new_n460), .A2(new_n462), .ZN(new_n463));
  NAND2_X1  g326(.A1(G99gat), .A2(G106gat), .ZN(new_n464));
  INV_X1    g327(.A(G85gat), .ZN(new_n465));
  INV_X1    g328(.A(G92gat), .ZN(RLL_wire_A_94));
  XOR2_X1 RLL_XOR_94 (.A(RLL_wire_A_94), .B(KEYINPUT94), .Z(new_n466) );
  AOI22_X1  g329(.A1(KEYINPUT8), .A2(new_n464), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  XNOR2_X1  g330(.A(G99gat), .B(G106gat), .ZN(new_n468));
  NAND3_X1  g331(.A1(new_n463), .A2(new_n467), .A3(new_n468), .ZN(new_n469));
  INV_X1    g332(.A(new_n469), .ZN(new_n470));
  AOI21_X1  g333(.A(new_n468), .B1(new_n463), .B2(new_n467), .ZN(new_n471));
  NOR2_X1   g334(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  INV_X1    g335(.A(new_n472), .ZN(new_n473));
  NAND3_X1  g336(.A1(new_n396), .A2(new_n473), .A3(new_n407), .ZN(new_n474));
  AOI22_X1  g337(.A1(new_n394), .A2(new_n472), .B1(KEYINPUT41), .B2(new_n454), .ZN(new_n475));
  XNOR2_X1  g338(.A(G190gat), .B(G218gat), .ZN(new_n476));
  INV_X1    g339(.A(new_n476), .ZN(RLL_wire_A_95));
  XOR2_X1 RLL_XOR_95 (.A(RLL_wire_A_95), .B(KEYINPUT95), .Z(new_n477) );
  NAND3_X1  g340(.A1(new_n474), .A2(new_n475), .A3(new_n477), .ZN(new_n478));
  INV_X1    g341(.A(new_n478), .ZN(new_n479));
  AOI21_X1  g342(.A(new_n477), .B1(new_n474), .B2(new_n475), .ZN(RLL_wire_A_96));
  XNOR2_X1 RLL_XNOR_96 (.A(RLL_wire_A_96), .B(KEYINPUT96), .ZN(new_n480) );
  OAI21_X1  g343(.A(new_n458), .B1(new_n479), .B2(new_n480), .ZN(new_n481));
  INV_X1    g344(.A(new_n480), .ZN(new_n482));
  NAND3_X1  g345(.A1(new_n482), .A2(new_n457), .A3(new_n478), .ZN(RLL_wire_A_97));
  XOR2_X1 RLL_XOR_97 (.A(RLL_wire_A_97), .B(KEYINPUT97), .Z(new_n483) );
  AND2_X1   g346(.A1(new_n481), .A2(new_n483), .ZN(new_n484));
  NAND2_X1  g347(.A1(new_n453), .A2(new_n484), .ZN(new_n485));
  OAI21_X1  g348(.A(new_n440), .B1(new_n470), .B2(new_n471), .ZN(new_n486));
  NAND2_X1  g349(.A1(new_n463), .A2(new_n467), .ZN(RLL_wire_A_98));
  XNOR2_X1 RLL_XNOR_98 (.A(RLL_wire_A_98), .B(KEYINPUT98), .ZN(new_n487) );
  INV_X1    g350(.A(new_n468), .ZN(new_n488));
  NAND2_X1  g351(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  NAND4_X1  g352(.A1(new_n489), .A2(new_n469), .A3(new_n431), .A4(new_n439), .ZN(new_n490));
  INV_X1    g353(.A(KEYINPUT10), .ZN(new_n491));
  NAND3_X1  g354(.A1(new_n486), .A2(new_n490), .A3(new_n491), .ZN(new_n492));
  NAND3_X1  g355(.A1(new_n472), .A2(KEYINPUT10), .A3(new_n449), .ZN(new_n493));
  NAND2_X1  g356(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  NAND2_X1  g357(.A1(G230gat), .A2(G233gat), .ZN(new_n495));
  NAND2_X1  g358(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  AOI21_X1  g359(.A(new_n495), .B1(new_n486), .B2(new_n490), .ZN(new_n497));
  INV_X1    g360(.A(new_n497), .ZN(new_n498));
  XNOR2_X1  g361(.A(G120gat), .B(G148gat), .ZN(new_n499));
  XNOR2_X1  g362(.A(G176gat), .B(G204gat), .ZN(new_n500));
  XOR2_X1   g363(.A(new_n499), .B(new_n500), .Z(new_n501));
  NAND3_X1  g364(.A1(new_n496), .A2(new_n498), .A3(new_n501), .ZN(new_n502));
  INV_X1    g365(.A(new_n501), .ZN(new_n503));
  INV_X1    g366(.A(new_n495), .ZN(new_n504));
  AOI21_X1  g367(.A(new_n504), .B1(new_n492), .B2(new_n493), .ZN(new_n505));
  OAI21_X1  g368(.A(new_n503), .B1(new_n505), .B2(new_n497), .ZN(new_n506));
  NAND2_X1  g369(.A1(new_n502), .A2(new_n506), .ZN(new_n507));
  NOR2_X1   g370(.A1(new_n485), .A2(new_n507), .ZN(new_n508));
  AND2_X1   g371(.A1(new_n425), .A2(new_n508), .ZN(new_n509));
  NOR2_X1   g372(.A1(new_n304), .A2(new_n305), .ZN(new_n510));
  NAND2_X1  g373(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  XNOR2_X1  g374(.A(new_n511), .B(G1gat), .ZN(RLL_wire_A_99));
  XOR2_X1 RLL_XOR_99 (.A(RLL_wire_A_99), .B(KEYINPUT99), .Z(G1324gat) );
  INV_X1    g375(.A(KEYINPUT42), .ZN(new_n513));
  NAND2_X1  g376(.A1(new_n509), .A2(new_n334), .ZN(new_n514));
  XOR2_X1   g377(.A(KEYINPUT16), .B(G8gat), .Z(new_n515));
  INV_X1    g378(.A(new_n515), .ZN(new_n516));
  OAI21_X1  g379(.A(new_n513), .B1(new_n514), .B2(new_n516), .ZN(RLL_wire_A_100));
  XNOR2_X1 RLL_XNOR_100 (.A(RLL_wire_A_100), .B(KEYINPUT100), .ZN(new_n517) );
  NAND2_X1  g380(.A1(new_n514), .A2(G8gat), .ZN(new_n518));
  NAND4_X1  g381(.A1(new_n509), .A2(KEYINPUT42), .A3(new_n334), .A4(new_n515), .ZN(new_n519));
  NAND3_X1  g382(.A1(new_n517), .A2(new_n518), .A3(new_n519), .ZN(G1325gat));
  AOI21_X1  g383(.A(G15gat), .B1(new_n509), .B2(new_n362), .ZN(new_n521));
  NAND2_X1  g384(.A1(new_n222), .A2(new_n218), .ZN(new_n522));
  INV_X1    g385(.A(new_n522), .ZN(new_n523));
  AND2_X1   g386(.A1(new_n523), .A2(G15gat), .ZN(new_n524));
  AOI21_X1  g387(.A(new_n521), .B1(new_n509), .B2(new_n524), .ZN(G1326gat));
  NAND2_X1  g388(.A1(new_n509), .A2(new_n332), .ZN(RLL_wire_A_101));
  XNOR2_X1 RLL_XNOR_101 (.A(RLL_wire_A_101), .B(KEYINPUT101), .ZN(new_n526) );
  XNOR2_X1  g389(.A(KEYINPUT43), .B(G22gat), .ZN(new_n527));
  XNOR2_X1  g390(.A(new_n526), .B(new_n527), .ZN(G1327gat));
  NOR3_X1   g391(.A1(new_n453), .A2(new_n484), .A3(new_n507), .ZN(new_n529));
  NAND4_X1  g392(.A1(new_n425), .A2(new_n379), .A3(new_n510), .A4(new_n529), .ZN(new_n530));
  XNOR2_X1  g393(.A(new_n530), .B(KEYINPUT45), .ZN(new_n531));
  NAND2_X1  g394(.A1(new_n421), .A2(new_n423), .ZN(new_n532));
  INV_X1    g395(.A(new_n453), .ZN(new_n533));
  INV_X1    g396(.A(new_n507), .ZN(new_n534));
  NAND3_X1  g397(.A1(new_n532), .A2(new_n533), .A3(new_n534), .ZN(new_n535));
  OAI21_X1  g398(.A(KEYINPUT44), .B1(new_n367), .B2(new_n484), .ZN(new_n536));
  NAND2_X1  g399(.A1(new_n306), .A2(new_n332), .ZN(new_n537));
  NAND3_X1  g400(.A1(new_n360), .A2(new_n537), .A3(new_n522), .ZN(RLL_wire_A_102));
  XNOR2_X1 RLL_XNOR_102 (.A(RLL_wire_A_102), .B(KEYINPUT102), .ZN(new_n538) );
  NAND2_X1  g401(.A1(new_n364), .A2(new_n366), .ZN(new_n539));
  NAND2_X1  g402(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  INV_X1    g403(.A(KEYINPUT44), .ZN(new_n541));
  INV_X1    g404(.A(new_n484), .ZN(new_n542));
  NAND3_X1  g405(.A1(new_n540), .A2(new_n541), .A3(new_n542), .ZN(new_n543));
  AOI21_X1  g406(.A(new_n535), .B1(new_n536), .B2(new_n543), .ZN(new_n544));
  AND2_X1   g407(.A1(new_n544), .A2(new_n510), .ZN(new_n545));
  OAI21_X1  g408(.A(new_n531), .B1(new_n545), .B2(new_n379), .ZN(G1328gat));
  NAND4_X1  g409(.A1(new_n425), .A2(new_n380), .A3(new_n334), .A4(new_n529), .ZN(new_n547));
  NAND2_X1  g410(.A1(new_n547), .A2(KEYINPUT46), .ZN(new_n548));
  OR2_X1    g411(.A1(new_n547), .A2(KEYINPUT46), .ZN(new_n549));
  AND2_X1   g412(.A1(new_n544), .A2(new_n334), .ZN(new_n550));
  OAI211_X1 g413(.A(new_n548), .B(new_n549), .C1(new_n550), .C2(new_n380), .ZN(G1329gat));
  INV_X1    g414(.A(KEYINPUT47), .ZN(RLL_wire_A_103));
  XOR2_X1 RLL_XOR_103 (.A(RLL_wire_A_103), .B(KEYINPUT103), .Z(new_n552) );
  AOI21_X1  g415(.A(new_n385), .B1(new_n544), .B2(new_n523), .ZN(new_n553));
  NAND4_X1  g416(.A1(new_n425), .A2(new_n385), .A3(new_n362), .A4(new_n529), .ZN(new_n554));
  INV_X1    g417(.A(new_n554), .ZN(new_n555));
  OAI21_X1  g418(.A(new_n552), .B1(new_n553), .B2(new_n555), .ZN(new_n556));
  AOI211_X1 g419(.A(new_n522), .B(new_n535), .C1(new_n536), .C2(new_n543), .ZN(new_n557));
  OAI211_X1 g420(.A(KEYINPUT47), .B(new_n554), .C1(new_n557), .C2(new_n385), .ZN(new_n558));
  NAND2_X1  g421(.A1(new_n556), .A2(new_n558), .ZN(RLL_wire_A_104));
  XNOR2_X1 RLL_XNOR_104 (.A(RLL_wire_A_104), .B(KEYINPUT104), .ZN(G1330gat) );
  INV_X1    g422(.A(KEYINPUT48), .ZN(new_n560));
  AOI21_X1  g423(.A(new_n387), .B1(new_n544), .B2(new_n332), .ZN(new_n561));
  NAND2_X1  g424(.A1(new_n425), .A2(new_n529), .ZN(new_n562));
  NAND2_X1  g425(.A1(new_n332), .A2(new_n387), .ZN(new_n563));
  NOR2_X1   g426(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  OAI21_X1  g427(.A(new_n560), .B1(new_n561), .B2(new_n564), .ZN(new_n565));
  OR2_X1    g428(.A1(new_n562), .A2(new_n563), .ZN(RLL_wire_A_105));
  XNOR2_X1 RLL_XNOR_105 (.A(RLL_wire_A_105), .B(KEYINPUT105), .ZN(new_n566) );
  AOI211_X1 g429(.A(new_n331), .B(new_n535), .C1(new_n536), .C2(new_n543), .ZN(RLL_wire_A_106));
  XNOR2_X1 RLL_XNOR_106 (.A(RLL_wire_A_106), .B(KEYINPUT106), .ZN(new_n567) );
  OAI211_X1 g430(.A(new_n566), .B(KEYINPUT48), .C1(new_n567), .C2(new_n387), .ZN(new_n568));
  NAND2_X1  g431(.A1(new_n565), .A2(new_n568), .ZN(G1331gat));
  NOR3_X1   g432(.A1(new_n485), .A2(new_n532), .A3(new_n534), .ZN(new_n570));
  NAND2_X1  g433(.A1(new_n540), .A2(new_n570), .ZN(new_n571));
  INV_X1    g434(.A(new_n510), .ZN(new_n572));
  NOR2_X1   g435(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  XNOR2_X1  g436(.A(new_n573), .B(new_n432), .ZN(G1332gat));
  INV_X1    g437(.A(new_n571), .ZN(new_n575));
  INV_X1    g438(.A(new_n334), .ZN(new_n576));
  AOI21_X1  g439(.A(new_n576), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n577));
  NAND2_X1  g440(.A1(new_n575), .A2(new_n577), .ZN(new_n578));
  NOR2_X1   g441(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n579));
  XOR2_X1   g442(.A(new_n578), .B(new_n579), .Z(G1333gat));
  NAND3_X1  g443(.A1(new_n575), .A2(G71gat), .A3(new_n523), .ZN(new_n581));
  INV_X1    g444(.A(new_n362), .ZN(new_n582));
  NOR2_X1   g445(.A1(new_n571), .A2(new_n582), .ZN(new_n583));
  OAI21_X1  g446(.A(new_n581), .B1(G71gat), .B2(new_n583), .ZN(new_n584));
  XNOR2_X1  g447(.A(new_n584), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g448(.A1(new_n575), .A2(new_n332), .ZN(new_n586));
  XNOR2_X1  g449(.A(new_n586), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g450(.A1(new_n453), .A2(new_n532), .ZN(new_n588));
  NAND2_X1  g451(.A1(new_n588), .A2(new_n507), .ZN(new_n589));
  AOI21_X1  g452(.A(new_n589), .B1(new_n536), .B2(new_n543), .ZN(new_n590));
  AND2_X1   g453(.A1(new_n590), .A2(new_n510), .ZN(new_n591));
  AOI21_X1  g454(.A(new_n484), .B1(new_n538), .B2(new_n539), .ZN(new_n592));
  NAND3_X1  g455(.A1(new_n592), .A2(KEYINPUT51), .A3(new_n588), .ZN(new_n593));
  INV_X1    g456(.A(new_n593), .ZN(new_n594));
  AOI21_X1  g457(.A(KEYINPUT51), .B1(new_n592), .B2(new_n588), .ZN(new_n595));
  NOR2_X1   g458(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  NAND3_X1  g459(.A1(new_n510), .A2(new_n465), .A3(new_n507), .ZN(RLL_wire_A_107));
  XNOR2_X1 RLL_XNOR_107 (.A(RLL_wire_A_107), .B(KEYINPUT107), .ZN(new_n597) );
  OAI22_X1  g460(.A1(new_n591), .A2(new_n465), .B1(new_n596), .B2(new_n597), .ZN(G1336gat));
  AOI21_X1  g461(.A(new_n466), .B1(new_n590), .B2(new_n334), .ZN(new_n599));
  NOR3_X1   g462(.A1(new_n576), .A2(G92gat), .A3(new_n534), .ZN(new_n600));
  INV_X1    g463(.A(new_n600), .ZN(new_n601));
  NAND2_X1  g464(.A1(new_n592), .A2(new_n588), .ZN(new_n602));
  INV_X1    g465(.A(KEYINPUT51), .ZN(new_n603));
  NAND2_X1  g466(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  AOI21_X1  g467(.A(new_n601), .B1(new_n604), .B2(new_n593), .ZN(RLL_wire_A_108));
  XNOR2_X1 RLL_XNOR_108 (.A(RLL_wire_A_108), .B(KEYINPUT108), .ZN(new_n605) );
  OAI21_X1  g468(.A(KEYINPUT52), .B1(new_n599), .B2(new_n605), .ZN(new_n606));
  OAI21_X1  g469(.A(new_n600), .B1(new_n594), .B2(new_n595), .ZN(RLL_wire_A_109));
  XNOR2_X1 RLL_XNOR_109 (.A(RLL_wire_A_109), .B(KEYINPUT109), .ZN(new_n607) );
  INV_X1    g470(.A(KEYINPUT52), .ZN(new_n608));
  AOI211_X1 g471(.A(new_n576), .B(new_n589), .C1(new_n536), .C2(new_n543), .ZN(new_n609));
  OAI211_X1 g472(.A(new_n607), .B(new_n608), .C1(new_n609), .C2(new_n466), .ZN(new_n610));
  NAND2_X1  g473(.A1(new_n606), .A2(new_n610), .ZN(G1337gat));
  AND2_X1   g474(.A1(new_n590), .A2(new_n523), .ZN(new_n612));
  INV_X1    g475(.A(G99gat), .ZN(new_n613));
  NAND3_X1  g476(.A1(new_n362), .A2(new_n613), .A3(new_n507), .ZN(new_n614));
  OAI22_X1  g477(.A1(new_n612), .A2(new_n613), .B1(new_n596), .B2(new_n614), .ZN(G1338gat));
  INV_X1    g478(.A(G106gat), .ZN(new_n616));
  AOI21_X1  g479(.A(new_n616), .B1(new_n590), .B2(new_n332), .ZN(RLL_wire_A_110));
  XNOR2_X1 RLL_XNOR_110 (.A(RLL_wire_A_110), .B(KEYINPUT110), .ZN(new_n617) );
  NOR3_X1   g480(.A1(new_n331), .A2(G106gat), .A3(new_n534), .ZN(new_n618));
  INV_X1    g481(.A(new_n618), .ZN(new_n619));
  AOI21_X1  g482(.A(new_n619), .B1(new_n604), .B2(new_n593), .ZN(new_n620));
  OAI21_X1  g483(.A(KEYINPUT53), .B1(new_n617), .B2(new_n620), .ZN(new_n621));
  OAI21_X1  g484(.A(new_n618), .B1(new_n594), .B2(new_n595), .ZN(new_n622));
  INV_X1    g485(.A(KEYINPUT53), .ZN(new_n623));
  AOI211_X1 g486(.A(new_n331), .B(new_n589), .C1(new_n536), .C2(new_n543), .ZN(new_n624));
  OAI211_X1 g487(.A(new_n622), .B(new_n623), .C1(new_n624), .C2(new_n616), .ZN(new_n625));
  NAND2_X1  g488(.A1(new_n621), .A2(new_n625), .ZN(G1339gat));
  NOR3_X1   g489(.A1(new_n485), .A2(new_n532), .A3(new_n507), .ZN(new_n627));
  NAND3_X1  g490(.A1(new_n492), .A2(new_n504), .A3(new_n493), .ZN(new_n628));
  NAND3_X1  g491(.A1(new_n496), .A2(KEYINPUT54), .A3(new_n628), .ZN(new_n629));
  INV_X1    g492(.A(KEYINPUT54), .ZN(new_n630));
  AOI21_X1  g493(.A(new_n501), .B1(new_n505), .B2(new_n630), .ZN(new_n631));
  NAND3_X1  g494(.A1(new_n629), .A2(KEYINPUT55), .A3(new_n631), .ZN(new_n632));
  NAND2_X1  g495(.A1(new_n632), .A2(new_n502), .ZN(new_n633));
  AOI21_X1  g496(.A(KEYINPUT55), .B1(new_n629), .B2(new_n631), .ZN(RLL_wire_A_111));
  XNOR2_X1 RLL_XNOR_111 (.A(RLL_wire_A_111), .B(KEYINPUT111), .ZN(new_n634) );
  NOR2_X1   g497(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  AOI21_X1  g498(.A(new_n409), .B1(new_n408), .B2(new_n411), .ZN(RLL_wire_A_112));
  XOR2_X1 RLL_XOR_112 (.A(RLL_wire_A_112), .B(KEYINPUT112), .Z(new_n636) );
  NOR3_X1   g499(.A1(new_n417), .A2(new_n418), .A3(new_n416), .ZN(new_n637));
  OAI21_X1  g500(.A(new_n371), .B1(new_n636), .B2(new_n637), .ZN(new_n638));
  AND2_X1   g501(.A1(new_n423), .A2(new_n638), .ZN(new_n639));
  NAND3_X1  g502(.A1(new_n635), .A2(new_n542), .A3(new_n639), .ZN(new_n640));
  AND3_X1   g503(.A1(new_n423), .A2(new_n507), .A3(new_n638), .ZN(new_n641));
  AOI21_X1  g504(.A(new_n641), .B1(new_n635), .B2(new_n532), .ZN(new_n642));
  OAI21_X1  g505(.A(new_n640), .B1(new_n642), .B2(new_n542), .ZN(new_n643));
  AOI21_X1  g506(.A(new_n627), .B1(new_n643), .B2(new_n533), .ZN(RLL_wire_A_113));
  XOR2_X1 RLL_XOR_113 (.A(RLL_wire_A_113), .B(KEYINPUT113), .Z(new_n644) );
  NOR2_X1   g507(.A1(new_n644), .A2(new_n332), .ZN(new_n645));
  NAND4_X1  g508(.A1(new_n645), .A2(new_n510), .A3(new_n576), .A4(new_n362), .ZN(new_n646));
  OAI21_X1  g509(.A(G113gat), .B1(new_n646), .B2(new_n424), .ZN(new_n647));
  NOR3_X1   g510(.A1(new_n644), .A2(new_n572), .A3(new_n365), .ZN(new_n648));
  NAND2_X1  g511(.A1(new_n648), .A2(new_n576), .ZN(new_n649));
  NAND2_X1  g512(.A1(new_n532), .A2(new_n190), .ZN(new_n650));
  OAI21_X1  g513(.A(new_n647), .B1(new_n649), .B2(new_n650), .ZN(G1340gat));
  OAI21_X1  g514(.A(G120gat), .B1(new_n646), .B2(new_n534), .ZN(new_n652));
  NAND2_X1  g515(.A1(new_n507), .A2(new_n188), .ZN(new_n653));
  OAI21_X1  g516(.A(new_n652), .B1(new_n649), .B2(new_n653), .ZN(G1341gat));
  NOR3_X1   g517(.A1(new_n646), .A2(new_n183), .A3(new_n533), .ZN(new_n655));
  NAND3_X1  g518(.A1(new_n648), .A2(new_n576), .A3(new_n453), .ZN(new_n656));
  AOI21_X1  g519(.A(new_n655), .B1(new_n183), .B2(new_n656), .ZN(G1342gat));
  NOR2_X1   g520(.A1(new_n484), .A2(new_n334), .ZN(new_n658));
  NAND3_X1  g521(.A1(new_n648), .A2(new_n181), .A3(new_n658), .ZN(new_n659));
  OR2_X1    g522(.A1(new_n659), .A2(KEYINPUT56), .ZN(new_n660));
  OAI21_X1  g523(.A(G134gat), .B1(new_n646), .B2(new_n484), .ZN(new_n661));
  NAND2_X1  g524(.A1(new_n659), .A2(KEYINPUT56), .ZN(new_n662));
  NAND3_X1  g525(.A1(new_n660), .A2(new_n661), .A3(new_n662), .ZN(RLL_wire_A_114));
  XNOR2_X1 RLL_XNOR_114 (.A(RLL_wire_A_114), .B(KEYINPUT114), .ZN(G1343gat) );
  NAND3_X1  g526(.A1(new_n522), .A2(new_n510), .A3(new_n576), .ZN(new_n664));
  INV_X1    g527(.A(KEYINPUT57), .ZN(new_n665));
  OAI21_X1  g528(.A(new_n665), .B1(new_n644), .B2(new_n331), .ZN(new_n666));
  NAND3_X1  g529(.A1(new_n423), .A2(new_n507), .A3(new_n638), .ZN(RLL_wire_A_115));
  XNOR2_X1 RLL_XNOR_115 (.A(RLL_wire_A_115), .B(KEYINPUT115), .ZN(new_n667) );
  NAND2_X1  g530(.A1(new_n629), .A2(new_n631), .ZN(new_n668));
  INV_X1    g531(.A(KEYINPUT55), .ZN(new_n669));
  NAND2_X1  g532(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  NAND3_X1  g533(.A1(new_n670), .A2(new_n502), .A3(new_n632), .ZN(new_n671));
  OAI21_X1  g534(.A(new_n667), .B1(new_n424), .B2(new_n671), .ZN(new_n672));
  NAND2_X1  g535(.A1(new_n672), .A2(new_n484), .ZN(new_n673));
  AOI21_X1  g536(.A(new_n453), .B1(new_n673), .B2(new_n640), .ZN(RLL_wire_A_116));
  XOR2_X1 RLL_XOR_116 (.A(RLL_wire_A_116), .B(KEYINPUT116), .Z(new_n674) );
  OAI211_X1 g537(.A(KEYINPUT57), .B(new_n332), .C1(new_n674), .C2(new_n627), .ZN(new_n675));
  AOI21_X1  g538(.A(new_n664), .B1(new_n666), .B2(new_n675), .ZN(new_n676));
  AOI21_X1  g539(.A(new_n264), .B1(new_n676), .B2(new_n532), .ZN(RLL_wire_A_117));
  XNOR2_X1 RLL_XNOR_117 (.A(RLL_wire_A_117), .B(KEYINPUT117), .ZN(new_n677) );
  NOR2_X1   g540(.A1(new_n644), .A2(new_n572), .ZN(new_n678));
  NOR2_X1   g541(.A1(new_n523), .A2(new_n331), .ZN(new_n679));
  NOR2_X1   g542(.A1(new_n424), .A2(G141gat), .ZN(RLL_wire_A_118));
  XOR2_X1 RLL_XOR_118 (.A(RLL_wire_A_118), .B(KEYINPUT118), .Z(new_n680) );
  AND4_X1   g543(.A1(new_n576), .A2(new_n678), .A3(new_n679), .A4(new_n680), .ZN(RLL_wire_A_119));
  XNOR2_X1 RLL_XNOR_119 (.A(RLL_wire_A_119), .B(KEYINPUT119), .ZN(new_n681) );
  OAI21_X1  g544(.A(KEYINPUT58), .B1(new_n677), .B2(new_n681), .ZN(new_n682));
  AND2_X1   g545(.A1(new_n678), .A2(new_n679), .ZN(new_n683));
  NAND3_X1  g546(.A1(new_n683), .A2(new_n576), .A3(new_n680), .ZN(new_n684));
  INV_X1    g547(.A(KEYINPUT58), .ZN(new_n685));
  AOI211_X1 g548(.A(new_n424), .B(new_n664), .C1(new_n666), .C2(new_n675), .ZN(new_n686));
  OAI211_X1 g549(.A(new_n684), .B(new_n685), .C1(new_n686), .C2(new_n264), .ZN(new_n687));
  NAND2_X1  g550(.A1(new_n682), .A2(new_n687), .ZN(G1344gat));
  NAND4_X1  g551(.A1(new_n683), .A2(new_n266), .A3(new_n576), .A4(new_n507), .ZN(new_n689));
  AOI211_X1 g552(.A(KEYINPUT59), .B(new_n266), .C1(new_n676), .C2(new_n507), .ZN(new_n690));
  INV_X1    g553(.A(KEYINPUT59), .ZN(new_n691));
  INV_X1    g554(.A(new_n664), .ZN(new_n692));
  NOR3_X1   g555(.A1(new_n644), .A2(new_n665), .A3(new_n331), .ZN(new_n693));
  NAND2_X1  g556(.A1(new_n508), .A2(new_n424), .ZN(RLL_wire_A_120));
  XNOR2_X1 RLL_XNOR_120 (.A(RLL_wire_A_120), .B(KEYINPUT120), .ZN(new_n694) );
  NOR3_X1   g557(.A1(new_n484), .A2(new_n633), .A3(new_n634), .ZN(new_n695));
  AOI22_X1  g558(.A1(new_n672), .A2(new_n484), .B1(new_n639), .B2(new_n695), .ZN(new_n696));
  OAI21_X1  g559(.A(new_n694), .B1(new_n696), .B2(new_n453), .ZN(new_n697));
  AOI21_X1  g560(.A(KEYINPUT57), .B1(new_n697), .B2(new_n332), .ZN(new_n698));
  OAI211_X1 g561(.A(new_n507), .B(new_n692), .C1(new_n693), .C2(new_n698), .ZN(new_n699));
  AOI21_X1  g562(.A(new_n691), .B1(new_n699), .B2(G148gat), .ZN(RLL_wire_A_121));
  XNOR2_X1 RLL_XNOR_121 (.A(RLL_wire_A_121), .B(KEYINPUT121), .ZN(new_n700) );
  OAI21_X1  g563(.A(new_n689), .B1(new_n690), .B2(new_n700), .ZN(G1345gat));
  NAND3_X1  g564(.A1(new_n683), .A2(new_n576), .A3(new_n453), .ZN(new_n702));
  NOR2_X1   g565(.A1(new_n533), .A2(new_n270), .ZN(RLL_wire_A_122));
  XNOR2_X1 RLL_XNOR_122 (.A(RLL_wire_A_122), .B(KEYINPUT122), .ZN(new_n703) );
  AOI22_X1  g566(.A1(new_n702), .A2(new_n270), .B1(new_n676), .B2(new_n703), .ZN(G1346gat));
  NAND3_X1  g567(.A1(new_n683), .A2(new_n271), .A3(new_n658), .ZN(new_n705));
  AND2_X1   g568(.A1(new_n676), .A2(new_n542), .ZN(new_n706));
  OAI21_X1  g569(.A(new_n705), .B1(new_n706), .B2(new_n271), .ZN(G1347gat));
  NOR2_X1   g570(.A1(new_n644), .A2(new_n510), .ZN(new_n708));
  NOR2_X1   g571(.A1(new_n365), .A2(new_n576), .ZN(new_n709));
  AND2_X1   g572(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  NAND3_X1  g573(.A1(new_n710), .A2(new_n145), .A3(new_n532), .ZN(new_n711));
  NAND2_X1  g574(.A1(new_n572), .A2(new_n334), .ZN(new_n712));
  NOR2_X1   g575(.A1(new_n712), .A2(new_n582), .ZN(new_n713));
  NAND2_X1  g576(.A1(new_n645), .A2(new_n713), .ZN(new_n714));
  OAI21_X1  g577(.A(G169gat), .B1(new_n714), .B2(new_n424), .ZN(new_n715));
  NAND2_X1  g578(.A1(new_n711), .A2(new_n715), .ZN(G1348gat));
  AOI21_X1  g579(.A(G176gat), .B1(new_n710), .B2(new_n507), .ZN(new_n717));
  NOR3_X1   g580(.A1(new_n714), .A2(new_n146), .A3(new_n534), .ZN(new_n718));
  NOR2_X1   g581(.A1(new_n717), .A2(new_n718), .ZN(G1349gat));
  NAND4_X1  g582(.A1(new_n708), .A2(new_n172), .A3(new_n453), .A4(new_n709), .ZN(new_n720));
  NOR2_X1   g583(.A1(new_n714), .A2(new_n533), .ZN(new_n721));
  OAI21_X1  g584(.A(new_n720), .B1(new_n721), .B2(new_n160), .ZN(new_n722));
  NAND2_X1  g585(.A1(new_n722), .A2(KEYINPUT60), .ZN(new_n723));
  INV_X1    g586(.A(KEYINPUT60), .ZN(new_n724));
  OAI211_X1 g587(.A(new_n724), .B(new_n720), .C1(new_n721), .C2(new_n160), .ZN(new_n725));
  NAND2_X1  g588(.A1(new_n723), .A2(new_n725), .ZN(RLL_wire_A_123));
  XOR2_X1 RLL_XOR_123 (.A(RLL_wire_A_123), .B(KEYINPUT123), .Z(G1350gat) );
  NAND3_X1  g589(.A1(new_n710), .A2(new_n161), .A3(new_n542), .ZN(new_n727));
  OAI21_X1  g590(.A(G190gat), .B1(new_n714), .B2(new_n484), .ZN(RLL_wire_A_124));
  XOR2_X1 RLL_XOR_124 (.A(RLL_wire_A_124), .B(KEYINPUT124), .Z(new_n728) );
  AND2_X1   g591(.A1(new_n728), .A2(KEYINPUT61), .ZN(new_n729));
  NOR2_X1   g592(.A1(new_n728), .A2(KEYINPUT61), .ZN(new_n730));
  OAI21_X1  g593(.A(new_n727), .B1(new_n729), .B2(new_n730), .ZN(G1351gat));
  NOR3_X1   g594(.A1(new_n523), .A2(new_n331), .A3(new_n576), .ZN(new_n732));
  AND2_X1   g595(.A1(new_n708), .A2(new_n732), .ZN(new_n733));
  INV_X1    g596(.A(G197gat), .ZN(new_n734));
  NAND3_X1  g597(.A1(new_n733), .A2(new_n734), .A3(new_n532), .ZN(new_n735));
  NOR2_X1   g598(.A1(new_n693), .A2(new_n698), .ZN(new_n736));
  NOR2_X1   g599(.A1(new_n523), .A2(new_n712), .ZN(new_n737));
  INV_X1    g600(.A(new_n737), .ZN(new_n738));
  NOR3_X1   g601(.A1(new_n736), .A2(new_n424), .A3(new_n738), .ZN(new_n739));
  OAI21_X1  g602(.A(new_n735), .B1(new_n739), .B2(new_n734), .ZN(G1352gat));
  INV_X1    g603(.A(G204gat), .ZN(new_n741));
  NAND4_X1  g604(.A1(new_n708), .A2(new_n741), .A3(new_n507), .A4(new_n732), .ZN(new_n742));
  NAND2_X1  g605(.A1(new_n742), .A2(KEYINPUT62), .ZN(new_n743));
  OR2_X1    g606(.A1(new_n742), .A2(KEYINPUT62), .ZN(new_n744));
  NOR3_X1   g607(.A1(new_n736), .A2(new_n534), .A3(new_n738), .ZN(new_n745));
  OAI211_X1 g608(.A(new_n743), .B(new_n744), .C1(new_n745), .C2(new_n741), .ZN(G1353gat));
  NAND3_X1  g609(.A1(new_n733), .A2(new_n225), .A3(new_n453), .ZN(new_n747));
  OAI211_X1 g610(.A(new_n453), .B(new_n737), .C1(new_n693), .C2(new_n698), .ZN(RLL_wire_A_125));
  XNOR2_X1 RLL_XNOR_125 (.A(RLL_wire_A_125), .B(KEYINPUT125), .ZN(new_n748) );
  AND3_X1   g611(.A1(new_n748), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n749));
  AOI21_X1  g612(.A(KEYINPUT63), .B1(new_n748), .B2(G211gat), .ZN(new_n750));
  OAI21_X1  g613(.A(new_n747), .B1(new_n749), .B2(new_n750), .ZN(G1354gat));
  AOI21_X1  g614(.A(G218gat), .B1(new_n733), .B2(new_n542), .ZN(new_n752));
  NOR2_X1   g615(.A1(new_n736), .A2(new_n738), .ZN(new_n753));
  NOR2_X1   g616(.A1(new_n484), .A2(new_n226), .ZN(RLL_wire_A_126));
  XOR2_X1 RLL_XOR_126 (.A(RLL_wire_A_126), .B(KEYINPUT126), .Z(new_n754) );
  AOI21_X1  g617(.A(new_n752), .B1(new_n753), .B2(new_n754), .ZN(RLL_wire_A_127));
  XOR2_X1 RLL_XOR_127 (.A(RLL_wire_A_127), .B(KEYINPUT127), .Z(G1355gat) );

endmodule
