//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 0 0 1 1 1 0 0 0 1 1 0 0 1 0 1 1 0 0 0 0 1 1 1 1 1 0 1 1 1 1 0 1 0 0 0 1 1 0 0 1 1 0 0 0 0 1 1 0 0 1 0 0 0 0 1 0 1 1 1 1 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:32:24 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n437, new_n448, new_n452, new_n453, new_n454, new_n455,
    new_n456, new_n459, new_n460, new_n461, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n496,
    new_n497, new_n498, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n521, new_n522, new_n523, new_n524, new_n525, new_n526,
    new_n529, new_n530, new_n531, new_n532, new_n533, new_n534, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n550, new_n551, new_n552, new_n554,
    new_n555, new_n556, new_n557, new_n558, new_n559, new_n560, new_n561,
    new_n562, new_n563, new_n565, new_n566, new_n567, new_n569, new_n570,
    new_n571, new_n572, new_n573, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n605, new_n606, new_n607, new_n608, new_n611,
    new_n613, new_n614, new_n615, new_n616, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n837, new_n838, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1195, new_n1196;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(new_n436));
  INV_X1    g011(.A(KEYINPUT64), .ZN(new_n437));
  XNOR2_X1  g012(.A(new_n436), .B(new_n437), .ZN(G220));
  INV_X1    g013(.A(G96), .ZN(G221));
  INV_X1    g014(.A(G69), .ZN(G235));
  INV_X1    g015(.A(G120), .ZN(G236));
  INV_X1    g016(.A(G57), .ZN(G237));
  INV_X1    g017(.A(G108), .ZN(G238));
  NAND4_X1  g018(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g019(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g020(.A(G452), .Z(G391));
  AND2_X1   g021(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XOR2_X1   g023(.A(new_n448), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g024(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g025(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g026(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n452));
  XOR2_X1   g027(.A(KEYINPUT65), .B(KEYINPUT2), .Z(new_n453));
  XNOR2_X1  g028(.A(new_n452), .B(new_n453), .ZN(new_n454));
  NOR4_X1   g029(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n455));
  INV_X1    g030(.A(new_n455), .ZN(new_n456));
  NOR2_X1   g031(.A1(new_n454), .A2(new_n456), .ZN(G325));
  INV_X1    g032(.A(G325), .ZN(G261));
  NAND2_X1  g033(.A1(new_n454), .A2(G2106), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n456), .A2(G567), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  INV_X1    g036(.A(new_n461), .ZN(G319));
  XNOR2_X1  g037(.A(KEYINPUT3), .B(G2104), .ZN(new_n463));
  INV_X1    g038(.A(G2105), .ZN(new_n464));
  AND2_X1   g039(.A1(new_n464), .A2(G137), .ZN(new_n465));
  AND2_X1   g040(.A1(new_n464), .A2(G2104), .ZN(new_n466));
  AOI22_X1  g041(.A1(new_n463), .A2(new_n465), .B1(new_n466), .B2(G101), .ZN(new_n467));
  AOI22_X1  g042(.A1(new_n463), .A2(G125), .B1(G113), .B2(G2104), .ZN(new_n468));
  OAI21_X1  g043(.A(new_n467), .B1(new_n468), .B2(new_n464), .ZN(new_n469));
  INV_X1    g044(.A(new_n469), .ZN(G160));
  XNOR2_X1  g045(.A(new_n463), .B(KEYINPUT66), .ZN(new_n471));
  NOR2_X1   g046(.A1(new_n471), .A2(new_n464), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n472), .A2(G124), .ZN(new_n473));
  OR2_X1    g048(.A1(G100), .A2(G2105), .ZN(new_n474));
  OAI211_X1 g049(.A(new_n474), .B(G2104), .C1(G112), .C2(new_n464), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n473), .A2(new_n475), .ZN(new_n476));
  NOR2_X1   g051(.A1(new_n471), .A2(G2105), .ZN(new_n477));
  AOI21_X1  g052(.A(new_n476), .B1(G136), .B2(new_n477), .ZN(G162));
  OAI21_X1  g053(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n479));
  INV_X1    g054(.A(new_n479), .ZN(new_n480));
  INV_X1    g055(.A(G114), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n481), .A2(G2105), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n480), .A2(new_n482), .ZN(new_n483));
  AND2_X1   g058(.A1(G126), .A2(G2105), .ZN(new_n484));
  AND2_X1   g059(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n485));
  NOR2_X1   g060(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n486));
  OAI21_X1  g061(.A(new_n484), .B1(new_n485), .B2(new_n486), .ZN(new_n487));
  NAND2_X1  g062(.A1(new_n483), .A2(new_n487), .ZN(new_n488));
  INV_X1    g063(.A(G138), .ZN(new_n489));
  NOR2_X1   g064(.A1(new_n489), .A2(G2105), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n463), .A2(new_n490), .ZN(new_n491));
  NAND2_X1  g066(.A1(new_n491), .A2(KEYINPUT4), .ZN(new_n492));
  INV_X1    g067(.A(KEYINPUT4), .ZN(new_n493));
  OAI211_X1 g068(.A(new_n490), .B(new_n493), .C1(new_n486), .C2(new_n485), .ZN(new_n494));
  AOI21_X1  g069(.A(new_n488), .B1(new_n492), .B2(new_n494), .ZN(G164));
  INV_X1    g070(.A(KEYINPUT67), .ZN(new_n496));
  INV_X1    g071(.A(G543), .ZN(new_n497));
  OAI21_X1  g072(.A(new_n496), .B1(new_n497), .B2(KEYINPUT5), .ZN(new_n498));
  INV_X1    g073(.A(KEYINPUT5), .ZN(new_n499));
  NAND3_X1  g074(.A1(new_n499), .A2(KEYINPUT67), .A3(G543), .ZN(new_n500));
  NAND2_X1  g075(.A1(new_n498), .A2(new_n500), .ZN(new_n501));
  NAND2_X1  g076(.A1(new_n497), .A2(KEYINPUT5), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  AND2_X1   g078(.A1(KEYINPUT6), .A2(G651), .ZN(new_n504));
  NOR2_X1   g079(.A1(KEYINPUT6), .A2(G651), .ZN(new_n505));
  NOR2_X1   g080(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  OAI21_X1  g081(.A(KEYINPUT68), .B1(new_n503), .B2(new_n506), .ZN(new_n507));
  AOI22_X1  g082(.A1(new_n498), .A2(new_n500), .B1(KEYINPUT5), .B2(new_n497), .ZN(new_n508));
  INV_X1    g083(.A(KEYINPUT68), .ZN(new_n509));
  OAI211_X1 g084(.A(new_n508), .B(new_n509), .C1(new_n505), .C2(new_n504), .ZN(new_n510));
  AND2_X1   g085(.A1(new_n507), .A2(new_n510), .ZN(new_n511));
  XNOR2_X1  g086(.A(KEYINPUT69), .B(G88), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  NAND2_X1  g088(.A1(G75), .A2(G543), .ZN(new_n514));
  INV_X1    g089(.A(G62), .ZN(new_n515));
  OAI21_X1  g090(.A(new_n514), .B1(new_n503), .B2(new_n515), .ZN(new_n516));
  NOR2_X1   g091(.A1(new_n506), .A2(new_n497), .ZN(new_n517));
  AOI22_X1  g092(.A1(new_n516), .A2(G651), .B1(G50), .B2(new_n517), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n513), .A2(new_n518), .ZN(G303));
  INV_X1    g094(.A(G303), .ZN(G166));
  NAND3_X1  g095(.A1(new_n508), .A2(G63), .A3(G651), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n517), .A2(G51), .ZN(new_n522));
  NAND3_X1  g097(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n523));
  XNOR2_X1  g098(.A(new_n523), .B(KEYINPUT7), .ZN(new_n524));
  AND3_X1   g099(.A1(new_n521), .A2(new_n522), .A3(new_n524), .ZN(new_n525));
  NAND3_X1  g100(.A1(new_n507), .A2(new_n510), .A3(G89), .ZN(new_n526));
  NAND2_X1  g101(.A1(new_n525), .A2(new_n526), .ZN(G286));
  INV_X1    g102(.A(G286), .ZN(G168));
  NAND2_X1  g103(.A1(G77), .A2(G543), .ZN(new_n529));
  INV_X1    g104(.A(G64), .ZN(new_n530));
  OAI21_X1  g105(.A(new_n529), .B1(new_n503), .B2(new_n530), .ZN(new_n531));
  AOI22_X1  g106(.A1(new_n531), .A2(G651), .B1(G52), .B2(new_n517), .ZN(new_n532));
  INV_X1    g107(.A(G90), .ZN(new_n533));
  NAND2_X1  g108(.A1(new_n507), .A2(new_n510), .ZN(new_n534));
  OAI21_X1  g109(.A(new_n532), .B1(new_n533), .B2(new_n534), .ZN(G301));
  INV_X1    g110(.A(G301), .ZN(G171));
  NAND2_X1  g111(.A1(G68), .A2(G543), .ZN(new_n537));
  INV_X1    g112(.A(G56), .ZN(new_n538));
  OAI21_X1  g113(.A(new_n537), .B1(new_n503), .B2(new_n538), .ZN(new_n539));
  INV_X1    g114(.A(KEYINPUT70), .ZN(new_n540));
  NAND2_X1  g115(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  OAI211_X1 g116(.A(KEYINPUT70), .B(new_n537), .C1(new_n503), .C2(new_n538), .ZN(new_n542));
  NAND3_X1  g117(.A1(new_n541), .A2(G651), .A3(new_n542), .ZN(new_n543));
  NAND2_X1  g118(.A1(new_n517), .A2(G43), .ZN(new_n544));
  NAND3_X1  g119(.A1(new_n507), .A2(new_n510), .A3(G81), .ZN(new_n545));
  NAND3_X1  g120(.A1(new_n543), .A2(new_n544), .A3(new_n545), .ZN(new_n546));
  INV_X1    g121(.A(new_n546), .ZN(new_n547));
  NAND2_X1  g122(.A1(new_n547), .A2(G860), .ZN(G153));
  NAND4_X1  g123(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  XOR2_X1   g124(.A(KEYINPUT71), .B(KEYINPUT8), .Z(new_n550));
  NAND2_X1  g125(.A1(G1), .A2(G3), .ZN(new_n551));
  XNOR2_X1  g126(.A(new_n550), .B(new_n551), .ZN(new_n552));
  NAND4_X1  g127(.A1(G319), .A2(G483), .A3(G661), .A4(new_n552), .ZN(G188));
  NAND2_X1  g128(.A1(new_n517), .A2(G53), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n554), .A2(KEYINPUT9), .ZN(new_n555));
  INV_X1    g130(.A(KEYINPUT9), .ZN(new_n556));
  NAND3_X1  g131(.A1(new_n517), .A2(new_n556), .A3(G53), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n555), .A2(new_n557), .ZN(new_n558));
  NAND2_X1  g133(.A1(G78), .A2(G543), .ZN(new_n559));
  INV_X1    g134(.A(G65), .ZN(new_n560));
  OAI21_X1  g135(.A(new_n559), .B1(new_n503), .B2(new_n560), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n561), .A2(G651), .ZN(new_n562));
  INV_X1    g137(.A(G91), .ZN(new_n563));
  OAI211_X1 g138(.A(new_n558), .B(new_n562), .C1(new_n563), .C2(new_n534), .ZN(G299));
  OR2_X1    g139(.A1(new_n508), .A2(G74), .ZN(new_n565));
  AOI22_X1  g140(.A1(new_n565), .A2(G651), .B1(G49), .B2(new_n517), .ZN(new_n566));
  NAND3_X1  g141(.A1(new_n507), .A2(new_n510), .A3(G87), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n566), .A2(new_n567), .ZN(G288));
  NAND2_X1  g143(.A1(G73), .A2(G543), .ZN(new_n569));
  INV_X1    g144(.A(G61), .ZN(new_n570));
  OAI21_X1  g145(.A(new_n569), .B1(new_n503), .B2(new_n570), .ZN(new_n571));
  AOI22_X1  g146(.A1(new_n571), .A2(G651), .B1(G48), .B2(new_n517), .ZN(new_n572));
  INV_X1    g147(.A(G86), .ZN(new_n573));
  OAI21_X1  g148(.A(new_n572), .B1(new_n573), .B2(new_n534), .ZN(G305));
  XOR2_X1   g149(.A(KEYINPUT72), .B(G47), .Z(new_n575));
  NAND2_X1  g150(.A1(new_n517), .A2(new_n575), .ZN(new_n576));
  INV_X1    g151(.A(G651), .ZN(new_n577));
  AOI22_X1  g152(.A1(new_n508), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n578));
  INV_X1    g153(.A(G85), .ZN(new_n579));
  OAI221_X1 g154(.A(new_n576), .B1(new_n577), .B2(new_n578), .C1(new_n534), .C2(new_n579), .ZN(G290));
  INV_X1    g155(.A(G868), .ZN(new_n581));
  NOR2_X1   g156(.A1(G301), .A2(new_n581), .ZN(new_n582));
  INV_X1    g157(.A(KEYINPUT10), .ZN(new_n583));
  NAND3_X1  g158(.A1(new_n511), .A2(new_n583), .A3(G92), .ZN(new_n584));
  INV_X1    g159(.A(G92), .ZN(new_n585));
  OAI21_X1  g160(.A(KEYINPUT10), .B1(new_n534), .B2(new_n585), .ZN(new_n586));
  NAND2_X1  g161(.A1(new_n584), .A2(new_n586), .ZN(new_n587));
  NAND2_X1  g162(.A1(G79), .A2(G543), .ZN(new_n588));
  INV_X1    g163(.A(G66), .ZN(new_n589));
  OAI21_X1  g164(.A(new_n588), .B1(new_n503), .B2(new_n589), .ZN(new_n590));
  NAND2_X1  g165(.A1(new_n590), .A2(KEYINPUT73), .ZN(new_n591));
  INV_X1    g166(.A(KEYINPUT73), .ZN(new_n592));
  OAI211_X1 g167(.A(new_n592), .B(new_n588), .C1(new_n503), .C2(new_n589), .ZN(new_n593));
  NAND3_X1  g168(.A1(new_n591), .A2(G651), .A3(new_n593), .ZN(new_n594));
  NAND2_X1  g169(.A1(new_n517), .A2(G54), .ZN(new_n595));
  NAND2_X1  g170(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  OAI21_X1  g171(.A(KEYINPUT74), .B1(new_n587), .B2(new_n596), .ZN(new_n597));
  AND2_X1   g172(.A1(new_n594), .A2(new_n595), .ZN(new_n598));
  INV_X1    g173(.A(KEYINPUT74), .ZN(new_n599));
  NAND4_X1  g174(.A1(new_n598), .A2(new_n599), .A3(new_n586), .A4(new_n584), .ZN(new_n600));
  NAND2_X1  g175(.A1(new_n597), .A2(new_n600), .ZN(new_n601));
  INV_X1    g176(.A(new_n601), .ZN(new_n602));
  AOI21_X1  g177(.A(new_n582), .B1(new_n602), .B2(new_n581), .ZN(G284));
  AOI21_X1  g178(.A(new_n582), .B1(new_n602), .B2(new_n581), .ZN(G321));
  NAND2_X1  g179(.A1(G286), .A2(G868), .ZN(new_n605));
  NOR2_X1   g180(.A1(new_n605), .A2(KEYINPUT75), .ZN(new_n606));
  AND2_X1   g181(.A1(new_n605), .A2(KEYINPUT75), .ZN(new_n607));
  NAND2_X1  g182(.A1(G299), .A2(new_n581), .ZN(new_n608));
  AOI21_X1  g183(.A(new_n606), .B1(new_n607), .B2(new_n608), .ZN(G297));
  AOI21_X1  g184(.A(new_n606), .B1(new_n607), .B2(new_n608), .ZN(G280));
  INV_X1    g185(.A(G559), .ZN(new_n611));
  OAI21_X1  g186(.A(new_n602), .B1(new_n611), .B2(G860), .ZN(G148));
  INV_X1    g187(.A(KEYINPUT76), .ZN(new_n613));
  OAI21_X1  g188(.A(new_n613), .B1(new_n601), .B2(G559), .ZN(new_n614));
  NAND4_X1  g189(.A1(new_n597), .A2(new_n600), .A3(KEYINPUT76), .A4(new_n611), .ZN(new_n615));
  NAND2_X1  g190(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  MUX2_X1   g191(.A(new_n546), .B(new_n616), .S(G868), .Z(G323));
  XNOR2_X1  g192(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g193(.A1(new_n463), .A2(new_n466), .ZN(new_n619));
  XOR2_X1   g194(.A(new_n619), .B(KEYINPUT12), .Z(new_n620));
  XNOR2_X1  g195(.A(new_n620), .B(KEYINPUT13), .ZN(new_n621));
  XOR2_X1   g196(.A(new_n621), .B(G2100), .Z(new_n622));
  NAND2_X1  g197(.A1(new_n477), .A2(G135), .ZN(new_n623));
  NAND2_X1  g198(.A1(new_n472), .A2(G123), .ZN(new_n624));
  OR2_X1    g199(.A1(G99), .A2(G2105), .ZN(new_n625));
  OAI211_X1 g200(.A(new_n625), .B(G2104), .C1(G111), .C2(new_n464), .ZN(new_n626));
  AND3_X1   g201(.A1(new_n623), .A2(new_n624), .A3(new_n626), .ZN(new_n627));
  INV_X1    g202(.A(new_n627), .ZN(new_n628));
  OR2_X1    g203(.A1(new_n628), .A2(G2096), .ZN(new_n629));
  NAND2_X1  g204(.A1(new_n628), .A2(G2096), .ZN(new_n630));
  NAND3_X1  g205(.A1(new_n622), .A2(new_n629), .A3(new_n630), .ZN(G156));
  XNOR2_X1  g206(.A(G2427), .B(G2438), .ZN(new_n632));
  XNOR2_X1  g207(.A(new_n632), .B(G2430), .ZN(new_n633));
  XNOR2_X1  g208(.A(KEYINPUT15), .B(G2435), .ZN(new_n634));
  OR2_X1    g209(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  NAND2_X1  g210(.A1(new_n633), .A2(new_n634), .ZN(new_n636));
  NAND3_X1  g211(.A1(new_n635), .A2(KEYINPUT14), .A3(new_n636), .ZN(new_n637));
  XOR2_X1   g212(.A(KEYINPUT77), .B(KEYINPUT16), .Z(new_n638));
  XNOR2_X1  g213(.A(new_n637), .B(new_n638), .ZN(new_n639));
  XOR2_X1   g214(.A(G2451), .B(G2454), .Z(new_n640));
  XNOR2_X1  g215(.A(G2443), .B(G2446), .ZN(new_n641));
  XNOR2_X1  g216(.A(new_n640), .B(new_n641), .ZN(new_n642));
  XNOR2_X1  g217(.A(new_n639), .B(new_n642), .ZN(new_n643));
  XNOR2_X1  g218(.A(G1341), .B(G1348), .ZN(new_n644));
  INV_X1    g219(.A(new_n644), .ZN(new_n645));
  NAND2_X1  g220(.A1(new_n643), .A2(new_n645), .ZN(new_n646));
  XOR2_X1   g221(.A(new_n646), .B(KEYINPUT78), .Z(new_n647));
  OAI21_X1  g222(.A(G14), .B1(new_n643), .B2(new_n645), .ZN(new_n648));
  NOR2_X1   g223(.A1(new_n647), .A2(new_n648), .ZN(G401));
  XOR2_X1   g224(.A(G2072), .B(G2078), .Z(new_n650));
  XOR2_X1   g225(.A(G2084), .B(G2090), .Z(new_n651));
  XNOR2_X1  g226(.A(G2067), .B(G2678), .ZN(new_n652));
  NAND2_X1  g227(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  AOI21_X1  g228(.A(new_n650), .B1(new_n653), .B2(KEYINPUT18), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n654), .B(KEYINPUT79), .ZN(new_n655));
  XOR2_X1   g230(.A(KEYINPUT80), .B(G2100), .Z(new_n656));
  XNOR2_X1  g231(.A(new_n655), .B(new_n656), .ZN(new_n657));
  INV_X1    g232(.A(KEYINPUT18), .ZN(new_n658));
  NAND2_X1  g233(.A1(new_n653), .A2(KEYINPUT17), .ZN(new_n659));
  NOR2_X1   g234(.A1(new_n651), .A2(new_n652), .ZN(new_n660));
  OAI21_X1  g235(.A(new_n658), .B1(new_n659), .B2(new_n660), .ZN(new_n661));
  XNOR2_X1  g236(.A(new_n661), .B(G2096), .ZN(new_n662));
  XNOR2_X1  g237(.A(new_n657), .B(new_n662), .ZN(G227));
  XOR2_X1   g238(.A(G1961), .B(G1966), .Z(new_n664));
  XNOR2_X1  g239(.A(new_n664), .B(KEYINPUT81), .ZN(new_n665));
  XOR2_X1   g240(.A(G1956), .B(G2474), .Z(new_n666));
  NAND2_X1  g241(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  INV_X1    g242(.A(KEYINPUT82), .ZN(new_n668));
  NAND2_X1  g243(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  NAND3_X1  g244(.A1(new_n665), .A2(KEYINPUT82), .A3(new_n666), .ZN(new_n670));
  XNOR2_X1  g245(.A(G1971), .B(G1976), .ZN(new_n671));
  XOR2_X1   g246(.A(new_n671), .B(KEYINPUT19), .Z(new_n672));
  NAND3_X1  g247(.A1(new_n669), .A2(new_n670), .A3(new_n672), .ZN(new_n673));
  XNOR2_X1  g248(.A(new_n673), .B(KEYINPUT20), .ZN(new_n674));
  OR2_X1    g249(.A1(new_n665), .A2(new_n666), .ZN(new_n675));
  INV_X1    g250(.A(new_n672), .ZN(new_n676));
  NAND3_X1  g251(.A1(new_n675), .A2(new_n667), .A3(new_n676), .ZN(new_n677));
  OAI211_X1 g252(.A(new_n674), .B(new_n677), .C1(new_n676), .C2(new_n675), .ZN(new_n678));
  XNOR2_X1  g253(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n679));
  XNOR2_X1  g254(.A(new_n678), .B(new_n679), .ZN(new_n680));
  XNOR2_X1  g255(.A(G1991), .B(G1996), .ZN(new_n681));
  XNOR2_X1  g256(.A(new_n680), .B(new_n681), .ZN(new_n682));
  XNOR2_X1  g257(.A(G1981), .B(G1986), .ZN(new_n683));
  INV_X1    g258(.A(new_n683), .ZN(new_n684));
  NAND2_X1  g259(.A1(new_n682), .A2(new_n684), .ZN(new_n685));
  OR2_X1    g260(.A1(new_n680), .A2(new_n681), .ZN(new_n686));
  NAND2_X1  g261(.A1(new_n680), .A2(new_n681), .ZN(new_n687));
  NAND3_X1  g262(.A1(new_n686), .A2(new_n683), .A3(new_n687), .ZN(new_n688));
  AND2_X1   g263(.A1(new_n685), .A2(new_n688), .ZN(G229));
  NAND2_X1  g264(.A1(new_n477), .A2(G131), .ZN(new_n690));
  NAND2_X1  g265(.A1(new_n472), .A2(G119), .ZN(new_n691));
  NOR2_X1   g266(.A1(new_n464), .A2(G107), .ZN(new_n692));
  OAI21_X1  g267(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n693));
  OAI211_X1 g268(.A(new_n690), .B(new_n691), .C1(new_n692), .C2(new_n693), .ZN(new_n694));
  XNOR2_X1  g269(.A(new_n694), .B(KEYINPUT84), .ZN(new_n695));
  INV_X1    g270(.A(G29), .ZN(new_n696));
  OR2_X1    g271(.A1(new_n696), .A2(KEYINPUT83), .ZN(new_n697));
  NAND2_X1  g272(.A1(new_n696), .A2(KEYINPUT83), .ZN(new_n698));
  AND2_X1   g273(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  NOR2_X1   g274(.A1(new_n695), .A2(new_n699), .ZN(new_n700));
  AOI21_X1  g275(.A(new_n700), .B1(G25), .B2(new_n699), .ZN(new_n701));
  XOR2_X1   g276(.A(KEYINPUT35), .B(G1991), .Z(new_n702));
  AND2_X1   g277(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  NOR2_X1   g278(.A1(new_n701), .A2(new_n702), .ZN(new_n704));
  MUX2_X1   g279(.A(G24), .B(G290), .S(G16), .Z(new_n705));
  XNOR2_X1  g280(.A(new_n705), .B(G1986), .ZN(new_n706));
  NOR3_X1   g281(.A1(new_n703), .A2(new_n704), .A3(new_n706), .ZN(new_n707));
  INV_X1    g282(.A(G16), .ZN(new_n708));
  NAND2_X1  g283(.A1(new_n708), .A2(G22), .ZN(new_n709));
  OAI21_X1  g284(.A(new_n709), .B1(G166), .B2(new_n708), .ZN(new_n710));
  INV_X1    g285(.A(G1971), .ZN(new_n711));
  XNOR2_X1  g286(.A(new_n710), .B(new_n711), .ZN(new_n712));
  NOR2_X1   g287(.A1(G16), .A2(G23), .ZN(new_n713));
  XNOR2_X1  g288(.A(new_n713), .B(KEYINPUT85), .ZN(new_n714));
  OAI21_X1  g289(.A(new_n714), .B1(G288), .B2(new_n708), .ZN(new_n715));
  XOR2_X1   g290(.A(KEYINPUT33), .B(G1976), .Z(new_n716));
  XNOR2_X1  g291(.A(new_n715), .B(new_n716), .ZN(new_n717));
  MUX2_X1   g292(.A(G6), .B(G305), .S(G16), .Z(new_n718));
  XOR2_X1   g293(.A(KEYINPUT32), .B(G1981), .Z(new_n719));
  XNOR2_X1  g294(.A(new_n718), .B(new_n719), .ZN(new_n720));
  NAND3_X1  g295(.A1(new_n712), .A2(new_n717), .A3(new_n720), .ZN(new_n721));
  NAND2_X1  g296(.A1(new_n721), .A2(KEYINPUT34), .ZN(new_n722));
  OR2_X1    g297(.A1(new_n721), .A2(KEYINPUT34), .ZN(new_n723));
  NAND3_X1  g298(.A1(new_n707), .A2(new_n722), .A3(new_n723), .ZN(new_n724));
  XOR2_X1   g299(.A(new_n724), .B(KEYINPUT36), .Z(new_n725));
  INV_X1    g300(.A(KEYINPUT99), .ZN(new_n726));
  NAND2_X1  g301(.A1(new_n699), .A2(G26), .ZN(new_n727));
  XOR2_X1   g302(.A(new_n727), .B(KEYINPUT28), .Z(new_n728));
  NAND2_X1  g303(.A1(new_n472), .A2(G128), .ZN(new_n729));
  XNOR2_X1  g304(.A(new_n729), .B(KEYINPUT86), .ZN(new_n730));
  OAI21_X1  g305(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n731));
  INV_X1    g306(.A(G116), .ZN(new_n732));
  AOI21_X1  g307(.A(new_n731), .B1(new_n732), .B2(G2105), .ZN(new_n733));
  INV_X1    g308(.A(KEYINPUT87), .ZN(new_n734));
  OR2_X1    g309(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  NAND2_X1  g310(.A1(new_n733), .A2(new_n734), .ZN(new_n736));
  AOI22_X1  g311(.A1(new_n477), .A2(G140), .B1(new_n735), .B2(new_n736), .ZN(new_n737));
  NAND2_X1  g312(.A1(new_n730), .A2(new_n737), .ZN(new_n738));
  AOI21_X1  g313(.A(new_n728), .B1(new_n738), .B2(G29), .ZN(new_n739));
  XNOR2_X1  g314(.A(KEYINPUT88), .B(G2067), .ZN(new_n740));
  XNOR2_X1  g315(.A(new_n739), .B(new_n740), .ZN(new_n741));
  NAND2_X1  g316(.A1(new_n708), .A2(G19), .ZN(new_n742));
  OAI21_X1  g317(.A(new_n742), .B1(new_n547), .B2(new_n708), .ZN(new_n743));
  NAND2_X1  g318(.A1(new_n743), .A2(G1341), .ZN(new_n744));
  OR2_X1    g319(.A1(new_n743), .A2(G1341), .ZN(new_n745));
  AND3_X1   g320(.A1(new_n741), .A2(new_n744), .A3(new_n745), .ZN(new_n746));
  NAND2_X1  g321(.A1(new_n708), .A2(G4), .ZN(new_n747));
  OAI21_X1  g322(.A(new_n747), .B1(new_n602), .B2(new_n708), .ZN(new_n748));
  OR2_X1    g323(.A1(new_n748), .A2(G1348), .ZN(new_n749));
  NAND2_X1  g324(.A1(new_n748), .A2(G1348), .ZN(new_n750));
  NAND3_X1  g325(.A1(new_n746), .A2(new_n749), .A3(new_n750), .ZN(new_n751));
  INV_X1    g326(.A(KEYINPUT89), .ZN(new_n752));
  XNOR2_X1  g327(.A(new_n751), .B(new_n752), .ZN(new_n753));
  INV_X1    g328(.A(new_n699), .ZN(new_n754));
  INV_X1    g329(.A(KEYINPUT24), .ZN(new_n755));
  NOR2_X1   g330(.A1(new_n755), .A2(G34), .ZN(new_n756));
  OR3_X1    g331(.A1(new_n754), .A2(KEYINPUT93), .A3(new_n756), .ZN(new_n757));
  OAI21_X1  g332(.A(KEYINPUT93), .B1(new_n754), .B2(new_n756), .ZN(new_n758));
  NAND2_X1  g333(.A1(new_n755), .A2(G34), .ZN(new_n759));
  NAND3_X1  g334(.A1(new_n757), .A2(new_n758), .A3(new_n759), .ZN(new_n760));
  OAI21_X1  g335(.A(new_n760), .B1(new_n696), .B2(new_n469), .ZN(new_n761));
  INV_X1    g336(.A(G2084), .ZN(new_n762));
  OR2_X1    g337(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  NAND2_X1  g338(.A1(new_n699), .A2(G27), .ZN(new_n764));
  OAI21_X1  g339(.A(new_n764), .B1(G164), .B2(new_n699), .ZN(new_n765));
  AOI22_X1  g340(.A1(new_n627), .A2(new_n754), .B1(G2078), .B2(new_n765), .ZN(new_n766));
  INV_X1    g341(.A(KEYINPUT30), .ZN(new_n767));
  AND2_X1   g342(.A1(new_n767), .A2(G28), .ZN(new_n768));
  OAI21_X1  g343(.A(new_n696), .B1(new_n767), .B2(G28), .ZN(new_n769));
  AND2_X1   g344(.A1(KEYINPUT31), .A2(G11), .ZN(new_n770));
  NOR2_X1   g345(.A1(KEYINPUT31), .A2(G11), .ZN(new_n771));
  OAI22_X1  g346(.A1(new_n768), .A2(new_n769), .B1(new_n770), .B2(new_n771), .ZN(new_n772));
  AOI21_X1  g347(.A(new_n772), .B1(new_n761), .B2(new_n762), .ZN(new_n773));
  OR2_X1    g348(.A1(new_n765), .A2(G2078), .ZN(new_n774));
  NAND4_X1  g349(.A1(new_n763), .A2(new_n766), .A3(new_n773), .A4(new_n774), .ZN(new_n775));
  NOR2_X1   g350(.A1(G5), .A2(G16), .ZN(new_n776));
  XOR2_X1   g351(.A(new_n776), .B(KEYINPUT97), .Z(new_n777));
  OAI21_X1  g352(.A(new_n777), .B1(G301), .B2(new_n708), .ZN(new_n778));
  INV_X1    g353(.A(G1961), .ZN(new_n779));
  NOR2_X1   g354(.A1(new_n778), .A2(new_n779), .ZN(new_n780));
  AND2_X1   g355(.A1(new_n778), .A2(new_n779), .ZN(new_n781));
  OR3_X1    g356(.A1(new_n775), .A2(new_n780), .A3(new_n781), .ZN(new_n782));
  NOR2_X1   g357(.A1(G29), .A2(G33), .ZN(new_n783));
  XOR2_X1   g358(.A(new_n783), .B(KEYINPUT90), .Z(new_n784));
  NAND2_X1  g359(.A1(new_n477), .A2(G139), .ZN(new_n785));
  XNOR2_X1  g360(.A(new_n785), .B(KEYINPUT92), .ZN(new_n786));
  NAND3_X1  g361(.A1(new_n464), .A2(G103), .A3(G2104), .ZN(new_n787));
  XNOR2_X1  g362(.A(new_n787), .B(KEYINPUT91), .ZN(new_n788));
  XOR2_X1   g363(.A(new_n788), .B(KEYINPUT25), .Z(new_n789));
  NAND2_X1  g364(.A1(new_n463), .A2(G127), .ZN(new_n790));
  NAND2_X1  g365(.A1(G115), .A2(G2104), .ZN(new_n791));
  AOI21_X1  g366(.A(new_n464), .B1(new_n790), .B2(new_n791), .ZN(new_n792));
  NOR2_X1   g367(.A1(new_n789), .A2(new_n792), .ZN(new_n793));
  NAND2_X1  g368(.A1(new_n786), .A2(new_n793), .ZN(new_n794));
  OAI21_X1  g369(.A(new_n784), .B1(new_n794), .B2(new_n696), .ZN(new_n795));
  XOR2_X1   g370(.A(new_n795), .B(G2072), .Z(new_n796));
  INV_X1    g371(.A(G21), .ZN(new_n797));
  AOI21_X1  g372(.A(KEYINPUT96), .B1(new_n708), .B2(new_n797), .ZN(new_n798));
  NAND2_X1  g373(.A1(G168), .A2(G16), .ZN(new_n799));
  MUX2_X1   g374(.A(KEYINPUT96), .B(new_n798), .S(new_n799), .Z(new_n800));
  AOI211_X1 g375(.A(new_n782), .B(new_n796), .C1(G1966), .C2(new_n800), .ZN(new_n801));
  NOR2_X1   g376(.A1(new_n754), .A2(G35), .ZN(new_n802));
  AOI21_X1  g377(.A(new_n802), .B1(G162), .B2(new_n754), .ZN(new_n803));
  XOR2_X1   g378(.A(new_n803), .B(KEYINPUT29), .Z(new_n804));
  INV_X1    g379(.A(G2090), .ZN(new_n805));
  NAND2_X1  g380(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  INV_X1    g381(.A(KEYINPUT98), .ZN(new_n807));
  XNOR2_X1  g382(.A(new_n806), .B(new_n807), .ZN(new_n808));
  NAND2_X1  g383(.A1(new_n477), .A2(G141), .ZN(new_n809));
  NAND2_X1  g384(.A1(new_n472), .A2(G129), .ZN(new_n810));
  NAND3_X1  g385(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n811));
  INV_X1    g386(.A(KEYINPUT26), .ZN(new_n812));
  OR2_X1    g387(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  NAND2_X1  g388(.A1(new_n811), .A2(new_n812), .ZN(new_n814));
  AOI22_X1  g389(.A1(new_n813), .A2(new_n814), .B1(G105), .B2(new_n466), .ZN(new_n815));
  NAND3_X1  g390(.A1(new_n809), .A2(new_n810), .A3(new_n815), .ZN(new_n816));
  XOR2_X1   g391(.A(new_n816), .B(KEYINPUT94), .Z(new_n817));
  NAND2_X1  g392(.A1(new_n817), .A2(G29), .ZN(new_n818));
  OR2_X1    g393(.A1(new_n818), .A2(KEYINPUT95), .ZN(new_n819));
  OAI211_X1 g394(.A(new_n818), .B(KEYINPUT95), .C1(G29), .C2(G32), .ZN(new_n820));
  NAND2_X1  g395(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  XNOR2_X1  g396(.A(KEYINPUT27), .B(G1996), .ZN(new_n822));
  XNOR2_X1  g397(.A(new_n821), .B(new_n822), .ZN(new_n823));
  NOR2_X1   g398(.A1(new_n804), .A2(new_n805), .ZN(new_n824));
  NAND2_X1  g399(.A1(new_n708), .A2(G20), .ZN(new_n825));
  XNOR2_X1  g400(.A(new_n825), .B(KEYINPUT23), .ZN(new_n826));
  INV_X1    g401(.A(G299), .ZN(new_n827));
  OAI21_X1  g402(.A(new_n826), .B1(new_n827), .B2(new_n708), .ZN(new_n828));
  XNOR2_X1  g403(.A(new_n828), .B(G1956), .ZN(new_n829));
  NOR2_X1   g404(.A1(new_n800), .A2(G1966), .ZN(new_n830));
  NOR3_X1   g405(.A1(new_n824), .A2(new_n829), .A3(new_n830), .ZN(new_n831));
  AND4_X1   g406(.A1(new_n801), .A2(new_n808), .A3(new_n823), .A4(new_n831), .ZN(new_n832));
  AOI21_X1  g407(.A(new_n726), .B1(new_n753), .B2(new_n832), .ZN(new_n833));
  INV_X1    g408(.A(new_n833), .ZN(new_n834));
  NAND3_X1  g409(.A1(new_n753), .A2(new_n832), .A3(new_n726), .ZN(new_n835));
  AOI21_X1  g410(.A(new_n725), .B1(new_n834), .B2(new_n835), .ZN(G311));
  INV_X1    g411(.A(new_n725), .ZN(new_n837));
  INV_X1    g412(.A(new_n835), .ZN(new_n838));
  OAI21_X1  g413(.A(new_n837), .B1(new_n838), .B2(new_n833), .ZN(G150));
  NAND2_X1  g414(.A1(new_n546), .A2(KEYINPUT101), .ZN(new_n840));
  INV_X1    g415(.A(KEYINPUT101), .ZN(new_n841));
  NAND4_X1  g416(.A1(new_n543), .A2(new_n841), .A3(new_n544), .A4(new_n545), .ZN(new_n842));
  XNOR2_X1  g417(.A(KEYINPUT100), .B(G93), .ZN(new_n843));
  NOR2_X1   g418(.A1(new_n534), .A2(new_n843), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n517), .A2(G55), .ZN(new_n845));
  AOI22_X1  g420(.A1(new_n508), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n846));
  OAI21_X1  g421(.A(new_n845), .B1(new_n846), .B2(new_n577), .ZN(new_n847));
  NOR2_X1   g422(.A1(new_n844), .A2(new_n847), .ZN(new_n848));
  NAND3_X1  g423(.A1(new_n840), .A2(new_n842), .A3(new_n848), .ZN(new_n849));
  OAI211_X1 g424(.A(new_n546), .B(KEYINPUT101), .C1(new_n844), .C2(new_n847), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n849), .A2(new_n850), .ZN(new_n851));
  XOR2_X1   g426(.A(new_n851), .B(KEYINPUT38), .Z(new_n852));
  NOR2_X1   g427(.A1(new_n601), .A2(new_n611), .ZN(new_n853));
  XNOR2_X1  g428(.A(new_n852), .B(new_n853), .ZN(new_n854));
  INV_X1    g429(.A(KEYINPUT39), .ZN(new_n855));
  AOI21_X1  g430(.A(G860), .B1(new_n854), .B2(new_n855), .ZN(new_n856));
  OAI21_X1  g431(.A(new_n856), .B1(new_n855), .B2(new_n854), .ZN(new_n857));
  OAI21_X1  g432(.A(G860), .B1(new_n844), .B2(new_n847), .ZN(new_n858));
  XOR2_X1   g433(.A(new_n858), .B(KEYINPUT37), .Z(new_n859));
  NAND2_X1  g434(.A1(new_n857), .A2(new_n859), .ZN(G145));
  XNOR2_X1  g435(.A(new_n627), .B(G160), .ZN(new_n861));
  XOR2_X1   g436(.A(new_n861), .B(G162), .Z(new_n862));
  AOI22_X1  g437(.A1(new_n463), .A2(new_n484), .B1(new_n480), .B2(new_n482), .ZN(new_n863));
  INV_X1    g438(.A(new_n494), .ZN(new_n864));
  AOI21_X1  g439(.A(new_n493), .B1(new_n463), .B2(new_n490), .ZN(new_n865));
  OAI21_X1  g440(.A(new_n863), .B1(new_n864), .B2(new_n865), .ZN(new_n866));
  XNOR2_X1  g441(.A(new_n738), .B(new_n866), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n477), .A2(G142), .ZN(new_n868));
  NAND2_X1  g443(.A1(new_n472), .A2(G130), .ZN(new_n869));
  OR2_X1    g444(.A1(G106), .A2(G2105), .ZN(new_n870));
  OAI211_X1 g445(.A(new_n870), .B(G2104), .C1(G118), .C2(new_n464), .ZN(new_n871));
  NAND3_X1  g446(.A1(new_n868), .A2(new_n869), .A3(new_n871), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n867), .A2(new_n872), .ZN(new_n873));
  INV_X1    g448(.A(new_n873), .ZN(new_n874));
  NOR2_X1   g449(.A1(new_n867), .A2(new_n872), .ZN(new_n875));
  OR2_X1    g450(.A1(new_n695), .A2(KEYINPUT102), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n695), .A2(KEYINPUT102), .ZN(new_n877));
  INV_X1    g452(.A(new_n620), .ZN(new_n878));
  AND3_X1   g453(.A1(new_n876), .A2(new_n877), .A3(new_n878), .ZN(new_n879));
  AOI21_X1  g454(.A(new_n878), .B1(new_n876), .B2(new_n877), .ZN(new_n880));
  OAI22_X1  g455(.A1(new_n874), .A2(new_n875), .B1(new_n879), .B2(new_n880), .ZN(new_n881));
  INV_X1    g456(.A(new_n875), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n876), .A2(new_n877), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n883), .A2(new_n620), .ZN(new_n884));
  NAND3_X1  g459(.A1(new_n876), .A2(new_n877), .A3(new_n878), .ZN(new_n885));
  NAND4_X1  g460(.A1(new_n882), .A2(new_n884), .A3(new_n885), .A4(new_n873), .ZN(new_n886));
  INV_X1    g461(.A(new_n816), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n794), .A2(new_n887), .ZN(new_n888));
  OAI21_X1  g463(.A(new_n888), .B1(new_n817), .B2(new_n794), .ZN(new_n889));
  AND3_X1   g464(.A1(new_n881), .A2(new_n886), .A3(new_n889), .ZN(new_n890));
  AOI21_X1  g465(.A(new_n889), .B1(new_n881), .B2(new_n886), .ZN(new_n891));
  OAI21_X1  g466(.A(new_n862), .B1(new_n890), .B2(new_n891), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n881), .A2(new_n886), .ZN(new_n893));
  INV_X1    g468(.A(new_n889), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  INV_X1    g470(.A(new_n862), .ZN(new_n896));
  NAND3_X1  g471(.A1(new_n881), .A2(new_n886), .A3(new_n889), .ZN(new_n897));
  NAND3_X1  g472(.A1(new_n895), .A2(new_n896), .A3(new_n897), .ZN(new_n898));
  INV_X1    g473(.A(G37), .ZN(new_n899));
  NAND3_X1  g474(.A1(new_n892), .A2(new_n898), .A3(new_n899), .ZN(new_n900));
  XNOR2_X1  g475(.A(new_n900), .B(KEYINPUT40), .ZN(G395));
  AND3_X1   g476(.A1(new_n614), .A2(KEYINPUT103), .A3(new_n615), .ZN(new_n902));
  AOI21_X1  g477(.A(KEYINPUT103), .B1(new_n614), .B2(new_n615), .ZN(new_n903));
  OAI21_X1  g478(.A(new_n851), .B1(new_n902), .B2(new_n903), .ZN(new_n904));
  INV_X1    g479(.A(KEYINPUT103), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n616), .A2(new_n905), .ZN(new_n906));
  INV_X1    g481(.A(new_n851), .ZN(new_n907));
  NAND3_X1  g482(.A1(new_n614), .A2(KEYINPUT103), .A3(new_n615), .ZN(new_n908));
  NAND3_X1  g483(.A1(new_n906), .A2(new_n907), .A3(new_n908), .ZN(new_n909));
  NAND3_X1  g484(.A1(new_n598), .A2(new_n586), .A3(new_n584), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n910), .A2(G299), .ZN(new_n911));
  NOR2_X1   g486(.A1(new_n587), .A2(new_n596), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n912), .A2(new_n827), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n911), .A2(new_n913), .ZN(new_n914));
  INV_X1    g489(.A(KEYINPUT41), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  NAND3_X1  g491(.A1(new_n911), .A2(new_n913), .A3(KEYINPUT41), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  AND3_X1   g493(.A1(new_n904), .A2(new_n909), .A3(new_n918), .ZN(new_n919));
  AND2_X1   g494(.A1(new_n911), .A2(new_n913), .ZN(new_n920));
  AOI21_X1  g495(.A(new_n920), .B1(new_n904), .B2(new_n909), .ZN(new_n921));
  OAI21_X1  g496(.A(KEYINPUT42), .B1(new_n919), .B2(new_n921), .ZN(new_n922));
  INV_X1    g497(.A(KEYINPUT42), .ZN(new_n923));
  NAND3_X1  g498(.A1(new_n904), .A2(new_n909), .A3(new_n918), .ZN(new_n924));
  AND2_X1   g499(.A1(new_n904), .A2(new_n909), .ZN(new_n925));
  OAI211_X1 g500(.A(new_n923), .B(new_n924), .C1(new_n925), .C2(new_n920), .ZN(new_n926));
  XOR2_X1   g501(.A(G303), .B(G290), .Z(new_n927));
  INV_X1    g502(.A(G288), .ZN(new_n928));
  XNOR2_X1  g503(.A(new_n928), .B(G305), .ZN(new_n929));
  XNOR2_X1  g504(.A(new_n927), .B(new_n929), .ZN(new_n930));
  INV_X1    g505(.A(new_n930), .ZN(new_n931));
  AND3_X1   g506(.A1(new_n922), .A2(new_n926), .A3(new_n931), .ZN(new_n932));
  AOI21_X1  g507(.A(new_n931), .B1(new_n922), .B2(new_n926), .ZN(new_n933));
  OAI21_X1  g508(.A(G868), .B1(new_n932), .B2(new_n933), .ZN(new_n934));
  OAI21_X1  g509(.A(new_n581), .B1(new_n844), .B2(new_n847), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n934), .A2(new_n935), .ZN(G295));
  NAND2_X1  g511(.A1(new_n934), .A2(new_n935), .ZN(G331));
  INV_X1    g512(.A(KEYINPUT44), .ZN(new_n938));
  AND2_X1   g513(.A1(new_n916), .A2(new_n917), .ZN(new_n939));
  NOR2_X1   g514(.A1(G301), .A2(G286), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n511), .A2(G90), .ZN(new_n941));
  AOI22_X1  g516(.A1(new_n941), .A2(new_n532), .B1(new_n525), .B2(new_n526), .ZN(new_n942));
  NOR2_X1   g517(.A1(new_n940), .A2(new_n942), .ZN(new_n943));
  NAND3_X1  g518(.A1(new_n849), .A2(new_n943), .A3(new_n850), .ZN(new_n944));
  INV_X1    g519(.A(KEYINPUT105), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n944), .A2(new_n945), .ZN(new_n946));
  INV_X1    g521(.A(new_n943), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n851), .A2(new_n947), .ZN(new_n948));
  NAND4_X1  g523(.A1(new_n849), .A2(new_n943), .A3(KEYINPUT105), .A4(new_n850), .ZN(new_n949));
  NAND3_X1  g524(.A1(new_n946), .A2(new_n948), .A3(new_n949), .ZN(new_n950));
  AOI21_X1  g525(.A(new_n943), .B1(new_n849), .B2(new_n850), .ZN(new_n951));
  NOR2_X1   g526(.A1(new_n951), .A2(new_n914), .ZN(new_n952));
  INV_X1    g527(.A(KEYINPUT104), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n944), .A2(new_n953), .ZN(new_n954));
  NAND4_X1  g529(.A1(new_n849), .A2(new_n943), .A3(KEYINPUT104), .A4(new_n850), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n954), .A2(new_n955), .ZN(new_n956));
  AOI22_X1  g531(.A1(new_n939), .A2(new_n950), .B1(new_n952), .B2(new_n956), .ZN(new_n957));
  OAI21_X1  g532(.A(new_n899), .B1(new_n957), .B2(new_n930), .ZN(new_n958));
  INV_X1    g533(.A(new_n958), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n956), .A2(new_n948), .ZN(new_n960));
  NAND2_X1  g535(.A1(new_n960), .A2(new_n939), .ZN(new_n961));
  INV_X1    g536(.A(KEYINPUT106), .ZN(new_n962));
  NAND4_X1  g537(.A1(new_n946), .A2(new_n948), .A3(new_n920), .A4(new_n949), .ZN(new_n963));
  NAND4_X1  g538(.A1(new_n961), .A2(new_n962), .A3(new_n930), .A4(new_n963), .ZN(new_n964));
  AOI21_X1  g539(.A(new_n951), .B1(new_n954), .B2(new_n955), .ZN(new_n965));
  OAI211_X1 g540(.A(new_n930), .B(new_n963), .C1(new_n965), .C2(new_n918), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n966), .A2(KEYINPUT106), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n964), .A2(new_n967), .ZN(new_n968));
  INV_X1    g543(.A(KEYINPUT43), .ZN(new_n969));
  NAND3_X1  g544(.A1(new_n959), .A2(new_n968), .A3(new_n969), .ZN(new_n970));
  OAI21_X1  g545(.A(new_n963), .B1(new_n965), .B2(new_n918), .ZN(new_n971));
  AOI21_X1  g546(.A(G37), .B1(new_n971), .B2(new_n931), .ZN(new_n972));
  AOI21_X1  g547(.A(new_n969), .B1(new_n968), .B2(new_n972), .ZN(new_n973));
  INV_X1    g548(.A(KEYINPUT107), .ZN(new_n974));
  OAI21_X1  g549(.A(new_n970), .B1(new_n973), .B2(new_n974), .ZN(new_n975));
  AOI211_X1 g550(.A(KEYINPUT107), .B(new_n969), .C1(new_n968), .C2(new_n972), .ZN(new_n976));
  OAI21_X1  g551(.A(new_n938), .B1(new_n975), .B2(new_n976), .ZN(new_n977));
  NAND3_X1  g552(.A1(new_n968), .A2(new_n969), .A3(new_n972), .ZN(new_n978));
  AOI21_X1  g553(.A(new_n958), .B1(new_n967), .B2(new_n964), .ZN(new_n979));
  INV_X1    g554(.A(KEYINPUT108), .ZN(new_n980));
  OAI21_X1  g555(.A(KEYINPUT43), .B1(new_n979), .B2(new_n980), .ZN(new_n981));
  AND3_X1   g556(.A1(new_n959), .A2(new_n968), .A3(new_n980), .ZN(new_n982));
  OAI211_X1 g557(.A(KEYINPUT44), .B(new_n978), .C1(new_n981), .C2(new_n982), .ZN(new_n983));
  NAND2_X1  g558(.A1(new_n977), .A2(new_n983), .ZN(G397));
  INV_X1    g559(.A(KEYINPUT50), .ZN(new_n985));
  INV_X1    g560(.A(G1384), .ZN(new_n986));
  NAND3_X1  g561(.A1(new_n866), .A2(new_n985), .A3(new_n986), .ZN(new_n987));
  INV_X1    g562(.A(KEYINPUT111), .ZN(new_n988));
  NAND2_X1  g563(.A1(new_n987), .A2(new_n988), .ZN(new_n989));
  NAND4_X1  g564(.A1(new_n866), .A2(KEYINPUT111), .A3(new_n985), .A4(new_n986), .ZN(new_n990));
  OAI211_X1 g565(.A(G40), .B(new_n467), .C1(new_n468), .C2(new_n464), .ZN(new_n991));
  INV_X1    g566(.A(new_n991), .ZN(new_n992));
  OAI21_X1  g567(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n993));
  NAND4_X1  g568(.A1(new_n989), .A2(new_n990), .A3(new_n992), .A4(new_n993), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n994), .A2(KEYINPUT119), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n866), .A2(new_n986), .ZN(new_n996));
  AOI21_X1  g571(.A(new_n991), .B1(new_n996), .B2(KEYINPUT50), .ZN(new_n997));
  INV_X1    g572(.A(KEYINPUT119), .ZN(new_n998));
  NAND4_X1  g573(.A1(new_n997), .A2(new_n989), .A3(new_n998), .A4(new_n990), .ZN(new_n999));
  NAND3_X1  g574(.A1(new_n995), .A2(new_n779), .A3(new_n999), .ZN(new_n1000));
  INV_X1    g575(.A(KEYINPUT124), .ZN(new_n1001));
  INV_X1    g576(.A(KEYINPUT45), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n996), .A2(new_n1002), .ZN(new_n1003));
  NAND3_X1  g578(.A1(new_n866), .A2(KEYINPUT45), .A3(new_n986), .ZN(new_n1004));
  NAND3_X1  g579(.A1(new_n1003), .A2(new_n992), .A3(new_n1004), .ZN(new_n1005));
  NOR2_X1   g580(.A1(new_n1005), .A2(G2078), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n1006), .A2(KEYINPUT53), .ZN(new_n1007));
  NAND3_X1  g582(.A1(new_n1000), .A2(new_n1001), .A3(new_n1007), .ZN(new_n1008));
  OR2_X1    g583(.A1(new_n1006), .A2(KEYINPUT53), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n1008), .A2(new_n1009), .ZN(new_n1010));
  AOI21_X1  g585(.A(new_n1001), .B1(new_n1000), .B2(new_n1007), .ZN(new_n1011));
  OAI21_X1  g586(.A(G171), .B1(new_n1010), .B2(new_n1011), .ZN(new_n1012));
  INV_X1    g587(.A(KEYINPUT125), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n1012), .A2(new_n1013), .ZN(new_n1014));
  OAI211_X1 g589(.A(KEYINPUT125), .B(G171), .C1(new_n1010), .C2(new_n1011), .ZN(new_n1015));
  NAND3_X1  g590(.A1(new_n1009), .A2(new_n1000), .A3(new_n1007), .ZN(new_n1016));
  OR2_X1    g591(.A1(new_n1016), .A2(G171), .ZN(new_n1017));
  NAND3_X1  g592(.A1(new_n1014), .A2(new_n1015), .A3(new_n1017), .ZN(new_n1018));
  INV_X1    g593(.A(KEYINPUT54), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n1018), .A2(new_n1019), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n1020), .A2(KEYINPUT126), .ZN(new_n1021));
  INV_X1    g596(.A(KEYINPUT126), .ZN(new_n1022));
  NAND3_X1  g597(.A1(new_n1018), .A2(new_n1022), .A3(new_n1019), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n993), .A2(new_n992), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n1024), .A2(KEYINPUT115), .ZN(new_n1025));
  INV_X1    g600(.A(KEYINPUT115), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n997), .A2(new_n1026), .ZN(new_n1027));
  NAND3_X1  g602(.A1(new_n1025), .A2(new_n987), .A3(new_n1027), .ZN(new_n1028));
  INV_X1    g603(.A(G1956), .ZN(new_n1029));
  NAND2_X1  g604(.A1(new_n1028), .A2(new_n1029), .ZN(new_n1030));
  INV_X1    g605(.A(KEYINPUT57), .ZN(new_n1031));
  OAI21_X1  g606(.A(new_n1031), .B1(new_n827), .B2(KEYINPUT118), .ZN(new_n1032));
  INV_X1    g607(.A(KEYINPUT118), .ZN(new_n1033));
  NAND3_X1  g608(.A1(G299), .A2(new_n1033), .A3(KEYINPUT57), .ZN(new_n1034));
  INV_X1    g609(.A(new_n1005), .ZN(new_n1035));
  XNOR2_X1  g610(.A(KEYINPUT56), .B(G2072), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n1035), .A2(new_n1036), .ZN(new_n1037));
  NAND4_X1  g612(.A1(new_n1030), .A2(new_n1032), .A3(new_n1034), .A4(new_n1037), .ZN(new_n1038));
  INV_X1    g613(.A(G1348), .ZN(new_n1039));
  NAND3_X1  g614(.A1(new_n995), .A2(new_n1039), .A3(new_n999), .ZN(new_n1040));
  NOR2_X1   g615(.A1(new_n996), .A2(new_n991), .ZN(new_n1041));
  INV_X1    g616(.A(G2067), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n1041), .A2(new_n1042), .ZN(new_n1043));
  AND3_X1   g618(.A1(new_n1040), .A2(KEYINPUT120), .A3(new_n1043), .ZN(new_n1044));
  AOI21_X1  g619(.A(KEYINPUT120), .B1(new_n1040), .B2(new_n1043), .ZN(new_n1045));
  NOR3_X1   g620(.A1(new_n1044), .A2(new_n1045), .A3(new_n910), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n1032), .A2(new_n1034), .ZN(new_n1047));
  INV_X1    g622(.A(new_n1037), .ZN(new_n1048));
  INV_X1    g623(.A(new_n987), .ZN(new_n1049));
  AOI21_X1  g624(.A(new_n1049), .B1(new_n1024), .B2(KEYINPUT115), .ZN(new_n1050));
  AOI21_X1  g625(.A(G1956), .B1(new_n1050), .B2(new_n1027), .ZN(new_n1051));
  OAI21_X1  g626(.A(new_n1047), .B1(new_n1048), .B2(new_n1051), .ZN(new_n1052));
  INV_X1    g627(.A(new_n1052), .ZN(new_n1053));
  OAI21_X1  g628(.A(new_n1038), .B1(new_n1046), .B2(new_n1053), .ZN(new_n1054));
  NAND2_X1  g629(.A1(new_n1038), .A2(new_n1052), .ZN(new_n1055));
  XNOR2_X1  g630(.A(KEYINPUT121), .B(KEYINPUT61), .ZN(new_n1056));
  XNOR2_X1  g631(.A(KEYINPUT58), .B(G1341), .ZN(new_n1057));
  OAI22_X1  g632(.A1(new_n1005), .A2(G1996), .B1(new_n1041), .B2(new_n1057), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n1058), .A2(new_n547), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n1059), .A2(KEYINPUT59), .ZN(new_n1060));
  OR2_X1    g635(.A1(new_n1059), .A2(KEYINPUT59), .ZN(new_n1061));
  AOI22_X1  g636(.A1(new_n1055), .A2(new_n1056), .B1(new_n1060), .B2(new_n1061), .ZN(new_n1062));
  INV_X1    g637(.A(KEYINPUT122), .ZN(new_n1063));
  INV_X1    g638(.A(KEYINPUT61), .ZN(new_n1064));
  OAI21_X1  g639(.A(new_n1063), .B1(new_n1055), .B2(new_n1064), .ZN(new_n1065));
  OAI211_X1 g640(.A(KEYINPUT60), .B(new_n910), .C1(new_n1044), .C2(new_n1045), .ZN(new_n1066));
  NAND4_X1  g641(.A1(new_n1038), .A2(new_n1052), .A3(KEYINPUT122), .A4(KEYINPUT61), .ZN(new_n1067));
  NAND4_X1  g642(.A1(new_n1062), .A2(new_n1065), .A3(new_n1066), .A4(new_n1067), .ZN(new_n1068));
  OAI21_X1  g643(.A(KEYINPUT60), .B1(new_n1044), .B2(new_n1045), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n1069), .A2(new_n912), .ZN(new_n1070));
  NOR3_X1   g645(.A1(new_n1044), .A2(new_n1045), .A3(KEYINPUT60), .ZN(new_n1071));
  NOR2_X1   g646(.A1(new_n1070), .A2(new_n1071), .ZN(new_n1072));
  OAI21_X1  g647(.A(new_n1054), .B1(new_n1068), .B2(new_n1072), .ZN(new_n1073));
  NAND2_X1  g648(.A1(G305), .A2(G1981), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n511), .A2(G86), .ZN(new_n1075));
  INV_X1    g650(.A(G1981), .ZN(new_n1076));
  NAND3_X1  g651(.A1(new_n1075), .A2(new_n1076), .A3(new_n572), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n1074), .A2(new_n1077), .ZN(new_n1078));
  NOR2_X1   g653(.A1(KEYINPUT114), .A2(KEYINPUT49), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n1078), .A2(new_n1079), .ZN(new_n1080));
  INV_X1    g655(.A(G8), .ZN(new_n1081));
  NOR2_X1   g656(.A1(new_n1041), .A2(new_n1081), .ZN(new_n1082));
  OAI211_X1 g657(.A(new_n1074), .B(new_n1077), .C1(KEYINPUT114), .C2(KEYINPUT49), .ZN(new_n1083));
  NAND3_X1  g658(.A1(new_n1080), .A2(new_n1082), .A3(new_n1083), .ZN(new_n1084));
  INV_X1    g659(.A(KEYINPUT52), .ZN(new_n1085));
  NAND3_X1  g660(.A1(new_n566), .A2(G1976), .A3(new_n567), .ZN(new_n1086));
  AOI21_X1  g661(.A(new_n1085), .B1(new_n1082), .B2(new_n1086), .ZN(new_n1087));
  AND2_X1   g662(.A1(new_n1082), .A2(new_n1086), .ZN(new_n1088));
  INV_X1    g663(.A(G1976), .ZN(new_n1089));
  AOI21_X1  g664(.A(KEYINPUT52), .B1(G288), .B2(new_n1089), .ZN(new_n1090));
  AOI21_X1  g665(.A(new_n1087), .B1(new_n1088), .B2(new_n1090), .ZN(new_n1091));
  NAND3_X1  g666(.A1(new_n1050), .A2(new_n805), .A3(new_n1027), .ZN(new_n1092));
  NAND2_X1  g667(.A1(new_n1005), .A2(new_n711), .ZN(new_n1093));
  AOI21_X1  g668(.A(new_n1081), .B1(new_n1092), .B2(new_n1093), .ZN(new_n1094));
  NAND2_X1  g669(.A1(G303), .A2(G8), .ZN(new_n1095));
  INV_X1    g670(.A(KEYINPUT55), .ZN(new_n1096));
  NAND2_X1  g671(.A1(new_n1095), .A2(new_n1096), .ZN(new_n1097));
  NAND3_X1  g672(.A1(G303), .A2(KEYINPUT55), .A3(G8), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n1097), .A2(new_n1098), .ZN(new_n1099));
  OAI211_X1 g674(.A(new_n1084), .B(new_n1091), .C1(new_n1094), .C2(new_n1099), .ZN(new_n1100));
  NAND4_X1  g675(.A1(new_n997), .A2(new_n989), .A3(new_n805), .A4(new_n990), .ZN(new_n1101));
  INV_X1    g676(.A(KEYINPUT112), .ZN(new_n1102));
  OR2_X1    g677(.A1(new_n1101), .A2(new_n1102), .ZN(new_n1103));
  AOI22_X1  g678(.A1(new_n1101), .A2(new_n1102), .B1(new_n1005), .B2(new_n711), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n1103), .A2(new_n1104), .ZN(new_n1105));
  NAND3_X1  g680(.A1(new_n1105), .A2(G8), .A3(new_n1099), .ZN(new_n1106));
  INV_X1    g681(.A(KEYINPUT113), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n1106), .A2(new_n1107), .ZN(new_n1108));
  AOI21_X1  g683(.A(new_n1081), .B1(new_n1103), .B2(new_n1104), .ZN(new_n1109));
  NAND3_X1  g684(.A1(new_n1109), .A2(KEYINPUT113), .A3(new_n1099), .ZN(new_n1110));
  AOI21_X1  g685(.A(new_n1100), .B1(new_n1108), .B2(new_n1110), .ZN(new_n1111));
  INV_X1    g686(.A(G1966), .ZN(new_n1112));
  NAND2_X1  g687(.A1(new_n1005), .A2(new_n1112), .ZN(new_n1113));
  NAND4_X1  g688(.A1(new_n997), .A2(new_n989), .A3(new_n762), .A4(new_n990), .ZN(new_n1114));
  AOI211_X1 g689(.A(new_n1081), .B(G168), .C1(new_n1113), .C2(new_n1114), .ZN(new_n1115));
  NAND3_X1  g690(.A1(new_n1113), .A2(G168), .A3(new_n1114), .ZN(new_n1116));
  AOI21_X1  g691(.A(KEYINPUT51), .B1(new_n1116), .B2(G8), .ZN(new_n1117));
  INV_X1    g692(.A(KEYINPUT123), .ZN(new_n1118));
  AOI21_X1  g693(.A(new_n1115), .B1(new_n1117), .B2(new_n1118), .ZN(new_n1119));
  OR2_X1    g694(.A1(new_n1117), .A2(new_n1118), .ZN(new_n1120));
  AND3_X1   g695(.A1(new_n1116), .A2(KEYINPUT51), .A3(G8), .ZN(new_n1121));
  OAI21_X1  g696(.A(new_n1119), .B1(new_n1120), .B2(new_n1121), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n1111), .A2(new_n1122), .ZN(new_n1123));
  INV_X1    g698(.A(new_n1011), .ZN(new_n1124));
  NAND4_X1  g699(.A1(new_n1124), .A2(G301), .A3(new_n1008), .A4(new_n1009), .ZN(new_n1125));
  OR2_X1    g700(.A1(new_n1125), .A2(KEYINPUT127), .ZN(new_n1126));
  NAND2_X1  g701(.A1(new_n1016), .A2(G171), .ZN(new_n1127));
  NAND2_X1  g702(.A1(new_n1127), .A2(KEYINPUT54), .ZN(new_n1128));
  AOI21_X1  g703(.A(new_n1128), .B1(new_n1125), .B2(KEYINPUT127), .ZN(new_n1129));
  AOI21_X1  g704(.A(new_n1123), .B1(new_n1126), .B2(new_n1129), .ZN(new_n1130));
  NAND4_X1  g705(.A1(new_n1021), .A2(new_n1023), .A3(new_n1073), .A4(new_n1130), .ZN(new_n1131));
  INV_X1    g706(.A(KEYINPUT63), .ZN(new_n1132));
  NAND2_X1  g707(.A1(new_n1092), .A2(new_n1093), .ZN(new_n1133));
  AOI21_X1  g708(.A(new_n1099), .B1(new_n1133), .B2(G8), .ZN(new_n1134));
  NAND2_X1  g709(.A1(new_n1084), .A2(new_n1091), .ZN(new_n1135));
  NOR2_X1   g710(.A1(new_n1134), .A2(new_n1135), .ZN(new_n1136));
  AOI211_X1 g711(.A(new_n1081), .B(G286), .C1(new_n1113), .C2(new_n1114), .ZN(new_n1137));
  INV_X1    g712(.A(new_n1110), .ZN(new_n1138));
  AOI21_X1  g713(.A(KEYINPUT113), .B1(new_n1109), .B2(new_n1099), .ZN(new_n1139));
  OAI211_X1 g714(.A(new_n1136), .B(new_n1137), .C1(new_n1138), .C2(new_n1139), .ZN(new_n1140));
  OAI21_X1  g715(.A(new_n1132), .B1(new_n1140), .B2(KEYINPUT116), .ZN(new_n1141));
  INV_X1    g716(.A(KEYINPUT116), .ZN(new_n1142));
  AOI21_X1  g717(.A(new_n1142), .B1(new_n1111), .B2(new_n1137), .ZN(new_n1143));
  OAI21_X1  g718(.A(KEYINPUT117), .B1(new_n1141), .B2(new_n1143), .ZN(new_n1144));
  NAND2_X1  g719(.A1(new_n1140), .A2(KEYINPUT116), .ZN(new_n1145));
  NAND3_X1  g720(.A1(new_n1111), .A2(new_n1142), .A3(new_n1137), .ZN(new_n1146));
  INV_X1    g721(.A(KEYINPUT117), .ZN(new_n1147));
  NAND4_X1  g722(.A1(new_n1145), .A2(new_n1146), .A3(new_n1147), .A4(new_n1132), .ZN(new_n1148));
  NAND2_X1  g723(.A1(new_n1108), .A2(new_n1110), .ZN(new_n1149));
  AND4_X1   g724(.A1(KEYINPUT63), .A2(new_n1084), .A3(new_n1091), .A4(new_n1137), .ZN(new_n1150));
  OAI211_X1 g725(.A(new_n1149), .B(new_n1150), .C1(new_n1099), .C2(new_n1109), .ZN(new_n1151));
  NAND3_X1  g726(.A1(new_n1144), .A2(new_n1148), .A3(new_n1151), .ZN(new_n1152));
  AND3_X1   g727(.A1(new_n1084), .A2(new_n1089), .A3(new_n928), .ZN(new_n1153));
  NOR2_X1   g728(.A1(G305), .A2(G1981), .ZN(new_n1154));
  OAI21_X1  g729(.A(new_n1082), .B1(new_n1153), .B2(new_n1154), .ZN(new_n1155));
  OAI21_X1  g730(.A(new_n1155), .B1(new_n1149), .B2(new_n1135), .ZN(new_n1156));
  XOR2_X1   g731(.A(new_n1122), .B(KEYINPUT62), .Z(new_n1157));
  INV_X1    g732(.A(new_n1111), .ZN(new_n1158));
  AOI21_X1  g733(.A(new_n1158), .B1(new_n1015), .B2(new_n1014), .ZN(new_n1159));
  AOI21_X1  g734(.A(new_n1156), .B1(new_n1157), .B2(new_n1159), .ZN(new_n1160));
  NAND3_X1  g735(.A1(new_n1131), .A2(new_n1152), .A3(new_n1160), .ZN(new_n1161));
  NAND2_X1  g736(.A1(new_n738), .A2(G2067), .ZN(new_n1162));
  NAND3_X1  g737(.A1(new_n730), .A2(new_n1042), .A3(new_n737), .ZN(new_n1163));
  NAND2_X1  g738(.A1(new_n1162), .A2(new_n1163), .ZN(new_n1164));
  XNOR2_X1  g739(.A(new_n1164), .B(KEYINPUT110), .ZN(new_n1165));
  INV_X1    g740(.A(G1996), .ZN(new_n1166));
  OAI21_X1  g741(.A(new_n1165), .B1(new_n1166), .B2(new_n887), .ZN(new_n1167));
  NOR2_X1   g742(.A1(new_n1003), .A2(new_n991), .ZN(new_n1168));
  XOR2_X1   g743(.A(new_n1168), .B(KEYINPUT109), .Z(new_n1169));
  NAND2_X1  g744(.A1(new_n1167), .A2(new_n1169), .ZN(new_n1170));
  AND2_X1   g745(.A1(new_n695), .A2(new_n702), .ZN(new_n1171));
  NOR2_X1   g746(.A1(new_n695), .A2(new_n702), .ZN(new_n1172));
  OAI21_X1  g747(.A(new_n1169), .B1(new_n1171), .B2(new_n1172), .ZN(new_n1173));
  INV_X1    g748(.A(new_n1168), .ZN(new_n1174));
  NOR2_X1   g749(.A1(new_n1174), .A2(G1996), .ZN(new_n1175));
  NAND2_X1  g750(.A1(new_n817), .A2(new_n1175), .ZN(new_n1176));
  NAND3_X1  g751(.A1(new_n1170), .A2(new_n1173), .A3(new_n1176), .ZN(new_n1177));
  XNOR2_X1  g752(.A(G290), .B(G1986), .ZN(new_n1178));
  AOI21_X1  g753(.A(new_n1177), .B1(new_n1168), .B2(new_n1178), .ZN(new_n1179));
  NAND2_X1  g754(.A1(new_n1161), .A2(new_n1179), .ZN(new_n1180));
  XNOR2_X1  g755(.A(new_n1175), .B(KEYINPUT46), .ZN(new_n1181));
  NAND2_X1  g756(.A1(new_n1165), .A2(new_n887), .ZN(new_n1182));
  AOI21_X1  g757(.A(new_n1181), .B1(new_n1182), .B2(new_n1169), .ZN(new_n1183));
  INV_X1    g758(.A(KEYINPUT47), .ZN(new_n1184));
  AND2_X1   g759(.A1(new_n1183), .A2(new_n1184), .ZN(new_n1185));
  NOR2_X1   g760(.A1(new_n1183), .A2(new_n1184), .ZN(new_n1186));
  NOR3_X1   g761(.A1(new_n1174), .A2(G1986), .A3(G290), .ZN(new_n1187));
  XNOR2_X1  g762(.A(new_n1187), .B(KEYINPUT48), .ZN(new_n1188));
  OAI22_X1  g763(.A1(new_n1185), .A2(new_n1186), .B1(new_n1177), .B2(new_n1188), .ZN(new_n1189));
  NAND3_X1  g764(.A1(new_n1170), .A2(new_n1171), .A3(new_n1176), .ZN(new_n1190));
  NAND2_X1  g765(.A1(new_n1190), .A2(new_n1163), .ZN(new_n1191));
  AOI21_X1  g766(.A(new_n1189), .B1(new_n1169), .B2(new_n1191), .ZN(new_n1192));
  NAND2_X1  g767(.A1(new_n1180), .A2(new_n1192), .ZN(G329));
  assign    G231 = 1'b0;
  OR2_X1    g768(.A1(G227), .A2(new_n461), .ZN(new_n1195));
  AOI211_X1 g769(.A(new_n1195), .B(G401), .C1(new_n685), .C2(new_n688), .ZN(new_n1196));
  OAI211_X1 g770(.A(new_n900), .B(new_n1196), .C1(new_n975), .C2(new_n976), .ZN(G225));
  INV_X1    g771(.A(G225), .ZN(G308));
endmodule


