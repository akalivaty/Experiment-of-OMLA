//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 0 0 1 1 0 0 1 0 0 0 0 1 1 0 1 1 1 0 0 0 0 0 0 0 1 1 1 1 1 0 1 0 1 0 0 0 0 1 0 1 0 1 0 1 0 1 1 1 1 0 0 0 0 0 0 1 0 0 0 0 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:25:00 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n697, new_n698, new_n699, new_n700, new_n701, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n714, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n726, new_n727, new_n728,
    new_n729, new_n730, new_n731, new_n732, new_n733, new_n734, new_n735,
    new_n736, new_n737, new_n738, new_n739, new_n740, new_n742, new_n743,
    new_n744, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n784, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n808, new_n809, new_n810,
    new_n811, new_n812, new_n813, new_n814, new_n815, new_n816, new_n817,
    new_n818, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n934, new_n935, new_n936, new_n937, new_n938,
    new_n939, new_n940, new_n941, new_n942, new_n943, new_n944, new_n945,
    new_n946, new_n947, new_n948, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n972, new_n973, new_n974, new_n975, new_n976,
    new_n977, new_n979, new_n980, new_n981, new_n982, new_n983, new_n984,
    new_n985, new_n986, new_n987, new_n988, new_n989, new_n990, new_n991,
    new_n992, new_n993, new_n994, new_n995, new_n996, new_n997, new_n999,
    new_n1000, new_n1001, new_n1002, new_n1003, new_n1004, new_n1005,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1022, new_n1023, new_n1024,
    new_n1025, new_n1026, new_n1027, new_n1028, new_n1029, new_n1030,
    new_n1032, new_n1033, new_n1034, new_n1035, new_n1036, new_n1037,
    new_n1038, new_n1039, new_n1040, new_n1041;
  INV_X1    g000(.A(KEYINPUT20), .ZN(new_n187));
  NOR2_X1   g001(.A1(G475), .A2(G902), .ZN(new_n188));
  XNOR2_X1  g002(.A(G113), .B(G122), .ZN(new_n189));
  XNOR2_X1  g003(.A(KEYINPUT85), .B(G104), .ZN(new_n190));
  XOR2_X1   g004(.A(new_n189), .B(new_n190), .Z(new_n191));
  INV_X1    g005(.A(new_n191), .ZN(new_n192));
  INV_X1    g006(.A(KEYINPUT65), .ZN(new_n193));
  INV_X1    g007(.A(G953), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n193), .A2(new_n194), .ZN(new_n195));
  INV_X1    g009(.A(G237), .ZN(new_n196));
  NAND2_X1  g010(.A1(KEYINPUT65), .A2(G953), .ZN(new_n197));
  NAND4_X1  g011(.A1(new_n195), .A2(G214), .A3(new_n196), .A4(new_n197), .ZN(new_n198));
  INV_X1    g012(.A(G143), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n198), .A2(new_n199), .ZN(new_n200));
  AND2_X1   g014(.A1(KEYINPUT65), .A2(G953), .ZN(new_n201));
  NOR2_X1   g015(.A1(KEYINPUT65), .A2(G953), .ZN(new_n202));
  NOR2_X1   g016(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NAND4_X1  g017(.A1(new_n203), .A2(G143), .A3(G214), .A4(new_n196), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n200), .A2(new_n204), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n205), .A2(G131), .ZN(new_n206));
  INV_X1    g020(.A(G131), .ZN(new_n207));
  NAND3_X1  g021(.A1(new_n200), .A2(new_n204), .A3(new_n207), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n206), .A2(new_n208), .ZN(new_n209));
  XNOR2_X1  g023(.A(KEYINPUT72), .B(G125), .ZN(new_n210));
  INV_X1    g024(.A(KEYINPUT16), .ZN(new_n211));
  INV_X1    g025(.A(G140), .ZN(new_n212));
  NAND3_X1  g026(.A1(new_n210), .A2(new_n211), .A3(new_n212), .ZN(new_n213));
  NOR2_X1   g027(.A1(G125), .A2(G140), .ZN(new_n214));
  AOI21_X1  g028(.A(new_n214), .B1(new_n210), .B2(G140), .ZN(new_n215));
  OAI211_X1 g029(.A(G146), .B(new_n213), .C1(new_n215), .C2(new_n211), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n215), .A2(KEYINPUT19), .ZN(new_n217));
  INV_X1    g031(.A(G146), .ZN(new_n218));
  XNOR2_X1  g032(.A(G125), .B(G140), .ZN(new_n219));
  INV_X1    g033(.A(KEYINPUT19), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  NAND3_X1  g035(.A1(new_n217), .A2(new_n218), .A3(new_n221), .ZN(new_n222));
  NAND3_X1  g036(.A1(new_n209), .A2(new_n216), .A3(new_n222), .ZN(new_n223));
  NAND2_X1  g037(.A1(KEYINPUT18), .A2(G131), .ZN(new_n224));
  XNOR2_X1  g038(.A(new_n224), .B(KEYINPUT82), .ZN(new_n225));
  NAND3_X1  g039(.A1(new_n200), .A2(new_n204), .A3(new_n225), .ZN(new_n226));
  AND2_X1   g040(.A1(KEYINPUT72), .A2(G125), .ZN(new_n227));
  NOR2_X1   g041(.A1(KEYINPUT72), .A2(G125), .ZN(new_n228));
  OAI21_X1  g042(.A(G140), .B1(new_n227), .B2(new_n228), .ZN(new_n229));
  INV_X1    g043(.A(new_n214), .ZN(new_n230));
  NAND3_X1  g044(.A1(new_n229), .A2(G146), .A3(new_n230), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n219), .A2(new_n218), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n231), .A2(new_n232), .ZN(new_n233));
  XNOR2_X1  g047(.A(new_n198), .B(G143), .ZN(new_n234));
  OAI211_X1 g048(.A(new_n226), .B(new_n233), .C1(new_n234), .C2(new_n224), .ZN(new_n235));
  INV_X1    g049(.A(KEYINPUT83), .ZN(new_n236));
  NOR2_X1   g050(.A1(new_n235), .A2(new_n236), .ZN(new_n237));
  INV_X1    g051(.A(new_n224), .ZN(new_n238));
  AOI22_X1  g052(.A1(new_n205), .A2(new_n238), .B1(new_n232), .B2(new_n231), .ZN(new_n239));
  AOI21_X1  g053(.A(KEYINPUT83), .B1(new_n239), .B2(new_n226), .ZN(new_n240));
  OAI21_X1  g054(.A(new_n223), .B1(new_n237), .B2(new_n240), .ZN(new_n241));
  INV_X1    g055(.A(KEYINPUT84), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n241), .A2(new_n242), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n235), .A2(new_n236), .ZN(new_n244));
  NAND3_X1  g058(.A1(new_n239), .A2(KEYINPUT83), .A3(new_n226), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n244), .A2(new_n245), .ZN(new_n246));
  NAND3_X1  g060(.A1(new_n246), .A2(KEYINPUT84), .A3(new_n223), .ZN(new_n247));
  AOI21_X1  g061(.A(new_n192), .B1(new_n243), .B2(new_n247), .ZN(new_n248));
  INV_X1    g062(.A(KEYINPUT17), .ZN(new_n249));
  NAND3_X1  g063(.A1(new_n206), .A2(new_n249), .A3(new_n208), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n250), .A2(KEYINPUT86), .ZN(new_n251));
  AOI21_X1  g065(.A(new_n211), .B1(new_n229), .B2(new_n230), .ZN(new_n252));
  NOR2_X1   g066(.A1(new_n227), .A2(new_n228), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n211), .A2(new_n212), .ZN(new_n254));
  NOR2_X1   g068(.A1(new_n253), .A2(new_n254), .ZN(new_n255));
  OAI21_X1  g069(.A(new_n218), .B1(new_n252), .B2(new_n255), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n256), .A2(new_n216), .ZN(new_n257));
  INV_X1    g071(.A(new_n257), .ZN(new_n258));
  INV_X1    g072(.A(KEYINPUT86), .ZN(new_n259));
  NAND4_X1  g073(.A1(new_n206), .A2(new_n259), .A3(new_n249), .A4(new_n208), .ZN(new_n260));
  NAND3_X1  g074(.A1(new_n205), .A2(KEYINPUT17), .A3(G131), .ZN(new_n261));
  NAND4_X1  g075(.A1(new_n251), .A2(new_n258), .A3(new_n260), .A4(new_n261), .ZN(new_n262));
  NAND3_X1  g076(.A1(new_n262), .A2(new_n192), .A3(new_n246), .ZN(new_n263));
  INV_X1    g077(.A(new_n263), .ZN(new_n264));
  OAI211_X1 g078(.A(new_n187), .B(new_n188), .C1(new_n248), .C2(new_n264), .ZN(new_n265));
  INV_X1    g079(.A(new_n188), .ZN(new_n266));
  AND3_X1   g080(.A1(new_n246), .A2(KEYINPUT84), .A3(new_n223), .ZN(new_n267));
  AOI21_X1  g081(.A(KEYINPUT84), .B1(new_n246), .B2(new_n223), .ZN(new_n268));
  OAI21_X1  g082(.A(new_n191), .B1(new_n267), .B2(new_n268), .ZN(new_n269));
  AOI21_X1  g083(.A(new_n266), .B1(new_n269), .B2(new_n263), .ZN(new_n270));
  XOR2_X1   g084(.A(KEYINPUT81), .B(KEYINPUT20), .Z(new_n271));
  OAI21_X1  g085(.A(new_n265), .B1(new_n270), .B2(new_n271), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n262), .A2(new_n246), .ZN(new_n273));
  NOR2_X1   g087(.A1(new_n192), .A2(KEYINPUT87), .ZN(new_n274));
  INV_X1    g088(.A(new_n274), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n273), .A2(new_n275), .ZN(new_n276));
  INV_X1    g090(.A(G902), .ZN(new_n277));
  NAND3_X1  g091(.A1(new_n262), .A2(new_n246), .A3(new_n274), .ZN(new_n278));
  NAND3_X1  g092(.A1(new_n276), .A2(new_n277), .A3(new_n278), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n279), .A2(G475), .ZN(new_n280));
  INV_X1    g094(.A(G116), .ZN(new_n281));
  OAI21_X1  g095(.A(KEYINPUT14), .B1(new_n281), .B2(G122), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n282), .A2(G107), .ZN(new_n283));
  XNOR2_X1  g097(.A(G116), .B(G122), .ZN(new_n284));
  OR2_X1    g098(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n283), .A2(new_n284), .ZN(new_n286));
  INV_X1    g100(.A(KEYINPUT88), .ZN(new_n287));
  OAI21_X1  g101(.A(new_n287), .B1(new_n199), .B2(G128), .ZN(new_n288));
  INV_X1    g102(.A(G128), .ZN(new_n289));
  NAND3_X1  g103(.A1(new_n289), .A2(KEYINPUT88), .A3(G143), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n288), .A2(new_n290), .ZN(new_n291));
  INV_X1    g105(.A(G134), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n199), .A2(G128), .ZN(new_n293));
  NAND3_X1  g107(.A1(new_n291), .A2(new_n292), .A3(new_n293), .ZN(new_n294));
  INV_X1    g108(.A(new_n294), .ZN(new_n295));
  AOI21_X1  g109(.A(new_n292), .B1(new_n291), .B2(new_n293), .ZN(new_n296));
  OAI211_X1 g110(.A(new_n285), .B(new_n286), .C1(new_n295), .C2(new_n296), .ZN(new_n297));
  INV_X1    g111(.A(KEYINPUT13), .ZN(new_n298));
  AOI22_X1  g112(.A1(new_n288), .A2(new_n290), .B1(new_n293), .B2(new_n298), .ZN(new_n299));
  INV_X1    g113(.A(new_n293), .ZN(new_n300));
  AOI22_X1  g114(.A1(new_n299), .A2(KEYINPUT89), .B1(KEYINPUT13), .B2(new_n300), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n293), .A2(new_n298), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n291), .A2(new_n302), .ZN(new_n303));
  INV_X1    g117(.A(KEYINPUT89), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  AOI21_X1  g119(.A(new_n292), .B1(new_n301), .B2(new_n305), .ZN(new_n306));
  OR2_X1    g120(.A1(new_n284), .A2(G107), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n284), .A2(G107), .ZN(new_n308));
  NAND3_X1  g122(.A1(new_n307), .A2(new_n294), .A3(new_n308), .ZN(new_n309));
  OAI21_X1  g123(.A(new_n297), .B1(new_n306), .B2(new_n309), .ZN(new_n310));
  XNOR2_X1  g124(.A(KEYINPUT9), .B(G234), .ZN(new_n311));
  INV_X1    g125(.A(G217), .ZN(new_n312));
  NOR3_X1   g126(.A1(new_n311), .A2(new_n312), .A3(G953), .ZN(new_n313));
  INV_X1    g127(.A(new_n313), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n310), .A2(new_n314), .ZN(new_n315));
  OAI211_X1 g129(.A(new_n297), .B(new_n313), .C1(new_n306), .C2(new_n309), .ZN(new_n316));
  AOI21_X1  g130(.A(G902), .B1(new_n315), .B2(new_n316), .ZN(new_n317));
  INV_X1    g131(.A(new_n317), .ZN(new_n318));
  INV_X1    g132(.A(G478), .ZN(new_n319));
  NOR2_X1   g133(.A1(new_n319), .A2(KEYINPUT15), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n318), .A2(new_n320), .ZN(new_n321));
  OAI21_X1  g135(.A(new_n317), .B1(KEYINPUT15), .B2(new_n319), .ZN(new_n322));
  INV_X1    g136(.A(G952), .ZN(new_n323));
  NOR2_X1   g137(.A1(new_n323), .A2(G953), .ZN(new_n324));
  INV_X1    g138(.A(G234), .ZN(new_n325));
  OAI21_X1  g139(.A(new_n324), .B1(new_n325), .B2(new_n196), .ZN(new_n326));
  INV_X1    g140(.A(new_n326), .ZN(new_n327));
  AOI211_X1 g141(.A(new_n277), .B(new_n203), .C1(G234), .C2(G237), .ZN(new_n328));
  XNOR2_X1  g142(.A(KEYINPUT21), .B(G898), .ZN(new_n329));
  AOI21_X1  g143(.A(new_n327), .B1(new_n328), .B2(new_n329), .ZN(new_n330));
  INV_X1    g144(.A(new_n330), .ZN(new_n331));
  NAND3_X1  g145(.A1(new_n321), .A2(new_n322), .A3(new_n331), .ZN(new_n332));
  INV_X1    g146(.A(new_n332), .ZN(new_n333));
  NAND3_X1  g147(.A1(new_n272), .A2(new_n280), .A3(new_n333), .ZN(new_n334));
  XOR2_X1   g148(.A(G110), .B(G140), .Z(new_n335));
  XNOR2_X1  g149(.A(new_n335), .B(KEYINPUT74), .ZN(new_n336));
  AND2_X1   g150(.A1(new_n203), .A2(G227), .ZN(new_n337));
  XNOR2_X1  g151(.A(new_n336), .B(new_n337), .ZN(new_n338));
  INV_X1    g152(.A(KEYINPUT11), .ZN(new_n339));
  OAI21_X1  g153(.A(new_n339), .B1(new_n292), .B2(G137), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n292), .A2(G137), .ZN(new_n341));
  INV_X1    g155(.A(G137), .ZN(new_n342));
  NAND3_X1  g156(.A1(new_n342), .A2(KEYINPUT11), .A3(G134), .ZN(new_n343));
  NAND3_X1  g157(.A1(new_n340), .A2(new_n341), .A3(new_n343), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n344), .A2(G131), .ZN(new_n345));
  NAND4_X1  g159(.A1(new_n340), .A2(new_n343), .A3(new_n207), .A4(new_n341), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n345), .A2(new_n346), .ZN(new_n347));
  INV_X1    g161(.A(new_n347), .ZN(new_n348));
  INV_X1    g162(.A(G104), .ZN(new_n349));
  OAI21_X1  g163(.A(KEYINPUT3), .B1(new_n349), .B2(G107), .ZN(new_n350));
  INV_X1    g164(.A(KEYINPUT3), .ZN(new_n351));
  INV_X1    g165(.A(G107), .ZN(new_n352));
  NAND3_X1  g166(.A1(new_n351), .A2(new_n352), .A3(G104), .ZN(new_n353));
  INV_X1    g167(.A(G101), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n349), .A2(G107), .ZN(new_n355));
  NAND4_X1  g169(.A1(new_n350), .A2(new_n353), .A3(new_n354), .A4(new_n355), .ZN(new_n356));
  NOR2_X1   g170(.A1(new_n349), .A2(G107), .ZN(new_n357));
  NOR2_X1   g171(.A1(new_n352), .A2(G104), .ZN(new_n358));
  OAI21_X1  g172(.A(G101), .B1(new_n357), .B2(new_n358), .ZN(new_n359));
  INV_X1    g173(.A(KEYINPUT1), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n218), .A2(G143), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n199), .A2(G146), .ZN(new_n362));
  AND4_X1   g176(.A1(new_n360), .A2(new_n361), .A3(new_n362), .A4(G128), .ZN(new_n363));
  OAI21_X1  g177(.A(KEYINPUT1), .B1(new_n199), .B2(G146), .ZN(new_n364));
  AOI22_X1  g178(.A1(new_n364), .A2(G128), .B1(new_n361), .B2(new_n362), .ZN(new_n365));
  OAI211_X1 g179(.A(new_n356), .B(new_n359), .C1(new_n363), .C2(new_n365), .ZN(new_n366));
  INV_X1    g180(.A(KEYINPUT75), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n366), .A2(new_n367), .ZN(new_n368));
  INV_X1    g182(.A(KEYINPUT10), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n368), .A2(new_n369), .ZN(new_n370));
  NAND3_X1  g184(.A1(new_n366), .A2(new_n367), .A3(KEYINPUT10), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  NAND3_X1  g186(.A1(new_n350), .A2(new_n353), .A3(new_n355), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n373), .A2(G101), .ZN(new_n374));
  NAND3_X1  g188(.A1(new_n374), .A2(KEYINPUT4), .A3(new_n356), .ZN(new_n375));
  NOR2_X1   g189(.A1(KEYINPUT0), .A2(G128), .ZN(new_n376));
  XNOR2_X1  g190(.A(G143), .B(G146), .ZN(new_n377));
  NAND2_X1  g191(.A1(KEYINPUT0), .A2(G128), .ZN(new_n378));
  AOI21_X1  g192(.A(new_n376), .B1(new_n377), .B2(new_n378), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n361), .A2(new_n362), .ZN(new_n380));
  NAND3_X1  g194(.A1(new_n380), .A2(KEYINPUT0), .A3(G128), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n379), .A2(new_n381), .ZN(new_n382));
  INV_X1    g196(.A(KEYINPUT4), .ZN(new_n383));
  NAND3_X1  g197(.A1(new_n373), .A2(new_n383), .A3(G101), .ZN(new_n384));
  NAND3_X1  g198(.A1(new_n375), .A2(new_n382), .A3(new_n384), .ZN(new_n385));
  AOI21_X1  g199(.A(new_n348), .B1(new_n372), .B2(new_n385), .ZN(new_n386));
  AND3_X1   g200(.A1(new_n366), .A2(new_n367), .A3(KEYINPUT10), .ZN(new_n387));
  AOI21_X1  g201(.A(KEYINPUT10), .B1(new_n366), .B2(new_n367), .ZN(new_n388));
  OAI211_X1 g202(.A(new_n348), .B(new_n385), .C1(new_n387), .C2(new_n388), .ZN(new_n389));
  INV_X1    g203(.A(new_n389), .ZN(new_n390));
  OAI21_X1  g204(.A(new_n338), .B1(new_n386), .B2(new_n390), .ZN(new_n391));
  NOR2_X1   g205(.A1(new_n363), .A2(new_n365), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n356), .A2(new_n359), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n392), .A2(new_n393), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n394), .A2(new_n366), .ZN(new_n395));
  AND3_X1   g209(.A1(new_n395), .A2(KEYINPUT12), .A3(new_n347), .ZN(new_n396));
  AOI21_X1  g210(.A(KEYINPUT12), .B1(new_n395), .B2(new_n347), .ZN(new_n397));
  OR2_X1    g211(.A1(new_n396), .A2(new_n397), .ZN(new_n398));
  INV_X1    g212(.A(new_n338), .ZN(new_n399));
  NAND3_X1  g213(.A1(new_n389), .A2(KEYINPUT76), .A3(new_n399), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n398), .A2(new_n400), .ZN(new_n401));
  AOI21_X1  g215(.A(KEYINPUT76), .B1(new_n389), .B2(new_n399), .ZN(new_n402));
  OAI21_X1  g216(.A(new_n391), .B1(new_n401), .B2(new_n402), .ZN(new_n403));
  INV_X1    g217(.A(G469), .ZN(new_n404));
  NAND3_X1  g218(.A1(new_n403), .A2(new_n404), .A3(new_n277), .ZN(new_n405));
  OAI21_X1  g219(.A(new_n385), .B1(new_n387), .B2(new_n388), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n406), .A2(new_n347), .ZN(new_n407));
  AND2_X1   g221(.A1(new_n389), .A2(new_n399), .ZN(new_n408));
  OAI21_X1  g222(.A(new_n389), .B1(new_n396), .B2(new_n397), .ZN(new_n409));
  AOI22_X1  g223(.A1(new_n407), .A2(new_n408), .B1(new_n409), .B2(new_n338), .ZN(new_n410));
  OAI21_X1  g224(.A(G469), .B1(new_n410), .B2(G902), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n405), .A2(new_n411), .ZN(new_n412));
  XNOR2_X1  g226(.A(G110), .B(G122), .ZN(new_n413));
  INV_X1    g227(.A(G119), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n414), .A2(G116), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n281), .A2(G119), .ZN(new_n416));
  NAND3_X1  g230(.A1(new_n415), .A2(new_n416), .A3(KEYINPUT5), .ZN(new_n417));
  OR3_X1    g231(.A1(new_n281), .A2(KEYINPUT5), .A3(G119), .ZN(new_n418));
  NAND3_X1  g232(.A1(new_n417), .A2(new_n418), .A3(G113), .ZN(new_n419));
  NAND2_X1  g233(.A1(KEYINPUT2), .A2(G113), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n420), .A2(KEYINPUT64), .ZN(new_n421));
  INV_X1    g235(.A(KEYINPUT64), .ZN(new_n422));
  NAND3_X1  g236(.A1(new_n422), .A2(KEYINPUT2), .A3(G113), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n421), .A2(new_n423), .ZN(new_n424));
  OR2_X1    g238(.A1(KEYINPUT2), .A2(G113), .ZN(new_n425));
  XNOR2_X1  g239(.A(G116), .B(G119), .ZN(new_n426));
  NAND3_X1  g240(.A1(new_n424), .A2(new_n425), .A3(new_n426), .ZN(new_n427));
  NAND4_X1  g241(.A1(new_n419), .A2(new_n427), .A3(new_n356), .A4(new_n359), .ZN(new_n428));
  AND3_X1   g242(.A1(new_n424), .A2(new_n425), .A3(new_n426), .ZN(new_n429));
  AOI21_X1  g243(.A(new_n426), .B1(new_n424), .B2(new_n425), .ZN(new_n430));
  OAI21_X1  g244(.A(new_n384), .B1(new_n429), .B2(new_n430), .ZN(new_n431));
  AND3_X1   g245(.A1(new_n374), .A2(KEYINPUT4), .A3(new_n356), .ZN(new_n432));
  OAI211_X1 g246(.A(new_n413), .B(new_n428), .C1(new_n431), .C2(new_n432), .ZN(new_n433));
  XNOR2_X1  g247(.A(new_n413), .B(KEYINPUT8), .ZN(new_n434));
  AND4_X1   g248(.A1(new_n427), .A2(new_n419), .A3(new_n356), .A4(new_n359), .ZN(new_n435));
  AOI22_X1  g249(.A1(new_n419), .A2(new_n427), .B1(new_n356), .B2(new_n359), .ZN(new_n436));
  OAI21_X1  g250(.A(new_n434), .B1(new_n435), .B2(new_n436), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n382), .A2(new_n210), .ZN(new_n438));
  OAI21_X1  g252(.A(new_n253), .B1(new_n363), .B2(new_n365), .ZN(new_n439));
  INV_X1    g253(.A(KEYINPUT7), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n194), .A2(G224), .ZN(new_n441));
  XNOR2_X1  g255(.A(new_n441), .B(KEYINPUT79), .ZN(new_n442));
  OAI211_X1 g256(.A(new_n438), .B(new_n439), .C1(new_n440), .C2(new_n442), .ZN(new_n443));
  NOR2_X1   g257(.A1(new_n442), .A2(new_n440), .ZN(new_n444));
  AOI21_X1  g258(.A(new_n253), .B1(new_n379), .B2(new_n381), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n364), .A2(G128), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n446), .A2(new_n380), .ZN(new_n447));
  NAND3_X1  g261(.A1(new_n377), .A2(G128), .A3(new_n364), .ZN(new_n448));
  AOI21_X1  g262(.A(new_n210), .B1(new_n447), .B2(new_n448), .ZN(new_n449));
  OAI21_X1  g263(.A(new_n444), .B1(new_n445), .B2(new_n449), .ZN(new_n450));
  NAND4_X1  g264(.A1(new_n433), .A2(new_n437), .A3(new_n443), .A4(new_n450), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n451), .A2(new_n277), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n452), .A2(KEYINPUT80), .ZN(new_n453));
  OAI21_X1  g267(.A(new_n428), .B1(new_n431), .B2(new_n432), .ZN(new_n454));
  INV_X1    g268(.A(new_n413), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  INV_X1    g270(.A(KEYINPUT78), .ZN(new_n457));
  INV_X1    g271(.A(KEYINPUT6), .ZN(new_n458));
  NOR2_X1   g272(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  NAND3_X1  g273(.A1(new_n456), .A2(new_n433), .A3(new_n459), .ZN(new_n460));
  OAI211_X1 g274(.A(new_n454), .B(new_n455), .C1(new_n457), .C2(new_n458), .ZN(new_n461));
  NOR2_X1   g275(.A1(new_n445), .A2(new_n449), .ZN(new_n462));
  XNOR2_X1  g276(.A(new_n462), .B(new_n442), .ZN(new_n463));
  NAND3_X1  g277(.A1(new_n460), .A2(new_n461), .A3(new_n463), .ZN(new_n464));
  INV_X1    g278(.A(KEYINPUT80), .ZN(new_n465));
  NAND3_X1  g279(.A1(new_n451), .A2(new_n465), .A3(new_n277), .ZN(new_n466));
  NAND3_X1  g280(.A1(new_n453), .A2(new_n464), .A3(new_n466), .ZN(new_n467));
  OAI21_X1  g281(.A(G210), .B1(G237), .B2(G902), .ZN(new_n468));
  INV_X1    g282(.A(new_n468), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n467), .A2(new_n469), .ZN(new_n470));
  NAND4_X1  g284(.A1(new_n453), .A2(new_n464), .A3(new_n468), .A4(new_n466), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  OAI21_X1  g286(.A(G214), .B1(G237), .B2(G902), .ZN(new_n473));
  XNOR2_X1  g287(.A(new_n473), .B(KEYINPUT77), .ZN(new_n474));
  OAI21_X1  g288(.A(G221), .B1(new_n311), .B2(G902), .ZN(new_n475));
  NAND4_X1  g289(.A1(new_n412), .A2(new_n472), .A3(new_n474), .A4(new_n475), .ZN(new_n476));
  NOR2_X1   g290(.A1(new_n334), .A2(new_n476), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n347), .A2(new_n382), .ZN(new_n478));
  NOR2_X1   g292(.A1(new_n429), .A2(new_n430), .ZN(new_n479));
  NOR2_X1   g293(.A1(new_n292), .A2(G137), .ZN(new_n480));
  NOR2_X1   g294(.A1(new_n342), .A2(G134), .ZN(new_n481));
  OAI21_X1  g295(.A(G131), .B1(new_n480), .B2(new_n481), .ZN(new_n482));
  OAI211_X1 g296(.A(new_n346), .B(new_n482), .C1(new_n363), .C2(new_n365), .ZN(new_n483));
  AND3_X1   g297(.A1(new_n478), .A2(new_n479), .A3(new_n483), .ZN(new_n484));
  AOI21_X1  g298(.A(new_n479), .B1(new_n478), .B2(new_n483), .ZN(new_n485));
  OAI21_X1  g299(.A(KEYINPUT28), .B1(new_n484), .B2(new_n485), .ZN(new_n486));
  NAND3_X1  g300(.A1(new_n478), .A2(new_n479), .A3(new_n483), .ZN(new_n487));
  INV_X1    g301(.A(KEYINPUT28), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n489), .A2(KEYINPUT66), .ZN(new_n490));
  NAND4_X1  g304(.A1(new_n195), .A2(G210), .A3(new_n196), .A4(new_n197), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n491), .A2(KEYINPUT27), .ZN(new_n492));
  INV_X1    g306(.A(KEYINPUT27), .ZN(new_n493));
  NAND4_X1  g307(.A1(new_n203), .A2(new_n493), .A3(G210), .A4(new_n196), .ZN(new_n494));
  XNOR2_X1  g308(.A(KEYINPUT26), .B(G101), .ZN(new_n495));
  AND3_X1   g309(.A1(new_n492), .A2(new_n494), .A3(new_n495), .ZN(new_n496));
  AOI21_X1  g310(.A(new_n495), .B1(new_n492), .B2(new_n494), .ZN(new_n497));
  NOR2_X1   g311(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  INV_X1    g312(.A(KEYINPUT66), .ZN(new_n499));
  NAND3_X1  g313(.A1(new_n487), .A2(new_n499), .A3(new_n488), .ZN(new_n500));
  NAND4_X1  g314(.A1(new_n486), .A2(new_n490), .A3(new_n498), .A4(new_n500), .ZN(new_n501));
  INV_X1    g315(.A(KEYINPUT29), .ZN(new_n502));
  OR2_X1    g316(.A1(new_n496), .A2(new_n497), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n346), .A2(new_n482), .ZN(new_n504));
  NOR2_X1   g318(.A1(new_n392), .A2(new_n504), .ZN(new_n505));
  AOI22_X1  g319(.A1(new_n346), .A2(new_n345), .B1(new_n379), .B2(new_n381), .ZN(new_n506));
  OAI21_X1  g320(.A(KEYINPUT30), .B1(new_n505), .B2(new_n506), .ZN(new_n507));
  INV_X1    g321(.A(KEYINPUT30), .ZN(new_n508));
  NAND3_X1  g322(.A1(new_n478), .A2(new_n508), .A3(new_n483), .ZN(new_n509));
  AOI21_X1  g323(.A(new_n479), .B1(new_n507), .B2(new_n509), .ZN(new_n510));
  OAI21_X1  g324(.A(new_n503), .B1(new_n510), .B2(new_n484), .ZN(new_n511));
  NAND3_X1  g325(.A1(new_n501), .A2(new_n502), .A3(new_n511), .ZN(new_n512));
  NOR2_X1   g326(.A1(new_n503), .A2(new_n502), .ZN(new_n513));
  NAND4_X1  g327(.A1(new_n486), .A2(new_n490), .A3(new_n500), .A4(new_n513), .ZN(new_n514));
  INV_X1    g328(.A(KEYINPUT69), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  OR2_X1    g330(.A1(new_n429), .A2(new_n430), .ZN(new_n517));
  OAI21_X1  g331(.A(new_n517), .B1(new_n505), .B2(new_n506), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n518), .A2(new_n487), .ZN(new_n519));
  AOI22_X1  g333(.A1(new_n519), .A2(KEYINPUT28), .B1(new_n489), .B2(KEYINPUT66), .ZN(new_n520));
  NAND4_X1  g334(.A1(new_n520), .A2(KEYINPUT69), .A3(new_n500), .A4(new_n513), .ZN(new_n521));
  NAND4_X1  g335(.A1(new_n512), .A2(new_n516), .A3(new_n277), .A4(new_n521), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n522), .A2(G472), .ZN(new_n523));
  INV_X1    g337(.A(KEYINPUT70), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  NAND3_X1  g339(.A1(new_n522), .A2(KEYINPUT70), .A3(G472), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  NOR2_X1   g341(.A1(G472), .A2(G902), .ZN(new_n528));
  INV_X1    g342(.A(new_n528), .ZN(new_n529));
  INV_X1    g343(.A(KEYINPUT31), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n487), .A2(new_n498), .ZN(new_n531));
  OAI21_X1  g345(.A(new_n530), .B1(new_n510), .B2(new_n531), .ZN(new_n532));
  AND3_X1   g346(.A1(new_n478), .A2(new_n508), .A3(new_n483), .ZN(new_n533));
  AOI21_X1  g347(.A(new_n508), .B1(new_n478), .B2(new_n483), .ZN(new_n534));
  OAI21_X1  g348(.A(new_n517), .B1(new_n533), .B2(new_n534), .ZN(new_n535));
  INV_X1    g349(.A(new_n531), .ZN(new_n536));
  NAND3_X1  g350(.A1(new_n535), .A2(KEYINPUT31), .A3(new_n536), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n532), .A2(new_n537), .ZN(new_n538));
  NAND3_X1  g352(.A1(new_n486), .A2(new_n490), .A3(new_n500), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n539), .A2(new_n503), .ZN(new_n540));
  AOI21_X1  g354(.A(new_n529), .B1(new_n538), .B2(new_n540), .ZN(new_n541));
  AOI21_X1  g355(.A(KEYINPUT71), .B1(new_n541), .B2(KEYINPUT32), .ZN(new_n542));
  INV_X1    g356(.A(new_n542), .ZN(new_n543));
  NAND3_X1  g357(.A1(new_n541), .A2(KEYINPUT71), .A3(KEYINPUT32), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  INV_X1    g359(.A(KEYINPUT68), .ZN(new_n546));
  XOR2_X1   g360(.A(KEYINPUT67), .B(KEYINPUT32), .Z(new_n547));
  OAI21_X1  g361(.A(new_n546), .B1(new_n541), .B2(new_n547), .ZN(new_n548));
  INV_X1    g362(.A(new_n547), .ZN(new_n549));
  AOI22_X1  g363(.A1(new_n532), .A2(new_n537), .B1(new_n539), .B2(new_n503), .ZN(new_n550));
  OAI211_X1 g364(.A(KEYINPUT68), .B(new_n549), .C1(new_n550), .C2(new_n529), .ZN(new_n551));
  AND2_X1   g365(.A1(new_n548), .A2(new_n551), .ZN(new_n552));
  NAND3_X1  g366(.A1(new_n527), .A2(new_n545), .A3(new_n552), .ZN(new_n553));
  INV_X1    g367(.A(KEYINPUT23), .ZN(new_n554));
  OAI21_X1  g368(.A(new_n554), .B1(new_n414), .B2(G128), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n414), .A2(G128), .ZN(new_n556));
  NAND3_X1  g370(.A1(new_n289), .A2(KEYINPUT23), .A3(G119), .ZN(new_n557));
  NAND3_X1  g371(.A1(new_n555), .A2(new_n556), .A3(new_n557), .ZN(new_n558));
  NOR2_X1   g372(.A1(new_n558), .A2(G110), .ZN(new_n559));
  XOR2_X1   g373(.A(KEYINPUT24), .B(G110), .Z(new_n560));
  XNOR2_X1  g374(.A(G119), .B(G128), .ZN(new_n561));
  NOR2_X1   g375(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  OAI211_X1 g376(.A(new_n216), .B(new_n232), .C1(new_n559), .C2(new_n562), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n558), .A2(G110), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n560), .A2(new_n561), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  INV_X1    g380(.A(new_n566), .ZN(new_n567));
  AOI21_X1  g381(.A(KEYINPUT73), .B1(new_n257), .B2(new_n567), .ZN(new_n568));
  INV_X1    g382(.A(KEYINPUT73), .ZN(new_n569));
  AOI211_X1 g383(.A(new_n569), .B(new_n566), .C1(new_n256), .C2(new_n216), .ZN(new_n570));
  OAI21_X1  g384(.A(new_n563), .B1(new_n568), .B2(new_n570), .ZN(new_n571));
  NAND3_X1  g385(.A1(new_n203), .A2(G221), .A3(G234), .ZN(new_n572));
  XNOR2_X1  g386(.A(KEYINPUT22), .B(G137), .ZN(new_n573));
  XNOR2_X1  g387(.A(new_n572), .B(new_n573), .ZN(new_n574));
  INV_X1    g388(.A(new_n574), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n571), .A2(new_n575), .ZN(new_n576));
  OAI211_X1 g390(.A(new_n563), .B(new_n574), .C1(new_n568), .C2(new_n570), .ZN(new_n577));
  AOI21_X1  g391(.A(new_n312), .B1(G234), .B2(new_n277), .ZN(new_n578));
  NOR2_X1   g392(.A1(new_n578), .A2(G902), .ZN(new_n579));
  AND3_X1   g393(.A1(new_n576), .A2(new_n577), .A3(new_n579), .ZN(new_n580));
  NAND3_X1  g394(.A1(new_n576), .A2(new_n277), .A3(new_n577), .ZN(new_n581));
  INV_X1    g395(.A(KEYINPUT25), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  NAND4_X1  g397(.A1(new_n576), .A2(KEYINPUT25), .A3(new_n277), .A4(new_n577), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  AOI21_X1  g399(.A(new_n580), .B1(new_n585), .B2(new_n578), .ZN(new_n586));
  NAND3_X1  g400(.A1(new_n477), .A2(new_n553), .A3(new_n586), .ZN(new_n587));
  XNOR2_X1  g401(.A(KEYINPUT90), .B(G101), .ZN(new_n588));
  XNOR2_X1  g402(.A(new_n587), .B(new_n588), .ZN(G3));
  INV_X1    g403(.A(KEYINPUT91), .ZN(new_n590));
  AOI21_X1  g404(.A(new_n590), .B1(new_n472), .B2(new_n473), .ZN(new_n591));
  INV_X1    g405(.A(new_n473), .ZN(new_n592));
  AOI211_X1 g406(.A(KEYINPUT91), .B(new_n592), .C1(new_n470), .C2(new_n471), .ZN(new_n593));
  NOR2_X1   g407(.A1(new_n591), .A2(new_n593), .ZN(new_n594));
  NOR2_X1   g408(.A1(new_n319), .A2(G902), .ZN(new_n595));
  INV_X1    g409(.A(new_n316), .ZN(new_n596));
  NAND3_X1  g410(.A1(new_n291), .A2(KEYINPUT89), .A3(new_n302), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n300), .A2(KEYINPUT13), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  NOR2_X1   g413(.A1(new_n299), .A2(KEYINPUT89), .ZN(new_n600));
  OAI21_X1  g414(.A(G134), .B1(new_n599), .B2(new_n600), .ZN(new_n601));
  INV_X1    g415(.A(new_n309), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  AOI21_X1  g417(.A(new_n313), .B1(new_n603), .B2(new_n297), .ZN(new_n604));
  OAI21_X1  g418(.A(KEYINPUT92), .B1(new_n596), .B2(new_n604), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n310), .A2(KEYINPUT33), .ZN(new_n606));
  INV_X1    g420(.A(KEYINPUT33), .ZN(new_n607));
  AND2_X1   g421(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  NOR2_X1   g422(.A1(new_n605), .A2(new_n608), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n606), .A2(new_n607), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n315), .A2(new_n316), .ZN(new_n611));
  AOI21_X1  g425(.A(new_n610), .B1(KEYINPUT92), .B2(new_n611), .ZN(new_n612));
  OAI21_X1  g426(.A(new_n595), .B1(new_n609), .B2(new_n612), .ZN(new_n613));
  INV_X1    g427(.A(KEYINPUT93), .ZN(new_n614));
  NOR2_X1   g428(.A1(new_n317), .A2(G478), .ZN(new_n615));
  INV_X1    g429(.A(new_n615), .ZN(new_n616));
  NAND3_X1  g430(.A1(new_n613), .A2(new_n614), .A3(new_n616), .ZN(new_n617));
  INV_X1    g431(.A(new_n595), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n605), .A2(new_n608), .ZN(new_n619));
  NAND3_X1  g433(.A1(new_n611), .A2(new_n610), .A3(KEYINPUT92), .ZN(new_n620));
  AOI21_X1  g434(.A(new_n618), .B1(new_n619), .B2(new_n620), .ZN(new_n621));
  OAI21_X1  g435(.A(KEYINPUT93), .B1(new_n621), .B2(new_n615), .ZN(new_n622));
  AOI22_X1  g436(.A1(new_n272), .A2(new_n280), .B1(new_n617), .B2(new_n622), .ZN(new_n623));
  NAND3_X1  g437(.A1(new_n594), .A2(new_n331), .A3(new_n623), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n538), .A2(new_n540), .ZN(new_n625));
  NAND2_X1  g439(.A1(new_n625), .A2(new_n277), .ZN(new_n626));
  AOI21_X1  g440(.A(new_n541), .B1(new_n626), .B2(G472), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n586), .A2(new_n627), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n412), .A2(new_n475), .ZN(new_n629));
  NOR2_X1   g443(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  INV_X1    g444(.A(new_n630), .ZN(new_n631));
  NOR2_X1   g445(.A1(new_n624), .A2(new_n631), .ZN(new_n632));
  XNOR2_X1  g446(.A(KEYINPUT34), .B(G104), .ZN(new_n633));
  XNOR2_X1  g447(.A(new_n632), .B(new_n633), .ZN(G6));
  NAND2_X1  g448(.A1(new_n321), .A2(new_n322), .ZN(new_n635));
  INV_X1    g449(.A(new_n635), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n270), .A2(new_n271), .ZN(new_n637));
  OAI21_X1  g451(.A(new_n188), .B1(new_n248), .B2(new_n264), .ZN(new_n638));
  INV_X1    g452(.A(new_n271), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  AOI21_X1  g454(.A(new_n636), .B1(new_n637), .B2(new_n640), .ZN(new_n641));
  INV_X1    g455(.A(G475), .ZN(new_n642));
  AOI21_X1  g456(.A(G902), .B1(new_n273), .B2(new_n275), .ZN(new_n643));
  AOI21_X1  g457(.A(new_n642), .B1(new_n643), .B2(new_n278), .ZN(new_n644));
  XOR2_X1   g458(.A(new_n330), .B(KEYINPUT94), .Z(new_n645));
  INV_X1    g459(.A(new_n645), .ZN(new_n646));
  NOR2_X1   g460(.A1(new_n644), .A2(new_n646), .ZN(new_n647));
  NAND3_X1  g461(.A1(new_n594), .A2(new_n641), .A3(new_n647), .ZN(new_n648));
  NOR2_X1   g462(.A1(new_n648), .A2(new_n631), .ZN(new_n649));
  XNOR2_X1  g463(.A(KEYINPUT35), .B(G107), .ZN(new_n650));
  XNOR2_X1  g464(.A(new_n649), .B(new_n650), .ZN(G9));
  INV_X1    g465(.A(new_n627), .ZN(new_n652));
  INV_X1    g466(.A(new_n578), .ZN(new_n653));
  AOI21_X1  g467(.A(new_n653), .B1(new_n583), .B2(new_n584), .ZN(new_n654));
  OR3_X1    g468(.A1(new_n571), .A2(KEYINPUT36), .A3(new_n575), .ZN(new_n655));
  OAI21_X1  g469(.A(new_n571), .B1(KEYINPUT36), .B2(new_n575), .ZN(new_n656));
  AND3_X1   g470(.A1(new_n655), .A2(new_n579), .A3(new_n656), .ZN(new_n657));
  NOR2_X1   g471(.A1(new_n654), .A2(new_n657), .ZN(new_n658));
  NOR2_X1   g472(.A1(new_n652), .A2(new_n658), .ZN(new_n659));
  NAND2_X1  g473(.A1(new_n477), .A2(new_n659), .ZN(new_n660));
  XOR2_X1   g474(.A(KEYINPUT37), .B(G110), .Z(new_n661));
  XNOR2_X1  g475(.A(new_n660), .B(new_n661), .ZN(G12));
  NOR3_X1   g476(.A1(new_n629), .A2(new_n591), .A3(new_n593), .ZN(new_n663));
  INV_X1    g477(.A(new_n328), .ZN(new_n664));
  OAI21_X1  g478(.A(new_n326), .B1(new_n664), .B2(G900), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n280), .A2(new_n665), .ZN(new_n666));
  AOI211_X1 g480(.A(new_n636), .B(new_n666), .C1(new_n640), .C2(new_n637), .ZN(new_n667));
  INV_X1    g481(.A(new_n658), .ZN(new_n668));
  NAND4_X1  g482(.A1(new_n663), .A2(new_n553), .A3(new_n667), .A4(new_n668), .ZN(new_n669));
  XNOR2_X1  g483(.A(new_n669), .B(G128), .ZN(G30));
  NAND2_X1  g484(.A1(new_n548), .A2(new_n551), .ZN(new_n671));
  AOI21_X1  g485(.A(new_n671), .B1(new_n543), .B2(new_n544), .ZN(new_n672));
  NOR2_X1   g486(.A1(new_n510), .A2(new_n484), .ZN(new_n673));
  NOR2_X1   g487(.A1(new_n673), .A2(new_n503), .ZN(new_n674));
  OAI21_X1  g488(.A(new_n277), .B1(new_n519), .B2(new_n498), .ZN(new_n675));
  OAI21_X1  g489(.A(G472), .B1(new_n674), .B2(new_n675), .ZN(new_n676));
  NAND3_X1  g490(.A1(new_n672), .A2(KEYINPUT95), .A3(new_n676), .ZN(new_n677));
  INV_X1    g491(.A(KEYINPUT95), .ZN(new_n678));
  AND3_X1   g492(.A1(new_n541), .A2(KEYINPUT71), .A3(KEYINPUT32), .ZN(new_n679));
  OAI211_X1 g493(.A(new_n548), .B(new_n551), .C1(new_n679), .C2(new_n542), .ZN(new_n680));
  INV_X1    g494(.A(new_n676), .ZN(new_n681));
  OAI21_X1  g495(.A(new_n678), .B1(new_n680), .B2(new_n681), .ZN(new_n682));
  NAND2_X1  g496(.A1(new_n677), .A2(new_n682), .ZN(new_n683));
  INV_X1    g497(.A(new_n683), .ZN(new_n684));
  XOR2_X1   g498(.A(new_n472), .B(KEYINPUT38), .Z(new_n685));
  OR2_X1    g499(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  INV_X1    g500(.A(new_n629), .ZN(new_n687));
  XNOR2_X1  g501(.A(new_n665), .B(KEYINPUT39), .ZN(new_n688));
  NAND2_X1  g502(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  XNOR2_X1  g503(.A(new_n689), .B(KEYINPUT40), .ZN(new_n690));
  AOI21_X1  g504(.A(new_n636), .B1(new_n272), .B2(new_n280), .ZN(new_n691));
  NAND3_X1  g505(.A1(new_n691), .A2(new_n473), .A3(new_n658), .ZN(new_n692));
  XNOR2_X1  g506(.A(new_n692), .B(KEYINPUT96), .ZN(new_n693));
  NOR3_X1   g507(.A1(new_n686), .A2(new_n690), .A3(new_n693), .ZN(new_n694));
  XNOR2_X1  g508(.A(KEYINPUT97), .B(G143), .ZN(new_n695));
  XNOR2_X1  g509(.A(new_n694), .B(new_n695), .ZN(G45));
  NAND2_X1  g510(.A1(new_n272), .A2(new_n280), .ZN(new_n697));
  NAND2_X1  g511(.A1(new_n617), .A2(new_n622), .ZN(new_n698));
  NAND3_X1  g512(.A1(new_n697), .A2(new_n698), .A3(new_n665), .ZN(new_n699));
  INV_X1    g513(.A(new_n699), .ZN(new_n700));
  NAND4_X1  g514(.A1(new_n700), .A2(new_n663), .A3(new_n553), .A4(new_n668), .ZN(new_n701));
  XNOR2_X1  g515(.A(new_n701), .B(G146), .ZN(G48));
  NAND2_X1  g516(.A1(new_n403), .A2(new_n277), .ZN(new_n703));
  NAND2_X1  g517(.A1(new_n703), .A2(G469), .ZN(new_n704));
  NAND3_X1  g518(.A1(new_n704), .A2(new_n475), .A3(new_n405), .ZN(new_n705));
  INV_X1    g519(.A(new_n705), .ZN(new_n706));
  AND3_X1   g520(.A1(new_n522), .A2(KEYINPUT70), .A3(G472), .ZN(new_n707));
  AOI21_X1  g521(.A(KEYINPUT70), .B1(new_n522), .B2(G472), .ZN(new_n708));
  NOR2_X1   g522(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  OAI211_X1 g523(.A(new_n586), .B(new_n706), .C1(new_n680), .C2(new_n709), .ZN(new_n710));
  NOR2_X1   g524(.A1(new_n710), .A2(new_n624), .ZN(new_n711));
  XOR2_X1   g525(.A(KEYINPUT41), .B(G113), .Z(new_n712));
  XNOR2_X1  g526(.A(new_n711), .B(new_n712), .ZN(G15));
  NOR2_X1   g527(.A1(new_n710), .A2(new_n648), .ZN(new_n714));
  XNOR2_X1  g528(.A(new_n714), .B(new_n281), .ZN(G18));
  AOI21_X1  g529(.A(new_n658), .B1(new_n672), .B2(new_n527), .ZN(new_n716));
  INV_X1    g530(.A(KEYINPUT98), .ZN(new_n717));
  AOI211_X1 g531(.A(new_n644), .B(new_n332), .C1(new_n640), .C2(new_n265), .ZN(new_n718));
  NOR3_X1   g532(.A1(new_n705), .A2(new_n591), .A3(new_n593), .ZN(new_n719));
  NAND4_X1  g533(.A1(new_n716), .A2(new_n717), .A3(new_n718), .A4(new_n719), .ZN(new_n720));
  OAI211_X1 g534(.A(new_n718), .B(new_n668), .C1(new_n709), .C2(new_n680), .ZN(new_n721));
  NAND2_X1  g535(.A1(new_n594), .A2(new_n706), .ZN(new_n722));
  OAI21_X1  g536(.A(KEYINPUT98), .B1(new_n721), .B2(new_n722), .ZN(new_n723));
  NAND2_X1  g537(.A1(new_n720), .A2(new_n723), .ZN(new_n724));
  XNOR2_X1  g538(.A(new_n724), .B(G119), .ZN(G21));
  NOR2_X1   g539(.A1(new_n705), .A2(new_n646), .ZN(new_n726));
  NAND2_X1  g540(.A1(new_n539), .A2(KEYINPUT99), .ZN(new_n727));
  INV_X1    g541(.A(KEYINPUT99), .ZN(new_n728));
  NAND3_X1  g542(.A1(new_n520), .A2(new_n728), .A3(new_n500), .ZN(new_n729));
  NAND3_X1  g543(.A1(new_n727), .A2(new_n729), .A3(new_n503), .ZN(new_n730));
  AOI21_X1  g544(.A(new_n529), .B1(new_n730), .B2(new_n538), .ZN(new_n731));
  INV_X1    g545(.A(G472), .ZN(new_n732));
  AOI21_X1  g546(.A(new_n732), .B1(new_n625), .B2(new_n277), .ZN(new_n733));
  NOR2_X1   g547(.A1(new_n731), .A2(new_n733), .ZN(new_n734));
  INV_X1    g548(.A(KEYINPUT100), .ZN(new_n735));
  AND3_X1   g549(.A1(new_n734), .A2(new_n586), .A3(new_n735), .ZN(new_n736));
  AOI21_X1  g550(.A(new_n735), .B1(new_n734), .B2(new_n586), .ZN(new_n737));
  OAI21_X1  g551(.A(new_n726), .B1(new_n736), .B2(new_n737), .ZN(new_n738));
  NAND2_X1  g552(.A1(new_n594), .A2(new_n691), .ZN(new_n739));
  NOR2_X1   g553(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  XOR2_X1   g554(.A(new_n740), .B(G122), .Z(G24));
  NAND2_X1  g555(.A1(new_n668), .A2(new_n734), .ZN(new_n742));
  INV_X1    g556(.A(new_n742), .ZN(new_n743));
  NAND3_X1  g557(.A1(new_n700), .A2(new_n743), .A3(new_n719), .ZN(new_n744));
  XNOR2_X1  g558(.A(new_n744), .B(G125), .ZN(G27));
  NAND3_X1  g559(.A1(new_n470), .A2(new_n471), .A3(new_n473), .ZN(new_n746));
  INV_X1    g560(.A(KEYINPUT102), .ZN(new_n747));
  NAND2_X1  g561(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  NAND2_X1  g562(.A1(G469), .A2(G902), .ZN(new_n749));
  NAND2_X1  g563(.A1(new_n409), .A2(new_n338), .ZN(new_n750));
  NAND3_X1  g564(.A1(new_n407), .A2(new_n389), .A3(new_n399), .ZN(new_n751));
  NAND2_X1  g565(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  OAI21_X1  g566(.A(KEYINPUT101), .B1(new_n752), .B2(new_n404), .ZN(new_n753));
  INV_X1    g567(.A(KEYINPUT101), .ZN(new_n754));
  NAND4_X1  g568(.A1(new_n750), .A2(new_n754), .A3(new_n751), .A4(G469), .ZN(new_n755));
  NAND4_X1  g569(.A1(new_n405), .A2(new_n749), .A3(new_n753), .A4(new_n755), .ZN(new_n756));
  NAND4_X1  g570(.A1(new_n470), .A2(KEYINPUT102), .A3(new_n471), .A4(new_n473), .ZN(new_n757));
  NAND4_X1  g571(.A1(new_n748), .A2(new_n756), .A3(new_n475), .A4(new_n757), .ZN(new_n758));
  NOR2_X1   g572(.A1(new_n699), .A2(new_n758), .ZN(new_n759));
  INV_X1    g573(.A(KEYINPUT104), .ZN(new_n760));
  NOR2_X1   g574(.A1(new_n541), .A2(KEYINPUT32), .ZN(new_n761));
  AND2_X1   g575(.A1(new_n532), .A2(new_n537), .ZN(new_n762));
  AOI21_X1  g576(.A(new_n498), .B1(new_n520), .B2(new_n500), .ZN(new_n763));
  OAI211_X1 g577(.A(KEYINPUT32), .B(new_n528), .C1(new_n762), .C2(new_n763), .ZN(new_n764));
  NAND2_X1  g578(.A1(new_n764), .A2(KEYINPUT103), .ZN(new_n765));
  INV_X1    g579(.A(KEYINPUT103), .ZN(new_n766));
  NAND3_X1  g580(.A1(new_n541), .A2(new_n766), .A3(KEYINPUT32), .ZN(new_n767));
  AOI21_X1  g581(.A(new_n761), .B1(new_n765), .B2(new_n767), .ZN(new_n768));
  NAND2_X1  g582(.A1(new_n527), .A2(new_n768), .ZN(new_n769));
  AOI21_X1  g583(.A(new_n760), .B1(new_n769), .B2(new_n586), .ZN(new_n770));
  NAND2_X1  g584(.A1(new_n585), .A2(new_n578), .ZN(new_n771));
  INV_X1    g585(.A(new_n580), .ZN(new_n772));
  NAND2_X1  g586(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  AOI211_X1 g587(.A(KEYINPUT104), .B(new_n773), .C1(new_n527), .C2(new_n768), .ZN(new_n774));
  OAI21_X1  g588(.A(new_n759), .B1(new_n770), .B2(new_n774), .ZN(new_n775));
  NAND2_X1  g589(.A1(new_n775), .A2(KEYINPUT42), .ZN(new_n776));
  NAND2_X1  g590(.A1(new_n553), .A2(new_n586), .ZN(new_n777));
  INV_X1    g591(.A(new_n777), .ZN(new_n778));
  NOR2_X1   g592(.A1(new_n699), .A2(KEYINPUT42), .ZN(new_n779));
  INV_X1    g593(.A(new_n758), .ZN(new_n780));
  NAND3_X1  g594(.A1(new_n778), .A2(new_n779), .A3(new_n780), .ZN(new_n781));
  NAND2_X1  g595(.A1(new_n776), .A2(new_n781), .ZN(new_n782));
  XNOR2_X1  g596(.A(new_n782), .B(new_n207), .ZN(G33));
  NAND4_X1  g597(.A1(new_n780), .A2(new_n553), .A3(new_n667), .A4(new_n586), .ZN(new_n784));
  XNOR2_X1  g598(.A(new_n784), .B(G134), .ZN(G36));
  AOI21_X1  g599(.A(new_n644), .B1(new_n640), .B2(new_n265), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n786), .A2(new_n698), .ZN(new_n787));
  INV_X1    g601(.A(KEYINPUT106), .ZN(new_n788));
  NAND2_X1  g602(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  XNOR2_X1  g603(.A(new_n789), .B(KEYINPUT43), .ZN(new_n790));
  XNOR2_X1  g604(.A(new_n790), .B(KEYINPUT107), .ZN(new_n791));
  NAND3_X1  g605(.A1(new_n791), .A2(new_n652), .A3(new_n668), .ZN(new_n792));
  INV_X1    g606(.A(KEYINPUT44), .ZN(new_n793));
  NAND2_X1  g607(.A1(new_n792), .A2(new_n793), .ZN(new_n794));
  AND2_X1   g608(.A1(new_n748), .A2(new_n757), .ZN(new_n795));
  NAND4_X1  g609(.A1(new_n791), .A2(KEYINPUT44), .A3(new_n652), .A4(new_n668), .ZN(new_n796));
  OR2_X1    g610(.A1(new_n410), .A2(KEYINPUT45), .ZN(new_n797));
  NAND2_X1  g611(.A1(new_n410), .A2(KEYINPUT45), .ZN(new_n798));
  NAND3_X1  g612(.A1(new_n797), .A2(G469), .A3(new_n798), .ZN(new_n799));
  NAND2_X1  g613(.A1(new_n799), .A2(new_n749), .ZN(new_n800));
  INV_X1    g614(.A(KEYINPUT46), .ZN(new_n801));
  OAI21_X1  g615(.A(new_n405), .B1(new_n800), .B2(new_n801), .ZN(new_n802));
  AOI22_X1  g616(.A1(new_n802), .A2(KEYINPUT105), .B1(new_n801), .B2(new_n800), .ZN(new_n803));
  OAI21_X1  g617(.A(new_n803), .B1(KEYINPUT105), .B2(new_n802), .ZN(new_n804));
  AND3_X1   g618(.A1(new_n804), .A2(new_n475), .A3(new_n688), .ZN(new_n805));
  NAND4_X1  g619(.A1(new_n794), .A2(new_n795), .A3(new_n796), .A4(new_n805), .ZN(new_n806));
  XNOR2_X1  g620(.A(new_n806), .B(G137), .ZN(G39));
  NAND2_X1  g621(.A1(new_n804), .A2(new_n475), .ZN(new_n808));
  NAND2_X1  g622(.A1(new_n808), .A2(KEYINPUT108), .ZN(new_n809));
  INV_X1    g623(.A(KEYINPUT108), .ZN(new_n810));
  NAND3_X1  g624(.A1(new_n804), .A2(new_n810), .A3(new_n475), .ZN(new_n811));
  XNOR2_X1  g625(.A(KEYINPUT109), .B(KEYINPUT47), .ZN(new_n812));
  AND3_X1   g626(.A1(new_n809), .A2(new_n811), .A3(new_n812), .ZN(new_n813));
  AOI22_X1  g627(.A1(new_n809), .A2(new_n811), .B1(KEYINPUT109), .B2(KEYINPUT47), .ZN(new_n814));
  NOR2_X1   g628(.A1(new_n813), .A2(new_n814), .ZN(new_n815));
  INV_X1    g629(.A(new_n795), .ZN(new_n816));
  NOR3_X1   g630(.A1(new_n816), .A2(new_n553), .A3(new_n586), .ZN(new_n817));
  NAND3_X1  g631(.A1(new_n815), .A2(new_n700), .A3(new_n817), .ZN(new_n818));
  XNOR2_X1  g632(.A(new_n818), .B(G140), .ZN(G42));
  INV_X1    g633(.A(KEYINPUT51), .ZN(new_n820));
  OR2_X1    g634(.A1(new_n736), .A2(new_n737), .ZN(new_n821));
  INV_X1    g635(.A(new_n821), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n790), .A2(new_n327), .ZN(new_n823));
  INV_X1    g637(.A(KEYINPUT114), .ZN(new_n824));
  NAND2_X1  g638(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  NAND3_X1  g639(.A1(new_n790), .A2(KEYINPUT114), .A3(new_n327), .ZN(new_n826));
  AOI21_X1  g640(.A(new_n822), .B1(new_n825), .B2(new_n826), .ZN(new_n827));
  NAND2_X1  g641(.A1(new_n827), .A2(new_n795), .ZN(new_n828));
  INV_X1    g642(.A(KEYINPUT115), .ZN(new_n829));
  NAND2_X1  g643(.A1(new_n828), .A2(new_n829), .ZN(new_n830));
  NAND3_X1  g644(.A1(new_n827), .A2(KEYINPUT115), .A3(new_n795), .ZN(new_n831));
  AND2_X1   g645(.A1(new_n704), .A2(new_n405), .ZN(new_n832));
  INV_X1    g646(.A(new_n475), .ZN(new_n833));
  NAND2_X1  g647(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  OAI21_X1  g648(.A(new_n834), .B1(new_n813), .B2(new_n814), .ZN(new_n835));
  AND3_X1   g649(.A1(new_n830), .A2(new_n831), .A3(new_n835), .ZN(new_n836));
  NOR2_X1   g650(.A1(new_n816), .A2(new_n705), .ZN(new_n837));
  NAND4_X1  g651(.A1(new_n684), .A2(new_n586), .A3(new_n327), .A4(new_n837), .ZN(new_n838));
  NOR3_X1   g652(.A1(new_n838), .A2(new_n697), .A3(new_n698), .ZN(new_n839));
  INV_X1    g653(.A(new_n837), .ZN(new_n840));
  AOI21_X1  g654(.A(new_n840), .B1(new_n825), .B2(new_n826), .ZN(new_n841));
  AOI21_X1  g655(.A(new_n839), .B1(new_n841), .B2(new_n743), .ZN(new_n842));
  AND3_X1   g656(.A1(new_n685), .A2(new_n592), .A3(new_n706), .ZN(new_n843));
  AND3_X1   g657(.A1(new_n827), .A2(KEYINPUT50), .A3(new_n843), .ZN(new_n844));
  AOI21_X1  g658(.A(KEYINPUT50), .B1(new_n827), .B2(new_n843), .ZN(new_n845));
  OAI21_X1  g659(.A(new_n842), .B1(new_n844), .B2(new_n845), .ZN(new_n846));
  OAI21_X1  g660(.A(new_n820), .B1(new_n836), .B2(new_n846), .ZN(new_n847));
  OR2_X1    g661(.A1(new_n844), .A2(new_n845), .ZN(new_n848));
  NAND3_X1  g662(.A1(new_n830), .A2(new_n835), .A3(new_n831), .ZN(new_n849));
  NAND4_X1  g663(.A1(new_n848), .A2(new_n849), .A3(KEYINPUT51), .A4(new_n842), .ZN(new_n850));
  NAND2_X1  g664(.A1(new_n827), .A2(new_n719), .ZN(new_n851));
  INV_X1    g665(.A(new_n623), .ZN(new_n852));
  OAI211_X1 g666(.A(new_n851), .B(new_n324), .C1(new_n852), .C2(new_n838), .ZN(new_n853));
  NOR2_X1   g667(.A1(new_n764), .A2(KEYINPUT103), .ZN(new_n854));
  AOI21_X1  g668(.A(new_n766), .B1(new_n541), .B2(KEYINPUT32), .ZN(new_n855));
  OAI22_X1  g669(.A1(new_n854), .A2(new_n855), .B1(KEYINPUT32), .B2(new_n541), .ZN(new_n856));
  OAI21_X1  g670(.A(new_n586), .B1(new_n856), .B2(new_n709), .ZN(new_n857));
  NAND2_X1  g671(.A1(new_n857), .A2(KEYINPUT104), .ZN(new_n858));
  NAND3_X1  g672(.A1(new_n769), .A2(new_n760), .A3(new_n586), .ZN(new_n859));
  NAND2_X1  g673(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  NAND2_X1  g674(.A1(new_n841), .A2(new_n860), .ZN(new_n861));
  OR2_X1    g675(.A1(new_n861), .A2(KEYINPUT48), .ZN(new_n862));
  NAND2_X1  g676(.A1(new_n861), .A2(KEYINPUT48), .ZN(new_n863));
  AOI21_X1  g677(.A(new_n853), .B1(new_n862), .B2(new_n863), .ZN(new_n864));
  NAND3_X1  g678(.A1(new_n847), .A2(new_n850), .A3(new_n864), .ZN(new_n865));
  AOI21_X1  g679(.A(new_n710), .B1(new_n624), .B2(new_n648), .ZN(new_n866));
  NOR2_X1   g680(.A1(new_n866), .A2(new_n740), .ZN(new_n867));
  AOI21_X1  g681(.A(new_n754), .B1(new_n410), .B2(G469), .ZN(new_n868));
  NAND2_X1  g682(.A1(new_n755), .A2(new_n749), .ZN(new_n869));
  NOR2_X1   g683(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  AOI21_X1  g684(.A(new_n833), .B1(new_n870), .B2(new_n405), .ZN(new_n871));
  NAND4_X1  g685(.A1(new_n795), .A2(new_n623), .A3(new_n665), .A4(new_n871), .ZN(new_n872));
  OAI21_X1  g686(.A(KEYINPUT111), .B1(new_n872), .B2(new_n742), .ZN(new_n873));
  INV_X1    g687(.A(KEYINPUT111), .ZN(new_n874));
  NAND3_X1  g688(.A1(new_n759), .A2(new_n874), .A3(new_n743), .ZN(new_n875));
  NAND2_X1  g689(.A1(new_n873), .A2(new_n875), .ZN(new_n876));
  AND2_X1   g690(.A1(new_n637), .A2(new_n640), .ZN(new_n877));
  INV_X1    g691(.A(KEYINPUT110), .ZN(new_n878));
  NAND2_X1  g692(.A1(new_n635), .A2(new_n878), .ZN(new_n879));
  NAND3_X1  g693(.A1(new_n321), .A2(KEYINPUT110), .A3(new_n322), .ZN(new_n880));
  NAND4_X1  g694(.A1(new_n879), .A2(new_n280), .A3(new_n880), .A4(new_n665), .ZN(new_n881));
  NOR3_X1   g695(.A1(new_n877), .A2(new_n658), .A3(new_n881), .ZN(new_n882));
  NAND4_X1  g696(.A1(new_n882), .A2(new_n553), .A3(new_n687), .A4(new_n795), .ZN(new_n883));
  AND2_X1   g697(.A1(new_n883), .A2(new_n784), .ZN(new_n884));
  AND4_X1   g698(.A1(new_n724), .A2(new_n867), .A3(new_n876), .A4(new_n884), .ZN(new_n885));
  INV_X1    g699(.A(KEYINPUT52), .ZN(new_n886));
  NAND3_X1  g700(.A1(new_n701), .A2(new_n669), .A3(new_n744), .ZN(new_n887));
  AND2_X1   g701(.A1(new_n658), .A2(new_n665), .ZN(new_n888));
  NAND4_X1  g702(.A1(new_n594), .A2(new_n888), .A3(new_n691), .A4(new_n871), .ZN(new_n889));
  AOI21_X1  g703(.A(new_n889), .B1(new_n682), .B2(new_n677), .ZN(new_n890));
  OAI21_X1  g704(.A(new_n886), .B1(new_n887), .B2(new_n890), .ZN(new_n891));
  INV_X1    g705(.A(new_n889), .ZN(new_n892));
  NAND2_X1  g706(.A1(new_n683), .A2(new_n892), .ZN(new_n893));
  OAI211_X1 g707(.A(new_n716), .B(new_n663), .C1(new_n667), .C2(new_n700), .ZN(new_n894));
  NAND4_X1  g708(.A1(new_n893), .A2(new_n894), .A3(KEYINPUT52), .A4(new_n744), .ZN(new_n895));
  NAND2_X1  g709(.A1(new_n891), .A2(new_n895), .ZN(new_n896));
  NAND3_X1  g710(.A1(new_n472), .A2(new_n474), .A3(new_n645), .ZN(new_n897));
  NOR3_X1   g711(.A1(new_n628), .A2(new_n629), .A3(new_n897), .ZN(new_n898));
  NAND2_X1  g712(.A1(new_n879), .A2(new_n880), .ZN(new_n899));
  NAND3_X1  g713(.A1(new_n272), .A2(new_n280), .A3(new_n899), .ZN(new_n900));
  AND2_X1   g714(.A1(new_n617), .A2(new_n622), .ZN(new_n901));
  OAI21_X1  g715(.A(new_n900), .B1(new_n786), .B2(new_n901), .ZN(new_n902));
  NAND2_X1  g716(.A1(new_n898), .A2(new_n902), .ZN(new_n903));
  AND4_X1   g717(.A1(KEYINPUT53), .A2(new_n587), .A3(new_n903), .A4(new_n660), .ZN(new_n904));
  AND3_X1   g718(.A1(new_n776), .A2(new_n904), .A3(new_n781), .ZN(new_n905));
  NAND3_X1  g719(.A1(new_n885), .A2(new_n896), .A3(new_n905), .ZN(new_n906));
  NAND2_X1  g720(.A1(new_n906), .A2(KEYINPUT112), .ZN(new_n907));
  NAND4_X1  g721(.A1(new_n867), .A2(new_n724), .A3(new_n876), .A4(new_n884), .ZN(new_n908));
  NAND3_X1  g722(.A1(new_n776), .A2(new_n904), .A3(new_n781), .ZN(new_n909));
  NOR2_X1   g723(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  INV_X1    g724(.A(KEYINPUT112), .ZN(new_n911));
  NAND3_X1  g725(.A1(new_n910), .A2(new_n911), .A3(new_n896), .ZN(new_n912));
  NAND2_X1  g726(.A1(new_n907), .A2(new_n912), .ZN(new_n913));
  INV_X1    g727(.A(KEYINPUT54), .ZN(new_n914));
  INV_X1    g728(.A(new_n782), .ZN(new_n915));
  AND3_X1   g729(.A1(new_n587), .A2(new_n903), .A3(new_n660), .ZN(new_n916));
  AND3_X1   g730(.A1(new_n867), .A2(new_n724), .A3(new_n916), .ZN(new_n917));
  AND2_X1   g731(.A1(new_n876), .A2(new_n884), .ZN(new_n918));
  NAND4_X1  g732(.A1(new_n896), .A2(new_n915), .A3(new_n917), .A4(new_n918), .ZN(new_n919));
  INV_X1    g733(.A(KEYINPUT53), .ZN(new_n920));
  NAND2_X1  g734(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  NAND3_X1  g735(.A1(new_n913), .A2(new_n914), .A3(new_n921), .ZN(new_n922));
  INV_X1    g736(.A(KEYINPUT113), .ZN(new_n923));
  NAND2_X1  g737(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  NAND4_X1  g738(.A1(new_n913), .A2(KEYINPUT113), .A3(new_n914), .A4(new_n921), .ZN(new_n925));
  NAND2_X1  g739(.A1(new_n921), .A2(new_n906), .ZN(new_n926));
  NAND2_X1  g740(.A1(new_n926), .A2(KEYINPUT54), .ZN(new_n927));
  NAND3_X1  g741(.A1(new_n924), .A2(new_n925), .A3(new_n927), .ZN(new_n928));
  OAI22_X1  g742(.A1(new_n865), .A2(new_n928), .B1(G952), .B2(G953), .ZN(new_n929));
  XOR2_X1   g743(.A(new_n832), .B(KEYINPUT49), .Z(new_n930));
  NAND4_X1  g744(.A1(new_n685), .A2(new_n586), .A3(new_n474), .A4(new_n475), .ZN(new_n931));
  OR4_X1    g745(.A1(new_n683), .A2(new_n930), .A3(new_n931), .A4(new_n787), .ZN(new_n932));
  NAND2_X1  g746(.A1(new_n929), .A2(new_n932), .ZN(G75));
  INV_X1    g747(.A(new_n203), .ZN(new_n934));
  NAND2_X1  g748(.A1(new_n934), .A2(new_n323), .ZN(new_n935));
  XOR2_X1   g749(.A(new_n935), .B(KEYINPUT118), .Z(new_n936));
  XOR2_X1   g750(.A(new_n936), .B(KEYINPUT119), .Z(new_n937));
  AOI21_X1  g751(.A(new_n277), .B1(new_n913), .B2(new_n921), .ZN(new_n938));
  AOI21_X1  g752(.A(KEYINPUT56), .B1(new_n938), .B2(G210), .ZN(new_n939));
  NAND2_X1  g753(.A1(new_n460), .A2(new_n461), .ZN(new_n940));
  XNOR2_X1  g754(.A(new_n940), .B(KEYINPUT116), .ZN(new_n941));
  XOR2_X1   g755(.A(new_n941), .B(KEYINPUT55), .Z(new_n942));
  XNOR2_X1  g756(.A(new_n942), .B(new_n463), .ZN(new_n943));
  OAI21_X1  g757(.A(new_n937), .B1(new_n939), .B2(new_n943), .ZN(new_n944));
  NAND2_X1  g758(.A1(new_n939), .A2(new_n943), .ZN(new_n945));
  INV_X1    g759(.A(KEYINPUT117), .ZN(new_n946));
  NAND2_X1  g760(.A1(new_n945), .A2(new_n946), .ZN(new_n947));
  NAND3_X1  g761(.A1(new_n939), .A2(KEYINPUT117), .A3(new_n943), .ZN(new_n948));
  AOI21_X1  g762(.A(new_n944), .B1(new_n947), .B2(new_n948), .ZN(G51));
  INV_X1    g763(.A(new_n936), .ZN(new_n950));
  AND4_X1   g764(.A1(new_n911), .A2(new_n885), .A3(new_n896), .A4(new_n905), .ZN(new_n951));
  AOI21_X1  g765(.A(new_n911), .B1(new_n910), .B2(new_n896), .ZN(new_n952));
  OAI21_X1  g766(.A(new_n921), .B1(new_n951), .B2(new_n952), .ZN(new_n953));
  NAND2_X1  g767(.A1(new_n953), .A2(KEYINPUT54), .ZN(new_n954));
  INV_X1    g768(.A(KEYINPUT120), .ZN(new_n955));
  NAND3_X1  g769(.A1(new_n954), .A2(new_n955), .A3(new_n922), .ZN(new_n956));
  NAND3_X1  g770(.A1(new_n953), .A2(KEYINPUT120), .A3(KEYINPUT54), .ZN(new_n957));
  XOR2_X1   g771(.A(new_n749), .B(KEYINPUT57), .Z(new_n958));
  NAND3_X1  g772(.A1(new_n956), .A2(new_n957), .A3(new_n958), .ZN(new_n959));
  NAND2_X1  g773(.A1(new_n959), .A2(new_n403), .ZN(new_n960));
  INV_X1    g774(.A(new_n799), .ZN(new_n961));
  AND3_X1   g775(.A1(new_n938), .A2(KEYINPUT121), .A3(new_n961), .ZN(new_n962));
  AOI21_X1  g776(.A(KEYINPUT121), .B1(new_n938), .B2(new_n961), .ZN(new_n963));
  NOR2_X1   g777(.A1(new_n962), .A2(new_n963), .ZN(new_n964));
  AOI21_X1  g778(.A(new_n950), .B1(new_n960), .B2(new_n964), .ZN(G54));
  AND3_X1   g779(.A1(new_n938), .A2(KEYINPUT58), .A3(G475), .ZN(new_n966));
  NAND2_X1  g780(.A1(new_n269), .A2(new_n263), .ZN(new_n967));
  INV_X1    g781(.A(new_n967), .ZN(new_n968));
  OR2_X1    g782(.A1(new_n966), .A2(new_n968), .ZN(new_n969));
  NAND2_X1  g783(.A1(new_n966), .A2(new_n968), .ZN(new_n970));
  AOI21_X1  g784(.A(new_n950), .B1(new_n969), .B2(new_n970), .ZN(G60));
  NAND2_X1  g785(.A1(new_n619), .A2(new_n620), .ZN(new_n972));
  NAND2_X1  g786(.A1(G478), .A2(G902), .ZN(new_n973));
  XNOR2_X1  g787(.A(new_n973), .B(KEYINPUT59), .ZN(new_n974));
  NAND4_X1  g788(.A1(new_n956), .A2(new_n972), .A3(new_n957), .A4(new_n974), .ZN(new_n975));
  NAND2_X1  g789(.A1(new_n975), .A2(new_n937), .ZN(new_n976));
  AOI21_X1  g790(.A(new_n972), .B1(new_n928), .B2(new_n974), .ZN(new_n977));
  NOR2_X1   g791(.A1(new_n976), .A2(new_n977), .ZN(G63));
  INV_X1    g792(.A(KEYINPUT123), .ZN(new_n979));
  AND2_X1   g793(.A1(new_n576), .A2(new_n577), .ZN(new_n980));
  NAND2_X1  g794(.A1(G217), .A2(G902), .ZN(new_n981));
  XNOR2_X1  g795(.A(new_n981), .B(KEYINPUT60), .ZN(new_n982));
  INV_X1    g796(.A(new_n982), .ZN(new_n983));
  AOI21_X1  g797(.A(new_n980), .B1(new_n953), .B2(new_n983), .ZN(new_n984));
  INV_X1    g798(.A(new_n937), .ZN(new_n985));
  OAI21_X1  g799(.A(new_n979), .B1(new_n984), .B2(new_n985), .ZN(new_n986));
  OR2_X1    g800(.A1(KEYINPUT123), .A2(KEYINPUT61), .ZN(new_n987));
  AOI21_X1  g801(.A(new_n982), .B1(new_n913), .B2(new_n921), .ZN(new_n988));
  OAI211_X1 g802(.A(new_n937), .B(new_n987), .C1(new_n988), .C2(new_n980), .ZN(new_n989));
  INV_X1    g803(.A(KEYINPUT122), .ZN(new_n990));
  AND2_X1   g804(.A1(new_n655), .A2(new_n656), .ZN(new_n991));
  NAND3_X1  g805(.A1(new_n988), .A2(new_n990), .A3(new_n991), .ZN(new_n992));
  NAND3_X1  g806(.A1(new_n953), .A2(new_n991), .A3(new_n983), .ZN(new_n993));
  NAND2_X1  g807(.A1(new_n993), .A2(KEYINPUT122), .ZN(new_n994));
  NAND4_X1  g808(.A1(new_n986), .A2(new_n989), .A3(new_n992), .A4(new_n994), .ZN(new_n995));
  INV_X1    g809(.A(new_n993), .ZN(new_n996));
  OAI21_X1  g810(.A(KEYINPUT61), .B1(new_n989), .B2(new_n996), .ZN(new_n997));
  AND2_X1   g811(.A1(new_n995), .A2(new_n997), .ZN(G66));
  INV_X1    g812(.A(new_n329), .ZN(new_n999));
  AOI21_X1  g813(.A(new_n194), .B1(new_n999), .B2(G224), .ZN(new_n1000));
  XOR2_X1   g814(.A(new_n917), .B(KEYINPUT124), .Z(new_n1001));
  INV_X1    g815(.A(new_n1001), .ZN(new_n1002));
  AOI21_X1  g816(.A(new_n1000), .B1(new_n1002), .B2(new_n203), .ZN(new_n1003));
  INV_X1    g817(.A(G898), .ZN(new_n1004));
  AOI21_X1  g818(.A(new_n941), .B1(new_n1004), .B2(new_n934), .ZN(new_n1005));
  XNOR2_X1  g819(.A(new_n1003), .B(new_n1005), .ZN(G69));
  AOI21_X1  g820(.A(new_n203), .B1(G227), .B2(G900), .ZN(new_n1007));
  INV_X1    g821(.A(new_n1007), .ZN(new_n1008));
  NAND3_X1  g822(.A1(new_n894), .A2(new_n744), .A3(new_n784), .ZN(new_n1009));
  AOI21_X1  g823(.A(new_n739), .B1(new_n858), .B2(new_n859), .ZN(new_n1010));
  AOI211_X1 g824(.A(new_n1009), .B(new_n782), .C1(new_n805), .C2(new_n1010), .ZN(new_n1011));
  NAND4_X1  g825(.A1(new_n806), .A2(new_n818), .A3(new_n203), .A4(new_n1011), .ZN(new_n1012));
  NOR2_X1   g826(.A1(new_n533), .A2(new_n534), .ZN(new_n1013));
  NAND2_X1  g827(.A1(new_n217), .A2(new_n221), .ZN(new_n1014));
  XNOR2_X1  g828(.A(new_n1014), .B(KEYINPUT125), .ZN(new_n1015));
  XNOR2_X1  g829(.A(new_n1013), .B(new_n1015), .ZN(new_n1016));
  AOI21_X1  g830(.A(new_n1016), .B1(G900), .B2(new_n934), .ZN(new_n1017));
  NAND2_X1  g831(.A1(new_n1012), .A2(new_n1017), .ZN(new_n1018));
  NOR2_X1   g832(.A1(new_n694), .A2(new_n887), .ZN(new_n1019));
  XNOR2_X1  g833(.A(new_n1019), .B(KEYINPUT62), .ZN(new_n1020));
  AOI21_X1  g834(.A(new_n689), .B1(new_n852), .B2(new_n900), .ZN(new_n1021));
  NAND3_X1  g835(.A1(new_n778), .A2(new_n1021), .A3(new_n795), .ZN(new_n1022));
  NAND4_X1  g836(.A1(new_n1020), .A2(new_n806), .A3(new_n818), .A4(new_n1022), .ZN(new_n1023));
  AND2_X1   g837(.A1(new_n1023), .A2(new_n203), .ZN(new_n1024));
  XOR2_X1   g838(.A(new_n1016), .B(KEYINPUT126), .Z(new_n1025));
  INV_X1    g839(.A(new_n1025), .ZN(new_n1026));
  OAI211_X1 g840(.A(new_n1008), .B(new_n1018), .C1(new_n1024), .C2(new_n1026), .ZN(new_n1027));
  AOI21_X1  g841(.A(new_n1026), .B1(new_n1023), .B2(new_n203), .ZN(new_n1028));
  INV_X1    g842(.A(new_n1018), .ZN(new_n1029));
  OAI21_X1  g843(.A(new_n1007), .B1(new_n1028), .B2(new_n1029), .ZN(new_n1030));
  NAND2_X1  g844(.A1(new_n1027), .A2(new_n1030), .ZN(G72));
  XNOR2_X1  g845(.A(KEYINPUT127), .B(KEYINPUT63), .ZN(new_n1032));
  NAND2_X1  g846(.A1(G472), .A2(G902), .ZN(new_n1033));
  XNOR2_X1  g847(.A(new_n1032), .B(new_n1033), .ZN(new_n1034));
  OAI21_X1  g848(.A(new_n511), .B1(new_n510), .B2(new_n531), .ZN(new_n1035));
  NAND3_X1  g849(.A1(new_n926), .A2(new_n1034), .A3(new_n1035), .ZN(new_n1036));
  NAND2_X1  g850(.A1(new_n1036), .A2(new_n936), .ZN(new_n1037));
  NAND2_X1  g851(.A1(new_n673), .A2(new_n503), .ZN(new_n1038));
  NAND4_X1  g852(.A1(new_n806), .A2(new_n818), .A3(new_n1001), .A4(new_n1011), .ZN(new_n1039));
  AOI21_X1  g853(.A(new_n1038), .B1(new_n1039), .B2(new_n1034), .ZN(new_n1040));
  OAI21_X1  g854(.A(new_n1034), .B1(new_n1023), .B2(new_n1002), .ZN(new_n1041));
  AOI211_X1 g855(.A(new_n1037), .B(new_n1040), .C1(new_n1041), .C2(new_n674), .ZN(G57));
endmodule


