//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 0 1 0 1 1 0 1 0 0 0 1 1 0 1 0 1 0 1 1 0 1 1 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 1 1 1 0 0 1 0 0 1 0 1 1 0 0 1 1 1 0 1 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:18:23 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n690, new_n691, new_n692,
    new_n693, new_n695, new_n696, new_n697, new_n698, new_n699, new_n700,
    new_n701, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n716, new_n717, new_n718, new_n719, new_n720, new_n721, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n752,
    new_n753, new_n754, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n770, new_n771, new_n772, new_n773, new_n774, new_n775,
    new_n776, new_n777, new_n778, new_n779, new_n780, new_n781, new_n782,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n791,
    new_n792, new_n793, new_n794, new_n796, new_n797, new_n798, new_n799,
    new_n800, new_n802, new_n804, new_n805, new_n806, new_n807, new_n808,
    new_n809, new_n810, new_n811, new_n812, new_n813, new_n814, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n822, new_n823, new_n824,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n870, new_n871, new_n873, new_n874, new_n876, new_n877, new_n878,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n952, new_n953, new_n954, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n965, new_n966,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n981, new_n982,
    new_n984, new_n985, new_n986, new_n987, new_n988, new_n989, new_n991,
    new_n992, new_n993, new_n994, new_n995, new_n997, new_n998, new_n999,
    new_n1000, new_n1001, new_n1002, new_n1003, new_n1004, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1018, new_n1019;
  NAND2_X1  g000(.A1(G229gat), .A2(G233gat), .ZN(new_n202));
  XOR2_X1   g001(.A(new_n202), .B(KEYINPUT13), .Z(new_n203));
  INV_X1    g002(.A(new_n203), .ZN(new_n204));
  INV_X1    g003(.A(G1gat), .ZN(new_n205));
  NAND2_X1  g004(.A1(new_n205), .A2(KEYINPUT16), .ZN(new_n206));
  INV_X1    g005(.A(G15gat), .ZN(new_n207));
  NAND2_X1  g006(.A1(new_n207), .A2(G22gat), .ZN(new_n208));
  INV_X1    g007(.A(G22gat), .ZN(new_n209));
  NAND2_X1  g008(.A1(new_n209), .A2(G15gat), .ZN(new_n210));
  NAND3_X1  g009(.A1(new_n206), .A2(new_n208), .A3(new_n210), .ZN(new_n211));
  INV_X1    g010(.A(new_n211), .ZN(new_n212));
  AOI21_X1  g011(.A(G1gat), .B1(new_n208), .B2(new_n210), .ZN(new_n213));
  NOR3_X1   g012(.A1(new_n212), .A2(new_n213), .A3(G8gat), .ZN(new_n214));
  INV_X1    g013(.A(G8gat), .ZN(new_n215));
  INV_X1    g014(.A(new_n213), .ZN(new_n216));
  AOI21_X1  g015(.A(new_n215), .B1(new_n216), .B2(new_n211), .ZN(new_n217));
  OR2_X1    g016(.A1(new_n214), .A2(new_n217), .ZN(new_n218));
  INV_X1    g017(.A(G50gat), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n219), .A2(G43gat), .ZN(new_n220));
  INV_X1    g019(.A(G43gat), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n221), .A2(G50gat), .ZN(new_n222));
  NAND3_X1  g021(.A1(new_n220), .A2(new_n222), .A3(KEYINPUT15), .ZN(new_n223));
  INV_X1    g022(.A(new_n223), .ZN(new_n224));
  INV_X1    g023(.A(G29gat), .ZN(new_n225));
  INV_X1    g024(.A(G36gat), .ZN(new_n226));
  NAND3_X1  g025(.A1(new_n225), .A2(new_n226), .A3(KEYINPUT91), .ZN(new_n227));
  INV_X1    g026(.A(KEYINPUT91), .ZN(new_n228));
  OAI21_X1  g027(.A(new_n228), .B1(G29gat), .B2(G36gat), .ZN(new_n229));
  AND3_X1   g028(.A1(new_n227), .A2(new_n229), .A3(KEYINPUT14), .ZN(new_n230));
  OAI22_X1  g029(.A1(new_n229), .A2(KEYINPUT14), .B1(new_n225), .B2(new_n226), .ZN(new_n231));
  OAI21_X1  g030(.A(new_n224), .B1(new_n230), .B2(new_n231), .ZN(new_n232));
  AND2_X1   g031(.A1(G29gat), .A2(G36gat), .ZN(new_n233));
  AOI21_X1  g032(.A(KEYINPUT91), .B1(new_n225), .B2(new_n226), .ZN(new_n234));
  INV_X1    g033(.A(KEYINPUT14), .ZN(new_n235));
  AOI21_X1  g034(.A(new_n233), .B1(new_n234), .B2(new_n235), .ZN(new_n236));
  INV_X1    g035(.A(KEYINPUT15), .ZN(new_n237));
  NOR2_X1   g036(.A1(new_n221), .A2(G50gat), .ZN(new_n238));
  NOR2_X1   g037(.A1(new_n219), .A2(G43gat), .ZN(new_n239));
  OAI21_X1  g038(.A(new_n237), .B1(new_n238), .B2(new_n239), .ZN(new_n240));
  NAND3_X1  g039(.A1(new_n227), .A2(new_n229), .A3(KEYINPUT14), .ZN(new_n241));
  NAND4_X1  g040(.A1(new_n236), .A2(new_n240), .A3(new_n223), .A4(new_n241), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n232), .A2(new_n242), .ZN(new_n243));
  INV_X1    g042(.A(KEYINPUT92), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n243), .A2(new_n244), .ZN(new_n245));
  NAND3_X1  g044(.A1(new_n232), .A2(new_n242), .A3(KEYINPUT92), .ZN(new_n246));
  NAND3_X1  g045(.A1(new_n218), .A2(new_n245), .A3(new_n246), .ZN(new_n247));
  NOR2_X1   g046(.A1(new_n214), .A2(new_n217), .ZN(new_n248));
  AND3_X1   g047(.A1(new_n232), .A2(new_n242), .A3(KEYINPUT92), .ZN(new_n249));
  AOI21_X1  g048(.A(KEYINPUT92), .B1(new_n232), .B2(new_n242), .ZN(new_n250));
  OAI21_X1  g049(.A(new_n248), .B1(new_n249), .B2(new_n250), .ZN(new_n251));
  AOI21_X1  g050(.A(new_n204), .B1(new_n247), .B2(new_n251), .ZN(new_n252));
  XOR2_X1   g051(.A(KEYINPUT93), .B(KEYINPUT17), .Z(new_n253));
  NOR3_X1   g052(.A1(new_n249), .A2(new_n250), .A3(new_n253), .ZN(new_n254));
  NAND3_X1  g053(.A1(new_n232), .A2(new_n242), .A3(KEYINPUT17), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n248), .A2(new_n255), .ZN(new_n256));
  OAI211_X1 g055(.A(new_n202), .B(new_n247), .C1(new_n254), .C2(new_n256), .ZN(new_n257));
  AOI21_X1  g056(.A(KEYINPUT18), .B1(new_n257), .B2(KEYINPUT94), .ZN(new_n258));
  INV_X1    g057(.A(new_n256), .ZN(new_n259));
  INV_X1    g058(.A(new_n253), .ZN(new_n260));
  NAND3_X1  g059(.A1(new_n245), .A2(new_n246), .A3(new_n260), .ZN(new_n261));
  NOR2_X1   g060(.A1(new_n249), .A2(new_n250), .ZN(new_n262));
  AOI22_X1  g061(.A1(new_n259), .A2(new_n261), .B1(new_n262), .B2(new_n218), .ZN(new_n263));
  INV_X1    g062(.A(KEYINPUT94), .ZN(new_n264));
  NAND3_X1  g063(.A1(new_n263), .A2(new_n264), .A3(new_n202), .ZN(new_n265));
  AOI21_X1  g064(.A(new_n252), .B1(new_n258), .B2(new_n265), .ZN(new_n266));
  INV_X1    g065(.A(KEYINPUT95), .ZN(new_n267));
  INV_X1    g066(.A(KEYINPUT18), .ZN(new_n268));
  OAI21_X1  g067(.A(new_n267), .B1(new_n257), .B2(new_n268), .ZN(new_n269));
  NAND4_X1  g068(.A1(new_n263), .A2(KEYINPUT95), .A3(KEYINPUT18), .A4(new_n202), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n266), .A2(new_n271), .ZN(new_n272));
  XOR2_X1   g071(.A(G169gat), .B(G197gat), .Z(new_n273));
  XNOR2_X1  g072(.A(new_n273), .B(KEYINPUT90), .ZN(new_n274));
  XOR2_X1   g073(.A(G113gat), .B(G141gat), .Z(new_n275));
  XNOR2_X1  g074(.A(new_n274), .B(new_n275), .ZN(new_n276));
  XNOR2_X1  g075(.A(KEYINPUT89), .B(KEYINPUT11), .ZN(new_n277));
  XNOR2_X1  g076(.A(new_n276), .B(new_n277), .ZN(new_n278));
  XNOR2_X1  g077(.A(new_n278), .B(KEYINPUT12), .ZN(new_n279));
  INV_X1    g078(.A(new_n279), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n272), .A2(new_n280), .ZN(new_n281));
  NAND3_X1  g080(.A1(new_n266), .A2(new_n279), .A3(new_n271), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  AND2_X1   g082(.A1(G232gat), .A2(G233gat), .ZN(new_n284));
  NOR2_X1   g083(.A1(new_n284), .A2(KEYINPUT41), .ZN(new_n285));
  XNOR2_X1  g084(.A(G134gat), .B(G162gat), .ZN(new_n286));
  XOR2_X1   g085(.A(new_n285), .B(new_n286), .Z(new_n287));
  INV_X1    g086(.A(new_n287), .ZN(new_n288));
  INV_X1    g087(.A(G190gat), .ZN(new_n289));
  INV_X1    g088(.A(KEYINPUT101), .ZN(new_n290));
  NAND2_X1  g089(.A1(G99gat), .A2(G106gat), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n291), .A2(KEYINPUT8), .ZN(new_n292));
  OR2_X1    g091(.A1(G85gat), .A2(G92gat), .ZN(new_n293));
  AND3_X1   g092(.A1(new_n292), .A2(KEYINPUT100), .A3(new_n293), .ZN(new_n294));
  AOI21_X1  g093(.A(KEYINPUT100), .B1(new_n292), .B2(new_n293), .ZN(new_n295));
  NOR2_X1   g094(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  NAND2_X1  g095(.A1(G85gat), .A2(G92gat), .ZN(new_n297));
  INV_X1    g096(.A(KEYINPUT99), .ZN(new_n298));
  AOI21_X1  g097(.A(new_n297), .B1(new_n298), .B2(KEYINPUT7), .ZN(new_n299));
  NAND2_X1  g098(.A1(KEYINPUT98), .A2(KEYINPUT7), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n300), .A2(KEYINPUT99), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n299), .A2(new_n301), .ZN(new_n302));
  NAND3_X1  g101(.A1(new_n300), .A2(new_n297), .A3(KEYINPUT99), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  XNOR2_X1  g103(.A(G99gat), .B(G106gat), .ZN(new_n305));
  INV_X1    g104(.A(new_n305), .ZN(new_n306));
  NOR3_X1   g105(.A1(new_n296), .A2(new_n304), .A3(new_n306), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n292), .A2(new_n293), .ZN(new_n308));
  INV_X1    g107(.A(KEYINPUT100), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n308), .A2(new_n309), .ZN(new_n310));
  NAND3_X1  g109(.A1(new_n292), .A2(new_n293), .A3(KEYINPUT100), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  AND3_X1   g111(.A1(new_n300), .A2(new_n297), .A3(KEYINPUT99), .ZN(new_n313));
  AOI21_X1  g112(.A(new_n313), .B1(new_n301), .B2(new_n299), .ZN(new_n314));
  AOI21_X1  g113(.A(new_n305), .B1(new_n312), .B2(new_n314), .ZN(new_n315));
  OAI21_X1  g114(.A(new_n290), .B1(new_n307), .B2(new_n315), .ZN(new_n316));
  OAI21_X1  g115(.A(new_n306), .B1(new_n296), .B2(new_n304), .ZN(new_n317));
  NAND3_X1  g116(.A1(new_n312), .A2(new_n305), .A3(new_n314), .ZN(new_n318));
  NAND3_X1  g117(.A1(new_n317), .A2(KEYINPUT101), .A3(new_n318), .ZN(new_n319));
  NAND3_X1  g118(.A1(new_n262), .A2(new_n316), .A3(new_n319), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n284), .A2(KEYINPUT41), .ZN(new_n321));
  AND2_X1   g120(.A1(new_n320), .A2(new_n321), .ZN(new_n322));
  INV_X1    g121(.A(new_n319), .ZN(new_n323));
  AOI21_X1  g122(.A(KEYINPUT101), .B1(new_n317), .B2(new_n318), .ZN(new_n324));
  OAI211_X1 g123(.A(new_n261), .B(new_n255), .C1(new_n323), .C2(new_n324), .ZN(new_n325));
  AOI21_X1  g124(.A(KEYINPUT102), .B1(new_n322), .B2(new_n325), .ZN(new_n326));
  AND4_X1   g125(.A1(KEYINPUT102), .A2(new_n325), .A3(new_n320), .A4(new_n321), .ZN(new_n327));
  OAI21_X1  g126(.A(new_n289), .B1(new_n326), .B2(new_n327), .ZN(new_n328));
  INV_X1    g127(.A(KEYINPUT102), .ZN(new_n329));
  INV_X1    g128(.A(new_n325), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n320), .A2(new_n321), .ZN(new_n331));
  OAI21_X1  g130(.A(new_n329), .B1(new_n330), .B2(new_n331), .ZN(new_n332));
  NAND3_X1  g131(.A1(new_n322), .A2(KEYINPUT102), .A3(new_n325), .ZN(new_n333));
  NAND3_X1  g132(.A1(new_n332), .A2(new_n333), .A3(G190gat), .ZN(new_n334));
  NAND3_X1  g133(.A1(new_n328), .A2(G218gat), .A3(new_n334), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n335), .A2(KEYINPUT97), .ZN(new_n336));
  AOI21_X1  g135(.A(G218gat), .B1(new_n328), .B2(new_n334), .ZN(new_n337));
  OAI21_X1  g136(.A(new_n288), .B1(new_n336), .B2(new_n337), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n328), .A2(new_n334), .ZN(new_n339));
  INV_X1    g138(.A(G218gat), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  NAND4_X1  g140(.A1(new_n341), .A2(KEYINPUT97), .A3(new_n335), .A4(new_n287), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n338), .A2(new_n342), .ZN(new_n343));
  XOR2_X1   g142(.A(G57gat), .B(G64gat), .Z(new_n344));
  INV_X1    g143(.A(G71gat), .ZN(new_n345));
  INV_X1    g144(.A(G78gat), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n345), .A2(new_n346), .ZN(new_n347));
  NAND2_X1  g146(.A1(G71gat), .A2(G78gat), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n347), .A2(new_n348), .ZN(new_n349));
  INV_X1    g148(.A(KEYINPUT9), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n348), .A2(new_n350), .ZN(new_n351));
  NAND3_X1  g150(.A1(new_n344), .A2(new_n349), .A3(new_n351), .ZN(new_n352));
  XNOR2_X1  g151(.A(G57gat), .B(G64gat), .ZN(new_n353));
  OAI211_X1 g152(.A(new_n348), .B(new_n347), .C1(new_n353), .C2(new_n350), .ZN(new_n354));
  AND2_X1   g153(.A1(new_n352), .A2(new_n354), .ZN(new_n355));
  INV_X1    g154(.A(new_n355), .ZN(new_n356));
  XOR2_X1   g155(.A(KEYINPUT96), .B(KEYINPUT21), .Z(new_n357));
  NAND2_X1  g156(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  NAND2_X1  g157(.A1(G231gat), .A2(G233gat), .ZN(new_n359));
  XNOR2_X1  g158(.A(new_n358), .B(new_n359), .ZN(new_n360));
  XNOR2_X1  g159(.A(new_n360), .B(G127gat), .ZN(new_n361));
  AOI21_X1  g160(.A(new_n218), .B1(KEYINPUT21), .B2(new_n355), .ZN(new_n362));
  XOR2_X1   g161(.A(new_n361), .B(new_n362), .Z(new_n363));
  XNOR2_X1  g162(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n364));
  INV_X1    g163(.A(G155gat), .ZN(new_n365));
  XNOR2_X1  g164(.A(new_n364), .B(new_n365), .ZN(new_n366));
  XOR2_X1   g165(.A(G183gat), .B(G211gat), .Z(new_n367));
  XNOR2_X1  g166(.A(new_n366), .B(new_n367), .ZN(new_n368));
  XNOR2_X1  g167(.A(new_n363), .B(new_n368), .ZN(new_n369));
  NOR2_X1   g168(.A1(new_n343), .A2(new_n369), .ZN(new_n370));
  OR2_X1    g169(.A1(new_n305), .A2(KEYINPUT103), .ZN(new_n371));
  AND3_X1   g170(.A1(new_n352), .A2(new_n354), .A3(new_n371), .ZN(new_n372));
  INV_X1    g171(.A(new_n372), .ZN(new_n373));
  OAI21_X1  g172(.A(new_n373), .B1(new_n307), .B2(new_n315), .ZN(new_n374));
  INV_X1    g173(.A(KEYINPUT10), .ZN(new_n375));
  NAND3_X1  g174(.A1(new_n317), .A2(new_n372), .A3(new_n318), .ZN(new_n376));
  NAND3_X1  g175(.A1(new_n374), .A2(new_n375), .A3(new_n376), .ZN(new_n377));
  NOR2_X1   g176(.A1(new_n356), .A2(new_n375), .ZN(new_n378));
  NAND3_X1  g177(.A1(new_n316), .A2(new_n319), .A3(new_n378), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n377), .A2(new_n379), .ZN(new_n380));
  NAND2_X1  g179(.A1(G230gat), .A2(G233gat), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n380), .A2(new_n381), .ZN(new_n382));
  AOI21_X1  g181(.A(new_n381), .B1(new_n374), .B2(new_n376), .ZN(new_n383));
  INV_X1    g182(.A(new_n383), .ZN(new_n384));
  XNOR2_X1  g183(.A(G120gat), .B(G148gat), .ZN(new_n385));
  XNOR2_X1  g184(.A(G176gat), .B(G204gat), .ZN(new_n386));
  XOR2_X1   g185(.A(new_n385), .B(new_n386), .Z(new_n387));
  NAND3_X1  g186(.A1(new_n382), .A2(new_n384), .A3(new_n387), .ZN(new_n388));
  INV_X1    g187(.A(new_n387), .ZN(new_n389));
  INV_X1    g188(.A(new_n381), .ZN(new_n390));
  AOI21_X1  g189(.A(new_n390), .B1(new_n377), .B2(new_n379), .ZN(new_n391));
  OAI21_X1  g190(.A(new_n389), .B1(new_n391), .B2(new_n383), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n388), .A2(new_n392), .ZN(new_n393));
  INV_X1    g192(.A(KEYINPUT104), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n393), .A2(new_n394), .ZN(new_n395));
  NAND3_X1  g194(.A1(new_n388), .A2(KEYINPUT104), .A3(new_n392), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n395), .A2(new_n396), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n370), .A2(new_n397), .ZN(new_n398));
  INV_X1    g197(.A(new_n398), .ZN(new_n399));
  INV_X1    g198(.A(KEYINPUT36), .ZN(new_n400));
  INV_X1    g199(.A(KEYINPUT32), .ZN(new_n401));
  XNOR2_X1  g200(.A(G113gat), .B(G120gat), .ZN(new_n402));
  NOR2_X1   g201(.A1(new_n402), .A2(KEYINPUT1), .ZN(new_n403));
  INV_X1    g202(.A(G127gat), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n404), .A2(G134gat), .ZN(new_n405));
  INV_X1    g204(.A(new_n405), .ZN(new_n406));
  XOR2_X1   g205(.A(KEYINPUT69), .B(G134gat), .Z(new_n407));
  AOI21_X1  g206(.A(new_n406), .B1(new_n407), .B2(G127gat), .ZN(new_n408));
  AOI21_X1  g207(.A(new_n403), .B1(new_n408), .B2(KEYINPUT70), .ZN(new_n409));
  XNOR2_X1  g208(.A(KEYINPUT69), .B(G134gat), .ZN(new_n410));
  OAI21_X1  g209(.A(new_n405), .B1(new_n410), .B2(new_n404), .ZN(new_n411));
  INV_X1    g210(.A(KEYINPUT70), .ZN(new_n412));
  NAND2_X1  g211(.A1(new_n411), .A2(new_n412), .ZN(new_n413));
  INV_X1    g212(.A(G120gat), .ZN(new_n414));
  NAND3_X1  g213(.A1(new_n414), .A2(KEYINPUT71), .A3(G113gat), .ZN(new_n415));
  INV_X1    g214(.A(KEYINPUT1), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n415), .A2(new_n416), .ZN(new_n417));
  INV_X1    g216(.A(G134gat), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n418), .A2(G127gat), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n405), .A2(new_n419), .ZN(new_n420));
  AOI21_X1  g219(.A(new_n417), .B1(KEYINPUT72), .B2(new_n420), .ZN(new_n421));
  INV_X1    g220(.A(new_n420), .ZN(new_n422));
  INV_X1    g221(.A(KEYINPUT72), .ZN(new_n423));
  INV_X1    g222(.A(KEYINPUT71), .ZN(new_n424));
  AOI22_X1  g223(.A1(new_n422), .A2(new_n423), .B1(new_n424), .B2(new_n402), .ZN(new_n425));
  AOI22_X1  g224(.A1(new_n409), .A2(new_n413), .B1(new_n421), .B2(new_n425), .ZN(new_n426));
  NOR2_X1   g225(.A1(G169gat), .A2(G176gat), .ZN(new_n427));
  NAND2_X1  g226(.A1(G169gat), .A2(G176gat), .ZN(new_n428));
  AOI21_X1  g227(.A(new_n427), .B1(KEYINPUT23), .B2(new_n428), .ZN(new_n429));
  AND2_X1   g228(.A1(new_n427), .A2(KEYINPUT23), .ZN(new_n430));
  NOR2_X1   g229(.A1(new_n429), .A2(new_n430), .ZN(new_n431));
  OAI21_X1  g230(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n432));
  NAND2_X1  g231(.A1(G183gat), .A2(G190gat), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n432), .A2(new_n433), .ZN(new_n434));
  INV_X1    g233(.A(KEYINPUT64), .ZN(new_n435));
  NAND4_X1  g234(.A1(new_n435), .A2(KEYINPUT24), .A3(G183gat), .A4(G190gat), .ZN(new_n436));
  NAND3_X1  g235(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n437), .A2(KEYINPUT64), .ZN(new_n438));
  NAND3_X1  g237(.A1(new_n434), .A2(new_n436), .A3(new_n438), .ZN(new_n439));
  AOI21_X1  g238(.A(KEYINPUT25), .B1(new_n431), .B2(new_n439), .ZN(new_n440));
  INV_X1    g239(.A(KEYINPUT66), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n437), .A2(new_n441), .ZN(new_n442));
  NAND4_X1  g241(.A1(KEYINPUT66), .A2(KEYINPUT24), .A3(G183gat), .A4(G190gat), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  AOI21_X1  g243(.A(KEYINPUT67), .B1(new_n444), .B2(new_n434), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n427), .A2(KEYINPUT65), .ZN(new_n446));
  INV_X1    g245(.A(KEYINPUT65), .ZN(new_n447));
  OAI21_X1  g246(.A(new_n447), .B1(G169gat), .B2(G176gat), .ZN(new_n448));
  NAND3_X1  g247(.A1(new_n446), .A2(KEYINPUT23), .A3(new_n448), .ZN(new_n449));
  INV_X1    g248(.A(KEYINPUT25), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n428), .A2(KEYINPUT23), .ZN(new_n451));
  INV_X1    g250(.A(G169gat), .ZN(new_n452));
  INV_X1    g251(.A(G176gat), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  AOI21_X1  g253(.A(new_n450), .B1(new_n451), .B2(new_n454), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n449), .A2(new_n455), .ZN(new_n456));
  NOR2_X1   g255(.A1(new_n445), .A2(new_n456), .ZN(new_n457));
  AOI22_X1  g256(.A1(new_n442), .A2(new_n443), .B1(new_n433), .B2(new_n432), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n458), .A2(KEYINPUT67), .ZN(new_n459));
  AOI21_X1  g258(.A(new_n440), .B1(new_n457), .B2(new_n459), .ZN(new_n460));
  AOI21_X1  g259(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n461));
  OR3_X1    g260(.A1(new_n461), .A2(new_n427), .A3(KEYINPUT68), .ZN(new_n462));
  OAI21_X1  g261(.A(KEYINPUT68), .B1(new_n461), .B2(new_n427), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n446), .A2(new_n448), .ZN(new_n464));
  OAI211_X1 g263(.A(new_n462), .B(new_n463), .C1(KEYINPUT26), .C2(new_n464), .ZN(new_n465));
  XNOR2_X1  g264(.A(KEYINPUT27), .B(G183gat), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n466), .A2(new_n289), .ZN(new_n467));
  OR2_X1    g266(.A1(new_n467), .A2(KEYINPUT28), .ZN(new_n468));
  AOI22_X1  g267(.A1(new_n467), .A2(KEYINPUT28), .B1(G183gat), .B2(G190gat), .ZN(new_n469));
  AND3_X1   g268(.A1(new_n465), .A2(new_n468), .A3(new_n469), .ZN(new_n470));
  OAI21_X1  g269(.A(new_n426), .B1(new_n460), .B2(new_n470), .ZN(new_n471));
  INV_X1    g270(.A(G227gat), .ZN(new_n472));
  INV_X1    g271(.A(G233gat), .ZN(new_n473));
  NOR2_X1   g272(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n431), .A2(new_n439), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n475), .A2(new_n450), .ZN(new_n476));
  INV_X1    g275(.A(new_n459), .ZN(new_n477));
  OAI211_X1 g276(.A(new_n449), .B(new_n455), .C1(new_n458), .C2(KEYINPUT67), .ZN(new_n478));
  OAI21_X1  g277(.A(new_n476), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n425), .A2(new_n421), .ZN(new_n480));
  OAI22_X1  g279(.A1(new_n411), .A2(new_n412), .B1(KEYINPUT1), .B2(new_n402), .ZN(new_n481));
  NAND2_X1  g280(.A1(new_n407), .A2(G127gat), .ZN(new_n482));
  AOI21_X1  g281(.A(KEYINPUT70), .B1(new_n482), .B2(new_n405), .ZN(new_n483));
  OAI21_X1  g282(.A(new_n480), .B1(new_n481), .B2(new_n483), .ZN(new_n484));
  NAND3_X1  g283(.A1(new_n465), .A2(new_n468), .A3(new_n469), .ZN(new_n485));
  NAND3_X1  g284(.A1(new_n479), .A2(new_n484), .A3(new_n485), .ZN(new_n486));
  NAND3_X1  g285(.A1(new_n471), .A2(new_n474), .A3(new_n486), .ZN(new_n487));
  INV_X1    g286(.A(KEYINPUT73), .ZN(new_n488));
  NAND2_X1  g287(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  NAND4_X1  g288(.A1(new_n471), .A2(new_n486), .A3(KEYINPUT73), .A4(new_n474), .ZN(new_n490));
  AOI21_X1  g289(.A(new_n401), .B1(new_n489), .B2(new_n490), .ZN(new_n491));
  INV_X1    g290(.A(KEYINPUT33), .ZN(new_n492));
  XNOR2_X1  g291(.A(G15gat), .B(G43gat), .ZN(new_n493));
  XNOR2_X1  g292(.A(G71gat), .B(G99gat), .ZN(new_n494));
  XNOR2_X1  g293(.A(new_n493), .B(new_n494), .ZN(new_n495));
  OAI21_X1  g294(.A(new_n491), .B1(new_n492), .B2(new_n495), .ZN(new_n496));
  AOI21_X1  g295(.A(KEYINPUT33), .B1(new_n489), .B2(new_n490), .ZN(new_n497));
  INV_X1    g296(.A(KEYINPUT74), .ZN(new_n498));
  NOR4_X1   g297(.A1(new_n491), .A2(new_n497), .A3(new_n498), .A4(new_n495), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n489), .A2(new_n490), .ZN(new_n500));
  AOI21_X1  g299(.A(new_n495), .B1(new_n500), .B2(KEYINPUT32), .ZN(new_n501));
  INV_X1    g300(.A(new_n497), .ZN(new_n502));
  AOI21_X1  g301(.A(KEYINPUT74), .B1(new_n501), .B2(new_n502), .ZN(new_n503));
  OAI21_X1  g302(.A(new_n496), .B1(new_n499), .B2(new_n503), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n471), .A2(new_n486), .ZN(new_n505));
  OAI21_X1  g304(.A(new_n505), .B1(new_n472), .B2(new_n473), .ZN(new_n506));
  XOR2_X1   g305(.A(new_n506), .B(KEYINPUT34), .Z(new_n507));
  INV_X1    g306(.A(new_n507), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n504), .A2(new_n508), .ZN(new_n509));
  OAI211_X1 g308(.A(new_n507), .B(new_n496), .C1(new_n499), .C2(new_n503), .ZN(new_n510));
  AOI21_X1  g309(.A(new_n400), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  INV_X1    g310(.A(KEYINPUT75), .ZN(new_n512));
  NAND3_X1  g311(.A1(new_n509), .A2(new_n512), .A3(new_n510), .ZN(new_n513));
  NAND3_X1  g312(.A1(new_n504), .A2(KEYINPUT75), .A3(new_n508), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  AOI21_X1  g314(.A(new_n511), .B1(new_n515), .B2(new_n400), .ZN(new_n516));
  XOR2_X1   g315(.A(G8gat), .B(G36gat), .Z(new_n517));
  XNOR2_X1  g316(.A(G64gat), .B(G92gat), .ZN(new_n518));
  XNOR2_X1  g317(.A(new_n517), .B(new_n518), .ZN(new_n519));
  XNOR2_X1  g318(.A(KEYINPUT77), .B(KEYINPUT78), .ZN(new_n520));
  XOR2_X1   g319(.A(new_n519), .B(new_n520), .Z(new_n521));
  XNOR2_X1  g320(.A(G197gat), .B(G204gat), .ZN(new_n522));
  INV_X1    g321(.A(G211gat), .ZN(new_n523));
  NOR2_X1   g322(.A1(new_n523), .A2(new_n340), .ZN(new_n524));
  OAI21_X1  g323(.A(new_n522), .B1(KEYINPUT22), .B2(new_n524), .ZN(new_n525));
  INV_X1    g324(.A(KEYINPUT76), .ZN(new_n526));
  XOR2_X1   g325(.A(G211gat), .B(G218gat), .Z(new_n527));
  NAND3_X1  g326(.A1(new_n525), .A2(new_n526), .A3(new_n527), .ZN(new_n528));
  XNOR2_X1  g327(.A(new_n525), .B(new_n527), .ZN(new_n529));
  OAI21_X1  g328(.A(new_n528), .B1(new_n529), .B2(new_n526), .ZN(new_n530));
  INV_X1    g329(.A(G226gat), .ZN(new_n531));
  NOR2_X1   g330(.A1(new_n531), .A2(new_n473), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n479), .A2(new_n485), .ZN(new_n533));
  INV_X1    g332(.A(KEYINPUT29), .ZN(new_n534));
  AOI21_X1  g333(.A(new_n532), .B1(new_n533), .B2(new_n534), .ZN(new_n535));
  INV_X1    g334(.A(new_n535), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n533), .A2(new_n532), .ZN(new_n537));
  AOI21_X1  g336(.A(new_n530), .B1(new_n536), .B2(new_n537), .ZN(new_n538));
  INV_X1    g337(.A(new_n537), .ZN(new_n539));
  INV_X1    g338(.A(new_n530), .ZN(new_n540));
  NOR3_X1   g339(.A1(new_n539), .A2(new_n535), .A3(new_n540), .ZN(new_n541));
  OAI21_X1  g340(.A(new_n521), .B1(new_n538), .B2(new_n541), .ZN(new_n542));
  INV_X1    g341(.A(KEYINPUT30), .ZN(new_n543));
  NOR2_X1   g342(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  NAND3_X1  g343(.A1(new_n536), .A2(new_n530), .A3(new_n537), .ZN(new_n545));
  OAI21_X1  g344(.A(new_n540), .B1(new_n539), .B2(new_n535), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  NOR2_X1   g346(.A1(new_n547), .A2(new_n521), .ZN(new_n548));
  NOR2_X1   g347(.A1(new_n544), .A2(new_n548), .ZN(new_n549));
  INV_X1    g348(.A(KEYINPUT79), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n542), .A2(new_n550), .ZN(new_n551));
  NAND3_X1  g350(.A1(new_n547), .A2(KEYINPUT79), .A3(new_n521), .ZN(new_n552));
  NAND3_X1  g351(.A1(new_n551), .A2(new_n552), .A3(new_n543), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n549), .A2(new_n553), .ZN(new_n554));
  INV_X1    g353(.A(KEYINPUT80), .ZN(new_n555));
  XOR2_X1   g354(.A(G141gat), .B(G148gat), .Z(new_n556));
  INV_X1    g355(.A(G162gat), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n365), .A2(new_n557), .ZN(new_n558));
  NAND2_X1  g357(.A1(G155gat), .A2(G162gat), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n559), .A2(KEYINPUT2), .ZN(new_n561));
  NAND3_X1  g360(.A1(new_n556), .A2(new_n560), .A3(new_n561), .ZN(new_n562));
  XNOR2_X1  g361(.A(G141gat), .B(G148gat), .ZN(new_n563));
  OAI211_X1 g362(.A(new_n559), .B(new_n558), .C1(new_n563), .C2(KEYINPUT2), .ZN(new_n564));
  NAND2_X1  g363(.A1(new_n562), .A2(new_n564), .ZN(new_n565));
  OAI21_X1  g364(.A(new_n555), .B1(new_n565), .B2(KEYINPUT3), .ZN(new_n566));
  INV_X1    g365(.A(KEYINPUT3), .ZN(new_n567));
  NAND4_X1  g366(.A1(new_n562), .A2(new_n564), .A3(KEYINPUT80), .A4(new_n567), .ZN(new_n568));
  NAND2_X1  g367(.A1(new_n566), .A2(new_n568), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n565), .A2(KEYINPUT3), .ZN(new_n570));
  NAND3_X1  g369(.A1(new_n569), .A2(new_n570), .A3(new_n484), .ZN(new_n571));
  INV_X1    g370(.A(new_n565), .ZN(new_n572));
  NAND3_X1  g371(.A1(new_n426), .A2(KEYINPUT4), .A3(new_n572), .ZN(new_n573));
  INV_X1    g372(.A(KEYINPUT4), .ZN(new_n574));
  OAI21_X1  g373(.A(new_n574), .B1(new_n484), .B2(new_n565), .ZN(new_n575));
  NAND2_X1  g374(.A1(G225gat), .A2(G233gat), .ZN(new_n576));
  NAND4_X1  g375(.A1(new_n571), .A2(new_n573), .A3(new_n575), .A4(new_n576), .ZN(new_n577));
  NAND2_X1  g376(.A1(new_n577), .A2(KEYINPUT81), .ZN(new_n578));
  XNOR2_X1  g377(.A(new_n484), .B(new_n565), .ZN(new_n579));
  INV_X1    g378(.A(new_n576), .ZN(new_n580));
  NAND2_X1  g379(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  NAND3_X1  g380(.A1(new_n578), .A2(KEYINPUT5), .A3(new_n581), .ZN(new_n582));
  XNOR2_X1  g381(.A(new_n484), .B(new_n572), .ZN(new_n583));
  OAI21_X1  g382(.A(KEYINPUT5), .B1(new_n583), .B2(new_n576), .ZN(new_n584));
  NAND3_X1  g383(.A1(new_n584), .A2(KEYINPUT81), .A3(new_n577), .ZN(new_n585));
  XNOR2_X1  g384(.A(G1gat), .B(G29gat), .ZN(new_n586));
  XNOR2_X1  g385(.A(new_n586), .B(KEYINPUT0), .ZN(new_n587));
  XNOR2_X1  g386(.A(G57gat), .B(G85gat), .ZN(new_n588));
  XOR2_X1   g387(.A(new_n587), .B(new_n588), .Z(new_n589));
  INV_X1    g388(.A(new_n589), .ZN(new_n590));
  AND4_X1   g389(.A1(KEYINPUT6), .A2(new_n582), .A3(new_n585), .A4(new_n590), .ZN(new_n591));
  AND2_X1   g390(.A1(new_n582), .A2(new_n585), .ZN(new_n592));
  NAND2_X1  g391(.A1(new_n592), .A2(new_n590), .ZN(new_n593));
  NAND2_X1  g392(.A1(new_n582), .A2(new_n585), .ZN(new_n594));
  AOI21_X1  g393(.A(KEYINPUT6), .B1(new_n594), .B2(new_n589), .ZN(new_n595));
  AOI21_X1  g394(.A(new_n591), .B1(new_n593), .B2(new_n595), .ZN(new_n596));
  NOR2_X1   g395(.A1(new_n554), .A2(new_n596), .ZN(new_n597));
  NAND2_X1  g396(.A1(G228gat), .A2(G233gat), .ZN(new_n598));
  NAND2_X1  g397(.A1(new_n569), .A2(new_n534), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n599), .A2(new_n530), .ZN(new_n600));
  INV_X1    g399(.A(new_n600), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n529), .A2(new_n534), .ZN(new_n602));
  AOI21_X1  g401(.A(new_n572), .B1(new_n602), .B2(new_n567), .ZN(new_n603));
  OAI21_X1  g402(.A(new_n598), .B1(new_n601), .B2(new_n603), .ZN(new_n604));
  OAI21_X1  g403(.A(new_n567), .B1(new_n530), .B2(KEYINPUT29), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n605), .A2(new_n565), .ZN(new_n606));
  NAND4_X1  g405(.A1(new_n606), .A2(new_n600), .A3(G228gat), .A4(G233gat), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n604), .A2(new_n607), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n608), .A2(G22gat), .ZN(new_n609));
  NAND3_X1  g408(.A1(new_n604), .A2(new_n607), .A3(new_n209), .ZN(new_n610));
  NAND3_X1  g409(.A1(new_n609), .A2(KEYINPUT83), .A3(new_n610), .ZN(new_n611));
  XNOR2_X1  g410(.A(G78gat), .B(G106gat), .ZN(new_n612));
  XNOR2_X1  g411(.A(new_n612), .B(KEYINPUT82), .ZN(new_n613));
  XOR2_X1   g412(.A(KEYINPUT31), .B(G50gat), .Z(new_n614));
  XNOR2_X1  g413(.A(new_n613), .B(new_n614), .ZN(new_n615));
  AOI21_X1  g414(.A(new_n209), .B1(new_n604), .B2(new_n607), .ZN(new_n616));
  INV_X1    g415(.A(KEYINPUT83), .ZN(new_n617));
  AOI21_X1  g416(.A(new_n615), .B1(new_n616), .B2(new_n617), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n611), .A2(new_n618), .ZN(new_n619));
  NAND3_X1  g418(.A1(new_n609), .A2(new_n615), .A3(new_n610), .ZN(new_n620));
  INV_X1    g419(.A(KEYINPUT84), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  NAND4_X1  g421(.A1(new_n609), .A2(KEYINPUT84), .A3(new_n615), .A4(new_n610), .ZN(new_n623));
  NAND3_X1  g422(.A1(new_n619), .A2(new_n622), .A3(new_n623), .ZN(new_n624));
  NOR2_X1   g423(.A1(new_n597), .A2(new_n624), .ZN(new_n625));
  INV_X1    g424(.A(new_n625), .ZN(new_n626));
  AOI21_X1  g425(.A(KEYINPUT85), .B1(new_n516), .B2(new_n626), .ZN(new_n627));
  AOI21_X1  g426(.A(KEYINPUT36), .B1(new_n513), .B2(new_n514), .ZN(new_n628));
  INV_X1    g427(.A(KEYINPUT85), .ZN(new_n629));
  NOR4_X1   g428(.A1(new_n628), .A2(new_n629), .A3(new_n625), .A4(new_n511), .ZN(new_n630));
  NAND3_X1  g429(.A1(new_n571), .A2(new_n575), .A3(new_n573), .ZN(new_n631));
  NAND2_X1  g430(.A1(new_n631), .A2(new_n580), .ZN(new_n632));
  OR2_X1    g431(.A1(new_n632), .A2(KEYINPUT39), .ZN(new_n633));
  OAI211_X1 g432(.A(new_n632), .B(KEYINPUT39), .C1(new_n580), .C2(new_n579), .ZN(new_n634));
  XOR2_X1   g433(.A(new_n589), .B(KEYINPUT86), .Z(new_n635));
  INV_X1    g434(.A(new_n635), .ZN(new_n636));
  NAND3_X1  g435(.A1(new_n633), .A2(new_n634), .A3(new_n636), .ZN(new_n637));
  INV_X1    g436(.A(KEYINPUT40), .ZN(new_n638));
  NAND2_X1  g437(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n592), .A2(new_n635), .ZN(new_n640));
  OR2_X1    g439(.A1(new_n637), .A2(new_n638), .ZN(new_n641));
  NAND4_X1  g440(.A1(new_n554), .A2(new_n639), .A3(new_n640), .A4(new_n641), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n642), .A2(new_n624), .ZN(new_n643));
  INV_X1    g442(.A(KEYINPUT87), .ZN(new_n644));
  AOI21_X1  g443(.A(new_n591), .B1(new_n640), .B2(new_n595), .ZN(new_n645));
  INV_X1    g444(.A(new_n645), .ZN(new_n646));
  AND2_X1   g445(.A1(new_n551), .A2(new_n552), .ZN(new_n647));
  NOR2_X1   g446(.A1(new_n538), .A2(new_n541), .ZN(new_n648));
  AOI21_X1  g447(.A(new_n521), .B1(new_n648), .B2(KEYINPUT37), .ZN(new_n649));
  INV_X1    g448(.A(KEYINPUT38), .ZN(new_n650));
  INV_X1    g449(.A(KEYINPUT37), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n547), .A2(new_n651), .ZN(new_n652));
  NAND3_X1  g451(.A1(new_n649), .A2(new_n650), .A3(new_n652), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n647), .A2(new_n653), .ZN(new_n654));
  OAI21_X1  g453(.A(new_n644), .B1(new_n646), .B2(new_n654), .ZN(new_n655));
  NAND4_X1  g454(.A1(new_n645), .A2(KEYINPUT87), .A3(new_n647), .A4(new_n653), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  INV_X1    g456(.A(new_n649), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n658), .A2(KEYINPUT88), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n659), .A2(new_n652), .ZN(new_n660));
  NOR2_X1   g459(.A1(new_n658), .A2(KEYINPUT88), .ZN(new_n661));
  OAI21_X1  g460(.A(KEYINPUT38), .B1(new_n660), .B2(new_n661), .ZN(new_n662));
  AOI21_X1  g461(.A(new_n643), .B1(new_n657), .B2(new_n662), .ZN(new_n663));
  NOR3_X1   g462(.A1(new_n627), .A2(new_n630), .A3(new_n663), .ZN(new_n664));
  NAND4_X1  g463(.A1(new_n597), .A2(new_n509), .A3(new_n510), .A4(new_n624), .ZN(new_n665));
  AND2_X1   g464(.A1(new_n665), .A2(KEYINPUT35), .ZN(new_n666));
  INV_X1    g465(.A(new_n554), .ZN(new_n667));
  INV_X1    g466(.A(KEYINPUT35), .ZN(new_n668));
  NAND4_X1  g467(.A1(new_n667), .A2(new_n624), .A3(new_n646), .A4(new_n668), .ZN(new_n669));
  AOI21_X1  g468(.A(new_n669), .B1(new_n514), .B2(new_n513), .ZN(new_n670));
  NOR2_X1   g469(.A1(new_n666), .A2(new_n670), .ZN(new_n671));
  OAI211_X1 g470(.A(new_n283), .B(new_n399), .C1(new_n664), .C2(new_n671), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n672), .A2(KEYINPUT105), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n515), .A2(new_n400), .ZN(new_n674));
  INV_X1    g473(.A(new_n511), .ZN(new_n675));
  NAND3_X1  g474(.A1(new_n674), .A2(new_n626), .A3(new_n675), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n676), .A2(new_n629), .ZN(new_n677));
  NAND3_X1  g476(.A1(new_n516), .A2(KEYINPUT85), .A3(new_n626), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n657), .A2(new_n662), .ZN(new_n679));
  INV_X1    g478(.A(new_n643), .ZN(new_n680));
  NAND2_X1  g479(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  NAND3_X1  g480(.A1(new_n677), .A2(new_n678), .A3(new_n681), .ZN(new_n682));
  INV_X1    g481(.A(new_n671), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  INV_X1    g483(.A(KEYINPUT105), .ZN(new_n685));
  NAND4_X1  g484(.A1(new_n684), .A2(new_n685), .A3(new_n283), .A4(new_n399), .ZN(new_n686));
  NAND2_X1  g485(.A1(new_n673), .A2(new_n686), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n687), .A2(new_n596), .ZN(new_n688));
  XNOR2_X1  g487(.A(new_n688), .B(G1gat), .ZN(G1324gat));
  AOI21_X1  g488(.A(new_n215), .B1(new_n687), .B2(new_n554), .ZN(new_n690));
  XNOR2_X1  g489(.A(KEYINPUT16), .B(G8gat), .ZN(new_n691));
  AOI211_X1 g490(.A(new_n667), .B(new_n691), .C1(new_n673), .C2(new_n686), .ZN(new_n692));
  OAI21_X1  g491(.A(KEYINPUT42), .B1(new_n690), .B2(new_n692), .ZN(new_n693));
  OAI21_X1  g492(.A(new_n693), .B1(KEYINPUT42), .B2(new_n692), .ZN(G1325gat));
  NAND3_X1  g493(.A1(new_n687), .A2(new_n207), .A3(new_n515), .ZN(new_n695));
  INV_X1    g494(.A(KEYINPUT106), .ZN(new_n696));
  NAND2_X1  g495(.A1(new_n516), .A2(new_n696), .ZN(new_n697));
  OAI21_X1  g496(.A(KEYINPUT106), .B1(new_n628), .B2(new_n511), .ZN(new_n698));
  NAND2_X1  g497(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  INV_X1    g498(.A(new_n699), .ZN(new_n700));
  AOI21_X1  g499(.A(new_n700), .B1(new_n673), .B2(new_n686), .ZN(new_n701));
  OAI21_X1  g500(.A(new_n695), .B1(new_n701), .B2(new_n207), .ZN(G1326gat));
  INV_X1    g501(.A(KEYINPUT107), .ZN(new_n703));
  INV_X1    g502(.A(new_n624), .ZN(new_n704));
  AOI21_X1  g503(.A(new_n703), .B1(new_n687), .B2(new_n704), .ZN(new_n705));
  AOI211_X1 g504(.A(KEYINPUT107), .B(new_n624), .C1(new_n673), .C2(new_n686), .ZN(new_n706));
  XNOR2_X1  g505(.A(KEYINPUT43), .B(G22gat), .ZN(new_n707));
  INV_X1    g506(.A(new_n707), .ZN(new_n708));
  NOR3_X1   g507(.A1(new_n705), .A2(new_n706), .A3(new_n708), .ZN(new_n709));
  AND3_X1   g508(.A1(new_n266), .A2(new_n279), .A3(new_n271), .ZN(new_n710));
  AOI21_X1  g509(.A(new_n279), .B1(new_n266), .B2(new_n271), .ZN(new_n711));
  NOR2_X1   g510(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  AOI21_X1  g511(.A(new_n712), .B1(new_n682), .B2(new_n683), .ZN(new_n713));
  AOI21_X1  g512(.A(new_n685), .B1(new_n713), .B2(new_n399), .ZN(new_n714));
  AOI21_X1  g513(.A(new_n663), .B1(new_n676), .B2(new_n629), .ZN(new_n715));
  AOI21_X1  g514(.A(new_n671), .B1(new_n715), .B2(new_n678), .ZN(new_n716));
  NOR4_X1   g515(.A1(new_n716), .A2(KEYINPUT105), .A3(new_n712), .A4(new_n398), .ZN(new_n717));
  OAI21_X1  g516(.A(new_n704), .B1(new_n714), .B2(new_n717), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n718), .A2(KEYINPUT107), .ZN(new_n719));
  NAND3_X1  g518(.A1(new_n687), .A2(new_n703), .A3(new_n704), .ZN(new_n720));
  AOI21_X1  g519(.A(new_n707), .B1(new_n719), .B2(new_n720), .ZN(new_n721));
  NOR2_X1   g520(.A1(new_n709), .A2(new_n721), .ZN(G1327gat));
  NAND2_X1  g521(.A1(new_n369), .A2(new_n397), .ZN(new_n723));
  AND2_X1   g522(.A1(new_n338), .A2(new_n342), .ZN(new_n724));
  NOR2_X1   g523(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  AND2_X1   g524(.A1(new_n713), .A2(new_n725), .ZN(new_n726));
  NAND3_X1  g525(.A1(new_n726), .A2(new_n225), .A3(new_n596), .ZN(new_n727));
  XNOR2_X1  g526(.A(new_n727), .B(KEYINPUT45), .ZN(new_n728));
  NAND4_X1  g527(.A1(new_n697), .A2(new_n626), .A3(new_n681), .A4(new_n698), .ZN(new_n729));
  INV_X1    g528(.A(KEYINPUT109), .ZN(new_n730));
  OAI21_X1  g529(.A(new_n730), .B1(new_n666), .B2(new_n670), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n665), .A2(KEYINPUT35), .ZN(new_n732));
  INV_X1    g531(.A(new_n515), .ZN(new_n733));
  OAI211_X1 g532(.A(KEYINPUT109), .B(new_n732), .C1(new_n733), .C2(new_n669), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n731), .A2(new_n734), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n729), .A2(new_n735), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n736), .A2(new_n343), .ZN(new_n737));
  INV_X1    g536(.A(KEYINPUT44), .ZN(new_n738));
  NAND2_X1  g537(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  NAND3_X1  g538(.A1(new_n684), .A2(KEYINPUT44), .A3(new_n343), .ZN(new_n740));
  AND2_X1   g539(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  OAI21_X1  g540(.A(KEYINPUT108), .B1(new_n710), .B2(new_n711), .ZN(new_n742));
  INV_X1    g541(.A(KEYINPUT108), .ZN(new_n743));
  NAND3_X1  g542(.A1(new_n281), .A2(new_n743), .A3(new_n282), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n742), .A2(new_n744), .ZN(new_n745));
  INV_X1    g544(.A(new_n745), .ZN(new_n746));
  NOR2_X1   g545(.A1(new_n723), .A2(new_n746), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n741), .A2(new_n747), .ZN(new_n748));
  INV_X1    g547(.A(new_n596), .ZN(new_n749));
  OAI21_X1  g548(.A(G29gat), .B1(new_n748), .B2(new_n749), .ZN(new_n750));
  NAND2_X1  g549(.A1(new_n728), .A2(new_n750), .ZN(G1328gat));
  NAND3_X1  g550(.A1(new_n726), .A2(new_n226), .A3(new_n554), .ZN(new_n752));
  XOR2_X1   g551(.A(new_n752), .B(KEYINPUT46), .Z(new_n753));
  OAI21_X1  g552(.A(G36gat), .B1(new_n748), .B2(new_n667), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n753), .A2(new_n754), .ZN(G1329gat));
  NAND4_X1  g554(.A1(new_n739), .A2(new_n740), .A3(new_n699), .A4(new_n747), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n756), .A2(G43gat), .ZN(new_n757));
  INV_X1    g556(.A(KEYINPUT111), .ZN(new_n758));
  AOI21_X1  g557(.A(KEYINPUT47), .B1(new_n757), .B2(new_n758), .ZN(new_n759));
  NOR2_X1   g558(.A1(new_n733), .A2(G43gat), .ZN(new_n760));
  NAND3_X1  g559(.A1(new_n713), .A2(new_n725), .A3(new_n760), .ZN(new_n761));
  INV_X1    g560(.A(KEYINPUT110), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  NAND4_X1  g562(.A1(new_n713), .A2(KEYINPUT110), .A3(new_n725), .A4(new_n760), .ZN(new_n764));
  NAND2_X1  g563(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  NAND2_X1  g564(.A1(new_n757), .A2(new_n765), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n759), .A2(new_n766), .ZN(new_n767));
  OAI211_X1 g566(.A(new_n757), .B(new_n765), .C1(new_n758), .C2(KEYINPUT47), .ZN(new_n768));
  NAND2_X1  g567(.A1(new_n767), .A2(new_n768), .ZN(G1330gat));
  NOR2_X1   g568(.A1(new_n624), .A2(new_n219), .ZN(new_n770));
  NAND4_X1  g569(.A1(new_n739), .A2(new_n740), .A3(new_n747), .A4(new_n770), .ZN(new_n771));
  NAND3_X1  g570(.A1(new_n713), .A2(new_n704), .A3(new_n725), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n772), .A2(new_n219), .ZN(new_n773));
  INV_X1    g572(.A(KEYINPUT48), .ZN(new_n774));
  NAND3_X1  g573(.A1(new_n771), .A2(new_n773), .A3(new_n774), .ZN(new_n775));
  INV_X1    g574(.A(KEYINPUT112), .ZN(new_n776));
  AND2_X1   g575(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  NOR2_X1   g576(.A1(new_n775), .A2(new_n776), .ZN(new_n778));
  NAND2_X1  g577(.A1(new_n771), .A2(new_n773), .ZN(new_n779));
  AOI21_X1  g578(.A(KEYINPUT113), .B1(new_n779), .B2(KEYINPUT48), .ZN(new_n780));
  INV_X1    g579(.A(KEYINPUT113), .ZN(new_n781));
  AOI211_X1 g580(.A(new_n781), .B(new_n774), .C1(new_n771), .C2(new_n773), .ZN(new_n782));
  OAI22_X1  g581(.A1(new_n777), .A2(new_n778), .B1(new_n780), .B2(new_n782), .ZN(G1331gat));
  INV_X1    g582(.A(new_n397), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n746), .A2(new_n784), .ZN(new_n785));
  NOR3_X1   g584(.A1(new_n785), .A2(new_n369), .A3(new_n343), .ZN(new_n786));
  NAND2_X1  g585(.A1(new_n736), .A2(new_n786), .ZN(new_n787));
  INV_X1    g586(.A(new_n787), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n788), .A2(new_n596), .ZN(new_n789));
  XNOR2_X1  g588(.A(new_n789), .B(G57gat), .ZN(G1332gat));
  NOR2_X1   g589(.A1(new_n787), .A2(new_n667), .ZN(new_n791));
  NOR2_X1   g590(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n792));
  AND2_X1   g591(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n793));
  OAI21_X1  g592(.A(new_n791), .B1(new_n792), .B2(new_n793), .ZN(new_n794));
  OAI21_X1  g593(.A(new_n794), .B1(new_n791), .B2(new_n792), .ZN(G1333gat));
  NAND3_X1  g594(.A1(new_n788), .A2(G71gat), .A3(new_n699), .ZN(new_n796));
  NOR2_X1   g595(.A1(new_n787), .A2(new_n733), .ZN(new_n797));
  AND2_X1   g596(.A1(new_n797), .A2(KEYINPUT114), .ZN(new_n798));
  OAI21_X1  g597(.A(new_n345), .B1(new_n797), .B2(KEYINPUT114), .ZN(new_n799));
  OAI21_X1  g598(.A(new_n796), .B1(new_n798), .B2(new_n799), .ZN(new_n800));
  XNOR2_X1  g599(.A(new_n800), .B(KEYINPUT50), .ZN(G1334gat));
  NOR2_X1   g600(.A1(new_n787), .A2(new_n624), .ZN(new_n802));
  XNOR2_X1  g601(.A(new_n802), .B(new_n346), .ZN(G1335gat));
  INV_X1    g602(.A(new_n369), .ZN(new_n804));
  NOR2_X1   g603(.A1(new_n785), .A2(new_n804), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n741), .A2(new_n805), .ZN(new_n806));
  OAI21_X1  g605(.A(G85gat), .B1(new_n806), .B2(new_n749), .ZN(new_n807));
  AOI21_X1  g606(.A(new_n724), .B1(new_n729), .B2(new_n735), .ZN(new_n808));
  NOR2_X1   g607(.A1(new_n804), .A2(new_n745), .ZN(new_n809));
  AND3_X1   g608(.A1(new_n808), .A2(KEYINPUT51), .A3(new_n809), .ZN(new_n810));
  AOI21_X1  g609(.A(KEYINPUT51), .B1(new_n808), .B2(new_n809), .ZN(new_n811));
  OR2_X1    g610(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  NOR3_X1   g611(.A1(new_n749), .A2(G85gat), .A3(new_n397), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n812), .A2(new_n813), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n807), .A2(new_n814), .ZN(G1336gat));
  NAND4_X1  g614(.A1(new_n739), .A2(new_n740), .A3(new_n554), .A4(new_n805), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n816), .A2(G92gat), .ZN(new_n817));
  NOR3_X1   g616(.A1(new_n667), .A2(G92gat), .A3(new_n397), .ZN(new_n818));
  OAI21_X1  g617(.A(new_n818), .B1(new_n810), .B2(new_n811), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n817), .A2(new_n819), .ZN(new_n820));
  XNOR2_X1  g619(.A(new_n820), .B(KEYINPUT52), .ZN(G1337gat));
  OAI21_X1  g620(.A(G99gat), .B1(new_n806), .B2(new_n700), .ZN(new_n822));
  NOR3_X1   g621(.A1(new_n733), .A2(G99gat), .A3(new_n397), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n812), .A2(new_n823), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n822), .A2(new_n824), .ZN(G1338gat));
  NAND4_X1  g624(.A1(new_n739), .A2(new_n740), .A3(new_n704), .A4(new_n805), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n826), .A2(G106gat), .ZN(new_n827));
  NOR3_X1   g626(.A1(new_n624), .A2(G106gat), .A3(new_n397), .ZN(new_n828));
  OAI21_X1  g627(.A(new_n828), .B1(new_n810), .B2(new_n811), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n827), .A2(new_n829), .ZN(new_n830));
  XNOR2_X1  g629(.A(new_n830), .B(KEYINPUT53), .ZN(G1339gat));
  NOR2_X1   g630(.A1(new_n263), .A2(new_n202), .ZN(new_n832));
  AND3_X1   g631(.A1(new_n247), .A2(new_n251), .A3(new_n204), .ZN(new_n833));
  OAI21_X1  g632(.A(new_n278), .B1(new_n832), .B2(new_n833), .ZN(new_n834));
  NAND2_X1  g633(.A1(new_n282), .A2(new_n834), .ZN(new_n835));
  INV_X1    g634(.A(new_n835), .ZN(new_n836));
  NAND3_X1  g635(.A1(new_n377), .A2(new_n379), .A3(new_n390), .ZN(new_n837));
  NAND3_X1  g636(.A1(new_n382), .A2(KEYINPUT54), .A3(new_n837), .ZN(new_n838));
  INV_X1    g637(.A(KEYINPUT54), .ZN(new_n839));
  AOI21_X1  g638(.A(new_n387), .B1(new_n391), .B2(new_n839), .ZN(new_n840));
  NAND3_X1  g639(.A1(new_n838), .A2(KEYINPUT55), .A3(new_n840), .ZN(new_n841));
  AND2_X1   g640(.A1(new_n841), .A2(new_n388), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n838), .A2(new_n840), .ZN(new_n843));
  INV_X1    g642(.A(KEYINPUT55), .ZN(new_n844));
  AOI21_X1  g643(.A(KEYINPUT115), .B1(new_n843), .B2(new_n844), .ZN(new_n845));
  INV_X1    g644(.A(KEYINPUT115), .ZN(new_n846));
  AOI211_X1 g645(.A(new_n846), .B(KEYINPUT55), .C1(new_n838), .C2(new_n840), .ZN(new_n847));
  OAI21_X1  g646(.A(new_n842), .B1(new_n845), .B2(new_n847), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n848), .A2(KEYINPUT116), .ZN(new_n849));
  INV_X1    g648(.A(KEYINPUT116), .ZN(new_n850));
  OAI211_X1 g649(.A(new_n842), .B(new_n850), .C1(new_n845), .C2(new_n847), .ZN(new_n851));
  AND4_X1   g650(.A1(new_n343), .A2(new_n836), .A3(new_n849), .A4(new_n851), .ZN(new_n852));
  NAND3_X1  g651(.A1(new_n849), .A2(new_n745), .A3(new_n851), .ZN(new_n853));
  NAND4_X1  g652(.A1(new_n395), .A2(new_n282), .A3(new_n396), .A4(new_n834), .ZN(new_n854));
  AOI21_X1  g653(.A(new_n343), .B1(new_n853), .B2(new_n854), .ZN(new_n855));
  OAI21_X1  g654(.A(new_n369), .B1(new_n852), .B2(new_n855), .ZN(new_n856));
  NAND3_X1  g655(.A1(new_n370), .A2(new_n397), .A3(new_n746), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  NAND2_X1  g657(.A1(new_n509), .A2(new_n510), .ZN(new_n859));
  NOR4_X1   g658(.A1(new_n859), .A2(new_n704), .A3(new_n749), .A4(new_n554), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n858), .A2(new_n860), .ZN(new_n861));
  INV_X1    g660(.A(new_n861), .ZN(new_n862));
  AOI21_X1  g661(.A(G113gat), .B1(new_n862), .B2(new_n745), .ZN(new_n863));
  AOI211_X1 g662(.A(new_n704), .B(new_n733), .C1(new_n856), .C2(new_n857), .ZN(new_n864));
  NOR2_X1   g663(.A1(new_n749), .A2(new_n554), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  INV_X1    g665(.A(new_n866), .ZN(new_n867));
  AND2_X1   g666(.A1(new_n283), .A2(G113gat), .ZN(new_n868));
  AOI21_X1  g667(.A(new_n863), .B1(new_n867), .B2(new_n868), .ZN(G1340gat));
  AOI21_X1  g668(.A(G120gat), .B1(new_n862), .B2(new_n784), .ZN(new_n870));
  NOR2_X1   g669(.A1(new_n397), .A2(new_n414), .ZN(new_n871));
  AOI21_X1  g670(.A(new_n870), .B1(new_n867), .B2(new_n871), .ZN(G1341gat));
  OAI21_X1  g671(.A(G127gat), .B1(new_n866), .B2(new_n369), .ZN(new_n873));
  NAND3_X1  g672(.A1(new_n862), .A2(new_n404), .A3(new_n804), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n873), .A2(new_n874), .ZN(G1342gat));
  NOR3_X1   g674(.A1(new_n861), .A2(new_n410), .A3(new_n724), .ZN(new_n876));
  XNOR2_X1  g675(.A(new_n876), .B(KEYINPUT56), .ZN(new_n877));
  OAI21_X1  g676(.A(G134gat), .B1(new_n866), .B2(new_n724), .ZN(new_n878));
  NAND2_X1  g677(.A1(new_n877), .A2(new_n878), .ZN(G1343gat));
  INV_X1    g678(.A(KEYINPUT121), .ZN(new_n880));
  AND3_X1   g679(.A1(new_n697), .A2(new_n698), .A3(new_n865), .ZN(new_n881));
  INV_X1    g680(.A(KEYINPUT119), .ZN(new_n882));
  INV_X1    g681(.A(KEYINPUT57), .ZN(new_n883));
  NOR2_X1   g682(.A1(new_n624), .A2(new_n883), .ZN(new_n884));
  INV_X1    g683(.A(KEYINPUT118), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n843), .A2(new_n844), .ZN(new_n886));
  NAND3_X1  g685(.A1(new_n886), .A2(new_n388), .A3(new_n841), .ZN(new_n887));
  OAI21_X1  g686(.A(new_n854), .B1(new_n712), .B2(new_n887), .ZN(new_n888));
  NAND2_X1  g687(.A1(new_n888), .A2(KEYINPUT117), .ZN(new_n889));
  INV_X1    g688(.A(KEYINPUT117), .ZN(new_n890));
  OAI211_X1 g689(.A(new_n890), .B(new_n854), .C1(new_n712), .C2(new_n887), .ZN(new_n891));
  AOI21_X1  g690(.A(new_n343), .B1(new_n889), .B2(new_n891), .ZN(new_n892));
  OAI211_X1 g691(.A(new_n885), .B(new_n369), .C1(new_n852), .C2(new_n892), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n893), .A2(new_n857), .ZN(new_n894));
  NAND3_X1  g693(.A1(new_n283), .A2(new_n842), .A3(new_n886), .ZN(new_n895));
  AOI21_X1  g694(.A(new_n890), .B1(new_n895), .B2(new_n854), .ZN(new_n896));
  INV_X1    g695(.A(new_n891), .ZN(new_n897));
  OAI21_X1  g696(.A(new_n724), .B1(new_n896), .B2(new_n897), .ZN(new_n898));
  AND2_X1   g697(.A1(new_n849), .A2(new_n851), .ZN(new_n899));
  AOI21_X1  g698(.A(new_n835), .B1(new_n338), .B2(new_n342), .ZN(new_n900));
  NAND2_X1  g699(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  NAND2_X1  g700(.A1(new_n898), .A2(new_n901), .ZN(new_n902));
  AOI21_X1  g701(.A(new_n885), .B1(new_n902), .B2(new_n369), .ZN(new_n903));
  OAI211_X1 g702(.A(new_n882), .B(new_n884), .C1(new_n894), .C2(new_n903), .ZN(new_n904));
  NAND2_X1  g703(.A1(new_n853), .A2(new_n854), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n905), .A2(new_n724), .ZN(new_n906));
  AOI21_X1  g705(.A(new_n804), .B1(new_n906), .B2(new_n901), .ZN(new_n907));
  INV_X1    g706(.A(new_n857), .ZN(new_n908));
  OAI21_X1  g707(.A(new_n704), .B1(new_n907), .B2(new_n908), .ZN(new_n909));
  NAND2_X1  g708(.A1(new_n909), .A2(new_n883), .ZN(new_n910));
  NAND2_X1  g709(.A1(new_n904), .A2(new_n910), .ZN(new_n911));
  NAND2_X1  g710(.A1(new_n889), .A2(new_n891), .ZN(new_n912));
  AOI22_X1  g711(.A1(new_n912), .A2(new_n724), .B1(new_n899), .B2(new_n900), .ZN(new_n913));
  OAI21_X1  g712(.A(KEYINPUT118), .B1(new_n913), .B2(new_n804), .ZN(new_n914));
  NAND3_X1  g713(.A1(new_n914), .A2(new_n857), .A3(new_n893), .ZN(new_n915));
  AOI21_X1  g714(.A(new_n882), .B1(new_n915), .B2(new_n884), .ZN(new_n916));
  OAI211_X1 g715(.A(new_n745), .B(new_n881), .C1(new_n911), .C2(new_n916), .ZN(new_n917));
  NAND2_X1  g716(.A1(new_n917), .A2(G141gat), .ZN(new_n918));
  AOI21_X1  g717(.A(new_n624), .B1(new_n856), .B2(new_n857), .ZN(new_n919));
  NOR2_X1   g718(.A1(new_n712), .A2(G141gat), .ZN(new_n920));
  NAND3_X1  g719(.A1(new_n881), .A2(new_n919), .A3(new_n920), .ZN(new_n921));
  INV_X1    g720(.A(KEYINPUT120), .ZN(new_n922));
  NAND2_X1  g721(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  NAND4_X1  g722(.A1(new_n881), .A2(KEYINPUT120), .A3(new_n919), .A4(new_n920), .ZN(new_n924));
  NAND2_X1  g723(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  INV_X1    g724(.A(new_n925), .ZN(new_n926));
  NAND2_X1  g725(.A1(new_n918), .A2(new_n926), .ZN(new_n927));
  AOI21_X1  g726(.A(new_n880), .B1(new_n927), .B2(KEYINPUT58), .ZN(new_n928));
  AOI21_X1  g727(.A(new_n925), .B1(new_n917), .B2(G141gat), .ZN(new_n929));
  INV_X1    g728(.A(KEYINPUT58), .ZN(new_n930));
  NOR3_X1   g729(.A1(new_n929), .A2(KEYINPUT121), .A3(new_n930), .ZN(new_n931));
  NAND2_X1  g730(.A1(new_n921), .A2(new_n930), .ZN(new_n932));
  OAI211_X1 g731(.A(new_n283), .B(new_n881), .C1(new_n911), .C2(new_n916), .ZN(new_n933));
  AOI21_X1  g732(.A(new_n932), .B1(new_n933), .B2(G141gat), .ZN(new_n934));
  INV_X1    g733(.A(KEYINPUT122), .ZN(new_n935));
  NOR2_X1   g734(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  AOI211_X1 g735(.A(KEYINPUT122), .B(new_n932), .C1(new_n933), .C2(G141gat), .ZN(new_n937));
  OAI22_X1  g736(.A1(new_n928), .A2(new_n931), .B1(new_n936), .B2(new_n937), .ZN(G1344gat));
  INV_X1    g737(.A(new_n881), .ZN(new_n939));
  NOR2_X1   g738(.A1(new_n939), .A2(new_n909), .ZN(new_n940));
  INV_X1    g739(.A(G148gat), .ZN(new_n941));
  NAND3_X1  g740(.A1(new_n940), .A2(new_n941), .A3(new_n784), .ZN(new_n942));
  XOR2_X1   g741(.A(new_n942), .B(KEYINPUT123), .Z(new_n943));
  NOR2_X1   g742(.A1(new_n911), .A2(new_n916), .ZN(new_n944));
  NOR2_X1   g743(.A1(new_n944), .A2(new_n939), .ZN(new_n945));
  AOI211_X1 g744(.A(KEYINPUT59), .B(new_n941), .C1(new_n945), .C2(new_n784), .ZN(new_n946));
  INV_X1    g745(.A(KEYINPUT59), .ZN(new_n947));
  NAND2_X1  g746(.A1(new_n399), .A2(new_n712), .ZN(new_n948));
  NOR3_X1   g747(.A1(new_n724), .A2(new_n835), .A3(new_n848), .ZN(new_n949));
  OAI21_X1  g748(.A(new_n369), .B1(new_n949), .B2(new_n892), .ZN(new_n950));
  AOI211_X1 g749(.A(KEYINPUT57), .B(new_n624), .C1(new_n948), .C2(new_n950), .ZN(new_n951));
  AOI21_X1  g750(.A(new_n951), .B1(KEYINPUT57), .B2(new_n909), .ZN(new_n952));
  NAND3_X1  g751(.A1(new_n952), .A2(new_n784), .A3(new_n881), .ZN(new_n953));
  AOI21_X1  g752(.A(new_n947), .B1(new_n953), .B2(G148gat), .ZN(new_n954));
  OAI21_X1  g753(.A(new_n943), .B1(new_n946), .B2(new_n954), .ZN(G1345gat));
  NAND2_X1  g754(.A1(new_n945), .A2(new_n804), .ZN(new_n956));
  NAND2_X1  g755(.A1(new_n956), .A2(G155gat), .ZN(new_n957));
  INV_X1    g756(.A(KEYINPUT124), .ZN(new_n958));
  NOR4_X1   g757(.A1(new_n939), .A2(G155gat), .A3(new_n909), .A4(new_n369), .ZN(new_n959));
  INV_X1    g758(.A(new_n959), .ZN(new_n960));
  NAND3_X1  g759(.A1(new_n957), .A2(new_n958), .A3(new_n960), .ZN(new_n961));
  AOI21_X1  g760(.A(new_n365), .B1(new_n945), .B2(new_n804), .ZN(new_n962));
  OAI21_X1  g761(.A(KEYINPUT124), .B1(new_n962), .B2(new_n959), .ZN(new_n963));
  NAND2_X1  g762(.A1(new_n961), .A2(new_n963), .ZN(G1346gat));
  AOI21_X1  g763(.A(G162gat), .B1(new_n940), .B2(new_n343), .ZN(new_n965));
  NOR2_X1   g764(.A1(new_n724), .A2(new_n557), .ZN(new_n966));
  AOI21_X1  g765(.A(new_n965), .B1(new_n945), .B2(new_n966), .ZN(G1347gat));
  NOR2_X1   g766(.A1(new_n667), .A2(new_n596), .ZN(new_n968));
  NAND2_X1  g767(.A1(new_n864), .A2(new_n968), .ZN(new_n969));
  OR2_X1    g768(.A1(new_n969), .A2(KEYINPUT126), .ZN(new_n970));
  NAND2_X1  g769(.A1(new_n969), .A2(KEYINPUT126), .ZN(new_n971));
  NAND2_X1  g770(.A1(new_n970), .A2(new_n971), .ZN(new_n972));
  OAI21_X1  g771(.A(G169gat), .B1(new_n972), .B2(new_n712), .ZN(new_n973));
  INV_X1    g772(.A(new_n968), .ZN(new_n974));
  NOR3_X1   g773(.A1(new_n974), .A2(new_n859), .A3(new_n704), .ZN(new_n975));
  NAND2_X1  g774(.A1(new_n858), .A2(new_n975), .ZN(new_n976));
  INV_X1    g775(.A(new_n976), .ZN(new_n977));
  NAND3_X1  g776(.A1(new_n977), .A2(new_n452), .A3(new_n745), .ZN(new_n978));
  XNOR2_X1  g777(.A(new_n978), .B(KEYINPUT125), .ZN(new_n979));
  NAND2_X1  g778(.A1(new_n973), .A2(new_n979), .ZN(G1348gat));
  OAI21_X1  g779(.A(G176gat), .B1(new_n972), .B2(new_n397), .ZN(new_n981));
  NAND3_X1  g780(.A1(new_n977), .A2(new_n453), .A3(new_n784), .ZN(new_n982));
  NAND2_X1  g781(.A1(new_n981), .A2(new_n982), .ZN(G1349gat));
  OAI21_X1  g782(.A(G183gat), .B1(new_n972), .B2(new_n369), .ZN(new_n984));
  NAND3_X1  g783(.A1(new_n977), .A2(new_n466), .A3(new_n804), .ZN(new_n985));
  NAND2_X1  g784(.A1(new_n984), .A2(new_n985), .ZN(new_n986));
  NAND2_X1  g785(.A1(new_n986), .A2(KEYINPUT60), .ZN(new_n987));
  INV_X1    g786(.A(KEYINPUT60), .ZN(new_n988));
  NAND3_X1  g787(.A1(new_n984), .A2(new_n988), .A3(new_n985), .ZN(new_n989));
  NAND2_X1  g788(.A1(new_n987), .A2(new_n989), .ZN(G1350gat));
  NAND3_X1  g789(.A1(new_n977), .A2(new_n289), .A3(new_n343), .ZN(new_n991));
  NAND3_X1  g790(.A1(new_n970), .A2(new_n343), .A3(new_n971), .ZN(new_n992));
  INV_X1    g791(.A(KEYINPUT61), .ZN(new_n993));
  AND3_X1   g792(.A1(new_n992), .A2(new_n993), .A3(G190gat), .ZN(new_n994));
  AOI21_X1  g793(.A(new_n993), .B1(new_n992), .B2(G190gat), .ZN(new_n995));
  OAI21_X1  g794(.A(new_n991), .B1(new_n994), .B2(new_n995), .ZN(G1351gat));
  NOR2_X1   g795(.A1(new_n699), .A2(new_n974), .ZN(new_n997));
  XOR2_X1   g796(.A(new_n997), .B(KEYINPUT127), .Z(new_n998));
  NAND2_X1  g797(.A1(new_n998), .A2(new_n952), .ZN(new_n999));
  INV_X1    g798(.A(G197gat), .ZN(new_n1000));
  NOR3_X1   g799(.A1(new_n999), .A2(new_n1000), .A3(new_n712), .ZN(new_n1001));
  NAND2_X1  g800(.A1(new_n997), .A2(new_n919), .ZN(new_n1002));
  INV_X1    g801(.A(new_n1002), .ZN(new_n1003));
  AOI21_X1  g802(.A(G197gat), .B1(new_n1003), .B2(new_n745), .ZN(new_n1004));
  NOR2_X1   g803(.A1(new_n1001), .A2(new_n1004), .ZN(G1352gat));
  NAND3_X1  g804(.A1(new_n998), .A2(new_n784), .A3(new_n952), .ZN(new_n1006));
  NAND2_X1  g805(.A1(new_n1006), .A2(G204gat), .ZN(new_n1007));
  NOR3_X1   g806(.A1(new_n1002), .A2(G204gat), .A3(new_n397), .ZN(new_n1008));
  INV_X1    g807(.A(KEYINPUT62), .ZN(new_n1009));
  OR2_X1    g808(.A1(new_n1008), .A2(new_n1009), .ZN(new_n1010));
  NAND2_X1  g809(.A1(new_n1008), .A2(new_n1009), .ZN(new_n1011));
  NAND3_X1  g810(.A1(new_n1007), .A2(new_n1010), .A3(new_n1011), .ZN(G1353gat));
  NAND3_X1  g811(.A1(new_n1003), .A2(new_n523), .A3(new_n804), .ZN(new_n1013));
  NAND3_X1  g812(.A1(new_n998), .A2(new_n804), .A3(new_n952), .ZN(new_n1014));
  AND3_X1   g813(.A1(new_n1014), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n1015));
  AOI21_X1  g814(.A(KEYINPUT63), .B1(new_n1014), .B2(G211gat), .ZN(new_n1016));
  OAI21_X1  g815(.A(new_n1013), .B1(new_n1015), .B2(new_n1016), .ZN(G1354gat));
  OAI21_X1  g816(.A(G218gat), .B1(new_n999), .B2(new_n724), .ZN(new_n1018));
  NAND3_X1  g817(.A1(new_n1003), .A2(new_n340), .A3(new_n343), .ZN(new_n1019));
  NAND2_X1  g818(.A1(new_n1018), .A2(new_n1019), .ZN(G1355gat));
endmodule


