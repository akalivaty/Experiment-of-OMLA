//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 0 1 1 1 1 0 0 0 0 1 0 0 0 1 0 0 1 0 0 0 0 1 1 0 1 0 0 1 0 0 1 1 0 0 1 1 0 0 1 0 1 0 1 0 1 1 1 1 1 1 1 1 0 1 0 1 1 0 0 1 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:26:23 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n680, new_n681, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n716, new_n717, new_n718, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n741, new_n742, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n751, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n774, new_n775, new_n776, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n802, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n825, new_n826, new_n827, new_n828, new_n829, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n947, new_n948, new_n949, new_n950, new_n951, new_n952,
    new_n953, new_n954, new_n955, new_n956, new_n957, new_n958, new_n959,
    new_n960, new_n961, new_n962, new_n963, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n972, new_n973, new_n974, new_n975,
    new_n977, new_n978, new_n979, new_n980, new_n981, new_n982, new_n983,
    new_n984, new_n985, new_n986, new_n987, new_n988, new_n989, new_n990,
    new_n992, new_n993, new_n994, new_n995, new_n996, new_n997, new_n998,
    new_n999, new_n1000, new_n1001, new_n1002, new_n1003, new_n1004,
    new_n1005, new_n1006, new_n1007, new_n1008, new_n1009, new_n1010,
    new_n1012, new_n1013, new_n1014, new_n1015, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1022, new_n1023, new_n1024,
    new_n1025, new_n1026, new_n1027, new_n1028, new_n1029, new_n1030,
    new_n1031, new_n1032, new_n1033, new_n1034, new_n1035, new_n1036,
    new_n1037, new_n1039, new_n1040, new_n1041, new_n1042, new_n1043,
    new_n1044, new_n1045, new_n1046, new_n1047, new_n1048, new_n1049,
    new_n1050, new_n1051;
  INV_X1    g000(.A(G146), .ZN(new_n187));
  NOR2_X1   g001(.A1(new_n187), .A2(G143), .ZN(new_n188));
  INV_X1    g002(.A(new_n188), .ZN(new_n189));
  XNOR2_X1  g003(.A(KEYINPUT64), .B(G143), .ZN(new_n190));
  OAI21_X1  g004(.A(new_n189), .B1(new_n190), .B2(G146), .ZN(new_n191));
  AND2_X1   g005(.A1(KEYINPUT0), .A2(G128), .ZN(new_n192));
  NOR2_X1   g006(.A1(KEYINPUT0), .A2(G128), .ZN(new_n193));
  NOR2_X1   g007(.A1(new_n192), .A2(new_n193), .ZN(new_n194));
  INV_X1    g008(.A(G143), .ZN(new_n195));
  NOR2_X1   g009(.A1(new_n195), .A2(G146), .ZN(new_n196));
  AOI21_X1  g010(.A(new_n196), .B1(new_n190), .B2(G146), .ZN(new_n197));
  AOI22_X1  g011(.A1(new_n191), .A2(new_n194), .B1(new_n197), .B2(new_n192), .ZN(new_n198));
  INV_X1    g012(.A(G104), .ZN(new_n199));
  OAI21_X1  g013(.A(KEYINPUT3), .B1(new_n199), .B2(G107), .ZN(new_n200));
  INV_X1    g014(.A(KEYINPUT3), .ZN(new_n201));
  INV_X1    g015(.A(G107), .ZN(new_n202));
  NAND3_X1  g016(.A1(new_n201), .A2(new_n202), .A3(G104), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n199), .A2(G107), .ZN(new_n204));
  NAND3_X1  g018(.A1(new_n200), .A2(new_n203), .A3(new_n204), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n205), .A2(G101), .ZN(new_n206));
  INV_X1    g020(.A(G101), .ZN(new_n207));
  NAND4_X1  g021(.A1(new_n200), .A2(new_n203), .A3(new_n207), .A4(new_n204), .ZN(new_n208));
  NAND3_X1  g022(.A1(new_n206), .A2(KEYINPUT4), .A3(new_n208), .ZN(new_n209));
  INV_X1    g023(.A(KEYINPUT4), .ZN(new_n210));
  NAND3_X1  g024(.A1(new_n205), .A2(new_n210), .A3(G101), .ZN(new_n211));
  AND3_X1   g025(.A1(new_n198), .A2(new_n209), .A3(new_n211), .ZN(new_n212));
  INV_X1    g026(.A(KEYINPUT1), .ZN(new_n213));
  OAI21_X1  g027(.A(G128), .B1(new_n196), .B2(new_n213), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n195), .A2(KEYINPUT64), .ZN(new_n215));
  INV_X1    g029(.A(KEYINPUT64), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n216), .A2(G143), .ZN(new_n217));
  AOI21_X1  g031(.A(G146), .B1(new_n215), .B2(new_n217), .ZN(new_n218));
  OAI21_X1  g032(.A(new_n214), .B1(new_n218), .B2(new_n188), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n219), .A2(KEYINPUT66), .ZN(new_n220));
  INV_X1    g034(.A(KEYINPUT66), .ZN(new_n221));
  NAND3_X1  g035(.A1(new_n191), .A2(new_n221), .A3(new_n214), .ZN(new_n222));
  INV_X1    g036(.A(G128), .ZN(new_n223));
  NOR2_X1   g037(.A1(new_n223), .A2(KEYINPUT1), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n197), .A2(new_n224), .ZN(new_n225));
  NAND3_X1  g039(.A1(new_n220), .A2(new_n222), .A3(new_n225), .ZN(new_n226));
  NOR2_X1   g040(.A1(new_n199), .A2(G107), .ZN(new_n227));
  NOR2_X1   g041(.A1(new_n202), .A2(G104), .ZN(new_n228));
  OAI21_X1  g042(.A(G101), .B1(new_n227), .B2(new_n228), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n208), .A2(new_n229), .ZN(new_n230));
  INV_X1    g044(.A(KEYINPUT10), .ZN(new_n231));
  NOR2_X1   g045(.A1(new_n230), .A2(new_n231), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n226), .A2(new_n232), .ZN(new_n233));
  INV_X1    g047(.A(KEYINPUT76), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n233), .A2(new_n234), .ZN(new_n235));
  NAND3_X1  g049(.A1(new_n226), .A2(KEYINPUT76), .A3(new_n232), .ZN(new_n236));
  AOI21_X1  g050(.A(new_n212), .B1(new_n235), .B2(new_n236), .ZN(new_n237));
  INV_X1    g051(.A(KEYINPUT75), .ZN(new_n238));
  NOR2_X1   g052(.A1(new_n216), .A2(G143), .ZN(new_n239));
  NOR2_X1   g053(.A1(new_n195), .A2(KEYINPUT64), .ZN(new_n240));
  OAI21_X1  g054(.A(new_n187), .B1(new_n239), .B2(new_n240), .ZN(new_n241));
  AOI21_X1  g055(.A(new_n223), .B1(new_n241), .B2(KEYINPUT1), .ZN(new_n242));
  OAI21_X1  g056(.A(KEYINPUT74), .B1(new_n242), .B2(new_n197), .ZN(new_n243));
  INV_X1    g057(.A(KEYINPUT74), .ZN(new_n244));
  INV_X1    g058(.A(new_n196), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n215), .A2(new_n217), .ZN(new_n246));
  OAI21_X1  g060(.A(new_n245), .B1(new_n246), .B2(new_n187), .ZN(new_n247));
  AOI21_X1  g061(.A(new_n213), .B1(new_n246), .B2(new_n187), .ZN(new_n248));
  OAI211_X1 g062(.A(new_n244), .B(new_n247), .C1(new_n248), .C2(new_n223), .ZN(new_n249));
  NAND3_X1  g063(.A1(new_n243), .A2(new_n225), .A3(new_n249), .ZN(new_n250));
  INV_X1    g064(.A(new_n230), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n250), .A2(new_n251), .ZN(new_n252));
  AOI21_X1  g066(.A(new_n238), .B1(new_n252), .B2(new_n231), .ZN(new_n253));
  AOI211_X1 g067(.A(KEYINPUT75), .B(KEYINPUT10), .C1(new_n250), .C2(new_n251), .ZN(new_n254));
  OAI21_X1  g068(.A(new_n237), .B1(new_n253), .B2(new_n254), .ZN(new_n255));
  INV_X1    g069(.A(G137), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n256), .A2(G134), .ZN(new_n257));
  INV_X1    g071(.A(G134), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n258), .A2(G137), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n257), .A2(new_n259), .ZN(new_n260));
  NOR2_X1   g074(.A1(KEYINPUT65), .A2(KEYINPUT11), .ZN(new_n261));
  INV_X1    g075(.A(new_n261), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n260), .A2(new_n262), .ZN(new_n263));
  NAND2_X1  g077(.A1(KEYINPUT65), .A2(KEYINPUT11), .ZN(new_n264));
  INV_X1    g078(.A(new_n264), .ZN(new_n265));
  OAI21_X1  g079(.A(new_n257), .B1(new_n265), .B2(new_n261), .ZN(new_n266));
  INV_X1    g080(.A(G131), .ZN(new_n267));
  NAND3_X1  g081(.A1(new_n263), .A2(new_n266), .A3(new_n267), .ZN(new_n268));
  INV_X1    g082(.A(new_n268), .ZN(new_n269));
  AOI21_X1  g083(.A(new_n267), .B1(new_n263), .B2(new_n266), .ZN(new_n270));
  NOR2_X1   g084(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  INV_X1    g085(.A(new_n271), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n255), .A2(new_n272), .ZN(new_n273));
  INV_X1    g087(.A(KEYINPUT78), .ZN(new_n274));
  OAI211_X1 g088(.A(new_n237), .B(new_n271), .C1(new_n253), .C2(new_n254), .ZN(new_n275));
  NAND3_X1  g089(.A1(new_n273), .A2(new_n274), .A3(new_n275), .ZN(new_n276));
  INV_X1    g090(.A(G953), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n277), .A2(G227), .ZN(new_n278));
  XNOR2_X1  g092(.A(new_n278), .B(G140), .ZN(new_n279));
  XNOR2_X1  g093(.A(KEYINPUT73), .B(G110), .ZN(new_n280));
  XNOR2_X1  g094(.A(new_n279), .B(new_n280), .ZN(new_n281));
  NAND3_X1  g095(.A1(new_n255), .A2(KEYINPUT78), .A3(new_n272), .ZN(new_n282));
  NAND3_X1  g096(.A1(new_n276), .A2(new_n281), .A3(new_n282), .ZN(new_n283));
  INV_X1    g097(.A(KEYINPUT12), .ZN(new_n284));
  AOI21_X1  g098(.A(new_n271), .B1(KEYINPUT77), .B2(new_n284), .ZN(new_n285));
  OAI21_X1  g099(.A(new_n247), .B1(new_n248), .B2(new_n223), .ZN(new_n286));
  AOI22_X1  g100(.A1(new_n286), .A2(KEYINPUT74), .B1(new_n197), .B2(new_n224), .ZN(new_n287));
  AOI21_X1  g101(.A(new_n230), .B1(new_n287), .B2(new_n249), .ZN(new_n288));
  NOR2_X1   g102(.A1(new_n226), .A2(new_n251), .ZN(new_n289));
  OAI21_X1  g103(.A(new_n285), .B1(new_n288), .B2(new_n289), .ZN(new_n290));
  INV_X1    g104(.A(KEYINPUT77), .ZN(new_n291));
  NAND3_X1  g105(.A1(new_n290), .A2(new_n291), .A3(KEYINPUT12), .ZN(new_n292));
  OAI221_X1 g106(.A(new_n285), .B1(KEYINPUT77), .B2(new_n284), .C1(new_n288), .C2(new_n289), .ZN(new_n293));
  NAND3_X1  g107(.A1(new_n275), .A2(new_n292), .A3(new_n293), .ZN(new_n294));
  OR2_X1    g108(.A1(new_n294), .A2(new_n281), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n283), .A2(new_n295), .ZN(new_n296));
  INV_X1    g110(.A(G469), .ZN(new_n297));
  INV_X1    g111(.A(G902), .ZN(new_n298));
  NAND3_X1  g112(.A1(new_n296), .A2(new_n297), .A3(new_n298), .ZN(new_n299));
  NOR2_X1   g113(.A1(new_n297), .A2(new_n298), .ZN(new_n300));
  INV_X1    g114(.A(new_n300), .ZN(new_n301));
  INV_X1    g115(.A(new_n281), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n275), .A2(new_n274), .ZN(new_n303));
  OAI21_X1  g117(.A(KEYINPUT75), .B1(new_n288), .B2(KEYINPUT10), .ZN(new_n304));
  NAND3_X1  g118(.A1(new_n252), .A2(new_n238), .A3(new_n231), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  AOI21_X1  g120(.A(new_n271), .B1(new_n306), .B2(new_n237), .ZN(new_n307));
  NOR2_X1   g121(.A1(new_n303), .A2(new_n307), .ZN(new_n308));
  INV_X1    g122(.A(new_n282), .ZN(new_n309));
  OAI21_X1  g123(.A(new_n302), .B1(new_n308), .B2(new_n309), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n294), .A2(new_n281), .ZN(new_n311));
  NAND3_X1  g125(.A1(new_n310), .A2(G469), .A3(new_n311), .ZN(new_n312));
  NAND3_X1  g126(.A1(new_n299), .A2(new_n301), .A3(new_n312), .ZN(new_n313));
  XNOR2_X1  g127(.A(KEYINPUT9), .B(G234), .ZN(new_n314));
  INV_X1    g128(.A(G217), .ZN(new_n315));
  NOR3_X1   g129(.A1(new_n314), .A2(new_n315), .A3(G953), .ZN(new_n316));
  INV_X1    g130(.A(new_n316), .ZN(new_n317));
  NAND3_X1  g131(.A1(new_n215), .A2(new_n217), .A3(G128), .ZN(new_n318));
  INV_X1    g132(.A(KEYINPUT91), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n318), .A2(new_n319), .ZN(new_n320));
  NAND3_X1  g134(.A1(new_n190), .A2(KEYINPUT91), .A3(G128), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n320), .A2(new_n321), .ZN(new_n322));
  INV_X1    g136(.A(KEYINPUT13), .ZN(new_n323));
  NOR2_X1   g137(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  NOR2_X1   g138(.A1(new_n195), .A2(G128), .ZN(new_n325));
  AOI21_X1  g139(.A(new_n325), .B1(new_n322), .B2(new_n323), .ZN(new_n326));
  AOI21_X1  g140(.A(new_n324), .B1(new_n326), .B2(KEYINPUT92), .ZN(new_n327));
  INV_X1    g141(.A(KEYINPUT92), .ZN(new_n328));
  AOI21_X1  g142(.A(KEYINPUT13), .B1(new_n320), .B2(new_n321), .ZN(new_n329));
  OAI21_X1  g143(.A(new_n328), .B1(new_n329), .B2(new_n325), .ZN(new_n330));
  AOI21_X1  g144(.A(new_n258), .B1(new_n327), .B2(new_n330), .ZN(new_n331));
  INV_X1    g145(.A(new_n325), .ZN(new_n332));
  AOI21_X1  g146(.A(KEYINPUT93), .B1(new_n322), .B2(new_n332), .ZN(new_n333));
  INV_X1    g147(.A(KEYINPUT93), .ZN(new_n334));
  AOI211_X1 g148(.A(new_n334), .B(new_n325), .C1(new_n320), .C2(new_n321), .ZN(new_n335));
  OAI21_X1  g149(.A(new_n258), .B1(new_n333), .B2(new_n335), .ZN(new_n336));
  INV_X1    g150(.A(KEYINPUT89), .ZN(new_n337));
  INV_X1    g151(.A(G116), .ZN(new_n338));
  OAI21_X1  g152(.A(new_n337), .B1(new_n338), .B2(G122), .ZN(new_n339));
  INV_X1    g153(.A(G122), .ZN(new_n340));
  NAND3_X1  g154(.A1(new_n340), .A2(KEYINPUT89), .A3(G116), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n339), .A2(new_n341), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n338), .A2(G122), .ZN(new_n343));
  NAND3_X1  g157(.A1(new_n342), .A2(KEYINPUT90), .A3(new_n343), .ZN(new_n344));
  INV_X1    g158(.A(new_n344), .ZN(new_n345));
  AOI21_X1  g159(.A(KEYINPUT90), .B1(new_n342), .B2(new_n343), .ZN(new_n346));
  OAI21_X1  g160(.A(new_n202), .B1(new_n345), .B2(new_n346), .ZN(new_n347));
  INV_X1    g161(.A(new_n346), .ZN(new_n348));
  NAND3_X1  g162(.A1(new_n348), .A2(G107), .A3(new_n344), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n347), .A2(new_n349), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n336), .A2(new_n350), .ZN(new_n351));
  NOR2_X1   g165(.A1(new_n331), .A2(new_n351), .ZN(new_n352));
  XOR2_X1   g166(.A(new_n343), .B(KEYINPUT14), .Z(new_n353));
  NAND2_X1  g167(.A1(new_n353), .A2(new_n342), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n354), .A2(G107), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n355), .A2(new_n347), .ZN(new_n356));
  AOI21_X1  g170(.A(KEYINPUT91), .B1(new_n190), .B2(G128), .ZN(new_n357));
  AND4_X1   g171(.A1(KEYINPUT91), .A2(new_n215), .A3(new_n217), .A4(G128), .ZN(new_n358));
  OAI21_X1  g172(.A(new_n332), .B1(new_n357), .B2(new_n358), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n359), .A2(new_n334), .ZN(new_n360));
  NAND3_X1  g174(.A1(new_n322), .A2(KEYINPUT93), .A3(new_n332), .ZN(new_n361));
  NAND3_X1  g175(.A1(new_n360), .A2(G134), .A3(new_n361), .ZN(new_n362));
  AOI21_X1  g176(.A(new_n356), .B1(new_n336), .B2(new_n362), .ZN(new_n363));
  OAI21_X1  g177(.A(KEYINPUT94), .B1(new_n352), .B2(new_n363), .ZN(new_n364));
  INV_X1    g178(.A(new_n324), .ZN(new_n365));
  OAI21_X1  g179(.A(new_n323), .B1(new_n357), .B2(new_n358), .ZN(new_n366));
  NAND3_X1  g180(.A1(new_n366), .A2(KEYINPUT92), .A3(new_n332), .ZN(new_n367));
  NAND3_X1  g181(.A1(new_n330), .A2(new_n365), .A3(new_n367), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n368), .A2(G134), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n360), .A2(new_n361), .ZN(new_n370));
  AOI22_X1  g184(.A1(new_n370), .A2(new_n258), .B1(new_n349), .B2(new_n347), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n369), .A2(new_n371), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n336), .A2(new_n362), .ZN(new_n373));
  INV_X1    g187(.A(new_n356), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n373), .A2(new_n374), .ZN(new_n375));
  INV_X1    g189(.A(KEYINPUT94), .ZN(new_n376));
  NAND3_X1  g190(.A1(new_n372), .A2(new_n375), .A3(new_n376), .ZN(new_n377));
  AOI21_X1  g191(.A(new_n317), .B1(new_n364), .B2(new_n377), .ZN(new_n378));
  AOI21_X1  g192(.A(new_n363), .B1(new_n369), .B2(new_n371), .ZN(new_n379));
  AOI21_X1  g193(.A(new_n316), .B1(new_n379), .B2(new_n376), .ZN(new_n380));
  OAI21_X1  g194(.A(new_n298), .B1(new_n378), .B2(new_n380), .ZN(new_n381));
  INV_X1    g195(.A(G478), .ZN(new_n382));
  NOR2_X1   g196(.A1(new_n382), .A2(KEYINPUT15), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n381), .A2(new_n383), .ZN(new_n384));
  INV_X1    g198(.A(KEYINPUT87), .ZN(new_n385));
  XNOR2_X1  g199(.A(G113), .B(G122), .ZN(new_n386));
  XNOR2_X1  g200(.A(new_n386), .B(G104), .ZN(new_n387));
  INV_X1    g201(.A(KEYINPUT16), .ZN(new_n388));
  INV_X1    g202(.A(G140), .ZN(new_n389));
  NAND3_X1  g203(.A1(new_n388), .A2(new_n389), .A3(G125), .ZN(new_n390));
  INV_X1    g204(.A(G125), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n391), .A2(G140), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n389), .A2(G125), .ZN(new_n393));
  INV_X1    g207(.A(KEYINPUT71), .ZN(new_n394));
  NAND3_X1  g208(.A1(new_n392), .A2(new_n393), .A3(new_n394), .ZN(new_n395));
  NAND3_X1  g209(.A1(new_n391), .A2(KEYINPUT71), .A3(G140), .ZN(new_n396));
  AOI21_X1  g210(.A(new_n388), .B1(new_n395), .B2(new_n396), .ZN(new_n397));
  INV_X1    g211(.A(KEYINPUT72), .ZN(new_n398));
  OAI21_X1  g212(.A(new_n390), .B1(new_n397), .B2(new_n398), .ZN(new_n399));
  AOI211_X1 g213(.A(KEYINPUT72), .B(new_n388), .C1(new_n395), .C2(new_n396), .ZN(new_n400));
  OAI21_X1  g214(.A(new_n187), .B1(new_n399), .B2(new_n400), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n395), .A2(new_n396), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n402), .A2(KEYINPUT16), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n403), .A2(KEYINPUT72), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n397), .A2(new_n398), .ZN(new_n405));
  NAND4_X1  g219(.A1(new_n404), .A2(G146), .A3(new_n405), .A4(new_n390), .ZN(new_n406));
  INV_X1    g220(.A(G214), .ZN(new_n407));
  NOR3_X1   g221(.A1(new_n407), .A2(G237), .A3(G953), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n408), .A2(G143), .ZN(new_n409));
  OAI21_X1  g223(.A(new_n409), .B1(new_n246), .B2(new_n408), .ZN(new_n410));
  NAND3_X1  g224(.A1(new_n410), .A2(KEYINPUT17), .A3(G131), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n410), .A2(G131), .ZN(new_n412));
  INV_X1    g226(.A(KEYINPUT17), .ZN(new_n413));
  OAI211_X1 g227(.A(new_n409), .B(new_n267), .C1(new_n246), .C2(new_n408), .ZN(new_n414));
  NAND3_X1  g228(.A1(new_n412), .A2(new_n413), .A3(new_n414), .ZN(new_n415));
  NAND4_X1  g229(.A1(new_n401), .A2(new_n406), .A3(new_n411), .A4(new_n415), .ZN(new_n416));
  OAI21_X1  g230(.A(KEYINPUT85), .B1(new_n402), .B2(new_n187), .ZN(new_n417));
  AND2_X1   g231(.A1(new_n392), .A2(new_n393), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n418), .A2(new_n187), .ZN(new_n419));
  INV_X1    g233(.A(KEYINPUT85), .ZN(new_n420));
  NAND4_X1  g234(.A1(new_n395), .A2(new_n420), .A3(G146), .A4(new_n396), .ZN(new_n421));
  NAND3_X1  g235(.A1(new_n417), .A2(new_n419), .A3(new_n421), .ZN(new_n422));
  AND2_X1   g236(.A1(KEYINPUT18), .A2(G131), .ZN(new_n423));
  INV_X1    g237(.A(new_n423), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n410), .A2(new_n424), .ZN(new_n425));
  OAI211_X1 g239(.A(new_n409), .B(new_n423), .C1(new_n246), .C2(new_n408), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n425), .A2(new_n426), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n422), .A2(new_n427), .ZN(new_n428));
  AOI21_X1  g242(.A(new_n387), .B1(new_n416), .B2(new_n428), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n428), .A2(new_n387), .ZN(new_n430));
  NOR2_X1   g244(.A1(new_n399), .A2(new_n400), .ZN(new_n431));
  AOI22_X1  g245(.A1(new_n431), .A2(G146), .B1(new_n412), .B2(new_n414), .ZN(new_n432));
  INV_X1    g246(.A(KEYINPUT86), .ZN(new_n433));
  NOR2_X1   g247(.A1(new_n418), .A2(KEYINPUT19), .ZN(new_n434));
  AOI21_X1  g248(.A(new_n434), .B1(new_n402), .B2(KEYINPUT19), .ZN(new_n435));
  OAI21_X1  g249(.A(new_n433), .B1(new_n435), .B2(G146), .ZN(new_n436));
  AND2_X1   g250(.A1(new_n402), .A2(KEYINPUT19), .ZN(new_n437));
  OAI211_X1 g251(.A(KEYINPUT86), .B(new_n187), .C1(new_n437), .C2(new_n434), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n436), .A2(new_n438), .ZN(new_n439));
  AOI21_X1  g253(.A(new_n430), .B1(new_n432), .B2(new_n439), .ZN(new_n440));
  NOR2_X1   g254(.A1(G475), .A2(G902), .ZN(new_n441));
  INV_X1    g255(.A(new_n441), .ZN(new_n442));
  NOR3_X1   g256(.A1(new_n429), .A2(new_n440), .A3(new_n442), .ZN(new_n443));
  INV_X1    g257(.A(KEYINPUT20), .ZN(new_n444));
  OAI21_X1  g258(.A(new_n385), .B1(new_n443), .B2(new_n444), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n416), .A2(new_n428), .ZN(new_n446));
  INV_X1    g260(.A(new_n387), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n446), .A2(new_n447), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n432), .A2(new_n439), .ZN(new_n449));
  NAND3_X1  g263(.A1(new_n449), .A2(new_n387), .A3(new_n428), .ZN(new_n450));
  NAND3_X1  g264(.A1(new_n448), .A2(new_n450), .A3(new_n441), .ZN(new_n451));
  NAND3_X1  g265(.A1(new_n451), .A2(KEYINPUT87), .A3(KEYINPUT20), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n443), .A2(new_n444), .ZN(new_n453));
  NAND3_X1  g267(.A1(new_n445), .A2(new_n452), .A3(new_n453), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n387), .A2(KEYINPUT88), .ZN(new_n455));
  AOI21_X1  g269(.A(G902), .B1(new_n446), .B2(new_n455), .ZN(new_n456));
  OAI21_X1  g270(.A(new_n456), .B1(new_n446), .B2(new_n455), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n457), .A2(G475), .ZN(new_n458));
  INV_X1    g272(.A(new_n383), .ZN(new_n459));
  OAI211_X1 g273(.A(new_n298), .B(new_n459), .C1(new_n378), .C2(new_n380), .ZN(new_n460));
  NAND4_X1  g274(.A1(new_n384), .A2(new_n454), .A3(new_n458), .A4(new_n460), .ZN(new_n461));
  OAI21_X1  g275(.A(G210), .B1(G237), .B2(G902), .ZN(new_n462));
  INV_X1    g276(.A(new_n462), .ZN(new_n463));
  INV_X1    g277(.A(G119), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n338), .A2(new_n464), .ZN(new_n465));
  NAND2_X1  g279(.A1(G116), .A2(G119), .ZN(new_n466));
  AND2_X1   g280(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  OR2_X1    g281(.A1(KEYINPUT2), .A2(G113), .ZN(new_n468));
  NAND2_X1  g282(.A1(KEYINPUT2), .A2(G113), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n467), .A2(new_n470), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n465), .A2(new_n466), .ZN(new_n472));
  NAND3_X1  g286(.A1(new_n472), .A2(new_n468), .A3(new_n469), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n471), .A2(new_n473), .ZN(new_n474));
  INV_X1    g288(.A(KEYINPUT67), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  NAND3_X1  g290(.A1(new_n471), .A2(new_n473), .A3(KEYINPUT67), .ZN(new_n477));
  NAND4_X1  g291(.A1(new_n476), .A2(new_n477), .A3(new_n211), .A4(new_n209), .ZN(new_n478));
  INV_X1    g292(.A(G113), .ZN(new_n479));
  XNOR2_X1  g293(.A(KEYINPUT80), .B(KEYINPUT5), .ZN(new_n480));
  NOR2_X1   g294(.A1(new_n338), .A2(G119), .ZN(new_n481));
  AOI21_X1  g295(.A(new_n479), .B1(new_n480), .B2(new_n481), .ZN(new_n482));
  OAI21_X1  g296(.A(new_n482), .B1(new_n467), .B2(new_n480), .ZN(new_n483));
  NAND3_X1  g297(.A1(new_n483), .A2(new_n251), .A3(new_n473), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n478), .A2(new_n484), .ZN(new_n485));
  XNOR2_X1  g299(.A(G110), .B(G122), .ZN(new_n486));
  INV_X1    g300(.A(new_n486), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n485), .A2(new_n487), .ZN(new_n488));
  NAND3_X1  g302(.A1(new_n478), .A2(new_n486), .A3(new_n484), .ZN(new_n489));
  NAND3_X1  g303(.A1(new_n488), .A2(KEYINPUT6), .A3(new_n489), .ZN(new_n490));
  NAND4_X1  g304(.A1(new_n220), .A2(new_n391), .A3(new_n222), .A4(new_n225), .ZN(new_n491));
  OAI211_X1 g305(.A(new_n245), .B(new_n192), .C1(new_n246), .C2(new_n187), .ZN(new_n492));
  NOR2_X1   g306(.A1(new_n218), .A2(new_n188), .ZN(new_n493));
  INV_X1    g307(.A(new_n194), .ZN(new_n494));
  OAI21_X1  g308(.A(new_n492), .B1(new_n493), .B2(new_n494), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n495), .A2(G125), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n491), .A2(new_n496), .ZN(new_n497));
  INV_X1    g311(.A(G224), .ZN(new_n498));
  NOR2_X1   g312(.A1(new_n498), .A2(G953), .ZN(new_n499));
  XNOR2_X1  g313(.A(new_n499), .B(KEYINPUT81), .ZN(new_n500));
  XOR2_X1   g314(.A(new_n500), .B(KEYINPUT82), .Z(new_n501));
  XNOR2_X1  g315(.A(new_n497), .B(new_n501), .ZN(new_n502));
  INV_X1    g316(.A(KEYINPUT6), .ZN(new_n503));
  NAND3_X1  g317(.A1(new_n485), .A2(new_n503), .A3(new_n487), .ZN(new_n504));
  AND3_X1   g318(.A1(new_n490), .A2(new_n502), .A3(new_n504), .ZN(new_n505));
  XNOR2_X1  g319(.A(new_n486), .B(KEYINPUT8), .ZN(new_n506));
  INV_X1    g320(.A(KEYINPUT5), .ZN(new_n507));
  OAI21_X1  g321(.A(new_n482), .B1(new_n507), .B2(new_n467), .ZN(new_n508));
  NAND3_X1  g322(.A1(new_n508), .A2(new_n251), .A3(new_n473), .ZN(new_n509));
  AOI21_X1  g323(.A(new_n251), .B1(new_n483), .B2(new_n473), .ZN(new_n510));
  INV_X1    g324(.A(KEYINPUT83), .ZN(new_n511));
  OAI21_X1  g325(.A(new_n509), .B1(new_n510), .B2(new_n511), .ZN(new_n512));
  AOI211_X1 g326(.A(KEYINPUT83), .B(new_n251), .C1(new_n473), .C2(new_n483), .ZN(new_n513));
  OAI21_X1  g327(.A(new_n506), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  OAI21_X1  g328(.A(KEYINPUT7), .B1(new_n498), .B2(G953), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n497), .A2(new_n515), .ZN(new_n516));
  INV_X1    g330(.A(new_n515), .ZN(new_n517));
  NAND3_X1  g331(.A1(new_n491), .A2(new_n496), .A3(new_n517), .ZN(new_n518));
  NAND4_X1  g332(.A1(new_n514), .A2(new_n489), .A3(new_n516), .A4(new_n518), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n519), .A2(new_n298), .ZN(new_n520));
  OAI21_X1  g334(.A(new_n463), .B1(new_n505), .B2(new_n520), .ZN(new_n521));
  INV_X1    g335(.A(KEYINPUT84), .ZN(new_n522));
  NAND3_X1  g336(.A1(new_n490), .A2(new_n502), .A3(new_n504), .ZN(new_n523));
  NAND4_X1  g337(.A1(new_n523), .A2(new_n298), .A3(new_n462), .A4(new_n519), .ZN(new_n524));
  NAND3_X1  g338(.A1(new_n521), .A2(new_n522), .A3(new_n524), .ZN(new_n525));
  OAI211_X1 g339(.A(KEYINPUT84), .B(new_n463), .C1(new_n505), .C2(new_n520), .ZN(new_n526));
  OAI21_X1  g340(.A(G214), .B1(G237), .B2(G902), .ZN(new_n527));
  XOR2_X1   g341(.A(new_n527), .B(KEYINPUT79), .Z(new_n528));
  NAND2_X1  g342(.A1(G234), .A2(G237), .ZN(new_n529));
  NAND3_X1  g343(.A1(new_n529), .A2(G952), .A3(new_n277), .ZN(new_n530));
  INV_X1    g344(.A(new_n530), .ZN(new_n531));
  NAND3_X1  g345(.A1(new_n529), .A2(G902), .A3(G953), .ZN(new_n532));
  INV_X1    g346(.A(new_n532), .ZN(new_n533));
  XNOR2_X1  g347(.A(KEYINPUT21), .B(G898), .ZN(new_n534));
  AOI21_X1  g348(.A(new_n531), .B1(new_n533), .B2(new_n534), .ZN(new_n535));
  NOR2_X1   g349(.A1(new_n528), .A2(new_n535), .ZN(new_n536));
  NAND3_X1  g350(.A1(new_n525), .A2(new_n526), .A3(new_n536), .ZN(new_n537));
  NOR2_X1   g351(.A1(new_n461), .A2(new_n537), .ZN(new_n538));
  OAI21_X1  g352(.A(G221), .B1(new_n314), .B2(G902), .ZN(new_n539));
  AND3_X1   g353(.A1(new_n313), .A2(new_n538), .A3(new_n539), .ZN(new_n540));
  INV_X1    g354(.A(KEYINPUT23), .ZN(new_n541));
  OAI21_X1  g355(.A(new_n541), .B1(new_n464), .B2(G128), .ZN(new_n542));
  NAND3_X1  g356(.A1(new_n223), .A2(KEYINPUT23), .A3(G119), .ZN(new_n543));
  OAI211_X1 g357(.A(new_n542), .B(new_n543), .C1(G119), .C2(new_n223), .ZN(new_n544));
  XNOR2_X1  g358(.A(KEYINPUT24), .B(G110), .ZN(new_n545));
  INV_X1    g359(.A(new_n545), .ZN(new_n546));
  XNOR2_X1  g360(.A(G119), .B(G128), .ZN(new_n547));
  OAI22_X1  g361(.A1(new_n544), .A2(G110), .B1(new_n546), .B2(new_n547), .ZN(new_n548));
  NAND3_X1  g362(.A1(new_n406), .A2(new_n419), .A3(new_n548), .ZN(new_n549));
  INV_X1    g363(.A(new_n549), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n544), .A2(G110), .ZN(new_n551));
  INV_X1    g365(.A(new_n547), .ZN(new_n552));
  OAI21_X1  g366(.A(new_n551), .B1(new_n552), .B2(new_n545), .ZN(new_n553));
  AOI21_X1  g367(.A(new_n553), .B1(new_n401), .B2(new_n406), .ZN(new_n554));
  NOR2_X1   g368(.A1(new_n550), .A2(new_n554), .ZN(new_n555));
  NAND3_X1  g369(.A1(new_n277), .A2(G221), .A3(G234), .ZN(new_n556));
  XNOR2_X1  g370(.A(new_n556), .B(KEYINPUT22), .ZN(new_n557));
  XNOR2_X1  g371(.A(new_n557), .B(G137), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n555), .A2(new_n558), .ZN(new_n559));
  INV_X1    g373(.A(new_n558), .ZN(new_n560));
  OAI21_X1  g374(.A(new_n560), .B1(new_n550), .B2(new_n554), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n559), .A2(new_n561), .ZN(new_n562));
  INV_X1    g376(.A(G234), .ZN(new_n563));
  OAI21_X1  g377(.A(G217), .B1(new_n563), .B2(G902), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n564), .A2(new_n298), .ZN(new_n565));
  NOR2_X1   g379(.A1(new_n562), .A2(new_n565), .ZN(new_n566));
  NAND3_X1  g380(.A1(new_n559), .A2(new_n298), .A3(new_n561), .ZN(new_n567));
  OR2_X1    g381(.A1(new_n567), .A2(KEYINPUT25), .ZN(new_n568));
  AOI21_X1  g382(.A(new_n564), .B1(new_n567), .B2(KEYINPUT25), .ZN(new_n569));
  AOI21_X1  g383(.A(new_n566), .B1(new_n568), .B2(new_n569), .ZN(new_n570));
  INV_X1    g384(.A(new_n570), .ZN(new_n571));
  INV_X1    g385(.A(KEYINPUT30), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n260), .A2(G131), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n268), .A2(new_n573), .ZN(new_n574));
  AOI22_X1  g388(.A1(new_n219), .A2(KEYINPUT66), .B1(new_n197), .B2(new_n224), .ZN(new_n575));
  AOI21_X1  g389(.A(new_n574), .B1(new_n575), .B2(new_n222), .ZN(new_n576));
  INV_X1    g390(.A(new_n270), .ZN(new_n577));
  AOI21_X1  g391(.A(new_n495), .B1(new_n268), .B2(new_n577), .ZN(new_n578));
  OAI21_X1  g392(.A(new_n572), .B1(new_n576), .B2(new_n578), .ZN(new_n579));
  INV_X1    g393(.A(new_n574), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n226), .A2(new_n580), .ZN(new_n581));
  OAI21_X1  g395(.A(new_n198), .B1(new_n269), .B2(new_n270), .ZN(new_n582));
  NAND3_X1  g396(.A1(new_n581), .A2(KEYINPUT30), .A3(new_n582), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n476), .A2(new_n477), .ZN(new_n584));
  INV_X1    g398(.A(new_n584), .ZN(new_n585));
  NAND3_X1  g399(.A1(new_n579), .A2(new_n583), .A3(new_n585), .ZN(new_n586));
  INV_X1    g400(.A(G237), .ZN(new_n587));
  NAND3_X1  g401(.A1(new_n587), .A2(new_n277), .A3(G210), .ZN(new_n588));
  XOR2_X1   g402(.A(new_n588), .B(KEYINPUT27), .Z(new_n589));
  XNOR2_X1  g403(.A(new_n589), .B(KEYINPUT26), .ZN(new_n590));
  XNOR2_X1  g404(.A(new_n590), .B(new_n207), .ZN(new_n591));
  NAND3_X1  g405(.A1(new_n581), .A2(new_n582), .A3(new_n584), .ZN(new_n592));
  NAND3_X1  g406(.A1(new_n586), .A2(new_n591), .A3(new_n592), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n593), .A2(KEYINPUT31), .ZN(new_n594));
  INV_X1    g408(.A(new_n591), .ZN(new_n595));
  INV_X1    g409(.A(KEYINPUT28), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n592), .A2(new_n596), .ZN(new_n597));
  INV_X1    g411(.A(new_n597), .ZN(new_n598));
  XNOR2_X1  g412(.A(KEYINPUT68), .B(KEYINPUT28), .ZN(new_n599));
  INV_X1    g413(.A(new_n599), .ZN(new_n600));
  OAI21_X1  g414(.A(new_n585), .B1(new_n576), .B2(new_n578), .ZN(new_n601));
  AOI21_X1  g415(.A(new_n600), .B1(new_n601), .B2(new_n592), .ZN(new_n602));
  OAI21_X1  g416(.A(new_n595), .B1(new_n598), .B2(new_n602), .ZN(new_n603));
  INV_X1    g417(.A(KEYINPUT31), .ZN(new_n604));
  NAND4_X1  g418(.A1(new_n586), .A2(new_n604), .A3(new_n591), .A4(new_n592), .ZN(new_n605));
  NAND3_X1  g419(.A1(new_n594), .A2(new_n603), .A3(new_n605), .ZN(new_n606));
  NOR2_X1   g420(.A1(G472), .A2(G902), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n608), .A2(KEYINPUT69), .ZN(new_n609));
  INV_X1    g423(.A(KEYINPUT32), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  NAND3_X1  g425(.A1(new_n608), .A2(KEYINPUT69), .A3(KEYINPUT32), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n586), .A2(new_n592), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n614), .A2(new_n595), .ZN(new_n615));
  AND3_X1   g429(.A1(new_n581), .A2(new_n582), .A3(new_n584), .ZN(new_n616));
  AOI21_X1  g430(.A(new_n584), .B1(new_n581), .B2(new_n582), .ZN(new_n617));
  OAI21_X1  g431(.A(new_n599), .B1(new_n616), .B2(new_n617), .ZN(new_n618));
  NAND3_X1  g432(.A1(new_n618), .A2(new_n591), .A3(new_n597), .ZN(new_n619));
  INV_X1    g433(.A(KEYINPUT29), .ZN(new_n620));
  NAND3_X1  g434(.A1(new_n615), .A2(new_n619), .A3(new_n620), .ZN(new_n621));
  NAND3_X1  g435(.A1(new_n601), .A2(new_n592), .A3(KEYINPUT70), .ZN(new_n622));
  OAI21_X1  g436(.A(new_n622), .B1(KEYINPUT70), .B2(new_n592), .ZN(new_n623));
  OAI21_X1  g437(.A(new_n597), .B1(new_n623), .B2(new_n596), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n591), .A2(KEYINPUT29), .ZN(new_n625));
  OAI211_X1 g439(.A(new_n621), .B(new_n298), .C1(new_n624), .C2(new_n625), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n626), .A2(G472), .ZN(new_n627));
  AOI21_X1  g441(.A(new_n571), .B1(new_n613), .B2(new_n627), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n540), .A2(new_n628), .ZN(new_n629));
  XNOR2_X1  g443(.A(new_n629), .B(G101), .ZN(G3));
  NAND2_X1  g444(.A1(new_n454), .A2(new_n458), .ZN(new_n631));
  NOR2_X1   g445(.A1(new_n382), .A2(G902), .ZN(new_n632));
  INV_X1    g446(.A(new_n632), .ZN(new_n633));
  AND3_X1   g447(.A1(new_n372), .A2(new_n376), .A3(new_n375), .ZN(new_n634));
  AOI21_X1  g448(.A(new_n376), .B1(new_n372), .B2(new_n375), .ZN(new_n635));
  OAI21_X1  g449(.A(new_n316), .B1(new_n634), .B2(new_n635), .ZN(new_n636));
  INV_X1    g450(.A(KEYINPUT33), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n377), .A2(new_n317), .ZN(new_n638));
  NAND3_X1  g452(.A1(new_n636), .A2(new_n637), .A3(new_n638), .ZN(new_n639));
  OAI21_X1  g453(.A(new_n379), .B1(KEYINPUT95), .B2(new_n316), .ZN(new_n640));
  NOR2_X1   g454(.A1(new_n316), .A2(KEYINPUT95), .ZN(new_n641));
  OAI21_X1  g455(.A(new_n641), .B1(new_n352), .B2(new_n363), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n640), .A2(new_n642), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n643), .A2(KEYINPUT33), .ZN(new_n644));
  AOI21_X1  g458(.A(new_n633), .B1(new_n639), .B2(new_n644), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n636), .A2(new_n638), .ZN(new_n646));
  AOI21_X1  g460(.A(G478), .B1(new_n646), .B2(new_n298), .ZN(new_n647));
  OAI21_X1  g461(.A(new_n631), .B1(new_n645), .B2(new_n647), .ZN(new_n648));
  INV_X1    g462(.A(KEYINPUT96), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  OAI211_X1 g464(.A(KEYINPUT96), .B(new_n631), .C1(new_n645), .C2(new_n647), .ZN(new_n651));
  NAND2_X1  g465(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  INV_X1    g466(.A(new_n527), .ZN(new_n653));
  AOI21_X1  g467(.A(new_n653), .B1(new_n521), .B2(new_n524), .ZN(new_n654));
  INV_X1    g468(.A(new_n654), .ZN(new_n655));
  NOR2_X1   g469(.A1(new_n655), .A2(new_n535), .ZN(new_n656));
  AND2_X1   g470(.A1(new_n652), .A2(new_n656), .ZN(new_n657));
  INV_X1    g471(.A(new_n539), .ZN(new_n658));
  INV_X1    g472(.A(G472), .ZN(new_n659));
  AOI21_X1  g473(.A(new_n659), .B1(new_n606), .B2(new_n298), .ZN(new_n660));
  INV_X1    g474(.A(new_n660), .ZN(new_n661));
  NAND3_X1  g475(.A1(new_n661), .A2(new_n570), .A3(new_n608), .ZN(new_n662));
  AND2_X1   g476(.A1(new_n294), .A2(new_n281), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n276), .A2(new_n282), .ZN(new_n664));
  AOI21_X1  g478(.A(new_n663), .B1(new_n664), .B2(new_n302), .ZN(new_n665));
  AOI21_X1  g479(.A(new_n300), .B1(new_n665), .B2(G469), .ZN(new_n666));
  AOI211_X1 g480(.A(new_n658), .B(new_n662), .C1(new_n666), .C2(new_n299), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n657), .A2(new_n667), .ZN(new_n668));
  XOR2_X1   g482(.A(new_n668), .B(KEYINPUT97), .Z(new_n669));
  XNOR2_X1  g483(.A(new_n669), .B(KEYINPUT34), .ZN(new_n670));
  XNOR2_X1  g484(.A(new_n670), .B(G104), .ZN(G6));
  AOI22_X1  g485(.A1(new_n384), .A2(new_n460), .B1(G475), .B2(new_n457), .ZN(new_n672));
  INV_X1    g486(.A(KEYINPUT98), .ZN(new_n673));
  NOR3_X1   g487(.A1(new_n443), .A2(new_n385), .A3(new_n444), .ZN(new_n674));
  AOI21_X1  g488(.A(KEYINPUT87), .B1(new_n451), .B2(KEYINPUT20), .ZN(new_n675));
  OAI21_X1  g489(.A(new_n673), .B1(new_n674), .B2(new_n675), .ZN(new_n676));
  NAND3_X1  g490(.A1(new_n445), .A2(KEYINPUT98), .A3(new_n452), .ZN(new_n677));
  NAND3_X1  g491(.A1(new_n676), .A2(new_n453), .A3(new_n677), .ZN(new_n678));
  AND3_X1   g492(.A1(new_n656), .A2(new_n672), .A3(new_n678), .ZN(new_n679));
  NAND2_X1  g493(.A1(new_n667), .A2(new_n679), .ZN(new_n680));
  XOR2_X1   g494(.A(KEYINPUT35), .B(G107), .Z(new_n681));
  XNOR2_X1  g495(.A(new_n680), .B(new_n681), .ZN(G9));
  AOI21_X1  g496(.A(new_n658), .B1(new_n666), .B2(new_n299), .ZN(new_n683));
  NAND2_X1  g497(.A1(new_n661), .A2(new_n608), .ZN(new_n684));
  INV_X1    g498(.A(new_n565), .ZN(new_n685));
  NOR2_X1   g499(.A1(new_n560), .A2(KEYINPUT36), .ZN(new_n686));
  XOR2_X1   g500(.A(new_n555), .B(new_n686), .Z(new_n687));
  AOI22_X1  g501(.A1(new_n568), .A2(new_n569), .B1(new_n685), .B2(new_n687), .ZN(new_n688));
  NOR2_X1   g502(.A1(new_n684), .A2(new_n688), .ZN(new_n689));
  NAND3_X1  g503(.A1(new_n683), .A2(new_n538), .A3(new_n689), .ZN(new_n690));
  XOR2_X1   g504(.A(KEYINPUT37), .B(G110), .Z(new_n691));
  XNOR2_X1  g505(.A(new_n690), .B(new_n691), .ZN(G12));
  NAND2_X1  g506(.A1(new_n312), .A2(new_n301), .ZN(new_n693));
  AOI211_X1 g507(.A(G469), .B(G902), .C1(new_n283), .C2(new_n295), .ZN(new_n694));
  OAI21_X1  g508(.A(new_n539), .B1(new_n693), .B2(new_n694), .ZN(new_n695));
  AOI21_X1  g509(.A(KEYINPUT32), .B1(new_n608), .B2(KEYINPUT69), .ZN(new_n696));
  INV_X1    g510(.A(KEYINPUT69), .ZN(new_n697));
  AOI211_X1 g511(.A(new_n697), .B(new_n610), .C1(new_n606), .C2(new_n607), .ZN(new_n698));
  OAI21_X1  g512(.A(new_n627), .B1(new_n696), .B2(new_n698), .ZN(new_n699));
  NOR2_X1   g513(.A1(new_n655), .A2(new_n688), .ZN(new_n700));
  NAND2_X1  g514(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  NOR2_X1   g515(.A1(new_n695), .A2(new_n701), .ZN(new_n702));
  INV_X1    g516(.A(KEYINPUT101), .ZN(new_n703));
  INV_X1    g517(.A(KEYINPUT100), .ZN(new_n704));
  INV_X1    g518(.A(G900), .ZN(new_n705));
  NAND2_X1  g519(.A1(new_n533), .A2(new_n705), .ZN(new_n706));
  AOI21_X1  g520(.A(new_n531), .B1(new_n706), .B2(KEYINPUT99), .ZN(new_n707));
  OAI21_X1  g521(.A(new_n707), .B1(KEYINPUT99), .B2(new_n706), .ZN(new_n708));
  NAND4_X1  g522(.A1(new_n672), .A2(new_n704), .A3(new_n678), .A4(new_n708), .ZN(new_n709));
  NAND2_X1  g523(.A1(new_n384), .A2(new_n460), .ZN(new_n710));
  NAND4_X1  g524(.A1(new_n710), .A2(new_n678), .A3(new_n458), .A4(new_n708), .ZN(new_n711));
  NAND2_X1  g525(.A1(new_n711), .A2(KEYINPUT100), .ZN(new_n712));
  NAND4_X1  g526(.A1(new_n702), .A2(new_n703), .A3(new_n709), .A4(new_n712), .ZN(new_n713));
  NAND2_X1  g527(.A1(new_n712), .A2(new_n709), .ZN(new_n714));
  NAND4_X1  g528(.A1(new_n313), .A2(new_n699), .A3(new_n539), .A4(new_n700), .ZN(new_n715));
  OAI21_X1  g529(.A(KEYINPUT101), .B1(new_n714), .B2(new_n715), .ZN(new_n716));
  NAND2_X1  g530(.A1(new_n713), .A2(new_n716), .ZN(new_n717));
  XNOR2_X1  g531(.A(new_n717), .B(KEYINPUT102), .ZN(new_n718));
  XNOR2_X1  g532(.A(new_n718), .B(new_n223), .ZN(G30));
  NAND2_X1  g533(.A1(new_n525), .A2(new_n526), .ZN(new_n720));
  XOR2_X1   g534(.A(new_n720), .B(KEYINPUT38), .Z(new_n721));
  NAND2_X1  g535(.A1(new_n623), .A2(new_n595), .ZN(new_n722));
  NAND2_X1  g536(.A1(new_n614), .A2(new_n591), .ZN(new_n723));
  NAND3_X1  g537(.A1(new_n722), .A2(new_n298), .A3(new_n723), .ZN(new_n724));
  NAND2_X1  g538(.A1(new_n724), .A2(G472), .ZN(new_n725));
  INV_X1    g539(.A(KEYINPUT103), .ZN(new_n726));
  XNOR2_X1  g540(.A(new_n725), .B(new_n726), .ZN(new_n727));
  NAND2_X1  g541(.A1(new_n613), .A2(new_n727), .ZN(new_n728));
  AND2_X1   g542(.A1(new_n710), .A2(new_n631), .ZN(new_n729));
  INV_X1    g543(.A(new_n688), .ZN(new_n730));
  NOR2_X1   g544(.A1(new_n730), .A2(new_n653), .ZN(new_n731));
  NAND4_X1  g545(.A1(new_n721), .A2(new_n728), .A3(new_n729), .A4(new_n731), .ZN(new_n732));
  XOR2_X1   g546(.A(new_n732), .B(KEYINPUT104), .Z(new_n733));
  XNOR2_X1  g547(.A(new_n708), .B(KEYINPUT39), .ZN(new_n734));
  NAND2_X1  g548(.A1(new_n683), .A2(new_n734), .ZN(new_n735));
  OR2_X1    g549(.A1(new_n735), .A2(KEYINPUT40), .ZN(new_n736));
  NAND2_X1  g550(.A1(new_n735), .A2(KEYINPUT40), .ZN(new_n737));
  NAND3_X1  g551(.A1(new_n733), .A2(new_n736), .A3(new_n737), .ZN(new_n738));
  XNOR2_X1  g552(.A(new_n738), .B(KEYINPUT105), .ZN(new_n739));
  XNOR2_X1  g553(.A(new_n739), .B(new_n190), .ZN(G45));
  OAI211_X1 g554(.A(new_n631), .B(new_n708), .C1(new_n645), .C2(new_n647), .ZN(new_n741));
  NOR2_X1   g555(.A1(new_n715), .A2(new_n741), .ZN(new_n742));
  XNOR2_X1  g556(.A(new_n742), .B(new_n187), .ZN(G48));
  AOI21_X1  g557(.A(new_n297), .B1(new_n296), .B2(new_n298), .ZN(new_n744));
  NOR3_X1   g558(.A1(new_n744), .A2(new_n694), .A3(new_n658), .ZN(new_n745));
  NAND4_X1  g559(.A1(new_n652), .A2(new_n745), .A3(new_n628), .A4(new_n656), .ZN(new_n746));
  XOR2_X1   g560(.A(new_n746), .B(KEYINPUT106), .Z(new_n747));
  XNOR2_X1  g561(.A(new_n747), .B(KEYINPUT107), .ZN(new_n748));
  XNOR2_X1  g562(.A(KEYINPUT41), .B(G113), .ZN(new_n749));
  XNOR2_X1  g563(.A(new_n748), .B(new_n749), .ZN(G15));
  NAND3_X1  g564(.A1(new_n679), .A2(new_n745), .A3(new_n628), .ZN(new_n751));
  XNOR2_X1  g565(.A(new_n751), .B(G116), .ZN(G18));
  NAND2_X1  g566(.A1(new_n296), .A2(new_n298), .ZN(new_n753));
  NAND2_X1  g567(.A1(new_n753), .A2(G469), .ZN(new_n754));
  NAND4_X1  g568(.A1(new_n754), .A2(new_n539), .A3(new_n299), .A4(new_n654), .ZN(new_n755));
  INV_X1    g569(.A(KEYINPUT108), .ZN(new_n756));
  NAND2_X1  g570(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  NOR2_X1   g571(.A1(new_n744), .A2(new_n694), .ZN(new_n758));
  NAND4_X1  g572(.A1(new_n758), .A2(KEYINPUT108), .A3(new_n539), .A4(new_n654), .ZN(new_n759));
  NAND2_X1  g573(.A1(new_n757), .A2(new_n759), .ZN(new_n760));
  INV_X1    g574(.A(new_n699), .ZN(new_n761));
  NOR4_X1   g575(.A1(new_n761), .A2(new_n461), .A3(new_n535), .A4(new_n688), .ZN(new_n762));
  NAND2_X1  g576(.A1(new_n760), .A2(new_n762), .ZN(new_n763));
  XNOR2_X1  g577(.A(new_n763), .B(G119), .ZN(G21));
  INV_X1    g578(.A(new_n607), .ZN(new_n765));
  NAND2_X1  g579(.A1(new_n624), .A2(new_n595), .ZN(new_n766));
  AND2_X1   g580(.A1(new_n594), .A2(new_n605), .ZN(new_n767));
  AOI21_X1  g581(.A(new_n765), .B1(new_n766), .B2(new_n767), .ZN(new_n768));
  NOR3_X1   g582(.A1(new_n571), .A2(new_n768), .A3(new_n660), .ZN(new_n769));
  NAND3_X1  g583(.A1(new_n729), .A2(new_n769), .A3(new_n656), .ZN(new_n770));
  NAND3_X1  g584(.A1(new_n754), .A2(new_n539), .A3(new_n299), .ZN(new_n771));
  NOR2_X1   g585(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  XNOR2_X1  g586(.A(new_n772), .B(new_n340), .ZN(G24));
  OR3_X1    g587(.A1(new_n688), .A2(new_n768), .A3(new_n660), .ZN(new_n774));
  NOR2_X1   g588(.A1(new_n774), .A2(new_n741), .ZN(new_n775));
  NAND2_X1  g589(.A1(new_n760), .A2(new_n775), .ZN(new_n776));
  XNOR2_X1  g590(.A(new_n776), .B(G125), .ZN(G27));
  INV_X1    g591(.A(new_n741), .ZN(new_n778));
  AOI21_X1  g592(.A(new_n653), .B1(new_n525), .B2(new_n526), .ZN(new_n779));
  AND2_X1   g593(.A1(new_n779), .A2(new_n539), .ZN(new_n780));
  INV_X1    g594(.A(KEYINPUT109), .ZN(new_n781));
  AOI21_X1  g595(.A(new_n781), .B1(new_n294), .B2(new_n281), .ZN(new_n782));
  INV_X1    g596(.A(new_n782), .ZN(new_n783));
  NAND3_X1  g597(.A1(new_n294), .A2(new_n781), .A3(new_n281), .ZN(new_n784));
  NAND4_X1  g598(.A1(new_n310), .A2(new_n783), .A3(G469), .A4(new_n784), .ZN(new_n785));
  NAND3_X1  g599(.A1(new_n299), .A2(new_n301), .A3(new_n785), .ZN(new_n786));
  NAND4_X1  g600(.A1(new_n628), .A2(new_n778), .A3(new_n780), .A4(new_n786), .ZN(new_n787));
  INV_X1    g601(.A(KEYINPUT42), .ZN(new_n788));
  NAND2_X1  g602(.A1(new_n779), .A2(new_n539), .ZN(new_n789));
  AOI21_X1  g603(.A(new_n281), .B1(new_n276), .B2(new_n282), .ZN(new_n790));
  AND3_X1   g604(.A1(new_n294), .A2(new_n781), .A3(new_n281), .ZN(new_n791));
  NOR3_X1   g605(.A1(new_n790), .A2(new_n791), .A3(new_n782), .ZN(new_n792));
  AOI21_X1  g606(.A(new_n300), .B1(new_n792), .B2(G469), .ZN(new_n793));
  AOI21_X1  g607(.A(new_n789), .B1(new_n793), .B2(new_n299), .ZN(new_n794));
  NAND3_X1  g608(.A1(new_n606), .A2(KEYINPUT32), .A3(new_n607), .ZN(new_n795));
  NAND2_X1  g609(.A1(new_n608), .A2(new_n610), .ZN(new_n796));
  NAND3_X1  g610(.A1(new_n627), .A2(new_n795), .A3(new_n796), .ZN(new_n797));
  NAND2_X1  g611(.A1(new_n797), .A2(new_n570), .ZN(new_n798));
  NOR3_X1   g612(.A1(new_n798), .A2(new_n788), .A3(new_n741), .ZN(new_n799));
  AOI22_X1  g613(.A1(new_n787), .A2(new_n788), .B1(new_n794), .B2(new_n799), .ZN(new_n800));
  XNOR2_X1  g614(.A(new_n800), .B(new_n267), .ZN(G33));
  NAND4_X1  g615(.A1(new_n794), .A2(new_n628), .A3(new_n709), .A4(new_n712), .ZN(new_n802));
  XNOR2_X1  g616(.A(new_n802), .B(G134), .ZN(G36));
  NAND2_X1  g617(.A1(new_n792), .A2(KEYINPUT45), .ZN(new_n804));
  OAI211_X1 g618(.A(new_n804), .B(G469), .C1(KEYINPUT45), .C2(new_n665), .ZN(new_n805));
  AOI21_X1  g619(.A(KEYINPUT46), .B1(new_n805), .B2(new_n301), .ZN(new_n806));
  NAND3_X1  g620(.A1(new_n805), .A2(KEYINPUT46), .A3(new_n301), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n807), .A2(new_n299), .ZN(new_n808));
  AOI21_X1  g622(.A(new_n806), .B1(new_n808), .B2(KEYINPUT110), .ZN(new_n809));
  INV_X1    g623(.A(KEYINPUT110), .ZN(new_n810));
  NAND3_X1  g624(.A1(new_n807), .A2(new_n810), .A3(new_n299), .ZN(new_n811));
  NAND2_X1  g625(.A1(new_n809), .A2(new_n811), .ZN(new_n812));
  AND3_X1   g626(.A1(new_n812), .A2(new_n539), .A3(new_n734), .ZN(new_n813));
  OAI211_X1 g627(.A(new_n454), .B(new_n458), .C1(new_n645), .C2(new_n647), .ZN(new_n814));
  OR2_X1    g628(.A1(new_n814), .A2(KEYINPUT43), .ZN(new_n815));
  NAND2_X1  g629(.A1(new_n814), .A2(KEYINPUT43), .ZN(new_n816));
  NAND4_X1  g630(.A1(new_n815), .A2(new_n684), .A3(new_n730), .A4(new_n816), .ZN(new_n817));
  INV_X1    g631(.A(KEYINPUT44), .ZN(new_n818));
  AND2_X1   g632(.A1(new_n817), .A2(new_n818), .ZN(new_n819));
  NOR2_X1   g633(.A1(new_n817), .A2(new_n818), .ZN(new_n820));
  INV_X1    g634(.A(new_n779), .ZN(new_n821));
  NOR3_X1   g635(.A1(new_n819), .A2(new_n820), .A3(new_n821), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n813), .A2(new_n822), .ZN(new_n823));
  XNOR2_X1  g637(.A(new_n823), .B(G137), .ZN(G39));
  AOI211_X1 g638(.A(KEYINPUT47), .B(new_n658), .C1(new_n809), .C2(new_n811), .ZN(new_n825));
  INV_X1    g639(.A(KEYINPUT47), .ZN(new_n826));
  AOI21_X1  g640(.A(new_n826), .B1(new_n812), .B2(new_n539), .ZN(new_n827));
  NAND3_X1  g641(.A1(new_n761), .A2(new_n571), .A3(new_n779), .ZN(new_n828));
  OR4_X1    g642(.A1(new_n741), .A2(new_n825), .A3(new_n827), .A4(new_n828), .ZN(new_n829));
  XNOR2_X1  g643(.A(new_n829), .B(G140), .ZN(G42));
  NAND2_X1  g644(.A1(new_n381), .A2(new_n382), .ZN(new_n831));
  AOI21_X1  g645(.A(new_n637), .B1(new_n640), .B2(new_n642), .ZN(new_n832));
  NAND2_X1  g646(.A1(new_n364), .A2(new_n377), .ZN(new_n833));
  AOI21_X1  g647(.A(new_n380), .B1(new_n833), .B2(new_n316), .ZN(new_n834));
  AOI21_X1  g648(.A(new_n832), .B1(new_n834), .B2(new_n637), .ZN(new_n835));
  OAI211_X1 g649(.A(new_n631), .B(new_n831), .C1(new_n835), .C2(new_n633), .ZN(new_n836));
  NAND3_X1  g650(.A1(new_n836), .A2(KEYINPUT111), .A3(new_n461), .ZN(new_n837));
  INV_X1    g651(.A(KEYINPUT111), .ZN(new_n838));
  NAND2_X1  g652(.A1(new_n648), .A2(new_n838), .ZN(new_n839));
  NAND2_X1  g653(.A1(new_n837), .A2(new_n839), .ZN(new_n840));
  INV_X1    g654(.A(new_n537), .ZN(new_n841));
  INV_X1    g655(.A(new_n662), .ZN(new_n842));
  NAND4_X1  g656(.A1(new_n840), .A2(new_n683), .A3(new_n841), .A4(new_n842), .ZN(new_n843));
  NAND4_X1  g657(.A1(new_n843), .A2(new_n746), .A3(new_n690), .A4(new_n751), .ZN(new_n844));
  AND3_X1   g658(.A1(new_n729), .A2(new_n769), .A3(new_n656), .ZN(new_n845));
  NAND2_X1  g659(.A1(new_n845), .A2(new_n745), .ZN(new_n846));
  NAND2_X1  g660(.A1(new_n629), .A2(new_n846), .ZN(new_n847));
  NOR2_X1   g661(.A1(new_n844), .A2(new_n847), .ZN(new_n848));
  AND2_X1   g662(.A1(new_n458), .A2(new_n708), .ZN(new_n849));
  NAND4_X1  g663(.A1(new_n678), .A2(new_n384), .A3(new_n460), .A4(new_n849), .ZN(new_n850));
  OAI21_X1  g664(.A(KEYINPUT112), .B1(new_n850), .B2(new_n821), .ZN(new_n851));
  AOI21_X1  g665(.A(new_n688), .B1(new_n613), .B2(new_n627), .ZN(new_n852));
  AND3_X1   g666(.A1(new_n384), .A2(new_n460), .A3(new_n849), .ZN(new_n853));
  INV_X1    g667(.A(KEYINPUT112), .ZN(new_n854));
  NAND4_X1  g668(.A1(new_n853), .A2(new_n854), .A3(new_n678), .A4(new_n779), .ZN(new_n855));
  NAND4_X1  g669(.A1(new_n851), .A2(new_n683), .A3(new_n852), .A4(new_n855), .ZN(new_n856));
  NAND2_X1  g670(.A1(new_n794), .A2(new_n775), .ZN(new_n857));
  NAND3_X1  g671(.A1(new_n802), .A2(new_n856), .A3(new_n857), .ZN(new_n858));
  NOR2_X1   g672(.A1(new_n858), .A2(new_n800), .ZN(new_n859));
  NAND3_X1  g673(.A1(new_n848), .A2(new_n859), .A3(new_n763), .ZN(new_n860));
  INV_X1    g674(.A(new_n728), .ZN(new_n861));
  AND3_X1   g675(.A1(new_n688), .A2(new_n539), .A3(new_n708), .ZN(new_n862));
  NAND4_X1  g676(.A1(new_n862), .A2(new_n631), .A3(new_n710), .A4(new_n654), .ZN(new_n863));
  NOR2_X1   g677(.A1(new_n861), .A2(new_n863), .ZN(new_n864));
  AOI22_X1  g678(.A1(new_n864), .A2(new_n786), .B1(new_n702), .B2(new_n778), .ZN(new_n865));
  NAND3_X1  g679(.A1(new_n717), .A2(new_n776), .A3(new_n865), .ZN(new_n866));
  INV_X1    g680(.A(KEYINPUT52), .ZN(new_n867));
  NAND2_X1  g681(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  AOI22_X1  g682(.A1(new_n713), .A2(new_n716), .B1(new_n760), .B2(new_n775), .ZN(new_n869));
  NAND3_X1  g683(.A1(new_n869), .A2(KEYINPUT52), .A3(new_n865), .ZN(new_n870));
  AOI21_X1  g684(.A(new_n860), .B1(new_n868), .B2(new_n870), .ZN(new_n871));
  OAI21_X1  g685(.A(KEYINPUT113), .B1(new_n871), .B2(KEYINPUT53), .ZN(new_n872));
  AND2_X1   g686(.A1(new_n746), .A2(new_n690), .ZN(new_n873));
  NAND2_X1  g687(.A1(new_n699), .A2(new_n570), .ZN(new_n874));
  NOR2_X1   g688(.A1(new_n771), .A2(new_n874), .ZN(new_n875));
  AOI21_X1  g689(.A(new_n537), .B1(new_n837), .B2(new_n839), .ZN(new_n876));
  AOI22_X1  g690(.A1(new_n679), .A2(new_n875), .B1(new_n876), .B2(new_n667), .ZN(new_n877));
  AOI22_X1  g691(.A1(new_n540), .A2(new_n628), .B1(new_n845), .B2(new_n745), .ZN(new_n878));
  NAND4_X1  g692(.A1(new_n873), .A2(new_n877), .A3(new_n763), .A4(new_n878), .ZN(new_n879));
  NAND4_X1  g693(.A1(new_n786), .A2(new_n780), .A3(new_n699), .A4(new_n570), .ZN(new_n880));
  OAI21_X1  g694(.A(new_n788), .B1(new_n880), .B2(new_n741), .ZN(new_n881));
  NAND2_X1  g695(.A1(new_n799), .A2(new_n794), .ZN(new_n882));
  NAND2_X1  g696(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  NAND4_X1  g697(.A1(new_n883), .A2(new_n802), .A3(new_n856), .A4(new_n857), .ZN(new_n884));
  NOR2_X1   g698(.A1(new_n879), .A2(new_n884), .ZN(new_n885));
  NOR2_X1   g699(.A1(new_n866), .A2(new_n867), .ZN(new_n886));
  AOI21_X1  g700(.A(KEYINPUT52), .B1(new_n869), .B2(new_n865), .ZN(new_n887));
  OAI21_X1  g701(.A(new_n885), .B1(new_n886), .B2(new_n887), .ZN(new_n888));
  INV_X1    g702(.A(KEYINPUT113), .ZN(new_n889));
  INV_X1    g703(.A(KEYINPUT53), .ZN(new_n890));
  NAND3_X1  g704(.A1(new_n888), .A2(new_n889), .A3(new_n890), .ZN(new_n891));
  NAND2_X1  g705(.A1(new_n872), .A2(new_n891), .ZN(new_n892));
  INV_X1    g706(.A(KEYINPUT54), .ZN(new_n893));
  OAI211_X1 g707(.A(KEYINPUT53), .B(new_n885), .C1(new_n886), .C2(new_n887), .ZN(new_n894));
  NAND2_X1  g708(.A1(new_n894), .A2(KEYINPUT114), .ZN(new_n895));
  NAND2_X1  g709(.A1(new_n868), .A2(new_n870), .ZN(new_n896));
  INV_X1    g710(.A(KEYINPUT114), .ZN(new_n897));
  NAND4_X1  g711(.A1(new_n896), .A2(new_n897), .A3(KEYINPUT53), .A4(new_n885), .ZN(new_n898));
  NAND2_X1  g712(.A1(new_n895), .A2(new_n898), .ZN(new_n899));
  AND3_X1   g713(.A1(new_n892), .A2(new_n893), .A3(new_n899), .ZN(new_n900));
  NAND2_X1  g714(.A1(new_n888), .A2(new_n890), .ZN(new_n901));
  AND2_X1   g715(.A1(new_n901), .A2(new_n894), .ZN(new_n902));
  NOR2_X1   g716(.A1(new_n902), .A2(new_n893), .ZN(new_n903));
  NOR2_X1   g717(.A1(new_n900), .A2(new_n903), .ZN(new_n904));
  AND3_X1   g718(.A1(new_n815), .A2(new_n531), .A3(new_n816), .ZN(new_n905));
  NAND2_X1  g719(.A1(new_n905), .A2(new_n769), .ZN(new_n906));
  OR2_X1    g720(.A1(new_n721), .A2(new_n527), .ZN(new_n907));
  NOR3_X1   g721(.A1(new_n906), .A2(new_n771), .A3(new_n907), .ZN(new_n908));
  XNOR2_X1  g722(.A(new_n908), .B(KEYINPUT50), .ZN(new_n909));
  INV_X1    g723(.A(KEYINPUT116), .ZN(new_n910));
  INV_X1    g724(.A(new_n758), .ZN(new_n911));
  NOR2_X1   g725(.A1(new_n911), .A2(new_n789), .ZN(new_n912));
  NAND2_X1  g726(.A1(new_n905), .A2(new_n912), .ZN(new_n913));
  NOR2_X1   g727(.A1(new_n913), .A2(new_n774), .ZN(new_n914));
  INV_X1    g728(.A(new_n912), .ZN(new_n915));
  NOR4_X1   g729(.A1(new_n915), .A2(new_n571), .A3(new_n530), .A4(new_n728), .ZN(new_n916));
  NOR3_X1   g730(.A1(new_n645), .A2(new_n631), .A3(new_n647), .ZN(new_n917));
  AOI21_X1  g731(.A(new_n914), .B1(new_n916), .B2(new_n917), .ZN(new_n918));
  AND3_X1   g732(.A1(new_n909), .A2(new_n910), .A3(new_n918), .ZN(new_n919));
  AOI21_X1  g733(.A(new_n910), .B1(new_n909), .B2(new_n918), .ZN(new_n920));
  NOR2_X1   g734(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  OAI22_X1  g735(.A1(new_n827), .A2(new_n825), .B1(new_n539), .B2(new_n911), .ZN(new_n922));
  NOR2_X1   g736(.A1(new_n906), .A2(new_n821), .ZN(new_n923));
  XNOR2_X1  g737(.A(new_n923), .B(KEYINPUT115), .ZN(new_n924));
  NAND2_X1  g738(.A1(new_n922), .A2(new_n924), .ZN(new_n925));
  AOI21_X1  g739(.A(KEYINPUT51), .B1(new_n921), .B2(new_n925), .ZN(new_n926));
  NOR2_X1   g740(.A1(new_n913), .A2(new_n798), .ZN(new_n927));
  XOR2_X1   g741(.A(new_n927), .B(KEYINPUT48), .Z(new_n928));
  NAND3_X1  g742(.A1(new_n760), .A2(new_n905), .A3(new_n769), .ZN(new_n929));
  INV_X1    g743(.A(G952), .ZN(new_n930));
  AOI211_X1 g744(.A(new_n930), .B(G953), .C1(new_n916), .C2(new_n652), .ZN(new_n931));
  AND3_X1   g745(.A1(new_n928), .A2(new_n929), .A3(new_n931), .ZN(new_n932));
  INV_X1    g746(.A(new_n925), .ZN(new_n933));
  INV_X1    g747(.A(KEYINPUT117), .ZN(new_n934));
  OR2_X1    g748(.A1(new_n918), .A2(new_n934), .ZN(new_n935));
  NAND2_X1  g749(.A1(new_n918), .A2(new_n934), .ZN(new_n936));
  NAND4_X1  g750(.A1(new_n935), .A2(KEYINPUT51), .A3(new_n909), .A4(new_n936), .ZN(new_n937));
  OAI21_X1  g751(.A(new_n932), .B1(new_n933), .B2(new_n937), .ZN(new_n938));
  NOR2_X1   g752(.A1(new_n926), .A2(new_n938), .ZN(new_n939));
  NAND2_X1  g753(.A1(new_n904), .A2(new_n939), .ZN(new_n940));
  AOI22_X1  g754(.A1(new_n940), .A2(KEYINPUT118), .B1(new_n930), .B2(new_n277), .ZN(new_n941));
  OAI21_X1  g755(.A(new_n941), .B1(KEYINPUT118), .B2(new_n940), .ZN(new_n942));
  OR4_X1    g756(.A1(new_n571), .A2(new_n721), .A3(new_n658), .A4(new_n528), .ZN(new_n943));
  XOR2_X1   g757(.A(new_n758), .B(KEYINPUT49), .Z(new_n944));
  OR4_X1    g758(.A1(new_n728), .A2(new_n943), .A3(new_n814), .A4(new_n944), .ZN(new_n945));
  NAND2_X1  g759(.A1(new_n942), .A2(new_n945), .ZN(G75));
  NOR2_X1   g760(.A1(new_n277), .A2(G952), .ZN(new_n947));
  INV_X1    g761(.A(new_n947), .ZN(new_n948));
  NOR3_X1   g762(.A1(new_n871), .A2(KEYINPUT113), .A3(KEYINPUT53), .ZN(new_n949));
  AOI21_X1  g763(.A(new_n889), .B1(new_n888), .B2(new_n890), .ZN(new_n950));
  NOR2_X1   g764(.A1(new_n949), .A2(new_n950), .ZN(new_n951));
  AND2_X1   g765(.A1(new_n895), .A2(new_n898), .ZN(new_n952));
  NOR2_X1   g766(.A1(new_n951), .A2(new_n952), .ZN(new_n953));
  NOR2_X1   g767(.A1(new_n953), .A2(new_n298), .ZN(new_n954));
  AOI21_X1  g768(.A(KEYINPUT56), .B1(new_n954), .B2(G210), .ZN(new_n955));
  NAND2_X1  g769(.A1(new_n490), .A2(new_n504), .ZN(new_n956));
  XNOR2_X1  g770(.A(new_n956), .B(new_n502), .ZN(new_n957));
  XNOR2_X1  g771(.A(new_n957), .B(KEYINPUT55), .ZN(new_n958));
  OAI21_X1  g772(.A(new_n948), .B1(new_n955), .B2(new_n958), .ZN(new_n959));
  NAND2_X1  g773(.A1(new_n955), .A2(new_n958), .ZN(new_n960));
  NAND2_X1  g774(.A1(new_n960), .A2(KEYINPUT119), .ZN(new_n961));
  INV_X1    g775(.A(KEYINPUT119), .ZN(new_n962));
  NAND3_X1  g776(.A1(new_n955), .A2(new_n962), .A3(new_n958), .ZN(new_n963));
  AOI21_X1  g777(.A(new_n959), .B1(new_n961), .B2(new_n963), .ZN(G51));
  AOI21_X1  g778(.A(new_n893), .B1(new_n892), .B2(new_n899), .ZN(new_n965));
  NOR2_X1   g779(.A1(new_n900), .A2(new_n965), .ZN(new_n966));
  XOR2_X1   g780(.A(new_n300), .B(KEYINPUT57), .Z(new_n967));
  OAI21_X1  g781(.A(new_n296), .B1(new_n966), .B2(new_n967), .ZN(new_n968));
  XNOR2_X1  g782(.A(new_n805), .B(KEYINPUT120), .ZN(new_n969));
  NAND2_X1  g783(.A1(new_n954), .A2(new_n969), .ZN(new_n970));
  AOI21_X1  g784(.A(new_n947), .B1(new_n968), .B2(new_n970), .ZN(G54));
  NAND3_X1  g785(.A1(new_n954), .A2(KEYINPUT58), .A3(G475), .ZN(new_n972));
  NAND2_X1  g786(.A1(new_n448), .A2(new_n450), .ZN(new_n973));
  AND2_X1   g787(.A1(new_n972), .A2(new_n973), .ZN(new_n974));
  NOR2_X1   g788(.A1(new_n972), .A2(new_n973), .ZN(new_n975));
  NOR3_X1   g789(.A1(new_n974), .A2(new_n975), .A3(new_n947), .ZN(G60));
  NAND2_X1  g790(.A1(G478), .A2(G902), .ZN(new_n977));
  XOR2_X1   g791(.A(new_n977), .B(KEYINPUT59), .Z(new_n978));
  OR2_X1    g792(.A1(new_n835), .A2(new_n978), .ZN(new_n979));
  OAI21_X1  g793(.A(KEYINPUT54), .B1(new_n951), .B2(new_n952), .ZN(new_n980));
  NAND3_X1  g794(.A1(new_n892), .A2(new_n893), .A3(new_n899), .ZN(new_n981));
  AOI21_X1  g795(.A(new_n979), .B1(new_n980), .B2(new_n981), .ZN(new_n982));
  OAI21_X1  g796(.A(KEYINPUT121), .B1(new_n982), .B2(new_n947), .ZN(new_n983));
  INV_X1    g797(.A(KEYINPUT121), .ZN(new_n984));
  OAI211_X1 g798(.A(new_n984), .B(new_n948), .C1(new_n966), .C2(new_n979), .ZN(new_n985));
  OAI21_X1  g799(.A(new_n835), .B1(new_n904), .B2(new_n978), .ZN(new_n986));
  NAND3_X1  g800(.A1(new_n983), .A2(new_n985), .A3(new_n986), .ZN(new_n987));
  INV_X1    g801(.A(KEYINPUT122), .ZN(new_n988));
  NAND2_X1  g802(.A1(new_n987), .A2(new_n988), .ZN(new_n989));
  NAND4_X1  g803(.A1(new_n983), .A2(new_n985), .A3(new_n986), .A4(KEYINPUT122), .ZN(new_n990));
  NAND2_X1  g804(.A1(new_n989), .A2(new_n990), .ZN(G63));
  NAND2_X1  g805(.A1(G217), .A2(G902), .ZN(new_n992));
  XNOR2_X1  g806(.A(new_n992), .B(KEYINPUT60), .ZN(new_n993));
  INV_X1    g807(.A(new_n993), .ZN(new_n994));
  OAI211_X1 g808(.A(new_n687), .B(new_n994), .C1(new_n951), .C2(new_n952), .ZN(new_n995));
  NAND3_X1  g809(.A1(new_n995), .A2(KEYINPUT123), .A3(new_n948), .ZN(new_n996));
  INV_X1    g810(.A(KEYINPUT124), .ZN(new_n997));
  AND3_X1   g811(.A1(new_n996), .A2(new_n997), .A3(KEYINPUT61), .ZN(new_n998));
  AOI21_X1  g812(.A(new_n997), .B1(new_n996), .B2(KEYINPUT61), .ZN(new_n999));
  OAI21_X1  g813(.A(new_n562), .B1(new_n953), .B2(new_n993), .ZN(new_n1000));
  NAND3_X1  g814(.A1(new_n1000), .A2(new_n948), .A3(new_n995), .ZN(new_n1001));
  NOR3_X1   g815(.A1(new_n998), .A2(new_n999), .A3(new_n1001), .ZN(new_n1002));
  AND3_X1   g816(.A1(new_n1000), .A2(new_n948), .A3(new_n995), .ZN(new_n1003));
  INV_X1    g817(.A(KEYINPUT123), .ZN(new_n1004));
  AOI21_X1  g818(.A(new_n993), .B1(new_n892), .B2(new_n899), .ZN(new_n1005));
  AOI211_X1 g819(.A(new_n1004), .B(new_n947), .C1(new_n1005), .C2(new_n687), .ZN(new_n1006));
  INV_X1    g820(.A(KEYINPUT61), .ZN(new_n1007));
  OAI21_X1  g821(.A(KEYINPUT124), .B1(new_n1006), .B2(new_n1007), .ZN(new_n1008));
  NAND3_X1  g822(.A1(new_n996), .A2(new_n997), .A3(KEYINPUT61), .ZN(new_n1009));
  AOI21_X1  g823(.A(new_n1003), .B1(new_n1008), .B2(new_n1009), .ZN(new_n1010));
  NOR2_X1   g824(.A1(new_n1002), .A2(new_n1010), .ZN(G66));
  NOR3_X1   g825(.A1(new_n534), .A2(new_n498), .A3(new_n277), .ZN(new_n1012));
  INV_X1    g826(.A(new_n879), .ZN(new_n1013));
  AOI21_X1  g827(.A(new_n1012), .B1(new_n1013), .B2(new_n277), .ZN(new_n1014));
  OAI21_X1  g828(.A(new_n956), .B1(G898), .B2(new_n277), .ZN(new_n1015));
  XNOR2_X1  g829(.A(new_n1014), .B(new_n1015), .ZN(G69));
  NAND3_X1  g830(.A1(G227), .A2(G900), .A3(G953), .ZN(new_n1017));
  NAND2_X1  g831(.A1(new_n579), .A2(new_n583), .ZN(new_n1018));
  XOR2_X1   g832(.A(new_n1018), .B(KEYINPUT125), .Z(new_n1019));
  XNOR2_X1  g833(.A(new_n1019), .B(new_n435), .ZN(new_n1020));
  INV_X1    g834(.A(new_n742), .ZN(new_n1021));
  NAND3_X1  g835(.A1(new_n738), .A2(new_n1021), .A3(new_n869), .ZN(new_n1022));
  XOR2_X1   g836(.A(new_n1022), .B(KEYINPUT62), .Z(new_n1023));
  NAND2_X1  g837(.A1(new_n1023), .A2(new_n829), .ZN(new_n1024));
  INV_X1    g838(.A(new_n735), .ZN(new_n1025));
  NAND4_X1  g839(.A1(new_n1025), .A2(new_n628), .A3(new_n779), .A4(new_n840), .ZN(new_n1026));
  AND2_X1   g840(.A1(new_n823), .A2(new_n1026), .ZN(new_n1027));
  NAND2_X1  g841(.A1(new_n1027), .A2(new_n277), .ZN(new_n1028));
  OAI211_X1 g842(.A(new_n1017), .B(new_n1020), .C1(new_n1024), .C2(new_n1028), .ZN(new_n1029));
  AND2_X1   g843(.A1(new_n729), .A2(new_n654), .ZN(new_n1030));
  NAND4_X1  g844(.A1(new_n813), .A2(new_n570), .A3(new_n797), .A4(new_n1030), .ZN(new_n1031));
  NAND4_X1  g845(.A1(new_n869), .A2(new_n1021), .A3(new_n883), .A4(new_n802), .ZN(new_n1032));
  AOI21_X1  g846(.A(new_n1032), .B1(new_n813), .B2(new_n822), .ZN(new_n1033));
  NAND3_X1  g847(.A1(new_n829), .A2(new_n1031), .A3(new_n1033), .ZN(new_n1034));
  AND2_X1   g848(.A1(new_n1034), .A2(new_n277), .ZN(new_n1035));
  NOR3_X1   g849(.A1(new_n705), .A2(new_n277), .A3(G227), .ZN(new_n1036));
  OR2_X1    g850(.A1(new_n1020), .A2(new_n1036), .ZN(new_n1037));
  OAI21_X1  g851(.A(new_n1029), .B1(new_n1035), .B2(new_n1037), .ZN(G72));
  XNOR2_X1  g852(.A(KEYINPUT126), .B(KEYINPUT63), .ZN(new_n1039));
  NOR2_X1   g853(.A1(new_n659), .A2(new_n298), .ZN(new_n1040));
  XNOR2_X1  g854(.A(new_n1039), .B(new_n1040), .ZN(new_n1041));
  OAI21_X1  g855(.A(new_n1041), .B1(new_n1034), .B2(new_n879), .ZN(new_n1042));
  NAND4_X1  g856(.A1(new_n1042), .A2(new_n595), .A3(new_n592), .A4(new_n586), .ZN(new_n1043));
  NAND2_X1  g857(.A1(new_n615), .A2(new_n593), .ZN(new_n1044));
  NAND2_X1  g858(.A1(new_n1044), .A2(new_n1041), .ZN(new_n1045));
  OAI211_X1 g859(.A(new_n1043), .B(new_n948), .C1(new_n902), .C2(new_n1045), .ZN(new_n1046));
  NAND2_X1  g860(.A1(new_n1027), .A2(new_n1013), .ZN(new_n1047));
  OAI21_X1  g861(.A(new_n1041), .B1(new_n1024), .B2(new_n1047), .ZN(new_n1048));
  NAND3_X1  g862(.A1(new_n1048), .A2(new_n591), .A3(new_n614), .ZN(new_n1049));
  OR2_X1    g863(.A1(new_n1049), .A2(KEYINPUT127), .ZN(new_n1050));
  NAND2_X1  g864(.A1(new_n1049), .A2(KEYINPUT127), .ZN(new_n1051));
  AOI21_X1  g865(.A(new_n1046), .B1(new_n1050), .B2(new_n1051), .ZN(G57));
endmodule


