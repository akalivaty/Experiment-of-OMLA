//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 1 1 1 0 0 0 1 0 0 0 1 1 0 1 1 1 0 0 0 0 0 0 1 1 0 0 1 1 0 0 1 1 0 1 0 1 0 1 1 0 1 0 0 0 0 1 0 0 0 0 1 0 1 1 0 1 0 1 0 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:29:43 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n437, new_n444, new_n445, new_n446, new_n451, new_n453,
    new_n456, new_n457, new_n458, new_n459, new_n460, new_n461, new_n464,
    new_n465, new_n466, new_n467, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n484, new_n485, new_n486,
    new_n487, new_n488, new_n489, new_n490, new_n491, new_n492, new_n493,
    new_n494, new_n495, new_n496, new_n497, new_n498, new_n499, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n533, new_n534, new_n535, new_n536, new_n537, new_n539,
    new_n540, new_n541, new_n542, new_n543, new_n544, new_n545, new_n546,
    new_n548, new_n549, new_n550, new_n551, new_n552, new_n553, new_n554,
    new_n555, new_n556, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n568, new_n569, new_n570, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n586, new_n587, new_n588, new_n589, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n597, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n618, new_n619, new_n622, new_n623, new_n625, new_n626,
    new_n627, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n824, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1131, new_n1132;
  BUF_X1    g000(.A(G452), .Z(G350));
  XNOR2_X1  g001(.A(KEYINPUT64), .B(G452), .ZN(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(new_n436));
  INV_X1    g011(.A(KEYINPUT65), .ZN(new_n437));
  XNOR2_X1  g012(.A(new_n436), .B(new_n437), .ZN(G220));
  INV_X1    g013(.A(G96), .ZN(G221));
  INV_X1    g014(.A(G69), .ZN(G235));
  INV_X1    g015(.A(G120), .ZN(G236));
  INV_X1    g016(.A(G57), .ZN(G237));
  XOR2_X1   g017(.A(KEYINPUT66), .B(G108), .Z(G238));
  INV_X1    g018(.A(G2072), .ZN(new_n444));
  INV_X1    g019(.A(G2078), .ZN(new_n445));
  NOR2_X1   g020(.A1(new_n444), .A2(new_n445), .ZN(new_n446));
  NAND3_X1  g021(.A1(new_n446), .A2(G2084), .A3(G2090), .ZN(G158));
  NAND3_X1  g022(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g023(.A(G452), .Z(G391));
  AND2_X1   g024(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g025(.A1(G7), .A2(G661), .ZN(new_n451));
  XOR2_X1   g026(.A(new_n451), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g027(.A1(G7), .A2(G567), .A3(G661), .ZN(new_n453));
  XNOR2_X1  g028(.A(new_n453), .B(KEYINPUT67), .ZN(G234));
  NAND3_X1  g029(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g030(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n456));
  XOR2_X1   g031(.A(KEYINPUT68), .B(KEYINPUT2), .Z(new_n457));
  XNOR2_X1  g032(.A(new_n456), .B(new_n457), .ZN(new_n458));
  NOR4_X1   g033(.A1(G238), .A2(G237), .A3(G235), .A4(G236), .ZN(new_n459));
  XOR2_X1   g034(.A(new_n459), .B(KEYINPUT69), .Z(new_n460));
  INV_X1    g035(.A(new_n460), .ZN(new_n461));
  NOR2_X1   g036(.A1(new_n458), .A2(new_n461), .ZN(G325));
  INV_X1    g037(.A(G325), .ZN(G261));
  NAND2_X1  g038(.A1(new_n461), .A2(G567), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n458), .A2(G2106), .ZN(new_n465));
  OAI21_X1  g040(.A(new_n464), .B1(new_n465), .B2(KEYINPUT70), .ZN(new_n466));
  AOI21_X1  g041(.A(new_n466), .B1(KEYINPUT70), .B2(new_n465), .ZN(new_n467));
  XOR2_X1   g042(.A(new_n467), .B(KEYINPUT71), .Z(G319));
  INV_X1    g043(.A(G2105), .ZN(new_n469));
  INV_X1    g044(.A(KEYINPUT3), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n470), .A2(G2104), .ZN(new_n471));
  INV_X1    g046(.A(G2104), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n472), .A2(KEYINPUT3), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n471), .A2(new_n473), .ZN(new_n474));
  INV_X1    g049(.A(new_n474), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n475), .A2(G125), .ZN(new_n476));
  NAND2_X1  g051(.A1(G113), .A2(G2104), .ZN(new_n477));
  AOI21_X1  g052(.A(new_n469), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  INV_X1    g053(.A(KEYINPUT74), .ZN(new_n479));
  INV_X1    g054(.A(KEYINPUT72), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n480), .A2(new_n472), .ZN(new_n481));
  NAND2_X1  g056(.A1(KEYINPUT72), .A2(G2104), .ZN(new_n482));
  NAND3_X1  g057(.A1(new_n481), .A2(KEYINPUT3), .A3(new_n482), .ZN(new_n483));
  NAND4_X1  g058(.A1(new_n483), .A2(G137), .A3(new_n469), .A4(new_n471), .ZN(new_n484));
  INV_X1    g059(.A(KEYINPUT73), .ZN(new_n485));
  NAND2_X1  g060(.A1(new_n481), .A2(new_n482), .ZN(new_n486));
  AOI21_X1  g061(.A(new_n485), .B1(new_n486), .B2(new_n469), .ZN(new_n487));
  AND2_X1   g062(.A1(KEYINPUT72), .A2(G2104), .ZN(new_n488));
  NOR2_X1   g063(.A1(KEYINPUT72), .A2(G2104), .ZN(new_n489));
  OAI211_X1 g064(.A(new_n485), .B(new_n469), .C1(new_n488), .C2(new_n489), .ZN(new_n490));
  INV_X1    g065(.A(new_n490), .ZN(new_n491));
  NOR2_X1   g066(.A1(new_n487), .A2(new_n491), .ZN(new_n492));
  INV_X1    g067(.A(G101), .ZN(new_n493));
  OAI211_X1 g068(.A(new_n479), .B(new_n484), .C1(new_n492), .C2(new_n493), .ZN(new_n494));
  OAI21_X1  g069(.A(new_n469), .B1(new_n488), .B2(new_n489), .ZN(new_n495));
  NAND2_X1  g070(.A1(new_n495), .A2(KEYINPUT73), .ZN(new_n496));
  AOI21_X1  g071(.A(new_n493), .B1(new_n496), .B2(new_n490), .ZN(new_n497));
  INV_X1    g072(.A(new_n484), .ZN(new_n498));
  OAI21_X1  g073(.A(KEYINPUT74), .B1(new_n497), .B2(new_n498), .ZN(new_n499));
  AOI21_X1  g074(.A(new_n478), .B1(new_n494), .B2(new_n499), .ZN(G160));
  NAND2_X1  g075(.A1(new_n483), .A2(new_n471), .ZN(new_n501));
  NOR2_X1   g076(.A1(new_n501), .A2(G2105), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n502), .A2(G136), .ZN(new_n503));
  NOR2_X1   g078(.A1(new_n501), .A2(new_n469), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n504), .A2(G124), .ZN(new_n505));
  OR2_X1    g080(.A1(G100), .A2(G2105), .ZN(new_n506));
  OAI211_X1 g081(.A(new_n506), .B(G2104), .C1(G112), .C2(new_n469), .ZN(new_n507));
  NAND3_X1  g082(.A1(new_n503), .A2(new_n505), .A3(new_n507), .ZN(new_n508));
  INV_X1    g083(.A(new_n508), .ZN(G162));
  NAND4_X1  g084(.A1(new_n483), .A2(G126), .A3(G2105), .A4(new_n471), .ZN(new_n510));
  OR2_X1    g085(.A1(G102), .A2(G2105), .ZN(new_n511));
  OAI211_X1 g086(.A(new_n511), .B(G2104), .C1(G114), .C2(new_n469), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n510), .A2(new_n512), .ZN(new_n513));
  INV_X1    g088(.A(G138), .ZN(new_n514));
  NOR4_X1   g089(.A1(new_n474), .A2(KEYINPUT4), .A3(new_n514), .A4(G2105), .ZN(new_n515));
  NOR2_X1   g090(.A1(new_n514), .A2(G2105), .ZN(new_n516));
  NAND3_X1  g091(.A1(new_n483), .A2(new_n471), .A3(new_n516), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n517), .A2(KEYINPUT4), .ZN(new_n518));
  AOI21_X1  g093(.A(new_n515), .B1(new_n518), .B2(KEYINPUT75), .ZN(new_n519));
  INV_X1    g094(.A(KEYINPUT75), .ZN(new_n520));
  NAND3_X1  g095(.A1(new_n517), .A2(new_n520), .A3(KEYINPUT4), .ZN(new_n521));
  AOI21_X1  g096(.A(new_n513), .B1(new_n519), .B2(new_n521), .ZN(G164));
  INV_X1    g097(.A(G50), .ZN(new_n523));
  AND2_X1   g098(.A1(KEYINPUT6), .A2(G651), .ZN(new_n524));
  NOR2_X1   g099(.A1(KEYINPUT6), .A2(G651), .ZN(new_n525));
  OR2_X1    g100(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  NAND2_X1  g101(.A1(new_n526), .A2(G543), .ZN(new_n527));
  XNOR2_X1  g102(.A(KEYINPUT5), .B(G543), .ZN(new_n528));
  NAND2_X1  g103(.A1(new_n526), .A2(new_n528), .ZN(new_n529));
  XOR2_X1   g104(.A(KEYINPUT76), .B(G88), .Z(new_n530));
  OAI22_X1  g105(.A1(new_n523), .A2(new_n527), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  INV_X1    g106(.A(KEYINPUT77), .ZN(new_n532));
  AOI22_X1  g107(.A1(new_n528), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n533));
  INV_X1    g108(.A(G651), .ZN(new_n534));
  NOR2_X1   g109(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  OR3_X1    g110(.A1(new_n531), .A2(new_n532), .A3(new_n535), .ZN(new_n536));
  OAI21_X1  g111(.A(new_n532), .B1(new_n531), .B2(new_n535), .ZN(new_n537));
  NAND2_X1  g112(.A1(new_n536), .A2(new_n537), .ZN(G166));
  NAND3_X1  g113(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n539));
  XNOR2_X1  g114(.A(new_n539), .B(KEYINPUT7), .ZN(new_n540));
  INV_X1    g115(.A(G51), .ZN(new_n541));
  OAI21_X1  g116(.A(new_n540), .B1(new_n527), .B2(new_n541), .ZN(new_n542));
  XOR2_X1   g117(.A(KEYINPUT5), .B(G543), .Z(new_n543));
  NAND2_X1  g118(.A1(new_n526), .A2(G89), .ZN(new_n544));
  NAND2_X1  g119(.A1(G63), .A2(G651), .ZN(new_n545));
  AOI21_X1  g120(.A(new_n543), .B1(new_n544), .B2(new_n545), .ZN(new_n546));
  NOR2_X1   g121(.A1(new_n542), .A2(new_n546), .ZN(G168));
  NAND2_X1  g122(.A1(G77), .A2(G543), .ZN(new_n548));
  INV_X1    g123(.A(G64), .ZN(new_n549));
  OAI21_X1  g124(.A(new_n548), .B1(new_n543), .B2(new_n549), .ZN(new_n550));
  AOI21_X1  g125(.A(new_n534), .B1(new_n550), .B2(KEYINPUT78), .ZN(new_n551));
  OAI21_X1  g126(.A(new_n551), .B1(KEYINPUT78), .B2(new_n550), .ZN(new_n552));
  INV_X1    g127(.A(new_n527), .ZN(new_n553));
  AND2_X1   g128(.A1(new_n526), .A2(new_n528), .ZN(new_n554));
  AOI22_X1  g129(.A1(G52), .A2(new_n553), .B1(new_n554), .B2(G90), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n552), .A2(new_n555), .ZN(new_n556));
  INV_X1    g131(.A(new_n556), .ZN(G171));
  AOI22_X1  g132(.A1(new_n528), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n558));
  OR2_X1    g133(.A1(new_n558), .A2(KEYINPUT79), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n558), .A2(KEYINPUT79), .ZN(new_n560));
  NAND3_X1  g135(.A1(new_n559), .A2(G651), .A3(new_n560), .ZN(new_n561));
  AOI22_X1  g136(.A1(G43), .A2(new_n553), .B1(new_n554), .B2(G81), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  XNOR2_X1  g138(.A(new_n563), .B(KEYINPUT80), .ZN(new_n564));
  INV_X1    g139(.A(new_n564), .ZN(new_n565));
  NAND2_X1  g140(.A1(new_n565), .A2(G860), .ZN(G153));
  NAND4_X1  g141(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g142(.A1(G1), .A2(G3), .ZN(new_n568));
  XNOR2_X1  g143(.A(new_n568), .B(KEYINPUT81), .ZN(new_n569));
  XNOR2_X1  g144(.A(new_n569), .B(KEYINPUT8), .ZN(new_n570));
  NAND4_X1  g145(.A1(G319), .A2(G483), .A3(G661), .A4(new_n570), .ZN(G188));
  INV_X1    g146(.A(KEYINPUT82), .ZN(new_n572));
  NAND2_X1  g147(.A1(new_n572), .A2(G53), .ZN(new_n573));
  OR3_X1    g148(.A1(new_n527), .A2(KEYINPUT9), .A3(new_n573), .ZN(new_n574));
  OAI21_X1  g149(.A(KEYINPUT9), .B1(new_n527), .B2(new_n573), .ZN(new_n575));
  AOI22_X1  g150(.A1(new_n574), .A2(new_n575), .B1(G91), .B2(new_n554), .ZN(new_n576));
  XNOR2_X1  g151(.A(new_n528), .B(KEYINPUT83), .ZN(new_n577));
  INV_X1    g152(.A(G65), .ZN(new_n578));
  NOR2_X1   g153(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  AND2_X1   g154(.A1(G78), .A2(G543), .ZN(new_n580));
  OAI21_X1  g155(.A(G651), .B1(new_n579), .B2(new_n580), .ZN(new_n581));
  NAND2_X1  g156(.A1(new_n576), .A2(new_n581), .ZN(G299));
  XOR2_X1   g157(.A(new_n556), .B(KEYINPUT84), .Z(G301));
  INV_X1    g158(.A(G168), .ZN(G286));
  INV_X1    g159(.A(G166), .ZN(G303));
  OAI211_X1 g160(.A(G49), .B(G543), .C1(new_n524), .C2(new_n525), .ZN(new_n586));
  XOR2_X1   g161(.A(new_n586), .B(KEYINPUT85), .Z(new_n587));
  OR2_X1    g162(.A1(new_n528), .A2(G74), .ZN(new_n588));
  AOI22_X1  g163(.A1(new_n554), .A2(G87), .B1(new_n588), .B2(G651), .ZN(new_n589));
  NAND2_X1  g164(.A1(new_n587), .A2(new_n589), .ZN(G288));
  INV_X1    g165(.A(G48), .ZN(new_n591));
  INV_X1    g166(.A(G86), .ZN(new_n592));
  OAI22_X1  g167(.A1(new_n591), .A2(new_n527), .B1(new_n529), .B2(new_n592), .ZN(new_n593));
  AOI22_X1  g168(.A1(new_n528), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n594));
  NOR2_X1   g169(.A1(new_n594), .A2(new_n534), .ZN(new_n595));
  NOR2_X1   g170(.A1(new_n593), .A2(new_n595), .ZN(new_n596));
  XOR2_X1   g171(.A(new_n596), .B(KEYINPUT86), .Z(new_n597));
  INV_X1    g172(.A(new_n597), .ZN(G305));
  AOI22_X1  g173(.A1(new_n528), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n599));
  NOR2_X1   g174(.A1(new_n599), .A2(new_n534), .ZN(new_n600));
  AOI22_X1  g175(.A1(G47), .A2(new_n553), .B1(new_n554), .B2(G85), .ZN(new_n601));
  INV_X1    g176(.A(KEYINPUT87), .ZN(new_n602));
  NOR2_X1   g177(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  INV_X1    g178(.A(new_n603), .ZN(new_n604));
  NAND2_X1  g179(.A1(new_n601), .A2(new_n602), .ZN(new_n605));
  AOI21_X1  g180(.A(new_n600), .B1(new_n604), .B2(new_n605), .ZN(new_n606));
  INV_X1    g181(.A(new_n606), .ZN(G290));
  NAND2_X1  g182(.A1(new_n554), .A2(G92), .ZN(new_n608));
  XNOR2_X1  g183(.A(new_n608), .B(KEYINPUT10), .ZN(new_n609));
  AOI21_X1  g184(.A(new_n609), .B1(G54), .B2(new_n553), .ZN(new_n610));
  INV_X1    g185(.A(G66), .ZN(new_n611));
  NOR2_X1   g186(.A1(new_n577), .A2(new_n611), .ZN(new_n612));
  AND2_X1   g187(.A1(G79), .A2(G543), .ZN(new_n613));
  OAI21_X1  g188(.A(G651), .B1(new_n612), .B2(new_n613), .ZN(new_n614));
  NAND2_X1  g189(.A1(new_n610), .A2(new_n614), .ZN(new_n615));
  MUX2_X1   g190(.A(new_n615), .B(G301), .S(G868), .Z(G284));
  MUX2_X1   g191(.A(new_n615), .B(G301), .S(G868), .Z(G321));
  INV_X1    g192(.A(G868), .ZN(new_n618));
  NAND2_X1  g193(.A1(G299), .A2(new_n618), .ZN(new_n619));
  OAI21_X1  g194(.A(new_n619), .B1(new_n618), .B2(G168), .ZN(G297));
  OAI21_X1  g195(.A(new_n619), .B1(new_n618), .B2(G168), .ZN(G280));
  INV_X1    g196(.A(new_n615), .ZN(new_n622));
  INV_X1    g197(.A(G559), .ZN(new_n623));
  OAI21_X1  g198(.A(new_n622), .B1(new_n623), .B2(G860), .ZN(G148));
  NAND2_X1  g199(.A1(new_n622), .A2(new_n623), .ZN(new_n625));
  XNOR2_X1  g200(.A(new_n625), .B(KEYINPUT88), .ZN(new_n626));
  NAND2_X1  g201(.A1(new_n626), .A2(G868), .ZN(new_n627));
  OAI21_X1  g202(.A(new_n627), .B1(G868), .B2(new_n565), .ZN(G323));
  XNOR2_X1  g203(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g204(.A1(new_n496), .A2(new_n490), .ZN(new_n630));
  NAND2_X1  g205(.A1(new_n630), .A2(new_n475), .ZN(new_n631));
  XOR2_X1   g206(.A(new_n631), .B(KEYINPUT12), .Z(new_n632));
  XOR2_X1   g207(.A(new_n632), .B(KEYINPUT13), .Z(new_n633));
  INV_X1    g208(.A(G2100), .ZN(new_n634));
  OR2_X1    g209(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  NAND2_X1  g210(.A1(new_n633), .A2(new_n634), .ZN(new_n636));
  NAND2_X1  g211(.A1(new_n502), .A2(G135), .ZN(new_n637));
  NAND2_X1  g212(.A1(new_n504), .A2(G123), .ZN(new_n638));
  OR2_X1    g213(.A1(G99), .A2(G2105), .ZN(new_n639));
  OAI211_X1 g214(.A(new_n639), .B(G2104), .C1(G111), .C2(new_n469), .ZN(new_n640));
  NAND3_X1  g215(.A1(new_n637), .A2(new_n638), .A3(new_n640), .ZN(new_n641));
  XOR2_X1   g216(.A(new_n641), .B(G2096), .Z(new_n642));
  NAND3_X1  g217(.A1(new_n635), .A2(new_n636), .A3(new_n642), .ZN(G156));
  XNOR2_X1  g218(.A(G2427), .B(G2438), .ZN(new_n644));
  XNOR2_X1  g219(.A(new_n644), .B(G2430), .ZN(new_n645));
  XNOR2_X1  g220(.A(KEYINPUT15), .B(G2435), .ZN(new_n646));
  OR2_X1    g221(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  NAND2_X1  g222(.A1(new_n645), .A2(new_n646), .ZN(new_n648));
  NAND3_X1  g223(.A1(new_n647), .A2(KEYINPUT14), .A3(new_n648), .ZN(new_n649));
  XOR2_X1   g224(.A(G1341), .B(G1348), .Z(new_n650));
  XNOR2_X1  g225(.A(G2443), .B(G2446), .ZN(new_n651));
  XNOR2_X1  g226(.A(new_n650), .B(new_n651), .ZN(new_n652));
  XNOR2_X1  g227(.A(new_n649), .B(new_n652), .ZN(new_n653));
  XOR2_X1   g228(.A(G2451), .B(G2454), .Z(new_n654));
  XNOR2_X1  g229(.A(KEYINPUT89), .B(KEYINPUT16), .ZN(new_n655));
  XNOR2_X1  g230(.A(new_n654), .B(new_n655), .ZN(new_n656));
  OR2_X1    g231(.A1(new_n653), .A2(new_n656), .ZN(new_n657));
  NAND2_X1  g232(.A1(new_n653), .A2(new_n656), .ZN(new_n658));
  NAND3_X1  g233(.A1(new_n657), .A2(G14), .A3(new_n658), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n659), .B(KEYINPUT90), .ZN(G401));
  XOR2_X1   g235(.A(G2084), .B(G2090), .Z(new_n661));
  XNOR2_X1  g236(.A(G2067), .B(G2678), .ZN(new_n662));
  XNOR2_X1  g237(.A(new_n662), .B(KEYINPUT91), .ZN(new_n663));
  XOR2_X1   g238(.A(G2072), .B(G2078), .Z(new_n664));
  AOI21_X1  g239(.A(new_n661), .B1(new_n663), .B2(new_n664), .ZN(new_n665));
  XNOR2_X1  g240(.A(new_n664), .B(KEYINPUT17), .ZN(new_n666));
  OAI21_X1  g241(.A(new_n665), .B1(new_n663), .B2(new_n666), .ZN(new_n667));
  XNOR2_X1  g242(.A(new_n667), .B(KEYINPUT92), .ZN(new_n668));
  INV_X1    g243(.A(new_n661), .ZN(new_n669));
  NOR3_X1   g244(.A1(new_n663), .A2(new_n664), .A3(new_n669), .ZN(new_n670));
  XNOR2_X1  g245(.A(new_n670), .B(KEYINPUT18), .ZN(new_n671));
  NAND3_X1  g246(.A1(new_n666), .A2(new_n663), .A3(new_n661), .ZN(new_n672));
  NAND3_X1  g247(.A1(new_n668), .A2(new_n671), .A3(new_n672), .ZN(new_n673));
  XNOR2_X1  g248(.A(new_n673), .B(KEYINPUT93), .ZN(new_n674));
  XOR2_X1   g249(.A(G2096), .B(G2100), .Z(new_n675));
  XNOR2_X1  g250(.A(new_n674), .B(new_n675), .ZN(G227));
  XNOR2_X1  g251(.A(G1956), .B(G2474), .ZN(new_n677));
  XNOR2_X1  g252(.A(new_n677), .B(KEYINPUT94), .ZN(new_n678));
  XNOR2_X1  g253(.A(G1961), .B(G1966), .ZN(new_n679));
  INV_X1    g254(.A(new_n679), .ZN(new_n680));
  NAND2_X1  g255(.A1(new_n678), .A2(new_n680), .ZN(new_n681));
  XNOR2_X1  g256(.A(G1971), .B(G1976), .ZN(new_n682));
  XNOR2_X1  g257(.A(new_n682), .B(KEYINPUT19), .ZN(new_n683));
  NOR2_X1   g258(.A1(new_n681), .A2(new_n683), .ZN(new_n684));
  XOR2_X1   g259(.A(new_n684), .B(KEYINPUT20), .Z(new_n685));
  NOR2_X1   g260(.A1(new_n678), .A2(new_n680), .ZN(new_n686));
  INV_X1    g261(.A(new_n686), .ZN(new_n687));
  NAND3_X1  g262(.A1(new_n687), .A2(new_n683), .A3(new_n681), .ZN(new_n688));
  OAI211_X1 g263(.A(new_n685), .B(new_n688), .C1(new_n683), .C2(new_n687), .ZN(new_n689));
  XNOR2_X1  g264(.A(new_n689), .B(KEYINPUT95), .ZN(new_n690));
  XOR2_X1   g265(.A(G1981), .B(G1986), .Z(new_n691));
  XNOR2_X1  g266(.A(G1991), .B(G1996), .ZN(new_n692));
  XNOR2_X1  g267(.A(new_n691), .B(new_n692), .ZN(new_n693));
  XOR2_X1   g268(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n694));
  XNOR2_X1  g269(.A(new_n693), .B(new_n694), .ZN(new_n695));
  XNOR2_X1  g270(.A(new_n690), .B(new_n695), .ZN(new_n696));
  INV_X1    g271(.A(new_n696), .ZN(G229));
  INV_X1    g272(.A(G16), .ZN(new_n698));
  NAND2_X1  g273(.A1(new_n698), .A2(G4), .ZN(new_n699));
  OAI21_X1  g274(.A(new_n699), .B1(new_n622), .B2(new_n698), .ZN(new_n700));
  XNOR2_X1  g275(.A(new_n700), .B(G1348), .ZN(new_n701));
  NAND2_X1  g276(.A1(new_n698), .A2(G19), .ZN(new_n702));
  OAI21_X1  g277(.A(new_n702), .B1(new_n565), .B2(new_n698), .ZN(new_n703));
  AOI21_X1  g278(.A(new_n701), .B1(G1341), .B2(new_n703), .ZN(new_n704));
  INV_X1    g279(.A(G29), .ZN(new_n705));
  NAND2_X1  g280(.A1(new_n705), .A2(G26), .ZN(new_n706));
  XNOR2_X1  g281(.A(new_n706), .B(KEYINPUT28), .ZN(new_n707));
  NAND2_X1  g282(.A1(new_n502), .A2(G140), .ZN(new_n708));
  NAND2_X1  g283(.A1(new_n504), .A2(G128), .ZN(new_n709));
  OR2_X1    g284(.A1(G104), .A2(G2105), .ZN(new_n710));
  OAI211_X1 g285(.A(new_n710), .B(G2104), .C1(G116), .C2(new_n469), .ZN(new_n711));
  NAND3_X1  g286(.A1(new_n708), .A2(new_n709), .A3(new_n711), .ZN(new_n712));
  INV_X1    g287(.A(new_n712), .ZN(new_n713));
  OAI21_X1  g288(.A(new_n707), .B1(new_n713), .B2(new_n705), .ZN(new_n714));
  XNOR2_X1  g289(.A(new_n714), .B(KEYINPUT100), .ZN(new_n715));
  XNOR2_X1  g290(.A(new_n715), .B(G2067), .ZN(new_n716));
  OAI211_X1 g291(.A(new_n704), .B(new_n716), .C1(G1341), .C2(new_n703), .ZN(new_n717));
  XOR2_X1   g292(.A(new_n717), .B(KEYINPUT101), .Z(new_n718));
  AOI22_X1  g293(.A1(new_n475), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n719));
  NOR2_X1   g294(.A1(new_n719), .A2(new_n469), .ZN(new_n720));
  NAND3_X1  g295(.A1(new_n469), .A2(G103), .A3(G2104), .ZN(new_n721));
  XNOR2_X1  g296(.A(new_n721), .B(KEYINPUT102), .ZN(new_n722));
  XOR2_X1   g297(.A(new_n722), .B(KEYINPUT25), .Z(new_n723));
  AOI211_X1 g298(.A(new_n720), .B(new_n723), .C1(G139), .C2(new_n502), .ZN(new_n724));
  NAND2_X1  g299(.A1(new_n724), .A2(G29), .ZN(new_n725));
  OAI21_X1  g300(.A(new_n725), .B1(G29), .B2(G33), .ZN(new_n726));
  NOR2_X1   g301(.A1(new_n726), .A2(new_n444), .ZN(new_n727));
  XOR2_X1   g302(.A(new_n727), .B(KEYINPUT103), .Z(new_n728));
  NAND2_X1  g303(.A1(new_n698), .A2(G5), .ZN(new_n729));
  OAI21_X1  g304(.A(new_n729), .B1(G171), .B2(new_n698), .ZN(new_n730));
  AOI22_X1  g305(.A1(new_n726), .A2(new_n444), .B1(new_n730), .B2(G1961), .ZN(new_n731));
  OAI211_X1 g306(.A(new_n728), .B(new_n731), .C1(G1961), .C2(new_n730), .ZN(new_n732));
  NOR2_X1   g307(.A1(G168), .A2(new_n698), .ZN(new_n733));
  AOI21_X1  g308(.A(new_n733), .B1(new_n698), .B2(G21), .ZN(new_n734));
  INV_X1    g309(.A(new_n734), .ZN(new_n735));
  NOR2_X1   g310(.A1(new_n735), .A2(G1966), .ZN(new_n736));
  XNOR2_X1  g311(.A(new_n736), .B(KEYINPUT105), .ZN(new_n737));
  NAND2_X1  g312(.A1(new_n705), .A2(G35), .ZN(new_n738));
  OAI21_X1  g313(.A(new_n738), .B1(G162), .B2(new_n705), .ZN(new_n739));
  XOR2_X1   g314(.A(KEYINPUT29), .B(G2090), .Z(new_n740));
  XNOR2_X1  g315(.A(new_n739), .B(new_n740), .ZN(new_n741));
  NAND2_X1  g316(.A1(new_n698), .A2(G20), .ZN(new_n742));
  XOR2_X1   g317(.A(new_n742), .B(KEYINPUT23), .Z(new_n743));
  AOI21_X1  g318(.A(new_n743), .B1(G299), .B2(G16), .ZN(new_n744));
  XNOR2_X1  g319(.A(new_n744), .B(G1956), .ZN(new_n745));
  INV_X1    g320(.A(G28), .ZN(new_n746));
  AOI21_X1  g321(.A(G29), .B1(new_n746), .B2(KEYINPUT30), .ZN(new_n747));
  OAI21_X1  g322(.A(new_n747), .B1(KEYINPUT30), .B2(new_n746), .ZN(new_n748));
  XNOR2_X1  g323(.A(KEYINPUT31), .B(G11), .ZN(new_n749));
  XNOR2_X1  g324(.A(new_n749), .B(KEYINPUT104), .ZN(new_n750));
  OAI211_X1 g325(.A(new_n748), .B(new_n750), .C1(new_n641), .C2(new_n705), .ZN(new_n751));
  AOI21_X1  g326(.A(new_n751), .B1(new_n735), .B2(G1966), .ZN(new_n752));
  NAND4_X1  g327(.A1(new_n737), .A2(new_n741), .A3(new_n745), .A4(new_n752), .ZN(new_n753));
  INV_X1    g328(.A(KEYINPUT24), .ZN(new_n754));
  OAI21_X1  g329(.A(new_n705), .B1(new_n754), .B2(G34), .ZN(new_n755));
  AOI21_X1  g330(.A(new_n755), .B1(new_n754), .B2(G34), .ZN(new_n756));
  AOI21_X1  g331(.A(new_n756), .B1(G160), .B2(G29), .ZN(new_n757));
  OR2_X1    g332(.A1(new_n757), .A2(G2084), .ZN(new_n758));
  NOR2_X1   g333(.A1(G27), .A2(G29), .ZN(new_n759));
  AOI21_X1  g334(.A(new_n759), .B1(G164), .B2(G29), .ZN(new_n760));
  NAND2_X1  g335(.A1(new_n760), .A2(G2078), .ZN(new_n761));
  OR2_X1    g336(.A1(new_n760), .A2(G2078), .ZN(new_n762));
  NAND2_X1  g337(.A1(new_n757), .A2(G2084), .ZN(new_n763));
  NAND4_X1  g338(.A1(new_n758), .A2(new_n761), .A3(new_n762), .A4(new_n763), .ZN(new_n764));
  NAND2_X1  g339(.A1(new_n705), .A2(G32), .ZN(new_n765));
  AOI22_X1  g340(.A1(G129), .A2(new_n504), .B1(new_n502), .B2(G141), .ZN(new_n766));
  NAND3_X1  g341(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n767));
  XNOR2_X1  g342(.A(new_n767), .B(KEYINPUT26), .ZN(new_n768));
  AOI21_X1  g343(.A(new_n768), .B1(new_n630), .B2(G105), .ZN(new_n769));
  NAND2_X1  g344(.A1(new_n766), .A2(new_n769), .ZN(new_n770));
  INV_X1    g345(.A(new_n770), .ZN(new_n771));
  OAI21_X1  g346(.A(new_n765), .B1(new_n771), .B2(new_n705), .ZN(new_n772));
  XNOR2_X1  g347(.A(new_n772), .B(KEYINPUT27), .ZN(new_n773));
  INV_X1    g348(.A(G1996), .ZN(new_n774));
  XNOR2_X1  g349(.A(new_n773), .B(new_n774), .ZN(new_n775));
  NOR4_X1   g350(.A1(new_n732), .A2(new_n753), .A3(new_n764), .A4(new_n775), .ZN(new_n776));
  NAND2_X1  g351(.A1(new_n718), .A2(new_n776), .ZN(new_n777));
  INV_X1    g352(.A(KEYINPUT98), .ZN(new_n778));
  NAND2_X1  g353(.A1(new_n778), .A2(KEYINPUT36), .ZN(new_n779));
  XOR2_X1   g354(.A(new_n779), .B(KEYINPUT99), .Z(new_n780));
  NAND2_X1  g355(.A1(new_n698), .A2(G23), .ZN(new_n781));
  NAND2_X1  g356(.A1(G288), .A2(KEYINPUT96), .ZN(new_n782));
  INV_X1    g357(.A(KEYINPUT96), .ZN(new_n783));
  NAND3_X1  g358(.A1(new_n587), .A2(new_n589), .A3(new_n783), .ZN(new_n784));
  NAND2_X1  g359(.A1(new_n782), .A2(new_n784), .ZN(new_n785));
  INV_X1    g360(.A(new_n785), .ZN(new_n786));
  OAI21_X1  g361(.A(new_n781), .B1(new_n786), .B2(new_n698), .ZN(new_n787));
  XNOR2_X1  g362(.A(new_n787), .B(KEYINPUT33), .ZN(new_n788));
  INV_X1    g363(.A(G1976), .ZN(new_n789));
  OR2_X1    g364(.A1(new_n788), .A2(new_n789), .ZN(new_n790));
  NAND2_X1  g365(.A1(new_n788), .A2(new_n789), .ZN(new_n791));
  NOR2_X1   g366(.A1(G6), .A2(G16), .ZN(new_n792));
  AOI21_X1  g367(.A(new_n792), .B1(new_n597), .B2(G16), .ZN(new_n793));
  XOR2_X1   g368(.A(KEYINPUT32), .B(G1981), .Z(new_n794));
  XNOR2_X1  g369(.A(new_n793), .B(new_n794), .ZN(new_n795));
  NOR2_X1   g370(.A1(G16), .A2(G22), .ZN(new_n796));
  AOI21_X1  g371(.A(new_n796), .B1(G166), .B2(G16), .ZN(new_n797));
  INV_X1    g372(.A(G1971), .ZN(new_n798));
  XNOR2_X1  g373(.A(new_n797), .B(new_n798), .ZN(new_n799));
  NAND4_X1  g374(.A1(new_n790), .A2(new_n791), .A3(new_n795), .A4(new_n799), .ZN(new_n800));
  NAND2_X1  g375(.A1(new_n800), .A2(KEYINPUT34), .ZN(new_n801));
  XNOR2_X1  g376(.A(new_n801), .B(KEYINPUT97), .ZN(new_n802));
  OR2_X1    g377(.A1(new_n800), .A2(KEYINPUT34), .ZN(new_n803));
  NAND2_X1  g378(.A1(new_n698), .A2(G24), .ZN(new_n804));
  OAI21_X1  g379(.A(new_n804), .B1(new_n606), .B2(new_n698), .ZN(new_n805));
  XNOR2_X1  g380(.A(new_n805), .B(G1986), .ZN(new_n806));
  NAND2_X1  g381(.A1(new_n502), .A2(G131), .ZN(new_n807));
  NAND2_X1  g382(.A1(new_n504), .A2(G119), .ZN(new_n808));
  NOR2_X1   g383(.A1(new_n469), .A2(G107), .ZN(new_n809));
  OAI21_X1  g384(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n810));
  OAI211_X1 g385(.A(new_n807), .B(new_n808), .C1(new_n809), .C2(new_n810), .ZN(new_n811));
  MUX2_X1   g386(.A(G25), .B(new_n811), .S(G29), .Z(new_n812));
  XOR2_X1   g387(.A(KEYINPUT35), .B(G1991), .Z(new_n813));
  INV_X1    g388(.A(new_n813), .ZN(new_n814));
  XNOR2_X1  g389(.A(new_n812), .B(new_n814), .ZN(new_n815));
  NOR2_X1   g390(.A1(new_n806), .A2(new_n815), .ZN(new_n816));
  NAND3_X1  g391(.A1(new_n802), .A2(new_n803), .A3(new_n816), .ZN(new_n817));
  NOR2_X1   g392(.A1(new_n778), .A2(KEYINPUT36), .ZN(new_n818));
  INV_X1    g393(.A(new_n818), .ZN(new_n819));
  AOI21_X1  g394(.A(new_n780), .B1(new_n817), .B2(new_n819), .ZN(new_n820));
  INV_X1    g395(.A(new_n820), .ZN(new_n821));
  NAND3_X1  g396(.A1(new_n817), .A2(new_n819), .A3(new_n780), .ZN(new_n822));
  AOI21_X1  g397(.A(new_n777), .B1(new_n821), .B2(new_n822), .ZN(G311));
  INV_X1    g398(.A(new_n822), .ZN(new_n824));
  OAI211_X1 g399(.A(new_n718), .B(new_n776), .C1(new_n824), .C2(new_n820), .ZN(G150));
  NAND2_X1  g400(.A1(new_n554), .A2(G93), .ZN(new_n826));
  AOI22_X1  g401(.A1(new_n528), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n827));
  XOR2_X1   g402(.A(KEYINPUT106), .B(G55), .Z(new_n828));
  OAI221_X1 g403(.A(new_n826), .B1(new_n534), .B2(new_n827), .C1(new_n527), .C2(new_n828), .ZN(new_n829));
  NAND2_X1  g404(.A1(new_n564), .A2(new_n829), .ZN(new_n830));
  OAI21_X1  g405(.A(new_n830), .B1(new_n563), .B2(new_n829), .ZN(new_n831));
  XOR2_X1   g406(.A(new_n831), .B(KEYINPUT38), .Z(new_n832));
  NAND2_X1  g407(.A1(new_n622), .A2(G559), .ZN(new_n833));
  XNOR2_X1  g408(.A(new_n832), .B(new_n833), .ZN(new_n834));
  AND2_X1   g409(.A1(new_n834), .A2(KEYINPUT39), .ZN(new_n835));
  NOR2_X1   g410(.A1(new_n834), .A2(KEYINPUT39), .ZN(new_n836));
  NOR3_X1   g411(.A1(new_n835), .A2(new_n836), .A3(G860), .ZN(new_n837));
  NAND2_X1  g412(.A1(new_n829), .A2(G860), .ZN(new_n838));
  XNOR2_X1  g413(.A(new_n838), .B(KEYINPUT37), .ZN(new_n839));
  OR2_X1    g414(.A1(new_n837), .A2(new_n839), .ZN(G145));
  INV_X1    g415(.A(KEYINPUT108), .ZN(new_n841));
  NAND2_X1  g416(.A1(new_n724), .A2(new_n841), .ZN(new_n842));
  XNOR2_X1  g417(.A(new_n842), .B(new_n771), .ZN(new_n843));
  NAND2_X1  g418(.A1(new_n504), .A2(G130), .ZN(new_n844));
  NOR2_X1   g419(.A1(new_n469), .A2(G118), .ZN(new_n845));
  OAI21_X1  g420(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n846));
  OAI21_X1  g421(.A(new_n844), .B1(new_n845), .B2(new_n846), .ZN(new_n847));
  AOI21_X1  g422(.A(new_n847), .B1(G142), .B2(new_n502), .ZN(new_n848));
  XNOR2_X1  g423(.A(new_n848), .B(new_n632), .ZN(new_n849));
  XNOR2_X1  g424(.A(new_n843), .B(new_n849), .ZN(new_n850));
  XNOR2_X1  g425(.A(G164), .B(new_n712), .ZN(new_n851));
  XNOR2_X1  g426(.A(new_n851), .B(new_n811), .ZN(new_n852));
  XNOR2_X1  g427(.A(new_n850), .B(new_n852), .ZN(new_n853));
  XNOR2_X1  g428(.A(new_n641), .B(KEYINPUT107), .ZN(new_n854));
  XNOR2_X1  g429(.A(new_n854), .B(G160), .ZN(new_n855));
  XNOR2_X1  g430(.A(new_n855), .B(G162), .ZN(new_n856));
  XNOR2_X1  g431(.A(new_n853), .B(new_n856), .ZN(new_n857));
  XNOR2_X1  g432(.A(KEYINPUT109), .B(G37), .ZN(new_n858));
  NAND2_X1  g433(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  XNOR2_X1  g434(.A(new_n859), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g435(.A1(new_n829), .A2(new_n618), .ZN(new_n861));
  XNOR2_X1  g436(.A(new_n626), .B(new_n831), .ZN(new_n862));
  XNOR2_X1  g437(.A(new_n615), .B(G299), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  XNOR2_X1  g439(.A(new_n863), .B(KEYINPUT41), .ZN(new_n865));
  OAI21_X1  g440(.A(new_n864), .B1(new_n862), .B2(new_n865), .ZN(new_n866));
  XNOR2_X1  g441(.A(new_n597), .B(new_n786), .ZN(new_n867));
  XNOR2_X1  g442(.A(new_n606), .B(G166), .ZN(new_n868));
  XNOR2_X1  g443(.A(new_n867), .B(new_n868), .ZN(new_n869));
  XOR2_X1   g444(.A(new_n869), .B(KEYINPUT42), .Z(new_n870));
  XNOR2_X1  g445(.A(new_n866), .B(new_n870), .ZN(new_n871));
  OAI21_X1  g446(.A(new_n861), .B1(new_n871), .B2(new_n618), .ZN(G295));
  OAI21_X1  g447(.A(new_n861), .B1(new_n871), .B2(new_n618), .ZN(G331));
  XNOR2_X1  g448(.A(KEYINPUT110), .B(KEYINPUT44), .ZN(new_n874));
  INV_X1    g449(.A(new_n858), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n556), .A2(G286), .ZN(new_n876));
  OAI21_X1  g451(.A(new_n876), .B1(G301), .B2(G286), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n831), .A2(new_n877), .ZN(new_n878));
  XNOR2_X1  g453(.A(new_n878), .B(KEYINPUT111), .ZN(new_n879));
  NOR2_X1   g454(.A1(new_n831), .A2(new_n877), .ZN(new_n880));
  INV_X1    g455(.A(new_n880), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n879), .A2(new_n881), .ZN(new_n882));
  NOR2_X1   g457(.A1(new_n880), .A2(new_n863), .ZN(new_n883));
  AOI22_X1  g458(.A1(new_n882), .A2(new_n865), .B1(new_n878), .B2(new_n883), .ZN(new_n884));
  AOI21_X1  g459(.A(new_n875), .B1(new_n884), .B2(new_n869), .ZN(new_n885));
  INV_X1    g460(.A(KEYINPUT43), .ZN(new_n886));
  INV_X1    g461(.A(new_n869), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n879), .A2(new_n883), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n881), .A2(new_n878), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n889), .A2(new_n865), .ZN(new_n890));
  OAI21_X1  g465(.A(new_n888), .B1(KEYINPUT112), .B2(new_n890), .ZN(new_n891));
  AND2_X1   g466(.A1(new_n890), .A2(KEYINPUT112), .ZN(new_n892));
  OAI21_X1  g467(.A(new_n887), .B1(new_n891), .B2(new_n892), .ZN(new_n893));
  NAND3_X1  g468(.A1(new_n885), .A2(new_n886), .A3(new_n893), .ZN(new_n894));
  AND2_X1   g469(.A1(new_n894), .A2(KEYINPUT113), .ZN(new_n895));
  INV_X1    g470(.A(G37), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n883), .A2(new_n878), .ZN(new_n897));
  INV_X1    g472(.A(KEYINPUT111), .ZN(new_n898));
  XNOR2_X1  g473(.A(new_n878), .B(new_n898), .ZN(new_n899));
  NOR2_X1   g474(.A1(new_n899), .A2(new_n880), .ZN(new_n900));
  INV_X1    g475(.A(new_n865), .ZN(new_n901));
  OAI21_X1  g476(.A(new_n897), .B1(new_n900), .B2(new_n901), .ZN(new_n902));
  OAI21_X1  g477(.A(new_n896), .B1(new_n902), .B2(new_n887), .ZN(new_n903));
  NOR2_X1   g478(.A1(new_n884), .A2(new_n869), .ZN(new_n904));
  OAI21_X1  g479(.A(KEYINPUT43), .B1(new_n903), .B2(new_n904), .ZN(new_n905));
  INV_X1    g480(.A(KEYINPUT113), .ZN(new_n906));
  NAND4_X1  g481(.A1(new_n885), .A2(new_n893), .A3(new_n906), .A4(new_n886), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n905), .A2(new_n907), .ZN(new_n908));
  OAI21_X1  g483(.A(new_n874), .B1(new_n895), .B2(new_n908), .ZN(new_n909));
  INV_X1    g484(.A(KEYINPUT44), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n885), .A2(new_n893), .ZN(new_n911));
  AOI21_X1  g486(.A(new_n910), .B1(new_n911), .B2(KEYINPUT43), .ZN(new_n912));
  NOR2_X1   g487(.A1(new_n903), .A2(new_n904), .ZN(new_n913));
  AOI21_X1  g488(.A(KEYINPUT114), .B1(new_n913), .B2(new_n886), .ZN(new_n914));
  INV_X1    g489(.A(KEYINPUT114), .ZN(new_n915));
  NOR4_X1   g490(.A1(new_n903), .A2(new_n904), .A3(new_n915), .A4(KEYINPUT43), .ZN(new_n916));
  OAI21_X1  g491(.A(new_n912), .B1(new_n914), .B2(new_n916), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n909), .A2(new_n917), .ZN(G397));
  XOR2_X1   g493(.A(new_n712), .B(G2067), .Z(new_n919));
  XNOR2_X1  g494(.A(new_n919), .B(KEYINPUT116), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n920), .A2(new_n771), .ZN(new_n921));
  INV_X1    g496(.A(KEYINPUT45), .ZN(new_n922));
  OAI21_X1  g497(.A(new_n922), .B1(G164), .B2(G1384), .ZN(new_n923));
  INV_X1    g498(.A(new_n923), .ZN(new_n924));
  INV_X1    g499(.A(G40), .ZN(new_n925));
  AOI211_X1 g500(.A(new_n925), .B(new_n478), .C1(new_n494), .C2(new_n499), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n924), .A2(new_n926), .ZN(new_n927));
  INV_X1    g502(.A(new_n927), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n921), .A2(new_n928), .ZN(new_n929));
  AOI21_X1  g504(.A(new_n929), .B1(new_n774), .B2(new_n920), .ZN(new_n930));
  NOR2_X1   g505(.A1(new_n927), .A2(G1996), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n931), .A2(new_n771), .ZN(new_n932));
  XNOR2_X1  g507(.A(new_n932), .B(KEYINPUT115), .ZN(new_n933));
  NOR2_X1   g508(.A1(new_n930), .A2(new_n933), .ZN(new_n934));
  AND2_X1   g509(.A1(new_n811), .A2(new_n814), .ZN(new_n935));
  NOR2_X1   g510(.A1(new_n811), .A2(new_n814), .ZN(new_n936));
  OAI21_X1  g511(.A(new_n928), .B1(new_n935), .B2(new_n936), .ZN(new_n937));
  AND2_X1   g512(.A1(new_n934), .A2(new_n937), .ZN(new_n938));
  XOR2_X1   g513(.A(new_n606), .B(G1986), .Z(new_n939));
  NAND2_X1  g514(.A1(new_n939), .A2(new_n928), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n938), .A2(new_n940), .ZN(new_n941));
  INV_X1    g516(.A(KEYINPUT63), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n518), .A2(KEYINPUT75), .ZN(new_n943));
  INV_X1    g518(.A(new_n515), .ZN(new_n944));
  NAND3_X1  g519(.A1(new_n943), .A2(new_n521), .A3(new_n944), .ZN(new_n945));
  INV_X1    g520(.A(new_n513), .ZN(new_n946));
  AOI21_X1  g521(.A(G1384), .B1(new_n945), .B2(new_n946), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n926), .A2(new_n947), .ZN(new_n948));
  NAND3_X1  g523(.A1(new_n782), .A2(G1976), .A3(new_n784), .ZN(new_n949));
  NAND3_X1  g524(.A1(new_n948), .A2(G8), .A3(new_n949), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n950), .A2(KEYINPUT52), .ZN(new_n951));
  INV_X1    g526(.A(G8), .ZN(new_n952));
  AOI21_X1  g527(.A(new_n952), .B1(new_n926), .B2(new_n947), .ZN(new_n953));
  AOI21_X1  g528(.A(KEYINPUT52), .B1(G288), .B2(new_n789), .ZN(new_n954));
  NAND3_X1  g529(.A1(new_n953), .A2(new_n949), .A3(new_n954), .ZN(new_n955));
  INV_X1    g530(.A(G1981), .ZN(new_n956));
  NOR2_X1   g531(.A1(new_n596), .A2(new_n956), .ZN(new_n957));
  INV_X1    g532(.A(KEYINPUT49), .ZN(new_n958));
  NOR3_X1   g533(.A1(new_n593), .A2(G1981), .A3(new_n595), .ZN(new_n959));
  OR3_X1    g534(.A1(new_n957), .A2(new_n958), .A3(new_n959), .ZN(new_n960));
  OAI21_X1  g535(.A(new_n958), .B1(new_n957), .B2(new_n959), .ZN(new_n961));
  NAND3_X1  g536(.A1(new_n953), .A2(new_n960), .A3(new_n961), .ZN(new_n962));
  NAND3_X1  g537(.A1(new_n951), .A2(new_n955), .A3(new_n962), .ZN(new_n963));
  INV_X1    g538(.A(G1384), .ZN(new_n964));
  AND3_X1   g539(.A1(new_n517), .A2(new_n520), .A3(KEYINPUT4), .ZN(new_n965));
  AOI21_X1  g540(.A(new_n520), .B1(new_n517), .B2(KEYINPUT4), .ZN(new_n966));
  NOR3_X1   g541(.A1(new_n965), .A2(new_n966), .A3(new_n515), .ZN(new_n967));
  OAI211_X1 g542(.A(KEYINPUT45), .B(new_n964), .C1(new_n967), .C2(new_n513), .ZN(new_n968));
  NAND3_X1  g543(.A1(new_n923), .A2(new_n926), .A3(new_n968), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n969), .A2(new_n798), .ZN(new_n970));
  XOR2_X1   g545(.A(KEYINPUT118), .B(KEYINPUT50), .Z(new_n971));
  INV_X1    g546(.A(new_n971), .ZN(new_n972));
  OAI21_X1  g547(.A(new_n972), .B1(G164), .B2(G1384), .ZN(new_n973));
  OAI21_X1  g548(.A(new_n964), .B1(new_n967), .B2(new_n513), .ZN(new_n974));
  OAI211_X1 g549(.A(new_n973), .B(new_n926), .C1(new_n974), .C2(KEYINPUT50), .ZN(new_n975));
  OAI21_X1  g550(.A(new_n970), .B1(G2090), .B2(new_n975), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n976), .A2(G8), .ZN(new_n977));
  NAND2_X1  g552(.A1(G303), .A2(G8), .ZN(new_n978));
  XNOR2_X1  g553(.A(new_n978), .B(KEYINPUT55), .ZN(new_n979));
  AOI21_X1  g554(.A(new_n963), .B1(new_n977), .B2(new_n979), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n970), .A2(KEYINPUT117), .ZN(new_n981));
  INV_X1    g556(.A(KEYINPUT117), .ZN(new_n982));
  NAND3_X1  g557(.A1(new_n969), .A2(new_n982), .A3(new_n798), .ZN(new_n983));
  INV_X1    g558(.A(new_n478), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n630), .A2(G101), .ZN(new_n985));
  AOI21_X1  g560(.A(new_n479), .B1(new_n985), .B2(new_n484), .ZN(new_n986));
  NOR3_X1   g561(.A1(new_n497), .A2(new_n498), .A3(KEYINPUT74), .ZN(new_n987));
  OAI211_X1 g562(.A(G40), .B(new_n984), .C1(new_n986), .C2(new_n987), .ZN(new_n988));
  AOI21_X1  g563(.A(new_n988), .B1(new_n947), .B2(new_n971), .ZN(new_n989));
  INV_X1    g564(.A(G2090), .ZN(new_n990));
  OAI211_X1 g565(.A(KEYINPUT119), .B(KEYINPUT50), .C1(G164), .C2(G1384), .ZN(new_n991));
  INV_X1    g566(.A(KEYINPUT119), .ZN(new_n992));
  INV_X1    g567(.A(KEYINPUT50), .ZN(new_n993));
  OAI21_X1  g568(.A(new_n992), .B1(new_n947), .B2(new_n993), .ZN(new_n994));
  NAND4_X1  g569(.A1(new_n989), .A2(new_n990), .A3(new_n991), .A4(new_n994), .ZN(new_n995));
  NAND3_X1  g570(.A1(new_n981), .A2(new_n983), .A3(new_n995), .ZN(new_n996));
  INV_X1    g571(.A(KEYINPUT55), .ZN(new_n997));
  XNOR2_X1  g572(.A(new_n978), .B(new_n997), .ZN(new_n998));
  NAND3_X1  g573(.A1(new_n996), .A2(G8), .A3(new_n998), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n980), .A2(new_n999), .ZN(new_n1000));
  INV_X1    g575(.A(G2084), .ZN(new_n1001));
  NAND4_X1  g576(.A1(new_n989), .A2(new_n1001), .A3(new_n991), .A4(new_n994), .ZN(new_n1002));
  INV_X1    g577(.A(G1966), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n969), .A2(new_n1003), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n1002), .A2(new_n1004), .ZN(new_n1005));
  NOR2_X1   g580(.A1(G286), .A2(new_n952), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n1005), .A2(new_n1006), .ZN(new_n1007));
  OAI21_X1  g582(.A(new_n942), .B1(new_n1000), .B2(new_n1007), .ZN(new_n1008));
  AOI21_X1  g583(.A(new_n998), .B1(new_n996), .B2(G8), .ZN(new_n1009));
  OAI21_X1  g584(.A(KEYINPUT121), .B1(new_n1009), .B2(new_n963), .ZN(new_n1010));
  AND3_X1   g585(.A1(new_n1005), .A2(KEYINPUT63), .A3(new_n1006), .ZN(new_n1011));
  AND2_X1   g586(.A1(new_n999), .A2(new_n1011), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n1010), .A2(new_n1012), .ZN(new_n1013));
  NOR3_X1   g588(.A1(new_n1009), .A2(KEYINPUT121), .A3(new_n963), .ZN(new_n1014));
  OAI21_X1  g589(.A(new_n1008), .B1(new_n1013), .B2(new_n1014), .ZN(new_n1015));
  AND4_X1   g590(.A1(new_n789), .A2(new_n962), .A3(new_n587), .A4(new_n589), .ZN(new_n1016));
  OAI21_X1  g591(.A(new_n953), .B1(new_n1016), .B2(new_n959), .ZN(new_n1017));
  OAI21_X1  g592(.A(new_n1017), .B1(new_n999), .B2(new_n963), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n1018), .A2(KEYINPUT120), .ZN(new_n1019));
  INV_X1    g594(.A(KEYINPUT120), .ZN(new_n1020));
  OAI211_X1 g595(.A(new_n1017), .B(new_n1020), .C1(new_n999), .C2(new_n963), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n1019), .A2(new_n1021), .ZN(new_n1022));
  AOI21_X1  g597(.A(KEYINPUT122), .B1(new_n1015), .B2(new_n1022), .ZN(new_n1023));
  NAND3_X1  g598(.A1(new_n1002), .A2(G168), .A3(new_n1004), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n1024), .A2(G8), .ZN(new_n1025));
  AOI21_X1  g600(.A(G168), .B1(new_n1002), .B2(new_n1004), .ZN(new_n1026));
  OAI21_X1  g601(.A(KEYINPUT51), .B1(new_n1025), .B2(new_n1026), .ZN(new_n1027));
  INV_X1    g602(.A(KEYINPUT51), .ZN(new_n1028));
  NAND3_X1  g603(.A1(new_n1024), .A2(new_n1028), .A3(G8), .ZN(new_n1029));
  NAND2_X1  g604(.A1(new_n1027), .A2(new_n1029), .ZN(new_n1030));
  NAND2_X1  g605(.A1(new_n1030), .A2(KEYINPUT62), .ZN(new_n1031));
  INV_X1    g606(.A(KEYINPUT62), .ZN(new_n1032));
  NAND3_X1  g607(.A1(new_n1027), .A2(new_n1032), .A3(new_n1029), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n947), .A2(new_n971), .ZN(new_n1034));
  NAND4_X1  g609(.A1(new_n994), .A2(new_n926), .A3(new_n991), .A4(new_n1034), .ZN(new_n1035));
  INV_X1    g610(.A(G1961), .ZN(new_n1036));
  INV_X1    g611(.A(KEYINPUT53), .ZN(new_n1037));
  NAND4_X1  g612(.A1(new_n923), .A2(new_n926), .A3(new_n968), .A4(new_n445), .ZN(new_n1038));
  AOI22_X1  g613(.A1(new_n1035), .A2(new_n1036), .B1(new_n1037), .B2(new_n1038), .ZN(new_n1039));
  OR2_X1    g614(.A1(new_n1038), .A2(new_n1037), .ZN(new_n1040));
  AOI21_X1  g615(.A(G301), .B1(new_n1039), .B2(new_n1040), .ZN(new_n1041));
  AND3_X1   g616(.A1(new_n980), .A2(new_n999), .A3(new_n1041), .ZN(new_n1042));
  NAND3_X1  g617(.A1(new_n1031), .A2(new_n1033), .A3(new_n1042), .ZN(new_n1043));
  NAND4_X1  g618(.A1(new_n923), .A2(new_n926), .A3(new_n968), .A4(new_n774), .ZN(new_n1044));
  XOR2_X1   g619(.A(KEYINPUT58), .B(G1341), .Z(new_n1045));
  OAI21_X1  g620(.A(new_n1045), .B1(new_n974), .B2(new_n988), .ZN(new_n1046));
  AOI21_X1  g621(.A(new_n564), .B1(new_n1044), .B2(new_n1046), .ZN(new_n1047));
  AOI21_X1  g622(.A(KEYINPUT124), .B1(new_n1047), .B2(KEYINPUT125), .ZN(new_n1048));
  INV_X1    g623(.A(KEYINPUT59), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n1048), .A2(new_n1049), .ZN(new_n1050));
  NAND2_X1  g625(.A1(new_n1047), .A2(KEYINPUT124), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n1051), .A2(KEYINPUT59), .ZN(new_n1052));
  OAI21_X1  g627(.A(new_n1050), .B1(new_n1052), .B2(new_n1048), .ZN(new_n1053));
  NOR3_X1   g628(.A1(new_n974), .A2(new_n988), .A3(G2067), .ZN(new_n1054));
  INV_X1    g629(.A(G1348), .ZN(new_n1055));
  AOI21_X1  g630(.A(new_n1054), .B1(new_n1035), .B2(new_n1055), .ZN(new_n1056));
  NOR2_X1   g631(.A1(new_n1056), .A2(KEYINPUT60), .ZN(new_n1057));
  INV_X1    g632(.A(KEYINPUT60), .ZN(new_n1058));
  AOI211_X1 g633(.A(new_n1058), .B(new_n1054), .C1(new_n1035), .C2(new_n1055), .ZN(new_n1059));
  NOR3_X1   g634(.A1(new_n1057), .A2(new_n1059), .A3(new_n615), .ZN(new_n1060));
  NOR2_X1   g635(.A1(new_n1053), .A2(new_n1060), .ZN(new_n1061));
  INV_X1    g636(.A(KEYINPUT61), .ZN(new_n1062));
  INV_X1    g637(.A(G1956), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n975), .A2(new_n1063), .ZN(new_n1064));
  XOR2_X1   g639(.A(G299), .B(KEYINPUT57), .Z(new_n1065));
  XNOR2_X1  g640(.A(KEYINPUT56), .B(G2072), .ZN(new_n1066));
  NAND4_X1  g641(.A1(new_n923), .A2(new_n926), .A3(new_n968), .A4(new_n1066), .ZN(new_n1067));
  NAND3_X1  g642(.A1(new_n1064), .A2(new_n1065), .A3(new_n1067), .ZN(new_n1068));
  INV_X1    g643(.A(new_n1068), .ZN(new_n1069));
  AOI21_X1  g644(.A(new_n1065), .B1(new_n1064), .B2(new_n1067), .ZN(new_n1070));
  OAI21_X1  g645(.A(new_n1062), .B1(new_n1069), .B2(new_n1070), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n1064), .A2(new_n1067), .ZN(new_n1072));
  INV_X1    g647(.A(new_n1065), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n1072), .A2(new_n1073), .ZN(new_n1074));
  NAND3_X1  g649(.A1(new_n1074), .A2(KEYINPUT61), .A3(new_n1068), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n1059), .A2(new_n615), .ZN(new_n1076));
  AND3_X1   g651(.A1(new_n1071), .A2(new_n1075), .A3(new_n1076), .ZN(new_n1077));
  INV_X1    g652(.A(new_n1056), .ZN(new_n1078));
  NAND3_X1  g653(.A1(new_n1078), .A2(KEYINPUT123), .A3(new_n622), .ZN(new_n1079));
  INV_X1    g654(.A(KEYINPUT123), .ZN(new_n1080));
  OAI21_X1  g655(.A(new_n1080), .B1(new_n1056), .B2(new_n615), .ZN(new_n1081));
  NAND3_X1  g656(.A1(new_n1079), .A2(new_n1081), .A3(new_n1074), .ZN(new_n1082));
  AOI22_X1  g657(.A1(new_n1061), .A2(new_n1077), .B1(new_n1068), .B2(new_n1082), .ZN(new_n1083));
  INV_X1    g658(.A(new_n1000), .ZN(new_n1084));
  INV_X1    g659(.A(KEYINPUT54), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n1039), .A2(new_n1040), .ZN(new_n1086));
  INV_X1    g661(.A(G301), .ZN(new_n1087));
  NOR2_X1   g662(.A1(new_n1086), .A2(new_n1087), .ZN(new_n1088));
  OAI21_X1  g663(.A(new_n1085), .B1(new_n1088), .B2(new_n1041), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n1086), .A2(G171), .ZN(new_n1090));
  OAI211_X1 g665(.A(new_n1090), .B(KEYINPUT54), .C1(new_n1087), .C2(new_n1086), .ZN(new_n1091));
  NAND4_X1  g666(.A1(new_n1084), .A2(new_n1089), .A3(new_n1091), .A4(new_n1030), .ZN(new_n1092));
  OAI21_X1  g667(.A(new_n1043), .B1(new_n1083), .B2(new_n1092), .ZN(new_n1093));
  NOR2_X1   g668(.A1(new_n1023), .A2(new_n1093), .ZN(new_n1094));
  INV_X1    g669(.A(KEYINPUT121), .ZN(new_n1095));
  INV_X1    g670(.A(new_n963), .ZN(new_n1096));
  AND2_X1   g671(.A1(new_n996), .A2(G8), .ZN(new_n1097));
  OAI211_X1 g672(.A(new_n1095), .B(new_n1096), .C1(new_n1097), .C2(new_n998), .ZN(new_n1098));
  NAND3_X1  g673(.A1(new_n1098), .A2(new_n1010), .A3(new_n1012), .ZN(new_n1099));
  AOI22_X1  g674(.A1(new_n1099), .A2(new_n1008), .B1(new_n1019), .B2(new_n1021), .ZN(new_n1100));
  NAND2_X1  g675(.A1(new_n1100), .A2(KEYINPUT122), .ZN(new_n1101));
  AOI21_X1  g676(.A(new_n941), .B1(new_n1094), .B2(new_n1101), .ZN(new_n1102));
  NOR3_X1   g677(.A1(new_n927), .A2(G290), .A3(G1986), .ZN(new_n1103));
  XOR2_X1   g678(.A(new_n1103), .B(KEYINPUT48), .Z(new_n1104));
  NAND2_X1  g679(.A1(new_n938), .A2(new_n1104), .ZN(new_n1105));
  XOR2_X1   g680(.A(new_n931), .B(KEYINPUT46), .Z(new_n1106));
  NAND2_X1  g681(.A1(new_n1106), .A2(new_n929), .ZN(new_n1107));
  XNOR2_X1  g682(.A(new_n1107), .B(KEYINPUT47), .ZN(new_n1108));
  NAND2_X1  g683(.A1(new_n1105), .A2(new_n1108), .ZN(new_n1109));
  INV_X1    g684(.A(G2067), .ZN(new_n1110));
  AOI22_X1  g685(.A1(new_n934), .A2(new_n936), .B1(new_n1110), .B2(new_n713), .ZN(new_n1111));
  NOR2_X1   g686(.A1(new_n1111), .A2(new_n927), .ZN(new_n1112));
  OR2_X1    g687(.A1(new_n1109), .A2(new_n1112), .ZN(new_n1113));
  OAI21_X1  g688(.A(KEYINPUT126), .B1(new_n1102), .B2(new_n1113), .ZN(new_n1114));
  INV_X1    g689(.A(new_n941), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n1082), .A2(new_n1068), .ZN(new_n1116));
  OAI21_X1  g691(.A(new_n622), .B1(new_n1078), .B2(new_n1058), .ZN(new_n1117));
  OAI221_X1 g692(.A(new_n1050), .B1(new_n1052), .B2(new_n1048), .C1(new_n1117), .C2(new_n1057), .ZN(new_n1118));
  NAND3_X1  g693(.A1(new_n1071), .A2(new_n1075), .A3(new_n1076), .ZN(new_n1119));
  OAI21_X1  g694(.A(new_n1116), .B1(new_n1118), .B2(new_n1119), .ZN(new_n1120));
  AND3_X1   g695(.A1(new_n1084), .A2(new_n1089), .A3(new_n1091), .ZN(new_n1121));
  NAND3_X1  g696(.A1(new_n1120), .A2(new_n1121), .A3(new_n1030), .ZN(new_n1122));
  OAI211_X1 g697(.A(new_n1122), .B(new_n1043), .C1(new_n1100), .C2(KEYINPUT122), .ZN(new_n1123));
  INV_X1    g698(.A(new_n1101), .ZN(new_n1124));
  OAI21_X1  g699(.A(new_n1115), .B1(new_n1123), .B2(new_n1124), .ZN(new_n1125));
  INV_X1    g700(.A(KEYINPUT126), .ZN(new_n1126));
  NOR2_X1   g701(.A1(new_n1109), .A2(new_n1112), .ZN(new_n1127));
  NAND3_X1  g702(.A1(new_n1125), .A2(new_n1126), .A3(new_n1127), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n1114), .A2(new_n1128), .ZN(G329));
  assign    G231 = 1'b0;
  NAND2_X1  g704(.A1(new_n467), .A2(new_n659), .ZN(new_n1131));
  NOR3_X1   g705(.A1(G229), .A2(G227), .A3(new_n1131), .ZN(new_n1132));
  OAI211_X1 g706(.A(new_n859), .B(new_n1132), .C1(new_n895), .C2(new_n908), .ZN(G225));
  INV_X1    g707(.A(G225), .ZN(G308));
endmodule


