//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 1 1 1 0 1 0 1 1 0 0 1 0 0 1 1 1 1 1 0 0 1 1 0 1 1 1 1 1 1 1 1 0 0 1 1 0 1 0 0 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 1 0 1 1 1 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:28:55 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n447, new_n451, new_n452, new_n453, new_n454, new_n457,
    new_n458, new_n459, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n527, new_n528, new_n529, new_n530, new_n531, new_n532,
    new_n533, new_n534, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n543, new_n544, new_n545, new_n546, new_n547, new_n548, new_n550,
    new_n552, new_n553, new_n555, new_n556, new_n557, new_n558, new_n559,
    new_n560, new_n561, new_n562, new_n563, new_n567, new_n568, new_n569,
    new_n570, new_n572, new_n573, new_n574, new_n575, new_n576, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n595,
    new_n596, new_n599, new_n601, new_n602, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n618, new_n619, new_n620, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n808,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n825, new_n826, new_n827, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n896, new_n897, new_n898,
    new_n899, new_n900, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1113, new_n1114, new_n1115, new_n1116, new_n1117, new_n1118,
    new_n1119;
  XOR2_X1   g000(.A(KEYINPUT64), .B(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  XNOR2_X1  g007(.A(KEYINPUT65), .B(G2066), .ZN(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  XOR2_X1   g009(.A(KEYINPUT66), .B(G132), .Z(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT67), .Z(new_n447));
  XNOR2_X1  g022(.A(new_n447), .B(KEYINPUT1), .ZN(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G219), .A2(G220), .A3(G218), .A4(G221), .ZN(new_n451));
  XNOR2_X1  g026(.A(new_n451), .B(KEYINPUT68), .ZN(new_n452));
  XOR2_X1   g027(.A(new_n452), .B(KEYINPUT2), .Z(new_n453));
  NAND4_X1  g028(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n454));
  NOR2_X1   g029(.A1(new_n453), .A2(new_n454), .ZN(G325));
  INV_X1    g030(.A(G325), .ZN(G261));
  NAND2_X1  g031(.A1(new_n453), .A2(G2106), .ZN(new_n457));
  NAND2_X1  g032(.A1(new_n454), .A2(G567), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  INV_X1    g034(.A(new_n459), .ZN(G319));
  INV_X1    g035(.A(G2104), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n461), .A2(KEYINPUT3), .ZN(new_n462));
  INV_X1    g037(.A(KEYINPUT3), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n463), .A2(G2104), .ZN(new_n464));
  NAND3_X1  g039(.A1(new_n462), .A2(new_n464), .A3(G125), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n465), .A2(KEYINPUT69), .ZN(new_n466));
  XNOR2_X1  g041(.A(KEYINPUT3), .B(G2104), .ZN(new_n467));
  INV_X1    g042(.A(KEYINPUT69), .ZN(new_n468));
  NAND3_X1  g043(.A1(new_n467), .A2(new_n468), .A3(G125), .ZN(new_n469));
  NAND3_X1  g044(.A1(KEYINPUT70), .A2(G113), .A3(G2104), .ZN(new_n470));
  INV_X1    g045(.A(KEYINPUT70), .ZN(new_n471));
  INV_X1    g046(.A(G113), .ZN(new_n472));
  OAI21_X1  g047(.A(new_n471), .B1(new_n472), .B2(new_n461), .ZN(new_n473));
  NAND4_X1  g048(.A1(new_n466), .A2(new_n469), .A3(new_n470), .A4(new_n473), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n474), .A2(G2105), .ZN(new_n475));
  INV_X1    g050(.A(G2105), .ZN(new_n476));
  AND3_X1   g051(.A1(new_n476), .A2(G101), .A3(G2104), .ZN(new_n477));
  NAND3_X1  g052(.A1(new_n467), .A2(G137), .A3(new_n476), .ZN(new_n478));
  INV_X1    g053(.A(KEYINPUT71), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  NAND4_X1  g055(.A1(new_n467), .A2(KEYINPUT71), .A3(G137), .A4(new_n476), .ZN(new_n481));
  AOI21_X1  g056(.A(new_n477), .B1(new_n480), .B2(new_n481), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n475), .A2(new_n482), .ZN(new_n483));
  INV_X1    g058(.A(new_n483), .ZN(G160));
  NAND2_X1  g059(.A1(new_n462), .A2(new_n464), .ZN(new_n485));
  NOR2_X1   g060(.A1(new_n485), .A2(new_n476), .ZN(new_n486));
  NAND2_X1  g061(.A1(new_n486), .A2(G124), .ZN(new_n487));
  NOR2_X1   g062(.A1(new_n485), .A2(G2105), .ZN(new_n488));
  NAND2_X1  g063(.A1(new_n488), .A2(G136), .ZN(new_n489));
  OR2_X1    g064(.A1(G100), .A2(G2105), .ZN(new_n490));
  OAI211_X1 g065(.A(new_n490), .B(G2104), .C1(G112), .C2(new_n476), .ZN(new_n491));
  NAND3_X1  g066(.A1(new_n487), .A2(new_n489), .A3(new_n491), .ZN(new_n492));
  INV_X1    g067(.A(new_n492), .ZN(G162));
  NAND2_X1  g068(.A1(new_n476), .A2(G2104), .ZN(new_n494));
  INV_X1    g069(.A(G102), .ZN(new_n495));
  NOR2_X1   g070(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  NAND2_X1  g071(.A1(G114), .A2(G2104), .ZN(new_n497));
  INV_X1    g072(.A(G126), .ZN(new_n498));
  OAI21_X1  g073(.A(new_n497), .B1(new_n485), .B2(new_n498), .ZN(new_n499));
  AOI21_X1  g074(.A(new_n496), .B1(new_n499), .B2(G2105), .ZN(new_n500));
  NAND4_X1  g075(.A1(new_n462), .A2(new_n464), .A3(G138), .A4(new_n476), .ZN(new_n501));
  NAND2_X1  g076(.A1(new_n501), .A2(KEYINPUT4), .ZN(new_n502));
  INV_X1    g077(.A(KEYINPUT4), .ZN(new_n503));
  NAND4_X1  g078(.A1(new_n467), .A2(new_n503), .A3(G138), .A4(new_n476), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n502), .A2(new_n504), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n500), .A2(new_n505), .ZN(new_n506));
  INV_X1    g081(.A(new_n506), .ZN(G164));
  INV_X1    g082(.A(KEYINPUT5), .ZN(new_n508));
  INV_X1    g083(.A(KEYINPUT72), .ZN(new_n509));
  INV_X1    g084(.A(G543), .ZN(new_n510));
  OAI21_X1  g085(.A(new_n508), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  NAND3_X1  g086(.A1(KEYINPUT72), .A2(KEYINPUT5), .A3(G543), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  AOI22_X1  g088(.A1(new_n513), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n514));
  INV_X1    g089(.A(G651), .ZN(new_n515));
  NOR2_X1   g090(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n515), .A2(KEYINPUT6), .ZN(new_n517));
  INV_X1    g092(.A(KEYINPUT6), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n518), .A2(G651), .ZN(new_n519));
  AND3_X1   g094(.A1(new_n517), .A2(new_n519), .A3(G543), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n520), .A2(G50), .ZN(new_n521));
  AND2_X1   g096(.A1(new_n517), .A2(new_n519), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n513), .A2(new_n522), .ZN(new_n523));
  INV_X1    g098(.A(G88), .ZN(new_n524));
  OAI21_X1  g099(.A(new_n521), .B1(new_n523), .B2(new_n524), .ZN(new_n525));
  NOR2_X1   g100(.A1(new_n516), .A2(new_n525), .ZN(G166));
  NAND3_X1  g101(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n527));
  XNOR2_X1  g102(.A(new_n527), .B(KEYINPUT73), .ZN(new_n528));
  XOR2_X1   g103(.A(new_n528), .B(KEYINPUT7), .Z(new_n529));
  NAND2_X1  g104(.A1(new_n520), .A2(G51), .ZN(new_n530));
  AOI22_X1  g105(.A1(new_n522), .A2(G89), .B1(G63), .B2(G651), .ZN(new_n531));
  INV_X1    g106(.A(new_n513), .ZN(new_n532));
  OAI21_X1  g107(.A(new_n530), .B1(new_n531), .B2(new_n532), .ZN(new_n533));
  NOR2_X1   g108(.A1(new_n529), .A2(new_n533), .ZN(new_n534));
  XNOR2_X1  g109(.A(new_n534), .B(KEYINPUT74), .ZN(G286));
  INV_X1    g110(.A(G286), .ZN(G168));
  AOI22_X1  g111(.A1(new_n513), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n537));
  NOR2_X1   g112(.A1(new_n537), .A2(new_n515), .ZN(new_n538));
  NAND2_X1  g113(.A1(new_n520), .A2(G52), .ZN(new_n539));
  INV_X1    g114(.A(G90), .ZN(new_n540));
  OAI21_X1  g115(.A(new_n539), .B1(new_n523), .B2(new_n540), .ZN(new_n541));
  NOR2_X1   g116(.A1(new_n538), .A2(new_n541), .ZN(G171));
  AOI22_X1  g117(.A1(new_n513), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n543));
  NOR2_X1   g118(.A1(new_n543), .A2(new_n515), .ZN(new_n544));
  NAND2_X1  g119(.A1(new_n520), .A2(G43), .ZN(new_n545));
  INV_X1    g120(.A(G81), .ZN(new_n546));
  OAI21_X1  g121(.A(new_n545), .B1(new_n523), .B2(new_n546), .ZN(new_n547));
  NOR2_X1   g122(.A1(new_n544), .A2(new_n547), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n548), .A2(G860), .ZN(G153));
  AND3_X1   g124(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n550), .A2(G36), .ZN(G176));
  NAND2_X1  g126(.A1(G1), .A2(G3), .ZN(new_n552));
  XNOR2_X1  g127(.A(new_n552), .B(KEYINPUT8), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n550), .A2(new_n553), .ZN(G188));
  NAND2_X1  g129(.A1(new_n522), .A2(G543), .ZN(new_n555));
  INV_X1    g130(.A(G53), .ZN(new_n556));
  OAI21_X1  g131(.A(KEYINPUT9), .B1(new_n555), .B2(new_n556), .ZN(new_n557));
  INV_X1    g132(.A(KEYINPUT9), .ZN(new_n558));
  NAND3_X1  g133(.A1(new_n520), .A2(new_n558), .A3(G53), .ZN(new_n559));
  INV_X1    g134(.A(new_n523), .ZN(new_n560));
  AOI22_X1  g135(.A1(new_n557), .A2(new_n559), .B1(new_n560), .B2(G91), .ZN(new_n561));
  AOI22_X1  g136(.A1(new_n513), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n562));
  OR2_X1    g137(.A1(new_n562), .A2(new_n515), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n561), .A2(new_n563), .ZN(G299));
  INV_X1    g139(.A(G171), .ZN(G301));
  INV_X1    g140(.A(G166), .ZN(G303));
  OAI21_X1  g141(.A(G651), .B1(new_n513), .B2(G74), .ZN(new_n567));
  INV_X1    g142(.A(G49), .ZN(new_n568));
  INV_X1    g143(.A(G87), .ZN(new_n569));
  OAI221_X1 g144(.A(new_n567), .B1(new_n555), .B2(new_n568), .C1(new_n569), .C2(new_n523), .ZN(new_n570));
  XOR2_X1   g145(.A(new_n570), .B(KEYINPUT75), .Z(G288));
  NAND2_X1  g146(.A1(new_n520), .A2(G48), .ZN(new_n572));
  XNOR2_X1  g147(.A(new_n572), .B(KEYINPUT76), .ZN(new_n573));
  AOI22_X1  g148(.A1(new_n513), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n574));
  OR2_X1    g149(.A1(new_n574), .A2(new_n515), .ZN(new_n575));
  NAND2_X1  g150(.A1(new_n560), .A2(G86), .ZN(new_n576));
  NAND3_X1  g151(.A1(new_n573), .A2(new_n575), .A3(new_n576), .ZN(G305));
  AOI22_X1  g152(.A1(new_n513), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n578));
  NOR2_X1   g153(.A1(new_n578), .A2(new_n515), .ZN(new_n579));
  NAND2_X1  g154(.A1(new_n520), .A2(G47), .ZN(new_n580));
  XNOR2_X1  g155(.A(KEYINPUT77), .B(G85), .ZN(new_n581));
  OAI21_X1  g156(.A(new_n580), .B1(new_n523), .B2(new_n581), .ZN(new_n582));
  NOR2_X1   g157(.A1(new_n579), .A2(new_n582), .ZN(new_n583));
  INV_X1    g158(.A(new_n583), .ZN(G290));
  NAND2_X1  g159(.A1(G301), .A2(G868), .ZN(new_n585));
  AND3_X1   g160(.A1(new_n513), .A2(new_n522), .A3(G92), .ZN(new_n586));
  XNOR2_X1  g161(.A(new_n586), .B(KEYINPUT10), .ZN(new_n587));
  NAND2_X1  g162(.A1(new_n520), .A2(G54), .ZN(new_n588));
  AOI22_X1  g163(.A1(new_n513), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n589));
  OR2_X1    g164(.A1(new_n589), .A2(new_n515), .ZN(new_n590));
  NAND3_X1  g165(.A1(new_n587), .A2(new_n588), .A3(new_n590), .ZN(new_n591));
  INV_X1    g166(.A(new_n591), .ZN(new_n592));
  OAI21_X1  g167(.A(new_n585), .B1(new_n592), .B2(G868), .ZN(G284));
  OAI21_X1  g168(.A(new_n585), .B1(new_n592), .B2(G868), .ZN(G321));
  NAND2_X1  g169(.A1(G286), .A2(G868), .ZN(new_n595));
  XNOR2_X1  g170(.A(G299), .B(KEYINPUT78), .ZN(new_n596));
  OAI21_X1  g171(.A(new_n595), .B1(G868), .B2(new_n596), .ZN(G297));
  OAI21_X1  g172(.A(new_n595), .B1(G868), .B2(new_n596), .ZN(G280));
  INV_X1    g173(.A(G559), .ZN(new_n599));
  OAI21_X1  g174(.A(new_n592), .B1(new_n599), .B2(G860), .ZN(G148));
  NAND2_X1  g175(.A1(new_n592), .A2(new_n599), .ZN(new_n601));
  NAND2_X1  g176(.A1(new_n601), .A2(G868), .ZN(new_n602));
  OAI21_X1  g177(.A(new_n602), .B1(G868), .B2(new_n548), .ZN(G323));
  XNOR2_X1  g178(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g179(.A1(new_n488), .A2(G2104), .ZN(new_n605));
  XNOR2_X1  g180(.A(new_n605), .B(KEYINPUT12), .ZN(new_n606));
  XNOR2_X1  g181(.A(new_n606), .B(G2100), .ZN(new_n607));
  XNOR2_X1  g182(.A(KEYINPUT79), .B(KEYINPUT13), .ZN(new_n608));
  XNOR2_X1  g183(.A(new_n607), .B(new_n608), .ZN(new_n609));
  NAND2_X1  g184(.A1(new_n486), .A2(G123), .ZN(new_n610));
  XNOR2_X1  g185(.A(new_n610), .B(KEYINPUT80), .ZN(new_n611));
  OR2_X1    g186(.A1(G99), .A2(G2105), .ZN(new_n612));
  OAI211_X1 g187(.A(new_n612), .B(G2104), .C1(G111), .C2(new_n476), .ZN(new_n613));
  NAND2_X1  g188(.A1(new_n488), .A2(G135), .ZN(new_n614));
  AND3_X1   g189(.A1(new_n611), .A2(new_n613), .A3(new_n614), .ZN(new_n615));
  XNOR2_X1  g190(.A(new_n615), .B(G2096), .ZN(new_n616));
  NAND2_X1  g191(.A1(new_n609), .A2(new_n616), .ZN(G156));
  INV_X1    g192(.A(KEYINPUT83), .ZN(new_n618));
  XNOR2_X1  g193(.A(KEYINPUT15), .B(G2435), .ZN(new_n619));
  INV_X1    g194(.A(G2438), .ZN(new_n620));
  XNOR2_X1  g195(.A(new_n619), .B(new_n620), .ZN(new_n621));
  XOR2_X1   g196(.A(G2427), .B(G2430), .Z(new_n622));
  OAI21_X1  g197(.A(KEYINPUT14), .B1(new_n621), .B2(new_n622), .ZN(new_n623));
  XOR2_X1   g198(.A(new_n623), .B(KEYINPUT82), .Z(new_n624));
  NAND2_X1  g199(.A1(new_n621), .A2(new_n622), .ZN(new_n625));
  NAND2_X1  g200(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  XNOR2_X1  g201(.A(G2451), .B(G2454), .ZN(new_n627));
  INV_X1    g202(.A(new_n627), .ZN(new_n628));
  XNOR2_X1  g203(.A(new_n626), .B(new_n628), .ZN(new_n629));
  XOR2_X1   g204(.A(KEYINPUT81), .B(KEYINPUT16), .Z(new_n630));
  NAND2_X1  g205(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  XNOR2_X1  g206(.A(new_n626), .B(new_n627), .ZN(new_n632));
  INV_X1    g207(.A(new_n630), .ZN(new_n633));
  NAND2_X1  g208(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  NAND2_X1  g209(.A1(new_n631), .A2(new_n634), .ZN(new_n635));
  XNOR2_X1  g210(.A(G2443), .B(G2446), .ZN(new_n636));
  INV_X1    g211(.A(new_n636), .ZN(new_n637));
  NAND2_X1  g212(.A1(new_n635), .A2(new_n637), .ZN(new_n638));
  NAND3_X1  g213(.A1(new_n631), .A2(new_n634), .A3(new_n636), .ZN(new_n639));
  NAND2_X1  g214(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  XOR2_X1   g215(.A(G1341), .B(G1348), .Z(new_n641));
  OAI21_X1  g216(.A(new_n618), .B1(new_n640), .B2(new_n641), .ZN(new_n642));
  NAND2_X1  g217(.A1(new_n640), .A2(new_n641), .ZN(new_n643));
  INV_X1    g218(.A(new_n641), .ZN(new_n644));
  NAND4_X1  g219(.A1(new_n638), .A2(KEYINPUT83), .A3(new_n644), .A4(new_n639), .ZN(new_n645));
  NAND4_X1  g220(.A1(new_n642), .A2(new_n643), .A3(G14), .A4(new_n645), .ZN(new_n646));
  INV_X1    g221(.A(new_n646), .ZN(G401));
  XOR2_X1   g222(.A(G2084), .B(G2090), .Z(new_n648));
  INV_X1    g223(.A(new_n648), .ZN(new_n649));
  XOR2_X1   g224(.A(G2067), .B(G2678), .Z(new_n650));
  OR2_X1    g225(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  NAND2_X1  g226(.A1(new_n649), .A2(new_n650), .ZN(new_n652));
  NAND3_X1  g227(.A1(new_n651), .A2(new_n652), .A3(KEYINPUT17), .ZN(new_n653));
  INV_X1    g228(.A(KEYINPUT18), .ZN(new_n654));
  NAND2_X1  g229(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  XOR2_X1   g230(.A(G2072), .B(G2078), .Z(new_n656));
  AOI21_X1  g231(.A(new_n656), .B1(new_n651), .B2(KEYINPUT18), .ZN(new_n657));
  XNOR2_X1  g232(.A(new_n655), .B(new_n657), .ZN(new_n658));
  XNOR2_X1  g233(.A(G2096), .B(G2100), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n658), .B(new_n659), .ZN(G227));
  XNOR2_X1  g235(.A(G1971), .B(G1976), .ZN(new_n661));
  XNOR2_X1  g236(.A(new_n661), .B(KEYINPUT84), .ZN(new_n662));
  XOR2_X1   g237(.A(new_n662), .B(KEYINPUT19), .Z(new_n663));
  XOR2_X1   g238(.A(G1956), .B(G2474), .Z(new_n664));
  XOR2_X1   g239(.A(G1961), .B(G1966), .Z(new_n665));
  NAND2_X1  g240(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  XOR2_X1   g241(.A(new_n666), .B(KEYINPUT85), .Z(new_n667));
  NOR2_X1   g242(.A1(new_n663), .A2(new_n667), .ZN(new_n668));
  INV_X1    g243(.A(new_n663), .ZN(new_n669));
  NOR2_X1   g244(.A1(new_n664), .A2(new_n665), .ZN(new_n670));
  AOI22_X1  g245(.A1(new_n668), .A2(KEYINPUT20), .B1(new_n669), .B2(new_n670), .ZN(new_n671));
  INV_X1    g246(.A(new_n670), .ZN(new_n672));
  NAND3_X1  g247(.A1(new_n663), .A2(new_n666), .A3(new_n672), .ZN(new_n673));
  OAI211_X1 g248(.A(new_n671), .B(new_n673), .C1(KEYINPUT20), .C2(new_n668), .ZN(new_n674));
  XOR2_X1   g249(.A(KEYINPUT86), .B(KEYINPUT87), .Z(new_n675));
  XNOR2_X1  g250(.A(new_n674), .B(new_n675), .ZN(new_n676));
  XOR2_X1   g251(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n677));
  XNOR2_X1  g252(.A(new_n677), .B(G1991), .ZN(new_n678));
  XNOR2_X1  g253(.A(new_n676), .B(new_n678), .ZN(new_n679));
  XNOR2_X1  g254(.A(G1981), .B(G1986), .ZN(new_n680));
  XNOR2_X1  g255(.A(new_n680), .B(G1996), .ZN(new_n681));
  INV_X1    g256(.A(new_n681), .ZN(new_n682));
  XNOR2_X1  g257(.A(new_n679), .B(new_n682), .ZN(new_n683));
  INV_X1    g258(.A(new_n683), .ZN(G229));
  INV_X1    g259(.A(G16), .ZN(new_n685));
  NAND2_X1  g260(.A1(new_n685), .A2(G24), .ZN(new_n686));
  OAI21_X1  g261(.A(new_n686), .B1(new_n583), .B2(new_n685), .ZN(new_n687));
  XNOR2_X1  g262(.A(new_n687), .B(G1986), .ZN(new_n688));
  MUX2_X1   g263(.A(G23), .B(new_n570), .S(G16), .Z(new_n689));
  XNOR2_X1  g264(.A(new_n689), .B(KEYINPUT33), .ZN(new_n690));
  XNOR2_X1  g265(.A(new_n690), .B(G1976), .ZN(new_n691));
  NAND2_X1  g266(.A1(new_n685), .A2(G22), .ZN(new_n692));
  OAI21_X1  g267(.A(new_n692), .B1(G166), .B2(new_n685), .ZN(new_n693));
  NAND2_X1  g268(.A1(new_n693), .A2(G1971), .ZN(new_n694));
  NAND2_X1  g269(.A1(new_n685), .A2(G6), .ZN(new_n695));
  INV_X1    g270(.A(G305), .ZN(new_n696));
  OAI21_X1  g271(.A(new_n695), .B1(new_n696), .B2(new_n685), .ZN(new_n697));
  XOR2_X1   g272(.A(KEYINPUT32), .B(G1981), .Z(new_n698));
  INV_X1    g273(.A(new_n698), .ZN(new_n699));
  OAI21_X1  g274(.A(new_n694), .B1(new_n697), .B2(new_n699), .ZN(new_n700));
  AOI21_X1  g275(.A(new_n700), .B1(new_n697), .B2(new_n699), .ZN(new_n701));
  OAI211_X1 g276(.A(new_n691), .B(new_n701), .C1(G1971), .C2(new_n693), .ZN(new_n702));
  AOI21_X1  g277(.A(new_n688), .B1(new_n702), .B2(KEYINPUT34), .ZN(new_n703));
  INV_X1    g278(.A(G29), .ZN(new_n704));
  NAND2_X1  g279(.A1(new_n704), .A2(G25), .ZN(new_n705));
  NAND2_X1  g280(.A1(new_n488), .A2(G131), .ZN(new_n706));
  XOR2_X1   g281(.A(new_n706), .B(KEYINPUT88), .Z(new_n707));
  OR2_X1    g282(.A1(G95), .A2(G2105), .ZN(new_n708));
  OAI211_X1 g283(.A(new_n708), .B(G2104), .C1(G107), .C2(new_n476), .ZN(new_n709));
  NAND2_X1  g284(.A1(new_n486), .A2(G119), .ZN(new_n710));
  NAND3_X1  g285(.A1(new_n707), .A2(new_n709), .A3(new_n710), .ZN(new_n711));
  INV_X1    g286(.A(new_n711), .ZN(new_n712));
  OAI21_X1  g287(.A(new_n705), .B1(new_n712), .B2(new_n704), .ZN(new_n713));
  XNOR2_X1  g288(.A(new_n713), .B(KEYINPUT89), .ZN(new_n714));
  XNOR2_X1  g289(.A(KEYINPUT35), .B(G1991), .ZN(new_n715));
  INV_X1    g290(.A(new_n715), .ZN(new_n716));
  XNOR2_X1  g291(.A(new_n714), .B(new_n716), .ZN(new_n717));
  OAI211_X1 g292(.A(new_n703), .B(new_n717), .C1(KEYINPUT34), .C2(new_n702), .ZN(new_n718));
  XNOR2_X1  g293(.A(new_n718), .B(KEYINPUT36), .ZN(new_n719));
  XNOR2_X1  g294(.A(KEYINPUT31), .B(G11), .ZN(new_n720));
  NAND2_X1  g295(.A1(new_n704), .A2(G35), .ZN(new_n721));
  OAI21_X1  g296(.A(new_n721), .B1(G162), .B2(new_n704), .ZN(new_n722));
  XOR2_X1   g297(.A(new_n722), .B(KEYINPUT98), .Z(new_n723));
  XNOR2_X1  g298(.A(new_n723), .B(KEYINPUT29), .ZN(new_n724));
  XOR2_X1   g299(.A(new_n724), .B(G2090), .Z(new_n725));
  NAND2_X1  g300(.A1(G160), .A2(G29), .ZN(new_n726));
  XNOR2_X1  g301(.A(KEYINPUT93), .B(KEYINPUT24), .ZN(new_n727));
  XNOR2_X1  g302(.A(new_n727), .B(G34), .ZN(new_n728));
  NAND2_X1  g303(.A1(new_n728), .A2(new_n704), .ZN(new_n729));
  AOI21_X1  g304(.A(G2084), .B1(new_n726), .B2(new_n729), .ZN(new_n730));
  NOR2_X1   g305(.A1(G4), .A2(G16), .ZN(new_n731));
  AOI21_X1  g306(.A(new_n731), .B1(new_n592), .B2(G16), .ZN(new_n732));
  AOI21_X1  g307(.A(new_n730), .B1(new_n732), .B2(G1348), .ZN(new_n733));
  INV_X1    g308(.A(KEYINPUT96), .ZN(new_n734));
  OAI21_X1  g309(.A(new_n734), .B1(G5), .B2(G16), .ZN(new_n735));
  OR3_X1    g310(.A1(new_n734), .A2(G5), .A3(G16), .ZN(new_n736));
  OAI211_X1 g311(.A(new_n735), .B(new_n736), .C1(G301), .C2(new_n685), .ZN(new_n737));
  XNOR2_X1  g312(.A(KEYINPUT97), .B(G1961), .ZN(new_n738));
  OR2_X1    g313(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  NOR2_X1   g314(.A1(G16), .A2(G19), .ZN(new_n740));
  AOI21_X1  g315(.A(new_n740), .B1(new_n548), .B2(G16), .ZN(new_n741));
  NAND2_X1  g316(.A1(new_n741), .A2(G1341), .ZN(new_n742));
  NAND2_X1  g317(.A1(new_n737), .A2(new_n738), .ZN(new_n743));
  NAND3_X1  g318(.A1(new_n739), .A2(new_n742), .A3(new_n743), .ZN(new_n744));
  NOR2_X1   g319(.A1(new_n741), .A2(G1341), .ZN(new_n745));
  NAND2_X1  g320(.A1(new_n704), .A2(G27), .ZN(new_n746));
  OAI21_X1  g321(.A(new_n746), .B1(G164), .B2(new_n704), .ZN(new_n747));
  XNOR2_X1  g322(.A(new_n747), .B(G2078), .ZN(new_n748));
  NAND2_X1  g323(.A1(new_n615), .A2(G29), .ZN(new_n749));
  OR2_X1    g324(.A1(G29), .A2(G33), .ZN(new_n750));
  NAND3_X1  g325(.A1(new_n476), .A2(G103), .A3(G2104), .ZN(new_n751));
  XOR2_X1   g326(.A(new_n751), .B(KEYINPUT25), .Z(new_n752));
  NAND2_X1  g327(.A1(new_n488), .A2(G139), .ZN(new_n753));
  AOI22_X1  g328(.A1(new_n467), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n754));
  OAI211_X1 g329(.A(new_n752), .B(new_n753), .C1(new_n476), .C2(new_n754), .ZN(new_n755));
  OAI21_X1  g330(.A(new_n750), .B1(new_n755), .B2(new_n704), .ZN(new_n756));
  INV_X1    g331(.A(G2072), .ZN(new_n757));
  OR2_X1    g332(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  NAND2_X1  g333(.A1(new_n756), .A2(new_n757), .ZN(new_n759));
  INV_X1    g334(.A(KEYINPUT30), .ZN(new_n760));
  OR2_X1    g335(.A1(new_n760), .A2(G28), .ZN(new_n761));
  NAND2_X1  g336(.A1(new_n760), .A2(G28), .ZN(new_n762));
  NAND3_X1  g337(.A1(new_n761), .A2(new_n762), .A3(new_n704), .ZN(new_n763));
  NAND4_X1  g338(.A1(new_n749), .A2(new_n758), .A3(new_n759), .A4(new_n763), .ZN(new_n764));
  NOR4_X1   g339(.A1(new_n744), .A2(new_n745), .A3(new_n748), .A4(new_n764), .ZN(new_n765));
  NAND3_X1  g340(.A1(new_n725), .A2(new_n733), .A3(new_n765), .ZN(new_n766));
  AOI22_X1  g341(.A1(G129), .A2(new_n486), .B1(new_n488), .B2(G141), .ZN(new_n767));
  XOR2_X1   g342(.A(KEYINPUT94), .B(KEYINPUT26), .Z(new_n768));
  NAND3_X1  g343(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n769));
  XNOR2_X1  g344(.A(new_n768), .B(new_n769), .ZN(new_n770));
  INV_X1    g345(.A(G105), .ZN(new_n771));
  OAI211_X1 g346(.A(new_n767), .B(new_n770), .C1(new_n771), .C2(new_n494), .ZN(new_n772));
  MUX2_X1   g347(.A(G32), .B(new_n772), .S(G29), .Z(new_n773));
  XOR2_X1   g348(.A(new_n773), .B(KEYINPUT95), .Z(new_n774));
  XOR2_X1   g349(.A(KEYINPUT27), .B(G1996), .Z(new_n775));
  INV_X1    g350(.A(new_n775), .ZN(new_n776));
  AND2_X1   g351(.A1(new_n774), .A2(new_n776), .ZN(new_n777));
  NOR2_X1   g352(.A1(new_n774), .A2(new_n776), .ZN(new_n778));
  NOR2_X1   g353(.A1(new_n732), .A2(G1348), .ZN(new_n779));
  NOR3_X1   g354(.A1(new_n777), .A2(new_n778), .A3(new_n779), .ZN(new_n780));
  NAND3_X1  g355(.A1(new_n726), .A2(G2084), .A3(new_n729), .ZN(new_n781));
  INV_X1    g356(.A(G299), .ZN(new_n782));
  OAI21_X1  g357(.A(KEYINPUT23), .B1(new_n782), .B2(new_n685), .ZN(new_n783));
  NAND2_X1  g358(.A1(new_n685), .A2(G20), .ZN(new_n784));
  MUX2_X1   g359(.A(KEYINPUT23), .B(new_n783), .S(new_n784), .Z(new_n785));
  NAND2_X1  g360(.A1(new_n785), .A2(G1956), .ZN(new_n786));
  OR2_X1    g361(.A1(new_n785), .A2(G1956), .ZN(new_n787));
  NAND4_X1  g362(.A1(new_n780), .A2(new_n781), .A3(new_n786), .A4(new_n787), .ZN(new_n788));
  NAND2_X1  g363(.A1(new_n704), .A2(G26), .ZN(new_n789));
  XOR2_X1   g364(.A(new_n789), .B(KEYINPUT92), .Z(new_n790));
  XNOR2_X1  g365(.A(new_n790), .B(KEYINPUT28), .ZN(new_n791));
  NAND2_X1  g366(.A1(new_n486), .A2(G128), .ZN(new_n792));
  XNOR2_X1  g367(.A(new_n792), .B(KEYINPUT91), .ZN(new_n793));
  OR2_X1    g368(.A1(G104), .A2(G2105), .ZN(new_n794));
  OAI211_X1 g369(.A(new_n794), .B(G2104), .C1(G116), .C2(new_n476), .ZN(new_n795));
  AND2_X1   g370(.A1(new_n793), .A2(new_n795), .ZN(new_n796));
  NAND2_X1  g371(.A1(new_n488), .A2(G140), .ZN(new_n797));
  XNOR2_X1  g372(.A(new_n797), .B(KEYINPUT90), .ZN(new_n798));
  NAND2_X1  g373(.A1(new_n796), .A2(new_n798), .ZN(new_n799));
  AOI21_X1  g374(.A(new_n791), .B1(new_n799), .B2(G29), .ZN(new_n800));
  INV_X1    g375(.A(G2067), .ZN(new_n801));
  XNOR2_X1  g376(.A(new_n800), .B(new_n801), .ZN(new_n802));
  NOR2_X1   g377(.A1(G16), .A2(G21), .ZN(new_n803));
  AOI21_X1  g378(.A(new_n803), .B1(G168), .B2(G16), .ZN(new_n804));
  XNOR2_X1  g379(.A(new_n804), .B(G1966), .ZN(new_n805));
  NOR4_X1   g380(.A1(new_n766), .A2(new_n788), .A3(new_n802), .A4(new_n805), .ZN(new_n806));
  NAND3_X1  g381(.A1(new_n719), .A2(new_n720), .A3(new_n806), .ZN(G150));
  INV_X1    g382(.A(KEYINPUT99), .ZN(new_n808));
  XNOR2_X1  g383(.A(G150), .B(new_n808), .ZN(G311));
  AOI22_X1  g384(.A1(new_n560), .A2(G93), .B1(G55), .B2(new_n520), .ZN(new_n810));
  AOI22_X1  g385(.A1(new_n513), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n811));
  OAI21_X1  g386(.A(new_n810), .B1(new_n515), .B2(new_n811), .ZN(new_n812));
  XNOR2_X1  g387(.A(KEYINPUT100), .B(G860), .ZN(new_n813));
  NAND2_X1  g388(.A1(new_n812), .A2(new_n813), .ZN(new_n814));
  XOR2_X1   g389(.A(new_n814), .B(KEYINPUT37), .Z(new_n815));
  XNOR2_X1  g390(.A(new_n812), .B(new_n548), .ZN(new_n816));
  XNOR2_X1  g391(.A(new_n816), .B(KEYINPUT38), .ZN(new_n817));
  NOR2_X1   g392(.A1(new_n591), .A2(new_n599), .ZN(new_n818));
  XNOR2_X1  g393(.A(new_n817), .B(new_n818), .ZN(new_n819));
  INV_X1    g394(.A(KEYINPUT39), .ZN(new_n820));
  OAI21_X1  g395(.A(new_n819), .B1(KEYINPUT101), .B2(new_n820), .ZN(new_n821));
  XNOR2_X1  g396(.A(KEYINPUT101), .B(KEYINPUT39), .ZN(new_n822));
  OAI21_X1  g397(.A(new_n821), .B1(new_n822), .B2(new_n819), .ZN(new_n823));
  OAI21_X1  g398(.A(new_n815), .B1(new_n823), .B2(new_n813), .ZN(G145));
  XNOR2_X1  g399(.A(new_n799), .B(new_n772), .ZN(new_n825));
  XNOR2_X1  g400(.A(new_n825), .B(new_n755), .ZN(new_n826));
  AOI22_X1  g401(.A1(new_n467), .A2(G126), .B1(G114), .B2(G2104), .ZN(new_n827));
  OAI22_X1  g402(.A1(new_n827), .A2(new_n476), .B1(new_n495), .B2(new_n494), .ZN(new_n828));
  INV_X1    g403(.A(KEYINPUT103), .ZN(new_n829));
  NAND2_X1  g404(.A1(new_n505), .A2(new_n829), .ZN(new_n830));
  NAND3_X1  g405(.A1(new_n502), .A2(new_n504), .A3(KEYINPUT103), .ZN(new_n831));
  AOI21_X1  g406(.A(new_n828), .B1(new_n830), .B2(new_n831), .ZN(new_n832));
  XNOR2_X1  g407(.A(new_n826), .B(new_n832), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n486), .A2(G130), .ZN(new_n834));
  XOR2_X1   g409(.A(new_n834), .B(KEYINPUT104), .Z(new_n835));
  NAND2_X1  g410(.A1(new_n488), .A2(G142), .ZN(new_n836));
  NOR2_X1   g411(.A1(G106), .A2(G2105), .ZN(new_n837));
  OAI21_X1  g412(.A(G2104), .B1(new_n476), .B2(G118), .ZN(new_n838));
  OAI211_X1 g413(.A(new_n835), .B(new_n836), .C1(new_n837), .C2(new_n838), .ZN(new_n839));
  XNOR2_X1  g414(.A(new_n839), .B(new_n606), .ZN(new_n840));
  XNOR2_X1  g415(.A(new_n840), .B(new_n711), .ZN(new_n841));
  OR2_X1    g416(.A1(new_n833), .A2(new_n841), .ZN(new_n842));
  XNOR2_X1  g417(.A(new_n492), .B(KEYINPUT102), .ZN(new_n843));
  XNOR2_X1  g418(.A(new_n843), .B(G160), .ZN(new_n844));
  XNOR2_X1  g419(.A(new_n844), .B(new_n615), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n833), .A2(new_n841), .ZN(new_n846));
  NAND3_X1  g421(.A1(new_n842), .A2(new_n845), .A3(new_n846), .ZN(new_n847));
  INV_X1    g422(.A(G37), .ZN(new_n848));
  INV_X1    g423(.A(KEYINPUT105), .ZN(new_n849));
  NAND2_X1  g424(.A1(new_n841), .A2(new_n849), .ZN(new_n850));
  XNOR2_X1  g425(.A(new_n833), .B(new_n850), .ZN(new_n851));
  OAI211_X1 g426(.A(new_n847), .B(new_n848), .C1(new_n851), .C2(new_n845), .ZN(new_n852));
  XNOR2_X1  g427(.A(new_n852), .B(KEYINPUT40), .ZN(G395));
  NOR2_X1   g428(.A1(new_n812), .A2(G868), .ZN(new_n854));
  XNOR2_X1  g429(.A(G166), .B(new_n570), .ZN(new_n855));
  XNOR2_X1  g430(.A(new_n855), .B(G290), .ZN(new_n856));
  XNOR2_X1  g431(.A(new_n856), .B(new_n696), .ZN(new_n857));
  XOR2_X1   g432(.A(new_n857), .B(KEYINPUT108), .Z(new_n858));
  XNOR2_X1  g433(.A(new_n858), .B(KEYINPUT42), .ZN(new_n859));
  INV_X1    g434(.A(new_n859), .ZN(new_n860));
  XNOR2_X1  g435(.A(new_n601), .B(new_n816), .ZN(new_n861));
  XNOR2_X1  g436(.A(new_n591), .B(G299), .ZN(new_n862));
  NOR2_X1   g437(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n862), .A2(KEYINPUT41), .ZN(new_n864));
  XOR2_X1   g439(.A(new_n864), .B(KEYINPUT107), .Z(new_n865));
  NOR2_X1   g440(.A1(new_n862), .A2(KEYINPUT41), .ZN(new_n866));
  XNOR2_X1  g441(.A(new_n866), .B(KEYINPUT106), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n865), .A2(new_n867), .ZN(new_n868));
  AOI21_X1  g443(.A(new_n863), .B1(new_n868), .B2(new_n861), .ZN(new_n869));
  OR2_X1    g444(.A1(new_n869), .A2(KEYINPUT109), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n869), .A2(KEYINPUT109), .ZN(new_n871));
  NAND3_X1  g446(.A1(new_n860), .A2(new_n870), .A3(new_n871), .ZN(new_n872));
  NAND3_X1  g447(.A1(new_n859), .A2(KEYINPUT109), .A3(new_n869), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  AOI21_X1  g449(.A(new_n854), .B1(new_n874), .B2(G868), .ZN(G295));
  AOI21_X1  g450(.A(new_n854), .B1(new_n874), .B2(G868), .ZN(G331));
  XNOR2_X1  g451(.A(G286), .B(new_n816), .ZN(new_n877));
  XNOR2_X1  g452(.A(new_n877), .B(G171), .ZN(new_n878));
  OR2_X1    g453(.A1(new_n878), .A2(new_n862), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n868), .A2(new_n878), .ZN(new_n880));
  NAND3_X1  g455(.A1(new_n879), .A2(new_n880), .A3(new_n857), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n881), .A2(new_n848), .ZN(new_n882));
  AOI21_X1  g457(.A(new_n857), .B1(new_n879), .B2(new_n880), .ZN(new_n883));
  OAI21_X1  g458(.A(KEYINPUT43), .B1(new_n882), .B2(new_n883), .ZN(new_n884));
  INV_X1    g459(.A(new_n864), .ZN(new_n885));
  OAI21_X1  g460(.A(new_n878), .B1(new_n885), .B2(new_n866), .ZN(new_n886));
  NAND3_X1  g461(.A1(new_n879), .A2(KEYINPUT110), .A3(new_n886), .ZN(new_n887));
  INV_X1    g462(.A(new_n857), .ZN(new_n888));
  OAI211_X1 g463(.A(new_n887), .B(new_n888), .C1(KEYINPUT110), .C2(new_n879), .ZN(new_n889));
  NAND3_X1  g464(.A1(new_n889), .A2(new_n848), .A3(new_n881), .ZN(new_n890));
  OAI21_X1  g465(.A(new_n884), .B1(new_n890), .B2(KEYINPUT43), .ZN(new_n891));
  INV_X1    g466(.A(KEYINPUT43), .ZN(new_n892));
  OAI21_X1  g467(.A(new_n892), .B1(new_n882), .B2(new_n883), .ZN(new_n893));
  OAI21_X1  g468(.A(new_n893), .B1(new_n890), .B2(new_n892), .ZN(new_n894));
  MUX2_X1   g469(.A(new_n891), .B(new_n894), .S(KEYINPUT44), .Z(G397));
  AND3_X1   g470(.A1(new_n502), .A2(new_n504), .A3(KEYINPUT103), .ZN(new_n896));
  AOI21_X1  g471(.A(KEYINPUT103), .B1(new_n502), .B2(new_n504), .ZN(new_n897));
  OAI21_X1  g472(.A(new_n500), .B1(new_n896), .B2(new_n897), .ZN(new_n898));
  INV_X1    g473(.A(G1384), .ZN(new_n899));
  AOI21_X1  g474(.A(KEYINPUT45), .B1(new_n898), .B2(new_n899), .ZN(new_n900));
  INV_X1    g475(.A(new_n900), .ZN(new_n901));
  NAND3_X1  g476(.A1(new_n475), .A2(new_n482), .A3(G40), .ZN(new_n902));
  OR3_X1    g477(.A1(new_n901), .A2(KEYINPUT111), .A3(new_n902), .ZN(new_n903));
  OAI21_X1  g478(.A(KEYINPUT111), .B1(new_n901), .B2(new_n902), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  INV_X1    g480(.A(new_n905), .ZN(new_n906));
  NAND2_X1  g481(.A1(new_n799), .A2(G2067), .ZN(new_n907));
  NAND3_X1  g482(.A1(new_n796), .A2(new_n801), .A3(new_n798), .ZN(new_n908));
  AND2_X1   g483(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  INV_X1    g484(.A(new_n909), .ZN(new_n910));
  OAI21_X1  g485(.A(new_n906), .B1(new_n910), .B2(new_n772), .ZN(new_n911));
  INV_X1    g486(.A(G1996), .ZN(new_n912));
  NAND3_X1  g487(.A1(new_n906), .A2(KEYINPUT46), .A3(new_n912), .ZN(new_n913));
  INV_X1    g488(.A(KEYINPUT46), .ZN(new_n914));
  OAI21_X1  g489(.A(new_n914), .B1(new_n905), .B2(G1996), .ZN(new_n915));
  NAND3_X1  g490(.A1(new_n911), .A2(new_n913), .A3(new_n915), .ZN(new_n916));
  XOR2_X1   g491(.A(new_n916), .B(KEYINPUT47), .Z(new_n917));
  NOR2_X1   g492(.A1(G290), .A2(G1986), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n906), .A2(new_n918), .ZN(new_n919));
  XOR2_X1   g494(.A(new_n919), .B(KEYINPUT48), .Z(new_n920));
  XNOR2_X1  g495(.A(new_n772), .B(new_n912), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n909), .A2(new_n921), .ZN(new_n922));
  INV_X1    g497(.A(new_n922), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n711), .A2(new_n715), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n712), .A2(new_n716), .ZN(new_n925));
  NAND3_X1  g500(.A1(new_n923), .A2(new_n924), .A3(new_n925), .ZN(new_n926));
  AOI21_X1  g501(.A(new_n920), .B1(new_n906), .B2(new_n926), .ZN(new_n927));
  OAI21_X1  g502(.A(new_n908), .B1(new_n922), .B2(new_n925), .ZN(new_n928));
  AOI211_X1 g503(.A(new_n917), .B(new_n927), .C1(new_n906), .C2(new_n928), .ZN(new_n929));
  INV_X1    g504(.A(KEYINPUT125), .ZN(new_n930));
  INV_X1    g505(.A(new_n926), .ZN(new_n931));
  INV_X1    g506(.A(G1986), .ZN(new_n932));
  OAI21_X1  g507(.A(new_n931), .B1(new_n932), .B2(new_n583), .ZN(new_n933));
  OAI21_X1  g508(.A(new_n906), .B1(new_n933), .B2(new_n918), .ZN(new_n934));
  INV_X1    g509(.A(KEYINPUT112), .ZN(new_n935));
  NAND3_X1  g510(.A1(new_n898), .A2(KEYINPUT45), .A3(new_n899), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n506), .A2(new_n899), .ZN(new_n937));
  INV_X1    g512(.A(KEYINPUT45), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  AND3_X1   g514(.A1(new_n475), .A2(G40), .A3(new_n482), .ZN(new_n940));
  NAND3_X1  g515(.A1(new_n936), .A2(new_n939), .A3(new_n940), .ZN(new_n941));
  INV_X1    g516(.A(G1971), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  INV_X1    g518(.A(new_n943), .ZN(new_n944));
  INV_X1    g519(.A(KEYINPUT50), .ZN(new_n945));
  NAND3_X1  g520(.A1(new_n898), .A2(new_n945), .A3(new_n899), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n937), .A2(KEYINPUT50), .ZN(new_n947));
  NAND3_X1  g522(.A1(new_n946), .A2(new_n947), .A3(new_n940), .ZN(new_n948));
  NOR2_X1   g523(.A1(new_n948), .A2(G2090), .ZN(new_n949));
  OAI21_X1  g524(.A(G8), .B1(new_n944), .B2(new_n949), .ZN(new_n950));
  NAND2_X1  g525(.A1(G303), .A2(G8), .ZN(new_n951));
  XNOR2_X1  g526(.A(new_n951), .B(KEYINPUT55), .ZN(new_n952));
  OAI21_X1  g527(.A(new_n935), .B1(new_n950), .B2(new_n952), .ZN(new_n953));
  INV_X1    g528(.A(G8), .ZN(new_n954));
  INV_X1    g529(.A(new_n949), .ZN(new_n955));
  AOI21_X1  g530(.A(new_n954), .B1(new_n955), .B2(new_n943), .ZN(new_n956));
  INV_X1    g531(.A(new_n952), .ZN(new_n957));
  NAND3_X1  g532(.A1(new_n956), .A2(KEYINPUT112), .A3(new_n957), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n953), .A2(new_n958), .ZN(new_n959));
  INV_X1    g534(.A(KEYINPUT113), .ZN(new_n960));
  NAND2_X1  g535(.A1(new_n898), .A2(new_n899), .ZN(new_n961));
  NOR2_X1   g536(.A1(new_n961), .A2(new_n902), .ZN(new_n962));
  OAI21_X1  g537(.A(new_n960), .B1(new_n962), .B2(new_n954), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n830), .A2(new_n831), .ZN(new_n964));
  AOI21_X1  g539(.A(G1384), .B1(new_n964), .B2(new_n500), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n965), .A2(new_n940), .ZN(new_n966));
  NAND3_X1  g541(.A1(new_n966), .A2(KEYINPUT113), .A3(G8), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n963), .A2(new_n967), .ZN(new_n968));
  INV_X1    g543(.A(G1976), .ZN(new_n969));
  OAI21_X1  g544(.A(new_n968), .B1(new_n969), .B2(new_n570), .ZN(new_n970));
  AND2_X1   g545(.A1(G305), .A2(G1981), .ZN(new_n971));
  NOR2_X1   g546(.A1(G305), .A2(G1981), .ZN(new_n972));
  OAI21_X1  g547(.A(KEYINPUT114), .B1(new_n971), .B2(new_n972), .ZN(new_n973));
  INV_X1    g548(.A(KEYINPUT49), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n973), .A2(new_n974), .ZN(new_n975));
  OAI211_X1 g550(.A(KEYINPUT114), .B(KEYINPUT49), .C1(new_n971), .C2(new_n972), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n975), .A2(new_n976), .ZN(new_n977));
  AOI22_X1  g552(.A1(KEYINPUT52), .A2(new_n970), .B1(new_n977), .B2(new_n968), .ZN(new_n978));
  NAND3_X1  g553(.A1(new_n506), .A2(new_n945), .A3(new_n899), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n940), .A2(new_n979), .ZN(new_n980));
  AOI21_X1  g555(.A(new_n945), .B1(new_n898), .B2(new_n899), .ZN(new_n981));
  NOR3_X1   g556(.A1(new_n980), .A2(new_n981), .A3(G2090), .ZN(new_n982));
  OAI21_X1  g557(.A(G8), .B1(new_n944), .B2(new_n982), .ZN(new_n983));
  NAND2_X1  g558(.A1(new_n983), .A2(new_n952), .ZN(new_n984));
  AOI21_X1  g559(.A(KEYINPUT52), .B1(G288), .B2(new_n969), .ZN(new_n985));
  OAI211_X1 g560(.A(new_n968), .B(new_n985), .C1(new_n969), .C2(new_n570), .ZN(new_n986));
  NAND4_X1  g561(.A1(new_n959), .A2(new_n978), .A3(new_n984), .A4(new_n986), .ZN(new_n987));
  INV_X1    g562(.A(KEYINPUT116), .ZN(new_n988));
  OAI21_X1  g563(.A(new_n988), .B1(new_n900), .B2(new_n902), .ZN(new_n989));
  OAI211_X1 g564(.A(KEYINPUT116), .B(new_n940), .C1(new_n965), .C2(KEYINPUT45), .ZN(new_n990));
  INV_X1    g565(.A(KEYINPUT53), .ZN(new_n991));
  NOR2_X1   g566(.A1(new_n991), .A2(G2078), .ZN(new_n992));
  NAND3_X1  g567(.A1(new_n506), .A2(KEYINPUT45), .A3(new_n899), .ZN(new_n993));
  NAND4_X1  g568(.A1(new_n989), .A2(new_n990), .A3(new_n992), .A4(new_n993), .ZN(new_n994));
  INV_X1    g569(.A(G2078), .ZN(new_n995));
  NAND4_X1  g570(.A1(new_n936), .A2(new_n939), .A3(new_n995), .A4(new_n940), .ZN(new_n996));
  INV_X1    g571(.A(G1961), .ZN(new_n997));
  AOI22_X1  g572(.A1(new_n996), .A2(new_n991), .B1(new_n948), .B2(new_n997), .ZN(new_n998));
  AOI21_X1  g573(.A(G301), .B1(new_n994), .B2(new_n998), .ZN(new_n999));
  INV_X1    g574(.A(new_n999), .ZN(new_n1000));
  OR2_X1    g575(.A1(new_n1000), .A2(KEYINPUT62), .ZN(new_n1001));
  AOI21_X1  g576(.A(KEYINPUT118), .B1(new_n557), .B2(new_n559), .ZN(new_n1002));
  NOR2_X1   g577(.A1(new_n1002), .A2(KEYINPUT57), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n1003), .A2(G299), .ZN(new_n1004));
  OAI211_X1 g579(.A(new_n561), .B(new_n563), .C1(new_n1002), .C2(KEYINPUT57), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n1004), .A2(new_n1005), .ZN(new_n1006));
  INV_X1    g581(.A(new_n1006), .ZN(new_n1007));
  XNOR2_X1  g582(.A(KEYINPUT56), .B(G2072), .ZN(new_n1008));
  NAND4_X1  g583(.A1(new_n936), .A2(new_n939), .A3(new_n940), .A4(new_n1008), .ZN(new_n1009));
  INV_X1    g584(.A(new_n1009), .ZN(new_n1010));
  AOI211_X1 g585(.A(KEYINPUT50), .B(G1384), .C1(new_n500), .C2(new_n505), .ZN(new_n1011));
  NOR2_X1   g586(.A1(new_n1011), .A2(new_n902), .ZN(new_n1012));
  OAI21_X1  g587(.A(KEYINPUT50), .B1(new_n832), .B2(G1384), .ZN(new_n1013));
  AOI21_X1  g588(.A(G1956), .B1(new_n1012), .B2(new_n1013), .ZN(new_n1014));
  OAI21_X1  g589(.A(new_n1007), .B1(new_n1010), .B2(new_n1014), .ZN(new_n1015));
  INV_X1    g590(.A(G1956), .ZN(new_n1016));
  OAI21_X1  g591(.A(new_n1016), .B1(new_n980), .B2(new_n981), .ZN(new_n1017));
  NAND3_X1  g592(.A1(new_n1017), .A2(new_n1006), .A3(new_n1009), .ZN(new_n1018));
  INV_X1    g593(.A(new_n1018), .ZN(new_n1019));
  AOI21_X1  g594(.A(new_n902), .B1(KEYINPUT50), .B2(new_n937), .ZN(new_n1020));
  AOI21_X1  g595(.A(G1348), .B1(new_n1020), .B2(new_n946), .ZN(new_n1021));
  NOR3_X1   g596(.A1(new_n961), .A2(G2067), .A3(new_n902), .ZN(new_n1022));
  OAI21_X1  g597(.A(new_n592), .B1(new_n1021), .B2(new_n1022), .ZN(new_n1023));
  OAI21_X1  g598(.A(new_n1015), .B1(new_n1019), .B2(new_n1023), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n1018), .A2(KEYINPUT120), .ZN(new_n1025));
  INV_X1    g600(.A(KEYINPUT120), .ZN(new_n1026));
  NAND4_X1  g601(.A1(new_n1017), .A2(new_n1026), .A3(new_n1006), .A4(new_n1009), .ZN(new_n1027));
  NAND3_X1  g602(.A1(new_n1025), .A2(KEYINPUT61), .A3(new_n1027), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n1028), .A2(KEYINPUT121), .ZN(new_n1029));
  INV_X1    g604(.A(KEYINPUT121), .ZN(new_n1030));
  NAND4_X1  g605(.A1(new_n1025), .A2(new_n1030), .A3(KEYINPUT61), .A4(new_n1027), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n1029), .A2(new_n1031), .ZN(new_n1032));
  INV_X1    g607(.A(G1348), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n948), .A2(new_n1033), .ZN(new_n1034));
  INV_X1    g609(.A(KEYINPUT60), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n962), .A2(new_n801), .ZN(new_n1036));
  NAND4_X1  g611(.A1(new_n1034), .A2(new_n1035), .A3(new_n1036), .A4(new_n592), .ZN(new_n1037));
  NAND2_X1  g612(.A1(KEYINPUT119), .A2(KEYINPUT59), .ZN(new_n1038));
  NAND4_X1  g613(.A1(new_n936), .A2(new_n939), .A3(new_n912), .A4(new_n940), .ZN(new_n1039));
  XOR2_X1   g614(.A(KEYINPUT58), .B(G1341), .Z(new_n1040));
  OAI21_X1  g615(.A(new_n1040), .B1(new_n961), .B2(new_n902), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n1039), .A2(new_n1041), .ZN(new_n1042));
  AOI21_X1  g617(.A(new_n1038), .B1(new_n1042), .B2(new_n548), .ZN(new_n1043));
  INV_X1    g618(.A(new_n548), .ZN(new_n1044));
  INV_X1    g619(.A(new_n1038), .ZN(new_n1045));
  AOI211_X1 g620(.A(new_n1044), .B(new_n1045), .C1(new_n1039), .C2(new_n1041), .ZN(new_n1046));
  OAI21_X1  g621(.A(new_n1037), .B1(new_n1043), .B2(new_n1046), .ZN(new_n1047));
  AOI21_X1  g622(.A(KEYINPUT61), .B1(new_n1015), .B2(new_n1018), .ZN(new_n1048));
  NAND3_X1  g623(.A1(new_n1034), .A2(new_n591), .A3(new_n1036), .ZN(new_n1049));
  AOI21_X1  g624(.A(new_n1035), .B1(new_n1023), .B2(new_n1049), .ZN(new_n1050));
  NOR3_X1   g625(.A1(new_n1047), .A2(new_n1048), .A3(new_n1050), .ZN(new_n1051));
  AOI21_X1  g626(.A(new_n1024), .B1(new_n1032), .B2(new_n1051), .ZN(new_n1052));
  XOR2_X1   g627(.A(KEYINPUT123), .B(KEYINPUT54), .Z(new_n1053));
  NAND3_X1  g628(.A1(new_n901), .A2(new_n936), .A3(new_n992), .ZN(new_n1054));
  XNOR2_X1  g629(.A(new_n902), .B(KEYINPUT124), .ZN(new_n1055));
  OAI21_X1  g630(.A(new_n998), .B1(new_n1054), .B2(new_n1055), .ZN(new_n1056));
  NOR2_X1   g631(.A1(new_n1056), .A2(G171), .ZN(new_n1057));
  OAI21_X1  g632(.A(new_n1053), .B1(new_n1057), .B2(new_n999), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n1056), .A2(G171), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n994), .A2(new_n998), .ZN(new_n1060));
  OAI211_X1 g635(.A(new_n1059), .B(KEYINPUT54), .C1(G171), .C2(new_n1060), .ZN(new_n1061));
  NAND2_X1  g636(.A1(new_n1058), .A2(new_n1061), .ZN(new_n1062));
  OAI21_X1  g637(.A(new_n1001), .B1(new_n1052), .B2(new_n1062), .ZN(new_n1063));
  NAND3_X1  g638(.A1(new_n989), .A2(new_n990), .A3(new_n993), .ZN(new_n1064));
  INV_X1    g639(.A(G1966), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n1064), .A2(new_n1065), .ZN(new_n1066));
  XOR2_X1   g641(.A(KEYINPUT117), .B(G2084), .Z(new_n1067));
  AND4_X1   g642(.A1(new_n940), .A2(new_n946), .A3(new_n947), .A4(new_n1067), .ZN(new_n1068));
  INV_X1    g643(.A(new_n1068), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n1066), .A2(new_n1069), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n1070), .A2(KEYINPUT122), .ZN(new_n1071));
  INV_X1    g646(.A(KEYINPUT122), .ZN(new_n1072));
  NAND3_X1  g647(.A1(new_n1066), .A2(new_n1072), .A3(new_n1069), .ZN(new_n1073));
  NOR2_X1   g648(.A1(G168), .A2(new_n954), .ZN(new_n1074));
  NAND3_X1  g649(.A1(new_n1071), .A2(new_n1073), .A3(new_n1074), .ZN(new_n1075));
  AOI21_X1  g650(.A(new_n1072), .B1(new_n1066), .B2(new_n1069), .ZN(new_n1076));
  AOI211_X1 g651(.A(KEYINPUT122), .B(new_n1068), .C1(new_n1064), .C2(new_n1065), .ZN(new_n1077));
  OAI21_X1  g652(.A(G168), .B1(new_n1076), .B2(new_n1077), .ZN(new_n1078));
  NAND4_X1  g653(.A1(new_n1075), .A2(new_n1078), .A3(KEYINPUT51), .A4(G8), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n1070), .A2(G8), .ZN(new_n1080));
  NOR2_X1   g655(.A1(new_n1074), .A2(KEYINPUT51), .ZN(new_n1081));
  NAND2_X1  g656(.A1(new_n1080), .A2(new_n1081), .ZN(new_n1082));
  AND2_X1   g657(.A1(new_n1079), .A2(new_n1082), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n1063), .A2(new_n1083), .ZN(new_n1084));
  AOI21_X1  g659(.A(new_n1000), .B1(new_n1079), .B2(new_n1082), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n1085), .A2(KEYINPUT62), .ZN(new_n1086));
  AOI21_X1  g661(.A(new_n987), .B1(new_n1084), .B2(new_n1086), .ZN(new_n1087));
  INV_X1    g662(.A(KEYINPUT63), .ZN(new_n1088));
  NOR2_X1   g663(.A1(new_n1080), .A2(G286), .ZN(new_n1089));
  INV_X1    g664(.A(new_n1089), .ZN(new_n1090));
  OAI21_X1  g665(.A(new_n1088), .B1(new_n987), .B2(new_n1090), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n978), .A2(new_n986), .ZN(new_n1092));
  INV_X1    g667(.A(new_n1092), .ZN(new_n1093));
  AOI21_X1  g668(.A(new_n1088), .B1(new_n950), .B2(new_n952), .ZN(new_n1094));
  NAND4_X1  g669(.A1(new_n1093), .A2(new_n959), .A3(new_n1089), .A4(new_n1094), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n1091), .A2(new_n1095), .ZN(new_n1096));
  NOR2_X1   g671(.A1(G288), .A2(G1976), .ZN(new_n1097));
  XNOR2_X1  g672(.A(new_n1097), .B(KEYINPUT115), .ZN(new_n1098));
  NAND3_X1  g673(.A1(new_n1098), .A2(new_n975), .A3(new_n976), .ZN(new_n1099));
  INV_X1    g674(.A(new_n972), .ZN(new_n1100));
  AOI22_X1  g675(.A1(new_n1099), .A2(new_n1100), .B1(new_n967), .B2(new_n963), .ZN(new_n1101));
  INV_X1    g676(.A(new_n1101), .ZN(new_n1102));
  OAI211_X1 g677(.A(new_n1096), .B(new_n1102), .C1(new_n959), .C2(new_n1092), .ZN(new_n1103));
  OAI211_X1 g678(.A(new_n930), .B(new_n934), .C1(new_n1087), .C2(new_n1103), .ZN(new_n1104));
  INV_X1    g679(.A(new_n1104), .ZN(new_n1105));
  NOR2_X1   g680(.A1(new_n1092), .A2(new_n959), .ZN(new_n1106));
  AOI211_X1 g681(.A(new_n1106), .B(new_n1101), .C1(new_n1091), .C2(new_n1095), .ZN(new_n1107));
  AOI22_X1  g682(.A1(new_n1063), .A2(new_n1083), .B1(new_n1085), .B2(KEYINPUT62), .ZN(new_n1108));
  OAI21_X1  g683(.A(new_n1107), .B1(new_n1108), .B2(new_n987), .ZN(new_n1109));
  AOI21_X1  g684(.A(new_n930), .B1(new_n1109), .B2(new_n934), .ZN(new_n1110));
  OAI21_X1  g685(.A(new_n929), .B1(new_n1105), .B2(new_n1110), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g686(.A1(G227), .A2(new_n459), .ZN(new_n1113));
  XOR2_X1   g687(.A(new_n1113), .B(KEYINPUT126), .Z(new_n1114));
  NAND3_X1  g688(.A1(new_n683), .A2(new_n646), .A3(new_n1114), .ZN(new_n1115));
  INV_X1    g689(.A(KEYINPUT127), .ZN(new_n1116));
  NAND2_X1  g690(.A1(new_n1115), .A2(new_n1116), .ZN(new_n1117));
  NAND4_X1  g691(.A1(new_n683), .A2(new_n646), .A3(KEYINPUT127), .A4(new_n1114), .ZN(new_n1118));
  NAND2_X1  g692(.A1(new_n1117), .A2(new_n1118), .ZN(new_n1119));
  AND3_X1   g693(.A1(new_n1119), .A2(new_n852), .A3(new_n891), .ZN(G308));
  NAND3_X1  g694(.A1(new_n1119), .A2(new_n852), .A3(new_n891), .ZN(G225));
endmodule


