

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598,
         n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609,
         n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620,
         n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631,
         n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642,
         n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653,
         n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664,
         n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675,
         n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686,
         n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697,
         n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708,
         n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719,
         n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730,
         n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741,
         n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752,
         n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, n763,
         n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, n774,
         n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, n785,
         n786, n787, n788, n789, n790, n791, n792, n793, n794, n795, n796,
         n797, n798, n799, n800, n801, n802, n803, n804, n805, n806, n807,
         n808, n809, n810, n811, n812, n813, n814, n815, n816, n817, n818,
         n819, n820, n821, n822, n823, n824, n825, n826, n827, n828, n829,
         n830, n831, n832, n833, n834, n835, n836, n837, n838, n839, n840,
         n841, n842, n843, n844, n845, n846, n847, n848, n849, n850, n851,
         n852, n853, n854, n855, n856, n857, n858, n859, n860, n861, n862,
         n863, n864, n865, n866, n867, n868, n869, n870, n871, n872, n873,
         n874, n875, n876, n877, n878, n879, n880, n881, n882, n883, n884,
         n885, n886, n887, n888, n889, n890, n891, n892, n893, n894, n895,
         n896, n897, n898, n899, n900, n901, n902, n903, n904, n905, n906,
         n907, n908, n909, n910, n911, n912, n913, n914, n915, n916, n917,
         n918, n919, n920, n921, n922, n923, n924, n925, n926, n927, n928,
         n929, n930, n931, n932, n933, n934, n935, n936, n937, n938, n939,
         n940, n941, n942, n943, n944, n945, n946, n947, n948, n949, n950,
         n951, n952, n953, n954, n955, n956, n957, n958, n959, n960, n961,
         n962, n963, n964, n965, n966, n967, n968, n969, n970, n971, n972,
         n973, n974, n975, n976, n977, n978, n979, n980, n981, n982, n983,
         n984, n985, n986, n987, n988, n989, n990, n991, n992, n993, n994,
         n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  AND2_X1 U544 ( .A1(G2105), .A2(n553), .ZN(n863) );
  INV_X1 U545 ( .A(KEYINPUT97), .ZN(n684) );
  XNOR2_X1 U546 ( .A(n685), .B(n684), .ZN(n686) );
  AND2_X1 U547 ( .A1(n753), .A2(n755), .ZN(n707) );
  INV_X1 U548 ( .A(KEYINPUT29), .ZN(n704) );
  XNOR2_X1 U549 ( .A(n705), .B(n704), .ZN(n712) );
  INV_X1 U550 ( .A(KEYINPUT99), .ZN(n725) );
  XNOR2_X1 U551 ( .A(n726), .B(n725), .ZN(n727) );
  OR2_X1 U552 ( .A1(n675), .A2(n674), .ZN(n676) );
  NOR2_X1 U553 ( .A1(n677), .A2(n676), .ZN(n753) );
  NOR2_X2 U554 ( .A1(G2105), .A2(n553), .ZN(n867) );
  NOR2_X1 U555 ( .A1(G651), .A2(n630), .ZN(n638) );
  NOR2_X1 U556 ( .A1(G651), .A2(G543), .ZN(n636) );
  NAND2_X1 U557 ( .A1(G89), .A2(n636), .ZN(n507) );
  XNOR2_X1 U558 ( .A(n507), .B(KEYINPUT80), .ZN(n508) );
  XNOR2_X1 U559 ( .A(n508), .B(KEYINPUT4), .ZN(n511) );
  XOR2_X1 U560 ( .A(G543), .B(KEYINPUT0), .Z(n630) );
  XNOR2_X1 U561 ( .A(KEYINPUT67), .B(G651), .ZN(n513) );
  NOR2_X1 U562 ( .A1(n630), .A2(n513), .ZN(n509) );
  XNOR2_X1 U563 ( .A(KEYINPUT68), .B(n509), .ZN(n637) );
  NAND2_X1 U564 ( .A1(G76), .A2(n637), .ZN(n510) );
  NAND2_X1 U565 ( .A1(n511), .A2(n510), .ZN(n512) );
  XNOR2_X1 U566 ( .A(KEYINPUT5), .B(n512), .ZN(n520) );
  XNOR2_X1 U567 ( .A(KEYINPUT81), .B(KEYINPUT6), .ZN(n518) );
  NAND2_X1 U568 ( .A1(n638), .A2(G51), .ZN(n516) );
  NOR2_X1 U569 ( .A1(G543), .A2(n513), .ZN(n514) );
  XOR2_X1 U570 ( .A(KEYINPUT1), .B(n514), .Z(n641) );
  NAND2_X1 U571 ( .A1(G63), .A2(n641), .ZN(n515) );
  NAND2_X1 U572 ( .A1(n516), .A2(n515), .ZN(n517) );
  XNOR2_X1 U573 ( .A(n518), .B(n517), .ZN(n519) );
  NAND2_X1 U574 ( .A1(n520), .A2(n519), .ZN(n521) );
  XNOR2_X1 U575 ( .A(KEYINPUT7), .B(n521), .ZN(G168) );
  XOR2_X1 U576 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U577 ( .A1(n638), .A2(G52), .ZN(n523) );
  NAND2_X1 U578 ( .A1(G64), .A2(n641), .ZN(n522) );
  NAND2_X1 U579 ( .A1(n523), .A2(n522), .ZN(n530) );
  NAND2_X1 U580 ( .A1(G90), .A2(n636), .ZN(n526) );
  NAND2_X1 U581 ( .A1(n637), .A2(G77), .ZN(n524) );
  XOR2_X1 U582 ( .A(KEYINPUT69), .B(n524), .Z(n525) );
  NAND2_X1 U583 ( .A1(n526), .A2(n525), .ZN(n527) );
  XNOR2_X1 U584 ( .A(n527), .B(KEYINPUT9), .ZN(n528) );
  XOR2_X1 U585 ( .A(KEYINPUT70), .B(n528), .Z(n529) );
  NOR2_X1 U586 ( .A1(n530), .A2(n529), .ZN(G171) );
  NAND2_X1 U587 ( .A1(n636), .A2(G85), .ZN(n532) );
  NAND2_X1 U588 ( .A1(G60), .A2(n641), .ZN(n531) );
  NAND2_X1 U589 ( .A1(n532), .A2(n531), .ZN(n536) );
  NAND2_X1 U590 ( .A1(G72), .A2(n637), .ZN(n534) );
  NAND2_X1 U591 ( .A1(G47), .A2(n638), .ZN(n533) );
  NAND2_X1 U592 ( .A1(n534), .A2(n533), .ZN(n535) );
  OR2_X1 U593 ( .A1(n536), .A2(n535), .ZN(G290) );
  XOR2_X1 U594 ( .A(G2435), .B(G2454), .Z(n538) );
  XNOR2_X1 U595 ( .A(G2430), .B(G2438), .ZN(n537) );
  XNOR2_X1 U596 ( .A(n538), .B(n537), .ZN(n545) );
  XOR2_X1 U597 ( .A(G2446), .B(KEYINPUT105), .Z(n540) );
  XNOR2_X1 U598 ( .A(G2451), .B(G2443), .ZN(n539) );
  XNOR2_X1 U599 ( .A(n540), .B(n539), .ZN(n541) );
  XOR2_X1 U600 ( .A(n541), .B(G2427), .Z(n543) );
  XNOR2_X1 U601 ( .A(G1348), .B(G1341), .ZN(n542) );
  XNOR2_X1 U602 ( .A(n543), .B(n542), .ZN(n544) );
  XNOR2_X1 U603 ( .A(n545), .B(n544), .ZN(n546) );
  AND2_X1 U604 ( .A1(n546), .A2(G14), .ZN(G401) );
  AND2_X1 U605 ( .A1(G2105), .A2(G2104), .ZN(n862) );
  NAND2_X1 U606 ( .A1(G111), .A2(n862), .ZN(n549) );
  NOR2_X1 U607 ( .A1(G2105), .A2(G2104), .ZN(n547) );
  XOR2_X2 U608 ( .A(KEYINPUT17), .B(n547), .Z(n866) );
  NAND2_X1 U609 ( .A1(G135), .A2(n866), .ZN(n548) );
  NAND2_X1 U610 ( .A1(n549), .A2(n548), .ZN(n552) );
  XOR2_X1 U611 ( .A(KEYINPUT64), .B(G2104), .Z(n553) );
  NAND2_X1 U612 ( .A1(n863), .A2(G123), .ZN(n550) );
  XOR2_X1 U613 ( .A(KEYINPUT18), .B(n550), .Z(n551) );
  NOR2_X1 U614 ( .A1(n552), .A2(n551), .ZN(n555) );
  NAND2_X1 U615 ( .A1(n867), .A2(G99), .ZN(n554) );
  NAND2_X1 U616 ( .A1(n555), .A2(n554), .ZN(n976) );
  XNOR2_X1 U617 ( .A(G2096), .B(n976), .ZN(n556) );
  OR2_X1 U618 ( .A1(G2100), .A2(n556), .ZN(G156) );
  INV_X1 U619 ( .A(G82), .ZN(G220) );
  NAND2_X1 U620 ( .A1(G138), .A2(n866), .ZN(n558) );
  NAND2_X1 U621 ( .A1(G102), .A2(n867), .ZN(n557) );
  NAND2_X1 U622 ( .A1(n558), .A2(n557), .ZN(n564) );
  INV_X1 U623 ( .A(KEYINPUT91), .ZN(n562) );
  NAND2_X1 U624 ( .A1(G114), .A2(n862), .ZN(n560) );
  NAND2_X1 U625 ( .A1(G126), .A2(n863), .ZN(n559) );
  NAND2_X1 U626 ( .A1(n560), .A2(n559), .ZN(n561) );
  XNOR2_X1 U627 ( .A(n562), .B(n561), .ZN(n563) );
  NOR2_X1 U628 ( .A1(n564), .A2(n563), .ZN(G164) );
  NAND2_X1 U629 ( .A1(n862), .A2(G113), .ZN(n565) );
  XOR2_X1 U630 ( .A(KEYINPUT65), .B(n565), .Z(n567) );
  NAND2_X1 U631 ( .A1(n866), .A2(G137), .ZN(n566) );
  NAND2_X1 U632 ( .A1(n567), .A2(n566), .ZN(n568) );
  XNOR2_X1 U633 ( .A(n568), .B(KEYINPUT66), .ZN(n570) );
  AND2_X1 U634 ( .A1(n863), .A2(G125), .ZN(n569) );
  OR2_X1 U635 ( .A1(n570), .A2(n569), .ZN(n677) );
  NAND2_X1 U636 ( .A1(G101), .A2(n867), .ZN(n571) );
  XNOR2_X1 U637 ( .A(KEYINPUT23), .B(n571), .ZN(n675) );
  NOR2_X1 U638 ( .A1(n677), .A2(n675), .ZN(G160) );
  NAND2_X1 U639 ( .A1(G94), .A2(G452), .ZN(n572) );
  XNOR2_X1 U640 ( .A(n572), .B(KEYINPUT71), .ZN(G173) );
  NAND2_X1 U641 ( .A1(G7), .A2(G661), .ZN(n573) );
  XNOR2_X1 U642 ( .A(n573), .B(KEYINPUT74), .ZN(n574) );
  XNOR2_X1 U643 ( .A(KEYINPUT10), .B(n574), .ZN(G223) );
  INV_X1 U644 ( .A(G223), .ZN(n811) );
  NAND2_X1 U645 ( .A1(n811), .A2(G567), .ZN(n575) );
  XOR2_X1 U646 ( .A(KEYINPUT11), .B(n575), .Z(G234) );
  NAND2_X1 U647 ( .A1(n641), .A2(G56), .ZN(n576) );
  XOR2_X1 U648 ( .A(KEYINPUT14), .B(n576), .Z(n582) );
  NAND2_X1 U649 ( .A1(n636), .A2(G81), .ZN(n577) );
  XNOR2_X1 U650 ( .A(n577), .B(KEYINPUT12), .ZN(n579) );
  NAND2_X1 U651 ( .A1(G68), .A2(n637), .ZN(n578) );
  NAND2_X1 U652 ( .A1(n579), .A2(n578), .ZN(n580) );
  XOR2_X1 U653 ( .A(KEYINPUT13), .B(n580), .Z(n581) );
  NOR2_X1 U654 ( .A1(n582), .A2(n581), .ZN(n584) );
  NAND2_X1 U655 ( .A1(n638), .A2(G43), .ZN(n583) );
  NAND2_X1 U656 ( .A1(n584), .A2(n583), .ZN(n909) );
  XNOR2_X1 U657 ( .A(G860), .B(KEYINPUT75), .ZN(n605) );
  OR2_X1 U658 ( .A1(n909), .A2(n605), .ZN(G153) );
  XOR2_X1 U659 ( .A(G171), .B(KEYINPUT76), .Z(G301) );
  NAND2_X1 U660 ( .A1(G92), .A2(n636), .ZN(n591) );
  NAND2_X1 U661 ( .A1(G79), .A2(n637), .ZN(n586) );
  NAND2_X1 U662 ( .A1(G54), .A2(n638), .ZN(n585) );
  NAND2_X1 U663 ( .A1(n586), .A2(n585), .ZN(n589) );
  NAND2_X1 U664 ( .A1(n641), .A2(G66), .ZN(n587) );
  XOR2_X1 U665 ( .A(KEYINPUT78), .B(n587), .Z(n588) );
  NOR2_X1 U666 ( .A1(n589), .A2(n588), .ZN(n590) );
  NAND2_X1 U667 ( .A1(n591), .A2(n590), .ZN(n592) );
  XNOR2_X1 U668 ( .A(n592), .B(KEYINPUT15), .ZN(n922) );
  NOR2_X1 U669 ( .A1(n922), .A2(G868), .ZN(n593) );
  XNOR2_X1 U670 ( .A(KEYINPUT79), .B(n593), .ZN(n596) );
  NAND2_X1 U671 ( .A1(G868), .A2(G301), .ZN(n594) );
  XOR2_X1 U672 ( .A(KEYINPUT77), .B(n594), .Z(n595) );
  NAND2_X1 U673 ( .A1(n596), .A2(n595), .ZN(G284) );
  NAND2_X1 U674 ( .A1(G78), .A2(n637), .ZN(n598) );
  NAND2_X1 U675 ( .A1(G53), .A2(n638), .ZN(n597) );
  NAND2_X1 U676 ( .A1(n598), .A2(n597), .ZN(n602) );
  NAND2_X1 U677 ( .A1(n636), .A2(G91), .ZN(n600) );
  NAND2_X1 U678 ( .A1(G65), .A2(n641), .ZN(n599) );
  NAND2_X1 U679 ( .A1(n600), .A2(n599), .ZN(n601) );
  NOR2_X1 U680 ( .A1(n602), .A2(n601), .ZN(n919) );
  INV_X1 U681 ( .A(n919), .ZN(G299) );
  INV_X1 U682 ( .A(G868), .ZN(n656) );
  NOR2_X1 U683 ( .A1(G286), .A2(n656), .ZN(n604) );
  NOR2_X1 U684 ( .A1(G868), .A2(G299), .ZN(n603) );
  NOR2_X1 U685 ( .A1(n604), .A2(n603), .ZN(G297) );
  NAND2_X1 U686 ( .A1(n605), .A2(G559), .ZN(n606) );
  NAND2_X1 U687 ( .A1(n606), .A2(n922), .ZN(n607) );
  XNOR2_X1 U688 ( .A(n607), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U689 ( .A1(G868), .A2(n909), .ZN(n610) );
  NAND2_X1 U690 ( .A1(G868), .A2(n922), .ZN(n608) );
  NOR2_X1 U691 ( .A1(G559), .A2(n608), .ZN(n609) );
  NOR2_X1 U692 ( .A1(n610), .A2(n609), .ZN(G282) );
  NAND2_X1 U693 ( .A1(n637), .A2(G80), .ZN(n612) );
  NAND2_X1 U694 ( .A1(G67), .A2(n641), .ZN(n611) );
  NAND2_X1 U695 ( .A1(n612), .A2(n611), .ZN(n615) );
  NAND2_X1 U696 ( .A1(G93), .A2(n636), .ZN(n613) );
  XNOR2_X1 U697 ( .A(KEYINPUT83), .B(n613), .ZN(n614) );
  NOR2_X1 U698 ( .A1(n615), .A2(n614), .ZN(n617) );
  NAND2_X1 U699 ( .A1(n638), .A2(G55), .ZN(n616) );
  NAND2_X1 U700 ( .A1(n617), .A2(n616), .ZN(n657) );
  XNOR2_X1 U701 ( .A(n909), .B(KEYINPUT82), .ZN(n619) );
  NAND2_X1 U702 ( .A1(n922), .A2(G559), .ZN(n618) );
  XNOR2_X1 U703 ( .A(n619), .B(n618), .ZN(n654) );
  NOR2_X1 U704 ( .A1(n654), .A2(G860), .ZN(n620) );
  XOR2_X1 U705 ( .A(n657), .B(n620), .Z(G145) );
  XOR2_X1 U706 ( .A(KEYINPUT2), .B(KEYINPUT85), .Z(n622) );
  NAND2_X1 U707 ( .A1(G73), .A2(n637), .ZN(n621) );
  XNOR2_X1 U708 ( .A(n622), .B(n621), .ZN(n629) );
  NAND2_X1 U709 ( .A1(n638), .A2(G48), .ZN(n624) );
  NAND2_X1 U710 ( .A1(G61), .A2(n641), .ZN(n623) );
  NAND2_X1 U711 ( .A1(n624), .A2(n623), .ZN(n627) );
  NAND2_X1 U712 ( .A1(n636), .A2(G86), .ZN(n625) );
  XOR2_X1 U713 ( .A(KEYINPUT84), .B(n625), .Z(n626) );
  NOR2_X1 U714 ( .A1(n627), .A2(n626), .ZN(n628) );
  NAND2_X1 U715 ( .A1(n629), .A2(n628), .ZN(G305) );
  NAND2_X1 U716 ( .A1(G87), .A2(n630), .ZN(n632) );
  NAND2_X1 U717 ( .A1(G74), .A2(G651), .ZN(n631) );
  NAND2_X1 U718 ( .A1(n632), .A2(n631), .ZN(n633) );
  NOR2_X1 U719 ( .A1(n641), .A2(n633), .ZN(n635) );
  NAND2_X1 U720 ( .A1(n638), .A2(G49), .ZN(n634) );
  NAND2_X1 U721 ( .A1(n635), .A2(n634), .ZN(G288) );
  NAND2_X1 U722 ( .A1(G88), .A2(n636), .ZN(n646) );
  NAND2_X1 U723 ( .A1(G75), .A2(n637), .ZN(n640) );
  NAND2_X1 U724 ( .A1(G50), .A2(n638), .ZN(n639) );
  NAND2_X1 U725 ( .A1(n640), .A2(n639), .ZN(n644) );
  NAND2_X1 U726 ( .A1(n641), .A2(G62), .ZN(n642) );
  XOR2_X1 U727 ( .A(KEYINPUT86), .B(n642), .Z(n643) );
  NOR2_X1 U728 ( .A1(n644), .A2(n643), .ZN(n645) );
  NAND2_X1 U729 ( .A1(n646), .A2(n645), .ZN(n647) );
  XNOR2_X1 U730 ( .A(n647), .B(KEYINPUT87), .ZN(G166) );
  XOR2_X1 U731 ( .A(G305), .B(G290), .Z(n648) );
  XNOR2_X1 U732 ( .A(n657), .B(n648), .ZN(n651) );
  XOR2_X1 U733 ( .A(KEYINPUT19), .B(KEYINPUT88), .Z(n649) );
  XNOR2_X1 U734 ( .A(G288), .B(n649), .ZN(n650) );
  XOR2_X1 U735 ( .A(n651), .B(n650), .Z(n653) );
  XNOR2_X1 U736 ( .A(n919), .B(G166), .ZN(n652) );
  XNOR2_X1 U737 ( .A(n653), .B(n652), .ZN(n878) );
  XNOR2_X1 U738 ( .A(n654), .B(n878), .ZN(n655) );
  NAND2_X1 U739 ( .A1(n655), .A2(G868), .ZN(n659) );
  NAND2_X1 U740 ( .A1(n657), .A2(n656), .ZN(n658) );
  NAND2_X1 U741 ( .A1(n659), .A2(n658), .ZN(G295) );
  NAND2_X1 U742 ( .A1(G2078), .A2(G2084), .ZN(n660) );
  XNOR2_X1 U743 ( .A(n660), .B(KEYINPUT20), .ZN(n661) );
  XNOR2_X1 U744 ( .A(KEYINPUT89), .B(n661), .ZN(n662) );
  NAND2_X1 U745 ( .A1(n662), .A2(G2090), .ZN(n663) );
  XNOR2_X1 U746 ( .A(KEYINPUT21), .B(n663), .ZN(n664) );
  NAND2_X1 U747 ( .A1(n664), .A2(G2072), .ZN(G158) );
  XOR2_X1 U748 ( .A(KEYINPUT72), .B(G57), .Z(G237) );
  XNOR2_X1 U749 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  XNOR2_X1 U750 ( .A(KEYINPUT73), .B(G132), .ZN(G219) );
  NAND2_X1 U751 ( .A1(G483), .A2(G661), .ZN(n672) );
  NAND2_X1 U752 ( .A1(G108), .A2(G120), .ZN(n665) );
  NOR2_X1 U753 ( .A1(G237), .A2(n665), .ZN(n666) );
  NAND2_X1 U754 ( .A1(G69), .A2(n666), .ZN(n815) );
  NAND2_X1 U755 ( .A1(n815), .A2(G567), .ZN(n671) );
  NOR2_X1 U756 ( .A1(G220), .A2(G219), .ZN(n667) );
  XOR2_X1 U757 ( .A(KEYINPUT22), .B(n667), .Z(n668) );
  NOR2_X1 U758 ( .A1(G218), .A2(n668), .ZN(n669) );
  NAND2_X1 U759 ( .A1(G96), .A2(n669), .ZN(n816) );
  NAND2_X1 U760 ( .A1(n816), .A2(G2106), .ZN(n670) );
  NAND2_X1 U761 ( .A1(n671), .A2(n670), .ZN(n817) );
  NOR2_X1 U762 ( .A1(n672), .A2(n817), .ZN(n673) );
  XNOR2_X1 U763 ( .A(n673), .B(KEYINPUT90), .ZN(n814) );
  NAND2_X1 U764 ( .A1(G36), .A2(n814), .ZN(G176) );
  XOR2_X1 U765 ( .A(KEYINPUT92), .B(G166), .Z(G303) );
  INV_X1 U766 ( .A(G40), .ZN(n674) );
  NOR2_X1 U767 ( .A1(G164), .A2(G1384), .ZN(n755) );
  NAND2_X1 U768 ( .A1(n753), .A2(n755), .ZN(n713) );
  NAND2_X1 U769 ( .A1(G8), .A2(n713), .ZN(n801) );
  NOR2_X1 U770 ( .A1(G1971), .A2(n801), .ZN(n679) );
  NOR2_X1 U771 ( .A1(G2090), .A2(n713), .ZN(n678) );
  NOR2_X1 U772 ( .A1(n679), .A2(n678), .ZN(n680) );
  NAND2_X1 U773 ( .A1(n680), .A2(G303), .ZN(n724) );
  NAND2_X1 U774 ( .A1(n707), .A2(G1996), .ZN(n681) );
  XNOR2_X1 U775 ( .A(n681), .B(KEYINPUT26), .ZN(n683) );
  NAND2_X1 U776 ( .A1(G1341), .A2(n713), .ZN(n682) );
  NAND2_X1 U777 ( .A1(n683), .A2(n682), .ZN(n685) );
  NOR2_X1 U778 ( .A1(n686), .A2(n909), .ZN(n691) );
  NAND2_X1 U779 ( .A1(n691), .A2(n922), .ZN(n690) );
  NOR2_X1 U780 ( .A1(G2067), .A2(n713), .ZN(n688) );
  NOR2_X1 U781 ( .A1(n707), .A2(G1348), .ZN(n687) );
  NOR2_X1 U782 ( .A1(n688), .A2(n687), .ZN(n689) );
  NAND2_X1 U783 ( .A1(n690), .A2(n689), .ZN(n693) );
  OR2_X1 U784 ( .A1(n922), .A2(n691), .ZN(n692) );
  NAND2_X1 U785 ( .A1(n693), .A2(n692), .ZN(n698) );
  NAND2_X1 U786 ( .A1(n707), .A2(G2072), .ZN(n694) );
  XNOR2_X1 U787 ( .A(n694), .B(KEYINPUT27), .ZN(n696) );
  INV_X1 U788 ( .A(G1956), .ZN(n918) );
  NOR2_X1 U789 ( .A1(n918), .A2(n707), .ZN(n695) );
  NOR2_X1 U790 ( .A1(n696), .A2(n695), .ZN(n699) );
  NAND2_X1 U791 ( .A1(n699), .A2(n919), .ZN(n697) );
  NAND2_X1 U792 ( .A1(n698), .A2(n697), .ZN(n703) );
  NOR2_X1 U793 ( .A1(n699), .A2(n919), .ZN(n701) );
  XOR2_X1 U794 ( .A(KEYINPUT96), .B(KEYINPUT28), .Z(n700) );
  XNOR2_X1 U795 ( .A(n701), .B(n700), .ZN(n702) );
  NAND2_X1 U796 ( .A1(n703), .A2(n702), .ZN(n705) );
  XOR2_X1 U797 ( .A(KEYINPUT25), .B(G2078), .Z(n889) );
  NOR2_X1 U798 ( .A1(n889), .A2(n713), .ZN(n706) );
  XNOR2_X1 U799 ( .A(n706), .B(KEYINPUT94), .ZN(n709) );
  NOR2_X1 U800 ( .A1(n707), .A2(G1961), .ZN(n708) );
  NOR2_X1 U801 ( .A1(n709), .A2(n708), .ZN(n710) );
  XNOR2_X1 U802 ( .A(KEYINPUT95), .B(n710), .ZN(n717) );
  NAND2_X1 U803 ( .A1(n717), .A2(G171), .ZN(n711) );
  NAND2_X1 U804 ( .A1(n712), .A2(n711), .ZN(n722) );
  NOR2_X1 U805 ( .A1(G1966), .A2(n801), .ZN(n732) );
  NOR2_X1 U806 ( .A1(G2084), .A2(n713), .ZN(n729) );
  NOR2_X1 U807 ( .A1(n732), .A2(n729), .ZN(n714) );
  NAND2_X1 U808 ( .A1(G8), .A2(n714), .ZN(n715) );
  XNOR2_X1 U809 ( .A(KEYINPUT30), .B(n715), .ZN(n716) );
  NOR2_X1 U810 ( .A1(G168), .A2(n716), .ZN(n719) );
  NOR2_X1 U811 ( .A1(G171), .A2(n717), .ZN(n718) );
  NOR2_X1 U812 ( .A1(n719), .A2(n718), .ZN(n720) );
  XOR2_X1 U813 ( .A(KEYINPUT31), .B(n720), .Z(n721) );
  NAND2_X1 U814 ( .A1(n722), .A2(n721), .ZN(n730) );
  NAND2_X1 U815 ( .A1(n730), .A2(G286), .ZN(n723) );
  NAND2_X1 U816 ( .A1(n724), .A2(n723), .ZN(n726) );
  NAND2_X1 U817 ( .A1(n727), .A2(G8), .ZN(n728) );
  XNOR2_X1 U818 ( .A(n728), .B(KEYINPUT32), .ZN(n736) );
  NAND2_X1 U819 ( .A1(G8), .A2(n729), .ZN(n734) );
  XOR2_X1 U820 ( .A(KEYINPUT98), .B(n730), .Z(n731) );
  NOR2_X1 U821 ( .A1(n732), .A2(n731), .ZN(n733) );
  NAND2_X1 U822 ( .A1(n734), .A2(n733), .ZN(n735) );
  NAND2_X1 U823 ( .A1(n736), .A2(n735), .ZN(n796) );
  NOR2_X1 U824 ( .A1(G2090), .A2(G303), .ZN(n737) );
  NAND2_X1 U825 ( .A1(G8), .A2(n737), .ZN(n738) );
  NAND2_X1 U826 ( .A1(n796), .A2(n738), .ZN(n739) );
  XNOR2_X1 U827 ( .A(n739), .B(KEYINPUT100), .ZN(n740) );
  NAND2_X1 U828 ( .A1(n740), .A2(n801), .ZN(n786) );
  NOR2_X1 U829 ( .A1(G1981), .A2(G305), .ZN(n741) );
  XOR2_X1 U830 ( .A(n741), .B(KEYINPUT24), .Z(n742) );
  NOR2_X1 U831 ( .A1(n801), .A2(n742), .ZN(n784) );
  NAND2_X1 U832 ( .A1(G140), .A2(n866), .ZN(n744) );
  NAND2_X1 U833 ( .A1(G104), .A2(n867), .ZN(n743) );
  NAND2_X1 U834 ( .A1(n744), .A2(n743), .ZN(n746) );
  XOR2_X1 U835 ( .A(KEYINPUT93), .B(KEYINPUT34), .Z(n745) );
  XNOR2_X1 U836 ( .A(n746), .B(n745), .ZN(n751) );
  NAND2_X1 U837 ( .A1(G116), .A2(n862), .ZN(n748) );
  NAND2_X1 U838 ( .A1(G128), .A2(n863), .ZN(n747) );
  NAND2_X1 U839 ( .A1(n748), .A2(n747), .ZN(n749) );
  XOR2_X1 U840 ( .A(KEYINPUT35), .B(n749), .Z(n750) );
  NOR2_X1 U841 ( .A1(n751), .A2(n750), .ZN(n752) );
  XNOR2_X1 U842 ( .A(KEYINPUT36), .B(n752), .ZN(n855) );
  XNOR2_X1 U843 ( .A(G2067), .B(KEYINPUT37), .ZN(n780) );
  NOR2_X1 U844 ( .A1(n855), .A2(n780), .ZN(n984) );
  INV_X1 U845 ( .A(n753), .ZN(n754) );
  NOR2_X1 U846 ( .A1(n755), .A2(n754), .ZN(n788) );
  NAND2_X1 U847 ( .A1(n984), .A2(n788), .ZN(n790) );
  NAND2_X1 U848 ( .A1(G105), .A2(n867), .ZN(n756) );
  XNOR2_X1 U849 ( .A(n756), .B(KEYINPUT38), .ZN(n758) );
  NAND2_X1 U850 ( .A1(n862), .A2(G117), .ZN(n757) );
  NAND2_X1 U851 ( .A1(n758), .A2(n757), .ZN(n762) );
  NAND2_X1 U852 ( .A1(G141), .A2(n866), .ZN(n760) );
  NAND2_X1 U853 ( .A1(G129), .A2(n863), .ZN(n759) );
  NAND2_X1 U854 ( .A1(n760), .A2(n759), .ZN(n761) );
  OR2_X1 U855 ( .A1(n762), .A2(n761), .ZN(n859) );
  NOR2_X1 U856 ( .A1(G1996), .A2(n859), .ZN(n974) );
  NAND2_X1 U857 ( .A1(G107), .A2(n862), .ZN(n764) );
  NAND2_X1 U858 ( .A1(G131), .A2(n866), .ZN(n763) );
  NAND2_X1 U859 ( .A1(n764), .A2(n763), .ZN(n768) );
  NAND2_X1 U860 ( .A1(G95), .A2(n867), .ZN(n766) );
  NAND2_X1 U861 ( .A1(G119), .A2(n863), .ZN(n765) );
  NAND2_X1 U862 ( .A1(n766), .A2(n765), .ZN(n767) );
  OR2_X1 U863 ( .A1(n768), .A2(n767), .ZN(n854) );
  NOR2_X1 U864 ( .A1(G1991), .A2(n854), .ZN(n979) );
  NOR2_X1 U865 ( .A1(G1986), .A2(G290), .ZN(n769) );
  XOR2_X1 U866 ( .A(n769), .B(KEYINPUT101), .Z(n770) );
  NOR2_X1 U867 ( .A1(n979), .A2(n770), .ZN(n774) );
  AND2_X1 U868 ( .A1(n854), .A2(G1991), .ZN(n772) );
  AND2_X1 U869 ( .A1(G1996), .A2(n859), .ZN(n771) );
  NOR2_X1 U870 ( .A1(n772), .A2(n771), .ZN(n986) );
  INV_X1 U871 ( .A(n986), .ZN(n773) );
  NOR2_X1 U872 ( .A1(n774), .A2(n773), .ZN(n775) );
  XNOR2_X1 U873 ( .A(n775), .B(KEYINPUT102), .ZN(n776) );
  NOR2_X1 U874 ( .A1(n974), .A2(n776), .ZN(n777) );
  XOR2_X1 U875 ( .A(n777), .B(KEYINPUT103), .Z(n778) );
  XNOR2_X1 U876 ( .A(KEYINPUT39), .B(n778), .ZN(n779) );
  NAND2_X1 U877 ( .A1(n790), .A2(n779), .ZN(n781) );
  NAND2_X1 U878 ( .A1(n855), .A2(n780), .ZN(n988) );
  NAND2_X1 U879 ( .A1(n781), .A2(n988), .ZN(n782) );
  NAND2_X1 U880 ( .A1(n782), .A2(n788), .ZN(n783) );
  XOR2_X1 U881 ( .A(KEYINPUT104), .B(n783), .Z(n787) );
  NOR2_X1 U882 ( .A1(n784), .A2(n787), .ZN(n785) );
  NAND2_X1 U883 ( .A1(n786), .A2(n785), .ZN(n794) );
  INV_X1 U884 ( .A(n787), .ZN(n793) );
  XOR2_X1 U885 ( .A(G1986), .B(G290), .Z(n923) );
  NAND2_X1 U886 ( .A1(n923), .A2(n986), .ZN(n789) );
  NAND2_X1 U887 ( .A1(n789), .A2(n788), .ZN(n791) );
  NAND2_X1 U888 ( .A1(n791), .A2(n790), .ZN(n792) );
  NAND2_X1 U889 ( .A1(n793), .A2(n792), .ZN(n805) );
  NAND2_X1 U890 ( .A1(n794), .A2(n805), .ZN(n809) );
  NOR2_X1 U891 ( .A1(G1976), .A2(G288), .ZN(n914) );
  NOR2_X1 U892 ( .A1(G303), .A2(G1971), .ZN(n926) );
  NOR2_X1 U893 ( .A1(n914), .A2(n926), .ZN(n795) );
  NAND2_X1 U894 ( .A1(n796), .A2(n795), .ZN(n799) );
  NAND2_X1 U895 ( .A1(G1976), .A2(G288), .ZN(n916) );
  INV_X1 U896 ( .A(n916), .ZN(n797) );
  NOR2_X1 U897 ( .A1(n801), .A2(n797), .ZN(n798) );
  AND2_X1 U898 ( .A1(n799), .A2(n798), .ZN(n800) );
  NOR2_X1 U899 ( .A1(KEYINPUT33), .A2(n800), .ZN(n804) );
  NAND2_X1 U900 ( .A1(n914), .A2(KEYINPUT33), .ZN(n802) );
  NOR2_X1 U901 ( .A1(n802), .A2(n801), .ZN(n803) );
  NOR2_X1 U902 ( .A1(n804), .A2(n803), .ZN(n807) );
  XOR2_X1 U903 ( .A(G1981), .B(G305), .Z(n930) );
  AND2_X1 U904 ( .A1(n930), .A2(n805), .ZN(n806) );
  NAND2_X1 U905 ( .A1(n807), .A2(n806), .ZN(n808) );
  AND2_X1 U906 ( .A1(n809), .A2(n808), .ZN(n810) );
  XOR2_X1 U907 ( .A(KEYINPUT40), .B(n810), .Z(G329) );
  NAND2_X1 U908 ( .A1(G2106), .A2(n811), .ZN(G217) );
  AND2_X1 U909 ( .A1(G15), .A2(G2), .ZN(n812) );
  NAND2_X1 U910 ( .A1(G661), .A2(n812), .ZN(G259) );
  NAND2_X1 U911 ( .A1(G3), .A2(G1), .ZN(n813) );
  NAND2_X1 U912 ( .A1(n814), .A2(n813), .ZN(G188) );
  NOR2_X1 U913 ( .A1(n816), .A2(n815), .ZN(G325) );
  XOR2_X1 U914 ( .A(KEYINPUT106), .B(G325), .Z(G261) );
  INV_X1 U916 ( .A(G120), .ZN(G236) );
  INV_X1 U917 ( .A(G108), .ZN(G238) );
  INV_X1 U918 ( .A(G96), .ZN(G221) );
  INV_X1 U919 ( .A(G69), .ZN(G235) );
  INV_X1 U920 ( .A(n817), .ZN(G319) );
  XOR2_X1 U921 ( .A(G2678), .B(G2090), .Z(n819) );
  XNOR2_X1 U922 ( .A(G2084), .B(G2078), .ZN(n818) );
  XNOR2_X1 U923 ( .A(n819), .B(n818), .ZN(n820) );
  XOR2_X1 U924 ( .A(n820), .B(G2100), .Z(n822) );
  XNOR2_X1 U925 ( .A(G2072), .B(G2067), .ZN(n821) );
  XNOR2_X1 U926 ( .A(n822), .B(n821), .ZN(n826) );
  XOR2_X1 U927 ( .A(G2096), .B(KEYINPUT107), .Z(n824) );
  XNOR2_X1 U928 ( .A(KEYINPUT42), .B(KEYINPUT43), .ZN(n823) );
  XNOR2_X1 U929 ( .A(n824), .B(n823), .ZN(n825) );
  XOR2_X1 U930 ( .A(n826), .B(n825), .Z(G227) );
  XOR2_X1 U931 ( .A(G1971), .B(G1956), .Z(n828) );
  XNOR2_X1 U932 ( .A(G1966), .B(G1961), .ZN(n827) );
  XNOR2_X1 U933 ( .A(n828), .B(n827), .ZN(n829) );
  XOR2_X1 U934 ( .A(n829), .B(G2474), .Z(n831) );
  XNOR2_X1 U935 ( .A(G1996), .B(G1991), .ZN(n830) );
  XNOR2_X1 U936 ( .A(n831), .B(n830), .ZN(n835) );
  XOR2_X1 U937 ( .A(KEYINPUT41), .B(G1986), .Z(n833) );
  XNOR2_X1 U938 ( .A(G1981), .B(G1976), .ZN(n832) );
  XNOR2_X1 U939 ( .A(n833), .B(n832), .ZN(n834) );
  XNOR2_X1 U940 ( .A(n835), .B(n834), .ZN(G229) );
  NAND2_X1 U941 ( .A1(n863), .A2(G124), .ZN(n836) );
  XNOR2_X1 U942 ( .A(n836), .B(KEYINPUT44), .ZN(n838) );
  NAND2_X1 U943 ( .A1(G136), .A2(n866), .ZN(n837) );
  NAND2_X1 U944 ( .A1(n838), .A2(n837), .ZN(n839) );
  XNOR2_X1 U945 ( .A(KEYINPUT108), .B(n839), .ZN(n843) );
  NAND2_X1 U946 ( .A1(G112), .A2(n862), .ZN(n841) );
  NAND2_X1 U947 ( .A1(G100), .A2(n867), .ZN(n840) );
  NAND2_X1 U948 ( .A1(n841), .A2(n840), .ZN(n842) );
  NOR2_X1 U949 ( .A1(n843), .A2(n842), .ZN(G162) );
  NAND2_X1 U950 ( .A1(G139), .A2(n866), .ZN(n845) );
  NAND2_X1 U951 ( .A1(G103), .A2(n867), .ZN(n844) );
  NAND2_X1 U952 ( .A1(n845), .A2(n844), .ZN(n850) );
  NAND2_X1 U953 ( .A1(G115), .A2(n862), .ZN(n847) );
  NAND2_X1 U954 ( .A1(G127), .A2(n863), .ZN(n846) );
  NAND2_X1 U955 ( .A1(n847), .A2(n846), .ZN(n848) );
  XOR2_X1 U956 ( .A(KEYINPUT47), .B(n848), .Z(n849) );
  NOR2_X1 U957 ( .A1(n850), .A2(n849), .ZN(n969) );
  XOR2_X1 U958 ( .A(KEYINPUT46), .B(KEYINPUT48), .Z(n852) );
  XNOR2_X1 U959 ( .A(KEYINPUT109), .B(KEYINPUT110), .ZN(n851) );
  XNOR2_X1 U960 ( .A(n852), .B(n851), .ZN(n853) );
  XNOR2_X1 U961 ( .A(n969), .B(n853), .ZN(n857) );
  XOR2_X1 U962 ( .A(n855), .B(n854), .Z(n856) );
  XNOR2_X1 U963 ( .A(n857), .B(n856), .ZN(n858) );
  XNOR2_X1 U964 ( .A(n976), .B(n858), .ZN(n861) );
  XOR2_X1 U965 ( .A(G160), .B(n859), .Z(n860) );
  XNOR2_X1 U966 ( .A(n861), .B(n860), .ZN(n874) );
  NAND2_X1 U967 ( .A1(G118), .A2(n862), .ZN(n865) );
  NAND2_X1 U968 ( .A1(G130), .A2(n863), .ZN(n864) );
  NAND2_X1 U969 ( .A1(n865), .A2(n864), .ZN(n872) );
  NAND2_X1 U970 ( .A1(G142), .A2(n866), .ZN(n869) );
  NAND2_X1 U971 ( .A1(G106), .A2(n867), .ZN(n868) );
  NAND2_X1 U972 ( .A1(n869), .A2(n868), .ZN(n870) );
  XOR2_X1 U973 ( .A(KEYINPUT45), .B(n870), .Z(n871) );
  NOR2_X1 U974 ( .A1(n872), .A2(n871), .ZN(n873) );
  XOR2_X1 U975 ( .A(n874), .B(n873), .Z(n876) );
  XNOR2_X1 U976 ( .A(G164), .B(G162), .ZN(n875) );
  XNOR2_X1 U977 ( .A(n876), .B(n875), .ZN(n877) );
  NOR2_X1 U978 ( .A1(G37), .A2(n877), .ZN(G395) );
  XNOR2_X1 U979 ( .A(n909), .B(n878), .ZN(n880) );
  XNOR2_X1 U980 ( .A(G171), .B(n922), .ZN(n879) );
  XNOR2_X1 U981 ( .A(n880), .B(n879), .ZN(n881) );
  XOR2_X1 U982 ( .A(G286), .B(n881), .Z(n882) );
  NOR2_X1 U983 ( .A1(G37), .A2(n882), .ZN(G397) );
  NOR2_X1 U984 ( .A1(G227), .A2(G229), .ZN(n883) );
  XNOR2_X1 U985 ( .A(n883), .B(KEYINPUT49), .ZN(n884) );
  NOR2_X1 U986 ( .A1(G401), .A2(n884), .ZN(n885) );
  NAND2_X1 U987 ( .A1(G319), .A2(n885), .ZN(n886) );
  XNOR2_X1 U988 ( .A(KEYINPUT111), .B(n886), .ZN(n888) );
  NOR2_X1 U989 ( .A1(G395), .A2(G397), .ZN(n887) );
  NAND2_X1 U990 ( .A1(n888), .A2(n887), .ZN(G225) );
  INV_X1 U991 ( .A(G225), .ZN(G308) );
  XNOR2_X1 U992 ( .A(G27), .B(n889), .ZN(n890) );
  XNOR2_X1 U993 ( .A(n890), .B(KEYINPUT117), .ZN(n900) );
  XOR2_X1 U994 ( .A(G1991), .B(G25), .Z(n891) );
  NAND2_X1 U995 ( .A1(n891), .A2(G28), .ZN(n892) );
  XNOR2_X1 U996 ( .A(n892), .B(KEYINPUT116), .ZN(n898) );
  XOR2_X1 U997 ( .A(G32), .B(G1996), .Z(n896) );
  XNOR2_X1 U998 ( .A(G2072), .B(G33), .ZN(n894) );
  XNOR2_X1 U999 ( .A(G2067), .B(G26), .ZN(n893) );
  NOR2_X1 U1000 ( .A1(n894), .A2(n893), .ZN(n895) );
  NAND2_X1 U1001 ( .A1(n896), .A2(n895), .ZN(n897) );
  NOR2_X1 U1002 ( .A1(n898), .A2(n897), .ZN(n899) );
  NAND2_X1 U1003 ( .A1(n900), .A2(n899), .ZN(n901) );
  XNOR2_X1 U1004 ( .A(KEYINPUT53), .B(n901), .ZN(n905) );
  XOR2_X1 U1005 ( .A(KEYINPUT118), .B(G34), .Z(n903) );
  XNOR2_X1 U1006 ( .A(G2084), .B(KEYINPUT54), .ZN(n902) );
  XNOR2_X1 U1007 ( .A(n903), .B(n902), .ZN(n904) );
  NAND2_X1 U1008 ( .A1(n905), .A2(n904), .ZN(n907) );
  XNOR2_X1 U1009 ( .A(G35), .B(G2090), .ZN(n906) );
  NOR2_X1 U1010 ( .A1(n907), .A2(n906), .ZN(n1002) );
  NAND2_X1 U1011 ( .A1(KEYINPUT55), .A2(n1002), .ZN(n908) );
  NAND2_X1 U1012 ( .A1(G11), .A2(n908), .ZN(n1001) );
  XNOR2_X1 U1013 ( .A(G16), .B(KEYINPUT56), .ZN(n938) );
  NAND2_X1 U1014 ( .A1(G303), .A2(G1971), .ZN(n911) );
  XOR2_X1 U1015 ( .A(G1341), .B(n909), .Z(n910) );
  NAND2_X1 U1016 ( .A1(n911), .A2(n910), .ZN(n913) );
  XOR2_X1 U1017 ( .A(G171), .B(G1961), .Z(n912) );
  NOR2_X1 U1018 ( .A1(n913), .A2(n912), .ZN(n936) );
  INV_X1 U1019 ( .A(n914), .ZN(n915) );
  NAND2_X1 U1020 ( .A1(n916), .A2(n915), .ZN(n917) );
  XNOR2_X1 U1021 ( .A(n917), .B(KEYINPUT120), .ZN(n921) );
  XNOR2_X1 U1022 ( .A(n919), .B(n918), .ZN(n920) );
  NOR2_X1 U1023 ( .A1(n921), .A2(n920), .ZN(n928) );
  XNOR2_X1 U1024 ( .A(G1348), .B(n922), .ZN(n924) );
  NAND2_X1 U1025 ( .A1(n924), .A2(n923), .ZN(n925) );
  NOR2_X1 U1026 ( .A1(n926), .A2(n925), .ZN(n927) );
  NAND2_X1 U1027 ( .A1(n928), .A2(n927), .ZN(n934) );
  XOR2_X1 U1028 ( .A(G1966), .B(G168), .Z(n929) );
  XNOR2_X1 U1029 ( .A(KEYINPUT119), .B(n929), .ZN(n931) );
  NAND2_X1 U1030 ( .A1(n931), .A2(n930), .ZN(n932) );
  XOR2_X1 U1031 ( .A(KEYINPUT57), .B(n932), .Z(n933) );
  NOR2_X1 U1032 ( .A1(n934), .A2(n933), .ZN(n935) );
  NAND2_X1 U1033 ( .A1(n936), .A2(n935), .ZN(n937) );
  NAND2_X1 U1034 ( .A1(n938), .A2(n937), .ZN(n967) );
  XOR2_X1 U1035 ( .A(G1986), .B(G24), .Z(n941) );
  XNOR2_X1 U1036 ( .A(G1971), .B(KEYINPUT125), .ZN(n939) );
  XNOR2_X1 U1037 ( .A(n939), .B(G22), .ZN(n940) );
  NAND2_X1 U1038 ( .A1(n941), .A2(n940), .ZN(n943) );
  XNOR2_X1 U1039 ( .A(G23), .B(G1976), .ZN(n942) );
  NOR2_X1 U1040 ( .A1(n943), .A2(n942), .ZN(n944) );
  XOR2_X1 U1041 ( .A(KEYINPUT58), .B(n944), .Z(n962) );
  XOR2_X1 U1042 ( .A(G1961), .B(G5), .Z(n947) );
  XNOR2_X1 U1043 ( .A(G1966), .B(G21), .ZN(n945) );
  XNOR2_X1 U1044 ( .A(n945), .B(KEYINPUT123), .ZN(n946) );
  NAND2_X1 U1045 ( .A1(n947), .A2(n946), .ZN(n959) );
  XNOR2_X1 U1046 ( .A(KEYINPUT59), .B(G4), .ZN(n948) );
  XNOR2_X1 U1047 ( .A(n948), .B(KEYINPUT121), .ZN(n949) );
  XNOR2_X1 U1048 ( .A(G1348), .B(n949), .ZN(n951) );
  XNOR2_X1 U1049 ( .A(G1341), .B(G19), .ZN(n950) );
  NOR2_X1 U1050 ( .A1(n951), .A2(n950), .ZN(n955) );
  XNOR2_X1 U1051 ( .A(G1956), .B(G20), .ZN(n953) );
  XNOR2_X1 U1052 ( .A(G1981), .B(G6), .ZN(n952) );
  NOR2_X1 U1053 ( .A1(n953), .A2(n952), .ZN(n954) );
  NAND2_X1 U1054 ( .A1(n955), .A2(n954), .ZN(n956) );
  XNOR2_X1 U1055 ( .A(n956), .B(KEYINPUT60), .ZN(n957) );
  XNOR2_X1 U1056 ( .A(n957), .B(KEYINPUT122), .ZN(n958) );
  NOR2_X1 U1057 ( .A1(n959), .A2(n958), .ZN(n960) );
  XOR2_X1 U1058 ( .A(KEYINPUT124), .B(n960), .Z(n961) );
  NOR2_X1 U1059 ( .A1(n962), .A2(n961), .ZN(n963) );
  XOR2_X1 U1060 ( .A(KEYINPUT61), .B(n963), .Z(n964) );
  NOR2_X1 U1061 ( .A1(G16), .A2(n964), .ZN(n965) );
  XOR2_X1 U1062 ( .A(KEYINPUT126), .B(n965), .Z(n966) );
  NAND2_X1 U1063 ( .A1(n967), .A2(n966), .ZN(n968) );
  XNOR2_X1 U1064 ( .A(n968), .B(KEYINPUT127), .ZN(n999) );
  XOR2_X1 U1065 ( .A(G2072), .B(n969), .Z(n971) );
  XOR2_X1 U1066 ( .A(G164), .B(G2078), .Z(n970) );
  NOR2_X1 U1067 ( .A1(n971), .A2(n970), .ZN(n972) );
  XNOR2_X1 U1068 ( .A(KEYINPUT50), .B(n972), .ZN(n992) );
  XOR2_X1 U1069 ( .A(G2090), .B(G162), .Z(n973) );
  NOR2_X1 U1070 ( .A1(n974), .A2(n973), .ZN(n975) );
  XOR2_X1 U1071 ( .A(KEYINPUT51), .B(n975), .Z(n982) );
  XNOR2_X1 U1072 ( .A(G160), .B(G2084), .ZN(n977) );
  NAND2_X1 U1073 ( .A1(n977), .A2(n976), .ZN(n978) );
  NOR2_X1 U1074 ( .A1(n979), .A2(n978), .ZN(n980) );
  XNOR2_X1 U1075 ( .A(n980), .B(KEYINPUT112), .ZN(n981) );
  NAND2_X1 U1076 ( .A1(n982), .A2(n981), .ZN(n983) );
  NOR2_X1 U1077 ( .A1(n984), .A2(n983), .ZN(n985) );
  NAND2_X1 U1078 ( .A1(n986), .A2(n985), .ZN(n987) );
  XNOR2_X1 U1079 ( .A(n987), .B(KEYINPUT113), .ZN(n989) );
  NAND2_X1 U1080 ( .A1(n989), .A2(n988), .ZN(n990) );
  XOR2_X1 U1081 ( .A(KEYINPUT114), .B(n990), .Z(n991) );
  NAND2_X1 U1082 ( .A1(n992), .A2(n991), .ZN(n993) );
  XNOR2_X1 U1083 ( .A(n993), .B(KEYINPUT115), .ZN(n994) );
  XNOR2_X1 U1084 ( .A(KEYINPUT52), .B(n994), .ZN(n996) );
  INV_X1 U1085 ( .A(KEYINPUT55), .ZN(n995) );
  NAND2_X1 U1086 ( .A1(n996), .A2(n995), .ZN(n997) );
  NAND2_X1 U1087 ( .A1(n997), .A2(G29), .ZN(n998) );
  NAND2_X1 U1088 ( .A1(n999), .A2(n998), .ZN(n1000) );
  NOR2_X1 U1089 ( .A1(n1001), .A2(n1000), .ZN(n1006) );
  INV_X1 U1090 ( .A(n1002), .ZN(n1004) );
  NOR2_X1 U1091 ( .A1(G29), .A2(KEYINPUT55), .ZN(n1003) );
  NAND2_X1 U1092 ( .A1(n1004), .A2(n1003), .ZN(n1005) );
  NAND2_X1 U1093 ( .A1(n1006), .A2(n1005), .ZN(n1007) );
  XOR2_X1 U1094 ( .A(KEYINPUT62), .B(n1007), .Z(G311) );
  INV_X1 U1095 ( .A(G311), .ZN(G150) );
endmodule

