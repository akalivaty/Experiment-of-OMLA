//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 1 0 1 1 0 1 1 0 1 0 0 1 1 1 1 1 0 1 1 0 1 1 0 1 0 0 0 0 0 0 1 1 1 1 1 0 0 1 0 0 0 1 1 1 0 0 1 1 1 1 0 0 1 1 1 0 0 1 0 0 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:23:10 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n716, new_n717,
    new_n718, new_n719, new_n720, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n729, new_n731, new_n732, new_n734, new_n735,
    new_n736, new_n737, new_n738, new_n739, new_n740, new_n742, new_n743,
    new_n744, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n755, new_n756, new_n757, new_n758, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n790, new_n791, new_n792, new_n793, new_n794, new_n795, new_n796,
    new_n797, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n912, new_n913, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n937, new_n938, new_n939, new_n940, new_n941,
    new_n942, new_n943, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n951, new_n952, new_n954, new_n955, new_n956, new_n957,
    new_n958, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1021;
  XNOR2_X1  g000(.A(KEYINPUT9), .B(G234), .ZN(new_n187));
  OAI21_X1  g001(.A(G221), .B1(new_n187), .B2(G902), .ZN(new_n188));
  XNOR2_X1  g002(.A(new_n188), .B(KEYINPUT76), .ZN(new_n189));
  INV_X1    g003(.A(G902), .ZN(new_n190));
  XNOR2_X1  g004(.A(G110), .B(G140), .ZN(new_n191));
  INV_X1    g005(.A(G953), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n192), .A2(G227), .ZN(new_n193));
  XOR2_X1   g007(.A(new_n191), .B(new_n193), .Z(new_n194));
  INV_X1    g008(.A(new_n194), .ZN(new_n195));
  INV_X1    g009(.A(G146), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n196), .A2(G143), .ZN(new_n197));
  INV_X1    g011(.A(G143), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n198), .A2(G146), .ZN(new_n199));
  NAND4_X1  g013(.A1(new_n197), .A2(new_n199), .A3(KEYINPUT0), .A4(G128), .ZN(new_n200));
  XNOR2_X1  g014(.A(G143), .B(G146), .ZN(new_n201));
  XNOR2_X1  g015(.A(KEYINPUT0), .B(G128), .ZN(new_n202));
  OAI21_X1  g016(.A(new_n200), .B1(new_n201), .B2(new_n202), .ZN(new_n203));
  INV_X1    g017(.A(new_n203), .ZN(new_n204));
  INV_X1    g018(.A(KEYINPUT4), .ZN(new_n205));
  INV_X1    g019(.A(KEYINPUT77), .ZN(new_n206));
  INV_X1    g020(.A(G104), .ZN(new_n207));
  OAI22_X1  g021(.A1(new_n206), .A2(KEYINPUT3), .B1(new_n207), .B2(G107), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n207), .A2(G107), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  INV_X1    g024(.A(G107), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n211), .A2(G104), .ZN(new_n212));
  INV_X1    g026(.A(KEYINPUT3), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n213), .A2(KEYINPUT77), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n206), .A2(KEYINPUT3), .ZN(new_n215));
  AOI21_X1  g029(.A(new_n212), .B1(new_n214), .B2(new_n215), .ZN(new_n216));
  OAI211_X1 g030(.A(new_n205), .B(G101), .C1(new_n210), .C2(new_n216), .ZN(new_n217));
  NOR2_X1   g031(.A1(new_n211), .A2(G104), .ZN(new_n218));
  AOI21_X1  g032(.A(new_n218), .B1(new_n212), .B2(new_n214), .ZN(new_n219));
  NOR2_X1   g033(.A1(new_n207), .A2(G107), .ZN(new_n220));
  NOR2_X1   g034(.A1(new_n206), .A2(KEYINPUT3), .ZN(new_n221));
  NOR2_X1   g035(.A1(new_n213), .A2(KEYINPUT77), .ZN(new_n222));
  OAI21_X1  g036(.A(new_n220), .B1(new_n221), .B2(new_n222), .ZN(new_n223));
  INV_X1    g037(.A(G101), .ZN(new_n224));
  NAND3_X1  g038(.A1(new_n219), .A2(new_n223), .A3(new_n224), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n225), .A2(KEYINPUT4), .ZN(new_n226));
  AOI21_X1  g040(.A(new_n224), .B1(new_n219), .B2(new_n223), .ZN(new_n227));
  OAI211_X1 g041(.A(new_n204), .B(new_n217), .C1(new_n226), .C2(new_n227), .ZN(new_n228));
  INV_X1    g042(.A(G128), .ZN(new_n229));
  OAI211_X1 g043(.A(new_n197), .B(new_n199), .C1(KEYINPUT1), .C2(new_n229), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n197), .A2(new_n199), .ZN(new_n231));
  OAI21_X1  g045(.A(KEYINPUT1), .B1(new_n198), .B2(G146), .ZN(new_n232));
  NAND3_X1  g046(.A1(new_n231), .A2(G128), .A3(new_n232), .ZN(new_n233));
  AOI21_X1  g047(.A(new_n224), .B1(new_n212), .B2(new_n209), .ZN(new_n234));
  INV_X1    g048(.A(new_n234), .ZN(new_n235));
  NAND4_X1  g049(.A1(new_n225), .A2(new_n230), .A3(new_n233), .A4(new_n235), .ZN(new_n236));
  XOR2_X1   g050(.A(KEYINPUT78), .B(KEYINPUT10), .Z(new_n237));
  NAND2_X1  g051(.A1(new_n236), .A2(new_n237), .ZN(new_n238));
  INV_X1    g052(.A(KEYINPUT11), .ZN(new_n239));
  NOR2_X1   g053(.A1(new_n239), .A2(KEYINPUT65), .ZN(new_n240));
  INV_X1    g054(.A(G134), .ZN(new_n241));
  NOR2_X1   g055(.A1(new_n241), .A2(G137), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n239), .A2(KEYINPUT65), .ZN(new_n243));
  AOI21_X1  g057(.A(new_n240), .B1(new_n242), .B2(new_n243), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n241), .A2(G137), .ZN(new_n245));
  INV_X1    g059(.A(KEYINPUT65), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n246), .A2(KEYINPUT11), .ZN(new_n247));
  INV_X1    g061(.A(G137), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n248), .A2(G134), .ZN(new_n249));
  OAI21_X1  g063(.A(new_n245), .B1(new_n247), .B2(new_n249), .ZN(new_n250));
  OAI21_X1  g064(.A(G131), .B1(new_n244), .B2(new_n250), .ZN(new_n251));
  NOR2_X1   g065(.A1(new_n248), .A2(G134), .ZN(new_n252));
  AOI21_X1  g066(.A(new_n252), .B1(new_n240), .B2(new_n242), .ZN(new_n253));
  INV_X1    g067(.A(G131), .ZN(new_n254));
  NOR2_X1   g068(.A1(new_n246), .A2(KEYINPUT11), .ZN(new_n255));
  OAI21_X1  g069(.A(new_n247), .B1(new_n255), .B2(new_n249), .ZN(new_n256));
  NAND3_X1  g070(.A1(new_n253), .A2(new_n254), .A3(new_n256), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n251), .A2(new_n257), .ZN(new_n258));
  INV_X1    g072(.A(new_n258), .ZN(new_n259));
  AND2_X1   g073(.A1(new_n233), .A2(new_n230), .ZN(new_n260));
  NAND4_X1  g074(.A1(new_n260), .A2(KEYINPUT10), .A3(new_n225), .A4(new_n235), .ZN(new_n261));
  NAND4_X1  g075(.A1(new_n228), .A2(new_n238), .A3(new_n259), .A4(new_n261), .ZN(new_n262));
  INV_X1    g076(.A(KEYINPUT79), .ZN(new_n263));
  AND2_X1   g077(.A1(new_n263), .A2(KEYINPUT12), .ZN(new_n264));
  NOR2_X1   g078(.A1(new_n264), .A2(KEYINPUT12), .ZN(new_n265));
  INV_X1    g079(.A(new_n265), .ZN(new_n266));
  AOI21_X1  g080(.A(new_n263), .B1(new_n251), .B2(new_n257), .ZN(new_n267));
  NOR3_X1   g081(.A1(new_n210), .A2(new_n216), .A3(G101), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n233), .A2(new_n230), .ZN(new_n269));
  NOR3_X1   g083(.A1(new_n268), .A2(new_n269), .A3(new_n234), .ZN(new_n270));
  AOI22_X1  g084(.A1(new_n225), .A2(new_n235), .B1(new_n230), .B2(new_n233), .ZN(new_n271));
  OAI211_X1 g085(.A(new_n266), .B(new_n267), .C1(new_n270), .C2(new_n271), .ZN(new_n272));
  INV_X1    g086(.A(new_n272), .ZN(new_n273));
  OAI21_X1  g087(.A(new_n269), .B1(new_n268), .B2(new_n234), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n274), .A2(new_n236), .ZN(new_n275));
  AOI21_X1  g089(.A(new_n266), .B1(new_n275), .B2(new_n267), .ZN(new_n276));
  OAI21_X1  g090(.A(new_n262), .B1(new_n273), .B2(new_n276), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n277), .A2(KEYINPUT80), .ZN(new_n278));
  INV_X1    g092(.A(KEYINPUT80), .ZN(new_n279));
  OAI211_X1 g093(.A(new_n279), .B(new_n262), .C1(new_n273), .C2(new_n276), .ZN(new_n280));
  AOI21_X1  g094(.A(new_n195), .B1(new_n278), .B2(new_n280), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n262), .A2(new_n195), .ZN(new_n282));
  NAND3_X1  g096(.A1(new_n228), .A2(new_n238), .A3(new_n261), .ZN(new_n283));
  AOI21_X1  g097(.A(new_n282), .B1(new_n258), .B2(new_n283), .ZN(new_n284));
  OAI21_X1  g098(.A(new_n190), .B1(new_n281), .B2(new_n284), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n285), .A2(G469), .ZN(new_n286));
  INV_X1    g100(.A(G469), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n275), .A2(new_n267), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n288), .A2(new_n265), .ZN(new_n289));
  AOI21_X1  g103(.A(new_n282), .B1(new_n272), .B2(new_n289), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n283), .A2(new_n258), .ZN(new_n291));
  AOI21_X1  g105(.A(new_n195), .B1(new_n291), .B2(new_n262), .ZN(new_n292));
  OAI211_X1 g106(.A(new_n287), .B(new_n190), .C1(new_n290), .C2(new_n292), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n293), .A2(KEYINPUT81), .ZN(new_n294));
  OAI211_X1 g108(.A(new_n195), .B(new_n262), .C1(new_n273), .C2(new_n276), .ZN(new_n295));
  AND2_X1   g109(.A1(new_n291), .A2(new_n262), .ZN(new_n296));
  OAI21_X1  g110(.A(new_n295), .B1(new_n296), .B2(new_n195), .ZN(new_n297));
  INV_X1    g111(.A(KEYINPUT81), .ZN(new_n298));
  NAND4_X1  g112(.A1(new_n297), .A2(new_n298), .A3(new_n287), .A4(new_n190), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n294), .A2(new_n299), .ZN(new_n300));
  AOI21_X1  g114(.A(new_n189), .B1(new_n286), .B2(new_n300), .ZN(new_n301));
  INV_X1    g115(.A(G140), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n302), .A2(G125), .ZN(new_n303));
  INV_X1    g117(.A(G125), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n304), .A2(G140), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n303), .A2(new_n305), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n306), .A2(G146), .ZN(new_n307));
  NAND3_X1  g121(.A1(new_n303), .A2(new_n305), .A3(new_n196), .ZN(new_n308));
  INV_X1    g122(.A(KEYINPUT87), .ZN(new_n309));
  AND3_X1   g123(.A1(new_n307), .A2(new_n308), .A3(new_n309), .ZN(new_n310));
  AOI21_X1  g124(.A(new_n309), .B1(new_n307), .B2(new_n308), .ZN(new_n311));
  INV_X1    g125(.A(G237), .ZN(new_n312));
  NAND3_X1  g126(.A1(new_n312), .A2(new_n192), .A3(G214), .ZN(new_n313));
  INV_X1    g127(.A(KEYINPUT86), .ZN(new_n314));
  NOR2_X1   g128(.A1(new_n314), .A2(G143), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n313), .A2(new_n315), .ZN(new_n316));
  NOR2_X1   g130(.A1(G237), .A2(G953), .ZN(new_n317));
  OAI211_X1 g131(.A(new_n317), .B(G214), .C1(new_n314), .C2(G143), .ZN(new_n318));
  AND4_X1   g132(.A1(KEYINPUT18), .A2(new_n316), .A3(new_n318), .A4(G131), .ZN(new_n319));
  AOI22_X1  g133(.A1(new_n316), .A2(new_n318), .B1(KEYINPUT18), .B2(G131), .ZN(new_n320));
  OAI22_X1  g134(.A1(new_n310), .A2(new_n311), .B1(new_n319), .B2(new_n320), .ZN(new_n321));
  AND3_X1   g135(.A1(new_n303), .A2(new_n305), .A3(KEYINPUT19), .ZN(new_n322));
  AOI21_X1  g136(.A(KEYINPUT19), .B1(new_n303), .B2(new_n305), .ZN(new_n323));
  NOR2_X1   g137(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  OAI21_X1  g138(.A(KEYINPUT88), .B1(new_n324), .B2(G146), .ZN(new_n325));
  INV_X1    g139(.A(KEYINPUT88), .ZN(new_n326));
  OAI211_X1 g140(.A(new_n326), .B(new_n196), .C1(new_n322), .C2(new_n323), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n325), .A2(new_n327), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n316), .A2(new_n318), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n329), .A2(G131), .ZN(new_n330));
  NAND3_X1  g144(.A1(new_n316), .A2(new_n318), .A3(new_n254), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n330), .A2(new_n331), .ZN(new_n332));
  NAND3_X1  g146(.A1(new_n303), .A2(new_n305), .A3(KEYINPUT16), .ZN(new_n333));
  OR3_X1    g147(.A1(new_n304), .A2(KEYINPUT16), .A3(G140), .ZN(new_n334));
  NAND3_X1  g148(.A1(new_n333), .A2(new_n334), .A3(G146), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n332), .A2(new_n335), .ZN(new_n336));
  OAI21_X1  g150(.A(new_n321), .B1(new_n328), .B2(new_n336), .ZN(new_n337));
  XNOR2_X1  g151(.A(G113), .B(G122), .ZN(new_n338));
  XNOR2_X1  g152(.A(new_n338), .B(new_n207), .ZN(new_n339));
  INV_X1    g153(.A(new_n339), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n337), .A2(new_n340), .ZN(new_n341));
  INV_X1    g155(.A(new_n335), .ZN(new_n342));
  AOI21_X1  g156(.A(G146), .B1(new_n333), .B2(new_n334), .ZN(new_n343));
  OAI21_X1  g157(.A(KEYINPUT89), .B1(new_n342), .B2(new_n343), .ZN(new_n344));
  INV_X1    g158(.A(new_n343), .ZN(new_n345));
  INV_X1    g159(.A(KEYINPUT89), .ZN(new_n346));
  NAND3_X1  g160(.A1(new_n345), .A2(new_n346), .A3(new_n335), .ZN(new_n347));
  INV_X1    g161(.A(KEYINPUT17), .ZN(new_n348));
  NAND3_X1  g162(.A1(new_n330), .A2(new_n348), .A3(new_n331), .ZN(new_n349));
  NAND3_X1  g163(.A1(new_n329), .A2(KEYINPUT17), .A3(G131), .ZN(new_n350));
  NAND4_X1  g164(.A1(new_n344), .A2(new_n347), .A3(new_n349), .A4(new_n350), .ZN(new_n351));
  NAND3_X1  g165(.A1(new_n351), .A2(new_n339), .A3(new_n321), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n341), .A2(new_n352), .ZN(new_n353));
  INV_X1    g167(.A(KEYINPUT20), .ZN(new_n354));
  NOR2_X1   g168(.A1(G475), .A2(G902), .ZN(new_n355));
  NAND3_X1  g169(.A1(new_n353), .A2(new_n354), .A3(new_n355), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n356), .A2(KEYINPUT90), .ZN(new_n357));
  INV_X1    g171(.A(KEYINPUT90), .ZN(new_n358));
  NAND4_X1  g172(.A1(new_n353), .A2(new_n358), .A3(new_n354), .A4(new_n355), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n353), .A2(new_n355), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n360), .A2(KEYINPUT20), .ZN(new_n361));
  NAND3_X1  g175(.A1(new_n357), .A2(new_n359), .A3(new_n361), .ZN(new_n362));
  AND3_X1   g176(.A1(new_n351), .A2(new_n339), .A3(new_n321), .ZN(new_n363));
  AOI21_X1  g177(.A(new_n339), .B1(new_n351), .B2(new_n321), .ZN(new_n364));
  OAI21_X1  g178(.A(new_n190), .B1(new_n363), .B2(new_n364), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n365), .A2(G475), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n362), .A2(new_n366), .ZN(new_n367));
  INV_X1    g181(.A(G122), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n368), .A2(G116), .ZN(new_n369));
  INV_X1    g183(.A(G116), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n370), .A2(G122), .ZN(new_n371));
  NAND3_X1  g185(.A1(new_n369), .A2(new_n371), .A3(new_n211), .ZN(new_n372));
  XNOR2_X1  g186(.A(G128), .B(G143), .ZN(new_n373));
  OAI21_X1  g187(.A(new_n372), .B1(new_n373), .B2(G134), .ZN(new_n374));
  AOI21_X1  g188(.A(new_n374), .B1(G134), .B2(new_n373), .ZN(new_n375));
  INV_X1    g189(.A(KEYINPUT94), .ZN(new_n376));
  INV_X1    g190(.A(KEYINPUT93), .ZN(new_n377));
  NOR2_X1   g191(.A1(new_n368), .A2(G116), .ZN(new_n378));
  INV_X1    g192(.A(KEYINPUT14), .ZN(new_n379));
  OAI21_X1  g193(.A(new_n377), .B1(new_n378), .B2(new_n379), .ZN(new_n380));
  OAI211_X1 g194(.A(KEYINPUT93), .B(KEYINPUT14), .C1(new_n368), .C2(G116), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n380), .A2(new_n381), .ZN(new_n382));
  NOR2_X1   g196(.A1(new_n370), .A2(G122), .ZN(new_n383));
  AOI21_X1  g197(.A(new_n383), .B1(new_n379), .B2(new_n378), .ZN(new_n384));
  AOI211_X1 g198(.A(new_n376), .B(new_n211), .C1(new_n382), .C2(new_n384), .ZN(new_n385));
  AOI21_X1  g199(.A(KEYINPUT93), .B1(new_n371), .B2(KEYINPUT14), .ZN(new_n386));
  INV_X1    g200(.A(new_n381), .ZN(new_n387));
  OAI21_X1  g201(.A(new_n384), .B1(new_n386), .B2(new_n387), .ZN(new_n388));
  AOI21_X1  g202(.A(KEYINPUT94), .B1(new_n388), .B2(G107), .ZN(new_n389));
  OAI21_X1  g203(.A(new_n375), .B1(new_n385), .B2(new_n389), .ZN(new_n390));
  INV_X1    g204(.A(KEYINPUT91), .ZN(new_n391));
  AND3_X1   g205(.A1(new_n369), .A2(new_n371), .A3(new_n211), .ZN(new_n392));
  AOI21_X1  g206(.A(new_n211), .B1(new_n369), .B2(new_n371), .ZN(new_n393));
  OAI21_X1  g207(.A(new_n391), .B1(new_n392), .B2(new_n393), .ZN(new_n394));
  OAI21_X1  g208(.A(G107), .B1(new_n383), .B2(new_n378), .ZN(new_n395));
  NAND3_X1  g209(.A1(new_n395), .A2(KEYINPUT91), .A3(new_n372), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n394), .A2(new_n396), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n229), .A2(G143), .ZN(new_n398));
  INV_X1    g212(.A(KEYINPUT13), .ZN(new_n399));
  AOI21_X1  g213(.A(new_n241), .B1(new_n398), .B2(new_n399), .ZN(new_n400));
  XNOR2_X1  g214(.A(new_n373), .B(new_n400), .ZN(new_n401));
  AND3_X1   g215(.A1(new_n397), .A2(new_n401), .A3(KEYINPUT92), .ZN(new_n402));
  AOI21_X1  g216(.A(KEYINPUT92), .B1(new_n397), .B2(new_n401), .ZN(new_n403));
  OAI21_X1  g217(.A(new_n390), .B1(new_n402), .B2(new_n403), .ZN(new_n404));
  INV_X1    g218(.A(G217), .ZN(new_n405));
  NOR3_X1   g219(.A1(new_n187), .A2(new_n405), .A3(G953), .ZN(new_n406));
  INV_X1    g220(.A(new_n406), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n404), .A2(new_n407), .ZN(new_n408));
  INV_X1    g222(.A(KEYINPUT95), .ZN(new_n409));
  OAI211_X1 g223(.A(new_n390), .B(new_n406), .C1(new_n402), .C2(new_n403), .ZN(new_n410));
  NAND3_X1  g224(.A1(new_n408), .A2(new_n409), .A3(new_n410), .ZN(new_n411));
  NAND3_X1  g225(.A1(new_n404), .A2(KEYINPUT95), .A3(new_n407), .ZN(new_n412));
  NAND3_X1  g226(.A1(new_n411), .A2(new_n190), .A3(new_n412), .ZN(new_n413));
  INV_X1    g227(.A(G478), .ZN(new_n414));
  NOR2_X1   g228(.A1(new_n414), .A2(KEYINPUT15), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n413), .A2(new_n415), .ZN(new_n416));
  INV_X1    g230(.A(new_n415), .ZN(new_n417));
  NAND4_X1  g231(.A1(new_n411), .A2(new_n190), .A3(new_n412), .A4(new_n417), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n416), .A2(new_n418), .ZN(new_n419));
  NAND2_X1  g233(.A1(G234), .A2(G237), .ZN(new_n420));
  NAND3_X1  g234(.A1(new_n420), .A2(G952), .A3(new_n192), .ZN(new_n421));
  XNOR2_X1  g235(.A(new_n421), .B(KEYINPUT96), .ZN(new_n422));
  XNOR2_X1  g236(.A(KEYINPUT21), .B(G898), .ZN(new_n423));
  INV_X1    g237(.A(new_n423), .ZN(new_n424));
  NAND3_X1  g238(.A1(new_n420), .A2(G902), .A3(G953), .ZN(new_n425));
  OAI21_X1  g239(.A(new_n422), .B1(new_n424), .B2(new_n425), .ZN(new_n426));
  INV_X1    g240(.A(new_n426), .ZN(new_n427));
  NOR3_X1   g241(.A1(new_n367), .A2(new_n419), .A3(new_n427), .ZN(new_n428));
  AND2_X1   g242(.A1(new_n301), .A2(new_n428), .ZN(new_n429));
  INV_X1    g243(.A(KEYINPUT75), .ZN(new_n430));
  INV_X1    g244(.A(KEYINPUT23), .ZN(new_n431));
  INV_X1    g245(.A(G119), .ZN(new_n432));
  OAI21_X1  g246(.A(new_n431), .B1(new_n432), .B2(G128), .ZN(new_n433));
  NAND3_X1  g247(.A1(new_n229), .A2(KEYINPUT23), .A3(G119), .ZN(new_n434));
  INV_X1    g248(.A(G110), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n432), .A2(G128), .ZN(new_n436));
  NAND4_X1  g250(.A1(new_n433), .A2(new_n434), .A3(new_n435), .A4(new_n436), .ZN(new_n437));
  XOR2_X1   g251(.A(KEYINPUT24), .B(G110), .Z(new_n438));
  XNOR2_X1  g252(.A(G119), .B(G128), .ZN(new_n439));
  OAI22_X1  g253(.A1(new_n437), .A2(KEYINPUT73), .B1(new_n438), .B2(new_n439), .ZN(new_n440));
  AND2_X1   g254(.A1(new_n437), .A2(KEYINPUT73), .ZN(new_n441));
  OAI211_X1 g255(.A(new_n335), .B(new_n308), .C1(new_n440), .C2(new_n441), .ZN(new_n442));
  NAND3_X1  g256(.A1(new_n433), .A2(new_n434), .A3(new_n436), .ZN(new_n443));
  AOI22_X1  g257(.A1(G110), .A2(new_n443), .B1(new_n438), .B2(new_n439), .ZN(new_n444));
  OAI21_X1  g258(.A(new_n444), .B1(new_n342), .B2(new_n343), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n442), .A2(new_n445), .ZN(new_n446));
  NAND3_X1  g260(.A1(new_n192), .A2(G221), .A3(G234), .ZN(new_n447));
  XNOR2_X1  g261(.A(new_n447), .B(KEYINPUT74), .ZN(new_n448));
  XNOR2_X1  g262(.A(KEYINPUT22), .B(G137), .ZN(new_n449));
  XNOR2_X1  g263(.A(new_n448), .B(new_n449), .ZN(new_n450));
  INV_X1    g264(.A(new_n450), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n446), .A2(new_n451), .ZN(new_n452));
  NAND3_X1  g266(.A1(new_n442), .A2(new_n450), .A3(new_n445), .ZN(new_n453));
  NAND3_X1  g267(.A1(new_n452), .A2(new_n190), .A3(new_n453), .ZN(new_n454));
  INV_X1    g268(.A(KEYINPUT25), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  NAND4_X1  g270(.A1(new_n452), .A2(KEYINPUT25), .A3(new_n190), .A4(new_n453), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  AOI21_X1  g272(.A(new_n405), .B1(G234), .B2(new_n190), .ZN(new_n459));
  AOI21_X1  g273(.A(new_n430), .B1(new_n458), .B2(new_n459), .ZN(new_n460));
  INV_X1    g274(.A(new_n459), .ZN(new_n461));
  AOI211_X1 g275(.A(KEYINPUT75), .B(new_n461), .C1(new_n456), .C2(new_n457), .ZN(new_n462));
  NOR2_X1   g276(.A1(new_n460), .A2(new_n462), .ZN(new_n463));
  AND3_X1   g277(.A1(new_n442), .A2(new_n450), .A3(new_n445), .ZN(new_n464));
  AOI21_X1  g278(.A(new_n450), .B1(new_n442), .B2(new_n445), .ZN(new_n465));
  NOR2_X1   g279(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  NOR2_X1   g280(.A1(new_n459), .A2(G902), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n463), .A2(new_n468), .ZN(new_n469));
  XOR2_X1   g283(.A(KEYINPUT64), .B(KEYINPUT30), .Z(new_n470));
  NAND2_X1  g284(.A1(new_n258), .A2(new_n204), .ZN(new_n471));
  INV_X1    g285(.A(KEYINPUT67), .ZN(new_n472));
  XNOR2_X1  g286(.A(G134), .B(G137), .ZN(new_n473));
  OAI21_X1  g287(.A(KEYINPUT66), .B1(new_n473), .B2(new_n254), .ZN(new_n474));
  INV_X1    g288(.A(KEYINPUT66), .ZN(new_n475));
  OAI211_X1 g289(.A(new_n475), .B(G131), .C1(new_n242), .C2(new_n252), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n474), .A2(new_n476), .ZN(new_n477));
  NAND4_X1  g291(.A1(new_n260), .A2(new_n472), .A3(new_n257), .A4(new_n477), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n471), .A2(new_n478), .ZN(new_n479));
  NOR2_X1   g293(.A1(new_n244), .A2(new_n250), .ZN(new_n480));
  AOI22_X1  g294(.A1(new_n480), .A2(new_n254), .B1(new_n476), .B2(new_n474), .ZN(new_n481));
  AOI21_X1  g295(.A(new_n472), .B1(new_n481), .B2(new_n260), .ZN(new_n482));
  OAI21_X1  g296(.A(new_n470), .B1(new_n479), .B2(new_n482), .ZN(new_n483));
  INV_X1    g297(.A(KEYINPUT68), .ZN(new_n484));
  NOR2_X1   g298(.A1(new_n370), .A2(G119), .ZN(new_n485));
  NOR2_X1   g299(.A1(new_n432), .A2(G116), .ZN(new_n486));
  OAI21_X1  g300(.A(new_n484), .B1(new_n485), .B2(new_n486), .ZN(new_n487));
  XNOR2_X1  g301(.A(KEYINPUT2), .B(G113), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n432), .A2(G116), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n370), .A2(G119), .ZN(new_n490));
  NAND3_X1  g304(.A1(new_n489), .A2(new_n490), .A3(KEYINPUT68), .ZN(new_n491));
  NAND3_X1  g305(.A1(new_n487), .A2(new_n488), .A3(new_n491), .ZN(new_n492));
  INV_X1    g306(.A(KEYINPUT69), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n489), .A2(new_n490), .ZN(new_n495));
  INV_X1    g309(.A(new_n495), .ZN(new_n496));
  INV_X1    g310(.A(new_n488), .ZN(new_n497));
  NAND3_X1  g311(.A1(new_n496), .A2(new_n497), .A3(KEYINPUT70), .ZN(new_n498));
  INV_X1    g312(.A(KEYINPUT70), .ZN(new_n499));
  OAI21_X1  g313(.A(new_n499), .B1(new_n495), .B2(new_n488), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n498), .A2(new_n500), .ZN(new_n501));
  NAND4_X1  g315(.A1(new_n487), .A2(KEYINPUT69), .A3(new_n488), .A4(new_n491), .ZN(new_n502));
  NAND3_X1  g316(.A1(new_n494), .A2(new_n501), .A3(new_n502), .ZN(new_n503));
  NAND3_X1  g317(.A1(new_n260), .A2(new_n257), .A3(new_n477), .ZN(new_n504));
  NAND3_X1  g318(.A1(new_n471), .A2(KEYINPUT30), .A3(new_n504), .ZN(new_n505));
  NAND3_X1  g319(.A1(new_n483), .A2(new_n503), .A3(new_n505), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n471), .A2(new_n504), .ZN(new_n507));
  NOR2_X1   g321(.A1(new_n507), .A2(new_n503), .ZN(new_n508));
  XNOR2_X1  g322(.A(KEYINPUT26), .B(G101), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n317), .A2(G210), .ZN(new_n510));
  XNOR2_X1  g324(.A(new_n509), .B(new_n510), .ZN(new_n511));
  XNOR2_X1  g325(.A(KEYINPUT71), .B(KEYINPUT27), .ZN(new_n512));
  XNOR2_X1  g326(.A(new_n511), .B(new_n512), .ZN(new_n513));
  INV_X1    g327(.A(new_n513), .ZN(new_n514));
  NOR2_X1   g328(.A1(new_n508), .A2(new_n514), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n506), .A2(new_n515), .ZN(new_n516));
  INV_X1    g330(.A(KEYINPUT31), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  NAND3_X1  g332(.A1(new_n506), .A2(KEYINPUT31), .A3(new_n515), .ZN(new_n519));
  AND3_X1   g333(.A1(new_n494), .A2(new_n501), .A3(new_n502), .ZN(new_n520));
  NAND3_X1  g334(.A1(new_n520), .A2(new_n471), .A3(new_n504), .ZN(new_n521));
  INV_X1    g335(.A(KEYINPUT28), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n504), .A2(KEYINPUT67), .ZN(new_n524));
  NAND3_X1  g338(.A1(new_n524), .A2(new_n471), .A3(new_n478), .ZN(new_n525));
  AOI21_X1  g339(.A(new_n508), .B1(new_n503), .B2(new_n525), .ZN(new_n526));
  OAI21_X1  g340(.A(new_n523), .B1(new_n526), .B2(new_n522), .ZN(new_n527));
  AOI22_X1  g341(.A1(new_n518), .A2(new_n519), .B1(new_n527), .B2(new_n514), .ZN(new_n528));
  NOR2_X1   g342(.A1(G472), .A2(G902), .ZN(new_n529));
  INV_X1    g343(.A(new_n529), .ZN(new_n530));
  OAI21_X1  g344(.A(KEYINPUT32), .B1(new_n528), .B2(new_n530), .ZN(new_n531));
  OAI21_X1  g345(.A(new_n503), .B1(new_n479), .B2(new_n482), .ZN(new_n532));
  AOI21_X1  g346(.A(new_n522), .B1(new_n532), .B2(new_n521), .ZN(new_n533));
  INV_X1    g347(.A(new_n523), .ZN(new_n534));
  OAI21_X1  g348(.A(new_n514), .B1(new_n533), .B2(new_n534), .ZN(new_n535));
  INV_X1    g349(.A(new_n519), .ZN(new_n536));
  AOI21_X1  g350(.A(KEYINPUT31), .B1(new_n506), .B2(new_n515), .ZN(new_n537));
  OAI21_X1  g351(.A(new_n535), .B1(new_n536), .B2(new_n537), .ZN(new_n538));
  INV_X1    g352(.A(KEYINPUT32), .ZN(new_n539));
  NAND3_X1  g353(.A1(new_n538), .A2(new_n539), .A3(new_n529), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n531), .A2(new_n540), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n506), .A2(new_n521), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n542), .A2(new_n514), .ZN(new_n543));
  INV_X1    g357(.A(KEYINPUT29), .ZN(new_n544));
  AOI21_X1  g358(.A(new_n514), .B1(new_n521), .B2(new_n522), .ZN(new_n545));
  OAI21_X1  g359(.A(new_n545), .B1(new_n526), .B2(new_n522), .ZN(new_n546));
  NAND4_X1  g360(.A1(new_n543), .A2(KEYINPUT72), .A3(new_n544), .A4(new_n546), .ZN(new_n547));
  INV_X1    g361(.A(KEYINPUT72), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n523), .A2(new_n513), .ZN(new_n549));
  OAI21_X1  g363(.A(new_n544), .B1(new_n533), .B2(new_n549), .ZN(new_n550));
  AOI21_X1  g364(.A(new_n513), .B1(new_n506), .B2(new_n521), .ZN(new_n551));
  OAI21_X1  g365(.A(new_n548), .B1(new_n550), .B2(new_n551), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n507), .A2(new_n503), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n553), .A2(new_n521), .ZN(new_n554));
  AOI21_X1  g368(.A(new_n534), .B1(new_n554), .B2(KEYINPUT28), .ZN(new_n555));
  NOR2_X1   g369(.A1(new_n514), .A2(new_n544), .ZN(new_n556));
  AOI21_X1  g370(.A(G902), .B1(new_n555), .B2(new_n556), .ZN(new_n557));
  NAND3_X1  g371(.A1(new_n547), .A2(new_n552), .A3(new_n557), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n558), .A2(G472), .ZN(new_n559));
  AOI21_X1  g373(.A(new_n469), .B1(new_n541), .B2(new_n559), .ZN(new_n560));
  NOR2_X1   g374(.A1(new_n268), .A2(new_n234), .ZN(new_n561));
  INV_X1    g375(.A(KEYINPUT5), .ZN(new_n562));
  NAND3_X1  g376(.A1(new_n562), .A2(new_n432), .A3(G116), .ZN(new_n563));
  OAI21_X1  g377(.A(G113), .B1(new_n563), .B2(KEYINPUT82), .ZN(new_n564));
  AOI21_X1  g378(.A(new_n564), .B1(KEYINPUT82), .B2(new_n563), .ZN(new_n565));
  INV_X1    g379(.A(new_n491), .ZN(new_n566));
  AOI21_X1  g380(.A(KEYINPUT68), .B1(new_n489), .B2(new_n490), .ZN(new_n567));
  OAI21_X1  g381(.A(KEYINPUT5), .B1(new_n566), .B2(new_n567), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n565), .A2(new_n568), .ZN(new_n569));
  NAND3_X1  g383(.A1(new_n561), .A2(new_n569), .A3(new_n501), .ZN(new_n570));
  OAI21_X1  g384(.A(new_n217), .B1(new_n226), .B2(new_n227), .ZN(new_n571));
  OAI21_X1  g385(.A(new_n570), .B1(new_n520), .B2(new_n571), .ZN(new_n572));
  XNOR2_X1  g386(.A(G110), .B(G122), .ZN(new_n573));
  INV_X1    g387(.A(KEYINPUT83), .ZN(new_n574));
  XNOR2_X1  g388(.A(new_n573), .B(new_n574), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n572), .A2(new_n575), .ZN(new_n576));
  XNOR2_X1  g390(.A(new_n573), .B(KEYINPUT83), .ZN(new_n577));
  OAI211_X1 g391(.A(new_n570), .B(new_n577), .C1(new_n520), .C2(new_n571), .ZN(new_n578));
  NAND3_X1  g392(.A1(new_n576), .A2(KEYINPUT6), .A3(new_n578), .ZN(new_n579));
  INV_X1    g393(.A(KEYINPUT6), .ZN(new_n580));
  NAND3_X1  g394(.A1(new_n572), .A2(new_n580), .A3(new_n575), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n203), .A2(G125), .ZN(new_n582));
  INV_X1    g396(.A(new_n582), .ZN(new_n583));
  AOI21_X1  g397(.A(G125), .B1(new_n233), .B2(new_n230), .ZN(new_n584));
  NOR2_X1   g398(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  INV_X1    g399(.A(G224), .ZN(new_n586));
  NOR2_X1   g400(.A1(new_n586), .A2(G953), .ZN(new_n587));
  XOR2_X1   g401(.A(new_n585), .B(new_n587), .Z(new_n588));
  NAND3_X1  g402(.A1(new_n579), .A2(new_n581), .A3(new_n588), .ZN(new_n589));
  INV_X1    g403(.A(KEYINPUT7), .ZN(new_n590));
  OAI22_X1  g404(.A1(new_n583), .A2(new_n584), .B1(new_n590), .B2(new_n587), .ZN(new_n591));
  NOR2_X1   g405(.A1(new_n587), .A2(new_n590), .ZN(new_n592));
  OAI211_X1 g406(.A(new_n582), .B(new_n592), .C1(new_n260), .C2(G125), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n591), .A2(new_n593), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n575), .A2(KEYINPUT8), .ZN(new_n595));
  INV_X1    g409(.A(KEYINPUT8), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n577), .A2(new_n596), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n595), .A2(new_n597), .ZN(new_n598));
  OAI21_X1  g412(.A(new_n565), .B1(new_n562), .B2(new_n495), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n599), .A2(new_n501), .ZN(new_n600));
  AOI21_X1  g414(.A(new_n598), .B1(new_n600), .B2(new_n561), .ZN(new_n601));
  OAI211_X1 g415(.A(new_n569), .B(new_n501), .C1(new_n268), .C2(new_n234), .ZN(new_n602));
  AOI21_X1  g416(.A(new_n594), .B1(new_n601), .B2(new_n602), .ZN(new_n603));
  AOI21_X1  g417(.A(G902), .B1(new_n603), .B2(new_n578), .ZN(new_n604));
  OAI21_X1  g418(.A(G210), .B1(G237), .B2(G902), .ZN(new_n605));
  NAND3_X1  g419(.A1(new_n589), .A2(new_n604), .A3(new_n605), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n589), .A2(new_n604), .ZN(new_n607));
  XOR2_X1   g421(.A(new_n605), .B(KEYINPUT84), .Z(new_n608));
  AOI21_X1  g422(.A(KEYINPUT85), .B1(new_n607), .B2(new_n608), .ZN(new_n609));
  INV_X1    g423(.A(KEYINPUT85), .ZN(new_n610));
  INV_X1    g424(.A(new_n608), .ZN(new_n611));
  AOI211_X1 g425(.A(new_n610), .B(new_n611), .C1(new_n589), .C2(new_n604), .ZN(new_n612));
  OAI21_X1  g426(.A(new_n606), .B1(new_n609), .B2(new_n612), .ZN(new_n613));
  OAI21_X1  g427(.A(G214), .B1(G237), .B2(G902), .ZN(new_n614));
  AND2_X1   g428(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  NAND3_X1  g429(.A1(new_n429), .A2(new_n560), .A3(new_n615), .ZN(new_n616));
  XNOR2_X1  g430(.A(new_n616), .B(G101), .ZN(G3));
  AND3_X1   g431(.A1(new_n589), .A2(new_n604), .A3(new_n605), .ZN(new_n618));
  AOI21_X1  g432(.A(new_n605), .B1(new_n589), .B2(new_n604), .ZN(new_n619));
  OAI211_X1 g433(.A(new_n614), .B(new_n426), .C1(new_n618), .C2(new_n619), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n413), .A2(new_n414), .ZN(new_n621));
  XNOR2_X1  g435(.A(KEYINPUT97), .B(KEYINPUT33), .ZN(new_n622));
  INV_X1    g436(.A(new_n622), .ZN(new_n623));
  NAND3_X1  g437(.A1(new_n411), .A2(new_n412), .A3(new_n623), .ZN(new_n624));
  NAND3_X1  g438(.A1(new_n408), .A2(KEYINPUT33), .A3(new_n410), .ZN(new_n625));
  NAND2_X1  g439(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n190), .A2(G478), .ZN(new_n627));
  OAI21_X1  g441(.A(new_n621), .B1(new_n626), .B2(new_n627), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n628), .A2(new_n367), .ZN(new_n629));
  INV_X1    g443(.A(KEYINPUT98), .ZN(new_n630));
  NAND2_X1  g444(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  NAND3_X1  g445(.A1(new_n628), .A2(KEYINPUT98), .A3(new_n367), .ZN(new_n632));
  AOI21_X1  g446(.A(new_n620), .B1(new_n631), .B2(new_n632), .ZN(new_n633));
  INV_X1    g447(.A(G472), .ZN(new_n634));
  AOI21_X1  g448(.A(new_n634), .B1(new_n538), .B2(new_n190), .ZN(new_n635));
  NOR2_X1   g449(.A1(new_n528), .A2(new_n530), .ZN(new_n636));
  NOR2_X1   g450(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  AOI22_X1  g451(.A1(new_n285), .A2(G469), .B1(new_n294), .B2(new_n299), .ZN(new_n638));
  NOR3_X1   g452(.A1(new_n638), .A2(new_n469), .A3(new_n189), .ZN(new_n639));
  NAND3_X1  g453(.A1(new_n633), .A2(new_n637), .A3(new_n639), .ZN(new_n640));
  XOR2_X1   g454(.A(KEYINPUT34), .B(G104), .Z(new_n641));
  XNOR2_X1  g455(.A(new_n640), .B(new_n641), .ZN(G6));
  INV_X1    g456(.A(KEYINPUT99), .ZN(new_n643));
  AOI21_X1  g457(.A(new_n354), .B1(new_n353), .B2(new_n355), .ZN(new_n644));
  INV_X1    g458(.A(new_n355), .ZN(new_n645));
  AOI211_X1 g459(.A(KEYINPUT20), .B(new_n645), .C1(new_n341), .C2(new_n352), .ZN(new_n646));
  OAI21_X1  g460(.A(new_n366), .B1(new_n644), .B2(new_n646), .ZN(new_n647));
  INV_X1    g461(.A(new_n647), .ZN(new_n648));
  NAND2_X1  g462(.A1(new_n419), .A2(new_n648), .ZN(new_n649));
  OAI21_X1  g463(.A(new_n643), .B1(new_n620), .B2(new_n649), .ZN(new_n650));
  INV_X1    g464(.A(new_n614), .ZN(new_n651));
  INV_X1    g465(.A(new_n605), .ZN(new_n652));
  NAND2_X1  g466(.A1(new_n607), .A2(new_n652), .ZN(new_n653));
  AOI21_X1  g467(.A(new_n651), .B1(new_n653), .B2(new_n606), .ZN(new_n654));
  AOI21_X1  g468(.A(new_n647), .B1(new_n416), .B2(new_n418), .ZN(new_n655));
  NAND4_X1  g469(.A1(new_n654), .A2(KEYINPUT99), .A3(new_n426), .A4(new_n655), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n650), .A2(new_n656), .ZN(new_n657));
  NAND3_X1  g471(.A1(new_n657), .A2(new_n637), .A3(new_n639), .ZN(new_n658));
  XOR2_X1   g472(.A(KEYINPUT35), .B(G107), .Z(new_n659));
  XNOR2_X1  g473(.A(new_n658), .B(new_n659), .ZN(G9));
  NOR2_X1   g474(.A1(new_n451), .A2(KEYINPUT36), .ZN(new_n661));
  XOR2_X1   g475(.A(new_n661), .B(new_n446), .Z(new_n662));
  INV_X1    g476(.A(new_n467), .ZN(new_n663));
  OR2_X1    g477(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  NAND3_X1  g478(.A1(new_n463), .A2(KEYINPUT100), .A3(new_n664), .ZN(new_n665));
  AOI21_X1  g479(.A(KEYINPUT25), .B1(new_n466), .B2(new_n190), .ZN(new_n666));
  INV_X1    g480(.A(new_n457), .ZN(new_n667));
  OAI21_X1  g481(.A(new_n459), .B1(new_n666), .B2(new_n667), .ZN(new_n668));
  NAND2_X1  g482(.A1(new_n668), .A2(KEYINPUT75), .ZN(new_n669));
  NAND3_X1  g483(.A1(new_n458), .A2(new_n430), .A3(new_n459), .ZN(new_n670));
  NAND3_X1  g484(.A1(new_n669), .A2(new_n670), .A3(new_n664), .ZN(new_n671));
  INV_X1    g485(.A(KEYINPUT100), .ZN(new_n672));
  NAND2_X1  g486(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  NAND2_X1  g487(.A1(new_n665), .A2(new_n673), .ZN(new_n674));
  OAI21_X1  g488(.A(G472), .B1(new_n528), .B2(G902), .ZN(new_n675));
  OAI21_X1  g489(.A(new_n675), .B1(new_n530), .B2(new_n528), .ZN(new_n676));
  NOR2_X1   g490(.A1(new_n674), .A2(new_n676), .ZN(new_n677));
  NAND3_X1  g491(.A1(new_n429), .A2(new_n677), .A3(new_n615), .ZN(new_n678));
  XOR2_X1   g492(.A(KEYINPUT37), .B(G110), .Z(new_n679));
  XNOR2_X1  g493(.A(new_n678), .B(new_n679), .ZN(G12));
  AOI22_X1  g494(.A1(new_n531), .A2(new_n540), .B1(new_n558), .B2(G472), .ZN(new_n681));
  NOR2_X1   g495(.A1(new_n681), .A2(new_n674), .ZN(new_n682));
  INV_X1    g496(.A(KEYINPUT103), .ZN(new_n683));
  NOR2_X1   g497(.A1(new_n192), .A2(G900), .ZN(new_n684));
  NAND3_X1  g498(.A1(new_n684), .A2(G902), .A3(new_n420), .ZN(new_n685));
  XOR2_X1   g499(.A(new_n685), .B(KEYINPUT101), .Z(new_n686));
  NAND2_X1  g500(.A1(new_n686), .A2(new_n422), .ZN(new_n687));
  XNOR2_X1  g501(.A(new_n687), .B(KEYINPUT102), .ZN(new_n688));
  INV_X1    g502(.A(new_n688), .ZN(new_n689));
  NAND3_X1  g503(.A1(new_n419), .A2(new_n648), .A3(new_n689), .ZN(new_n690));
  OAI21_X1  g504(.A(new_n614), .B1(new_n618), .B2(new_n619), .ZN(new_n691));
  OAI21_X1  g505(.A(new_n683), .B1(new_n690), .B2(new_n691), .ZN(new_n692));
  NAND4_X1  g506(.A1(new_n654), .A2(KEYINPUT103), .A3(new_n655), .A4(new_n689), .ZN(new_n693));
  NAND2_X1  g507(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  NAND3_X1  g508(.A1(new_n682), .A2(new_n694), .A3(new_n301), .ZN(new_n695));
  XNOR2_X1  g509(.A(new_n695), .B(G128), .ZN(G30));
  INV_X1    g510(.A(new_n542), .ZN(new_n697));
  NOR2_X1   g511(.A1(new_n697), .A2(new_n514), .ZN(new_n698));
  OAI21_X1  g512(.A(new_n190), .B1(new_n554), .B2(new_n513), .ZN(new_n699));
  OAI21_X1  g513(.A(G472), .B1(new_n698), .B2(new_n699), .ZN(new_n700));
  NAND2_X1  g514(.A1(new_n541), .A2(new_n700), .ZN(new_n701));
  INV_X1    g515(.A(KEYINPUT104), .ZN(new_n702));
  XNOR2_X1  g516(.A(new_n701), .B(new_n702), .ZN(new_n703));
  INV_X1    g517(.A(new_n671), .ZN(new_n704));
  AOI21_X1  g518(.A(new_n651), .B1(new_n416), .B2(new_n418), .ZN(new_n705));
  NAND3_X1  g519(.A1(new_n704), .A2(new_n367), .A3(new_n705), .ZN(new_n706));
  XOR2_X1   g520(.A(new_n688), .B(KEYINPUT39), .Z(new_n707));
  NAND2_X1  g521(.A1(new_n301), .A2(new_n707), .ZN(new_n708));
  AOI21_X1  g522(.A(new_n706), .B1(new_n708), .B2(KEYINPUT40), .ZN(new_n709));
  OR2_X1    g523(.A1(new_n708), .A2(KEYINPUT40), .ZN(new_n710));
  OR2_X1    g524(.A1(new_n613), .A2(KEYINPUT38), .ZN(new_n711));
  NAND2_X1  g525(.A1(new_n613), .A2(KEYINPUT38), .ZN(new_n712));
  NAND2_X1  g526(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  NAND4_X1  g527(.A1(new_n703), .A2(new_n709), .A3(new_n710), .A4(new_n713), .ZN(new_n714));
  XNOR2_X1  g528(.A(new_n714), .B(G143), .ZN(G45));
  NAND2_X1  g529(.A1(new_n541), .A2(new_n559), .ZN(new_n716));
  AND2_X1   g530(.A1(new_n665), .A2(new_n673), .ZN(new_n717));
  NAND3_X1  g531(.A1(new_n628), .A2(new_n367), .A3(new_n689), .ZN(new_n718));
  NOR2_X1   g532(.A1(new_n718), .A2(new_n691), .ZN(new_n719));
  NAND4_X1  g533(.A1(new_n716), .A2(new_n717), .A3(new_n719), .A4(new_n301), .ZN(new_n720));
  XNOR2_X1  g534(.A(new_n720), .B(G146), .ZN(G48));
  INV_X1    g535(.A(new_n297), .ZN(new_n722));
  OAI21_X1  g536(.A(G469), .B1(new_n722), .B2(G902), .ZN(new_n723));
  NAND2_X1  g537(.A1(new_n300), .A2(new_n723), .ZN(new_n724));
  NOR2_X1   g538(.A1(new_n724), .A2(new_n189), .ZN(new_n725));
  NAND3_X1  g539(.A1(new_n633), .A2(new_n560), .A3(new_n725), .ZN(new_n726));
  XNOR2_X1  g540(.A(KEYINPUT41), .B(G113), .ZN(new_n727));
  XNOR2_X1  g541(.A(new_n726), .B(new_n727), .ZN(G15));
  NAND3_X1  g542(.A1(new_n657), .A2(new_n560), .A3(new_n725), .ZN(new_n729));
  XNOR2_X1  g543(.A(new_n729), .B(G116), .ZN(G18));
  NOR3_X1   g544(.A1(new_n724), .A2(new_n189), .A3(new_n691), .ZN(new_n731));
  NAND4_X1  g545(.A1(new_n731), .A2(new_n716), .A3(new_n717), .A4(new_n428), .ZN(new_n732));
  XNOR2_X1  g546(.A(new_n732), .B(G119), .ZN(G21));
  OR2_X1    g547(.A1(new_n555), .A2(new_n513), .ZN(new_n734));
  NAND2_X1  g548(.A1(new_n518), .A2(new_n519), .ZN(new_n735));
  AOI21_X1  g549(.A(new_n530), .B1(new_n734), .B2(new_n735), .ZN(new_n736));
  NOR3_X1   g550(.A1(new_n469), .A2(new_n635), .A3(new_n736), .ZN(new_n737));
  NAND2_X1  g551(.A1(new_n653), .A2(new_n606), .ZN(new_n738));
  AND3_X1   g552(.A1(new_n738), .A2(new_n367), .A3(new_n705), .ZN(new_n739));
  NAND4_X1  g553(.A1(new_n737), .A2(new_n725), .A3(new_n426), .A4(new_n739), .ZN(new_n740));
  XNOR2_X1  g554(.A(new_n740), .B(G122), .ZN(G24));
  NOR3_X1   g555(.A1(new_n704), .A2(new_n635), .A3(new_n736), .ZN(new_n742));
  INV_X1    g556(.A(new_n718), .ZN(new_n743));
  NAND3_X1  g557(.A1(new_n731), .A2(new_n742), .A3(new_n743), .ZN(new_n744));
  XNOR2_X1  g558(.A(new_n744), .B(G125), .ZN(G27));
  AND2_X1   g559(.A1(new_n606), .A2(new_n614), .ZN(new_n746));
  OAI21_X1  g560(.A(new_n746), .B1(new_n609), .B2(new_n612), .ZN(new_n747));
  NOR3_X1   g561(.A1(new_n747), .A2(new_n638), .A3(new_n189), .ZN(new_n748));
  NAND3_X1  g562(.A1(new_n748), .A2(new_n560), .A3(new_n743), .ZN(new_n749));
  INV_X1    g563(.A(KEYINPUT42), .ZN(new_n750));
  NAND2_X1  g564(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  NAND4_X1  g565(.A1(new_n748), .A2(new_n560), .A3(KEYINPUT42), .A4(new_n743), .ZN(new_n752));
  NAND2_X1  g566(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  XNOR2_X1  g567(.A(new_n753), .B(G131), .ZN(G33));
  AND4_X1   g568(.A1(KEYINPUT105), .A2(new_n419), .A3(new_n648), .A4(new_n689), .ZN(new_n755));
  AOI21_X1  g569(.A(KEYINPUT105), .B1(new_n655), .B2(new_n689), .ZN(new_n756));
  NOR2_X1   g570(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  NAND3_X1  g571(.A1(new_n748), .A2(new_n560), .A3(new_n757), .ZN(new_n758));
  XNOR2_X1  g572(.A(new_n758), .B(G134), .ZN(G36));
  INV_X1    g573(.A(new_n707), .ZN(new_n760));
  NAND2_X1  g574(.A1(new_n278), .A2(new_n280), .ZN(new_n761));
  AOI21_X1  g575(.A(new_n284), .B1(new_n761), .B2(new_n194), .ZN(new_n762));
  NAND2_X1  g576(.A1(new_n762), .A2(KEYINPUT45), .ZN(new_n763));
  INV_X1    g577(.A(KEYINPUT45), .ZN(new_n764));
  OAI21_X1  g578(.A(new_n764), .B1(new_n281), .B2(new_n284), .ZN(new_n765));
  NAND3_X1  g579(.A1(new_n763), .A2(G469), .A3(new_n765), .ZN(new_n766));
  NAND2_X1  g580(.A1(G469), .A2(G902), .ZN(new_n767));
  NAND2_X1  g581(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  INV_X1    g582(.A(KEYINPUT46), .ZN(new_n769));
  AOI22_X1  g583(.A1(new_n768), .A2(new_n769), .B1(new_n294), .B2(new_n299), .ZN(new_n770));
  NAND3_X1  g584(.A1(new_n766), .A2(KEYINPUT46), .A3(new_n767), .ZN(new_n771));
  AOI211_X1 g585(.A(new_n189), .B(new_n760), .C1(new_n770), .C2(new_n771), .ZN(new_n772));
  INV_X1    g586(.A(KEYINPUT44), .ZN(new_n773));
  AND2_X1   g587(.A1(new_n362), .A2(new_n366), .ZN(new_n774));
  NAND2_X1  g588(.A1(new_n774), .A2(new_n628), .ZN(new_n775));
  XNOR2_X1  g589(.A(KEYINPUT106), .B(KEYINPUT43), .ZN(new_n776));
  NOR2_X1   g590(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  INV_X1    g591(.A(KEYINPUT106), .ZN(new_n778));
  AOI22_X1  g592(.A1(new_n774), .A2(new_n628), .B1(new_n778), .B2(KEYINPUT43), .ZN(new_n779));
  NOR2_X1   g593(.A1(new_n777), .A2(new_n779), .ZN(new_n780));
  NAND2_X1  g594(.A1(new_n676), .A2(new_n671), .ZN(new_n781));
  OAI21_X1  g595(.A(new_n773), .B1(new_n780), .B2(new_n781), .ZN(new_n782));
  NOR2_X1   g596(.A1(new_n637), .A2(new_n704), .ZN(new_n783));
  OAI211_X1 g597(.A(new_n783), .B(KEYINPUT44), .C1(new_n777), .C2(new_n779), .ZN(new_n784));
  INV_X1    g598(.A(new_n747), .ZN(new_n785));
  AND3_X1   g599(.A1(new_n784), .A2(KEYINPUT107), .A3(new_n785), .ZN(new_n786));
  AOI21_X1  g600(.A(KEYINPUT107), .B1(new_n784), .B2(new_n785), .ZN(new_n787));
  OAI211_X1 g601(.A(new_n772), .B(new_n782), .C1(new_n786), .C2(new_n787), .ZN(new_n788));
  XNOR2_X1  g602(.A(new_n788), .B(G137), .ZN(G39));
  NAND3_X1  g603(.A1(new_n785), .A2(new_n743), .A3(new_n469), .ZN(new_n790));
  NOR2_X1   g604(.A1(new_n790), .A2(new_n716), .ZN(new_n791));
  NAND2_X1  g605(.A1(new_n770), .A2(new_n771), .ZN(new_n792));
  INV_X1    g606(.A(new_n189), .ZN(new_n793));
  AOI21_X1  g607(.A(KEYINPUT47), .B1(new_n792), .B2(new_n793), .ZN(new_n794));
  INV_X1    g608(.A(KEYINPUT47), .ZN(new_n795));
  AOI211_X1 g609(.A(new_n795), .B(new_n189), .C1(new_n770), .C2(new_n771), .ZN(new_n796));
  OAI21_X1  g610(.A(new_n791), .B1(new_n794), .B2(new_n796), .ZN(new_n797));
  XNOR2_X1  g611(.A(new_n797), .B(G140), .ZN(G42));
  NOR4_X1   g612(.A1(new_n775), .A2(new_n469), .A3(new_n651), .A4(new_n189), .ZN(new_n799));
  XOR2_X1   g613(.A(new_n799), .B(KEYINPUT108), .Z(new_n800));
  XNOR2_X1  g614(.A(new_n724), .B(KEYINPUT49), .ZN(new_n801));
  OR4_X1    g615(.A1(new_n703), .A2(new_n800), .A3(new_n713), .A4(new_n801), .ZN(new_n802));
  INV_X1    g616(.A(KEYINPUT53), .ZN(new_n803));
  INV_X1    g617(.A(KEYINPUT109), .ZN(new_n804));
  NAND4_X1  g618(.A1(new_n301), .A2(new_n614), .A3(new_n613), .A4(new_n428), .ZN(new_n805));
  INV_X1    g619(.A(new_n469), .ZN(new_n806));
  NAND2_X1  g620(.A1(new_n716), .A2(new_n806), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n717), .A2(new_n637), .ZN(new_n808));
  AOI21_X1  g622(.A(new_n805), .B1(new_n807), .B2(new_n808), .ZN(new_n809));
  NAND3_X1  g623(.A1(new_n419), .A2(new_n366), .A3(new_n362), .ZN(new_n810));
  AOI21_X1  g624(.A(new_n427), .B1(new_n629), .B2(new_n810), .ZN(new_n811));
  NAND3_X1  g625(.A1(new_n811), .A2(new_n614), .A3(new_n613), .ZN(new_n812));
  NAND3_X1  g626(.A1(new_n301), .A2(new_n637), .A3(new_n806), .ZN(new_n813));
  NOR2_X1   g627(.A1(new_n812), .A2(new_n813), .ZN(new_n814));
  OAI21_X1  g628(.A(new_n804), .B1(new_n809), .B2(new_n814), .ZN(new_n815));
  NAND4_X1  g629(.A1(new_n639), .A2(new_n615), .A3(new_n637), .A4(new_n811), .ZN(new_n816));
  NAND4_X1  g630(.A1(new_n616), .A2(new_n678), .A3(new_n816), .A4(KEYINPUT109), .ZN(new_n817));
  NAND2_X1  g631(.A1(new_n815), .A2(new_n817), .ZN(new_n818));
  AND4_X1   g632(.A1(new_n726), .A2(new_n729), .A3(new_n732), .A4(new_n740), .ZN(new_n819));
  NAND4_X1  g633(.A1(new_n648), .A2(new_n416), .A3(new_n418), .A4(new_n689), .ZN(new_n820));
  NOR2_X1   g634(.A1(new_n747), .A2(new_n820), .ZN(new_n821));
  NAND4_X1  g635(.A1(new_n716), .A2(new_n821), .A3(new_n717), .A4(new_n301), .ZN(new_n822));
  NAND4_X1  g636(.A1(new_n742), .A2(new_n785), .A3(new_n301), .A4(new_n743), .ZN(new_n823));
  NAND3_X1  g637(.A1(new_n758), .A2(new_n822), .A3(new_n823), .ZN(new_n824));
  AOI21_X1  g638(.A(new_n824), .B1(new_n751), .B2(new_n752), .ZN(new_n825));
  NAND3_X1  g639(.A1(new_n818), .A2(new_n819), .A3(new_n825), .ZN(new_n826));
  NOR2_X1   g640(.A1(new_n671), .A2(new_n688), .ZN(new_n827));
  NAND4_X1  g641(.A1(new_n701), .A2(new_n301), .A3(new_n739), .A4(new_n827), .ZN(new_n828));
  NAND4_X1  g642(.A1(new_n695), .A2(new_n720), .A3(new_n744), .A4(new_n828), .ZN(new_n829));
  XNOR2_X1  g643(.A(new_n829), .B(KEYINPUT52), .ZN(new_n830));
  OAI21_X1  g644(.A(new_n803), .B1(new_n826), .B2(new_n830), .ZN(new_n831));
  INV_X1    g645(.A(KEYINPUT110), .ZN(new_n832));
  INV_X1    g646(.A(KEYINPUT52), .ZN(new_n833));
  XNOR2_X1  g647(.A(new_n829), .B(new_n833), .ZN(new_n834));
  INV_X1    g648(.A(new_n824), .ZN(new_n835));
  AND3_X1   g649(.A1(new_n819), .A2(new_n753), .A3(new_n835), .ZN(new_n836));
  NAND4_X1  g650(.A1(new_n834), .A2(new_n836), .A3(KEYINPUT53), .A4(new_n818), .ZN(new_n837));
  NAND3_X1  g651(.A1(new_n831), .A2(new_n832), .A3(new_n837), .ZN(new_n838));
  OAI211_X1 g652(.A(KEYINPUT110), .B(new_n803), .C1(new_n826), .C2(new_n830), .ZN(new_n839));
  NAND3_X1  g653(.A1(new_n838), .A2(KEYINPUT54), .A3(new_n839), .ZN(new_n840));
  INV_X1    g654(.A(KEYINPUT54), .ZN(new_n841));
  NAND3_X1  g655(.A1(new_n831), .A2(new_n841), .A3(new_n837), .ZN(new_n842));
  AND3_X1   g656(.A1(new_n840), .A2(KEYINPUT111), .A3(new_n842), .ZN(new_n843));
  AOI21_X1  g657(.A(KEYINPUT111), .B1(new_n840), .B2(new_n842), .ZN(new_n844));
  NAND4_X1  g658(.A1(new_n711), .A2(new_n651), .A3(new_n712), .A4(new_n725), .ZN(new_n845));
  INV_X1    g659(.A(new_n422), .ZN(new_n846));
  OAI211_X1 g660(.A(new_n737), .B(new_n846), .C1(new_n777), .C2(new_n779), .ZN(new_n847));
  INV_X1    g661(.A(KEYINPUT50), .ZN(new_n848));
  OR3_X1    g662(.A1(new_n845), .A2(new_n847), .A3(new_n848), .ZN(new_n849));
  OAI21_X1  g663(.A(new_n848), .B1(new_n845), .B2(new_n847), .ZN(new_n850));
  NAND2_X1  g664(.A1(new_n849), .A2(new_n850), .ZN(new_n851));
  NOR2_X1   g665(.A1(new_n703), .A2(new_n469), .ZN(new_n852));
  NAND2_X1  g666(.A1(new_n725), .A2(new_n785), .ZN(new_n853));
  NAND2_X1  g667(.A1(new_n853), .A2(KEYINPUT113), .ZN(new_n854));
  INV_X1    g668(.A(KEYINPUT113), .ZN(new_n855));
  NAND3_X1  g669(.A1(new_n725), .A2(new_n785), .A3(new_n855), .ZN(new_n856));
  AND3_X1   g670(.A1(new_n854), .A2(new_n846), .A3(new_n856), .ZN(new_n857));
  NOR2_X1   g671(.A1(new_n628), .A2(new_n367), .ZN(new_n858));
  NAND3_X1  g672(.A1(new_n852), .A2(new_n857), .A3(new_n858), .ZN(new_n859));
  INV_X1    g673(.A(new_n780), .ZN(new_n860));
  NAND3_X1  g674(.A1(new_n857), .A2(new_n742), .A3(new_n860), .ZN(new_n861));
  NAND3_X1  g675(.A1(new_n851), .A2(new_n859), .A3(new_n861), .ZN(new_n862));
  INV_X1    g676(.A(new_n862), .ZN(new_n863));
  INV_X1    g677(.A(new_n847), .ZN(new_n864));
  NAND2_X1  g678(.A1(new_n792), .A2(new_n793), .ZN(new_n865));
  NAND2_X1  g679(.A1(new_n865), .A2(new_n795), .ZN(new_n866));
  NAND3_X1  g680(.A1(new_n792), .A2(KEYINPUT47), .A3(new_n793), .ZN(new_n867));
  NAND2_X1  g681(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  OR2_X1    g682(.A1(new_n724), .A2(KEYINPUT112), .ZN(new_n869));
  NAND2_X1  g683(.A1(new_n724), .A2(KEYINPUT112), .ZN(new_n870));
  AND3_X1   g684(.A1(new_n869), .A2(new_n189), .A3(new_n870), .ZN(new_n871));
  OAI211_X1 g685(.A(new_n785), .B(new_n864), .C1(new_n868), .C2(new_n871), .ZN(new_n872));
  NAND3_X1  g686(.A1(new_n863), .A2(new_n872), .A3(KEYINPUT51), .ZN(new_n873));
  INV_X1    g687(.A(KEYINPUT51), .ZN(new_n874));
  NAND2_X1  g688(.A1(new_n864), .A2(new_n785), .ZN(new_n875));
  NOR2_X1   g689(.A1(new_n794), .A2(new_n796), .ZN(new_n876));
  INV_X1    g690(.A(new_n871), .ZN(new_n877));
  AOI21_X1  g691(.A(new_n875), .B1(new_n876), .B2(new_n877), .ZN(new_n878));
  OAI21_X1  g692(.A(new_n874), .B1(new_n878), .B2(new_n862), .ZN(new_n879));
  NAND4_X1  g693(.A1(new_n860), .A2(new_n854), .A3(new_n846), .A4(new_n856), .ZN(new_n880));
  NOR2_X1   g694(.A1(new_n880), .A2(new_n807), .ZN(new_n881));
  NAND3_X1  g695(.A1(new_n881), .A2(KEYINPUT114), .A3(KEYINPUT48), .ZN(new_n882));
  XOR2_X1   g696(.A(KEYINPUT114), .B(KEYINPUT48), .Z(new_n883));
  OAI21_X1  g697(.A(new_n883), .B1(new_n880), .B2(new_n807), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n631), .A2(new_n632), .ZN(new_n885));
  NAND3_X1  g699(.A1(new_n852), .A2(new_n857), .A3(new_n885), .ZN(new_n886));
  NAND2_X1  g700(.A1(new_n192), .A2(G952), .ZN(new_n887));
  AOI21_X1  g701(.A(new_n887), .B1(new_n864), .B2(new_n731), .ZN(new_n888));
  AND4_X1   g702(.A1(new_n882), .A2(new_n884), .A3(new_n886), .A4(new_n888), .ZN(new_n889));
  NAND3_X1  g703(.A1(new_n873), .A2(new_n879), .A3(new_n889), .ZN(new_n890));
  NAND2_X1  g704(.A1(new_n890), .A2(KEYINPUT115), .ZN(new_n891));
  INV_X1    g705(.A(KEYINPUT115), .ZN(new_n892));
  NAND4_X1  g706(.A1(new_n873), .A2(new_n879), .A3(new_n892), .A4(new_n889), .ZN(new_n893));
  NAND2_X1  g707(.A1(new_n891), .A2(new_n893), .ZN(new_n894));
  NOR3_X1   g708(.A1(new_n843), .A2(new_n844), .A3(new_n894), .ZN(new_n895));
  NOR2_X1   g709(.A1(G952), .A2(G953), .ZN(new_n896));
  OAI21_X1  g710(.A(new_n802), .B1(new_n895), .B2(new_n896), .ZN(G75));
  NOR2_X1   g711(.A1(new_n192), .A2(G952), .ZN(new_n898));
  INV_X1    g712(.A(new_n898), .ZN(new_n899));
  NAND2_X1  g713(.A1(new_n831), .A2(new_n837), .ZN(new_n900));
  NAND2_X1  g714(.A1(new_n900), .A2(G902), .ZN(new_n901));
  NOR2_X1   g715(.A1(new_n901), .A2(new_n611), .ZN(new_n902));
  NAND2_X1  g716(.A1(new_n579), .A2(new_n581), .ZN(new_n903));
  XNOR2_X1  g717(.A(new_n903), .B(new_n588), .ZN(new_n904));
  XOR2_X1   g718(.A(new_n904), .B(KEYINPUT55), .Z(new_n905));
  XOR2_X1   g719(.A(KEYINPUT117), .B(KEYINPUT56), .Z(new_n906));
  OR2_X1    g720(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  OAI21_X1  g721(.A(new_n899), .B1(new_n902), .B2(new_n907), .ZN(new_n908));
  INV_X1    g722(.A(G210), .ZN(new_n909));
  OR3_X1    g723(.A1(new_n901), .A2(KEYINPUT116), .A3(new_n909), .ZN(new_n910));
  INV_X1    g724(.A(KEYINPUT56), .ZN(new_n911));
  OAI21_X1  g725(.A(KEYINPUT116), .B1(new_n901), .B2(new_n909), .ZN(new_n912));
  NAND3_X1  g726(.A1(new_n910), .A2(new_n911), .A3(new_n912), .ZN(new_n913));
  AOI21_X1  g727(.A(new_n908), .B1(new_n913), .B2(new_n905), .ZN(G51));
  INV_X1    g728(.A(KEYINPUT118), .ZN(new_n915));
  NOR2_X1   g729(.A1(new_n901), .A2(new_n766), .ZN(new_n916));
  XOR2_X1   g730(.A(new_n767), .B(KEYINPUT57), .Z(new_n917));
  AND3_X1   g731(.A1(new_n831), .A2(new_n841), .A3(new_n837), .ZN(new_n918));
  AOI21_X1  g732(.A(new_n841), .B1(new_n831), .B2(new_n837), .ZN(new_n919));
  OAI21_X1  g733(.A(new_n917), .B1(new_n918), .B2(new_n919), .ZN(new_n920));
  AOI21_X1  g734(.A(new_n916), .B1(new_n297), .B2(new_n920), .ZN(new_n921));
  OAI21_X1  g735(.A(new_n915), .B1(new_n921), .B2(new_n898), .ZN(new_n922));
  NAND2_X1  g736(.A1(new_n900), .A2(KEYINPUT54), .ZN(new_n923));
  NAND2_X1  g737(.A1(new_n923), .A2(new_n842), .ZN(new_n924));
  AOI21_X1  g738(.A(new_n722), .B1(new_n924), .B2(new_n917), .ZN(new_n925));
  OAI211_X1 g739(.A(KEYINPUT118), .B(new_n899), .C1(new_n925), .C2(new_n916), .ZN(new_n926));
  NAND2_X1  g740(.A1(new_n922), .A2(new_n926), .ZN(G54));
  INV_X1    g741(.A(KEYINPUT119), .ZN(new_n928));
  INV_X1    g742(.A(new_n901), .ZN(new_n929));
  AND2_X1   g743(.A1(KEYINPUT58), .A2(G475), .ZN(new_n930));
  NAND2_X1  g744(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  INV_X1    g745(.A(new_n353), .ZN(new_n932));
  OAI21_X1  g746(.A(new_n928), .B1(new_n931), .B2(new_n932), .ZN(new_n933));
  AOI21_X1  g747(.A(new_n898), .B1(new_n931), .B2(new_n932), .ZN(new_n934));
  NAND4_X1  g748(.A1(new_n929), .A2(KEYINPUT119), .A3(new_n353), .A4(new_n930), .ZN(new_n935));
  AND3_X1   g749(.A1(new_n933), .A2(new_n934), .A3(new_n935), .ZN(G60));
  INV_X1    g750(.A(new_n924), .ZN(new_n937));
  NAND2_X1  g751(.A1(G478), .A2(G902), .ZN(new_n938));
  XOR2_X1   g752(.A(new_n938), .B(KEYINPUT59), .Z(new_n939));
  INV_X1    g753(.A(new_n939), .ZN(new_n940));
  NAND3_X1  g754(.A1(new_n624), .A2(new_n625), .A3(new_n940), .ZN(new_n941));
  OAI21_X1  g755(.A(new_n899), .B1(new_n937), .B2(new_n941), .ZN(new_n942));
  OAI21_X1  g756(.A(new_n940), .B1(new_n843), .B2(new_n844), .ZN(new_n943));
  AOI21_X1  g757(.A(new_n942), .B1(new_n943), .B2(new_n626), .ZN(G63));
  XNOR2_X1  g758(.A(KEYINPUT120), .B(KEYINPUT60), .ZN(new_n945));
  NOR2_X1   g759(.A1(new_n405), .A2(new_n190), .ZN(new_n946));
  XNOR2_X1  g760(.A(new_n945), .B(new_n946), .ZN(new_n947));
  NAND2_X1  g761(.A1(new_n900), .A2(new_n947), .ZN(new_n948));
  INV_X1    g762(.A(new_n466), .ZN(new_n949));
  AOI21_X1  g763(.A(new_n898), .B1(new_n948), .B2(new_n949), .ZN(new_n950));
  OAI21_X1  g764(.A(new_n950), .B1(new_n662), .B2(new_n948), .ZN(new_n951));
  XNOR2_X1  g765(.A(KEYINPUT121), .B(KEYINPUT61), .ZN(new_n952));
  XNOR2_X1  g766(.A(new_n951), .B(new_n952), .ZN(G66));
  OAI21_X1  g767(.A(G953), .B1(new_n423), .B2(new_n586), .ZN(new_n954));
  AND2_X1   g768(.A1(new_n818), .A2(new_n819), .ZN(new_n955));
  OAI21_X1  g769(.A(new_n954), .B1(new_n955), .B2(G953), .ZN(new_n956));
  OAI21_X1  g770(.A(new_n903), .B1(G898), .B2(new_n192), .ZN(new_n957));
  XOR2_X1   g771(.A(new_n957), .B(KEYINPUT122), .Z(new_n958));
  XNOR2_X1  g772(.A(new_n956), .B(new_n958), .ZN(G69));
  AOI21_X1  g773(.A(new_n192), .B1(G227), .B2(G900), .ZN(new_n960));
  INV_X1    g774(.A(new_n791), .ZN(new_n961));
  AOI21_X1  g775(.A(new_n961), .B1(new_n866), .B2(new_n867), .ZN(new_n962));
  NAND3_X1  g776(.A1(new_n695), .A2(new_n720), .A3(new_n744), .ZN(new_n963));
  INV_X1    g777(.A(new_n963), .ZN(new_n964));
  NAND2_X1  g778(.A1(new_n964), .A2(new_n714), .ZN(new_n965));
  INV_X1    g779(.A(KEYINPUT62), .ZN(new_n966));
  NAND2_X1  g780(.A1(new_n965), .A2(new_n966), .ZN(new_n967));
  NAND3_X1  g781(.A1(new_n964), .A2(new_n714), .A3(KEYINPUT62), .ZN(new_n968));
  AOI21_X1  g782(.A(new_n962), .B1(new_n967), .B2(new_n968), .ZN(new_n969));
  INV_X1    g783(.A(KEYINPUT124), .ZN(new_n970));
  AOI21_X1  g784(.A(new_n747), .B1(new_n629), .B2(new_n810), .ZN(new_n971));
  NAND3_X1  g785(.A1(new_n971), .A2(new_n301), .A3(new_n707), .ZN(new_n972));
  NOR2_X1   g786(.A1(new_n972), .A2(new_n807), .ZN(new_n973));
  INV_X1    g787(.A(new_n973), .ZN(new_n974));
  AND3_X1   g788(.A1(new_n788), .A2(new_n970), .A3(new_n974), .ZN(new_n975));
  AOI21_X1  g789(.A(new_n970), .B1(new_n788), .B2(new_n974), .ZN(new_n976));
  OAI211_X1 g790(.A(new_n969), .B(KEYINPUT125), .C1(new_n975), .C2(new_n976), .ZN(new_n977));
  INV_X1    g791(.A(new_n977), .ZN(new_n978));
  NAND4_X1  g792(.A1(new_n782), .A2(new_n792), .A3(new_n793), .A4(new_n707), .ZN(new_n979));
  INV_X1    g793(.A(new_n787), .ZN(new_n980));
  NAND3_X1  g794(.A1(new_n784), .A2(KEYINPUT107), .A3(new_n785), .ZN(new_n981));
  AOI21_X1  g795(.A(new_n979), .B1(new_n980), .B2(new_n981), .ZN(new_n982));
  OAI21_X1  g796(.A(KEYINPUT124), .B1(new_n982), .B2(new_n973), .ZN(new_n983));
  NAND3_X1  g797(.A1(new_n788), .A2(new_n970), .A3(new_n974), .ZN(new_n984));
  NAND2_X1  g798(.A1(new_n983), .A2(new_n984), .ZN(new_n985));
  AOI21_X1  g799(.A(KEYINPUT125), .B1(new_n985), .B2(new_n969), .ZN(new_n986));
  OAI21_X1  g800(.A(new_n192), .B1(new_n978), .B2(new_n986), .ZN(new_n987));
  NAND2_X1  g801(.A1(new_n483), .A2(new_n505), .ZN(new_n988));
  XNOR2_X1  g802(.A(new_n988), .B(new_n324), .ZN(new_n989));
  XOR2_X1   g803(.A(new_n989), .B(KEYINPUT123), .Z(new_n990));
  NAND2_X1  g804(.A1(new_n987), .A2(new_n990), .ZN(new_n991));
  AND2_X1   g805(.A1(new_n560), .A2(new_n739), .ZN(new_n992));
  NAND2_X1  g806(.A1(new_n772), .A2(new_n992), .ZN(new_n993));
  NAND4_X1  g807(.A1(new_n993), .A2(new_n753), .A3(new_n758), .A4(new_n964), .ZN(new_n994));
  INV_X1    g808(.A(new_n994), .ZN(new_n995));
  NAND4_X1  g809(.A1(new_n995), .A2(KEYINPUT126), .A3(new_n788), .A4(new_n797), .ZN(new_n996));
  INV_X1    g810(.A(KEYINPUT126), .ZN(new_n997));
  NAND2_X1  g811(.A1(new_n788), .A2(new_n797), .ZN(new_n998));
  OAI21_X1  g812(.A(new_n997), .B1(new_n998), .B2(new_n994), .ZN(new_n999));
  AOI21_X1  g813(.A(G953), .B1(new_n996), .B2(new_n999), .ZN(new_n1000));
  OAI21_X1  g814(.A(new_n989), .B1(new_n1000), .B2(new_n684), .ZN(new_n1001));
  AOI21_X1  g815(.A(new_n960), .B1(new_n991), .B2(new_n1001), .ZN(new_n1002));
  OAI21_X1  g816(.A(new_n969), .B1(new_n975), .B2(new_n976), .ZN(new_n1003));
  INV_X1    g817(.A(KEYINPUT125), .ZN(new_n1004));
  NAND2_X1  g818(.A1(new_n1003), .A2(new_n1004), .ZN(new_n1005));
  AOI21_X1  g819(.A(G953), .B1(new_n1005), .B2(new_n977), .ZN(new_n1006));
  INV_X1    g820(.A(new_n990), .ZN(new_n1007));
  OAI211_X1 g821(.A(new_n1001), .B(new_n960), .C1(new_n1006), .C2(new_n1007), .ZN(new_n1008));
  INV_X1    g822(.A(new_n1008), .ZN(new_n1009));
  NOR2_X1   g823(.A1(new_n1002), .A2(new_n1009), .ZN(G72));
  AND3_X1   g824(.A1(new_n996), .A2(new_n999), .A3(new_n955), .ZN(new_n1011));
  NAND2_X1  g825(.A1(G472), .A2(G902), .ZN(new_n1012));
  XOR2_X1   g826(.A(new_n1012), .B(KEYINPUT63), .Z(new_n1013));
  INV_X1    g827(.A(new_n1013), .ZN(new_n1014));
  OAI211_X1 g828(.A(new_n514), .B(new_n697), .C1(new_n1011), .C2(new_n1014), .ZN(new_n1015));
  AOI21_X1  g829(.A(new_n1014), .B1(new_n543), .B2(new_n516), .ZN(new_n1016));
  XNOR2_X1  g830(.A(new_n1016), .B(KEYINPUT127), .ZN(new_n1017));
  NAND3_X1  g831(.A1(new_n838), .A2(new_n839), .A3(new_n1017), .ZN(new_n1018));
  NAND3_X1  g832(.A1(new_n1015), .A2(new_n899), .A3(new_n1018), .ZN(new_n1019));
  NAND3_X1  g833(.A1(new_n1005), .A2(new_n955), .A3(new_n977), .ZN(new_n1020));
  NAND2_X1  g834(.A1(new_n1020), .A2(new_n1013), .ZN(new_n1021));
  AOI21_X1  g835(.A(new_n1019), .B1(new_n698), .B2(new_n1021), .ZN(G57));
endmodule


