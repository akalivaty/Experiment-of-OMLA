//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 0 0 0 1 1 1 0 0 0 1 1 1 0 0 1 0 0 0 0 0 0 1 0 1 1 1 0 1 1 0 0 0 1 1 0 1 1 1 0 0 1 1 1 0 1 0 0 0 1 1 1 0 0 0 1 1 0 0 1 1 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:33:09 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n447, new_n448, new_n450, new_n453, new_n454, new_n455,
    new_n456, new_n457, new_n458, new_n459, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n484, new_n485, new_n486,
    new_n487, new_n488, new_n489, new_n490, new_n491, new_n492, new_n493,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n533, new_n534, new_n535, new_n536, new_n537, new_n538,
    new_n541, new_n542, new_n543, new_n544, new_n545, new_n546, new_n547,
    new_n548, new_n549, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n557, new_n558, new_n559, new_n560, new_n561, new_n562, new_n563,
    new_n564, new_n565, new_n567, new_n568, new_n570, new_n571, new_n573,
    new_n574, new_n575, new_n576, new_n577, new_n578, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n589, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n619, new_n622, new_n623, new_n624, new_n626,
    new_n627, new_n628, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1197, new_n1198;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  XOR2_X1   g012(.A(KEYINPUT64), .B(G96), .Z(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  XNOR2_X1  g021(.A(KEYINPUT65), .B(KEYINPUT1), .ZN(new_n447));
  NAND2_X1  g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XNOR2_X1  g023(.A(new_n447), .B(new_n448), .ZN(G223));
  INV_X1    g024(.A(new_n448), .ZN(new_n450));
  NAND2_X1  g025(.A1(new_n450), .A2(G567), .ZN(G234));
  NAND2_X1  g026(.A1(new_n450), .A2(G2106), .ZN(G217));
  NOR4_X1   g027(.A1(G220), .A2(G221), .A3(G218), .A4(G219), .ZN(new_n453));
  XNOR2_X1  g028(.A(KEYINPUT66), .B(KEYINPUT2), .ZN(new_n454));
  XOR2_X1   g029(.A(new_n453), .B(new_n454), .Z(new_n455));
  INV_X1    g030(.A(new_n455), .ZN(new_n456));
  NAND4_X1  g031(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n457));
  XNOR2_X1  g032(.A(new_n457), .B(KEYINPUT67), .ZN(new_n458));
  INV_X1    g033(.A(new_n458), .ZN(new_n459));
  NOR2_X1   g034(.A1(new_n456), .A2(new_n459), .ZN(G325));
  INV_X1    g035(.A(G325), .ZN(G261));
  AOI22_X1  g036(.A1(new_n456), .A2(G2106), .B1(G567), .B2(new_n459), .ZN(G319));
  INV_X1    g037(.A(G2104), .ZN(new_n463));
  NAND3_X1  g038(.A1(new_n463), .A2(KEYINPUT70), .A3(KEYINPUT3), .ZN(new_n464));
  INV_X1    g039(.A(new_n464), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n463), .A2(KEYINPUT3), .ZN(new_n466));
  INV_X1    g041(.A(KEYINPUT3), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n467), .A2(G2104), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n468), .A2(KEYINPUT70), .ZN(new_n469));
  AOI21_X1  g044(.A(new_n465), .B1(new_n466), .B2(new_n469), .ZN(new_n470));
  INV_X1    g045(.A(G2105), .ZN(new_n471));
  NAND4_X1  g046(.A1(new_n470), .A2(KEYINPUT71), .A3(G137), .A4(new_n471), .ZN(new_n472));
  NOR2_X1   g047(.A1(new_n463), .A2(KEYINPUT3), .ZN(new_n473));
  INV_X1    g048(.A(KEYINPUT70), .ZN(new_n474));
  OAI21_X1  g049(.A(new_n466), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  NAND4_X1  g050(.A1(new_n475), .A2(G137), .A3(new_n471), .A4(new_n464), .ZN(new_n476));
  INV_X1    g051(.A(KEYINPUT71), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  AND2_X1   g053(.A1(new_n472), .A2(new_n478), .ZN(new_n479));
  NOR2_X1   g054(.A1(new_n463), .A2(G2105), .ZN(new_n480));
  INV_X1    g055(.A(new_n480), .ZN(new_n481));
  INV_X1    g056(.A(G101), .ZN(new_n482));
  NOR2_X1   g057(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  INV_X1    g058(.A(new_n483), .ZN(new_n484));
  INV_X1    g059(.A(KEYINPUT68), .ZN(new_n485));
  AND3_X1   g060(.A1(new_n466), .A2(new_n468), .A3(new_n485), .ZN(new_n486));
  AOI21_X1  g061(.A(new_n485), .B1(new_n466), .B2(new_n468), .ZN(new_n487));
  OAI21_X1  g062(.A(G125), .B1(new_n486), .B2(new_n487), .ZN(new_n488));
  NAND2_X1  g063(.A1(G113), .A2(G2104), .ZN(new_n489));
  XNOR2_X1  g064(.A(new_n489), .B(KEYINPUT69), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n488), .A2(new_n490), .ZN(new_n491));
  NAND2_X1  g066(.A1(new_n491), .A2(G2105), .ZN(new_n492));
  NAND3_X1  g067(.A1(new_n479), .A2(new_n484), .A3(new_n492), .ZN(new_n493));
  INV_X1    g068(.A(new_n493), .ZN(G160));
  NAND3_X1  g069(.A1(new_n475), .A2(new_n471), .A3(new_n464), .ZN(new_n495));
  INV_X1    g070(.A(G136), .ZN(new_n496));
  OR3_X1    g071(.A1(new_n495), .A2(KEYINPUT72), .A3(new_n496), .ZN(new_n497));
  NAND3_X1  g072(.A1(new_n475), .A2(G2105), .A3(new_n464), .ZN(new_n498));
  INV_X1    g073(.A(new_n498), .ZN(new_n499));
  NAND2_X1  g074(.A1(new_n499), .A2(G124), .ZN(new_n500));
  OAI21_X1  g075(.A(KEYINPUT72), .B1(new_n495), .B2(new_n496), .ZN(new_n501));
  OR2_X1    g076(.A1(G100), .A2(G2105), .ZN(new_n502));
  OAI211_X1 g077(.A(new_n502), .B(G2104), .C1(G112), .C2(new_n471), .ZN(new_n503));
  NAND4_X1  g078(.A1(new_n497), .A2(new_n500), .A3(new_n501), .A4(new_n503), .ZN(new_n504));
  INV_X1    g079(.A(new_n504), .ZN(G162));
  NAND4_X1  g080(.A1(new_n475), .A2(G126), .A3(G2105), .A4(new_n464), .ZN(new_n506));
  OR2_X1    g081(.A1(G102), .A2(G2105), .ZN(new_n507));
  OAI211_X1 g082(.A(new_n507), .B(G2104), .C1(G114), .C2(new_n471), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n506), .A2(new_n508), .ZN(new_n509));
  AND2_X1   g084(.A1(new_n471), .A2(G138), .ZN(new_n510));
  AOI21_X1  g085(.A(new_n474), .B1(new_n467), .B2(G2104), .ZN(new_n511));
  NOR2_X1   g086(.A1(new_n467), .A2(G2104), .ZN(new_n512));
  OAI211_X1 g087(.A(new_n464), .B(new_n510), .C1(new_n511), .C2(new_n512), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n513), .A2(KEYINPUT73), .ZN(new_n514));
  INV_X1    g089(.A(KEYINPUT73), .ZN(new_n515));
  NAND4_X1  g090(.A1(new_n475), .A2(new_n515), .A3(new_n464), .A4(new_n510), .ZN(new_n516));
  NAND3_X1  g091(.A1(new_n514), .A2(KEYINPUT4), .A3(new_n516), .ZN(new_n517));
  INV_X1    g092(.A(KEYINPUT4), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n510), .A2(new_n518), .ZN(new_n519));
  OAI21_X1  g094(.A(KEYINPUT68), .B1(new_n512), .B2(new_n473), .ZN(new_n520));
  NAND3_X1  g095(.A1(new_n466), .A2(new_n468), .A3(new_n485), .ZN(new_n521));
  AOI21_X1  g096(.A(new_n519), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  INV_X1    g097(.A(new_n522), .ZN(new_n523));
  AOI21_X1  g098(.A(new_n509), .B1(new_n517), .B2(new_n523), .ZN(G164));
  INV_X1    g099(.A(G543), .ZN(new_n525));
  NAND2_X1  g100(.A1(new_n525), .A2(KEYINPUT5), .ZN(new_n526));
  INV_X1    g101(.A(KEYINPUT5), .ZN(new_n527));
  NAND2_X1  g102(.A1(new_n527), .A2(G543), .ZN(new_n528));
  AND2_X1   g103(.A1(new_n526), .A2(new_n528), .ZN(new_n529));
  AOI22_X1  g104(.A1(new_n529), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n530));
  INV_X1    g105(.A(G651), .ZN(new_n531));
  NOR2_X1   g106(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  XNOR2_X1  g107(.A(KEYINPUT6), .B(G651), .ZN(new_n533));
  NAND2_X1  g108(.A1(new_n529), .A2(new_n533), .ZN(new_n534));
  INV_X1    g109(.A(G88), .ZN(new_n535));
  NAND2_X1  g110(.A1(new_n533), .A2(G543), .ZN(new_n536));
  INV_X1    g111(.A(G50), .ZN(new_n537));
  OAI22_X1  g112(.A1(new_n534), .A2(new_n535), .B1(new_n536), .B2(new_n537), .ZN(new_n538));
  OR2_X1    g113(.A1(new_n532), .A2(new_n538), .ZN(G303));
  INV_X1    g114(.A(G303), .ZN(G166));
  INV_X1    g115(.A(G89), .ZN(new_n541));
  INV_X1    g116(.A(G51), .ZN(new_n542));
  OAI22_X1  g117(.A1(new_n534), .A2(new_n541), .B1(new_n536), .B2(new_n542), .ZN(new_n543));
  NAND3_X1  g118(.A1(new_n529), .A2(G63), .A3(G651), .ZN(new_n544));
  NAND3_X1  g119(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n545));
  INV_X1    g120(.A(KEYINPUT7), .ZN(new_n546));
  OR2_X1    g121(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  NAND2_X1  g122(.A1(new_n545), .A2(new_n546), .ZN(new_n548));
  NAND3_X1  g123(.A1(new_n544), .A2(new_n547), .A3(new_n548), .ZN(new_n549));
  NOR2_X1   g124(.A1(new_n543), .A2(new_n549), .ZN(G168));
  AOI22_X1  g125(.A1(new_n529), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n551));
  NOR2_X1   g126(.A1(new_n551), .A2(new_n531), .ZN(new_n552));
  INV_X1    g127(.A(G90), .ZN(new_n553));
  INV_X1    g128(.A(G52), .ZN(new_n554));
  OAI22_X1  g129(.A1(new_n534), .A2(new_n553), .B1(new_n536), .B2(new_n554), .ZN(new_n555));
  NOR2_X1   g130(.A1(new_n552), .A2(new_n555), .ZN(G171));
  AOI22_X1  g131(.A1(new_n529), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n557));
  INV_X1    g132(.A(KEYINPUT74), .ZN(new_n558));
  AOI21_X1  g133(.A(new_n531), .B1(new_n557), .B2(new_n558), .ZN(new_n559));
  OAI21_X1  g134(.A(new_n559), .B1(new_n558), .B2(new_n557), .ZN(new_n560));
  AND2_X1   g135(.A1(new_n529), .A2(new_n533), .ZN(new_n561));
  INV_X1    g136(.A(new_n536), .ZN(new_n562));
  AOI22_X1  g137(.A1(new_n561), .A2(G81), .B1(new_n562), .B2(G43), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n560), .A2(new_n563), .ZN(new_n564));
  INV_X1    g139(.A(new_n564), .ZN(new_n565));
  NAND2_X1  g140(.A1(new_n565), .A2(G860), .ZN(G153));
  AND3_X1   g141(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n567), .A2(G36), .ZN(new_n568));
  XNOR2_X1  g143(.A(new_n568), .B(KEYINPUT75), .ZN(G176));
  NAND2_X1  g144(.A1(G1), .A2(G3), .ZN(new_n570));
  XNOR2_X1  g145(.A(new_n570), .B(KEYINPUT8), .ZN(new_n571));
  NAND2_X1  g146(.A1(new_n567), .A2(new_n571), .ZN(G188));
  NAND2_X1  g147(.A1(new_n562), .A2(G53), .ZN(new_n573));
  XOR2_X1   g148(.A(new_n573), .B(KEYINPUT9), .Z(new_n574));
  AOI22_X1  g149(.A1(new_n529), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n575));
  INV_X1    g150(.A(G91), .ZN(new_n576));
  OAI22_X1  g151(.A1(new_n575), .A2(new_n531), .B1(new_n576), .B2(new_n534), .ZN(new_n577));
  NOR2_X1   g152(.A1(new_n574), .A2(new_n577), .ZN(new_n578));
  INV_X1    g153(.A(new_n578), .ZN(G299));
  OR2_X1    g154(.A1(new_n552), .A2(new_n555), .ZN(G301));
  INV_X1    g155(.A(G168), .ZN(G286));
  NAND2_X1  g156(.A1(new_n561), .A2(G87), .ZN(new_n582));
  NAND3_X1  g157(.A1(new_n562), .A2(KEYINPUT76), .A3(G49), .ZN(new_n583));
  INV_X1    g158(.A(KEYINPUT76), .ZN(new_n584));
  INV_X1    g159(.A(G49), .ZN(new_n585));
  OAI21_X1  g160(.A(new_n584), .B1(new_n536), .B2(new_n585), .ZN(new_n586));
  OAI21_X1  g161(.A(G651), .B1(new_n529), .B2(G74), .ZN(new_n587));
  NAND4_X1  g162(.A1(new_n582), .A2(new_n583), .A3(new_n586), .A4(new_n587), .ZN(G288));
  AOI22_X1  g163(.A1(new_n529), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n589));
  NOR2_X1   g164(.A1(new_n589), .A2(new_n531), .ZN(new_n590));
  INV_X1    g165(.A(G86), .ZN(new_n591));
  INV_X1    g166(.A(G48), .ZN(new_n592));
  OAI22_X1  g167(.A1(new_n534), .A2(new_n591), .B1(new_n536), .B2(new_n592), .ZN(new_n593));
  NOR2_X1   g168(.A1(new_n590), .A2(new_n593), .ZN(new_n594));
  INV_X1    g169(.A(new_n594), .ZN(G305));
  AOI22_X1  g170(.A1(new_n529), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n596));
  NOR2_X1   g171(.A1(new_n596), .A2(new_n531), .ZN(new_n597));
  INV_X1    g172(.A(G85), .ZN(new_n598));
  INV_X1    g173(.A(G47), .ZN(new_n599));
  OAI22_X1  g174(.A1(new_n534), .A2(new_n598), .B1(new_n536), .B2(new_n599), .ZN(new_n600));
  NOR2_X1   g175(.A1(new_n597), .A2(new_n600), .ZN(new_n601));
  INV_X1    g176(.A(new_n601), .ZN(G290));
  NAND2_X1  g177(.A1(G301), .A2(G868), .ZN(new_n603));
  NAND2_X1  g178(.A1(G79), .A2(G543), .ZN(new_n604));
  NAND2_X1  g179(.A1(new_n526), .A2(new_n528), .ZN(new_n605));
  INV_X1    g180(.A(G66), .ZN(new_n606));
  OAI21_X1  g181(.A(new_n604), .B1(new_n605), .B2(new_n606), .ZN(new_n607));
  INV_X1    g182(.A(KEYINPUT77), .ZN(new_n608));
  OR2_X1    g183(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  AOI21_X1  g184(.A(new_n531), .B1(new_n607), .B2(new_n608), .ZN(new_n610));
  AOI22_X1  g185(.A1(new_n609), .A2(new_n610), .B1(G54), .B2(new_n562), .ZN(new_n611));
  INV_X1    g186(.A(KEYINPUT78), .ZN(new_n612));
  XNOR2_X1  g187(.A(new_n611), .B(new_n612), .ZN(new_n613));
  NAND2_X1  g188(.A1(new_n561), .A2(G92), .ZN(new_n614));
  XOR2_X1   g189(.A(new_n614), .B(KEYINPUT10), .Z(new_n615));
  AND2_X1   g190(.A1(new_n613), .A2(new_n615), .ZN(new_n616));
  OAI21_X1  g191(.A(new_n603), .B1(new_n616), .B2(G868), .ZN(G321));
  XOR2_X1   g192(.A(G321), .B(KEYINPUT79), .Z(G284));
  NAND2_X1  g193(.A1(G286), .A2(G868), .ZN(new_n619));
  OAI21_X1  g194(.A(new_n619), .B1(new_n578), .B2(G868), .ZN(G297));
  OAI21_X1  g195(.A(new_n619), .B1(new_n578), .B2(G868), .ZN(G280));
  NAND2_X1  g196(.A1(new_n613), .A2(new_n615), .ZN(new_n622));
  INV_X1    g197(.A(G860), .ZN(new_n623));
  AOI21_X1  g198(.A(new_n622), .B1(G559), .B2(new_n623), .ZN(new_n624));
  XOR2_X1   g199(.A(new_n624), .B(KEYINPUT80), .Z(G148));
  INV_X1    g200(.A(G868), .ZN(new_n626));
  NAND2_X1  g201(.A1(new_n564), .A2(new_n626), .ZN(new_n627));
  NOR2_X1   g202(.A1(new_n622), .A2(G559), .ZN(new_n628));
  OAI21_X1  g203(.A(new_n627), .B1(new_n628), .B2(new_n626), .ZN(G323));
  XNOR2_X1  g204(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g205(.A1(new_n520), .A2(new_n521), .ZN(new_n631));
  NAND2_X1  g206(.A1(new_n631), .A2(new_n480), .ZN(new_n632));
  XNOR2_X1  g207(.A(new_n632), .B(KEYINPUT12), .ZN(new_n633));
  XNOR2_X1  g208(.A(new_n633), .B(KEYINPUT13), .ZN(new_n634));
  XNOR2_X1  g209(.A(new_n634), .B(G2100), .ZN(new_n635));
  INV_X1    g210(.A(G123), .ZN(new_n636));
  OR3_X1    g211(.A1(new_n498), .A2(KEYINPUT81), .A3(new_n636), .ZN(new_n637));
  INV_X1    g212(.A(new_n495), .ZN(new_n638));
  NAND2_X1  g213(.A1(new_n638), .A2(G135), .ZN(new_n639));
  OAI21_X1  g214(.A(KEYINPUT81), .B1(new_n498), .B2(new_n636), .ZN(new_n640));
  OAI21_X1  g215(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n641));
  INV_X1    g216(.A(KEYINPUT82), .ZN(new_n642));
  INV_X1    g217(.A(G111), .ZN(new_n643));
  AOI22_X1  g218(.A1(new_n641), .A2(new_n642), .B1(new_n643), .B2(G2105), .ZN(new_n644));
  OAI21_X1  g219(.A(new_n644), .B1(new_n642), .B2(new_n641), .ZN(new_n645));
  NAND4_X1  g220(.A1(new_n637), .A2(new_n639), .A3(new_n640), .A4(new_n645), .ZN(new_n646));
  XOR2_X1   g221(.A(new_n646), .B(G2096), .Z(new_n647));
  NAND2_X1  g222(.A1(new_n635), .A2(new_n647), .ZN(G156));
  XNOR2_X1  g223(.A(KEYINPUT15), .B(G2435), .ZN(new_n649));
  XNOR2_X1  g224(.A(KEYINPUT84), .B(G2438), .ZN(new_n650));
  XNOR2_X1  g225(.A(new_n649), .B(new_n650), .ZN(new_n651));
  XOR2_X1   g226(.A(G2427), .B(G2430), .Z(new_n652));
  OR2_X1    g227(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  NAND2_X1  g228(.A1(new_n651), .A2(new_n652), .ZN(new_n654));
  NAND3_X1  g229(.A1(new_n653), .A2(KEYINPUT14), .A3(new_n654), .ZN(new_n655));
  XNOR2_X1  g230(.A(new_n655), .B(KEYINPUT85), .ZN(new_n656));
  XOR2_X1   g231(.A(G2443), .B(G2446), .Z(new_n657));
  XNOR2_X1  g232(.A(new_n656), .B(new_n657), .ZN(new_n658));
  XOR2_X1   g233(.A(G2451), .B(G2454), .Z(new_n659));
  XNOR2_X1  g234(.A(KEYINPUT83), .B(KEYINPUT16), .ZN(new_n660));
  XNOR2_X1  g235(.A(new_n659), .B(new_n660), .ZN(new_n661));
  XNOR2_X1  g236(.A(new_n658), .B(new_n661), .ZN(new_n662));
  XNOR2_X1  g237(.A(G1341), .B(G1348), .ZN(new_n663));
  OR3_X1    g238(.A1(new_n662), .A2(KEYINPUT86), .A3(new_n663), .ZN(new_n664));
  OAI21_X1  g239(.A(KEYINPUT86), .B1(new_n662), .B2(new_n663), .ZN(new_n665));
  INV_X1    g240(.A(G14), .ZN(new_n666));
  AOI21_X1  g241(.A(new_n666), .B1(new_n662), .B2(new_n663), .ZN(new_n667));
  NAND3_X1  g242(.A1(new_n664), .A2(new_n665), .A3(new_n667), .ZN(new_n668));
  INV_X1    g243(.A(new_n668), .ZN(G401));
  XOR2_X1   g244(.A(G2072), .B(G2078), .Z(new_n670));
  XOR2_X1   g245(.A(G2084), .B(G2090), .Z(new_n671));
  INV_X1    g246(.A(new_n671), .ZN(new_n672));
  XOR2_X1   g247(.A(G2067), .B(G2678), .Z(new_n673));
  OR2_X1    g248(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  XNOR2_X1  g249(.A(KEYINPUT87), .B(KEYINPUT18), .ZN(new_n675));
  AOI21_X1  g250(.A(new_n670), .B1(new_n674), .B2(new_n675), .ZN(new_n676));
  XOR2_X1   g251(.A(G2096), .B(G2100), .Z(new_n677));
  XNOR2_X1  g252(.A(new_n676), .B(new_n677), .ZN(new_n678));
  INV_X1    g253(.A(KEYINPUT17), .ZN(new_n679));
  AOI21_X1  g254(.A(new_n679), .B1(new_n672), .B2(new_n673), .ZN(new_n680));
  AOI21_X1  g255(.A(new_n675), .B1(new_n674), .B2(new_n680), .ZN(new_n681));
  XNOR2_X1  g256(.A(new_n678), .B(new_n681), .ZN(G227));
  XNOR2_X1  g257(.A(G1971), .B(G1976), .ZN(new_n683));
  XNOR2_X1  g258(.A(new_n683), .B(KEYINPUT19), .ZN(new_n684));
  INV_X1    g259(.A(new_n684), .ZN(new_n685));
  XOR2_X1   g260(.A(G1956), .B(G2474), .Z(new_n686));
  XOR2_X1   g261(.A(G1961), .B(G1966), .Z(new_n687));
  AND2_X1   g262(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  NOR2_X1   g263(.A1(new_n686), .A2(new_n687), .ZN(new_n689));
  OR3_X1    g264(.A1(new_n685), .A2(new_n688), .A3(new_n689), .ZN(new_n690));
  NAND2_X1  g265(.A1(new_n685), .A2(new_n689), .ZN(new_n691));
  INV_X1    g266(.A(KEYINPUT20), .ZN(new_n692));
  OR2_X1    g267(.A1(new_n688), .A2(KEYINPUT88), .ZN(new_n693));
  NAND2_X1  g268(.A1(new_n688), .A2(KEYINPUT88), .ZN(new_n694));
  NAND3_X1  g269(.A1(new_n693), .A2(new_n685), .A3(new_n694), .ZN(new_n695));
  OAI211_X1 g270(.A(new_n690), .B(new_n691), .C1(new_n692), .C2(new_n695), .ZN(new_n696));
  AOI21_X1  g271(.A(new_n696), .B1(new_n692), .B2(new_n695), .ZN(new_n697));
  XNOR2_X1  g272(.A(KEYINPUT89), .B(KEYINPUT90), .ZN(new_n698));
  XNOR2_X1  g273(.A(new_n697), .B(new_n698), .ZN(new_n699));
  XOR2_X1   g274(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n700));
  XNOR2_X1  g275(.A(G1981), .B(G1986), .ZN(new_n701));
  XNOR2_X1  g276(.A(new_n700), .B(new_n701), .ZN(new_n702));
  XNOR2_X1  g277(.A(G1991), .B(G1996), .ZN(new_n703));
  XNOR2_X1  g278(.A(new_n702), .B(new_n703), .ZN(new_n704));
  XNOR2_X1  g279(.A(new_n699), .B(new_n704), .ZN(G229));
  INV_X1    g280(.A(KEYINPUT92), .ZN(new_n706));
  XNOR2_X1  g281(.A(G288), .B(new_n706), .ZN(new_n707));
  MUX2_X1   g282(.A(G23), .B(new_n707), .S(G16), .Z(new_n708));
  XOR2_X1   g283(.A(KEYINPUT33), .B(G1976), .Z(new_n709));
  OR2_X1    g284(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  NAND2_X1  g285(.A1(new_n708), .A2(new_n709), .ZN(new_n711));
  INV_X1    g286(.A(G16), .ZN(new_n712));
  NAND2_X1  g287(.A1(new_n712), .A2(G22), .ZN(new_n713));
  OAI21_X1  g288(.A(new_n713), .B1(G166), .B2(new_n712), .ZN(new_n714));
  INV_X1    g289(.A(G1971), .ZN(new_n715));
  XNOR2_X1  g290(.A(new_n714), .B(new_n715), .ZN(new_n716));
  NAND2_X1  g291(.A1(new_n712), .A2(G6), .ZN(new_n717));
  OAI21_X1  g292(.A(new_n717), .B1(new_n594), .B2(new_n712), .ZN(new_n718));
  XOR2_X1   g293(.A(KEYINPUT32), .B(G1981), .Z(new_n719));
  XNOR2_X1  g294(.A(new_n718), .B(new_n719), .ZN(new_n720));
  NAND4_X1  g295(.A1(new_n710), .A2(new_n711), .A3(new_n716), .A4(new_n720), .ZN(new_n721));
  XOR2_X1   g296(.A(new_n721), .B(KEYINPUT34), .Z(new_n722));
  INV_X1    g297(.A(G29), .ZN(new_n723));
  NAND2_X1  g298(.A1(new_n723), .A2(G25), .ZN(new_n724));
  NAND2_X1  g299(.A1(new_n499), .A2(G119), .ZN(new_n725));
  NAND2_X1  g300(.A1(new_n638), .A2(G131), .ZN(new_n726));
  OR2_X1    g301(.A1(G95), .A2(G2105), .ZN(new_n727));
  OAI211_X1 g302(.A(new_n727), .B(G2104), .C1(G107), .C2(new_n471), .ZN(new_n728));
  NAND3_X1  g303(.A1(new_n725), .A2(new_n726), .A3(new_n728), .ZN(new_n729));
  INV_X1    g304(.A(new_n729), .ZN(new_n730));
  OAI21_X1  g305(.A(new_n724), .B1(new_n730), .B2(new_n723), .ZN(new_n731));
  XNOR2_X1  g306(.A(new_n731), .B(KEYINPUT91), .ZN(new_n732));
  XOR2_X1   g307(.A(KEYINPUT35), .B(G1991), .Z(new_n733));
  XNOR2_X1  g308(.A(new_n732), .B(new_n733), .ZN(new_n734));
  NAND2_X1  g309(.A1(new_n712), .A2(G24), .ZN(new_n735));
  OAI21_X1  g310(.A(new_n735), .B1(new_n601), .B2(new_n712), .ZN(new_n736));
  OAI21_X1  g311(.A(KEYINPUT93), .B1(new_n736), .B2(G1986), .ZN(new_n737));
  AOI21_X1  g312(.A(new_n737), .B1(G1986), .B2(new_n736), .ZN(new_n738));
  NAND3_X1  g313(.A1(new_n722), .A2(new_n734), .A3(new_n738), .ZN(new_n739));
  INV_X1    g314(.A(KEYINPUT36), .ZN(new_n740));
  AND2_X1   g315(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  INV_X1    g316(.A(KEYINPUT23), .ZN(new_n742));
  AND2_X1   g317(.A1(new_n712), .A2(G20), .ZN(new_n743));
  AOI211_X1 g318(.A(new_n742), .B(new_n743), .C1(G299), .C2(G16), .ZN(new_n744));
  AOI21_X1  g319(.A(new_n744), .B1(new_n742), .B2(new_n743), .ZN(new_n745));
  XOR2_X1   g320(.A(KEYINPUT99), .B(G1956), .Z(new_n746));
  XNOR2_X1  g321(.A(new_n745), .B(new_n746), .ZN(new_n747));
  NOR2_X1   g322(.A1(G27), .A2(G29), .ZN(new_n748));
  AOI21_X1  g323(.A(new_n748), .B1(G164), .B2(G29), .ZN(new_n749));
  XOR2_X1   g324(.A(KEYINPUT98), .B(G2078), .Z(new_n750));
  XNOR2_X1  g325(.A(new_n749), .B(new_n750), .ZN(new_n751));
  NAND2_X1  g326(.A1(new_n723), .A2(G33), .ZN(new_n752));
  NAND2_X1  g327(.A1(new_n631), .A2(G127), .ZN(new_n753));
  NAND2_X1  g328(.A1(G115), .A2(G2104), .ZN(new_n754));
  AOI21_X1  g329(.A(new_n471), .B1(new_n753), .B2(new_n754), .ZN(new_n755));
  NAND2_X1  g330(.A1(new_n480), .A2(G103), .ZN(new_n756));
  INV_X1    g331(.A(KEYINPUT25), .ZN(new_n757));
  XNOR2_X1  g332(.A(new_n756), .B(new_n757), .ZN(new_n758));
  INV_X1    g333(.A(G139), .ZN(new_n759));
  OAI21_X1  g334(.A(new_n758), .B1(new_n759), .B2(new_n495), .ZN(new_n760));
  NOR2_X1   g335(.A1(new_n755), .A2(new_n760), .ZN(new_n761));
  OAI21_X1  g336(.A(new_n752), .B1(new_n761), .B2(new_n723), .ZN(new_n762));
  XOR2_X1   g337(.A(new_n762), .B(G2072), .Z(new_n763));
  NAND2_X1  g338(.A1(new_n712), .A2(G19), .ZN(new_n764));
  OAI21_X1  g339(.A(new_n764), .B1(new_n565), .B2(new_n712), .ZN(new_n765));
  XNOR2_X1  g340(.A(new_n765), .B(G1341), .ZN(new_n766));
  NOR2_X1   g341(.A1(G5), .A2(G16), .ZN(new_n767));
  AOI21_X1  g342(.A(new_n767), .B1(G171), .B2(G16), .ZN(new_n768));
  INV_X1    g343(.A(G1961), .ZN(new_n769));
  XNOR2_X1  g344(.A(new_n768), .B(new_n769), .ZN(new_n770));
  OAI21_X1  g345(.A(new_n770), .B1(new_n723), .B2(new_n646), .ZN(new_n771));
  NOR2_X1   g346(.A1(G16), .A2(G21), .ZN(new_n772));
  AOI21_X1  g347(.A(new_n772), .B1(G168), .B2(G16), .ZN(new_n773));
  NOR2_X1   g348(.A1(new_n773), .A2(G1966), .ZN(new_n774));
  NAND2_X1  g349(.A1(new_n773), .A2(G1966), .ZN(new_n775));
  NOR2_X1   g350(.A1(KEYINPUT31), .A2(G11), .ZN(new_n776));
  AND2_X1   g351(.A1(KEYINPUT31), .A2(G11), .ZN(new_n777));
  INV_X1    g352(.A(KEYINPUT30), .ZN(new_n778));
  AND2_X1   g353(.A1(new_n778), .A2(G28), .ZN(new_n779));
  OAI21_X1  g354(.A(new_n723), .B1(new_n778), .B2(G28), .ZN(new_n780));
  OAI221_X1 g355(.A(new_n775), .B1(new_n776), .B2(new_n777), .C1(new_n779), .C2(new_n780), .ZN(new_n781));
  NOR4_X1   g356(.A1(new_n766), .A2(new_n771), .A3(new_n774), .A4(new_n781), .ZN(new_n782));
  NAND4_X1  g357(.A1(new_n747), .A2(new_n751), .A3(new_n763), .A4(new_n782), .ZN(new_n783));
  NAND3_X1  g358(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n784));
  INV_X1    g359(.A(KEYINPUT26), .ZN(new_n785));
  OR2_X1    g360(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  NAND2_X1  g361(.A1(new_n784), .A2(new_n785), .ZN(new_n787));
  AOI22_X1  g362(.A1(new_n786), .A2(new_n787), .B1(G105), .B2(new_n480), .ZN(new_n788));
  INV_X1    g363(.A(G141), .ZN(new_n789));
  INV_X1    g364(.A(G129), .ZN(new_n790));
  OAI221_X1 g365(.A(new_n788), .B1(new_n495), .B2(new_n789), .C1(new_n790), .C2(new_n498), .ZN(new_n791));
  MUX2_X1   g366(.A(G32), .B(new_n791), .S(G29), .Z(new_n792));
  XOR2_X1   g367(.A(new_n792), .B(KEYINPUT97), .Z(new_n793));
  XOR2_X1   g368(.A(KEYINPUT27), .B(G1996), .Z(new_n794));
  OR2_X1    g369(.A1(new_n793), .A2(new_n794), .ZN(new_n795));
  NAND2_X1  g370(.A1(new_n793), .A2(new_n794), .ZN(new_n796));
  NAND2_X1  g371(.A1(new_n723), .A2(G35), .ZN(new_n797));
  OAI21_X1  g372(.A(new_n797), .B1(G162), .B2(new_n723), .ZN(new_n798));
  XOR2_X1   g373(.A(KEYINPUT29), .B(G2090), .Z(new_n799));
  XNOR2_X1  g374(.A(new_n798), .B(new_n799), .ZN(new_n800));
  INV_X1    g375(.A(KEYINPUT24), .ZN(new_n801));
  OAI21_X1  g376(.A(new_n723), .B1(new_n801), .B2(G34), .ZN(new_n802));
  INV_X1    g377(.A(KEYINPUT95), .ZN(new_n803));
  AOI22_X1  g378(.A1(new_n802), .A2(new_n803), .B1(new_n801), .B2(G34), .ZN(new_n804));
  OAI21_X1  g379(.A(new_n804), .B1(new_n803), .B2(new_n802), .ZN(new_n805));
  XOR2_X1   g380(.A(new_n805), .B(KEYINPUT96), .Z(new_n806));
  OAI21_X1  g381(.A(new_n806), .B1(new_n493), .B2(new_n723), .ZN(new_n807));
  XNOR2_X1  g382(.A(new_n807), .B(G2084), .ZN(new_n808));
  NAND4_X1  g383(.A1(new_n795), .A2(new_n796), .A3(new_n800), .A4(new_n808), .ZN(new_n809));
  NOR2_X1   g384(.A1(new_n783), .A2(new_n809), .ZN(new_n810));
  NAND2_X1  g385(.A1(new_n723), .A2(G26), .ZN(new_n811));
  XNOR2_X1  g386(.A(new_n811), .B(KEYINPUT28), .ZN(new_n812));
  NAND2_X1  g387(.A1(new_n499), .A2(G128), .ZN(new_n813));
  NAND2_X1  g388(.A1(new_n638), .A2(G140), .ZN(new_n814));
  NOR2_X1   g389(.A1(new_n471), .A2(G116), .ZN(new_n815));
  OAI21_X1  g390(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n816));
  OAI211_X1 g391(.A(new_n813), .B(new_n814), .C1(new_n815), .C2(new_n816), .ZN(new_n817));
  NAND2_X1  g392(.A1(new_n817), .A2(G29), .ZN(new_n818));
  AND2_X1   g393(.A1(new_n818), .A2(KEYINPUT94), .ZN(new_n819));
  NOR2_X1   g394(.A1(new_n818), .A2(KEYINPUT94), .ZN(new_n820));
  OAI21_X1  g395(.A(new_n812), .B1(new_n819), .B2(new_n820), .ZN(new_n821));
  INV_X1    g396(.A(G2067), .ZN(new_n822));
  XNOR2_X1  g397(.A(new_n821), .B(new_n822), .ZN(new_n823));
  NAND2_X1  g398(.A1(new_n616), .A2(G16), .ZN(new_n824));
  OAI21_X1  g399(.A(new_n824), .B1(G4), .B2(G16), .ZN(new_n825));
  XNOR2_X1  g400(.A(new_n825), .B(G1348), .ZN(new_n826));
  NAND3_X1  g401(.A1(new_n810), .A2(new_n823), .A3(new_n826), .ZN(new_n827));
  NOR2_X1   g402(.A1(new_n739), .A2(new_n740), .ZN(new_n828));
  NOR3_X1   g403(.A1(new_n741), .A2(new_n827), .A3(new_n828), .ZN(G311));
  INV_X1    g404(.A(G311), .ZN(G150));
  NAND2_X1  g405(.A1(new_n616), .A2(G559), .ZN(new_n831));
  XOR2_X1   g406(.A(KEYINPUT38), .B(KEYINPUT39), .Z(new_n832));
  XOR2_X1   g407(.A(new_n831), .B(new_n832), .Z(new_n833));
  XOR2_X1   g408(.A(KEYINPUT100), .B(G55), .Z(new_n834));
  AOI22_X1  g409(.A1(new_n561), .A2(G93), .B1(new_n562), .B2(new_n834), .ZN(new_n835));
  XNOR2_X1  g410(.A(new_n835), .B(KEYINPUT101), .ZN(new_n836));
  AOI22_X1  g411(.A1(new_n529), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n837));
  OR2_X1    g412(.A1(new_n837), .A2(new_n531), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n836), .A2(new_n838), .ZN(new_n839));
  NAND2_X1  g414(.A1(new_n839), .A2(new_n565), .ZN(new_n840));
  NAND3_X1  g415(.A1(new_n836), .A2(new_n564), .A3(new_n838), .ZN(new_n841));
  NAND2_X1  g416(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  OR2_X1    g417(.A1(new_n833), .A2(new_n842), .ZN(new_n843));
  NAND2_X1  g418(.A1(new_n833), .A2(new_n842), .ZN(new_n844));
  NAND3_X1  g419(.A1(new_n843), .A2(new_n623), .A3(new_n844), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n839), .A2(G860), .ZN(new_n846));
  XOR2_X1   g421(.A(new_n846), .B(KEYINPUT37), .Z(new_n847));
  NAND2_X1  g422(.A1(new_n845), .A2(new_n847), .ZN(G145));
  XNOR2_X1  g423(.A(new_n761), .B(new_n791), .ZN(new_n849));
  XNOR2_X1  g424(.A(new_n817), .B(KEYINPUT104), .ZN(new_n850));
  XNOR2_X1  g425(.A(new_n849), .B(new_n850), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n517), .A2(new_n523), .ZN(new_n852));
  INV_X1    g427(.A(KEYINPUT103), .ZN(new_n853));
  INV_X1    g428(.A(new_n509), .ZN(new_n854));
  NAND3_X1  g429(.A1(new_n852), .A2(new_n853), .A3(new_n854), .ZN(new_n855));
  AOI21_X1  g430(.A(new_n518), .B1(new_n513), .B2(KEYINPUT73), .ZN(new_n856));
  AOI21_X1  g431(.A(new_n522), .B1(new_n856), .B2(new_n516), .ZN(new_n857));
  OAI21_X1  g432(.A(KEYINPUT103), .B1(new_n857), .B2(new_n509), .ZN(new_n858));
  NAND2_X1  g433(.A1(new_n855), .A2(new_n858), .ZN(new_n859));
  OR2_X1    g434(.A1(new_n851), .A2(new_n859), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n851), .A2(new_n859), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n638), .A2(G142), .ZN(new_n863));
  NOR2_X1   g438(.A1(new_n471), .A2(G118), .ZN(new_n864));
  OAI21_X1  g439(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n865));
  OAI21_X1  g440(.A(new_n863), .B1(new_n864), .B2(new_n865), .ZN(new_n866));
  AOI21_X1  g441(.A(new_n866), .B1(G130), .B2(new_n499), .ZN(new_n867));
  XOR2_X1   g442(.A(new_n867), .B(new_n633), .Z(new_n868));
  XNOR2_X1  g443(.A(new_n868), .B(new_n730), .ZN(new_n869));
  INV_X1    g444(.A(new_n869), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n862), .A2(new_n870), .ZN(new_n871));
  INV_X1    g446(.A(KEYINPUT105), .ZN(new_n872));
  NAND3_X1  g447(.A1(new_n869), .A2(new_n860), .A3(new_n861), .ZN(new_n873));
  NAND3_X1  g448(.A1(new_n871), .A2(new_n872), .A3(new_n873), .ZN(new_n874));
  XNOR2_X1  g449(.A(new_n493), .B(KEYINPUT102), .ZN(new_n875));
  XNOR2_X1  g450(.A(new_n875), .B(G162), .ZN(new_n876));
  XNOR2_X1  g451(.A(new_n876), .B(new_n646), .ZN(new_n877));
  AOI21_X1  g452(.A(new_n869), .B1(new_n860), .B2(new_n861), .ZN(new_n878));
  AOI21_X1  g453(.A(new_n877), .B1(new_n878), .B2(KEYINPUT105), .ZN(new_n879));
  AOI21_X1  g454(.A(G37), .B1(new_n874), .B2(new_n879), .ZN(new_n880));
  INV_X1    g455(.A(KEYINPUT106), .ZN(new_n881));
  AND2_X1   g456(.A1(new_n871), .A2(new_n873), .ZN(new_n882));
  AOI21_X1  g457(.A(new_n881), .B1(new_n882), .B2(new_n877), .ZN(new_n883));
  AND4_X1   g458(.A1(new_n881), .A2(new_n871), .A3(new_n873), .A4(new_n877), .ZN(new_n884));
  OAI21_X1  g459(.A(new_n880), .B1(new_n883), .B2(new_n884), .ZN(new_n885));
  XNOR2_X1  g460(.A(new_n885), .B(KEYINPUT40), .ZN(G395));
  XNOR2_X1  g461(.A(G305), .B(G303), .ZN(new_n887));
  XNOR2_X1  g462(.A(new_n707), .B(new_n601), .ZN(new_n888));
  INV_X1    g463(.A(KEYINPUT108), .ZN(new_n889));
  AND2_X1   g464(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  NOR2_X1   g465(.A1(new_n888), .A2(new_n889), .ZN(new_n891));
  OAI21_X1  g466(.A(new_n887), .B1(new_n890), .B2(new_n891), .ZN(new_n892));
  OAI21_X1  g467(.A(new_n892), .B1(new_n891), .B2(new_n887), .ZN(new_n893));
  INV_X1    g468(.A(KEYINPUT42), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n894), .A2(KEYINPUT109), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n893), .A2(new_n895), .ZN(new_n896));
  INV_X1    g471(.A(new_n896), .ZN(new_n897));
  NOR2_X1   g472(.A1(new_n894), .A2(KEYINPUT109), .ZN(new_n898));
  NOR2_X1   g473(.A1(new_n622), .A2(new_n578), .ZN(new_n899));
  INV_X1    g474(.A(new_n899), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n622), .A2(new_n578), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  INV_X1    g477(.A(KEYINPUT41), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  INV_X1    g479(.A(new_n901), .ZN(new_n905));
  NOR2_X1   g480(.A1(new_n905), .A2(new_n899), .ZN(new_n906));
  NAND2_X1  g481(.A1(new_n906), .A2(KEYINPUT41), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n842), .A2(KEYINPUT107), .ZN(new_n908));
  INV_X1    g483(.A(KEYINPUT107), .ZN(new_n909));
  NAND3_X1  g484(.A1(new_n840), .A2(new_n909), .A3(new_n841), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n908), .A2(new_n910), .ZN(new_n911));
  INV_X1    g486(.A(new_n628), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  NAND3_X1  g488(.A1(new_n908), .A2(new_n628), .A3(new_n910), .ZN(new_n914));
  AOI22_X1  g489(.A1(new_n904), .A2(new_n907), .B1(new_n913), .B2(new_n914), .ZN(new_n915));
  AND3_X1   g490(.A1(new_n913), .A2(new_n902), .A3(new_n914), .ZN(new_n916));
  OAI21_X1  g491(.A(new_n898), .B1(new_n915), .B2(new_n916), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n907), .A2(new_n904), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n913), .A2(new_n914), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  INV_X1    g495(.A(new_n898), .ZN(new_n921));
  NAND3_X1  g496(.A1(new_n913), .A2(new_n902), .A3(new_n914), .ZN(new_n922));
  NAND3_X1  g497(.A1(new_n920), .A2(new_n921), .A3(new_n922), .ZN(new_n923));
  NAND3_X1  g498(.A1(new_n897), .A2(new_n917), .A3(new_n923), .ZN(new_n924));
  INV_X1    g499(.A(new_n924), .ZN(new_n925));
  AOI21_X1  g500(.A(new_n897), .B1(new_n917), .B2(new_n923), .ZN(new_n926));
  OAI21_X1  g501(.A(G868), .B1(new_n925), .B2(new_n926), .ZN(new_n927));
  INV_X1    g502(.A(KEYINPUT110), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n839), .A2(new_n626), .ZN(new_n929));
  NAND3_X1  g504(.A1(new_n927), .A2(new_n928), .A3(new_n929), .ZN(new_n930));
  NOR3_X1   g505(.A1(new_n915), .A2(new_n916), .A3(new_n898), .ZN(new_n931));
  AOI21_X1  g506(.A(new_n921), .B1(new_n920), .B2(new_n922), .ZN(new_n932));
  OAI21_X1  g507(.A(new_n896), .B1(new_n931), .B2(new_n932), .ZN(new_n933));
  AOI21_X1  g508(.A(new_n626), .B1(new_n933), .B2(new_n924), .ZN(new_n934));
  INV_X1    g509(.A(new_n929), .ZN(new_n935));
  OAI21_X1  g510(.A(KEYINPUT110), .B1(new_n934), .B2(new_n935), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n930), .A2(new_n936), .ZN(G295));
  NAND2_X1  g512(.A1(new_n927), .A2(new_n929), .ZN(G331));
  INV_X1    g513(.A(new_n893), .ZN(new_n939));
  INV_X1    g514(.A(KEYINPUT111), .ZN(new_n940));
  OAI21_X1  g515(.A(G168), .B1(G301), .B2(new_n940), .ZN(new_n941));
  NOR2_X1   g516(.A1(G171), .A2(KEYINPUT111), .ZN(new_n942));
  XOR2_X1   g517(.A(new_n941), .B(new_n942), .Z(new_n943));
  NAND2_X1  g518(.A1(new_n943), .A2(new_n842), .ZN(new_n944));
  XNOR2_X1  g519(.A(new_n941), .B(new_n942), .ZN(new_n945));
  NAND3_X1  g520(.A1(new_n945), .A2(new_n840), .A3(new_n841), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n944), .A2(new_n946), .ZN(new_n947));
  INV_X1    g522(.A(KEYINPUT112), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n944), .A2(KEYINPUT112), .ZN(new_n950));
  NAND3_X1  g525(.A1(new_n949), .A2(new_n902), .A3(new_n950), .ZN(new_n951));
  INV_X1    g526(.A(new_n951), .ZN(new_n952));
  AOI22_X1  g527(.A1(new_n907), .A2(new_n904), .B1(new_n944), .B2(new_n946), .ZN(new_n953));
  OAI21_X1  g528(.A(new_n939), .B1(new_n952), .B2(new_n953), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n954), .A2(KEYINPUT113), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n918), .A2(new_n947), .ZN(new_n956));
  AOI21_X1  g531(.A(new_n893), .B1(new_n956), .B2(new_n951), .ZN(new_n957));
  INV_X1    g532(.A(KEYINPUT113), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n957), .A2(new_n958), .ZN(new_n959));
  INV_X1    g534(.A(KEYINPUT43), .ZN(new_n960));
  NOR2_X1   g535(.A1(new_n947), .A2(new_n906), .ZN(new_n961));
  NAND2_X1  g536(.A1(new_n949), .A2(new_n950), .ZN(new_n962));
  AOI21_X1  g537(.A(new_n961), .B1(new_n962), .B2(new_n918), .ZN(new_n963));
  AOI21_X1  g538(.A(G37), .B1(new_n963), .B2(new_n893), .ZN(new_n964));
  NAND4_X1  g539(.A1(new_n955), .A2(new_n959), .A3(new_n960), .A4(new_n964), .ZN(new_n965));
  AOI22_X1  g540(.A1(new_n949), .A2(new_n950), .B1(new_n907), .B2(new_n904), .ZN(new_n966));
  OAI21_X1  g541(.A(new_n939), .B1(new_n966), .B2(new_n961), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n964), .A2(new_n967), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n968), .A2(KEYINPUT43), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n965), .A2(new_n969), .ZN(new_n970));
  INV_X1    g545(.A(KEYINPUT44), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n970), .A2(new_n971), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n962), .A2(new_n918), .ZN(new_n973));
  INV_X1    g548(.A(new_n961), .ZN(new_n974));
  NAND3_X1  g549(.A1(new_n973), .A2(new_n893), .A3(new_n974), .ZN(new_n975));
  INV_X1    g550(.A(G37), .ZN(new_n976));
  OAI211_X1 g551(.A(new_n975), .B(new_n976), .C1(new_n957), .C2(new_n958), .ZN(new_n977));
  NOR2_X1   g552(.A1(new_n954), .A2(KEYINPUT113), .ZN(new_n978));
  OAI21_X1  g553(.A(KEYINPUT43), .B1(new_n977), .B2(new_n978), .ZN(new_n979));
  NAND3_X1  g554(.A1(new_n964), .A2(new_n960), .A3(new_n967), .ZN(new_n980));
  INV_X1    g555(.A(KEYINPUT114), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n980), .A2(new_n981), .ZN(new_n982));
  NAND4_X1  g557(.A1(new_n964), .A2(KEYINPUT114), .A3(new_n960), .A4(new_n967), .ZN(new_n983));
  NAND4_X1  g558(.A1(new_n979), .A2(new_n982), .A3(KEYINPUT44), .A4(new_n983), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n972), .A2(new_n984), .ZN(G397));
  AOI21_X1  g560(.A(G1384), .B1(new_n855), .B2(new_n858), .ZN(new_n986));
  NOR2_X1   g561(.A1(new_n986), .A2(KEYINPUT45), .ZN(new_n987));
  INV_X1    g562(.A(new_n987), .ZN(new_n988));
  NAND4_X1  g563(.A1(new_n479), .A2(G40), .A3(new_n484), .A4(new_n492), .ZN(new_n989));
  NOR2_X1   g564(.A1(new_n988), .A2(new_n989), .ZN(new_n990));
  INV_X1    g565(.A(new_n990), .ZN(new_n991));
  NOR2_X1   g566(.A1(G290), .A2(G1986), .ZN(new_n992));
  INV_X1    g567(.A(new_n992), .ZN(new_n993));
  NOR2_X1   g568(.A1(new_n991), .A2(new_n993), .ZN(new_n994));
  OR2_X1    g569(.A1(new_n994), .A2(KEYINPUT48), .ZN(new_n995));
  XNOR2_X1  g570(.A(new_n817), .B(new_n822), .ZN(new_n996));
  INV_X1    g571(.A(G1996), .ZN(new_n997));
  XNOR2_X1  g572(.A(new_n791), .B(new_n997), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n996), .A2(new_n998), .ZN(new_n999));
  XOR2_X1   g574(.A(new_n729), .B(new_n733), .Z(new_n1000));
  OAI21_X1  g575(.A(new_n990), .B1(new_n999), .B2(new_n1000), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n995), .A2(new_n1001), .ZN(new_n1002));
  AOI21_X1  g577(.A(new_n1002), .B1(KEYINPUT48), .B2(new_n994), .ZN(new_n1003));
  INV_X1    g578(.A(KEYINPUT46), .ZN(new_n1004));
  OAI21_X1  g579(.A(new_n1004), .B1(new_n991), .B2(G1996), .ZN(new_n1005));
  NAND3_X1  g580(.A1(new_n990), .A2(KEYINPUT46), .A3(new_n997), .ZN(new_n1006));
  INV_X1    g581(.A(new_n996), .ZN(new_n1007));
  OAI21_X1  g582(.A(new_n990), .B1(new_n791), .B2(new_n1007), .ZN(new_n1008));
  NAND3_X1  g583(.A1(new_n1005), .A2(new_n1006), .A3(new_n1008), .ZN(new_n1009));
  XOR2_X1   g584(.A(new_n1009), .B(KEYINPUT47), .Z(new_n1010));
  NAND2_X1  g585(.A1(new_n730), .A2(new_n733), .ZN(new_n1011));
  OAI22_X1  g586(.A1(new_n999), .A2(new_n1011), .B1(G2067), .B2(new_n817), .ZN(new_n1012));
  AOI211_X1 g587(.A(new_n1003), .B(new_n1010), .C1(new_n990), .C2(new_n1012), .ZN(new_n1013));
  AOI22_X1  g588(.A1(G303), .A2(G8), .B1(KEYINPUT117), .B2(KEYINPUT55), .ZN(new_n1014));
  NOR2_X1   g589(.A1(KEYINPUT117), .A2(KEYINPUT55), .ZN(new_n1015));
  XNOR2_X1  g590(.A(new_n1014), .B(new_n1015), .ZN(new_n1016));
  INV_X1    g591(.A(KEYINPUT45), .ZN(new_n1017));
  AOI211_X1 g592(.A(new_n1017), .B(G1384), .C1(new_n855), .C2(new_n858), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n472), .A2(new_n478), .ZN(new_n1019));
  AOI21_X1  g594(.A(new_n471), .B1(new_n488), .B2(new_n490), .ZN(new_n1020));
  INV_X1    g595(.A(G40), .ZN(new_n1021));
  NOR4_X1   g596(.A1(new_n1019), .A2(new_n1020), .A3(new_n1021), .A4(new_n483), .ZN(new_n1022));
  NOR2_X1   g597(.A1(G164), .A2(G1384), .ZN(new_n1023));
  OAI21_X1  g598(.A(new_n1022), .B1(new_n1023), .B2(KEYINPUT45), .ZN(new_n1024));
  OAI21_X1  g599(.A(KEYINPUT116), .B1(new_n1018), .B2(new_n1024), .ZN(new_n1025));
  INV_X1    g600(.A(G1384), .ZN(new_n1026));
  NOR2_X1   g601(.A1(G164), .A2(new_n853), .ZN(new_n1027));
  NOR3_X1   g602(.A1(new_n857), .A2(KEYINPUT103), .A3(new_n509), .ZN(new_n1028));
  OAI211_X1 g603(.A(KEYINPUT45), .B(new_n1026), .C1(new_n1027), .C2(new_n1028), .ZN(new_n1029));
  OAI21_X1  g604(.A(new_n1026), .B1(new_n857), .B2(new_n509), .ZN(new_n1030));
  AOI21_X1  g605(.A(new_n989), .B1(new_n1017), .B2(new_n1030), .ZN(new_n1031));
  INV_X1    g606(.A(KEYINPUT116), .ZN(new_n1032));
  NAND3_X1  g607(.A1(new_n1029), .A2(new_n1031), .A3(new_n1032), .ZN(new_n1033));
  AOI21_X1  g608(.A(G1971), .B1(new_n1025), .B2(new_n1033), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n1030), .A2(KEYINPUT50), .ZN(new_n1035));
  INV_X1    g610(.A(KEYINPUT50), .ZN(new_n1036));
  OAI211_X1 g611(.A(new_n1036), .B(new_n1026), .C1(new_n857), .C2(new_n509), .ZN(new_n1037));
  NAND3_X1  g612(.A1(new_n1035), .A2(new_n1022), .A3(new_n1037), .ZN(new_n1038));
  NOR2_X1   g613(.A1(new_n1038), .A2(G2090), .ZN(new_n1039));
  OAI211_X1 g614(.A(G8), .B(new_n1016), .C1(new_n1034), .C2(new_n1039), .ZN(new_n1040));
  INV_X1    g615(.A(G1981), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n594), .A2(new_n1041), .ZN(new_n1042));
  OAI21_X1  g617(.A(G1981), .B1(new_n590), .B2(new_n593), .ZN(new_n1043));
  AND3_X1   g618(.A1(new_n1042), .A2(KEYINPUT49), .A3(new_n1043), .ZN(new_n1044));
  AOI21_X1  g619(.A(KEYINPUT49), .B1(new_n1042), .B2(new_n1043), .ZN(new_n1045));
  NOR2_X1   g620(.A1(new_n1044), .A2(new_n1045), .ZN(new_n1046));
  INV_X1    g621(.A(KEYINPUT118), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n1022), .A2(new_n1023), .ZN(new_n1048));
  AOI21_X1  g623(.A(new_n1047), .B1(new_n1048), .B2(G8), .ZN(new_n1049));
  OAI211_X1 g624(.A(new_n1047), .B(G8), .C1(new_n989), .C2(new_n1030), .ZN(new_n1050));
  INV_X1    g625(.A(new_n1050), .ZN(new_n1051));
  OAI21_X1  g626(.A(new_n1046), .B1(new_n1049), .B2(new_n1051), .ZN(new_n1052));
  INV_X1    g627(.A(G1976), .ZN(new_n1053));
  NOR2_X1   g628(.A1(new_n707), .A2(new_n1053), .ZN(new_n1054));
  OAI21_X1  g629(.A(G8), .B1(new_n989), .B2(new_n1030), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n1055), .A2(KEYINPUT118), .ZN(new_n1056));
  AOI21_X1  g631(.A(new_n1054), .B1(new_n1056), .B2(new_n1050), .ZN(new_n1057));
  INV_X1    g632(.A(KEYINPUT52), .ZN(new_n1058));
  OAI21_X1  g633(.A(new_n1052), .B1(new_n1057), .B2(new_n1058), .ZN(new_n1059));
  NAND2_X1  g634(.A1(G288), .A2(new_n1053), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n1060), .A2(new_n1058), .ZN(new_n1061));
  AOI211_X1 g636(.A(new_n1061), .B(new_n1054), .C1(new_n1056), .C2(new_n1050), .ZN(new_n1062));
  NOR2_X1   g637(.A1(new_n1059), .A2(new_n1062), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n1040), .A2(new_n1063), .ZN(new_n1064));
  AND3_X1   g639(.A1(new_n1029), .A2(new_n1031), .A3(new_n1032), .ZN(new_n1065));
  AOI21_X1  g640(.A(new_n1032), .B1(new_n1029), .B2(new_n1031), .ZN(new_n1066));
  OAI21_X1  g641(.A(new_n715), .B1(new_n1065), .B2(new_n1066), .ZN(new_n1067));
  INV_X1    g642(.A(new_n1039), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n1067), .A2(new_n1068), .ZN(new_n1069));
  AOI21_X1  g644(.A(new_n1016), .B1(new_n1069), .B2(G8), .ZN(new_n1070));
  NOR2_X1   g645(.A1(new_n1064), .A2(new_n1070), .ZN(new_n1071));
  INV_X1    g646(.A(KEYINPUT51), .ZN(new_n1072));
  NAND3_X1  g647(.A1(new_n1023), .A2(KEYINPUT120), .A3(KEYINPUT45), .ZN(new_n1073));
  INV_X1    g648(.A(KEYINPUT120), .ZN(new_n1074));
  OAI21_X1  g649(.A(new_n1074), .B1(new_n1030), .B2(new_n1017), .ZN(new_n1075));
  NAND3_X1  g650(.A1(new_n1031), .A2(new_n1073), .A3(new_n1075), .ZN(new_n1076));
  INV_X1    g651(.A(G1966), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n1076), .A2(new_n1077), .ZN(new_n1078));
  INV_X1    g653(.A(new_n1038), .ZN(new_n1079));
  INV_X1    g654(.A(G2084), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1079), .A2(new_n1080), .ZN(new_n1081));
  NAND2_X1  g656(.A1(new_n1078), .A2(new_n1081), .ZN(new_n1082));
  OAI211_X1 g657(.A(new_n1072), .B(G8), .C1(new_n1082), .C2(G286), .ZN(new_n1083));
  INV_X1    g658(.A(G8), .ZN(new_n1084));
  NOR2_X1   g659(.A1(G168), .A2(new_n1084), .ZN(new_n1085));
  INV_X1    g660(.A(new_n1085), .ZN(new_n1086));
  AOI22_X1  g661(.A1(new_n1076), .A2(new_n1077), .B1(new_n1079), .B2(new_n1080), .ZN(new_n1087));
  OAI211_X1 g662(.A(KEYINPUT51), .B(new_n1086), .C1(new_n1087), .C2(new_n1084), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n1082), .A2(new_n1085), .ZN(new_n1089));
  NAND3_X1  g664(.A1(new_n1083), .A2(new_n1088), .A3(new_n1089), .ZN(new_n1090));
  NAND2_X1  g665(.A1(new_n1090), .A2(KEYINPUT62), .ZN(new_n1091));
  INV_X1    g666(.A(G2078), .ZN(new_n1092));
  NAND3_X1  g667(.A1(new_n1025), .A2(new_n1092), .A3(new_n1033), .ZN(new_n1093));
  INV_X1    g668(.A(KEYINPUT53), .ZN(new_n1094));
  AOI22_X1  g669(.A1(new_n1093), .A2(new_n1094), .B1(new_n769), .B2(new_n1038), .ZN(new_n1095));
  OR3_X1    g670(.A1(new_n1076), .A2(new_n1094), .A3(G2078), .ZN(new_n1096));
  AOI21_X1  g671(.A(G301), .B1(new_n1095), .B2(new_n1096), .ZN(new_n1097));
  INV_X1    g672(.A(KEYINPUT62), .ZN(new_n1098));
  NAND4_X1  g673(.A1(new_n1083), .A2(new_n1098), .A3(new_n1088), .A4(new_n1089), .ZN(new_n1099));
  NAND4_X1  g674(.A1(new_n1071), .A2(new_n1091), .A3(new_n1097), .A4(new_n1099), .ZN(new_n1100));
  NOR3_X1   g675(.A1(new_n1040), .A2(new_n1062), .A3(new_n1059), .ZN(new_n1101));
  NOR2_X1   g676(.A1(G288), .A2(G1976), .ZN(new_n1102));
  XOR2_X1   g677(.A(new_n1102), .B(KEYINPUT119), .Z(new_n1103));
  OAI21_X1  g678(.A(new_n1103), .B1(new_n1044), .B2(new_n1045), .ZN(new_n1104));
  AOI22_X1  g679(.A1(new_n1104), .A2(new_n1042), .B1(new_n1050), .B2(new_n1056), .ZN(new_n1105));
  NOR2_X1   g680(.A1(new_n1101), .A2(new_n1105), .ZN(new_n1106));
  NOR3_X1   g681(.A1(new_n1087), .A2(new_n1084), .A3(G286), .ZN(new_n1107));
  AOI21_X1  g682(.A(KEYINPUT63), .B1(new_n1071), .B2(new_n1107), .ZN(new_n1108));
  INV_X1    g683(.A(KEYINPUT63), .ZN(new_n1109));
  INV_X1    g684(.A(new_n1107), .ZN(new_n1110));
  NOR4_X1   g685(.A1(new_n1064), .A2(new_n1070), .A3(new_n1109), .A4(new_n1110), .ZN(new_n1111));
  OAI211_X1 g686(.A(new_n1100), .B(new_n1106), .C1(new_n1108), .C2(new_n1111), .ZN(new_n1112));
  INV_X1    g687(.A(KEYINPUT123), .ZN(new_n1113));
  INV_X1    g688(.A(KEYINPUT59), .ZN(new_n1114));
  NAND3_X1  g689(.A1(new_n1029), .A2(new_n1031), .A3(new_n997), .ZN(new_n1115));
  XOR2_X1   g690(.A(KEYINPUT58), .B(G1341), .Z(new_n1116));
  NAND2_X1  g691(.A1(new_n1048), .A2(new_n1116), .ZN(new_n1117));
  NAND2_X1  g692(.A1(new_n1115), .A2(new_n1117), .ZN(new_n1118));
  INV_X1    g693(.A(KEYINPUT122), .ZN(new_n1119));
  NAND2_X1  g694(.A1(new_n1118), .A2(new_n1119), .ZN(new_n1120));
  NAND3_X1  g695(.A1(new_n1115), .A2(KEYINPUT122), .A3(new_n1117), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n1120), .A2(new_n1121), .ZN(new_n1122));
  AOI21_X1  g697(.A(new_n1114), .B1(new_n1122), .B2(new_n565), .ZN(new_n1123));
  AND3_X1   g698(.A1(new_n1115), .A2(KEYINPUT122), .A3(new_n1117), .ZN(new_n1124));
  AOI21_X1  g699(.A(KEYINPUT122), .B1(new_n1115), .B2(new_n1117), .ZN(new_n1125));
  OAI211_X1 g700(.A(new_n1114), .B(new_n565), .C1(new_n1124), .C2(new_n1125), .ZN(new_n1126));
  INV_X1    g701(.A(new_n1126), .ZN(new_n1127));
  NOR2_X1   g702(.A1(new_n1123), .A2(new_n1127), .ZN(new_n1128));
  XNOR2_X1  g703(.A(KEYINPUT56), .B(G2072), .ZN(new_n1129));
  NAND3_X1  g704(.A1(new_n1029), .A2(new_n1031), .A3(new_n1129), .ZN(new_n1130));
  NAND2_X1  g705(.A1(new_n578), .A2(KEYINPUT57), .ZN(new_n1131));
  INV_X1    g706(.A(KEYINPUT57), .ZN(new_n1132));
  OAI21_X1  g707(.A(new_n1132), .B1(new_n574), .B2(new_n577), .ZN(new_n1133));
  NAND2_X1  g708(.A1(new_n1131), .A2(new_n1133), .ZN(new_n1134));
  INV_X1    g709(.A(G1956), .ZN(new_n1135));
  NAND2_X1  g710(.A1(new_n1038), .A2(new_n1135), .ZN(new_n1136));
  NAND3_X1  g711(.A1(new_n1130), .A2(new_n1134), .A3(new_n1136), .ZN(new_n1137));
  INV_X1    g712(.A(KEYINPUT121), .ZN(new_n1138));
  NAND2_X1  g713(.A1(new_n1137), .A2(new_n1138), .ZN(new_n1139));
  NAND2_X1  g714(.A1(new_n1130), .A2(new_n1136), .ZN(new_n1140));
  INV_X1    g715(.A(new_n1134), .ZN(new_n1141));
  NAND2_X1  g716(.A1(new_n1140), .A2(new_n1141), .ZN(new_n1142));
  NAND4_X1  g717(.A1(new_n1130), .A2(new_n1136), .A3(new_n1134), .A4(KEYINPUT121), .ZN(new_n1143));
  NAND3_X1  g718(.A1(new_n1139), .A2(new_n1142), .A3(new_n1143), .ZN(new_n1144));
  INV_X1    g719(.A(KEYINPUT61), .ZN(new_n1145));
  NAND2_X1  g720(.A1(new_n1144), .A2(new_n1145), .ZN(new_n1146));
  NAND3_X1  g721(.A1(new_n1142), .A2(KEYINPUT61), .A3(new_n1137), .ZN(new_n1147));
  NAND2_X1  g722(.A1(new_n1146), .A2(new_n1147), .ZN(new_n1148));
  OAI21_X1  g723(.A(new_n1113), .B1(new_n1128), .B2(new_n1148), .ZN(new_n1149));
  OAI21_X1  g724(.A(new_n565), .B1(new_n1124), .B2(new_n1125), .ZN(new_n1150));
  NAND2_X1  g725(.A1(new_n1150), .A2(KEYINPUT59), .ZN(new_n1151));
  NAND2_X1  g726(.A1(new_n1151), .A2(new_n1126), .ZN(new_n1152));
  NAND4_X1  g727(.A1(new_n1152), .A2(KEYINPUT123), .A3(new_n1147), .A4(new_n1146), .ZN(new_n1153));
  INV_X1    g728(.A(G1348), .ZN(new_n1154));
  NAND2_X1  g729(.A1(new_n1038), .A2(new_n1154), .ZN(new_n1155));
  NAND3_X1  g730(.A1(new_n1022), .A2(new_n1023), .A3(new_n822), .ZN(new_n1156));
  AND2_X1   g731(.A1(new_n1155), .A2(new_n1156), .ZN(new_n1157));
  NAND3_X1  g732(.A1(new_n1157), .A2(KEYINPUT124), .A3(KEYINPUT60), .ZN(new_n1158));
  INV_X1    g733(.A(KEYINPUT124), .ZN(new_n1159));
  NAND2_X1  g734(.A1(new_n1155), .A2(new_n1156), .ZN(new_n1160));
  INV_X1    g735(.A(KEYINPUT60), .ZN(new_n1161));
  OAI21_X1  g736(.A(new_n1159), .B1(new_n1160), .B2(new_n1161), .ZN(new_n1162));
  NAND2_X1  g737(.A1(new_n1158), .A2(new_n1162), .ZN(new_n1163));
  AOI21_X1  g738(.A(new_n622), .B1(new_n1160), .B2(new_n1161), .ZN(new_n1164));
  XNOR2_X1  g739(.A(new_n1163), .B(new_n1164), .ZN(new_n1165));
  NAND3_X1  g740(.A1(new_n1149), .A2(new_n1153), .A3(new_n1165), .ZN(new_n1166));
  OAI21_X1  g741(.A(new_n1142), .B1(new_n622), .B2(new_n1157), .ZN(new_n1167));
  NAND3_X1  g742(.A1(new_n1167), .A2(new_n1139), .A3(new_n1143), .ZN(new_n1168));
  NAND2_X1  g743(.A1(new_n1166), .A2(new_n1168), .ZN(new_n1169));
  INV_X1    g744(.A(KEYINPUT54), .ZN(new_n1170));
  NAND2_X1  g745(.A1(new_n1093), .A2(new_n1094), .ZN(new_n1171));
  INV_X1    g746(.A(KEYINPUT125), .ZN(new_n1172));
  NAND3_X1  g747(.A1(new_n988), .A2(new_n1172), .A3(new_n1022), .ZN(new_n1173));
  OAI21_X1  g748(.A(KEYINPUT125), .B1(new_n987), .B2(new_n989), .ZN(new_n1174));
  XOR2_X1   g749(.A(KEYINPUT126), .B(G2078), .Z(new_n1175));
  NOR3_X1   g750(.A1(new_n1018), .A2(new_n1094), .A3(new_n1175), .ZN(new_n1176));
  NAND3_X1  g751(.A1(new_n1173), .A2(new_n1174), .A3(new_n1176), .ZN(new_n1177));
  NAND2_X1  g752(.A1(new_n1038), .A2(new_n769), .ZN(new_n1178));
  NAND3_X1  g753(.A1(new_n1171), .A2(new_n1177), .A3(new_n1178), .ZN(new_n1179));
  NOR2_X1   g754(.A1(new_n1179), .A2(G171), .ZN(new_n1180));
  OAI21_X1  g755(.A(new_n1170), .B1(new_n1180), .B2(new_n1097), .ZN(new_n1181));
  NAND3_X1  g756(.A1(new_n1181), .A2(new_n1071), .A3(new_n1090), .ZN(new_n1182));
  AOI211_X1 g757(.A(KEYINPUT127), .B(G301), .C1(new_n1095), .C2(new_n1177), .ZN(new_n1183));
  NAND3_X1  g758(.A1(new_n1095), .A2(G301), .A3(new_n1096), .ZN(new_n1184));
  NAND2_X1  g759(.A1(new_n1184), .A2(KEYINPUT54), .ZN(new_n1185));
  INV_X1    g760(.A(KEYINPUT127), .ZN(new_n1186));
  AOI21_X1  g761(.A(new_n1186), .B1(new_n1179), .B2(G171), .ZN(new_n1187));
  NOR3_X1   g762(.A1(new_n1183), .A2(new_n1185), .A3(new_n1187), .ZN(new_n1188));
  NOR2_X1   g763(.A1(new_n1182), .A2(new_n1188), .ZN(new_n1189));
  AOI21_X1  g764(.A(new_n1112), .B1(new_n1169), .B2(new_n1189), .ZN(new_n1190));
  NAND2_X1  g765(.A1(new_n993), .A2(KEYINPUT115), .ZN(new_n1191));
  NAND2_X1  g766(.A1(G290), .A2(G1986), .ZN(new_n1192));
  XOR2_X1   g767(.A(new_n1191), .B(new_n1192), .Z(new_n1193));
  OAI21_X1  g768(.A(new_n1001), .B1(new_n1193), .B2(new_n991), .ZN(new_n1194));
  OAI21_X1  g769(.A(new_n1013), .B1(new_n1190), .B2(new_n1194), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g770(.A(G319), .ZN(new_n1197));
  NOR4_X1   g771(.A1(G401), .A2(new_n1197), .A3(G227), .A4(G229), .ZN(new_n1198));
  AND3_X1   g772(.A1(new_n970), .A2(new_n1198), .A3(new_n885), .ZN(G308));
  NAND3_X1  g773(.A1(new_n970), .A2(new_n1198), .A3(new_n885), .ZN(G225));
endmodule


