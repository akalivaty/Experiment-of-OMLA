

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n522, n523, n524, n525,
         n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536,
         n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547,
         n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558,
         n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569,
         n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580,
         n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591,
         n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602,
         n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613,
         n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624,
         n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635,
         n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646,
         n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657,
         n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668,
         n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679,
         n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690,
         n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701,
         n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712,
         n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723,
         n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734,
         n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745,
         n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756,
         n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n767,
         n768, n769, n770, n771, n772, n773, n774, n775, n776, n777, n778,
         n779, n780, n781, n782, n783, n784, n785, n786, n787, n788, n789,
         n790, n791, n792, n793, n794, n795, n796, n797, n798, n799, n800,
         n801, n802, n803, n804, n805, n806, n807, n808, n809, n810, n811,
         n812, n813, n814, n815, n816, n817, n818, n819, n820, n821, n822,
         n823, n824, n825, n826, n827, n828, n829, n830, n831, n832, n833,
         n834, n835, n836, n837, n838, n839, n840, n841, n842, n843, n844,
         n845, n846, n847, n848, n849, n850, n851, n852, n853, n854, n855,
         n856, n857, n858, n859, n860, n861, n862, n863, n864, n865, n866,
         n867, n868, n869, n870, n871, n872, n873, n874, n875, n876, n877,
         n878, n879, n880, n881, n882, n883, n884, n885, n886, n887, n888,
         n889, n890, n891, n892, n893, n894, n895, n896, n897, n898, n899,
         n900, n901, n902, n903, n904, n905, n906, n907, n908, n909, n910,
         n911, n912, n913, n914, n915, n916, n917, n918, n919, n920, n921,
         n922, n923, n924, n925, n926, n927, n928, n929, n930, n931, n932,
         n933, n934, n935, n936, n937, n938, n939, n940, n941, n942, n943,
         n944, n945, n946, n947, n948, n949, n950, n951, n952, n953, n954,
         n955, n956, n957, n958, n959, n960, n961, n962, n963, n964, n965,
         n966, n967, n968, n969, n970, n971, n972, n973, n974, n975, n976,
         n977, n978, n979, n980, n981, n982, n983, n984, n985, n986, n987,
         n988, n989, n990, n991, n992, n993, n994, n995, n996, n997, n998,
         n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008,
         n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018,
         n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028,
         n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038,
         n1039, n1040, n1041;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  OR2_X1 U556 ( .A1(n687), .A2(n686), .ZN(n688) );
  INV_X1 U557 ( .A(KEYINPUT29), .ZN(n653) );
  NOR2_X1 U558 ( .A1(n737), .A2(n736), .ZN(n739) );
  INV_X1 U559 ( .A(KEYINPUT94), .ZN(n696) );
  NOR2_X1 U560 ( .A1(G2105), .A2(G2104), .ZN(n526) );
  AND2_X1 U561 ( .A1(n731), .A2(n762), .ZN(n522) );
  NAND2_X1 U562 ( .A1(n700), .A2(n743), .ZN(n523) );
  NOR2_X1 U563 ( .A1(n997), .A2(n628), .ZN(n643) );
  INV_X1 U564 ( .A(KEYINPUT92), .ZN(n646) );
  BUF_X1 U565 ( .A(n660), .Z(n668) );
  NOR2_X1 U566 ( .A1(n666), .A2(n665), .ZN(n667) );
  NOR2_X1 U567 ( .A1(G1966), .A2(n737), .ZN(n684) );
  NAND2_X1 U568 ( .A1(n719), .A2(n601), .ZN(n660) );
  INV_X1 U569 ( .A(KEYINPUT64), .ZN(n738) );
  INV_X1 U570 ( .A(KEYINPUT33), .ZN(n740) );
  NOR2_X1 U571 ( .A1(G164), .A2(G1384), .ZN(n719) );
  INV_X1 U572 ( .A(KEYINPUT17), .ZN(n525) );
  NAND2_X1 U573 ( .A1(n908), .A2(G138), .ZN(n527) );
  NAND2_X1 U574 ( .A1(G2104), .A2(G2105), .ZN(n524) );
  XNOR2_X2 U575 ( .A(n524), .B(KEYINPUT67), .ZN(n903) );
  NAND2_X1 U576 ( .A1(G114), .A2(n903), .ZN(n528) );
  XNOR2_X2 U577 ( .A(n526), .B(n525), .ZN(n908) );
  NAND2_X1 U578 ( .A1(n528), .A2(n527), .ZN(n534) );
  XNOR2_X1 U579 ( .A(G2104), .B(KEYINPUT65), .ZN(n530) );
  NOR2_X1 U580 ( .A1(G2105), .A2(n530), .ZN(n592) );
  INV_X1 U581 ( .A(n592), .ZN(n529) );
  INV_X2 U582 ( .A(n529), .ZN(n907) );
  NAND2_X1 U583 ( .A1(G102), .A2(n907), .ZN(n532) );
  AND2_X1 U584 ( .A1(n530), .A2(G2105), .ZN(n904) );
  NAND2_X1 U585 ( .A1(G126), .A2(n904), .ZN(n531) );
  NAND2_X1 U586 ( .A1(n532), .A2(n531), .ZN(n533) );
  OR2_X1 U587 ( .A1(n534), .A2(n533), .ZN(n535) );
  XNOR2_X2 U588 ( .A(n535), .B(KEYINPUT83), .ZN(G164) );
  INV_X1 U589 ( .A(G651), .ZN(n543) );
  NOR2_X1 U590 ( .A1(G543), .A2(n543), .ZN(n536) );
  XOR2_X2 U591 ( .A(KEYINPUT1), .B(n536), .Z(n795) );
  NAND2_X1 U592 ( .A1(G65), .A2(n795), .ZN(n538) );
  XOR2_X1 U593 ( .A(G543), .B(KEYINPUT0), .Z(n582) );
  NOR2_X1 U594 ( .A1(G651), .A2(n582), .ZN(n797) );
  NAND2_X1 U595 ( .A1(G53), .A2(n797), .ZN(n537) );
  NAND2_X1 U596 ( .A1(n538), .A2(n537), .ZN(n539) );
  XNOR2_X1 U597 ( .A(KEYINPUT72), .B(n539), .ZN(n542) );
  NOR2_X1 U598 ( .A1(G651), .A2(G543), .ZN(n801) );
  NAND2_X1 U599 ( .A1(G91), .A2(n801), .ZN(n540) );
  XNOR2_X1 U600 ( .A(KEYINPUT71), .B(n540), .ZN(n541) );
  NOR2_X1 U601 ( .A1(n542), .A2(n541), .ZN(n546) );
  OR2_X1 U602 ( .A1(n543), .A2(n582), .ZN(n544) );
  XOR2_X1 U603 ( .A(KEYINPUT68), .B(n544), .Z(n608) );
  BUF_X1 U604 ( .A(n608), .Z(n802) );
  NAND2_X1 U605 ( .A1(G78), .A2(n802), .ZN(n545) );
  NAND2_X1 U606 ( .A1(n546), .A2(n545), .ZN(G299) );
  NAND2_X1 U607 ( .A1(G64), .A2(n795), .ZN(n548) );
  NAND2_X1 U608 ( .A1(G52), .A2(n797), .ZN(n547) );
  NAND2_X1 U609 ( .A1(n548), .A2(n547), .ZN(n554) );
  NAND2_X1 U610 ( .A1(G90), .A2(n801), .ZN(n550) );
  NAND2_X1 U611 ( .A1(G77), .A2(n802), .ZN(n549) );
  NAND2_X1 U612 ( .A1(n550), .A2(n549), .ZN(n551) );
  XOR2_X1 U613 ( .A(KEYINPUT70), .B(n551), .Z(n552) );
  XNOR2_X1 U614 ( .A(KEYINPUT9), .B(n552), .ZN(n553) );
  NOR2_X1 U615 ( .A1(n554), .A2(n553), .ZN(G171) );
  NAND2_X1 U616 ( .A1(n801), .A2(G89), .ZN(n555) );
  XNOR2_X1 U617 ( .A(n555), .B(KEYINPUT4), .ZN(n557) );
  NAND2_X1 U618 ( .A1(G76), .A2(n802), .ZN(n556) );
  NAND2_X1 U619 ( .A1(n557), .A2(n556), .ZN(n558) );
  XNOR2_X1 U620 ( .A(n558), .B(KEYINPUT5), .ZN(n563) );
  NAND2_X1 U621 ( .A1(G63), .A2(n795), .ZN(n560) );
  NAND2_X1 U622 ( .A1(G51), .A2(n797), .ZN(n559) );
  NAND2_X1 U623 ( .A1(n560), .A2(n559), .ZN(n561) );
  XOR2_X1 U624 ( .A(KEYINPUT6), .B(n561), .Z(n562) );
  NAND2_X1 U625 ( .A1(n563), .A2(n562), .ZN(n564) );
  XNOR2_X1 U626 ( .A(n564), .B(KEYINPUT7), .ZN(G168) );
  NAND2_X1 U627 ( .A1(n802), .A2(G75), .ZN(n565) );
  XNOR2_X1 U628 ( .A(n565), .B(KEYINPUT80), .ZN(n567) );
  NAND2_X1 U629 ( .A1(n801), .A2(G88), .ZN(n566) );
  NAND2_X1 U630 ( .A1(n567), .A2(n566), .ZN(n571) );
  NAND2_X1 U631 ( .A1(G62), .A2(n795), .ZN(n569) );
  NAND2_X1 U632 ( .A1(G50), .A2(n797), .ZN(n568) );
  NAND2_X1 U633 ( .A1(n569), .A2(n568), .ZN(n570) );
  NOR2_X1 U634 ( .A1(n571), .A2(n570), .ZN(G166) );
  INV_X1 U635 ( .A(G166), .ZN(G303) );
  XOR2_X1 U636 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U637 ( .A1(G86), .A2(n801), .ZN(n573) );
  NAND2_X1 U638 ( .A1(G48), .A2(n797), .ZN(n572) );
  NAND2_X1 U639 ( .A1(n573), .A2(n572), .ZN(n576) );
  NAND2_X1 U640 ( .A1(n802), .A2(G73), .ZN(n574) );
  XOR2_X1 U641 ( .A(KEYINPUT2), .B(n574), .Z(n575) );
  NOR2_X1 U642 ( .A1(n576), .A2(n575), .ZN(n578) );
  NAND2_X1 U643 ( .A1(n795), .A2(G61), .ZN(n577) );
  NAND2_X1 U644 ( .A1(n578), .A2(n577), .ZN(G305) );
  NAND2_X1 U645 ( .A1(G49), .A2(n797), .ZN(n580) );
  NAND2_X1 U646 ( .A1(G74), .A2(G651), .ZN(n579) );
  NAND2_X1 U647 ( .A1(n580), .A2(n579), .ZN(n581) );
  NOR2_X1 U648 ( .A1(n795), .A2(n581), .ZN(n584) );
  NAND2_X1 U649 ( .A1(n582), .A2(G87), .ZN(n583) );
  NAND2_X1 U650 ( .A1(n584), .A2(n583), .ZN(G288) );
  NAND2_X1 U651 ( .A1(G85), .A2(n801), .ZN(n586) );
  NAND2_X1 U652 ( .A1(G47), .A2(n797), .ZN(n585) );
  NAND2_X1 U653 ( .A1(n586), .A2(n585), .ZN(n589) );
  NAND2_X1 U654 ( .A1(G60), .A2(n795), .ZN(n587) );
  XNOR2_X1 U655 ( .A(KEYINPUT69), .B(n587), .ZN(n588) );
  NOR2_X1 U656 ( .A1(n589), .A2(n588), .ZN(n591) );
  NAND2_X1 U657 ( .A1(G72), .A2(n802), .ZN(n590) );
  NAND2_X1 U658 ( .A1(n591), .A2(n590), .ZN(G290) );
  NAND2_X1 U659 ( .A1(n592), .A2(G101), .ZN(n593) );
  XOR2_X1 U660 ( .A(n593), .B(KEYINPUT23), .Z(n595) );
  NAND2_X1 U661 ( .A1(n904), .A2(G125), .ZN(n594) );
  NAND2_X1 U662 ( .A1(n595), .A2(n594), .ZN(n596) );
  XNOR2_X1 U663 ( .A(n596), .B(KEYINPUT66), .ZN(n781) );
  NAND2_X1 U664 ( .A1(G113), .A2(n903), .ZN(n598) );
  NAND2_X1 U665 ( .A1(G137), .A2(n908), .ZN(n597) );
  NAND2_X1 U666 ( .A1(n598), .A2(n597), .ZN(n780) );
  INV_X1 U667 ( .A(G40), .ZN(n599) );
  OR2_X1 U668 ( .A1(n780), .A2(n599), .ZN(n600) );
  OR2_X1 U669 ( .A1(n781), .A2(n600), .ZN(n718) );
  INV_X1 U670 ( .A(n718), .ZN(n601) );
  INV_X1 U671 ( .A(n668), .ZN(n637) );
  NAND2_X1 U672 ( .A1(n637), .A2(G2072), .ZN(n602) );
  XNOR2_X1 U673 ( .A(n602), .B(KEYINPUT27), .ZN(n604) );
  INV_X1 U674 ( .A(G1956), .ZN(n1026) );
  NOR2_X1 U675 ( .A1(n1026), .A2(n637), .ZN(n603) );
  NOR2_X1 U676 ( .A1(n604), .A2(n603), .ZN(n648) );
  INV_X1 U677 ( .A(G299), .ZN(n1001) );
  NOR2_X1 U678 ( .A1(n648), .A2(n1001), .ZN(n606) );
  XNOR2_X1 U679 ( .A(KEYINPUT28), .B(KEYINPUT89), .ZN(n605) );
  XNOR2_X1 U680 ( .A(n606), .B(n605), .ZN(n652) );
  NAND2_X1 U681 ( .A1(n801), .A2(G81), .ZN(n607) );
  XNOR2_X1 U682 ( .A(KEYINPUT12), .B(n607), .ZN(n612) );
  NAND2_X1 U683 ( .A1(G68), .A2(n608), .ZN(n609) );
  XOR2_X1 U684 ( .A(n609), .B(KEYINPUT73), .Z(n613) );
  NAND2_X1 U685 ( .A1(n612), .A2(n613), .ZN(n610) );
  NAND2_X1 U686 ( .A1(n610), .A2(KEYINPUT13), .ZN(n616) );
  INV_X1 U687 ( .A(KEYINPUT13), .ZN(n611) );
  AND2_X1 U688 ( .A1(n612), .A2(n611), .ZN(n614) );
  NAND2_X1 U689 ( .A1(n614), .A2(n613), .ZN(n615) );
  NAND2_X1 U690 ( .A1(n616), .A2(n615), .ZN(n621) );
  AND2_X1 U691 ( .A1(G43), .A2(n797), .ZN(n619) );
  NAND2_X1 U692 ( .A1(n795), .A2(G56), .ZN(n617) );
  XOR2_X1 U693 ( .A(KEYINPUT14), .B(n617), .Z(n618) );
  NOR2_X1 U694 ( .A1(n619), .A2(n618), .ZN(n620) );
  AND2_X1 U695 ( .A1(n621), .A2(n620), .ZN(n622) );
  XOR2_X2 U696 ( .A(KEYINPUT74), .B(n622), .Z(n997) );
  INV_X1 U697 ( .A(n660), .ZN(n623) );
  NAND2_X1 U698 ( .A1(n623), .A2(G1996), .ZN(n624) );
  XNOR2_X1 U699 ( .A(n624), .B(KEYINPUT26), .ZN(n626) );
  NAND2_X1 U700 ( .A1(G1341), .A2(n668), .ZN(n625) );
  NAND2_X1 U701 ( .A1(n626), .A2(n625), .ZN(n627) );
  XNOR2_X1 U702 ( .A(n627), .B(KEYINPUT90), .ZN(n628) );
  NAND2_X1 U703 ( .A1(n802), .A2(G79), .ZN(n635) );
  NAND2_X1 U704 ( .A1(G66), .A2(n795), .ZN(n630) );
  NAND2_X1 U705 ( .A1(G92), .A2(n801), .ZN(n629) );
  NAND2_X1 U706 ( .A1(n630), .A2(n629), .ZN(n633) );
  NAND2_X1 U707 ( .A1(G54), .A2(n797), .ZN(n631) );
  XNOR2_X1 U708 ( .A(KEYINPUT75), .B(n631), .ZN(n632) );
  NOR2_X1 U709 ( .A1(n633), .A2(n632), .ZN(n634) );
  NAND2_X1 U710 ( .A1(n635), .A2(n634), .ZN(n636) );
  XNOR2_X1 U711 ( .A(n636), .B(KEYINPUT15), .ZN(n987) );
  NAND2_X1 U712 ( .A1(n643), .A2(n987), .ZN(n641) );
  NOR2_X1 U713 ( .A1(n637), .A2(G1348), .ZN(n639) );
  NOR2_X1 U714 ( .A1(G2067), .A2(n668), .ZN(n638) );
  NOR2_X1 U715 ( .A1(n639), .A2(n638), .ZN(n640) );
  NAND2_X1 U716 ( .A1(n641), .A2(n640), .ZN(n642) );
  XNOR2_X1 U717 ( .A(n642), .B(KEYINPUT91), .ZN(n645) );
  NOR2_X1 U718 ( .A1(n987), .A2(n643), .ZN(n644) );
  NOR2_X1 U719 ( .A1(n645), .A2(n644), .ZN(n647) );
  XNOR2_X1 U720 ( .A(n647), .B(n646), .ZN(n650) );
  NAND2_X1 U721 ( .A1(n648), .A2(n1001), .ZN(n649) );
  NAND2_X1 U722 ( .A1(n650), .A2(n649), .ZN(n651) );
  NAND2_X1 U723 ( .A1(n652), .A2(n651), .ZN(n654) );
  XNOR2_X1 U724 ( .A(n654), .B(n653), .ZN(n658) );
  XNOR2_X1 U725 ( .A(G2078), .B(KEYINPUT25), .ZN(n936) );
  NOR2_X1 U726 ( .A1(n668), .A2(n936), .ZN(n656) );
  AND2_X1 U727 ( .A1(n668), .A2(G1961), .ZN(n655) );
  NOR2_X1 U728 ( .A1(n656), .A2(n655), .ZN(n659) );
  NAND2_X1 U729 ( .A1(G171), .A2(n659), .ZN(n657) );
  NAND2_X1 U730 ( .A1(n658), .A2(n657), .ZN(n682) );
  NOR2_X1 U731 ( .A1(G171), .A2(n659), .ZN(n666) );
  NAND2_X1 U732 ( .A1(n660), .A2(G8), .ZN(n661) );
  XNOR2_X1 U733 ( .A(n661), .B(KEYINPUT87), .ZN(n743) );
  INV_X1 U734 ( .A(n743), .ZN(n737) );
  NOR2_X1 U735 ( .A1(G2084), .A2(n668), .ZN(n683) );
  NOR2_X1 U736 ( .A1(n684), .A2(n683), .ZN(n662) );
  NAND2_X1 U737 ( .A1(G8), .A2(n662), .ZN(n663) );
  XNOR2_X1 U738 ( .A(KEYINPUT30), .B(n663), .ZN(n664) );
  NOR2_X1 U739 ( .A1(G168), .A2(n664), .ZN(n665) );
  XOR2_X1 U740 ( .A(KEYINPUT31), .B(n667), .Z(n681) );
  INV_X1 U741 ( .A(G8), .ZN(n673) );
  NOR2_X1 U742 ( .A1(G1971), .A2(n737), .ZN(n670) );
  NOR2_X1 U743 ( .A1(G2090), .A2(n668), .ZN(n669) );
  NOR2_X1 U744 ( .A1(n670), .A2(n669), .ZN(n671) );
  NAND2_X1 U745 ( .A1(n671), .A2(G303), .ZN(n672) );
  OR2_X1 U746 ( .A1(n673), .A2(n672), .ZN(n675) );
  AND2_X1 U747 ( .A1(n681), .A2(n675), .ZN(n674) );
  NAND2_X1 U748 ( .A1(n682), .A2(n674), .ZN(n679) );
  INV_X1 U749 ( .A(n675), .ZN(n677) );
  AND2_X1 U750 ( .A1(G286), .A2(G8), .ZN(n676) );
  OR2_X1 U751 ( .A1(n677), .A2(n676), .ZN(n678) );
  NAND2_X1 U752 ( .A1(n679), .A2(n678), .ZN(n680) );
  XNOR2_X1 U753 ( .A(n680), .B(KEYINPUT32), .ZN(n689) );
  AND2_X1 U754 ( .A1(n682), .A2(n681), .ZN(n687) );
  AND2_X1 U755 ( .A1(G8), .A2(n683), .ZN(n685) );
  OR2_X1 U756 ( .A1(n685), .A2(n684), .ZN(n686) );
  NAND2_X1 U757 ( .A1(n689), .A2(n688), .ZN(n691) );
  INV_X1 U758 ( .A(KEYINPUT93), .ZN(n690) );
  XNOR2_X1 U759 ( .A(n691), .B(n690), .ZN(n734) );
  INV_X1 U760 ( .A(n734), .ZN(n694) );
  NAND2_X1 U761 ( .A1(G166), .A2(G8), .ZN(n692) );
  NOR2_X1 U762 ( .A1(G2090), .A2(n692), .ZN(n693) );
  NOR2_X1 U763 ( .A1(n694), .A2(n693), .ZN(n695) );
  NOR2_X1 U764 ( .A1(n695), .A2(n743), .ZN(n697) );
  XNOR2_X1 U765 ( .A(n697), .B(n696), .ZN(n701) );
  NOR2_X1 U766 ( .A1(G1981), .A2(G305), .ZN(n698) );
  XNOR2_X1 U767 ( .A(n698), .B(KEYINPUT88), .ZN(n699) );
  XNOR2_X1 U768 ( .A(n699), .B(KEYINPUT24), .ZN(n700) );
  NAND2_X1 U769 ( .A1(n701), .A2(n523), .ZN(n732) );
  NAND2_X1 U770 ( .A1(G95), .A2(n907), .ZN(n703) );
  NAND2_X1 U771 ( .A1(G131), .A2(n908), .ZN(n702) );
  NAND2_X1 U772 ( .A1(n703), .A2(n702), .ZN(n707) );
  NAND2_X1 U773 ( .A1(G107), .A2(n903), .ZN(n705) );
  NAND2_X1 U774 ( .A1(G119), .A2(n904), .ZN(n704) );
  NAND2_X1 U775 ( .A1(n705), .A2(n704), .ZN(n706) );
  OR2_X1 U776 ( .A1(n707), .A2(n706), .ZN(n887) );
  AND2_X1 U777 ( .A1(n887), .A2(G1991), .ZN(n717) );
  NAND2_X1 U778 ( .A1(n903), .A2(G117), .ZN(n714) );
  NAND2_X1 U779 ( .A1(G141), .A2(n908), .ZN(n709) );
  NAND2_X1 U780 ( .A1(G129), .A2(n904), .ZN(n708) );
  NAND2_X1 U781 ( .A1(n709), .A2(n708), .ZN(n712) );
  NAND2_X1 U782 ( .A1(n907), .A2(G105), .ZN(n710) );
  XOR2_X1 U783 ( .A(KEYINPUT38), .B(n710), .Z(n711) );
  NOR2_X1 U784 ( .A1(n712), .A2(n711), .ZN(n713) );
  NAND2_X1 U785 ( .A1(n714), .A2(n713), .ZN(n715) );
  XOR2_X1 U786 ( .A(KEYINPUT85), .B(n715), .Z(n893) );
  AND2_X1 U787 ( .A1(n893), .A2(G1996), .ZN(n716) );
  NOR2_X1 U788 ( .A1(n717), .A2(n716), .ZN(n960) );
  NOR2_X1 U789 ( .A1(n719), .A2(n718), .ZN(n766) );
  INV_X1 U790 ( .A(n766), .ZN(n720) );
  NOR2_X1 U791 ( .A1(n960), .A2(n720), .ZN(n756) );
  XOR2_X1 U792 ( .A(KEYINPUT86), .B(n756), .Z(n731) );
  NAND2_X1 U793 ( .A1(G104), .A2(n907), .ZN(n722) );
  NAND2_X1 U794 ( .A1(G140), .A2(n908), .ZN(n721) );
  NAND2_X1 U795 ( .A1(n722), .A2(n721), .ZN(n723) );
  XNOR2_X1 U796 ( .A(KEYINPUT34), .B(n723), .ZN(n728) );
  NAND2_X1 U797 ( .A1(G116), .A2(n903), .ZN(n725) );
  NAND2_X1 U798 ( .A1(G128), .A2(n904), .ZN(n724) );
  NAND2_X1 U799 ( .A1(n725), .A2(n724), .ZN(n726) );
  XOR2_X1 U800 ( .A(n726), .B(KEYINPUT35), .Z(n727) );
  NOR2_X1 U801 ( .A1(n728), .A2(n727), .ZN(n729) );
  XOR2_X1 U802 ( .A(KEYINPUT36), .B(n729), .Z(n730) );
  XOR2_X1 U803 ( .A(KEYINPUT84), .B(n730), .Z(n889) );
  XNOR2_X1 U804 ( .A(KEYINPUT37), .B(G2067), .ZN(n764) );
  NOR2_X1 U805 ( .A1(n889), .A2(n764), .ZN(n958) );
  NAND2_X1 U806 ( .A1(n766), .A2(n958), .ZN(n762) );
  NAND2_X1 U807 ( .A1(n732), .A2(n522), .ZN(n750) );
  NOR2_X1 U808 ( .A1(G1976), .A2(G288), .ZN(n742) );
  NOR2_X1 U809 ( .A1(G1971), .A2(G303), .ZN(n733) );
  NOR2_X1 U810 ( .A1(n742), .A2(n733), .ZN(n992) );
  NAND2_X1 U811 ( .A1(n992), .A2(n734), .ZN(n735) );
  NAND2_X1 U812 ( .A1(G1976), .A2(G288), .ZN(n991) );
  NAND2_X1 U813 ( .A1(n735), .A2(n991), .ZN(n736) );
  XNOR2_X1 U814 ( .A(n739), .B(n738), .ZN(n741) );
  NAND2_X1 U815 ( .A1(n741), .A2(n740), .ZN(n748) );
  XNOR2_X1 U816 ( .A(G1981), .B(G305), .ZN(n985) );
  AND2_X1 U817 ( .A1(n742), .A2(KEYINPUT33), .ZN(n744) );
  AND2_X1 U818 ( .A1(n744), .A2(n743), .ZN(n745) );
  NOR2_X1 U819 ( .A1(n985), .A2(n745), .ZN(n746) );
  AND2_X1 U820 ( .A1(n746), .A2(n522), .ZN(n747) );
  NAND2_X1 U821 ( .A1(n748), .A2(n747), .ZN(n749) );
  NAND2_X1 U822 ( .A1(n750), .A2(n749), .ZN(n752) );
  XNOR2_X1 U823 ( .A(G1986), .B(G290), .ZN(n1005) );
  NAND2_X1 U824 ( .A1(n1005), .A2(n766), .ZN(n751) );
  NAND2_X1 U825 ( .A1(n752), .A2(n751), .ZN(n769) );
  NOR2_X1 U826 ( .A1(G1996), .A2(n893), .ZN(n753) );
  XOR2_X1 U827 ( .A(KEYINPUT95), .B(n753), .Z(n962) );
  NOR2_X1 U828 ( .A1(G1991), .A2(n887), .ZN(n955) );
  NOR2_X1 U829 ( .A1(G1986), .A2(G290), .ZN(n754) );
  NOR2_X1 U830 ( .A1(n955), .A2(n754), .ZN(n755) );
  NOR2_X1 U831 ( .A1(n756), .A2(n755), .ZN(n757) );
  XNOR2_X1 U832 ( .A(n757), .B(KEYINPUT96), .ZN(n758) );
  NOR2_X1 U833 ( .A1(n962), .A2(n758), .ZN(n761) );
  XOR2_X1 U834 ( .A(KEYINPUT97), .B(KEYINPUT98), .Z(n759) );
  XNOR2_X1 U835 ( .A(KEYINPUT39), .B(n759), .ZN(n760) );
  XNOR2_X1 U836 ( .A(n761), .B(n760), .ZN(n763) );
  NAND2_X1 U837 ( .A1(n763), .A2(n762), .ZN(n765) );
  NAND2_X1 U838 ( .A1(n889), .A2(n764), .ZN(n967) );
  NAND2_X1 U839 ( .A1(n765), .A2(n967), .ZN(n767) );
  NAND2_X1 U840 ( .A1(n767), .A2(n766), .ZN(n768) );
  NAND2_X1 U841 ( .A1(n769), .A2(n768), .ZN(n770) );
  XNOR2_X1 U842 ( .A(n770), .B(KEYINPUT40), .ZN(G329) );
  AND2_X1 U843 ( .A1(G452), .A2(G94), .ZN(G173) );
  NAND2_X1 U844 ( .A1(G123), .A2(n904), .ZN(n771) );
  XNOR2_X1 U845 ( .A(n771), .B(KEYINPUT18), .ZN(n778) );
  NAND2_X1 U846 ( .A1(G99), .A2(n907), .ZN(n773) );
  NAND2_X1 U847 ( .A1(G135), .A2(n908), .ZN(n772) );
  NAND2_X1 U848 ( .A1(n773), .A2(n772), .ZN(n776) );
  NAND2_X1 U849 ( .A1(n903), .A2(G111), .ZN(n774) );
  XOR2_X1 U850 ( .A(KEYINPUT76), .B(n774), .Z(n775) );
  NOR2_X1 U851 ( .A1(n776), .A2(n775), .ZN(n777) );
  NAND2_X1 U852 ( .A1(n778), .A2(n777), .ZN(n952) );
  XNOR2_X1 U853 ( .A(G2096), .B(n952), .ZN(n779) );
  OR2_X1 U854 ( .A1(G2100), .A2(n779), .ZN(G156) );
  INV_X1 U855 ( .A(G860), .ZN(n789) );
  OR2_X1 U856 ( .A1(n789), .A2(n997), .ZN(G153) );
  INV_X1 U857 ( .A(G57), .ZN(G237) );
  INV_X1 U858 ( .A(G132), .ZN(G219) );
  INV_X1 U859 ( .A(G82), .ZN(G220) );
  NOR2_X1 U860 ( .A1(n781), .A2(n780), .ZN(G160) );
  NAND2_X1 U861 ( .A1(G7), .A2(G661), .ZN(n782) );
  XNOR2_X1 U862 ( .A(n782), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U863 ( .A(G223), .ZN(n834) );
  NAND2_X1 U864 ( .A1(n834), .A2(G567), .ZN(n783) );
  XOR2_X1 U865 ( .A(KEYINPUT11), .B(n783), .Z(G234) );
  INV_X1 U866 ( .A(G171), .ZN(G301) );
  NAND2_X1 U867 ( .A1(G868), .A2(G301), .ZN(n785) );
  OR2_X1 U868 ( .A1(n987), .A2(G868), .ZN(n784) );
  NAND2_X1 U869 ( .A1(n785), .A2(n784), .ZN(G284) );
  INV_X1 U870 ( .A(G868), .ZN(n786) );
  NOR2_X1 U871 ( .A1(G286), .A2(n786), .ZN(n788) );
  NOR2_X1 U872 ( .A1(G868), .A2(G299), .ZN(n787) );
  NOR2_X1 U873 ( .A1(n788), .A2(n787), .ZN(G297) );
  NAND2_X1 U874 ( .A1(n789), .A2(G559), .ZN(n790) );
  NAND2_X1 U875 ( .A1(n790), .A2(n987), .ZN(n791) );
  XNOR2_X1 U876 ( .A(n791), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U877 ( .A1(n997), .A2(G868), .ZN(n794) );
  NAND2_X1 U878 ( .A1(n987), .A2(G868), .ZN(n792) );
  NOR2_X1 U879 ( .A1(G559), .A2(n792), .ZN(n793) );
  NOR2_X1 U880 ( .A1(n794), .A2(n793), .ZN(G282) );
  NAND2_X1 U881 ( .A1(n795), .A2(G67), .ZN(n796) );
  XOR2_X1 U882 ( .A(KEYINPUT77), .B(n796), .Z(n799) );
  NAND2_X1 U883 ( .A1(n797), .A2(G55), .ZN(n798) );
  NAND2_X1 U884 ( .A1(n799), .A2(n798), .ZN(n800) );
  XNOR2_X1 U885 ( .A(KEYINPUT78), .B(n800), .ZN(n806) );
  NAND2_X1 U886 ( .A1(G93), .A2(n801), .ZN(n804) );
  NAND2_X1 U887 ( .A1(G80), .A2(n802), .ZN(n803) );
  NAND2_X1 U888 ( .A1(n804), .A2(n803), .ZN(n805) );
  NOR2_X1 U889 ( .A1(n806), .A2(n805), .ZN(n812) );
  NAND2_X1 U890 ( .A1(G559), .A2(n987), .ZN(n807) );
  XNOR2_X1 U891 ( .A(n807), .B(n997), .ZN(n817) );
  NOR2_X1 U892 ( .A1(n817), .A2(G860), .ZN(n808) );
  XOR2_X1 U893 ( .A(KEYINPUT79), .B(n808), .Z(n809) );
  XNOR2_X1 U894 ( .A(n812), .B(n809), .ZN(G145) );
  NOR2_X1 U895 ( .A1(G868), .A2(n812), .ZN(n810) );
  XOR2_X1 U896 ( .A(n810), .B(KEYINPUT82), .Z(n821) );
  XNOR2_X1 U897 ( .A(KEYINPUT19), .B(G290), .ZN(n811) );
  XNOR2_X1 U898 ( .A(n811), .B(G288), .ZN(n813) );
  XOR2_X1 U899 ( .A(n813), .B(n812), .Z(n815) );
  XNOR2_X1 U900 ( .A(G166), .B(n1001), .ZN(n814) );
  XNOR2_X1 U901 ( .A(n815), .B(n814), .ZN(n816) );
  XNOR2_X1 U902 ( .A(n816), .B(G305), .ZN(n918) );
  XNOR2_X1 U903 ( .A(n918), .B(n817), .ZN(n818) );
  XNOR2_X1 U904 ( .A(n818), .B(KEYINPUT81), .ZN(n819) );
  NAND2_X1 U905 ( .A1(G868), .A2(n819), .ZN(n820) );
  NAND2_X1 U906 ( .A1(n821), .A2(n820), .ZN(G295) );
  NAND2_X1 U907 ( .A1(G2078), .A2(G2084), .ZN(n822) );
  XOR2_X1 U908 ( .A(KEYINPUT20), .B(n822), .Z(n823) );
  NAND2_X1 U909 ( .A1(G2090), .A2(n823), .ZN(n824) );
  XNOR2_X1 U910 ( .A(KEYINPUT21), .B(n824), .ZN(n825) );
  NAND2_X1 U911 ( .A1(n825), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U912 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U913 ( .A1(G220), .A2(G219), .ZN(n826) );
  XOR2_X1 U914 ( .A(KEYINPUT22), .B(n826), .Z(n827) );
  NOR2_X1 U915 ( .A1(G218), .A2(n827), .ZN(n828) );
  NAND2_X1 U916 ( .A1(G96), .A2(n828), .ZN(n840) );
  NAND2_X1 U917 ( .A1(n840), .A2(G2106), .ZN(n832) );
  NAND2_X1 U918 ( .A1(G120), .A2(G108), .ZN(n829) );
  NOR2_X1 U919 ( .A1(G237), .A2(n829), .ZN(n830) );
  NAND2_X1 U920 ( .A1(G69), .A2(n830), .ZN(n841) );
  NAND2_X1 U921 ( .A1(n841), .A2(G567), .ZN(n831) );
  NAND2_X1 U922 ( .A1(n832), .A2(n831), .ZN(n855) );
  NAND2_X1 U923 ( .A1(G483), .A2(G661), .ZN(n833) );
  NOR2_X1 U924 ( .A1(n855), .A2(n833), .ZN(n838) );
  NAND2_X1 U925 ( .A1(n838), .A2(G36), .ZN(G176) );
  NAND2_X1 U926 ( .A1(G2106), .A2(n834), .ZN(G217) );
  NAND2_X1 U927 ( .A1(G15), .A2(G2), .ZN(n835) );
  XNOR2_X1 U928 ( .A(KEYINPUT103), .B(n835), .ZN(n836) );
  NAND2_X1 U929 ( .A1(n836), .A2(G661), .ZN(G259) );
  NAND2_X1 U930 ( .A1(G3), .A2(G1), .ZN(n837) );
  XNOR2_X1 U931 ( .A(KEYINPUT104), .B(n837), .ZN(n839) );
  NAND2_X1 U932 ( .A1(n839), .A2(n838), .ZN(G188) );
  XOR2_X1 U933 ( .A(G108), .B(KEYINPUT112), .Z(G238) );
  INV_X1 U935 ( .A(G120), .ZN(G236) );
  INV_X1 U936 ( .A(G96), .ZN(G221) );
  NOR2_X1 U937 ( .A1(n841), .A2(n840), .ZN(G325) );
  INV_X1 U938 ( .A(G325), .ZN(G261) );
  XOR2_X1 U939 ( .A(KEYINPUT100), .B(G2443), .Z(n843) );
  XNOR2_X1 U940 ( .A(G2451), .B(G2427), .ZN(n842) );
  XNOR2_X1 U941 ( .A(n843), .B(n842), .ZN(n844) );
  XOR2_X1 U942 ( .A(n844), .B(G2430), .Z(n846) );
  XNOR2_X1 U943 ( .A(G1341), .B(G1348), .ZN(n845) );
  XNOR2_X1 U944 ( .A(n846), .B(n845), .ZN(n850) );
  XOR2_X1 U945 ( .A(KEYINPUT101), .B(G2435), .Z(n848) );
  XNOR2_X1 U946 ( .A(G2438), .B(G2454), .ZN(n847) );
  XNOR2_X1 U947 ( .A(n848), .B(n847), .ZN(n849) );
  XOR2_X1 U948 ( .A(n850), .B(n849), .Z(n852) );
  XNOR2_X1 U949 ( .A(G2446), .B(KEYINPUT99), .ZN(n851) );
  XNOR2_X1 U950 ( .A(n852), .B(n851), .ZN(n853) );
  NAND2_X1 U951 ( .A1(G14), .A2(n853), .ZN(n854) );
  XOR2_X1 U952 ( .A(KEYINPUT102), .B(n854), .Z(G401) );
  INV_X1 U953 ( .A(n855), .ZN(G319) );
  XOR2_X1 U954 ( .A(G1961), .B(G1971), .Z(n857) );
  XNOR2_X1 U955 ( .A(G1986), .B(G1976), .ZN(n856) );
  XNOR2_X1 U956 ( .A(n857), .B(n856), .ZN(n858) );
  XOR2_X1 U957 ( .A(n858), .B(KEYINPUT41), .Z(n860) );
  XNOR2_X1 U958 ( .A(G1996), .B(G1991), .ZN(n859) );
  XNOR2_X1 U959 ( .A(n860), .B(n859), .ZN(n864) );
  XOR2_X1 U960 ( .A(G2474), .B(G1956), .Z(n862) );
  XNOR2_X1 U961 ( .A(G1981), .B(G1966), .ZN(n861) );
  XNOR2_X1 U962 ( .A(n862), .B(n861), .ZN(n863) );
  XNOR2_X1 U963 ( .A(n864), .B(n863), .ZN(G229) );
  XOR2_X1 U964 ( .A(G2096), .B(G2090), .Z(n866) );
  XNOR2_X1 U965 ( .A(G2067), .B(G2072), .ZN(n865) );
  XNOR2_X1 U966 ( .A(n866), .B(n865), .ZN(n876) );
  XOR2_X1 U967 ( .A(KEYINPUT42), .B(KEYINPUT107), .Z(n868) );
  XNOR2_X1 U968 ( .A(G2678), .B(KEYINPUT108), .ZN(n867) );
  XNOR2_X1 U969 ( .A(n868), .B(n867), .ZN(n872) );
  XOR2_X1 U970 ( .A(G2100), .B(KEYINPUT43), .Z(n870) );
  XNOR2_X1 U971 ( .A(KEYINPUT105), .B(KEYINPUT106), .ZN(n869) );
  XNOR2_X1 U972 ( .A(n870), .B(n869), .ZN(n871) );
  XOR2_X1 U973 ( .A(n872), .B(n871), .Z(n874) );
  XNOR2_X1 U974 ( .A(G2078), .B(G2084), .ZN(n873) );
  XNOR2_X1 U975 ( .A(n874), .B(n873), .ZN(n875) );
  XOR2_X1 U976 ( .A(n876), .B(n875), .Z(G227) );
  NAND2_X1 U977 ( .A1(G124), .A2(n904), .ZN(n877) );
  XOR2_X1 U978 ( .A(KEYINPUT44), .B(n877), .Z(n878) );
  XNOR2_X1 U979 ( .A(n878), .B(KEYINPUT109), .ZN(n880) );
  NAND2_X1 U980 ( .A1(G112), .A2(n903), .ZN(n879) );
  NAND2_X1 U981 ( .A1(n880), .A2(n879), .ZN(n884) );
  NAND2_X1 U982 ( .A1(G100), .A2(n907), .ZN(n882) );
  NAND2_X1 U983 ( .A1(G136), .A2(n908), .ZN(n881) );
  NAND2_X1 U984 ( .A1(n882), .A2(n881), .ZN(n883) );
  NOR2_X1 U985 ( .A1(n884), .A2(n883), .ZN(G162) );
  XNOR2_X1 U986 ( .A(KEYINPUT110), .B(KEYINPUT48), .ZN(n886) );
  XNOR2_X1 U987 ( .A(n952), .B(KEYINPUT46), .ZN(n885) );
  XNOR2_X1 U988 ( .A(n886), .B(n885), .ZN(n888) );
  XNOR2_X1 U989 ( .A(n888), .B(n887), .ZN(n891) );
  XNOR2_X1 U990 ( .A(G160), .B(n889), .ZN(n890) );
  XNOR2_X1 U991 ( .A(n891), .B(n890), .ZN(n892) );
  XOR2_X1 U992 ( .A(n892), .B(G162), .Z(n895) );
  XOR2_X1 U993 ( .A(G164), .B(n893), .Z(n894) );
  XNOR2_X1 U994 ( .A(n895), .B(n894), .ZN(n916) );
  NAND2_X1 U995 ( .A1(G103), .A2(n907), .ZN(n897) );
  NAND2_X1 U996 ( .A1(G139), .A2(n908), .ZN(n896) );
  NAND2_X1 U997 ( .A1(n897), .A2(n896), .ZN(n902) );
  NAND2_X1 U998 ( .A1(G115), .A2(n903), .ZN(n899) );
  NAND2_X1 U999 ( .A1(G127), .A2(n904), .ZN(n898) );
  NAND2_X1 U1000 ( .A1(n899), .A2(n898), .ZN(n900) );
  XOR2_X1 U1001 ( .A(KEYINPUT47), .B(n900), .Z(n901) );
  NOR2_X1 U1002 ( .A1(n902), .A2(n901), .ZN(n970) );
  NAND2_X1 U1003 ( .A1(G118), .A2(n903), .ZN(n906) );
  NAND2_X1 U1004 ( .A1(G130), .A2(n904), .ZN(n905) );
  NAND2_X1 U1005 ( .A1(n906), .A2(n905), .ZN(n913) );
  NAND2_X1 U1006 ( .A1(G106), .A2(n907), .ZN(n910) );
  NAND2_X1 U1007 ( .A1(G142), .A2(n908), .ZN(n909) );
  NAND2_X1 U1008 ( .A1(n910), .A2(n909), .ZN(n911) );
  XOR2_X1 U1009 ( .A(KEYINPUT45), .B(n911), .Z(n912) );
  NOR2_X1 U1010 ( .A1(n913), .A2(n912), .ZN(n914) );
  XOR2_X1 U1011 ( .A(n970), .B(n914), .Z(n915) );
  XNOR2_X1 U1012 ( .A(n916), .B(n915), .ZN(n917) );
  NOR2_X1 U1013 ( .A1(G37), .A2(n917), .ZN(G395) );
  XOR2_X1 U1014 ( .A(n918), .B(G286), .Z(n920) );
  XNOR2_X1 U1015 ( .A(G171), .B(n987), .ZN(n919) );
  XNOR2_X1 U1016 ( .A(n920), .B(n919), .ZN(n921) );
  XOR2_X1 U1017 ( .A(n997), .B(n921), .Z(n922) );
  NOR2_X1 U1018 ( .A1(G37), .A2(n922), .ZN(G397) );
  NOR2_X1 U1019 ( .A1(G229), .A2(G227), .ZN(n923) );
  XOR2_X1 U1020 ( .A(KEYINPUT49), .B(n923), .Z(n924) );
  NAND2_X1 U1021 ( .A1(G319), .A2(n924), .ZN(n925) );
  NOR2_X1 U1022 ( .A1(G401), .A2(n925), .ZN(n928) );
  NOR2_X1 U1023 ( .A1(G395), .A2(G397), .ZN(n926) );
  XOR2_X1 U1024 ( .A(KEYINPUT111), .B(n926), .Z(n927) );
  NAND2_X1 U1025 ( .A1(n928), .A2(n927), .ZN(G225) );
  INV_X1 U1026 ( .A(G225), .ZN(G308) );
  INV_X1 U1027 ( .A(G69), .ZN(G235) );
  XOR2_X1 U1028 ( .A(G2090), .B(G35), .Z(n932) );
  XNOR2_X1 U1029 ( .A(KEYINPUT54), .B(G34), .ZN(n929) );
  XNOR2_X1 U1030 ( .A(n929), .B(KEYINPUT119), .ZN(n930) );
  XNOR2_X1 U1031 ( .A(n930), .B(G2084), .ZN(n931) );
  NAND2_X1 U1032 ( .A1(n932), .A2(n931), .ZN(n947) );
  XNOR2_X1 U1033 ( .A(KEYINPUT117), .B(KEYINPUT118), .ZN(n933) );
  XNOR2_X1 U1034 ( .A(n933), .B(KEYINPUT53), .ZN(n945) );
  XNOR2_X1 U1035 ( .A(G2067), .B(G26), .ZN(n935) );
  XNOR2_X1 U1036 ( .A(G33), .B(G2072), .ZN(n934) );
  NOR2_X1 U1037 ( .A1(n935), .A2(n934), .ZN(n940) );
  XOR2_X1 U1038 ( .A(n936), .B(G27), .Z(n938) );
  XNOR2_X1 U1039 ( .A(G1996), .B(G32), .ZN(n937) );
  NOR2_X1 U1040 ( .A1(n938), .A2(n937), .ZN(n939) );
  NAND2_X1 U1041 ( .A1(n940), .A2(n939), .ZN(n943) );
  XOR2_X1 U1042 ( .A(G25), .B(G1991), .Z(n941) );
  NAND2_X1 U1043 ( .A1(n941), .A2(G28), .ZN(n942) );
  NOR2_X1 U1044 ( .A1(n943), .A2(n942), .ZN(n944) );
  XOR2_X1 U1045 ( .A(n945), .B(n944), .Z(n946) );
  NOR2_X1 U1046 ( .A1(n947), .A2(n946), .ZN(n948) );
  XNOR2_X1 U1047 ( .A(KEYINPUT55), .B(n948), .ZN(n950) );
  INV_X1 U1048 ( .A(G29), .ZN(n949) );
  NAND2_X1 U1049 ( .A1(n950), .A2(n949), .ZN(n951) );
  NAND2_X1 U1050 ( .A1(n951), .A2(G11), .ZN(n982) );
  XNOR2_X1 U1051 ( .A(G160), .B(G2084), .ZN(n953) );
  NAND2_X1 U1052 ( .A1(n953), .A2(n952), .ZN(n954) );
  NOR2_X1 U1053 ( .A1(n955), .A2(n954), .ZN(n956) );
  XNOR2_X1 U1054 ( .A(KEYINPUT113), .B(n956), .ZN(n957) );
  NOR2_X1 U1055 ( .A1(n958), .A2(n957), .ZN(n959) );
  NAND2_X1 U1056 ( .A1(n960), .A2(n959), .ZN(n965) );
  XOR2_X1 U1057 ( .A(G2090), .B(G162), .Z(n961) );
  NOR2_X1 U1058 ( .A1(n962), .A2(n961), .ZN(n963) );
  XNOR2_X1 U1059 ( .A(n963), .B(KEYINPUT51), .ZN(n964) );
  NOR2_X1 U1060 ( .A1(n965), .A2(n964), .ZN(n966) );
  XNOR2_X1 U1061 ( .A(n966), .B(KEYINPUT114), .ZN(n968) );
  NAND2_X1 U1062 ( .A1(n968), .A2(n967), .ZN(n969) );
  XOR2_X1 U1063 ( .A(KEYINPUT115), .B(n969), .Z(n975) );
  XOR2_X1 U1064 ( .A(G2072), .B(n970), .Z(n972) );
  XOR2_X1 U1065 ( .A(G164), .B(G2078), .Z(n971) );
  NOR2_X1 U1066 ( .A1(n972), .A2(n971), .ZN(n973) );
  XOR2_X1 U1067 ( .A(KEYINPUT50), .B(n973), .Z(n974) );
  NOR2_X1 U1068 ( .A1(n975), .A2(n974), .ZN(n976) );
  XNOR2_X1 U1069 ( .A(KEYINPUT52), .B(n976), .ZN(n978) );
  INV_X1 U1070 ( .A(KEYINPUT55), .ZN(n977) );
  NAND2_X1 U1071 ( .A1(n978), .A2(n977), .ZN(n979) );
  NAND2_X1 U1072 ( .A1(n979), .A2(G29), .ZN(n980) );
  XOR2_X1 U1073 ( .A(KEYINPUT116), .B(n980), .Z(n981) );
  NOR2_X1 U1074 ( .A1(n982), .A2(n981), .ZN(n1011) );
  XNOR2_X1 U1075 ( .A(G16), .B(KEYINPUT120), .ZN(n983) );
  XNOR2_X1 U1076 ( .A(n983), .B(KEYINPUT56), .ZN(n1009) );
  XOR2_X1 U1077 ( .A(G1966), .B(G168), .Z(n984) );
  NOR2_X1 U1078 ( .A1(n985), .A2(n984), .ZN(n986) );
  XOR2_X1 U1079 ( .A(KEYINPUT57), .B(n986), .Z(n996) );
  XOR2_X1 U1080 ( .A(G1348), .B(KEYINPUT121), .Z(n988) );
  XNOR2_X1 U1081 ( .A(n988), .B(n987), .ZN(n990) );
  NAND2_X1 U1082 ( .A1(G1971), .A2(G303), .ZN(n989) );
  NAND2_X1 U1083 ( .A1(n990), .A2(n989), .ZN(n994) );
  NAND2_X1 U1084 ( .A1(n992), .A2(n991), .ZN(n993) );
  NOR2_X1 U1085 ( .A1(n994), .A2(n993), .ZN(n995) );
  NAND2_X1 U1086 ( .A1(n996), .A2(n995), .ZN(n1000) );
  XNOR2_X1 U1087 ( .A(G1341), .B(n997), .ZN(n998) );
  XNOR2_X1 U1088 ( .A(KEYINPUT122), .B(n998), .ZN(n999) );
  NOR2_X1 U1089 ( .A1(n1000), .A2(n999), .ZN(n1007) );
  XNOR2_X1 U1090 ( .A(n1001), .B(G1956), .ZN(n1003) );
  XNOR2_X1 U1091 ( .A(G171), .B(G1961), .ZN(n1002) );
  NAND2_X1 U1092 ( .A1(n1003), .A2(n1002), .ZN(n1004) );
  NOR2_X1 U1093 ( .A1(n1005), .A2(n1004), .ZN(n1006) );
  NAND2_X1 U1094 ( .A1(n1007), .A2(n1006), .ZN(n1008) );
  NAND2_X1 U1095 ( .A1(n1009), .A2(n1008), .ZN(n1010) );
  NAND2_X1 U1096 ( .A1(n1011), .A2(n1010), .ZN(n1040) );
  XNOR2_X1 U1097 ( .A(G1961), .B(KEYINPUT123), .ZN(n1012) );
  XNOR2_X1 U1098 ( .A(n1012), .B(G5), .ZN(n1020) );
  XNOR2_X1 U1099 ( .A(G1976), .B(G23), .ZN(n1014) );
  XNOR2_X1 U1100 ( .A(G1971), .B(G22), .ZN(n1013) );
  NOR2_X1 U1101 ( .A1(n1014), .A2(n1013), .ZN(n1017) );
  XNOR2_X1 U1102 ( .A(G1986), .B(KEYINPUT127), .ZN(n1015) );
  XNOR2_X1 U1103 ( .A(n1015), .B(G24), .ZN(n1016) );
  NAND2_X1 U1104 ( .A1(n1017), .A2(n1016), .ZN(n1018) );
  XOR2_X1 U1105 ( .A(KEYINPUT58), .B(n1018), .Z(n1019) );
  NAND2_X1 U1106 ( .A1(n1020), .A2(n1019), .ZN(n1036) );
  XOR2_X1 U1107 ( .A(G1341), .B(G19), .Z(n1025) );
  XOR2_X1 U1108 ( .A(KEYINPUT125), .B(G4), .Z(n1022) );
  XNOR2_X1 U1109 ( .A(G1348), .B(KEYINPUT59), .ZN(n1021) );
  XNOR2_X1 U1110 ( .A(n1022), .B(n1021), .ZN(n1023) );
  XNOR2_X1 U1111 ( .A(KEYINPUT124), .B(n1023), .ZN(n1024) );
  NAND2_X1 U1112 ( .A1(n1025), .A2(n1024), .ZN(n1030) );
  XOR2_X1 U1113 ( .A(G1981), .B(G6), .Z(n1028) );
  XNOR2_X1 U1114 ( .A(n1026), .B(G20), .ZN(n1027) );
  NAND2_X1 U1115 ( .A1(n1028), .A2(n1027), .ZN(n1029) );
  NOR2_X1 U1116 ( .A1(n1030), .A2(n1029), .ZN(n1031) );
  XOR2_X1 U1117 ( .A(KEYINPUT60), .B(n1031), .Z(n1033) );
  XNOR2_X1 U1118 ( .A(G1966), .B(G21), .ZN(n1032) );
  NOR2_X1 U1119 ( .A1(n1033), .A2(n1032), .ZN(n1034) );
  XOR2_X1 U1120 ( .A(KEYINPUT126), .B(n1034), .Z(n1035) );
  NOR2_X1 U1121 ( .A1(n1036), .A2(n1035), .ZN(n1037) );
  XOR2_X1 U1122 ( .A(KEYINPUT61), .B(n1037), .Z(n1038) );
  NOR2_X1 U1123 ( .A1(G16), .A2(n1038), .ZN(n1039) );
  NOR2_X1 U1124 ( .A1(n1040), .A2(n1039), .ZN(n1041) );
  XNOR2_X1 U1125 ( .A(n1041), .B(KEYINPUT62), .ZN(G311) );
  INV_X1 U1126 ( .A(G311), .ZN(G150) );
endmodule

