

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300,
         n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311,
         n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322,
         n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333,
         n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344,
         n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581;

  XNOR2_X1 U322 ( .A(KEYINPUT121), .B(n471), .ZN(n562) );
  XNOR2_X1 U323 ( .A(n448), .B(n447), .ZN(n496) );
  XNOR2_X1 U324 ( .A(n413), .B(n412), .ZN(n517) );
  XOR2_X1 U325 ( .A(KEYINPUT25), .B(n434), .Z(n290) );
  XOR2_X1 U326 ( .A(KEYINPUT86), .B(KEYINPUT17), .Z(n291) );
  XNOR2_X1 U327 ( .A(n415), .B(n403), .ZN(n404) );
  XNOR2_X1 U328 ( .A(n405), .B(n404), .ZN(n406) );
  XNOR2_X1 U329 ( .A(n314), .B(n313), .ZN(n315) );
  XNOR2_X1 U330 ( .A(KEYINPUT48), .B(KEYINPUT64), .ZN(n463) );
  XNOR2_X1 U331 ( .A(n414), .B(n315), .ZN(n319) );
  XNOR2_X1 U332 ( .A(n464), .B(n463), .ZN(n527) );
  XNOR2_X1 U333 ( .A(n326), .B(n325), .ZN(n327) );
  XNOR2_X1 U334 ( .A(n328), .B(n327), .ZN(n571) );
  INV_X1 U335 ( .A(G36GAT), .ZN(n449) );
  XNOR2_X1 U336 ( .A(n473), .B(n472), .ZN(n474) );
  XNOR2_X1 U337 ( .A(n449), .B(KEYINPUT104), .ZN(n450) );
  XNOR2_X1 U338 ( .A(n475), .B(n474), .ZN(G1351GAT) );
  XNOR2_X1 U339 ( .A(n451), .B(n450), .ZN(G1329GAT) );
  XOR2_X1 U340 ( .A(KEYINPUT103), .B(KEYINPUT38), .Z(n448) );
  XOR2_X1 U341 ( .A(G8GAT), .B(KEYINPUT29), .Z(n293) );
  XNOR2_X1 U342 ( .A(KEYINPUT68), .B(KEYINPUT30), .ZN(n292) );
  XNOR2_X1 U343 ( .A(n293), .B(n292), .ZN(n311) );
  XOR2_X1 U344 ( .A(G22GAT), .B(G141GAT), .Z(n295) );
  XNOR2_X1 U345 ( .A(G50GAT), .B(G36GAT), .ZN(n294) );
  XNOR2_X1 U346 ( .A(n295), .B(n294), .ZN(n299) );
  XOR2_X1 U347 ( .A(G15GAT), .B(G113GAT), .Z(n297) );
  XNOR2_X1 U348 ( .A(G169GAT), .B(G197GAT), .ZN(n296) );
  XNOR2_X1 U349 ( .A(n297), .B(n296), .ZN(n298) );
  XOR2_X1 U350 ( .A(n299), .B(n298), .Z(n309) );
  XOR2_X1 U351 ( .A(KEYINPUT73), .B(KEYINPUT71), .Z(n301) );
  XNOR2_X1 U352 ( .A(KEYINPUT70), .B(KEYINPUT69), .ZN(n300) );
  XNOR2_X1 U353 ( .A(n301), .B(n300), .ZN(n307) );
  XOR2_X1 U354 ( .A(G29GAT), .B(G43GAT), .Z(n303) );
  XNOR2_X1 U355 ( .A(KEYINPUT8), .B(KEYINPUT7), .ZN(n302) );
  XNOR2_X1 U356 ( .A(n303), .B(n302), .ZN(n346) );
  XOR2_X1 U357 ( .A(KEYINPUT72), .B(G1GAT), .Z(n340) );
  XOR2_X1 U358 ( .A(n346), .B(n340), .Z(n305) );
  NAND2_X1 U359 ( .A1(G229GAT), .A2(G233GAT), .ZN(n304) );
  XNOR2_X1 U360 ( .A(n305), .B(n304), .ZN(n306) );
  XNOR2_X1 U361 ( .A(n307), .B(n306), .ZN(n308) );
  XNOR2_X1 U362 ( .A(n309), .B(n308), .ZN(n310) );
  XNOR2_X1 U363 ( .A(n311), .B(n310), .ZN(n555) );
  INV_X1 U364 ( .A(n555), .ZN(n567) );
  XNOR2_X1 U365 ( .A(G106GAT), .B(G78GAT), .ZN(n312) );
  XNOR2_X1 U366 ( .A(n312), .B(G148GAT), .ZN(n414) );
  NAND2_X1 U367 ( .A1(G230GAT), .A2(G233GAT), .ZN(n314) );
  INV_X1 U368 ( .A(KEYINPUT76), .ZN(n313) );
  XOR2_X1 U369 ( .A(KEYINPUT33), .B(KEYINPUT77), .Z(n317) );
  XNOR2_X1 U370 ( .A(KEYINPUT32), .B(KEYINPUT75), .ZN(n316) );
  XNOR2_X1 U371 ( .A(n317), .B(n316), .ZN(n318) );
  XOR2_X1 U372 ( .A(n319), .B(n318), .Z(n328) );
  XOR2_X1 U373 ( .A(KEYINPUT74), .B(KEYINPUT13), .Z(n321) );
  XNOR2_X1 U374 ( .A(G71GAT), .B(G57GAT), .ZN(n320) );
  XNOR2_X1 U375 ( .A(n321), .B(n320), .ZN(n333) );
  XOR2_X1 U376 ( .A(G64GAT), .B(G92GAT), .Z(n323) );
  XNOR2_X1 U377 ( .A(G176GAT), .B(G204GAT), .ZN(n322) );
  XNOR2_X1 U378 ( .A(n323), .B(n322), .ZN(n411) );
  XNOR2_X1 U379 ( .A(n333), .B(n411), .ZN(n326) );
  XNOR2_X1 U380 ( .A(G120GAT), .B(KEYINPUT31), .ZN(n324) );
  XNOR2_X1 U381 ( .A(G99GAT), .B(G85GAT), .ZN(n343) );
  XNOR2_X1 U382 ( .A(n324), .B(n343), .ZN(n325) );
  INV_X1 U383 ( .A(n571), .ZN(n460) );
  NOR2_X1 U384 ( .A1(n567), .A2(n460), .ZN(n480) );
  XNOR2_X1 U385 ( .A(G8GAT), .B(G183GAT), .ZN(n329) );
  XOR2_X1 U386 ( .A(n329), .B(G211GAT), .Z(n412) );
  XOR2_X1 U387 ( .A(G22GAT), .B(G155GAT), .Z(n418) );
  XNOR2_X1 U388 ( .A(n412), .B(n418), .ZN(n331) );
  NAND2_X1 U389 ( .A1(G231GAT), .A2(G233GAT), .ZN(n330) );
  XNOR2_X1 U390 ( .A(n331), .B(n330), .ZN(n332) );
  XOR2_X1 U391 ( .A(n332), .B(KEYINPUT12), .Z(n335) );
  XNOR2_X1 U392 ( .A(n333), .B(KEYINPUT15), .ZN(n334) );
  XNOR2_X1 U393 ( .A(n335), .B(n334), .ZN(n339) );
  XOR2_X1 U394 ( .A(KEYINPUT14), .B(KEYINPUT81), .Z(n337) );
  XNOR2_X1 U395 ( .A(G78GAT), .B(G64GAT), .ZN(n336) );
  XOR2_X1 U396 ( .A(n337), .B(n336), .Z(n338) );
  XNOR2_X1 U397 ( .A(n339), .B(n338), .ZN(n342) );
  XOR2_X1 U398 ( .A(G15GAT), .B(G127GAT), .Z(n393) );
  XNOR2_X1 U399 ( .A(n340), .B(n393), .ZN(n341) );
  XNOR2_X1 U400 ( .A(n342), .B(n341), .ZN(n476) );
  XOR2_X1 U401 ( .A(G36GAT), .B(G190GAT), .Z(n407) );
  XNOR2_X1 U402 ( .A(n407), .B(n343), .ZN(n345) );
  XOR2_X1 U403 ( .A(G50GAT), .B(G162GAT), .Z(n419) );
  XOR2_X1 U404 ( .A(G134GAT), .B(KEYINPUT80), .Z(n374) );
  XNOR2_X1 U405 ( .A(n419), .B(n374), .ZN(n344) );
  XNOR2_X1 U406 ( .A(n345), .B(n344), .ZN(n350) );
  XOR2_X1 U407 ( .A(G92GAT), .B(n346), .Z(n348) );
  NAND2_X1 U408 ( .A1(G232GAT), .A2(G233GAT), .ZN(n347) );
  XNOR2_X1 U409 ( .A(n348), .B(n347), .ZN(n349) );
  XOR2_X1 U410 ( .A(n350), .B(n349), .Z(n358) );
  XOR2_X1 U411 ( .A(KEYINPUT66), .B(KEYINPUT11), .Z(n352) );
  XNOR2_X1 U412 ( .A(G218GAT), .B(KEYINPUT78), .ZN(n351) );
  XNOR2_X1 U413 ( .A(n352), .B(n351), .ZN(n356) );
  XOR2_X1 U414 ( .A(KEYINPUT10), .B(KEYINPUT9), .Z(n354) );
  XNOR2_X1 U415 ( .A(G106GAT), .B(KEYINPUT79), .ZN(n353) );
  XNOR2_X1 U416 ( .A(n354), .B(n353), .ZN(n355) );
  XNOR2_X1 U417 ( .A(n356), .B(n355), .ZN(n357) );
  XNOR2_X1 U418 ( .A(n358), .B(n357), .ZN(n552) );
  XNOR2_X1 U419 ( .A(KEYINPUT36), .B(n552), .ZN(n578) );
  NOR2_X1 U420 ( .A1(n476), .A2(n578), .ZN(n445) );
  XOR2_X1 U421 ( .A(KEYINPUT0), .B(KEYINPUT83), .Z(n360) );
  XNOR2_X1 U422 ( .A(KEYINPUT82), .B(G120GAT), .ZN(n359) );
  XNOR2_X1 U423 ( .A(n360), .B(n359), .ZN(n361) );
  XOR2_X1 U424 ( .A(G113GAT), .B(n361), .Z(n400) );
  XOR2_X1 U425 ( .A(KEYINPUT1), .B(KEYINPUT95), .Z(n363) );
  XNOR2_X1 U426 ( .A(G1GAT), .B(G57GAT), .ZN(n362) );
  XNOR2_X1 U427 ( .A(n363), .B(n362), .ZN(n367) );
  XOR2_X1 U428 ( .A(KEYINPUT5), .B(KEYINPUT93), .Z(n365) );
  XNOR2_X1 U429 ( .A(KEYINPUT6), .B(KEYINPUT94), .ZN(n364) );
  XNOR2_X1 U430 ( .A(n365), .B(n364), .ZN(n366) );
  XOR2_X1 U431 ( .A(n367), .B(n366), .Z(n380) );
  XNOR2_X1 U432 ( .A(G141GAT), .B(KEYINPUT3), .ZN(n368) );
  XNOR2_X1 U433 ( .A(n368), .B(KEYINPUT2), .ZN(n427) );
  XOR2_X1 U434 ( .A(KEYINPUT4), .B(n427), .Z(n370) );
  NAND2_X1 U435 ( .A1(G225GAT), .A2(G233GAT), .ZN(n369) );
  XNOR2_X1 U436 ( .A(n370), .B(n369), .ZN(n378) );
  XOR2_X1 U437 ( .A(G155GAT), .B(G162GAT), .Z(n372) );
  XNOR2_X1 U438 ( .A(G127GAT), .B(G148GAT), .ZN(n371) );
  XNOR2_X1 U439 ( .A(n372), .B(n371), .ZN(n373) );
  XOR2_X1 U440 ( .A(n373), .B(G85GAT), .Z(n376) );
  XNOR2_X1 U441 ( .A(G29GAT), .B(n374), .ZN(n375) );
  XNOR2_X1 U442 ( .A(n376), .B(n375), .ZN(n377) );
  XNOR2_X1 U443 ( .A(n378), .B(n377), .ZN(n379) );
  XNOR2_X1 U444 ( .A(n380), .B(n379), .ZN(n381) );
  XNOR2_X1 U445 ( .A(n400), .B(n381), .ZN(n440) );
  INV_X1 U446 ( .A(n440), .ZN(n514) );
  XOR2_X1 U447 ( .A(G71GAT), .B(KEYINPUT20), .Z(n383) );
  XNOR2_X1 U448 ( .A(KEYINPUT85), .B(KEYINPUT84), .ZN(n382) );
  XNOR2_X1 U449 ( .A(n383), .B(n382), .ZN(n387) );
  XOR2_X1 U450 ( .A(G176GAT), .B(G183GAT), .Z(n385) );
  XNOR2_X1 U451 ( .A(KEYINPUT87), .B(KEYINPUT88), .ZN(n384) );
  XNOR2_X1 U452 ( .A(n385), .B(n384), .ZN(n386) );
  XOR2_X1 U453 ( .A(n387), .B(n386), .Z(n398) );
  XNOR2_X1 U454 ( .A(KEYINPUT19), .B(KEYINPUT18), .ZN(n388) );
  XNOR2_X1 U455 ( .A(n291), .B(n388), .ZN(n389) );
  XOR2_X1 U456 ( .A(G169GAT), .B(n389), .Z(n405) );
  XOR2_X1 U457 ( .A(G190GAT), .B(G134GAT), .Z(n391) );
  XNOR2_X1 U458 ( .A(G43GAT), .B(G99GAT), .ZN(n390) );
  XNOR2_X1 U459 ( .A(n391), .B(n390), .ZN(n392) );
  XOR2_X1 U460 ( .A(n393), .B(n392), .Z(n395) );
  NAND2_X1 U461 ( .A1(G227GAT), .A2(G233GAT), .ZN(n394) );
  XNOR2_X1 U462 ( .A(n395), .B(n394), .ZN(n396) );
  XNOR2_X1 U463 ( .A(n405), .B(n396), .ZN(n397) );
  XNOR2_X1 U464 ( .A(n398), .B(n397), .ZN(n399) );
  XNOR2_X1 U465 ( .A(n400), .B(n399), .ZN(n528) );
  INV_X1 U466 ( .A(n528), .ZN(n519) );
  XOR2_X1 U467 ( .A(KEYINPUT90), .B(KEYINPUT21), .Z(n402) );
  XNOR2_X1 U468 ( .A(G197GAT), .B(G218GAT), .ZN(n401) );
  XNOR2_X1 U469 ( .A(n402), .B(n401), .ZN(n415) );
  XOR2_X1 U470 ( .A(KEYINPUT96), .B(KEYINPUT97), .Z(n403) );
  XOR2_X1 U471 ( .A(n407), .B(n406), .Z(n409) );
  NAND2_X1 U472 ( .A1(G226GAT), .A2(G233GAT), .ZN(n408) );
  XNOR2_X1 U473 ( .A(n409), .B(n408), .ZN(n410) );
  XNOR2_X1 U474 ( .A(n411), .B(n410), .ZN(n413) );
  OR2_X1 U475 ( .A1(n519), .A2(n517), .ZN(n432) );
  XNOR2_X1 U476 ( .A(n415), .B(n414), .ZN(n431) );
  XOR2_X1 U477 ( .A(KEYINPUT22), .B(KEYINPUT92), .Z(n417) );
  XNOR2_X1 U478 ( .A(G211GAT), .B(G204GAT), .ZN(n416) );
  XNOR2_X1 U479 ( .A(n417), .B(n416), .ZN(n423) );
  XOR2_X1 U480 ( .A(KEYINPUT24), .B(KEYINPUT89), .Z(n421) );
  XNOR2_X1 U481 ( .A(n419), .B(n418), .ZN(n420) );
  XNOR2_X1 U482 ( .A(n421), .B(n420), .ZN(n422) );
  XOR2_X1 U483 ( .A(n423), .B(n422), .Z(n425) );
  NAND2_X1 U484 ( .A1(G228GAT), .A2(G233GAT), .ZN(n424) );
  XNOR2_X1 U485 ( .A(n425), .B(n424), .ZN(n426) );
  XOR2_X1 U486 ( .A(n426), .B(KEYINPUT91), .Z(n429) );
  XNOR2_X1 U487 ( .A(n427), .B(KEYINPUT23), .ZN(n428) );
  XNOR2_X1 U488 ( .A(n429), .B(n428), .ZN(n430) );
  XNOR2_X1 U489 ( .A(n431), .B(n430), .ZN(n468) );
  NAND2_X1 U490 ( .A1(n432), .A2(n468), .ZN(n433) );
  XNOR2_X1 U491 ( .A(n433), .B(KEYINPUT98), .ZN(n434) );
  XOR2_X1 U492 ( .A(KEYINPUT27), .B(n517), .Z(n439) );
  NOR2_X1 U493 ( .A1(n528), .A2(n468), .ZN(n435) );
  XNOR2_X1 U494 ( .A(n435), .B(KEYINPUT26), .ZN(n565) );
  NAND2_X1 U495 ( .A1(n439), .A2(n565), .ZN(n436) );
  NAND2_X1 U496 ( .A1(n290), .A2(n436), .ZN(n437) );
  NAND2_X1 U497 ( .A1(n514), .A2(n437), .ZN(n438) );
  XOR2_X1 U498 ( .A(KEYINPUT99), .B(n438), .Z(n444) );
  NAND2_X1 U499 ( .A1(n440), .A2(n439), .ZN(n526) );
  NOR2_X1 U500 ( .A1(n528), .A2(n526), .ZN(n442) );
  XOR2_X1 U501 ( .A(n468), .B(KEYINPUT67), .Z(n441) );
  XNOR2_X1 U502 ( .A(KEYINPUT28), .B(n441), .ZN(n531) );
  NAND2_X1 U503 ( .A1(n442), .A2(n531), .ZN(n443) );
  NAND2_X1 U504 ( .A1(n444), .A2(n443), .ZN(n479) );
  NAND2_X1 U505 ( .A1(n445), .A2(n479), .ZN(n446) );
  XNOR2_X1 U506 ( .A(KEYINPUT37), .B(n446), .ZN(n513) );
  NAND2_X1 U507 ( .A1(n480), .A2(n513), .ZN(n447) );
  NOR2_X1 U508 ( .A1(n496), .A2(n517), .ZN(n451) );
  XNOR2_X1 U509 ( .A(n476), .B(KEYINPUT114), .ZN(n561) );
  XOR2_X1 U510 ( .A(n571), .B(KEYINPUT41), .Z(n546) );
  INV_X1 U511 ( .A(n546), .ZN(n499) );
  NAND2_X1 U512 ( .A1(n499), .A2(n555), .ZN(n453) );
  XOR2_X1 U513 ( .A(KEYINPUT115), .B(KEYINPUT46), .Z(n452) );
  XOR2_X1 U514 ( .A(n453), .B(n452), .Z(n454) );
  NOR2_X1 U515 ( .A1(n561), .A2(n454), .ZN(n455) );
  NAND2_X1 U516 ( .A1(n455), .A2(n552), .ZN(n456) );
  XNOR2_X1 U517 ( .A(n456), .B(KEYINPUT47), .ZN(n462) );
  INV_X1 U518 ( .A(n476), .ZN(n574) );
  NOR2_X1 U519 ( .A1(n578), .A2(n574), .ZN(n457) );
  XNOR2_X1 U520 ( .A(KEYINPUT45), .B(n457), .ZN(n458) );
  NAND2_X1 U521 ( .A1(n458), .A2(n567), .ZN(n459) );
  NOR2_X1 U522 ( .A1(n460), .A2(n459), .ZN(n461) );
  NOR2_X1 U523 ( .A1(n462), .A2(n461), .ZN(n464) );
  NOR2_X1 U524 ( .A1(n527), .A2(n517), .ZN(n465) );
  XNOR2_X1 U525 ( .A(n465), .B(KEYINPUT54), .ZN(n466) );
  NAND2_X1 U526 ( .A1(n466), .A2(n514), .ZN(n467) );
  XNOR2_X1 U527 ( .A(n467), .B(KEYINPUT65), .ZN(n566) );
  NAND2_X1 U528 ( .A1(n468), .A2(n566), .ZN(n469) );
  XNOR2_X1 U529 ( .A(n469), .B(KEYINPUT55), .ZN(n470) );
  NAND2_X1 U530 ( .A1(n470), .A2(n528), .ZN(n471) );
  INV_X1 U531 ( .A(n552), .ZN(n539) );
  NAND2_X1 U532 ( .A1(n562), .A2(n539), .ZN(n475) );
  XOR2_X1 U533 ( .A(KEYINPUT124), .B(KEYINPUT58), .Z(n473) );
  INV_X1 U534 ( .A(G190GAT), .ZN(n472) );
  NAND2_X1 U535 ( .A1(n552), .A2(n476), .ZN(n477) );
  XOR2_X1 U536 ( .A(KEYINPUT16), .B(n477), .Z(n478) );
  AND2_X1 U537 ( .A1(n479), .A2(n478), .ZN(n501) );
  NAND2_X1 U538 ( .A1(n480), .A2(n501), .ZN(n489) );
  NOR2_X1 U539 ( .A1(n514), .A2(n489), .ZN(n482) );
  XNOR2_X1 U540 ( .A(KEYINPUT34), .B(KEYINPUT100), .ZN(n481) );
  XNOR2_X1 U541 ( .A(n482), .B(n481), .ZN(n483) );
  XOR2_X1 U542 ( .A(G1GAT), .B(n483), .Z(G1324GAT) );
  NOR2_X1 U543 ( .A1(n517), .A2(n489), .ZN(n485) );
  XNOR2_X1 U544 ( .A(G8GAT), .B(KEYINPUT101), .ZN(n484) );
  XNOR2_X1 U545 ( .A(n485), .B(n484), .ZN(G1325GAT) );
  NOR2_X1 U546 ( .A1(n519), .A2(n489), .ZN(n487) );
  XNOR2_X1 U547 ( .A(KEYINPUT102), .B(KEYINPUT35), .ZN(n486) );
  XNOR2_X1 U548 ( .A(n487), .B(n486), .ZN(n488) );
  XNOR2_X1 U549 ( .A(G15GAT), .B(n488), .ZN(G1326GAT) );
  NOR2_X1 U550 ( .A1(n531), .A2(n489), .ZN(n490) );
  XOR2_X1 U551 ( .A(G22GAT), .B(n490), .Z(G1327GAT) );
  NOR2_X1 U552 ( .A1(n514), .A2(n496), .ZN(n491) );
  XNOR2_X1 U553 ( .A(n491), .B(KEYINPUT39), .ZN(n492) );
  XNOR2_X1 U554 ( .A(G29GAT), .B(n492), .ZN(G1328GAT) );
  XNOR2_X1 U555 ( .A(KEYINPUT40), .B(KEYINPUT105), .ZN(n494) );
  NOR2_X1 U556 ( .A1(n519), .A2(n496), .ZN(n493) );
  XNOR2_X1 U557 ( .A(n494), .B(n493), .ZN(n495) );
  XNOR2_X1 U558 ( .A(G43GAT), .B(n495), .ZN(G1330GAT) );
  NOR2_X1 U559 ( .A1(n496), .A2(n531), .ZN(n497) );
  XOR2_X1 U560 ( .A(KEYINPUT106), .B(n497), .Z(n498) );
  XNOR2_X1 U561 ( .A(G50GAT), .B(n498), .ZN(G1331GAT) );
  NAND2_X1 U562 ( .A1(n499), .A2(n567), .ZN(n500) );
  XNOR2_X1 U563 ( .A(n500), .B(KEYINPUT107), .ZN(n512) );
  NAND2_X1 U564 ( .A1(n512), .A2(n501), .ZN(n509) );
  NOR2_X1 U565 ( .A1(n514), .A2(n509), .ZN(n503) );
  XNOR2_X1 U566 ( .A(KEYINPUT108), .B(KEYINPUT42), .ZN(n502) );
  XNOR2_X1 U567 ( .A(n503), .B(n502), .ZN(n504) );
  XOR2_X1 U568 ( .A(G57GAT), .B(n504), .Z(G1332GAT) );
  NOR2_X1 U569 ( .A1(n517), .A2(n509), .ZN(n506) );
  XNOR2_X1 U570 ( .A(G64GAT), .B(KEYINPUT109), .ZN(n505) );
  XNOR2_X1 U571 ( .A(n506), .B(n505), .ZN(G1333GAT) );
  NOR2_X1 U572 ( .A1(n519), .A2(n509), .ZN(n507) );
  XOR2_X1 U573 ( .A(KEYINPUT110), .B(n507), .Z(n508) );
  XNOR2_X1 U574 ( .A(G71GAT), .B(n508), .ZN(G1334GAT) );
  NOR2_X1 U575 ( .A1(n531), .A2(n509), .ZN(n511) );
  XNOR2_X1 U576 ( .A(G78GAT), .B(KEYINPUT43), .ZN(n510) );
  XNOR2_X1 U577 ( .A(n511), .B(n510), .ZN(G1335GAT) );
  NAND2_X1 U578 ( .A1(n513), .A2(n512), .ZN(n522) );
  NOR2_X1 U579 ( .A1(n514), .A2(n522), .ZN(n515) );
  XNOR2_X1 U580 ( .A(n515), .B(KEYINPUT111), .ZN(n516) );
  XNOR2_X1 U581 ( .A(G85GAT), .B(n516), .ZN(G1336GAT) );
  NOR2_X1 U582 ( .A1(n517), .A2(n522), .ZN(n518) );
  XOR2_X1 U583 ( .A(G92GAT), .B(n518), .Z(G1337GAT) );
  NOR2_X1 U584 ( .A1(n519), .A2(n522), .ZN(n520) );
  XOR2_X1 U585 ( .A(KEYINPUT112), .B(n520), .Z(n521) );
  XNOR2_X1 U586 ( .A(G99GAT), .B(n521), .ZN(G1338GAT) );
  NOR2_X1 U587 ( .A1(n531), .A2(n522), .ZN(n524) );
  XNOR2_X1 U588 ( .A(KEYINPUT44), .B(KEYINPUT113), .ZN(n523) );
  XNOR2_X1 U589 ( .A(n524), .B(n523), .ZN(n525) );
  XNOR2_X1 U590 ( .A(G106GAT), .B(n525), .ZN(G1339GAT) );
  NOR2_X1 U591 ( .A1(n527), .A2(n526), .ZN(n544) );
  NAND2_X1 U592 ( .A1(n544), .A2(n528), .ZN(n529) );
  XOR2_X1 U593 ( .A(KEYINPUT116), .B(n529), .Z(n530) );
  NAND2_X1 U594 ( .A1(n531), .A2(n530), .ZN(n532) );
  XNOR2_X1 U595 ( .A(n532), .B(KEYINPUT117), .ZN(n540) );
  NAND2_X1 U596 ( .A1(n540), .A2(n555), .ZN(n533) );
  XNOR2_X1 U597 ( .A(G113GAT), .B(n533), .ZN(G1340GAT) );
  XOR2_X1 U598 ( .A(KEYINPUT118), .B(KEYINPUT49), .Z(n535) );
  NAND2_X1 U599 ( .A1(n540), .A2(n499), .ZN(n534) );
  XNOR2_X1 U600 ( .A(n535), .B(n534), .ZN(n536) );
  XNOR2_X1 U601 ( .A(G120GAT), .B(n536), .ZN(G1341GAT) );
  NAND2_X1 U602 ( .A1(n561), .A2(n540), .ZN(n537) );
  XNOR2_X1 U603 ( .A(n537), .B(KEYINPUT50), .ZN(n538) );
  XNOR2_X1 U604 ( .A(G127GAT), .B(n538), .ZN(G1342GAT) );
  XOR2_X1 U605 ( .A(KEYINPUT51), .B(KEYINPUT119), .Z(n542) );
  NAND2_X1 U606 ( .A1(n540), .A2(n539), .ZN(n541) );
  XNOR2_X1 U607 ( .A(n542), .B(n541), .ZN(n543) );
  XOR2_X1 U608 ( .A(G134GAT), .B(n543), .Z(G1343GAT) );
  NAND2_X1 U609 ( .A1(n544), .A2(n565), .ZN(n551) );
  NOR2_X1 U610 ( .A1(n567), .A2(n551), .ZN(n545) );
  XOR2_X1 U611 ( .A(G141GAT), .B(n545), .Z(G1344GAT) );
  NOR2_X1 U612 ( .A1(n546), .A2(n551), .ZN(n548) );
  XNOR2_X1 U613 ( .A(KEYINPUT53), .B(KEYINPUT52), .ZN(n547) );
  XNOR2_X1 U614 ( .A(n548), .B(n547), .ZN(n549) );
  XNOR2_X1 U615 ( .A(G148GAT), .B(n549), .ZN(G1345GAT) );
  NOR2_X1 U616 ( .A1(n574), .A2(n551), .ZN(n550) );
  XOR2_X1 U617 ( .A(G155GAT), .B(n550), .Z(G1346GAT) );
  NOR2_X1 U618 ( .A1(n552), .A2(n551), .ZN(n553) );
  XOR2_X1 U619 ( .A(KEYINPUT120), .B(n553), .Z(n554) );
  XNOR2_X1 U620 ( .A(G162GAT), .B(n554), .ZN(G1347GAT) );
  NAND2_X1 U621 ( .A1(n555), .A2(n562), .ZN(n556) );
  XNOR2_X1 U622 ( .A(n556), .B(G169GAT), .ZN(G1348GAT) );
  NAND2_X1 U623 ( .A1(n562), .A2(n499), .ZN(n558) );
  XOR2_X1 U624 ( .A(KEYINPUT122), .B(KEYINPUT57), .Z(n557) );
  XNOR2_X1 U625 ( .A(n558), .B(n557), .ZN(n560) );
  XNOR2_X1 U626 ( .A(G176GAT), .B(KEYINPUT56), .ZN(n559) );
  XNOR2_X1 U627 ( .A(n560), .B(n559), .ZN(G1349GAT) );
  XOR2_X1 U628 ( .A(G183GAT), .B(KEYINPUT123), .Z(n564) );
  NAND2_X1 U629 ( .A1(n562), .A2(n561), .ZN(n563) );
  XNOR2_X1 U630 ( .A(n564), .B(n563), .ZN(G1350GAT) );
  NAND2_X1 U631 ( .A1(n566), .A2(n565), .ZN(n577) );
  NOR2_X1 U632 ( .A1(n567), .A2(n577), .ZN(n569) );
  XNOR2_X1 U633 ( .A(KEYINPUT60), .B(KEYINPUT59), .ZN(n568) );
  XNOR2_X1 U634 ( .A(n569), .B(n568), .ZN(n570) );
  XNOR2_X1 U635 ( .A(G197GAT), .B(n570), .ZN(G1352GAT) );
  NOR2_X1 U636 ( .A1(n571), .A2(n577), .ZN(n573) );
  XNOR2_X1 U637 ( .A(G204GAT), .B(KEYINPUT61), .ZN(n572) );
  XNOR2_X1 U638 ( .A(n573), .B(n572), .ZN(G1353GAT) );
  NOR2_X1 U639 ( .A1(n574), .A2(n577), .ZN(n576) );
  XNOR2_X1 U640 ( .A(G211GAT), .B(KEYINPUT125), .ZN(n575) );
  XNOR2_X1 U641 ( .A(n576), .B(n575), .ZN(G1354GAT) );
  NOR2_X1 U642 ( .A1(n578), .A2(n577), .ZN(n580) );
  XNOR2_X1 U643 ( .A(KEYINPUT62), .B(KEYINPUT126), .ZN(n579) );
  XNOR2_X1 U644 ( .A(n580), .B(n579), .ZN(n581) );
  XOR2_X1 U645 ( .A(G218GAT), .B(n581), .Z(G1355GAT) );
endmodule

