//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 0 0 1 0 1 0 1 1 0 1 1 0 1 0 0 0 1 1 1 0 1 0 1 1 1 1 0 1 0 0 0 1 1 1 1 1 0 0 1 0 0 0 1 0 0 1 1 0 1 0 0 1 1 1 0 0 1 0 0 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:19:54 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n684, new_n685, new_n686, new_n687,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n723, new_n724,
    new_n725, new_n726, new_n727, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n757, new_n758, new_n759, new_n761, new_n762, new_n763, new_n765,
    new_n766, new_n767, new_n768, new_n770, new_n771, new_n772, new_n773,
    new_n774, new_n775, new_n776, new_n777, new_n778, new_n779, new_n780,
    new_n781, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n794, new_n795, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n841,
    new_n842, new_n843, new_n845, new_n846, new_n847, new_n849, new_n850,
    new_n851, new_n852, new_n853, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n928, new_n929, new_n931,
    new_n932, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n946, new_n947,
    new_n948, new_n949, new_n951, new_n952, new_n953, new_n954, new_n955,
    new_n956, new_n957, new_n958, new_n960, new_n961, new_n962, new_n964,
    new_n965, new_n966, new_n967, new_n968, new_n969, new_n970, new_n971,
    new_n972, new_n974, new_n975, new_n976, new_n977, new_n979, new_n980,
    new_n981, new_n982, new_n983, new_n984, new_n985, new_n986, new_n987,
    new_n988, new_n990, new_n991;
  XNOR2_X1  g000(.A(G15gat), .B(G22gat), .ZN(new_n202));
  INV_X1    g001(.A(G1gat), .ZN(new_n203));
  NAND2_X1  g002(.A1(new_n203), .A2(KEYINPUT16), .ZN(new_n204));
  NAND2_X1  g003(.A1(new_n202), .A2(new_n204), .ZN(new_n205));
  OAI21_X1  g004(.A(new_n205), .B1(G1gat), .B2(new_n202), .ZN(new_n206));
  XNOR2_X1  g005(.A(new_n206), .B(G8gat), .ZN(new_n207));
  INV_X1    g006(.A(new_n207), .ZN(new_n208));
  INV_X1    g007(.A(KEYINPUT17), .ZN(new_n209));
  INV_X1    g008(.A(G29gat), .ZN(new_n210));
  NAND3_X1  g009(.A1(new_n210), .A2(KEYINPUT14), .A3(G36gat), .ZN(new_n211));
  XOR2_X1   g010(.A(KEYINPUT14), .B(G29gat), .Z(new_n212));
  OAI21_X1  g011(.A(new_n211), .B1(new_n212), .B2(G36gat), .ZN(new_n213));
  INV_X1    g012(.A(KEYINPUT15), .ZN(new_n214));
  INV_X1    g013(.A(G43gat), .ZN(new_n215));
  INV_X1    g014(.A(G50gat), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  NAND2_X1  g016(.A1(G43gat), .A2(G50gat), .ZN(new_n218));
  AOI21_X1  g017(.A(new_n214), .B1(new_n217), .B2(new_n218), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n213), .A2(new_n219), .ZN(new_n220));
  XNOR2_X1  g019(.A(KEYINPUT88), .B(G50gat), .ZN(new_n221));
  OAI211_X1 g020(.A(new_n214), .B(new_n218), .C1(new_n221), .C2(G43gat), .ZN(new_n222));
  AND2_X1   g021(.A1(new_n213), .A2(new_n222), .ZN(new_n223));
  OAI211_X1 g022(.A(new_n209), .B(new_n220), .C1(new_n223), .C2(new_n219), .ZN(new_n224));
  INV_X1    g023(.A(new_n220), .ZN(new_n225));
  AOI21_X1  g024(.A(new_n219), .B1(new_n213), .B2(new_n222), .ZN(new_n226));
  OAI21_X1  g025(.A(KEYINPUT17), .B1(new_n225), .B2(new_n226), .ZN(new_n227));
  NAND3_X1  g026(.A1(new_n208), .A2(new_n224), .A3(new_n227), .ZN(new_n228));
  NOR2_X1   g027(.A1(new_n225), .A2(new_n226), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n229), .A2(new_n207), .ZN(new_n230));
  NAND2_X1  g029(.A1(G229gat), .A2(G233gat), .ZN(new_n231));
  NAND3_X1  g030(.A1(new_n228), .A2(new_n230), .A3(new_n231), .ZN(new_n232));
  INV_X1    g031(.A(KEYINPUT18), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n232), .A2(new_n233), .ZN(new_n234));
  INV_X1    g033(.A(new_n234), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n235), .A2(KEYINPUT90), .ZN(new_n236));
  XNOR2_X1  g035(.A(G113gat), .B(G141gat), .ZN(new_n237));
  INV_X1    g036(.A(G197gat), .ZN(new_n238));
  XNOR2_X1  g037(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XNOR2_X1  g038(.A(KEYINPUT11), .B(G169gat), .ZN(new_n240));
  XNOR2_X1  g039(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XOR2_X1   g040(.A(new_n241), .B(KEYINPUT12), .Z(new_n242));
  INV_X1    g041(.A(new_n242), .ZN(new_n243));
  XNOR2_X1  g042(.A(new_n229), .B(new_n207), .ZN(new_n244));
  XOR2_X1   g043(.A(new_n231), .B(KEYINPUT13), .Z(new_n245));
  NAND2_X1  g044(.A1(new_n244), .A2(new_n245), .ZN(new_n246));
  NAND4_X1  g045(.A1(new_n228), .A2(KEYINPUT18), .A3(new_n230), .A4(new_n231), .ZN(new_n247));
  AND3_X1   g046(.A1(new_n243), .A2(new_n246), .A3(new_n247), .ZN(new_n248));
  INV_X1    g047(.A(KEYINPUT90), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n234), .A2(new_n249), .ZN(new_n250));
  NAND3_X1  g049(.A1(new_n236), .A2(new_n248), .A3(new_n250), .ZN(new_n251));
  INV_X1    g050(.A(KEYINPUT89), .ZN(new_n252));
  AND3_X1   g051(.A1(new_n246), .A2(new_n252), .A3(new_n247), .ZN(new_n253));
  AOI21_X1  g052(.A(new_n252), .B1(new_n246), .B2(new_n247), .ZN(new_n254));
  NOR3_X1   g053(.A1(new_n253), .A2(new_n254), .A3(new_n235), .ZN(new_n255));
  OAI21_X1  g054(.A(new_n251), .B1(new_n255), .B2(new_n243), .ZN(new_n256));
  INV_X1    g055(.A(new_n256), .ZN(new_n257));
  INV_X1    g056(.A(KEYINPUT25), .ZN(new_n258));
  NOR2_X1   g057(.A1(G169gat), .A2(G176gat), .ZN(new_n259));
  AOI21_X1  g058(.A(new_n258), .B1(new_n259), .B2(KEYINPUT23), .ZN(new_n260));
  INV_X1    g059(.A(KEYINPUT66), .ZN(new_n261));
  NAND3_X1  g060(.A1(new_n261), .A2(G169gat), .A3(G176gat), .ZN(new_n262));
  INV_X1    g061(.A(KEYINPUT23), .ZN(new_n263));
  OAI21_X1  g062(.A(new_n263), .B1(G169gat), .B2(G176gat), .ZN(new_n264));
  NAND2_X1  g063(.A1(G169gat), .A2(G176gat), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n265), .A2(KEYINPUT66), .ZN(new_n266));
  NAND4_X1  g065(.A1(new_n260), .A2(new_n262), .A3(new_n264), .A4(new_n266), .ZN(new_n267));
  NAND2_X1  g066(.A1(G183gat), .A2(G190gat), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n268), .A2(KEYINPUT24), .ZN(new_n269));
  INV_X1    g068(.A(KEYINPUT24), .ZN(new_n270));
  NAND3_X1  g069(.A1(new_n270), .A2(G183gat), .A3(G190gat), .ZN(new_n271));
  INV_X1    g070(.A(G183gat), .ZN(new_n272));
  INV_X1    g071(.A(G190gat), .ZN(new_n273));
  AOI22_X1  g072(.A1(new_n269), .A2(new_n271), .B1(new_n272), .B2(new_n273), .ZN(new_n274));
  OAI21_X1  g073(.A(KEYINPUT67), .B1(new_n267), .B2(new_n274), .ZN(new_n275));
  OAI21_X1  g074(.A(KEYINPUT65), .B1(G183gat), .B2(G190gat), .ZN(new_n276));
  INV_X1    g075(.A(KEYINPUT65), .ZN(new_n277));
  NAND3_X1  g076(.A1(new_n277), .A2(new_n272), .A3(new_n273), .ZN(new_n278));
  AOI22_X1  g077(.A1(new_n276), .A2(new_n278), .B1(new_n269), .B2(new_n271), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n259), .A2(KEYINPUT23), .ZN(new_n280));
  NAND3_X1  g079(.A1(new_n280), .A2(new_n264), .A3(new_n265), .ZN(new_n281));
  OAI21_X1  g080(.A(new_n258), .B1(new_n279), .B2(new_n281), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n269), .A2(new_n271), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n272), .A2(new_n273), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  AND3_X1   g084(.A1(new_n266), .A2(new_n264), .A3(new_n262), .ZN(new_n286));
  INV_X1    g085(.A(KEYINPUT67), .ZN(new_n287));
  NAND4_X1  g086(.A1(new_n285), .A2(new_n286), .A3(new_n287), .A4(new_n260), .ZN(new_n288));
  NAND3_X1  g087(.A1(new_n275), .A2(new_n282), .A3(new_n288), .ZN(new_n289));
  NOR3_X1   g088(.A1(KEYINPUT26), .A2(G169gat), .A3(G176gat), .ZN(new_n290));
  INV_X1    g089(.A(KEYINPUT26), .ZN(new_n291));
  OAI21_X1  g090(.A(new_n265), .B1(new_n259), .B2(new_n291), .ZN(new_n292));
  XNOR2_X1  g091(.A(KEYINPUT27), .B(G183gat), .ZN(new_n293));
  AND3_X1   g092(.A1(new_n293), .A2(KEYINPUT28), .A3(new_n273), .ZN(new_n294));
  AOI21_X1  g093(.A(KEYINPUT28), .B1(new_n293), .B2(new_n273), .ZN(new_n295));
  OAI221_X1 g094(.A(new_n268), .B1(new_n290), .B2(new_n292), .C1(new_n294), .C2(new_n295), .ZN(new_n296));
  NAND2_X1  g095(.A1(new_n289), .A2(new_n296), .ZN(new_n297));
  INV_X1    g096(.A(KEYINPUT70), .ZN(new_n298));
  NAND2_X1  g097(.A1(G127gat), .A2(G134gat), .ZN(new_n299));
  INV_X1    g098(.A(new_n299), .ZN(new_n300));
  NOR2_X1   g099(.A1(G127gat), .A2(G134gat), .ZN(new_n301));
  OAI21_X1  g100(.A(new_n298), .B1(new_n300), .B2(new_n301), .ZN(new_n302));
  INV_X1    g101(.A(KEYINPUT1), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  NOR3_X1   g103(.A1(new_n300), .A2(new_n301), .A3(new_n298), .ZN(new_n305));
  NOR2_X1   g104(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  INV_X1    g105(.A(G120gat), .ZN(new_n307));
  NOR2_X1   g106(.A1(new_n307), .A2(G113gat), .ZN(new_n308));
  INV_X1    g107(.A(new_n308), .ZN(new_n309));
  XOR2_X1   g108(.A(KEYINPUT69), .B(G120gat), .Z(new_n310));
  INV_X1    g109(.A(G113gat), .ZN(new_n311));
  OAI21_X1  g110(.A(new_n309), .B1(new_n310), .B2(new_n311), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n307), .A2(G113gat), .ZN(new_n313));
  NAND3_X1  g112(.A1(new_n309), .A2(new_n313), .A3(KEYINPUT68), .ZN(new_n314));
  INV_X1    g113(.A(KEYINPUT68), .ZN(new_n315));
  NOR2_X1   g114(.A1(new_n311), .A2(G120gat), .ZN(new_n316));
  OAI21_X1  g115(.A(new_n315), .B1(new_n308), .B2(new_n316), .ZN(new_n317));
  NAND3_X1  g116(.A1(new_n314), .A2(new_n317), .A3(new_n303), .ZN(new_n318));
  NOR2_X1   g117(.A1(new_n300), .A2(new_n301), .ZN(new_n319));
  AOI22_X1  g118(.A1(new_n306), .A2(new_n312), .B1(new_n318), .B2(new_n319), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n297), .A2(new_n320), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n306), .A2(new_n312), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n318), .A2(new_n319), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  NAND3_X1  g123(.A1(new_n324), .A2(new_n296), .A3(new_n289), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n321), .A2(new_n325), .ZN(new_n326));
  INV_X1    g125(.A(KEYINPUT34), .ZN(new_n327));
  NAND2_X1  g126(.A1(G227gat), .A2(G233gat), .ZN(new_n328));
  XOR2_X1   g127(.A(new_n328), .B(KEYINPUT64), .Z(new_n329));
  INV_X1    g128(.A(new_n329), .ZN(new_n330));
  NAND3_X1  g129(.A1(new_n326), .A2(new_n327), .A3(new_n330), .ZN(new_n331));
  INV_X1    g130(.A(new_n331), .ZN(new_n332));
  XOR2_X1   g131(.A(G15gat), .B(G43gat), .Z(new_n333));
  XNOR2_X1  g132(.A(G71gat), .B(G99gat), .ZN(new_n334));
  XNOR2_X1  g133(.A(new_n333), .B(new_n334), .ZN(new_n335));
  INV_X1    g134(.A(new_n335), .ZN(new_n336));
  NAND3_X1  g135(.A1(new_n321), .A2(new_n329), .A3(new_n325), .ZN(new_n337));
  INV_X1    g136(.A(KEYINPUT33), .ZN(new_n338));
  AOI21_X1  g137(.A(new_n336), .B1(new_n337), .B2(new_n338), .ZN(new_n339));
  AOI21_X1  g138(.A(new_n327), .B1(new_n326), .B2(new_n330), .ZN(new_n340));
  OR3_X1    g139(.A1(new_n332), .A2(new_n339), .A3(new_n340), .ZN(new_n341));
  AND2_X1   g140(.A1(new_n337), .A2(KEYINPUT32), .ZN(new_n342));
  OAI21_X1  g141(.A(new_n339), .B1(new_n332), .B2(new_n340), .ZN(new_n343));
  AND3_X1   g142(.A1(new_n341), .A2(new_n342), .A3(new_n343), .ZN(new_n344));
  AOI21_X1  g143(.A(new_n342), .B1(new_n341), .B2(new_n343), .ZN(new_n345));
  NOR2_X1   g144(.A1(new_n344), .A2(new_n345), .ZN(new_n346));
  INV_X1    g145(.A(KEYINPUT71), .ZN(new_n347));
  INV_X1    g146(.A(KEYINPUT36), .ZN(new_n348));
  NAND3_X1  g147(.A1(new_n346), .A2(new_n347), .A3(new_n348), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n347), .A2(new_n348), .ZN(new_n350));
  NAND2_X1  g149(.A1(KEYINPUT71), .A2(KEYINPUT36), .ZN(new_n351));
  OAI211_X1 g150(.A(new_n350), .B(new_n351), .C1(new_n344), .C2(new_n345), .ZN(new_n352));
  XNOR2_X1  g151(.A(G78gat), .B(G106gat), .ZN(new_n353));
  XNOR2_X1  g152(.A(new_n353), .B(new_n216), .ZN(new_n354));
  XNOR2_X1  g153(.A(new_n354), .B(G22gat), .ZN(new_n355));
  INV_X1    g154(.A(new_n355), .ZN(new_n356));
  NAND2_X1  g155(.A1(G228gat), .A2(G233gat), .ZN(new_n357));
  INV_X1    g156(.A(new_n357), .ZN(new_n358));
  NAND2_X1  g157(.A1(G155gat), .A2(G162gat), .ZN(new_n359));
  INV_X1    g158(.A(G155gat), .ZN(new_n360));
  INV_X1    g159(.A(G162gat), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  OAI21_X1  g161(.A(new_n359), .B1(new_n362), .B2(KEYINPUT2), .ZN(new_n363));
  AND2_X1   g162(.A1(G141gat), .A2(G148gat), .ZN(new_n364));
  NOR2_X1   g163(.A1(G141gat), .A2(G148gat), .ZN(new_n365));
  NOR2_X1   g164(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n363), .A2(new_n366), .ZN(new_n367));
  INV_X1    g166(.A(KEYINPUT77), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  NAND3_X1  g168(.A1(new_n363), .A2(new_n366), .A3(KEYINPUT77), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n369), .A2(new_n370), .ZN(new_n371));
  OAI21_X1  g170(.A(KEYINPUT75), .B1(new_n364), .B2(new_n365), .ZN(new_n372));
  INV_X1    g171(.A(G141gat), .ZN(new_n373));
  INV_X1    g172(.A(G148gat), .ZN(new_n374));
  NAND2_X1  g173(.A1(new_n373), .A2(new_n374), .ZN(new_n375));
  INV_X1    g174(.A(KEYINPUT75), .ZN(new_n376));
  NAND2_X1  g175(.A1(G141gat), .A2(G148gat), .ZN(new_n377));
  NAND3_X1  g176(.A1(new_n375), .A2(new_n376), .A3(new_n377), .ZN(new_n378));
  INV_X1    g177(.A(KEYINPUT2), .ZN(new_n379));
  NAND3_X1  g178(.A1(new_n372), .A2(new_n378), .A3(new_n379), .ZN(new_n380));
  INV_X1    g179(.A(KEYINPUT76), .ZN(new_n381));
  AND2_X1   g180(.A1(new_n362), .A2(new_n359), .ZN(new_n382));
  AND3_X1   g181(.A1(new_n380), .A2(new_n381), .A3(new_n382), .ZN(new_n383));
  AOI21_X1  g182(.A(new_n381), .B1(new_n380), .B2(new_n382), .ZN(new_n384));
  OAI21_X1  g183(.A(new_n371), .B1(new_n383), .B2(new_n384), .ZN(new_n385));
  INV_X1    g184(.A(new_n385), .ZN(new_n386));
  INV_X1    g185(.A(G211gat), .ZN(new_n387));
  INV_X1    g186(.A(G218gat), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n387), .A2(new_n388), .ZN(new_n389));
  NAND2_X1  g188(.A1(G211gat), .A2(G218gat), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n389), .A2(new_n390), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n391), .A2(KEYINPUT72), .ZN(new_n392));
  INV_X1    g191(.A(KEYINPUT72), .ZN(new_n393));
  NAND3_X1  g192(.A1(new_n389), .A2(new_n393), .A3(new_n390), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n392), .A2(new_n394), .ZN(new_n395));
  XNOR2_X1  g194(.A(G197gat), .B(G204gat), .ZN(new_n396));
  INV_X1    g195(.A(KEYINPUT22), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n390), .A2(new_n397), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n396), .A2(new_n398), .ZN(new_n399));
  INV_X1    g198(.A(new_n399), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n395), .A2(new_n400), .ZN(new_n401));
  NAND3_X1  g200(.A1(new_n392), .A2(new_n399), .A3(new_n394), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n401), .A2(new_n402), .ZN(new_n403));
  INV_X1    g202(.A(KEYINPUT29), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n403), .A2(new_n404), .ZN(new_n405));
  INV_X1    g204(.A(KEYINPUT82), .ZN(new_n406));
  AOI21_X1  g205(.A(KEYINPUT3), .B1(new_n405), .B2(new_n406), .ZN(new_n407));
  NAND3_X1  g206(.A1(new_n403), .A2(KEYINPUT82), .A3(new_n404), .ZN(new_n408));
  AOI21_X1  g207(.A(new_n386), .B1(new_n407), .B2(new_n408), .ZN(new_n409));
  INV_X1    g208(.A(KEYINPUT3), .ZN(new_n410));
  OAI211_X1 g209(.A(new_n371), .B(new_n410), .C1(new_n383), .C2(new_n384), .ZN(new_n411));
  AOI21_X1  g210(.A(new_n403), .B1(new_n411), .B2(new_n404), .ZN(new_n412));
  OAI21_X1  g211(.A(new_n358), .B1(new_n409), .B2(new_n412), .ZN(new_n413));
  NOR2_X1   g212(.A1(new_n403), .A2(KEYINPUT81), .ZN(new_n414));
  INV_X1    g213(.A(KEYINPUT81), .ZN(new_n415));
  OAI21_X1  g214(.A(new_n404), .B1(new_n401), .B2(new_n415), .ZN(new_n416));
  OAI21_X1  g215(.A(new_n410), .B1(new_n414), .B2(new_n416), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n417), .A2(new_n385), .ZN(new_n418));
  INV_X1    g217(.A(new_n412), .ZN(new_n419));
  NAND3_X1  g218(.A1(new_n418), .A2(new_n357), .A3(new_n419), .ZN(new_n420));
  XNOR2_X1  g219(.A(KEYINPUT80), .B(KEYINPUT31), .ZN(new_n421));
  INV_X1    g220(.A(new_n421), .ZN(new_n422));
  AND3_X1   g221(.A1(new_n413), .A2(new_n420), .A3(new_n422), .ZN(new_n423));
  AOI21_X1  g222(.A(new_n422), .B1(new_n413), .B2(new_n420), .ZN(new_n424));
  OAI21_X1  g223(.A(new_n356), .B1(new_n423), .B2(new_n424), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n413), .A2(new_n420), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n426), .A2(new_n421), .ZN(new_n427));
  NAND3_X1  g226(.A1(new_n413), .A2(new_n420), .A3(new_n422), .ZN(new_n428));
  NAND3_X1  g227(.A1(new_n427), .A2(new_n428), .A3(new_n355), .ZN(new_n429));
  AND2_X1   g228(.A1(new_n425), .A2(new_n429), .ZN(new_n430));
  NAND2_X1  g229(.A1(G225gat), .A2(G233gat), .ZN(new_n431));
  INV_X1    g230(.A(new_n431), .ZN(new_n432));
  NOR2_X1   g231(.A1(new_n385), .A2(new_n324), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n380), .A2(new_n382), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n434), .A2(KEYINPUT76), .ZN(new_n435));
  NAND3_X1  g234(.A1(new_n380), .A2(new_n381), .A3(new_n382), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n435), .A2(new_n436), .ZN(new_n437));
  AOI21_X1  g236(.A(new_n320), .B1(new_n437), .B2(new_n371), .ZN(new_n438));
  OAI21_X1  g237(.A(new_n432), .B1(new_n433), .B2(new_n438), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n439), .A2(KEYINPUT5), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n385), .A2(KEYINPUT3), .ZN(new_n441));
  NAND3_X1  g240(.A1(new_n441), .A2(new_n411), .A3(new_n324), .ZN(new_n442));
  INV_X1    g241(.A(KEYINPUT4), .ZN(new_n443));
  OAI21_X1  g242(.A(new_n443), .B1(new_n385), .B2(new_n324), .ZN(new_n444));
  NAND4_X1  g243(.A1(new_n437), .A2(new_n320), .A3(KEYINPUT4), .A4(new_n371), .ZN(new_n445));
  NAND4_X1  g244(.A1(new_n442), .A2(new_n431), .A3(new_n444), .A4(new_n445), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n440), .A2(new_n446), .ZN(new_n447));
  AND2_X1   g246(.A1(new_n444), .A2(new_n445), .ZN(new_n448));
  NAND4_X1  g247(.A1(new_n448), .A2(KEYINPUT5), .A3(new_n431), .A4(new_n442), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n447), .A2(new_n449), .ZN(new_n450));
  XOR2_X1   g249(.A(G1gat), .B(G29gat), .Z(new_n451));
  XNOR2_X1  g250(.A(KEYINPUT78), .B(KEYINPUT0), .ZN(new_n452));
  XNOR2_X1  g251(.A(new_n451), .B(new_n452), .ZN(new_n453));
  XNOR2_X1  g252(.A(G57gat), .B(G85gat), .ZN(new_n454));
  XNOR2_X1  g253(.A(new_n453), .B(new_n454), .ZN(new_n455));
  OAI21_X1  g254(.A(KEYINPUT79), .B1(new_n450), .B2(new_n455), .ZN(new_n456));
  AOI21_X1  g255(.A(KEYINPUT6), .B1(new_n450), .B2(new_n455), .ZN(new_n457));
  INV_X1    g256(.A(KEYINPUT79), .ZN(new_n458));
  INV_X1    g257(.A(new_n455), .ZN(new_n459));
  NAND4_X1  g258(.A1(new_n447), .A2(new_n458), .A3(new_n449), .A4(new_n459), .ZN(new_n460));
  NAND3_X1  g259(.A1(new_n456), .A2(new_n457), .A3(new_n460), .ZN(new_n461));
  NAND4_X1  g260(.A1(new_n447), .A2(KEYINPUT6), .A3(new_n449), .A4(new_n459), .ZN(new_n462));
  NAND2_X1  g261(.A1(G226gat), .A2(G233gat), .ZN(new_n463));
  INV_X1    g262(.A(new_n463), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n297), .A2(new_n464), .ZN(new_n465));
  AOI21_X1  g264(.A(KEYINPUT29), .B1(new_n289), .B2(new_n296), .ZN(new_n466));
  OAI211_X1 g265(.A(new_n465), .B(new_n403), .C1(new_n464), .C2(new_n466), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n467), .A2(KEYINPUT74), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n297), .A2(new_n404), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n469), .A2(new_n463), .ZN(new_n470));
  INV_X1    g269(.A(KEYINPUT74), .ZN(new_n471));
  NAND4_X1  g270(.A1(new_n470), .A2(new_n471), .A3(new_n403), .A4(new_n465), .ZN(new_n472));
  AOI21_X1  g271(.A(new_n464), .B1(new_n297), .B2(new_n404), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n465), .A2(KEYINPUT73), .ZN(new_n474));
  AOI21_X1  g273(.A(new_n463), .B1(new_n289), .B2(new_n296), .ZN(new_n475));
  INV_X1    g274(.A(KEYINPUT73), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  AOI21_X1  g276(.A(new_n473), .B1(new_n474), .B2(new_n477), .ZN(new_n478));
  OAI211_X1 g277(.A(new_n468), .B(new_n472), .C1(new_n478), .C2(new_n403), .ZN(new_n479));
  XNOR2_X1  g278(.A(G8gat), .B(G36gat), .ZN(new_n480));
  XNOR2_X1  g279(.A(G64gat), .B(G92gat), .ZN(new_n481));
  XOR2_X1   g280(.A(new_n480), .B(new_n481), .Z(new_n482));
  INV_X1    g281(.A(new_n482), .ZN(new_n483));
  OR3_X1    g282(.A1(new_n479), .A2(KEYINPUT30), .A3(new_n483), .ZN(new_n484));
  INV_X1    g283(.A(new_n403), .ZN(new_n485));
  NOR2_X1   g284(.A1(new_n475), .A2(new_n476), .ZN(new_n486));
  AOI211_X1 g285(.A(KEYINPUT73), .B(new_n463), .C1(new_n289), .C2(new_n296), .ZN(new_n487));
  OAI21_X1  g286(.A(new_n470), .B1(new_n486), .B2(new_n487), .ZN(new_n488));
  NOR3_X1   g287(.A1(new_n473), .A2(new_n485), .A3(new_n475), .ZN(new_n489));
  AOI22_X1  g288(.A1(new_n485), .A2(new_n488), .B1(new_n489), .B2(new_n471), .ZN(new_n490));
  NAND3_X1  g289(.A1(new_n490), .A2(new_n482), .A3(new_n468), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n479), .A2(new_n483), .ZN(new_n492));
  NAND3_X1  g291(.A1(new_n491), .A2(new_n492), .A3(KEYINPUT30), .ZN(new_n493));
  AOI22_X1  g292(.A1(new_n461), .A2(new_n462), .B1(new_n484), .B2(new_n493), .ZN(new_n494));
  OAI211_X1 g293(.A(new_n349), .B(new_n352), .C1(new_n430), .C2(new_n494), .ZN(new_n495));
  INV_X1    g294(.A(new_n495), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n450), .A2(KEYINPUT84), .ZN(new_n497));
  INV_X1    g296(.A(KEYINPUT84), .ZN(new_n498));
  NAND3_X1  g297(.A1(new_n447), .A2(new_n498), .A3(new_n449), .ZN(new_n499));
  NAND3_X1  g298(.A1(new_n497), .A2(new_n459), .A3(new_n499), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n500), .A2(new_n457), .ZN(new_n501));
  OAI21_X1  g300(.A(new_n483), .B1(new_n479), .B2(KEYINPUT37), .ZN(new_n502));
  INV_X1    g301(.A(KEYINPUT37), .ZN(new_n503));
  AOI21_X1  g302(.A(new_n503), .B1(new_n490), .B2(new_n468), .ZN(new_n504));
  OAI21_X1  g303(.A(KEYINPUT38), .B1(new_n502), .B2(new_n504), .ZN(new_n505));
  NAND4_X1  g304(.A1(new_n501), .A2(new_n462), .A3(new_n505), .A4(new_n491), .ZN(new_n506));
  NAND2_X1  g305(.A1(new_n483), .A2(KEYINPUT37), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n492), .A2(new_n507), .ZN(new_n508));
  INV_X1    g307(.A(KEYINPUT38), .ZN(new_n509));
  OAI211_X1 g308(.A(new_n470), .B(new_n403), .C1(new_n486), .C2(new_n487), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n510), .A2(KEYINPUT85), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n474), .A2(new_n477), .ZN(new_n512));
  INV_X1    g311(.A(KEYINPUT85), .ZN(new_n513));
  NAND4_X1  g312(.A1(new_n512), .A2(new_n513), .A3(new_n403), .A4(new_n470), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n470), .A2(new_n465), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n515), .A2(new_n485), .ZN(new_n516));
  NAND3_X1  g315(.A1(new_n511), .A2(new_n514), .A3(new_n516), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n517), .A2(KEYINPUT37), .ZN(new_n518));
  NAND4_X1  g317(.A1(new_n508), .A2(KEYINPUT86), .A3(new_n509), .A4(new_n518), .ZN(new_n519));
  INV_X1    g318(.A(KEYINPUT86), .ZN(new_n520));
  OAI211_X1 g319(.A(new_n509), .B(new_n483), .C1(new_n479), .C2(KEYINPUT37), .ZN(new_n521));
  AOI22_X1  g320(.A1(new_n510), .A2(KEYINPUT85), .B1(new_n485), .B2(new_n515), .ZN(new_n522));
  AOI21_X1  g321(.A(new_n503), .B1(new_n522), .B2(new_n514), .ZN(new_n523));
  OAI21_X1  g322(.A(new_n520), .B1(new_n521), .B2(new_n523), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n519), .A2(new_n524), .ZN(new_n525));
  NOR2_X1   g324(.A1(new_n506), .A2(new_n525), .ZN(new_n526));
  INV_X1    g325(.A(KEYINPUT87), .ZN(new_n527));
  INV_X1    g326(.A(KEYINPUT40), .ZN(new_n528));
  OR3_X1    g327(.A1(new_n433), .A2(new_n438), .A3(new_n432), .ZN(new_n529));
  NAND2_X1  g328(.A1(new_n529), .A2(KEYINPUT39), .ZN(new_n530));
  NAND2_X1  g329(.A1(new_n448), .A2(new_n442), .ZN(new_n531));
  AOI21_X1  g330(.A(new_n530), .B1(new_n432), .B2(new_n531), .ZN(new_n532));
  XOR2_X1   g331(.A(KEYINPUT83), .B(KEYINPUT39), .Z(new_n533));
  NAND3_X1  g332(.A1(new_n531), .A2(new_n432), .A3(new_n533), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n534), .A2(new_n455), .ZN(new_n535));
  OAI21_X1  g334(.A(new_n528), .B1(new_n532), .B2(new_n535), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n531), .A2(new_n432), .ZN(new_n537));
  NAND3_X1  g336(.A1(new_n537), .A2(KEYINPUT39), .A3(new_n529), .ZN(new_n538));
  NAND4_X1  g337(.A1(new_n538), .A2(KEYINPUT40), .A3(new_n455), .A4(new_n534), .ZN(new_n539));
  NAND3_X1  g338(.A1(new_n500), .A2(new_n536), .A3(new_n539), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n493), .A2(new_n484), .ZN(new_n541));
  OAI21_X1  g340(.A(new_n430), .B1(new_n540), .B2(new_n541), .ZN(new_n542));
  NOR3_X1   g341(.A1(new_n526), .A2(new_n527), .A3(new_n542), .ZN(new_n543));
  AND2_X1   g342(.A1(new_n519), .A2(new_n524), .ZN(new_n544));
  INV_X1    g343(.A(new_n462), .ZN(new_n545));
  INV_X1    g344(.A(new_n491), .ZN(new_n546));
  AOI211_X1 g345(.A(new_n545), .B(new_n546), .C1(new_n500), .C2(new_n457), .ZN(new_n547));
  NAND3_X1  g346(.A1(new_n544), .A2(new_n547), .A3(new_n505), .ZN(new_n548));
  INV_X1    g347(.A(new_n542), .ZN(new_n549));
  AOI21_X1  g348(.A(KEYINPUT87), .B1(new_n548), .B2(new_n549), .ZN(new_n550));
  OAI21_X1  g349(.A(new_n496), .B1(new_n543), .B2(new_n550), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n425), .A2(new_n429), .ZN(new_n552));
  NOR3_X1   g351(.A1(new_n552), .A2(new_n344), .A3(new_n345), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n553), .A2(new_n494), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n554), .A2(KEYINPUT35), .ZN(new_n555));
  AOI21_X1  g354(.A(new_n545), .B1(new_n500), .B2(new_n457), .ZN(new_n556));
  NOR2_X1   g355(.A1(new_n556), .A2(KEYINPUT35), .ZN(new_n557));
  NAND3_X1  g356(.A1(new_n557), .A2(new_n541), .A3(new_n553), .ZN(new_n558));
  NAND2_X1  g357(.A1(new_n555), .A2(new_n558), .ZN(new_n559));
  AOI21_X1  g358(.A(new_n257), .B1(new_n551), .B2(new_n559), .ZN(new_n560));
  NAND2_X1  g359(.A1(G71gat), .A2(G78gat), .ZN(new_n561));
  INV_X1    g360(.A(KEYINPUT91), .ZN(new_n562));
  NAND2_X1  g361(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  OR2_X1    g362(.A1(G71gat), .A2(G78gat), .ZN(new_n564));
  NAND3_X1  g363(.A1(KEYINPUT91), .A2(G71gat), .A3(G78gat), .ZN(new_n565));
  NAND3_X1  g364(.A1(new_n563), .A2(new_n564), .A3(new_n565), .ZN(new_n566));
  INV_X1    g365(.A(KEYINPUT92), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  NAND4_X1  g367(.A1(new_n563), .A2(new_n564), .A3(KEYINPUT92), .A4(new_n565), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  XOR2_X1   g369(.A(G57gat), .B(G64gat), .Z(new_n571));
  INV_X1    g370(.A(KEYINPUT9), .ZN(new_n572));
  NAND2_X1  g371(.A1(new_n561), .A2(new_n572), .ZN(new_n573));
  NAND2_X1  g372(.A1(new_n571), .A2(new_n573), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n570), .A2(new_n574), .ZN(new_n575));
  INV_X1    g374(.A(KEYINPUT93), .ZN(new_n576));
  NAND4_X1  g375(.A1(new_n571), .A2(KEYINPUT9), .A3(new_n561), .A4(new_n564), .ZN(new_n577));
  NAND3_X1  g376(.A1(new_n575), .A2(new_n576), .A3(new_n577), .ZN(new_n578));
  AOI22_X1  g377(.A1(new_n568), .A2(new_n569), .B1(new_n573), .B2(new_n571), .ZN(new_n579));
  INV_X1    g378(.A(new_n577), .ZN(new_n580));
  OAI21_X1  g379(.A(KEYINPUT93), .B1(new_n579), .B2(new_n580), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n578), .A2(new_n581), .ZN(new_n582));
  INV_X1    g381(.A(G231gat), .ZN(new_n583));
  INV_X1    g382(.A(G233gat), .ZN(new_n584));
  NOR2_X1   g383(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  OR3_X1    g384(.A1(new_n582), .A2(KEYINPUT21), .A3(new_n585), .ZN(new_n586));
  INV_X1    g385(.A(G127gat), .ZN(new_n587));
  OAI21_X1  g386(.A(new_n585), .B1(new_n582), .B2(KEYINPUT21), .ZN(new_n588));
  AND3_X1   g387(.A1(new_n586), .A2(new_n587), .A3(new_n588), .ZN(new_n589));
  AOI21_X1  g388(.A(new_n587), .B1(new_n586), .B2(new_n588), .ZN(new_n590));
  OR2_X1    g389(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  XOR2_X1   g390(.A(G183gat), .B(G211gat), .Z(new_n592));
  OR2_X1    g391(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  OAI21_X1  g392(.A(new_n592), .B1(new_n589), .B2(new_n590), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  AOI21_X1  g394(.A(new_n207), .B1(new_n582), .B2(KEYINPUT21), .ZN(new_n596));
  XNOR2_X1  g395(.A(new_n596), .B(KEYINPUT94), .ZN(new_n597));
  XNOR2_X1  g396(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n598));
  XNOR2_X1  g397(.A(new_n598), .B(new_n360), .ZN(new_n599));
  XNOR2_X1  g398(.A(new_n597), .B(new_n599), .ZN(new_n600));
  INV_X1    g399(.A(new_n600), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n595), .A2(new_n601), .ZN(new_n602));
  NAND3_X1  g401(.A1(new_n593), .A2(new_n594), .A3(new_n600), .ZN(new_n603));
  INV_X1    g402(.A(KEYINPUT97), .ZN(new_n604));
  NAND2_X1  g403(.A1(new_n604), .A2(KEYINPUT7), .ZN(new_n605));
  INV_X1    g404(.A(KEYINPUT7), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n606), .A2(KEYINPUT97), .ZN(new_n607));
  NAND4_X1  g406(.A1(new_n605), .A2(new_n607), .A3(G85gat), .A4(G92gat), .ZN(new_n608));
  INV_X1    g407(.A(G85gat), .ZN(new_n609));
  INV_X1    g408(.A(G92gat), .ZN(new_n610));
  OAI211_X1 g409(.A(KEYINPUT97), .B(new_n606), .C1(new_n609), .C2(new_n610), .ZN(new_n611));
  NAND2_X1  g410(.A1(G99gat), .A2(G106gat), .ZN(new_n612));
  AOI22_X1  g411(.A1(KEYINPUT8), .A2(new_n612), .B1(new_n609), .B2(new_n610), .ZN(new_n613));
  NAND3_X1  g412(.A1(new_n608), .A2(new_n611), .A3(new_n613), .ZN(new_n614));
  OR2_X1    g413(.A1(G99gat), .A2(G106gat), .ZN(new_n615));
  NAND3_X1  g414(.A1(new_n614), .A2(new_n612), .A3(new_n615), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n615), .A2(new_n612), .ZN(new_n617));
  NAND4_X1  g416(.A1(new_n608), .A2(new_n617), .A3(new_n611), .A4(new_n613), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n616), .A2(new_n618), .ZN(new_n619));
  INV_X1    g418(.A(new_n619), .ZN(new_n620));
  AND2_X1   g419(.A1(G232gat), .A2(G233gat), .ZN(new_n621));
  AOI22_X1  g420(.A1(new_n229), .A2(new_n620), .B1(KEYINPUT41), .B2(new_n621), .ZN(new_n622));
  NAND3_X1  g421(.A1(new_n224), .A2(new_n227), .A3(new_n619), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  XNOR2_X1  g423(.A(G190gat), .B(G218gat), .ZN(new_n625));
  XNOR2_X1  g424(.A(KEYINPUT98), .B(KEYINPUT99), .ZN(new_n626));
  XOR2_X1   g425(.A(new_n625), .B(new_n626), .Z(new_n627));
  XNOR2_X1  g426(.A(new_n624), .B(new_n627), .ZN(new_n628));
  XOR2_X1   g427(.A(G134gat), .B(G162gat), .Z(new_n629));
  NOR2_X1   g428(.A1(new_n621), .A2(KEYINPUT41), .ZN(new_n630));
  XNOR2_X1  g429(.A(new_n629), .B(new_n630), .ZN(new_n631));
  XOR2_X1   g430(.A(KEYINPUT95), .B(KEYINPUT96), .Z(new_n632));
  XNOR2_X1  g431(.A(new_n631), .B(new_n632), .ZN(new_n633));
  INV_X1    g432(.A(new_n633), .ZN(new_n634));
  OR2_X1    g433(.A1(new_n628), .A2(new_n634), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n628), .A2(new_n634), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  NAND3_X1  g436(.A1(new_n602), .A2(new_n603), .A3(new_n637), .ZN(new_n638));
  NAND2_X1  g437(.A1(new_n638), .A2(KEYINPUT100), .ZN(new_n639));
  INV_X1    g438(.A(KEYINPUT100), .ZN(new_n640));
  NAND4_X1  g439(.A1(new_n602), .A2(new_n603), .A3(new_n640), .A4(new_n637), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n639), .A2(new_n641), .ZN(new_n642));
  NAND3_X1  g441(.A1(new_n582), .A2(KEYINPUT10), .A3(new_n620), .ZN(new_n643));
  NOR3_X1   g442(.A1(new_n619), .A2(new_n579), .A3(new_n580), .ZN(new_n644));
  AOI21_X1  g443(.A(new_n644), .B1(new_n582), .B2(new_n619), .ZN(new_n645));
  OAI21_X1  g444(.A(new_n643), .B1(new_n645), .B2(KEYINPUT10), .ZN(new_n646));
  NAND2_X1  g445(.A1(G230gat), .A2(G233gat), .ZN(new_n647));
  NAND2_X1  g446(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  NAND2_X1  g447(.A1(new_n648), .A2(KEYINPUT101), .ZN(new_n649));
  INV_X1    g448(.A(KEYINPUT101), .ZN(new_n650));
  NAND3_X1  g449(.A1(new_n646), .A2(new_n650), .A3(new_n647), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n649), .A2(new_n651), .ZN(new_n652));
  INV_X1    g451(.A(new_n647), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n645), .A2(new_n653), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n652), .A2(new_n654), .ZN(new_n655));
  XNOR2_X1  g454(.A(G120gat), .B(G148gat), .ZN(new_n656));
  XNOR2_X1  g455(.A(G176gat), .B(G204gat), .ZN(new_n657));
  XOR2_X1   g456(.A(new_n656), .B(new_n657), .Z(new_n658));
  INV_X1    g457(.A(new_n658), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n655), .A2(new_n659), .ZN(new_n660));
  NAND3_X1  g459(.A1(new_n648), .A2(new_n654), .A3(new_n658), .ZN(new_n661));
  NAND2_X1  g460(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  NOR2_X1   g461(.A1(new_n642), .A2(new_n662), .ZN(new_n663));
  NAND2_X1  g462(.A1(new_n560), .A2(new_n663), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n461), .A2(new_n462), .ZN(new_n665));
  NOR2_X1   g464(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  XNOR2_X1  g465(.A(new_n666), .B(new_n203), .ZN(G1324gat));
  INV_X1    g466(.A(new_n664), .ZN(new_n668));
  INV_X1    g467(.A(new_n541), .ZN(new_n669));
  XOR2_X1   g468(.A(KEYINPUT16), .B(G8gat), .Z(new_n670));
  AND3_X1   g469(.A1(new_n668), .A2(new_n669), .A3(new_n670), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n668), .A2(new_n669), .ZN(new_n672));
  AOI22_X1  g471(.A1(new_n671), .A2(KEYINPUT42), .B1(G8gat), .B2(new_n672), .ZN(new_n673));
  NOR2_X1   g472(.A1(new_n671), .A2(KEYINPUT42), .ZN(new_n674));
  AND2_X1   g473(.A1(new_n674), .A2(KEYINPUT102), .ZN(new_n675));
  NOR2_X1   g474(.A1(new_n674), .A2(KEYINPUT102), .ZN(new_n676));
  OAI21_X1  g475(.A(new_n673), .B1(new_n675), .B2(new_n676), .ZN(G1325gat));
  NAND2_X1  g476(.A1(new_n349), .A2(new_n352), .ZN(new_n678));
  INV_X1    g477(.A(new_n678), .ZN(new_n679));
  OAI21_X1  g478(.A(G15gat), .B1(new_n664), .B2(new_n679), .ZN(new_n680));
  INV_X1    g479(.A(new_n346), .ZN(new_n681));
  OR2_X1    g480(.A1(new_n681), .A2(G15gat), .ZN(new_n682));
  OAI21_X1  g481(.A(new_n680), .B1(new_n664), .B2(new_n682), .ZN(G1326gat));
  NAND2_X1  g482(.A1(new_n560), .A2(new_n552), .ZN(new_n684));
  NOR3_X1   g483(.A1(new_n684), .A2(new_n642), .A3(new_n662), .ZN(new_n685));
  XNOR2_X1  g484(.A(new_n685), .B(KEYINPUT103), .ZN(new_n686));
  XNOR2_X1  g485(.A(KEYINPUT43), .B(G22gat), .ZN(new_n687));
  XNOR2_X1  g486(.A(new_n686), .B(new_n687), .ZN(G1327gat));
  NAND2_X1  g487(.A1(new_n551), .A2(KEYINPUT105), .ZN(new_n689));
  OAI21_X1  g488(.A(new_n527), .B1(new_n526), .B2(new_n542), .ZN(new_n690));
  NAND3_X1  g489(.A1(new_n548), .A2(KEYINPUT87), .A3(new_n549), .ZN(new_n691));
  AOI21_X1  g490(.A(new_n495), .B1(new_n690), .B2(new_n691), .ZN(new_n692));
  INV_X1    g491(.A(KEYINPUT105), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  INV_X1    g493(.A(KEYINPUT106), .ZN(new_n695));
  NAND3_X1  g494(.A1(new_n346), .A2(new_n430), .A3(new_n541), .ZN(new_n696));
  NOR3_X1   g495(.A1(new_n696), .A2(KEYINPUT35), .A3(new_n556), .ZN(new_n697));
  INV_X1    g496(.A(KEYINPUT35), .ZN(new_n698));
  AOI21_X1  g497(.A(new_n698), .B1(new_n553), .B2(new_n494), .ZN(new_n699));
  OAI21_X1  g498(.A(new_n695), .B1(new_n697), .B2(new_n699), .ZN(new_n700));
  NAND3_X1  g499(.A1(new_n555), .A2(KEYINPUT106), .A3(new_n558), .ZN(new_n701));
  NAND2_X1  g500(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  NAND3_X1  g501(.A1(new_n689), .A2(new_n694), .A3(new_n702), .ZN(new_n703));
  INV_X1    g502(.A(new_n637), .ZN(new_n704));
  AOI21_X1  g503(.A(KEYINPUT44), .B1(new_n703), .B2(new_n704), .ZN(new_n705));
  INV_X1    g504(.A(KEYINPUT44), .ZN(new_n706));
  AOI211_X1 g505(.A(new_n706), .B(new_n637), .C1(new_n551), .C2(new_n559), .ZN(new_n707));
  NOR2_X1   g506(.A1(new_n705), .A2(new_n707), .ZN(new_n708));
  XNOR2_X1  g507(.A(new_n662), .B(KEYINPUT104), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n602), .A2(new_n603), .ZN(new_n710));
  INV_X1    g509(.A(new_n710), .ZN(new_n711));
  NOR3_X1   g510(.A1(new_n709), .A2(new_n257), .A3(new_n711), .ZN(new_n712));
  NAND2_X1  g511(.A1(new_n708), .A2(new_n712), .ZN(new_n713));
  OAI21_X1  g512(.A(G29gat), .B1(new_n713), .B2(new_n665), .ZN(new_n714));
  INV_X1    g513(.A(KEYINPUT45), .ZN(new_n715));
  NOR3_X1   g514(.A1(new_n711), .A2(new_n637), .A3(new_n662), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n560), .A2(new_n716), .ZN(new_n717));
  NOR2_X1   g516(.A1(new_n665), .A2(G29gat), .ZN(new_n718));
  INV_X1    g517(.A(new_n718), .ZN(new_n719));
  OAI21_X1  g518(.A(new_n715), .B1(new_n717), .B2(new_n719), .ZN(new_n720));
  NAND4_X1  g519(.A1(new_n560), .A2(KEYINPUT45), .A3(new_n716), .A4(new_n718), .ZN(new_n721));
  NAND3_X1  g520(.A1(new_n714), .A2(new_n720), .A3(new_n721), .ZN(G1328gat));
  OAI21_X1  g521(.A(G36gat), .B1(new_n713), .B2(new_n541), .ZN(new_n723));
  NOR2_X1   g522(.A1(new_n541), .A2(G36gat), .ZN(new_n724));
  INV_X1    g523(.A(new_n724), .ZN(new_n725));
  OAI21_X1  g524(.A(KEYINPUT46), .B1(new_n717), .B2(new_n725), .ZN(new_n726));
  OR3_X1    g525(.A1(new_n717), .A2(KEYINPUT46), .A3(new_n725), .ZN(new_n727));
  NAND3_X1  g526(.A1(new_n723), .A2(new_n726), .A3(new_n727), .ZN(G1329gat));
  NAND4_X1  g527(.A1(new_n708), .A2(G43gat), .A3(new_n678), .A4(new_n712), .ZN(new_n729));
  OR2_X1    g528(.A1(KEYINPUT107), .A2(KEYINPUT47), .ZN(new_n730));
  NAND3_X1  g529(.A1(new_n560), .A2(new_n346), .A3(new_n716), .ZN(new_n731));
  AOI22_X1  g530(.A1(new_n731), .A2(new_n215), .B1(KEYINPUT107), .B2(KEYINPUT47), .ZN(new_n732));
  AND3_X1   g531(.A1(new_n729), .A2(new_n730), .A3(new_n732), .ZN(new_n733));
  AOI21_X1  g532(.A(new_n730), .B1(new_n729), .B2(new_n732), .ZN(new_n734));
  NOR2_X1   g533(.A1(new_n733), .A2(new_n734), .ZN(G1330gat));
  OAI21_X1  g534(.A(new_n702), .B1(new_n692), .B2(new_n693), .ZN(new_n736));
  AOI211_X1 g535(.A(KEYINPUT105), .B(new_n495), .C1(new_n690), .C2(new_n691), .ZN(new_n737));
  OAI21_X1  g536(.A(new_n704), .B1(new_n736), .B2(new_n737), .ZN(new_n738));
  NAND2_X1  g537(.A1(new_n738), .A2(new_n706), .ZN(new_n739));
  INV_X1    g538(.A(new_n707), .ZN(new_n740));
  NAND4_X1  g539(.A1(new_n739), .A2(new_n552), .A3(new_n740), .A4(new_n712), .ZN(new_n741));
  AOI21_X1  g540(.A(KEYINPUT108), .B1(new_n741), .B2(new_n221), .ZN(new_n742));
  INV_X1    g541(.A(new_n716), .ZN(new_n743));
  NOR3_X1   g542(.A1(new_n684), .A2(new_n221), .A3(new_n743), .ZN(new_n744));
  AOI21_X1  g543(.A(new_n744), .B1(new_n741), .B2(new_n221), .ZN(new_n745));
  INV_X1    g544(.A(KEYINPUT48), .ZN(new_n746));
  NOR3_X1   g545(.A1(new_n742), .A2(new_n745), .A3(new_n746), .ZN(new_n747));
  AOI221_X4 g546(.A(new_n744), .B1(KEYINPUT108), .B2(KEYINPUT48), .C1(new_n741), .C2(new_n221), .ZN(new_n748));
  NOR2_X1   g547(.A1(new_n747), .A2(new_n748), .ZN(G1331gat));
  INV_X1    g548(.A(new_n709), .ZN(new_n750));
  NOR3_X1   g549(.A1(new_n642), .A2(new_n750), .A3(new_n256), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n703), .A2(new_n751), .ZN(new_n752));
  INV_X1    g551(.A(new_n752), .ZN(new_n753));
  XNOR2_X1  g552(.A(new_n665), .B(KEYINPUT109), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  XNOR2_X1  g554(.A(new_n755), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g555(.A1(new_n753), .A2(new_n669), .ZN(new_n757));
  OAI21_X1  g556(.A(new_n757), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n758));
  XOR2_X1   g557(.A(KEYINPUT49), .B(G64gat), .Z(new_n759));
  OAI21_X1  g558(.A(new_n758), .B1(new_n757), .B2(new_n759), .ZN(G1333gat));
  OAI21_X1  g559(.A(G71gat), .B1(new_n752), .B2(new_n679), .ZN(new_n761));
  OR2_X1    g560(.A1(new_n681), .A2(G71gat), .ZN(new_n762));
  OAI21_X1  g561(.A(new_n761), .B1(new_n752), .B2(new_n762), .ZN(new_n763));
  XOR2_X1   g562(.A(new_n763), .B(KEYINPUT50), .Z(G1334gat));
  OR3_X1    g563(.A1(new_n752), .A2(KEYINPUT111), .A3(new_n430), .ZN(new_n765));
  OAI21_X1  g564(.A(KEYINPUT111), .B1(new_n752), .B2(new_n430), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  XNOR2_X1  g566(.A(KEYINPUT110), .B(G78gat), .ZN(new_n768));
  XOR2_X1   g567(.A(new_n767), .B(new_n768), .Z(G1335gat));
  NOR2_X1   g568(.A1(new_n711), .A2(new_n256), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n770), .A2(new_n662), .ZN(new_n771));
  INV_X1    g570(.A(new_n771), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n708), .A2(new_n772), .ZN(new_n773));
  OAI21_X1  g572(.A(G85gat), .B1(new_n773), .B2(new_n665), .ZN(new_n774));
  OAI211_X1 g573(.A(new_n704), .B(new_n770), .C1(new_n736), .C2(new_n737), .ZN(new_n775));
  INV_X1    g574(.A(KEYINPUT51), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  NAND4_X1  g576(.A1(new_n703), .A2(KEYINPUT51), .A3(new_n704), .A4(new_n770), .ZN(new_n778));
  NAND2_X1  g577(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  NAND2_X1  g578(.A1(new_n779), .A2(new_n662), .ZN(new_n780));
  NAND3_X1  g579(.A1(new_n461), .A2(new_n609), .A3(new_n462), .ZN(new_n781));
  OAI21_X1  g580(.A(new_n774), .B1(new_n780), .B2(new_n781), .ZN(G1336gat));
  INV_X1    g581(.A(KEYINPUT52), .ZN(new_n783));
  NAND3_X1  g582(.A1(new_n708), .A2(new_n669), .A3(new_n772), .ZN(new_n784));
  XOR2_X1   g583(.A(KEYINPUT112), .B(KEYINPUT51), .Z(new_n785));
  NAND2_X1  g584(.A1(new_n775), .A2(new_n785), .ZN(new_n786));
  NAND2_X1  g585(.A1(new_n786), .A2(new_n778), .ZN(new_n787));
  NOR3_X1   g586(.A1(new_n750), .A2(G92gat), .A3(new_n541), .ZN(new_n788));
  AOI22_X1  g587(.A1(new_n784), .A2(G92gat), .B1(new_n787), .B2(new_n788), .ZN(new_n789));
  AND2_X1   g588(.A1(new_n784), .A2(G92gat), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n779), .A2(new_n788), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n791), .A2(new_n783), .ZN(new_n792));
  OAI22_X1  g591(.A1(new_n783), .A2(new_n789), .B1(new_n790), .B2(new_n792), .ZN(G1337gat));
  OAI21_X1  g592(.A(G99gat), .B1(new_n773), .B2(new_n679), .ZN(new_n794));
  OR2_X1    g593(.A1(new_n681), .A2(G99gat), .ZN(new_n795));
  OAI21_X1  g594(.A(new_n794), .B1(new_n780), .B2(new_n795), .ZN(G1338gat));
  NOR4_X1   g595(.A1(new_n705), .A2(new_n430), .A3(new_n707), .A4(new_n771), .ZN(new_n797));
  INV_X1    g596(.A(G106gat), .ZN(new_n798));
  NOR3_X1   g597(.A1(new_n750), .A2(G106gat), .A3(new_n430), .ZN(new_n799));
  INV_X1    g598(.A(new_n799), .ZN(new_n800));
  AOI21_X1  g599(.A(new_n800), .B1(new_n786), .B2(new_n778), .ZN(new_n801));
  INV_X1    g600(.A(KEYINPUT113), .ZN(new_n802));
  OAI22_X1  g601(.A1(new_n797), .A2(new_n798), .B1(new_n801), .B2(new_n802), .ZN(new_n803));
  AND2_X1   g602(.A1(new_n801), .A2(new_n802), .ZN(new_n804));
  OAI21_X1  g603(.A(KEYINPUT53), .B1(new_n803), .B2(new_n804), .ZN(new_n805));
  AOI21_X1  g604(.A(KEYINPUT53), .B1(new_n779), .B2(new_n799), .ZN(new_n806));
  OAI21_X1  g605(.A(new_n806), .B1(new_n798), .B2(new_n797), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n805), .A2(new_n807), .ZN(G1339gat));
  INV_X1    g607(.A(new_n662), .ZN(new_n809));
  NAND4_X1  g608(.A1(new_n639), .A2(new_n257), .A3(new_n641), .A4(new_n809), .ZN(new_n810));
  INV_X1    g609(.A(KEYINPUT54), .ZN(new_n811));
  NAND3_X1  g610(.A1(new_n649), .A2(new_n811), .A3(new_n651), .ZN(new_n812));
  AOI21_X1  g611(.A(new_n811), .B1(new_n646), .B2(new_n647), .ZN(new_n813));
  OAI211_X1 g612(.A(new_n653), .B(new_n643), .C1(new_n645), .C2(KEYINPUT10), .ZN(new_n814));
  AOI21_X1  g613(.A(new_n658), .B1(new_n813), .B2(new_n814), .ZN(new_n815));
  NAND3_X1  g614(.A1(new_n812), .A2(KEYINPUT55), .A3(new_n815), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n816), .A2(new_n661), .ZN(new_n817));
  AOI21_X1  g616(.A(KEYINPUT55), .B1(new_n812), .B2(new_n815), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n228), .A2(new_n230), .ZN(new_n819));
  NAND3_X1  g618(.A1(new_n819), .A2(G229gat), .A3(G233gat), .ZN(new_n820));
  OAI21_X1  g619(.A(new_n820), .B1(new_n244), .B2(new_n245), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n821), .A2(new_n241), .ZN(new_n822));
  NAND2_X1  g621(.A1(new_n251), .A2(new_n822), .ZN(new_n823));
  NOR4_X1   g622(.A1(new_n817), .A2(new_n818), .A3(new_n637), .A4(new_n823), .ZN(new_n824));
  INV_X1    g623(.A(new_n823), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n662), .A2(new_n825), .ZN(new_n826));
  NAND3_X1  g625(.A1(new_n256), .A2(new_n816), .A3(new_n661), .ZN(new_n827));
  OAI21_X1  g626(.A(new_n826), .B1(new_n818), .B2(new_n827), .ZN(new_n828));
  AOI21_X1  g627(.A(new_n824), .B1(new_n828), .B2(new_n637), .ZN(new_n829));
  OAI21_X1  g628(.A(new_n810), .B1(new_n829), .B2(new_n711), .ZN(new_n830));
  AND2_X1   g629(.A1(new_n830), .A2(new_n754), .ZN(new_n831));
  INV_X1    g630(.A(new_n696), .ZN(new_n832));
  NAND2_X1  g631(.A1(new_n831), .A2(new_n832), .ZN(new_n833));
  INV_X1    g632(.A(new_n833), .ZN(new_n834));
  AOI21_X1  g633(.A(G113gat), .B1(new_n834), .B2(new_n256), .ZN(new_n835));
  AND2_X1   g634(.A1(new_n830), .A2(new_n430), .ZN(new_n836));
  NOR2_X1   g635(.A1(new_n665), .A2(new_n669), .ZN(new_n837));
  AND3_X1   g636(.A1(new_n836), .A2(new_n346), .A3(new_n837), .ZN(new_n838));
  NOR2_X1   g637(.A1(new_n257), .A2(new_n311), .ZN(new_n839));
  AOI21_X1  g638(.A(new_n835), .B1(new_n838), .B2(new_n839), .ZN(G1340gat));
  NOR3_X1   g639(.A1(new_n833), .A2(new_n310), .A3(new_n809), .ZN(new_n841));
  NAND2_X1  g640(.A1(new_n838), .A2(new_n709), .ZN(new_n842));
  AOI21_X1  g641(.A(new_n841), .B1(new_n842), .B2(G120gat), .ZN(new_n843));
  XOR2_X1   g642(.A(new_n843), .B(KEYINPUT114), .Z(G1341gat));
  NOR3_X1   g643(.A1(new_n833), .A2(G127gat), .A3(new_n710), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n838), .A2(new_n711), .ZN(new_n846));
  AOI21_X1  g645(.A(new_n845), .B1(new_n846), .B2(G127gat), .ZN(new_n847));
  XNOR2_X1  g646(.A(new_n847), .B(KEYINPUT115), .ZN(G1342gat));
  INV_X1    g647(.A(G134gat), .ZN(new_n849));
  NOR2_X1   g648(.A1(new_n669), .A2(new_n637), .ZN(new_n850));
  NAND4_X1  g649(.A1(new_n831), .A2(new_n849), .A3(new_n553), .A4(new_n850), .ZN(new_n851));
  XNOR2_X1  g650(.A(new_n851), .B(KEYINPUT56), .ZN(new_n852));
  AOI21_X1  g651(.A(new_n849), .B1(new_n838), .B2(new_n704), .ZN(new_n853));
  OR2_X1    g652(.A1(new_n852), .A2(new_n853), .ZN(G1343gat));
  NAND2_X1  g653(.A1(new_n679), .A2(new_n837), .ZN(new_n855));
  INV_X1    g654(.A(new_n855), .ZN(new_n856));
  INV_X1    g655(.A(KEYINPUT57), .ZN(new_n857));
  NOR2_X1   g656(.A1(new_n430), .A2(new_n857), .ZN(new_n858));
  INV_X1    g657(.A(KEYINPUT116), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n812), .A2(new_n815), .ZN(new_n860));
  INV_X1    g659(.A(KEYINPUT55), .ZN(new_n861));
  AOI21_X1  g660(.A(new_n859), .B1(new_n860), .B2(new_n861), .ZN(new_n862));
  AOI211_X1 g661(.A(KEYINPUT116), .B(KEYINPUT55), .C1(new_n812), .C2(new_n815), .ZN(new_n863));
  NOR3_X1   g662(.A1(new_n827), .A2(new_n862), .A3(new_n863), .ZN(new_n864));
  AOI21_X1  g663(.A(new_n823), .B1(new_n660), .B2(new_n661), .ZN(new_n865));
  OAI21_X1  g664(.A(new_n637), .B1(new_n864), .B2(new_n865), .ZN(new_n866));
  INV_X1    g665(.A(KEYINPUT117), .ZN(new_n867));
  AOI21_X1  g666(.A(new_n824), .B1(new_n866), .B2(new_n867), .ZN(new_n868));
  INV_X1    g667(.A(new_n862), .ZN(new_n869));
  AND3_X1   g668(.A1(new_n256), .A2(new_n816), .A3(new_n661), .ZN(new_n870));
  INV_X1    g669(.A(new_n863), .ZN(new_n871));
  NAND3_X1  g670(.A1(new_n869), .A2(new_n870), .A3(new_n871), .ZN(new_n872));
  AOI21_X1  g671(.A(new_n704), .B1(new_n872), .B2(new_n826), .ZN(new_n873));
  NAND2_X1  g672(.A1(new_n873), .A2(KEYINPUT117), .ZN(new_n874));
  AOI21_X1  g673(.A(new_n711), .B1(new_n868), .B2(new_n874), .ZN(new_n875));
  INV_X1    g674(.A(new_n810), .ZN(new_n876));
  OAI211_X1 g675(.A(KEYINPUT118), .B(new_n858), .C1(new_n875), .C2(new_n876), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n830), .A2(new_n552), .ZN(new_n878));
  NAND2_X1  g677(.A1(new_n878), .A2(new_n857), .ZN(new_n879));
  NAND2_X1  g678(.A1(new_n877), .A2(new_n879), .ZN(new_n880));
  INV_X1    g679(.A(new_n824), .ZN(new_n881));
  OAI21_X1  g680(.A(new_n881), .B1(new_n873), .B2(KEYINPUT117), .ZN(new_n882));
  NOR2_X1   g681(.A1(new_n866), .A2(new_n867), .ZN(new_n883));
  OAI21_X1  g682(.A(new_n710), .B1(new_n882), .B2(new_n883), .ZN(new_n884));
  NAND2_X1  g683(.A1(new_n884), .A2(new_n810), .ZN(new_n885));
  AOI21_X1  g684(.A(KEYINPUT118), .B1(new_n885), .B2(new_n858), .ZN(new_n886));
  OAI211_X1 g685(.A(new_n256), .B(new_n856), .C1(new_n880), .C2(new_n886), .ZN(new_n887));
  NAND2_X1  g686(.A1(new_n887), .A2(KEYINPUT121), .ZN(new_n888));
  INV_X1    g687(.A(KEYINPUT118), .ZN(new_n889));
  NAND2_X1  g688(.A1(new_n868), .A2(new_n874), .ZN(new_n890));
  AOI21_X1  g689(.A(new_n876), .B1(new_n890), .B2(new_n710), .ZN(new_n891));
  INV_X1    g690(.A(new_n858), .ZN(new_n892));
  OAI21_X1  g691(.A(new_n889), .B1(new_n891), .B2(new_n892), .ZN(new_n893));
  NAND3_X1  g692(.A1(new_n893), .A2(new_n879), .A3(new_n877), .ZN(new_n894));
  INV_X1    g693(.A(KEYINPUT121), .ZN(new_n895));
  NAND4_X1  g694(.A1(new_n894), .A2(new_n895), .A3(new_n256), .A4(new_n856), .ZN(new_n896));
  NAND3_X1  g695(.A1(new_n888), .A2(G141gat), .A3(new_n896), .ZN(new_n897));
  NOR2_X1   g696(.A1(new_n678), .A2(new_n430), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n831), .A2(new_n898), .ZN(new_n899));
  INV_X1    g698(.A(new_n899), .ZN(new_n900));
  NAND2_X1  g699(.A1(new_n900), .A2(KEYINPUT120), .ZN(new_n901));
  INV_X1    g700(.A(KEYINPUT120), .ZN(new_n902));
  NAND2_X1  g701(.A1(new_n899), .A2(new_n902), .ZN(new_n903));
  AND3_X1   g702(.A1(new_n901), .A2(new_n541), .A3(new_n903), .ZN(new_n904));
  NOR2_X1   g703(.A1(new_n257), .A2(G141gat), .ZN(new_n905));
  AOI21_X1  g704(.A(KEYINPUT58), .B1(new_n904), .B2(new_n905), .ZN(new_n906));
  NAND2_X1  g705(.A1(new_n897), .A2(new_n906), .ZN(new_n907));
  AND2_X1   g706(.A1(new_n887), .A2(G141gat), .ZN(new_n908));
  NAND2_X1  g707(.A1(new_n905), .A2(new_n541), .ZN(new_n909));
  OR2_X1    g708(.A1(new_n899), .A2(new_n909), .ZN(new_n910));
  INV_X1    g709(.A(KEYINPUT119), .ZN(new_n911));
  XNOR2_X1  g710(.A(new_n910), .B(new_n911), .ZN(new_n912));
  OAI21_X1  g711(.A(KEYINPUT58), .B1(new_n908), .B2(new_n912), .ZN(new_n913));
  NAND2_X1  g712(.A1(new_n907), .A2(new_n913), .ZN(G1344gat));
  NAND3_X1  g713(.A1(new_n904), .A2(new_n374), .A3(new_n662), .ZN(new_n915));
  NAND2_X1  g714(.A1(new_n894), .A2(new_n856), .ZN(new_n916));
  NOR2_X1   g715(.A1(new_n916), .A2(new_n809), .ZN(new_n917));
  INV_X1    g716(.A(KEYINPUT59), .ZN(new_n918));
  NAND2_X1  g717(.A1(new_n918), .A2(G148gat), .ZN(new_n919));
  NOR2_X1   g718(.A1(new_n917), .A2(new_n919), .ZN(new_n920));
  AOI21_X1  g719(.A(new_n711), .B1(new_n866), .B2(new_n881), .ZN(new_n921));
  OR2_X1    g720(.A1(new_n921), .A2(new_n876), .ZN(new_n922));
  NOR2_X1   g721(.A1(new_n430), .A2(KEYINPUT57), .ZN(new_n923));
  AOI22_X1  g722(.A1(new_n878), .A2(KEYINPUT57), .B1(new_n922), .B2(new_n923), .ZN(new_n924));
  NAND3_X1  g723(.A1(new_n924), .A2(new_n662), .A3(new_n856), .ZN(new_n925));
  AOI21_X1  g724(.A(new_n918), .B1(new_n925), .B2(G148gat), .ZN(new_n926));
  OAI21_X1  g725(.A(new_n915), .B1(new_n920), .B2(new_n926), .ZN(G1345gat));
  NAND3_X1  g726(.A1(new_n904), .A2(new_n360), .A3(new_n711), .ZN(new_n928));
  OAI21_X1  g727(.A(G155gat), .B1(new_n916), .B2(new_n710), .ZN(new_n929));
  NAND2_X1  g728(.A1(new_n928), .A2(new_n929), .ZN(G1346gat));
  OAI21_X1  g729(.A(G162gat), .B1(new_n916), .B2(new_n637), .ZN(new_n931));
  NAND4_X1  g730(.A1(new_n901), .A2(new_n361), .A3(new_n850), .A4(new_n903), .ZN(new_n932));
  NAND2_X1  g731(.A1(new_n931), .A2(new_n932), .ZN(G1347gat));
  AND2_X1   g732(.A1(new_n830), .A2(new_n665), .ZN(new_n934));
  NOR3_X1   g733(.A1(new_n681), .A2(new_n552), .A3(new_n541), .ZN(new_n935));
  AND2_X1   g734(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  INV_X1    g735(.A(G169gat), .ZN(new_n937));
  NAND3_X1  g736(.A1(new_n936), .A2(new_n937), .A3(new_n256), .ZN(new_n938));
  XNOR2_X1  g737(.A(new_n938), .B(KEYINPUT122), .ZN(new_n939));
  NOR2_X1   g738(.A1(new_n754), .A2(new_n541), .ZN(new_n940));
  NAND2_X1  g739(.A1(new_n940), .A2(new_n346), .ZN(new_n941));
  XNOR2_X1  g740(.A(new_n941), .B(KEYINPUT123), .ZN(new_n942));
  NAND2_X1  g741(.A1(new_n942), .A2(new_n836), .ZN(new_n943));
  OAI21_X1  g742(.A(G169gat), .B1(new_n943), .B2(new_n257), .ZN(new_n944));
  NAND2_X1  g743(.A1(new_n939), .A2(new_n944), .ZN(G1348gat));
  NAND4_X1  g744(.A1(new_n942), .A2(new_n836), .A3(G176gat), .A4(new_n709), .ZN(new_n946));
  AND2_X1   g745(.A1(new_n946), .A2(KEYINPUT124), .ZN(new_n947));
  AOI21_X1  g746(.A(G176gat), .B1(new_n936), .B2(new_n662), .ZN(new_n948));
  NOR2_X1   g747(.A1(new_n946), .A2(KEYINPUT124), .ZN(new_n949));
  NOR3_X1   g748(.A1(new_n947), .A2(new_n948), .A3(new_n949), .ZN(G1349gat));
  OR3_X1    g749(.A1(new_n943), .A2(KEYINPUT125), .A3(new_n710), .ZN(new_n951));
  OAI21_X1  g750(.A(KEYINPUT125), .B1(new_n943), .B2(new_n710), .ZN(new_n952));
  NAND3_X1  g751(.A1(new_n951), .A2(G183gat), .A3(new_n952), .ZN(new_n953));
  NAND3_X1  g752(.A1(new_n936), .A2(new_n293), .A3(new_n711), .ZN(new_n954));
  NAND2_X1  g753(.A1(new_n953), .A2(new_n954), .ZN(new_n955));
  NAND2_X1  g754(.A1(new_n955), .A2(KEYINPUT60), .ZN(new_n956));
  INV_X1    g755(.A(KEYINPUT60), .ZN(new_n957));
  NAND3_X1  g756(.A1(new_n953), .A2(new_n957), .A3(new_n954), .ZN(new_n958));
  NAND2_X1  g757(.A1(new_n956), .A2(new_n958), .ZN(G1350gat));
  OAI21_X1  g758(.A(G190gat), .B1(new_n943), .B2(new_n637), .ZN(new_n960));
  XNOR2_X1  g759(.A(new_n960), .B(KEYINPUT61), .ZN(new_n961));
  NAND3_X1  g760(.A1(new_n936), .A2(new_n273), .A3(new_n704), .ZN(new_n962));
  NAND2_X1  g761(.A1(new_n961), .A2(new_n962), .ZN(G1351gat));
  AND3_X1   g762(.A1(new_n934), .A2(new_n669), .A3(new_n898), .ZN(new_n964));
  AOI21_X1  g763(.A(G197gat), .B1(new_n964), .B2(new_n256), .ZN(new_n965));
  OR2_X1    g764(.A1(new_n924), .A2(KEYINPUT126), .ZN(new_n966));
  NAND2_X1  g765(.A1(new_n924), .A2(KEYINPUT126), .ZN(new_n967));
  NAND2_X1  g766(.A1(new_n940), .A2(new_n679), .ZN(new_n968));
  INV_X1    g767(.A(new_n968), .ZN(new_n969));
  NAND3_X1  g768(.A1(new_n966), .A2(new_n967), .A3(new_n969), .ZN(new_n970));
  INV_X1    g769(.A(new_n970), .ZN(new_n971));
  NOR2_X1   g770(.A1(new_n257), .A2(new_n238), .ZN(new_n972));
  AOI21_X1  g771(.A(new_n965), .B1(new_n971), .B2(new_n972), .ZN(G1352gat));
  OAI21_X1  g772(.A(G204gat), .B1(new_n970), .B2(new_n750), .ZN(new_n974));
  INV_X1    g773(.A(G204gat), .ZN(new_n975));
  NAND3_X1  g774(.A1(new_n964), .A2(new_n975), .A3(new_n662), .ZN(new_n976));
  XOR2_X1   g775(.A(new_n976), .B(KEYINPUT62), .Z(new_n977));
  NAND2_X1  g776(.A1(new_n974), .A2(new_n977), .ZN(G1353gat));
  NAND3_X1  g777(.A1(new_n964), .A2(new_n387), .A3(new_n711), .ZN(new_n979));
  INV_X1    g778(.A(KEYINPUT127), .ZN(new_n980));
  NOR2_X1   g779(.A1(new_n968), .A2(new_n710), .ZN(new_n981));
  NAND3_X1  g780(.A1(new_n924), .A2(new_n980), .A3(new_n981), .ZN(new_n982));
  NAND2_X1  g781(.A1(new_n982), .A2(G211gat), .ZN(new_n983));
  AOI21_X1  g782(.A(new_n980), .B1(new_n924), .B2(new_n981), .ZN(new_n984));
  NOR2_X1   g783(.A1(new_n983), .A2(new_n984), .ZN(new_n985));
  NOR2_X1   g784(.A1(new_n985), .A2(KEYINPUT63), .ZN(new_n986));
  INV_X1    g785(.A(KEYINPUT63), .ZN(new_n987));
  NOR3_X1   g786(.A1(new_n983), .A2(new_n987), .A3(new_n984), .ZN(new_n988));
  OAI21_X1  g787(.A(new_n979), .B1(new_n986), .B2(new_n988), .ZN(G1354gat));
  AOI21_X1  g788(.A(G218gat), .B1(new_n964), .B2(new_n704), .ZN(new_n990));
  NOR2_X1   g789(.A1(new_n637), .A2(new_n388), .ZN(new_n991));
  AOI21_X1  g790(.A(new_n990), .B1(new_n971), .B2(new_n991), .ZN(G1355gat));
endmodule


