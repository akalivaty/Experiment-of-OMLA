//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 1 0 0 0 0 1 1 0 0 0 0 1 1 1 0 0 0 0 1 0 1 1 0 1 0 1 1 1 1 1 0 0 1 1 1 0 0 0 0 1 0 1 0 1 1 0 1 0 0 1 1 1 1 1 1 1 1 1 1 0 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:30:53 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n437, new_n448, new_n452, new_n453, new_n454, new_n455,
    new_n458, new_n459, new_n460, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n533, new_n534, new_n535, new_n536, new_n537, new_n538,
    new_n539, new_n540, new_n541, new_n543, new_n544, new_n545, new_n546,
    new_n547, new_n550, new_n551, new_n552, new_n553, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n564, new_n566,
    new_n567, new_n569, new_n570, new_n571, new_n572, new_n573, new_n574,
    new_n575, new_n576, new_n579, new_n580, new_n581, new_n583, new_n584,
    new_n585, new_n586, new_n587, new_n588, new_n589, new_n590, new_n591,
    new_n592, new_n593, new_n595, new_n596, new_n597, new_n598, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n612, new_n613, new_n616, new_n618, new_n619,
    new_n620, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n837, new_n838, new_n839, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1144, new_n1145;
  XOR2_X1   g000(.A(KEYINPUT64), .B(G452), .Z(G350));
  XOR2_X1   g001(.A(KEYINPUT65), .B(G452), .Z(G335));
  XNOR2_X1  g002(.A(KEYINPUT66), .B(G452), .ZN(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(new_n436));
  XNOR2_X1  g011(.A(new_n436), .B(KEYINPUT67), .ZN(new_n437));
  INV_X1    g012(.A(new_n437), .ZN(G220));
  XNOR2_X1  g013(.A(KEYINPUT68), .B(G96), .ZN(G221));
  INV_X1    g014(.A(G69), .ZN(G235));
  INV_X1    g015(.A(G120), .ZN(G236));
  XNOR2_X1  g016(.A(KEYINPUT69), .B(G57), .ZN(G237));
  INV_X1    g017(.A(G108), .ZN(G238));
  NAND4_X1  g018(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g019(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g020(.A(G452), .Z(G391));
  AND2_X1   g021(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XOR2_X1   g023(.A(new_n448), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g024(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g025(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g026(.A1(G220), .A2(G218), .A3(G219), .A4(G221), .ZN(new_n452));
  XOR2_X1   g027(.A(new_n452), .B(KEYINPUT2), .Z(new_n453));
  NOR4_X1   g028(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n453), .A2(new_n455), .ZN(G325));
  XNOR2_X1  g031(.A(G325), .B(KEYINPUT70), .ZN(G261));
  NAND2_X1  g032(.A1(new_n453), .A2(G2106), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n455), .A2(G567), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  INV_X1    g035(.A(new_n460), .ZN(G319));
  NAND2_X1  g036(.A1(G113), .A2(G2104), .ZN(new_n462));
  INV_X1    g037(.A(KEYINPUT3), .ZN(new_n463));
  NOR2_X1   g038(.A1(new_n463), .A2(G2104), .ZN(new_n464));
  INV_X1    g039(.A(G2104), .ZN(new_n465));
  NOR2_X1   g040(.A1(new_n465), .A2(KEYINPUT3), .ZN(new_n466));
  OR2_X1    g041(.A1(new_n464), .A2(new_n466), .ZN(new_n467));
  INV_X1    g042(.A(G125), .ZN(new_n468));
  OAI21_X1  g043(.A(new_n462), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n469), .A2(G2105), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n465), .A2(KEYINPUT3), .ZN(new_n471));
  INV_X1    g046(.A(KEYINPUT71), .ZN(new_n472));
  OAI21_X1  g047(.A(new_n471), .B1(new_n466), .B2(new_n472), .ZN(new_n473));
  NAND3_X1  g048(.A1(new_n465), .A2(KEYINPUT71), .A3(KEYINPUT3), .ZN(new_n474));
  AND2_X1   g049(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  INV_X1    g050(.A(G2105), .ZN(new_n476));
  NAND3_X1  g051(.A1(new_n475), .A2(G137), .A3(new_n476), .ZN(new_n477));
  NAND3_X1  g052(.A1(new_n476), .A2(G101), .A3(G2104), .ZN(new_n478));
  AND3_X1   g053(.A1(new_n470), .A2(new_n477), .A3(new_n478), .ZN(G160));
  NAND2_X1  g054(.A1(new_n475), .A2(new_n476), .ZN(new_n480));
  INV_X1    g055(.A(new_n480), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n481), .A2(G136), .ZN(new_n482));
  NAND3_X1  g057(.A1(new_n473), .A2(G2105), .A3(new_n474), .ZN(new_n483));
  INV_X1    g058(.A(new_n483), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n484), .A2(G124), .ZN(new_n485));
  OR2_X1    g060(.A1(G100), .A2(G2105), .ZN(new_n486));
  OAI211_X1 g061(.A(new_n486), .B(G2104), .C1(G112), .C2(new_n476), .ZN(new_n487));
  NAND3_X1  g062(.A1(new_n482), .A2(new_n485), .A3(new_n487), .ZN(new_n488));
  INV_X1    g063(.A(new_n488), .ZN(G162));
  AND2_X1   g064(.A1(new_n476), .A2(G138), .ZN(new_n490));
  AOI21_X1  g065(.A(new_n472), .B1(new_n463), .B2(G2104), .ZN(new_n491));
  OAI211_X1 g066(.A(new_n474), .B(new_n490), .C1(new_n491), .C2(new_n464), .ZN(new_n492));
  NAND2_X1  g067(.A1(new_n492), .A2(KEYINPUT75), .ZN(new_n493));
  INV_X1    g068(.A(KEYINPUT75), .ZN(new_n494));
  NAND4_X1  g069(.A1(new_n473), .A2(new_n494), .A3(new_n474), .A4(new_n490), .ZN(new_n495));
  NAND3_X1  g070(.A1(new_n493), .A2(KEYINPUT4), .A3(new_n495), .ZN(new_n496));
  NOR2_X1   g071(.A1(new_n467), .A2(KEYINPUT4), .ZN(new_n497));
  NAND2_X1  g072(.A1(new_n497), .A2(new_n490), .ZN(new_n498));
  NAND2_X1  g073(.A1(new_n496), .A2(new_n498), .ZN(new_n499));
  NAND4_X1  g074(.A1(new_n473), .A2(G126), .A3(G2105), .A4(new_n474), .ZN(new_n500));
  INV_X1    g075(.A(KEYINPUT72), .ZN(new_n501));
  INV_X1    g076(.A(G114), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  NAND2_X1  g078(.A1(KEYINPUT72), .A2(G114), .ZN(new_n504));
  NAND3_X1  g079(.A1(new_n503), .A2(G2105), .A3(new_n504), .ZN(new_n505));
  OAI21_X1  g080(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n506));
  INV_X1    g081(.A(new_n506), .ZN(new_n507));
  AND3_X1   g082(.A1(new_n505), .A2(KEYINPUT73), .A3(new_n507), .ZN(new_n508));
  AOI21_X1  g083(.A(KEYINPUT73), .B1(new_n505), .B2(new_n507), .ZN(new_n509));
  OAI21_X1  g084(.A(new_n500), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  INV_X1    g085(.A(KEYINPUT74), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  OAI211_X1 g087(.A(KEYINPUT74), .B(new_n500), .C1(new_n508), .C2(new_n509), .ZN(new_n513));
  NAND3_X1  g088(.A1(new_n499), .A2(new_n512), .A3(new_n513), .ZN(new_n514));
  INV_X1    g089(.A(new_n514), .ZN(G164));
  INV_X1    g090(.A(KEYINPUT76), .ZN(new_n516));
  INV_X1    g091(.A(KEYINPUT6), .ZN(new_n517));
  OAI21_X1  g092(.A(new_n516), .B1(new_n517), .B2(G651), .ZN(new_n518));
  INV_X1    g093(.A(G651), .ZN(new_n519));
  NAND3_X1  g094(.A1(new_n519), .A2(KEYINPUT76), .A3(KEYINPUT6), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n518), .A2(new_n520), .ZN(new_n521));
  NAND2_X1  g096(.A1(KEYINPUT77), .A2(G543), .ZN(new_n522));
  INV_X1    g097(.A(KEYINPUT5), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  NAND3_X1  g099(.A1(KEYINPUT77), .A2(KEYINPUT5), .A3(G543), .ZN(new_n525));
  NAND2_X1  g100(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  NAND2_X1  g101(.A1(new_n517), .A2(G651), .ZN(new_n527));
  NAND3_X1  g102(.A1(new_n521), .A2(new_n526), .A3(new_n527), .ZN(new_n528));
  INV_X1    g103(.A(new_n528), .ZN(new_n529));
  NAND3_X1  g104(.A1(new_n521), .A2(G543), .A3(new_n527), .ZN(new_n530));
  INV_X1    g105(.A(new_n530), .ZN(new_n531));
  AOI22_X1  g106(.A1(G88), .A2(new_n529), .B1(new_n531), .B2(G50), .ZN(new_n532));
  NAND2_X1  g107(.A1(G75), .A2(G543), .ZN(new_n533));
  AND2_X1   g108(.A1(new_n524), .A2(new_n525), .ZN(new_n534));
  INV_X1    g109(.A(G62), .ZN(new_n535));
  OAI21_X1  g110(.A(new_n533), .B1(new_n534), .B2(new_n535), .ZN(new_n536));
  NAND2_X1  g111(.A1(new_n536), .A2(G651), .ZN(new_n537));
  NAND2_X1  g112(.A1(new_n532), .A2(new_n537), .ZN(new_n538));
  INV_X1    g113(.A(KEYINPUT78), .ZN(new_n539));
  NAND2_X1  g114(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  NAND3_X1  g115(.A1(new_n532), .A2(KEYINPUT78), .A3(new_n537), .ZN(new_n541));
  NAND2_X1  g116(.A1(new_n540), .A2(new_n541), .ZN(G166));
  NAND2_X1  g117(.A1(new_n529), .A2(G89), .ZN(new_n543));
  NAND2_X1  g118(.A1(new_n531), .A2(G51), .ZN(new_n544));
  NAND3_X1  g119(.A1(new_n526), .A2(G63), .A3(G651), .ZN(new_n545));
  NAND3_X1  g120(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n546));
  XNOR2_X1  g121(.A(new_n546), .B(KEYINPUT7), .ZN(new_n547));
  NAND4_X1  g122(.A1(new_n543), .A2(new_n544), .A3(new_n545), .A4(new_n547), .ZN(G286));
  INV_X1    g123(.A(G286), .ZN(G168));
  AOI22_X1  g124(.A1(new_n526), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n550));
  OR2_X1    g125(.A1(new_n550), .A2(new_n519), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n529), .A2(G90), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n531), .A2(G52), .ZN(new_n553));
  NAND3_X1  g128(.A1(new_n551), .A2(new_n552), .A3(new_n553), .ZN(G301));
  INV_X1    g129(.A(G301), .ZN(G171));
  AOI22_X1  g130(.A1(new_n526), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n556));
  OR2_X1    g131(.A1(new_n556), .A2(new_n519), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n529), .A2(G81), .ZN(new_n558));
  XNOR2_X1  g133(.A(KEYINPUT79), .B(G43), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n531), .A2(new_n559), .ZN(new_n560));
  AND3_X1   g135(.A1(new_n557), .A2(new_n558), .A3(new_n560), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n561), .A2(G860), .ZN(new_n562));
  XOR2_X1   g137(.A(new_n562), .B(KEYINPUT80), .Z(G153));
  AND3_X1   g138(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n564));
  NAND2_X1  g139(.A1(new_n564), .A2(G36), .ZN(G176));
  NAND2_X1  g140(.A1(G1), .A2(G3), .ZN(new_n566));
  XNOR2_X1  g141(.A(new_n566), .B(KEYINPUT8), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n564), .A2(new_n567), .ZN(G188));
  INV_X1    g143(.A(KEYINPUT81), .ZN(new_n569));
  NAND3_X1  g144(.A1(new_n531), .A2(new_n569), .A3(G53), .ZN(new_n570));
  XNOR2_X1  g145(.A(new_n570), .B(KEYINPUT9), .ZN(new_n571));
  NAND2_X1  g146(.A1(new_n529), .A2(G91), .ZN(new_n572));
  NAND2_X1  g147(.A1(G78), .A2(G543), .ZN(new_n573));
  XNOR2_X1  g148(.A(KEYINPUT82), .B(G65), .ZN(new_n574));
  OAI21_X1  g149(.A(new_n573), .B1(new_n534), .B2(new_n574), .ZN(new_n575));
  NAND2_X1  g150(.A1(new_n575), .A2(G651), .ZN(new_n576));
  NAND3_X1  g151(.A1(new_n571), .A2(new_n572), .A3(new_n576), .ZN(G299));
  INV_X1    g152(.A(G166), .ZN(G303));
  NAND2_X1  g153(.A1(new_n529), .A2(G87), .ZN(new_n579));
  NAND2_X1  g154(.A1(new_n531), .A2(G49), .ZN(new_n580));
  OAI21_X1  g155(.A(G651), .B1(new_n526), .B2(G74), .ZN(new_n581));
  NAND3_X1  g156(.A1(new_n579), .A2(new_n580), .A3(new_n581), .ZN(G288));
  NAND4_X1  g157(.A1(new_n521), .A2(new_n526), .A3(G86), .A4(new_n527), .ZN(new_n583));
  NAND4_X1  g158(.A1(new_n521), .A2(G48), .A3(G543), .A4(new_n527), .ZN(new_n584));
  AND2_X1   g159(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  NAND2_X1  g160(.A1(G73), .A2(G543), .ZN(new_n586));
  XNOR2_X1  g161(.A(new_n586), .B(KEYINPUT83), .ZN(new_n587));
  INV_X1    g162(.A(G61), .ZN(new_n588));
  AOI21_X1  g163(.A(new_n588), .B1(new_n524), .B2(new_n525), .ZN(new_n589));
  OAI21_X1  g164(.A(G651), .B1(new_n587), .B2(new_n589), .ZN(new_n590));
  INV_X1    g165(.A(KEYINPUT84), .ZN(new_n591));
  NAND2_X1  g166(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  OAI211_X1 g167(.A(KEYINPUT84), .B(G651), .C1(new_n587), .C2(new_n589), .ZN(new_n593));
  NAND3_X1  g168(.A1(new_n585), .A2(new_n592), .A3(new_n593), .ZN(G305));
  AOI22_X1  g169(.A1(new_n526), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n595));
  OR2_X1    g170(.A1(new_n595), .A2(new_n519), .ZN(new_n596));
  NAND2_X1  g171(.A1(new_n529), .A2(G85), .ZN(new_n597));
  NAND2_X1  g172(.A1(new_n531), .A2(G47), .ZN(new_n598));
  NAND3_X1  g173(.A1(new_n596), .A2(new_n597), .A3(new_n598), .ZN(G290));
  NAND2_X1  g174(.A1(G301), .A2(G868), .ZN(new_n600));
  NAND2_X1  g175(.A1(G79), .A2(G543), .ZN(new_n601));
  INV_X1    g176(.A(G66), .ZN(new_n602));
  OAI21_X1  g177(.A(new_n601), .B1(new_n534), .B2(new_n602), .ZN(new_n603));
  AOI22_X1  g178(.A1(new_n531), .A2(G54), .B1(new_n603), .B2(G651), .ZN(new_n604));
  INV_X1    g179(.A(G92), .ZN(new_n605));
  OAI21_X1  g180(.A(KEYINPUT10), .B1(new_n528), .B2(new_n605), .ZN(new_n606));
  OR3_X1    g181(.A1(new_n528), .A2(KEYINPUT10), .A3(new_n605), .ZN(new_n607));
  NAND3_X1  g182(.A1(new_n604), .A2(new_n606), .A3(new_n607), .ZN(new_n608));
  INV_X1    g183(.A(new_n608), .ZN(new_n609));
  OAI21_X1  g184(.A(new_n600), .B1(new_n609), .B2(G868), .ZN(G284));
  OAI21_X1  g185(.A(new_n600), .B1(new_n609), .B2(G868), .ZN(G321));
  NAND2_X1  g186(.A1(G286), .A2(G868), .ZN(new_n612));
  INV_X1    g187(.A(G299), .ZN(new_n613));
  OAI21_X1  g188(.A(new_n612), .B1(new_n613), .B2(G868), .ZN(G280));
  XOR2_X1   g189(.A(G280), .B(KEYINPUT85), .Z(G297));
  INV_X1    g190(.A(G559), .ZN(new_n616));
  OAI21_X1  g191(.A(new_n609), .B1(new_n616), .B2(G860), .ZN(G148));
  OAI21_X1  g192(.A(KEYINPUT86), .B1(new_n561), .B2(G868), .ZN(new_n618));
  NAND2_X1  g193(.A1(new_n609), .A2(new_n616), .ZN(new_n619));
  NAND2_X1  g194(.A1(new_n619), .A2(G868), .ZN(new_n620));
  MUX2_X1   g195(.A(KEYINPUT86), .B(new_n618), .S(new_n620), .Z(G323));
  XNOR2_X1  g196(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g197(.A1(new_n484), .A2(G123), .ZN(new_n623));
  OAI21_X1  g198(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n624));
  NOR2_X1   g199(.A1(new_n476), .A2(G111), .ZN(new_n625));
  INV_X1    g200(.A(G135), .ZN(new_n626));
  OAI221_X1 g201(.A(new_n623), .B1(new_n624), .B2(new_n625), .C1(new_n626), .C2(new_n480), .ZN(new_n627));
  INV_X1    g202(.A(KEYINPUT88), .ZN(new_n628));
  XNOR2_X1  g203(.A(new_n627), .B(new_n628), .ZN(new_n629));
  XOR2_X1   g204(.A(KEYINPUT89), .B(G2096), .Z(new_n630));
  XNOR2_X1  g205(.A(new_n629), .B(new_n630), .ZN(new_n631));
  XNOR2_X1  g206(.A(KEYINPUT87), .B(KEYINPUT12), .ZN(new_n632));
  NAND3_X1  g207(.A1(new_n476), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n633));
  XNOR2_X1  g208(.A(new_n632), .B(new_n633), .ZN(new_n634));
  XNOR2_X1  g209(.A(KEYINPUT13), .B(G2100), .ZN(new_n635));
  XNOR2_X1  g210(.A(new_n634), .B(new_n635), .ZN(new_n636));
  NAND2_X1  g211(.A1(new_n631), .A2(new_n636), .ZN(G156));
  XNOR2_X1  g212(.A(G2427), .B(G2438), .ZN(new_n638));
  XNOR2_X1  g213(.A(new_n638), .B(G2430), .ZN(new_n639));
  XNOR2_X1  g214(.A(new_n639), .B(KEYINPUT15), .ZN(new_n640));
  XOR2_X1   g215(.A(new_n640), .B(G2435), .Z(new_n641));
  NAND2_X1  g216(.A1(new_n641), .A2(KEYINPUT14), .ZN(new_n642));
  XNOR2_X1  g217(.A(G1341), .B(G1348), .ZN(new_n643));
  XNOR2_X1  g218(.A(new_n643), .B(KEYINPUT91), .ZN(new_n644));
  XOR2_X1   g219(.A(KEYINPUT90), .B(KEYINPUT16), .Z(new_n645));
  XNOR2_X1  g220(.A(new_n644), .B(new_n645), .ZN(new_n646));
  XNOR2_X1  g221(.A(G2443), .B(G2446), .ZN(new_n647));
  XNOR2_X1  g222(.A(G2451), .B(G2454), .ZN(new_n648));
  XOR2_X1   g223(.A(new_n647), .B(new_n648), .Z(new_n649));
  XNOR2_X1  g224(.A(new_n646), .B(new_n649), .ZN(new_n650));
  XNOR2_X1  g225(.A(new_n642), .B(new_n650), .ZN(new_n651));
  AND2_X1   g226(.A1(new_n651), .A2(G14), .ZN(G401));
  XNOR2_X1  g227(.A(G2067), .B(G2678), .ZN(new_n653));
  XOR2_X1   g228(.A(new_n653), .B(KEYINPUT92), .Z(new_n654));
  XOR2_X1   g229(.A(G2072), .B(G2078), .Z(new_n655));
  NAND2_X1  g230(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  XOR2_X1   g231(.A(G2084), .B(G2090), .Z(new_n657));
  INV_X1    g232(.A(new_n657), .ZN(new_n658));
  XNOR2_X1  g233(.A(new_n655), .B(KEYINPUT17), .ZN(new_n659));
  OAI211_X1 g234(.A(new_n656), .B(new_n658), .C1(new_n654), .C2(new_n659), .ZN(new_n660));
  INV_X1    g235(.A(new_n655), .ZN(new_n661));
  NAND3_X1  g236(.A1(new_n661), .A2(new_n653), .A3(new_n657), .ZN(new_n662));
  XOR2_X1   g237(.A(new_n662), .B(KEYINPUT18), .Z(new_n663));
  NAND3_X1  g238(.A1(new_n654), .A2(new_n659), .A3(new_n657), .ZN(new_n664));
  NAND3_X1  g239(.A1(new_n660), .A2(new_n663), .A3(new_n664), .ZN(new_n665));
  XOR2_X1   g240(.A(G2096), .B(G2100), .Z(new_n666));
  XNOR2_X1  g241(.A(new_n665), .B(new_n666), .ZN(G227));
  XNOR2_X1  g242(.A(G1971), .B(G1976), .ZN(new_n668));
  XNOR2_X1  g243(.A(new_n668), .B(KEYINPUT19), .ZN(new_n669));
  XOR2_X1   g244(.A(G1956), .B(G2474), .Z(new_n670));
  XOR2_X1   g245(.A(G1961), .B(G1966), .Z(new_n671));
  NAND2_X1  g246(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  NOR2_X1   g247(.A1(new_n669), .A2(new_n672), .ZN(new_n673));
  XNOR2_X1  g248(.A(new_n673), .B(KEYINPUT93), .ZN(new_n674));
  XOR2_X1   g249(.A(new_n674), .B(KEYINPUT20), .Z(new_n675));
  NOR2_X1   g250(.A1(new_n670), .A2(new_n671), .ZN(new_n676));
  INV_X1    g251(.A(new_n672), .ZN(new_n677));
  AOI21_X1  g252(.A(new_n676), .B1(new_n669), .B2(new_n677), .ZN(new_n678));
  NAND2_X1  g253(.A1(new_n669), .A2(KEYINPUT94), .ZN(new_n679));
  XNOR2_X1  g254(.A(new_n678), .B(new_n679), .ZN(new_n680));
  NAND2_X1  g255(.A1(new_n675), .A2(new_n680), .ZN(new_n681));
  XOR2_X1   g256(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n682));
  XNOR2_X1  g257(.A(new_n681), .B(new_n682), .ZN(new_n683));
  XNOR2_X1  g258(.A(G1991), .B(G1996), .ZN(new_n684));
  INV_X1    g259(.A(G1981), .ZN(new_n685));
  XNOR2_X1  g260(.A(new_n684), .B(new_n685), .ZN(new_n686));
  XNOR2_X1  g261(.A(new_n686), .B(G1986), .ZN(new_n687));
  XNOR2_X1  g262(.A(new_n683), .B(new_n687), .ZN(G229));
  NAND2_X1  g263(.A1(G166), .A2(G16), .ZN(new_n689));
  XOR2_X1   g264(.A(KEYINPUT96), .B(G1971), .Z(new_n690));
  NOR2_X1   g265(.A1(G16), .A2(G22), .ZN(new_n691));
  INV_X1    g266(.A(new_n691), .ZN(new_n692));
  NAND3_X1  g267(.A1(new_n689), .A2(new_n690), .A3(new_n692), .ZN(new_n693));
  INV_X1    g268(.A(new_n690), .ZN(new_n694));
  INV_X1    g269(.A(G16), .ZN(new_n695));
  AOI21_X1  g270(.A(new_n695), .B1(new_n540), .B2(new_n541), .ZN(new_n696));
  OAI21_X1  g271(.A(new_n694), .B1(new_n696), .B2(new_n691), .ZN(new_n697));
  AND2_X1   g272(.A1(new_n693), .A2(new_n697), .ZN(new_n698));
  INV_X1    g273(.A(KEYINPUT97), .ZN(new_n699));
  NAND2_X1  g274(.A1(new_n695), .A2(G23), .ZN(new_n700));
  INV_X1    g275(.A(G288), .ZN(new_n701));
  OAI21_X1  g276(.A(new_n700), .B1(new_n701), .B2(new_n695), .ZN(new_n702));
  XNOR2_X1  g277(.A(KEYINPUT33), .B(G1976), .ZN(new_n703));
  XNOR2_X1  g278(.A(new_n702), .B(new_n703), .ZN(new_n704));
  OR2_X1    g279(.A1(G6), .A2(G16), .ZN(new_n705));
  OAI21_X1  g280(.A(new_n705), .B1(G305), .B2(new_n695), .ZN(new_n706));
  XNOR2_X1  g281(.A(KEYINPUT32), .B(G1981), .ZN(new_n707));
  XNOR2_X1  g282(.A(new_n706), .B(new_n707), .ZN(new_n708));
  NAND4_X1  g283(.A1(new_n698), .A2(new_n699), .A3(new_n704), .A4(new_n708), .ZN(new_n709));
  NAND3_X1  g284(.A1(new_n693), .A2(new_n704), .A3(new_n697), .ZN(new_n710));
  INV_X1    g285(.A(new_n708), .ZN(new_n711));
  OAI21_X1  g286(.A(KEYINPUT97), .B1(new_n710), .B2(new_n711), .ZN(new_n712));
  NAND3_X1  g287(.A1(new_n709), .A2(new_n712), .A3(KEYINPUT34), .ZN(new_n713));
  AOI21_X1  g288(.A(KEYINPUT34), .B1(new_n709), .B2(new_n712), .ZN(new_n714));
  INV_X1    g289(.A(G29), .ZN(new_n715));
  NAND2_X1  g290(.A1(new_n715), .A2(G25), .ZN(new_n716));
  NAND2_X1  g291(.A1(new_n481), .A2(G131), .ZN(new_n717));
  NAND2_X1  g292(.A1(new_n484), .A2(G119), .ZN(new_n718));
  OR2_X1    g293(.A1(G95), .A2(G2105), .ZN(new_n719));
  OAI211_X1 g294(.A(new_n719), .B(G2104), .C1(G107), .C2(new_n476), .ZN(new_n720));
  NAND3_X1  g295(.A1(new_n717), .A2(new_n718), .A3(new_n720), .ZN(new_n721));
  INV_X1    g296(.A(new_n721), .ZN(new_n722));
  OAI21_X1  g297(.A(new_n716), .B1(new_n722), .B2(new_n715), .ZN(new_n723));
  XOR2_X1   g298(.A(KEYINPUT35), .B(G1991), .Z(new_n724));
  XNOR2_X1  g299(.A(new_n724), .B(KEYINPUT95), .ZN(new_n725));
  XOR2_X1   g300(.A(new_n723), .B(new_n725), .Z(new_n726));
  OR2_X1    g301(.A1(G16), .A2(G24), .ZN(new_n727));
  OAI21_X1  g302(.A(new_n727), .B1(G290), .B2(new_n695), .ZN(new_n728));
  INV_X1    g303(.A(G1986), .ZN(new_n729));
  XNOR2_X1  g304(.A(new_n728), .B(new_n729), .ZN(new_n730));
  NOR3_X1   g305(.A1(new_n714), .A2(new_n726), .A3(new_n730), .ZN(new_n731));
  NOR2_X1   g306(.A1(new_n731), .A2(KEYINPUT98), .ZN(new_n732));
  INV_X1    g307(.A(KEYINPUT98), .ZN(new_n733));
  NOR4_X1   g308(.A1(new_n714), .A2(new_n733), .A3(new_n726), .A4(new_n730), .ZN(new_n734));
  OAI21_X1  g309(.A(new_n713), .B1(new_n732), .B2(new_n734), .ZN(new_n735));
  NAND2_X1  g310(.A1(KEYINPUT99), .A2(KEYINPUT36), .ZN(new_n736));
  NAND2_X1  g311(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  NAND2_X1  g312(.A1(new_n695), .A2(G21), .ZN(new_n738));
  OAI21_X1  g313(.A(new_n738), .B1(G168), .B2(new_n695), .ZN(new_n739));
  XOR2_X1   g314(.A(new_n739), .B(KEYINPUT105), .Z(new_n740));
  INV_X1    g315(.A(G1966), .ZN(new_n741));
  NAND2_X1  g316(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  NAND2_X1  g317(.A1(new_n715), .A2(G26), .ZN(new_n743));
  NAND2_X1  g318(.A1(new_n481), .A2(G140), .ZN(new_n744));
  NAND2_X1  g319(.A1(new_n484), .A2(G128), .ZN(new_n745));
  OR2_X1    g320(.A1(G104), .A2(G2105), .ZN(new_n746));
  OAI211_X1 g321(.A(new_n746), .B(G2104), .C1(G116), .C2(new_n476), .ZN(new_n747));
  NAND3_X1  g322(.A1(new_n744), .A2(new_n745), .A3(new_n747), .ZN(new_n748));
  INV_X1    g323(.A(new_n748), .ZN(new_n749));
  OAI21_X1  g324(.A(new_n743), .B1(new_n749), .B2(new_n715), .ZN(new_n750));
  MUX2_X1   g325(.A(new_n743), .B(new_n750), .S(KEYINPUT28), .Z(new_n751));
  INV_X1    g326(.A(G2067), .ZN(new_n752));
  XNOR2_X1  g327(.A(new_n751), .B(new_n752), .ZN(new_n753));
  INV_X1    g328(.A(KEYINPUT24), .ZN(new_n754));
  OAI21_X1  g329(.A(new_n715), .B1(new_n754), .B2(G34), .ZN(new_n755));
  INV_X1    g330(.A(KEYINPUT102), .ZN(new_n756));
  OR2_X1    g331(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  NAND2_X1  g332(.A1(new_n754), .A2(G34), .ZN(new_n758));
  NAND2_X1  g333(.A1(new_n755), .A2(new_n756), .ZN(new_n759));
  NAND3_X1  g334(.A1(new_n757), .A2(new_n758), .A3(new_n759), .ZN(new_n760));
  NAND3_X1  g335(.A1(new_n470), .A2(new_n477), .A3(new_n478), .ZN(new_n761));
  OAI21_X1  g336(.A(new_n760), .B1(new_n761), .B2(new_n715), .ZN(new_n762));
  XNOR2_X1  g337(.A(new_n762), .B(G2084), .ZN(new_n763));
  NAND3_X1  g338(.A1(new_n695), .A2(KEYINPUT23), .A3(G20), .ZN(new_n764));
  INV_X1    g339(.A(KEYINPUT23), .ZN(new_n765));
  INV_X1    g340(.A(G20), .ZN(new_n766));
  OAI21_X1  g341(.A(new_n765), .B1(new_n766), .B2(G16), .ZN(new_n767));
  OAI211_X1 g342(.A(new_n764), .B(new_n767), .C1(new_n613), .C2(new_n695), .ZN(new_n768));
  INV_X1    g343(.A(G1956), .ZN(new_n769));
  XNOR2_X1  g344(.A(new_n768), .B(new_n769), .ZN(new_n770));
  NAND2_X1  g345(.A1(new_n695), .A2(G19), .ZN(new_n771));
  OAI21_X1  g346(.A(new_n771), .B1(new_n561), .B2(new_n695), .ZN(new_n772));
  XNOR2_X1  g347(.A(new_n772), .B(G1341), .ZN(new_n773));
  NOR2_X1   g348(.A1(G4), .A2(G16), .ZN(new_n774));
  AOI21_X1  g349(.A(new_n774), .B1(new_n609), .B2(G16), .ZN(new_n775));
  INV_X1    g350(.A(KEYINPUT31), .ZN(new_n776));
  OAI22_X1  g351(.A1(new_n775), .A2(G1348), .B1(new_n776), .B2(G11), .ZN(new_n777));
  NOR2_X1   g352(.A1(new_n773), .A2(new_n777), .ZN(new_n778));
  NAND4_X1  g353(.A1(new_n753), .A2(new_n763), .A3(new_n770), .A4(new_n778), .ZN(new_n779));
  XOR2_X1   g354(.A(KEYINPUT106), .B(KEYINPUT30), .Z(new_n780));
  XOR2_X1   g355(.A(new_n780), .B(G28), .Z(new_n781));
  NOR2_X1   g356(.A1(new_n781), .A2(G29), .ZN(new_n782));
  NAND2_X1  g357(.A1(new_n715), .A2(G32), .ZN(new_n783));
  NAND2_X1  g358(.A1(new_n484), .A2(G129), .ZN(new_n784));
  NAND3_X1  g359(.A1(new_n476), .A2(G105), .A3(G2104), .ZN(new_n785));
  INV_X1    g360(.A(G141), .ZN(new_n786));
  OAI211_X1 g361(.A(new_n784), .B(new_n785), .C1(new_n786), .C2(new_n480), .ZN(new_n787));
  NAND3_X1  g362(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n788));
  XNOR2_X1  g363(.A(new_n788), .B(KEYINPUT103), .ZN(new_n789));
  XOR2_X1   g364(.A(new_n789), .B(KEYINPUT26), .Z(new_n790));
  NOR2_X1   g365(.A1(new_n787), .A2(new_n790), .ZN(new_n791));
  INV_X1    g366(.A(KEYINPUT104), .ZN(new_n792));
  XNOR2_X1  g367(.A(new_n791), .B(new_n792), .ZN(new_n793));
  OAI21_X1  g368(.A(new_n783), .B1(new_n793), .B2(new_n715), .ZN(new_n794));
  XOR2_X1   g369(.A(KEYINPUT27), .B(G1996), .Z(new_n795));
  NOR2_X1   g370(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  AOI211_X1 g371(.A(new_n782), .B(new_n796), .C1(G1348), .C2(new_n775), .ZN(new_n797));
  INV_X1    g372(.A(new_n740), .ZN(new_n798));
  AOI22_X1  g373(.A1(new_n798), .A2(G1966), .B1(new_n795), .B2(new_n794), .ZN(new_n799));
  NAND2_X1  g374(.A1(new_n715), .A2(G27), .ZN(new_n800));
  OAI21_X1  g375(.A(new_n800), .B1(G164), .B2(new_n715), .ZN(new_n801));
  INV_X1    g376(.A(G2078), .ZN(new_n802));
  XNOR2_X1  g377(.A(new_n801), .B(new_n802), .ZN(new_n803));
  NOR2_X1   g378(.A1(new_n629), .A2(new_n715), .ZN(new_n804));
  NAND2_X1  g379(.A1(G171), .A2(G16), .ZN(new_n805));
  OAI21_X1  g380(.A(new_n805), .B1(G5), .B2(G16), .ZN(new_n806));
  INV_X1    g381(.A(G1961), .ZN(new_n807));
  AND2_X1   g382(.A1(new_n806), .A2(new_n807), .ZN(new_n808));
  NOR2_X1   g383(.A1(new_n806), .A2(new_n807), .ZN(new_n809));
  NOR3_X1   g384(.A1(new_n804), .A2(new_n808), .A3(new_n809), .ZN(new_n810));
  NAND4_X1  g385(.A1(new_n797), .A2(new_n799), .A3(new_n803), .A4(new_n810), .ZN(new_n811));
  AOI211_X1 g386(.A(new_n779), .B(new_n811), .C1(new_n776), .C2(G11), .ZN(new_n812));
  INV_X1    g387(.A(new_n736), .ZN(new_n813));
  OAI211_X1 g388(.A(new_n713), .B(new_n813), .C1(new_n732), .C2(new_n734), .ZN(new_n814));
  NAND4_X1  g389(.A1(new_n737), .A2(new_n742), .A3(new_n812), .A4(new_n814), .ZN(new_n815));
  NAND2_X1  g390(.A1(new_n715), .A2(G33), .ZN(new_n816));
  NAND2_X1  g391(.A1(new_n481), .A2(G139), .ZN(new_n817));
  XNOR2_X1  g392(.A(new_n817), .B(KEYINPUT100), .ZN(new_n818));
  NAND2_X1  g393(.A1(G115), .A2(G2104), .ZN(new_n819));
  INV_X1    g394(.A(G127), .ZN(new_n820));
  OAI21_X1  g395(.A(new_n819), .B1(new_n467), .B2(new_n820), .ZN(new_n821));
  NAND2_X1  g396(.A1(new_n821), .A2(G2105), .ZN(new_n822));
  NAND3_X1  g397(.A1(new_n476), .A2(G103), .A3(G2104), .ZN(new_n823));
  XOR2_X1   g398(.A(new_n823), .B(KEYINPUT25), .Z(new_n824));
  NAND3_X1  g399(.A1(new_n818), .A2(new_n822), .A3(new_n824), .ZN(new_n825));
  INV_X1    g400(.A(KEYINPUT101), .ZN(new_n826));
  NAND2_X1  g401(.A1(new_n825), .A2(new_n826), .ZN(new_n827));
  NAND4_X1  g402(.A1(new_n818), .A2(KEYINPUT101), .A3(new_n822), .A4(new_n824), .ZN(new_n828));
  AND2_X1   g403(.A1(new_n827), .A2(new_n828), .ZN(new_n829));
  OAI21_X1  g404(.A(new_n816), .B1(new_n829), .B2(new_n715), .ZN(new_n830));
  XNOR2_X1  g405(.A(new_n830), .B(G2072), .ZN(new_n831));
  NAND2_X1  g406(.A1(new_n715), .A2(G35), .ZN(new_n832));
  OAI21_X1  g407(.A(new_n832), .B1(G162), .B2(new_n715), .ZN(new_n833));
  XNOR2_X1  g408(.A(KEYINPUT29), .B(G2090), .ZN(new_n834));
  XNOR2_X1  g409(.A(new_n833), .B(new_n834), .ZN(new_n835));
  NOR3_X1   g410(.A1(new_n815), .A2(new_n831), .A3(new_n835), .ZN(G311));
  AND3_X1   g411(.A1(new_n737), .A2(new_n814), .A3(new_n812), .ZN(new_n837));
  INV_X1    g412(.A(new_n831), .ZN(new_n838));
  INV_X1    g413(.A(new_n835), .ZN(new_n839));
  NAND4_X1  g414(.A1(new_n837), .A2(new_n838), .A3(new_n839), .A4(new_n742), .ZN(G150));
  NAND2_X1  g415(.A1(new_n529), .A2(G93), .ZN(new_n841));
  NAND2_X1  g416(.A1(new_n531), .A2(G55), .ZN(new_n842));
  AOI22_X1  g417(.A1(new_n526), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n843));
  OAI211_X1 g418(.A(new_n841), .B(new_n842), .C1(new_n519), .C2(new_n843), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n844), .A2(G860), .ZN(new_n845));
  XOR2_X1   g420(.A(new_n845), .B(KEYINPUT37), .Z(new_n846));
  XNOR2_X1  g421(.A(new_n561), .B(new_n844), .ZN(new_n847));
  XNOR2_X1  g422(.A(new_n847), .B(KEYINPUT39), .ZN(new_n848));
  NAND2_X1  g423(.A1(new_n609), .A2(G559), .ZN(new_n849));
  XNOR2_X1  g424(.A(new_n849), .B(KEYINPUT38), .ZN(new_n850));
  XNOR2_X1  g425(.A(new_n848), .B(new_n850), .ZN(new_n851));
  OAI21_X1  g426(.A(new_n846), .B1(new_n851), .B2(G860), .ZN(G145));
  INV_X1    g427(.A(G142), .ZN(new_n853));
  OAI21_X1  g428(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n854));
  NOR2_X1   g429(.A1(new_n476), .A2(G118), .ZN(new_n855));
  OAI22_X1  g430(.A1(new_n480), .A2(new_n853), .B1(new_n854), .B2(new_n855), .ZN(new_n856));
  AOI21_X1  g431(.A(new_n856), .B1(G130), .B2(new_n484), .ZN(new_n857));
  XNOR2_X1  g432(.A(new_n722), .B(new_n857), .ZN(new_n858));
  XNOR2_X1  g433(.A(new_n858), .B(new_n634), .ZN(new_n859));
  XNOR2_X1  g434(.A(new_n791), .B(new_n748), .ZN(new_n860));
  INV_X1    g435(.A(new_n510), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n499), .A2(new_n861), .ZN(new_n862));
  XNOR2_X1  g437(.A(new_n860), .B(new_n862), .ZN(new_n863));
  INV_X1    g438(.A(KEYINPUT107), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n829), .A2(new_n864), .ZN(new_n865));
  NAND3_X1  g440(.A1(new_n827), .A2(new_n792), .A3(new_n828), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n866), .A2(KEYINPUT107), .ZN(new_n867));
  AOI21_X1  g442(.A(new_n863), .B1(new_n865), .B2(new_n867), .ZN(new_n868));
  AND2_X1   g443(.A1(new_n867), .A2(new_n863), .ZN(new_n869));
  OAI21_X1  g444(.A(new_n859), .B1(new_n868), .B2(new_n869), .ZN(new_n870));
  NOR3_X1   g445(.A1(new_n868), .A2(new_n869), .A3(new_n859), .ZN(new_n871));
  OAI21_X1  g446(.A(new_n870), .B1(new_n871), .B2(KEYINPUT108), .ZN(new_n872));
  XNOR2_X1  g447(.A(new_n629), .B(new_n761), .ZN(new_n873));
  XNOR2_X1  g448(.A(new_n873), .B(new_n488), .ZN(new_n874));
  INV_X1    g449(.A(new_n874), .ZN(new_n875));
  INV_X1    g450(.A(KEYINPUT108), .ZN(new_n876));
  OAI211_X1 g451(.A(new_n876), .B(new_n859), .C1(new_n868), .C2(new_n869), .ZN(new_n877));
  NAND3_X1  g452(.A1(new_n872), .A2(new_n875), .A3(new_n877), .ZN(new_n878));
  INV_X1    g453(.A(KEYINPUT109), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  INV_X1    g455(.A(new_n871), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n881), .A2(new_n870), .ZN(new_n882));
  AOI21_X1  g457(.A(G37), .B1(new_n882), .B2(new_n874), .ZN(new_n883));
  NAND4_X1  g458(.A1(new_n872), .A2(new_n877), .A3(KEYINPUT109), .A4(new_n875), .ZN(new_n884));
  NAND3_X1  g459(.A1(new_n880), .A2(new_n883), .A3(new_n884), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n885), .A2(KEYINPUT40), .ZN(new_n886));
  INV_X1    g461(.A(KEYINPUT40), .ZN(new_n887));
  NAND4_X1  g462(.A1(new_n880), .A2(new_n883), .A3(new_n887), .A4(new_n884), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n886), .A2(new_n888), .ZN(G395));
  XNOR2_X1  g464(.A(G166), .B(G290), .ZN(new_n890));
  XOR2_X1   g465(.A(G305), .B(G288), .Z(new_n891));
  XNOR2_X1  g466(.A(new_n890), .B(new_n891), .ZN(new_n892));
  NOR2_X1   g467(.A1(new_n892), .A2(KEYINPUT42), .ZN(new_n893));
  XNOR2_X1  g468(.A(new_n892), .B(KEYINPUT110), .ZN(new_n894));
  AOI21_X1  g469(.A(new_n893), .B1(new_n894), .B2(KEYINPUT42), .ZN(new_n895));
  XNOR2_X1  g470(.A(new_n847), .B(new_n619), .ZN(new_n896));
  XNOR2_X1  g471(.A(G299), .B(new_n608), .ZN(new_n897));
  NOR2_X1   g472(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n897), .A2(KEYINPUT41), .ZN(new_n899));
  XNOR2_X1  g474(.A(G299), .B(new_n609), .ZN(new_n900));
  INV_X1    g475(.A(KEYINPUT41), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n899), .A2(new_n902), .ZN(new_n903));
  AOI21_X1  g478(.A(new_n898), .B1(new_n903), .B2(new_n896), .ZN(new_n904));
  OR2_X1    g479(.A1(new_n895), .A2(new_n904), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n895), .A2(new_n904), .ZN(new_n906));
  NAND3_X1  g481(.A1(new_n905), .A2(G868), .A3(new_n906), .ZN(new_n907));
  INV_X1    g482(.A(KEYINPUT111), .ZN(new_n908));
  NOR2_X1   g483(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  INV_X1    g484(.A(G868), .ZN(new_n910));
  AOI21_X1  g485(.A(KEYINPUT111), .B1(new_n844), .B2(new_n910), .ZN(new_n911));
  AOI21_X1  g486(.A(new_n909), .B1(new_n911), .B2(new_n907), .ZN(G295));
  AOI21_X1  g487(.A(new_n909), .B1(new_n911), .B2(new_n907), .ZN(G331));
  XNOR2_X1  g488(.A(G171), .B(G286), .ZN(new_n914));
  AOI21_X1  g489(.A(KEYINPUT112), .B1(new_n914), .B2(new_n847), .ZN(new_n915));
  XNOR2_X1  g490(.A(new_n914), .B(new_n847), .ZN(new_n916));
  AOI21_X1  g491(.A(new_n915), .B1(new_n916), .B2(KEYINPUT112), .ZN(new_n917));
  INV_X1    g492(.A(new_n917), .ZN(new_n918));
  NAND3_X1  g493(.A1(new_n897), .A2(KEYINPUT113), .A3(KEYINPUT41), .ZN(new_n919));
  OAI211_X1 g494(.A(new_n918), .B(new_n919), .C1(new_n903), .C2(KEYINPUT113), .ZN(new_n920));
  OAI21_X1  g495(.A(new_n920), .B1(new_n897), .B2(new_n916), .ZN(new_n921));
  INV_X1    g496(.A(KEYINPUT110), .ZN(new_n922));
  XNOR2_X1  g497(.A(new_n892), .B(new_n922), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n921), .A2(new_n923), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n917), .A2(new_n900), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n903), .A2(new_n916), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  INV_X1    g502(.A(new_n927), .ZN(new_n928));
  AOI21_X1  g503(.A(G37), .B1(new_n894), .B2(new_n928), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n924), .A2(new_n929), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n930), .A2(KEYINPUT43), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n931), .A2(KEYINPUT114), .ZN(new_n932));
  INV_X1    g507(.A(KEYINPUT114), .ZN(new_n933));
  NAND3_X1  g508(.A1(new_n930), .A2(new_n933), .A3(KEYINPUT43), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n932), .A2(new_n934), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n923), .A2(new_n927), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n929), .A2(new_n936), .ZN(new_n937));
  OAI21_X1  g512(.A(KEYINPUT44), .B1(new_n937), .B2(KEYINPUT43), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n937), .A2(KEYINPUT43), .ZN(new_n939));
  INV_X1    g514(.A(KEYINPUT43), .ZN(new_n940));
  NAND3_X1  g515(.A1(new_n924), .A2(new_n929), .A3(new_n940), .ZN(new_n941));
  AND2_X1   g516(.A1(new_n939), .A2(new_n941), .ZN(new_n942));
  OAI22_X1  g517(.A1(new_n935), .A2(new_n938), .B1(KEYINPUT44), .B2(new_n942), .ZN(G397));
  AOI21_X1  g518(.A(new_n510), .B1(new_n496), .B2(new_n498), .ZN(new_n944));
  XNOR2_X1  g519(.A(KEYINPUT115), .B(G1384), .ZN(new_n945));
  NOR2_X1   g520(.A1(new_n944), .A2(new_n945), .ZN(new_n946));
  NOR2_X1   g521(.A1(new_n946), .A2(KEYINPUT45), .ZN(new_n947));
  INV_X1    g522(.A(G40), .ZN(new_n948));
  NOR2_X1   g523(.A1(new_n761), .A2(new_n948), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n947), .A2(new_n949), .ZN(new_n950));
  INV_X1    g525(.A(new_n950), .ZN(new_n951));
  XNOR2_X1  g526(.A(new_n748), .B(new_n752), .ZN(new_n952));
  XNOR2_X1  g527(.A(new_n952), .B(KEYINPUT116), .ZN(new_n953));
  INV_X1    g528(.A(G1996), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n793), .A2(new_n954), .ZN(new_n955));
  OAI21_X1  g530(.A(G1996), .B1(new_n787), .B2(new_n790), .ZN(new_n956));
  NAND3_X1  g531(.A1(new_n953), .A2(new_n955), .A3(new_n956), .ZN(new_n957));
  INV_X1    g532(.A(new_n957), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n722), .A2(new_n725), .ZN(new_n959));
  OR2_X1    g534(.A1(new_n722), .A2(new_n725), .ZN(new_n960));
  NAND3_X1  g535(.A1(new_n958), .A2(new_n959), .A3(new_n960), .ZN(new_n961));
  XNOR2_X1  g536(.A(G290), .B(G1986), .ZN(new_n962));
  OAI21_X1  g537(.A(new_n951), .B1(new_n961), .B2(new_n962), .ZN(new_n963));
  NAND2_X1  g538(.A1(G286), .A2(G8), .ZN(new_n964));
  INV_X1    g539(.A(G8), .ZN(new_n965));
  INV_X1    g540(.A(G2084), .ZN(new_n966));
  NAND2_X1  g541(.A1(G160), .A2(G40), .ZN(new_n967));
  NOR2_X1   g542(.A1(new_n944), .A2(G1384), .ZN(new_n968));
  INV_X1    g543(.A(KEYINPUT50), .ZN(new_n969));
  AOI21_X1  g544(.A(new_n967), .B1(new_n968), .B2(new_n969), .ZN(new_n970));
  INV_X1    g545(.A(KEYINPUT118), .ZN(new_n971));
  INV_X1    g546(.A(G1384), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n514), .A2(new_n972), .ZN(new_n973));
  AOI21_X1  g548(.A(new_n971), .B1(new_n973), .B2(KEYINPUT50), .ZN(new_n974));
  AOI211_X1 g549(.A(KEYINPUT118), .B(new_n969), .C1(new_n514), .C2(new_n972), .ZN(new_n975));
  OAI211_X1 g550(.A(new_n966), .B(new_n970), .C1(new_n974), .C2(new_n975), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n862), .A2(new_n972), .ZN(new_n977));
  INV_X1    g552(.A(KEYINPUT45), .ZN(new_n978));
  NAND2_X1  g553(.A1(new_n977), .A2(new_n978), .ZN(new_n979));
  OAI211_X1 g554(.A(new_n979), .B(new_n949), .C1(new_n978), .C2(new_n973), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n980), .A2(new_n741), .ZN(new_n981));
  AOI21_X1  g556(.A(new_n965), .B1(new_n976), .B2(new_n981), .ZN(new_n982));
  INV_X1    g557(.A(KEYINPUT51), .ZN(new_n983));
  NOR2_X1   g558(.A1(new_n983), .A2(KEYINPUT125), .ZN(new_n984));
  OAI21_X1  g559(.A(new_n964), .B1(new_n982), .B2(new_n984), .ZN(new_n985));
  AOI211_X1 g560(.A(KEYINPUT125), .B(new_n965), .C1(new_n976), .C2(new_n981), .ZN(new_n986));
  NOR2_X1   g561(.A1(new_n985), .A2(new_n986), .ZN(new_n987));
  NOR2_X1   g562(.A1(new_n983), .A2(KEYINPUT124), .ZN(new_n988));
  AOI21_X1  g563(.A(new_n988), .B1(new_n982), .B2(G286), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n983), .A2(KEYINPUT124), .ZN(new_n990));
  INV_X1    g565(.A(new_n990), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n976), .A2(new_n981), .ZN(new_n992));
  OAI211_X1 g567(.A(G8), .B(new_n991), .C1(new_n992), .C2(G286), .ZN(new_n993));
  NAND2_X1  g568(.A1(new_n989), .A2(new_n993), .ZN(new_n994));
  OAI21_X1  g569(.A(KEYINPUT62), .B1(new_n987), .B2(new_n994), .ZN(new_n995));
  OAI21_X1  g570(.A(new_n970), .B1(new_n974), .B2(new_n975), .ZN(new_n996));
  INV_X1    g571(.A(KEYINPUT53), .ZN(new_n997));
  AOI21_X1  g572(.A(new_n967), .B1(new_n946), .B2(KEYINPUT45), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n973), .A2(new_n978), .ZN(new_n999));
  NAND3_X1  g574(.A1(new_n998), .A2(new_n999), .A3(new_n802), .ZN(new_n1000));
  AOI22_X1  g575(.A1(new_n996), .A2(new_n807), .B1(new_n997), .B2(new_n1000), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n802), .A2(KEYINPUT53), .ZN(new_n1002));
  OR2_X1    g577(.A1(new_n980), .A2(new_n1002), .ZN(new_n1003));
  AOI21_X1  g578(.A(G301), .B1(new_n1001), .B2(new_n1003), .ZN(new_n1004));
  INV_X1    g579(.A(G1971), .ZN(new_n1005));
  INV_X1    g580(.A(new_n945), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n862), .A2(new_n1006), .ZN(new_n1007));
  OAI21_X1  g582(.A(new_n949), .B1(new_n1007), .B2(new_n978), .ZN(new_n1008));
  AOI21_X1  g583(.A(KEYINPUT45), .B1(new_n514), .B2(new_n972), .ZN(new_n1009));
  OAI21_X1  g584(.A(new_n1005), .B1(new_n1008), .B2(new_n1009), .ZN(new_n1010));
  NAND3_X1  g585(.A1(new_n514), .A2(new_n969), .A3(new_n972), .ZN(new_n1011));
  INV_X1    g586(.A(G2090), .ZN(new_n1012));
  OAI21_X1  g587(.A(KEYINPUT50), .B1(new_n944), .B2(G1384), .ZN(new_n1013));
  NAND4_X1  g588(.A1(new_n1011), .A2(new_n1012), .A3(new_n949), .A4(new_n1013), .ZN(new_n1014));
  AOI21_X1  g589(.A(new_n965), .B1(new_n1010), .B2(new_n1014), .ZN(new_n1015));
  NAND3_X1  g590(.A1(new_n540), .A2(G8), .A3(new_n541), .ZN(new_n1016));
  XNOR2_X1  g591(.A(new_n1016), .B(KEYINPUT55), .ZN(new_n1017));
  INV_X1    g592(.A(new_n1017), .ZN(new_n1018));
  OAI21_X1  g593(.A(KEYINPUT121), .B1(new_n1015), .B2(new_n1018), .ZN(new_n1019));
  AOI21_X1  g594(.A(G1971), .B1(new_n998), .B2(new_n999), .ZN(new_n1020));
  INV_X1    g595(.A(new_n1014), .ZN(new_n1021));
  OAI21_X1  g596(.A(G8), .B1(new_n1020), .B2(new_n1021), .ZN(new_n1022));
  INV_X1    g597(.A(KEYINPUT121), .ZN(new_n1023));
  NAND3_X1  g598(.A1(new_n1022), .A2(new_n1023), .A3(new_n1017), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n1019), .A2(new_n1024), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n1020), .A2(KEYINPUT117), .ZN(new_n1026));
  INV_X1    g601(.A(KEYINPUT117), .ZN(new_n1027));
  NAND2_X1  g602(.A1(new_n1010), .A2(new_n1027), .ZN(new_n1028));
  OAI211_X1 g603(.A(new_n1026), .B(new_n1028), .C1(G2090), .C2(new_n996), .ZN(new_n1029));
  NAND3_X1  g604(.A1(new_n1029), .A2(G8), .A3(new_n1018), .ZN(new_n1030));
  INV_X1    g605(.A(KEYINPUT49), .ZN(new_n1031));
  NAND2_X1  g606(.A1(G305), .A2(G1981), .ZN(new_n1032));
  NAND4_X1  g607(.A1(new_n585), .A2(new_n592), .A3(new_n685), .A4(new_n593), .ZN(new_n1033));
  NAND3_X1  g608(.A1(new_n1032), .A2(KEYINPUT119), .A3(new_n1033), .ZN(new_n1034));
  INV_X1    g609(.A(KEYINPUT119), .ZN(new_n1035));
  NAND3_X1  g610(.A1(G305), .A2(new_n1035), .A3(G1981), .ZN(new_n1036));
  AOI21_X1  g611(.A(new_n1031), .B1(new_n1034), .B2(new_n1036), .ZN(new_n1037));
  OR2_X1    g612(.A1(new_n1037), .A2(KEYINPUT120), .ZN(new_n1038));
  NAND3_X1  g613(.A1(new_n1034), .A2(new_n1031), .A3(new_n1036), .ZN(new_n1039));
  AOI21_X1  g614(.A(new_n965), .B1(new_n968), .B2(new_n949), .ZN(new_n1040));
  AND2_X1   g615(.A1(new_n1039), .A2(new_n1040), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n1037), .A2(KEYINPUT120), .ZN(new_n1042));
  NAND3_X1  g617(.A1(new_n1038), .A2(new_n1041), .A3(new_n1042), .ZN(new_n1043));
  INV_X1    g618(.A(G1976), .ZN(new_n1044));
  OAI21_X1  g619(.A(new_n1040), .B1(new_n1044), .B2(G288), .ZN(new_n1045));
  NOR2_X1   g620(.A1(new_n701), .A2(G1976), .ZN(new_n1046));
  OR3_X1    g621(.A1(new_n1045), .A2(KEYINPUT52), .A3(new_n1046), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n1045), .A2(KEYINPUT52), .ZN(new_n1048));
  AND3_X1   g623(.A1(new_n1043), .A2(new_n1047), .A3(new_n1048), .ZN(new_n1049));
  AND4_X1   g624(.A1(new_n1004), .A2(new_n1025), .A3(new_n1030), .A4(new_n1049), .ZN(new_n1050));
  INV_X1    g625(.A(KEYINPUT125), .ZN(new_n1051));
  NAND3_X1  g626(.A1(new_n992), .A2(new_n1051), .A3(G8), .ZN(new_n1052));
  OAI211_X1 g627(.A(new_n1052), .B(new_n964), .C1(new_n982), .C2(new_n984), .ZN(new_n1053));
  INV_X1    g628(.A(KEYINPUT62), .ZN(new_n1054));
  NAND4_X1  g629(.A1(new_n1053), .A2(new_n1054), .A3(new_n993), .A4(new_n989), .ZN(new_n1055));
  NAND3_X1  g630(.A1(new_n995), .A2(new_n1050), .A3(new_n1055), .ZN(new_n1056));
  INV_X1    g631(.A(KEYINPUT127), .ZN(new_n1057));
  NAND2_X1  g632(.A1(new_n1056), .A2(new_n1057), .ZN(new_n1058));
  NAND4_X1  g633(.A1(new_n995), .A2(new_n1050), .A3(new_n1055), .A4(KEYINPUT127), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n1058), .A2(new_n1059), .ZN(new_n1060));
  OR2_X1    g635(.A1(new_n1029), .A2(new_n1018), .ZN(new_n1061));
  NAND4_X1  g636(.A1(new_n1061), .A2(G168), .A3(new_n982), .A4(new_n1049), .ZN(new_n1062));
  NAND3_X1  g637(.A1(new_n1043), .A2(new_n1044), .A3(new_n701), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n1063), .A2(new_n1033), .ZN(new_n1064));
  AOI22_X1  g639(.A1(new_n1062), .A2(KEYINPUT63), .B1(new_n1040), .B2(new_n1064), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n1060), .A2(new_n1065), .ZN(new_n1066));
  INV_X1    g641(.A(new_n1049), .ZN(new_n1067));
  NOR2_X1   g642(.A1(new_n1004), .A2(KEYINPUT54), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n1000), .A2(new_n997), .ZN(new_n1069));
  OR3_X1    g644(.A1(new_n1008), .A2(new_n947), .A3(new_n1002), .ZN(new_n1070));
  OAI21_X1  g645(.A(new_n949), .B1(new_n977), .B2(KEYINPUT50), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n973), .A2(KEYINPUT50), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n1072), .A2(KEYINPUT118), .ZN(new_n1073));
  NAND3_X1  g648(.A1(new_n973), .A2(new_n971), .A3(KEYINPUT50), .ZN(new_n1074));
  AOI21_X1  g649(.A(new_n1071), .B1(new_n1073), .B2(new_n1074), .ZN(new_n1075));
  OAI211_X1 g650(.A(new_n1069), .B(new_n1070), .C1(new_n1075), .C2(G1961), .ZN(new_n1076));
  OAI21_X1  g651(.A(new_n1068), .B1(G171), .B2(new_n1076), .ZN(new_n1077));
  INV_X1    g652(.A(KEYINPUT126), .ZN(new_n1078));
  AND3_X1   g653(.A1(new_n1076), .A2(new_n1078), .A3(G171), .ZN(new_n1079));
  AOI21_X1  g654(.A(new_n1078), .B1(new_n1076), .B2(G171), .ZN(new_n1080));
  AND3_X1   g655(.A1(new_n1001), .A2(G301), .A3(new_n1003), .ZN(new_n1081));
  NOR3_X1   g656(.A1(new_n1079), .A2(new_n1080), .A3(new_n1081), .ZN(new_n1082));
  INV_X1    g657(.A(KEYINPUT54), .ZN(new_n1083));
  OAI21_X1  g658(.A(new_n1077), .B1(new_n1082), .B2(new_n1083), .ZN(new_n1084));
  NAND3_X1  g659(.A1(new_n1053), .A2(new_n993), .A3(new_n989), .ZN(new_n1085));
  AND2_X1   g660(.A1(new_n1025), .A2(new_n1030), .ZN(new_n1086));
  INV_X1    g661(.A(KEYINPUT57), .ZN(new_n1087));
  NAND2_X1  g662(.A1(G299), .A2(new_n1087), .ZN(new_n1088));
  NAND4_X1  g663(.A1(new_n571), .A2(KEYINPUT57), .A3(new_n572), .A4(new_n576), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n1088), .A2(new_n1089), .ZN(new_n1090));
  INV_X1    g665(.A(new_n1011), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n1013), .A2(new_n949), .ZN(new_n1092));
  OAI21_X1  g667(.A(new_n769), .B1(new_n1091), .B2(new_n1092), .ZN(new_n1093));
  XNOR2_X1  g668(.A(KEYINPUT56), .B(G2072), .ZN(new_n1094));
  NAND3_X1  g669(.A1(new_n998), .A2(new_n999), .A3(new_n1094), .ZN(new_n1095));
  AOI21_X1  g670(.A(new_n1090), .B1(new_n1093), .B2(new_n1095), .ZN(new_n1096));
  INV_X1    g671(.A(G1348), .ZN(new_n1097));
  NOR2_X1   g672(.A1(new_n977), .A2(new_n967), .ZN(new_n1098));
  AOI22_X1  g673(.A1(new_n996), .A2(new_n1097), .B1(new_n752), .B2(new_n1098), .ZN(new_n1099));
  AND3_X1   g674(.A1(new_n1093), .A2(new_n1090), .A3(new_n1095), .ZN(new_n1100));
  NOR2_X1   g675(.A1(new_n1099), .A2(new_n1100), .ZN(new_n1101));
  AOI21_X1  g676(.A(new_n1096), .B1(new_n1101), .B2(new_n609), .ZN(new_n1102));
  NOR3_X1   g677(.A1(new_n1008), .A2(G1996), .A3(new_n1009), .ZN(new_n1103));
  XNOR2_X1  g678(.A(KEYINPUT58), .B(G1341), .ZN(new_n1104));
  NOR2_X1   g679(.A1(new_n1098), .A2(new_n1104), .ZN(new_n1105));
  OAI21_X1  g680(.A(new_n561), .B1(new_n1103), .B2(new_n1105), .ZN(new_n1106));
  AND2_X1   g681(.A1(KEYINPUT122), .A2(KEYINPUT59), .ZN(new_n1107));
  XNOR2_X1  g682(.A(new_n1106), .B(new_n1107), .ZN(new_n1108));
  INV_X1    g683(.A(KEYINPUT60), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n608), .A2(new_n1109), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n1099), .A2(new_n1110), .ZN(new_n1111));
  NOR2_X1   g686(.A1(new_n608), .A2(new_n1109), .ZN(new_n1112));
  NAND2_X1  g687(.A1(new_n1111), .A2(new_n1112), .ZN(new_n1113));
  INV_X1    g688(.A(KEYINPUT123), .ZN(new_n1114));
  NOR2_X1   g689(.A1(new_n1114), .A2(KEYINPUT61), .ZN(new_n1115));
  OAI21_X1  g690(.A(new_n1115), .B1(new_n1100), .B2(new_n1096), .ZN(new_n1116));
  INV_X1    g691(.A(new_n1112), .ZN(new_n1117));
  NAND3_X1  g692(.A1(new_n1099), .A2(new_n1110), .A3(new_n1117), .ZN(new_n1118));
  NAND4_X1  g693(.A1(new_n1108), .A2(new_n1113), .A3(new_n1116), .A4(new_n1118), .ZN(new_n1119));
  OR2_X1    g694(.A1(new_n1100), .A2(new_n1096), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n1114), .A2(KEYINPUT61), .ZN(new_n1121));
  AOI21_X1  g696(.A(new_n1115), .B1(new_n1120), .B2(new_n1121), .ZN(new_n1122));
  OAI21_X1  g697(.A(new_n1102), .B1(new_n1119), .B2(new_n1122), .ZN(new_n1123));
  NAND4_X1  g698(.A1(new_n1084), .A2(new_n1085), .A3(new_n1086), .A4(new_n1123), .ZN(new_n1124));
  INV_X1    g699(.A(KEYINPUT63), .ZN(new_n1125));
  NAND4_X1  g700(.A1(new_n1025), .A2(new_n1125), .A3(G168), .A4(new_n982), .ZN(new_n1126));
  AND2_X1   g701(.A1(new_n1126), .A2(new_n1030), .ZN(new_n1127));
  AOI21_X1  g702(.A(new_n1067), .B1(new_n1124), .B2(new_n1127), .ZN(new_n1128));
  OAI21_X1  g703(.A(new_n963), .B1(new_n1066), .B2(new_n1128), .ZN(new_n1129));
  OR2_X1    g704(.A1(new_n957), .A2(new_n959), .ZN(new_n1130));
  NAND2_X1  g705(.A1(new_n749), .A2(new_n752), .ZN(new_n1131));
  AOI21_X1  g706(.A(new_n950), .B1(new_n1130), .B2(new_n1131), .ZN(new_n1132));
  AOI21_X1  g707(.A(new_n950), .B1(new_n953), .B2(new_n791), .ZN(new_n1133));
  AOI21_X1  g708(.A(KEYINPUT46), .B1(new_n951), .B2(new_n954), .ZN(new_n1134));
  AND3_X1   g709(.A1(new_n951), .A2(KEYINPUT46), .A3(new_n954), .ZN(new_n1135));
  NOR3_X1   g710(.A1(new_n1133), .A2(new_n1134), .A3(new_n1135), .ZN(new_n1136));
  XNOR2_X1  g711(.A(new_n1136), .B(KEYINPUT47), .ZN(new_n1137));
  NAND2_X1  g712(.A1(new_n961), .A2(new_n951), .ZN(new_n1138));
  NOR3_X1   g713(.A1(new_n950), .A2(G1986), .A3(G290), .ZN(new_n1139));
  XOR2_X1   g714(.A(new_n1139), .B(KEYINPUT48), .Z(new_n1140));
  AOI211_X1 g715(.A(new_n1132), .B(new_n1137), .C1(new_n1138), .C2(new_n1140), .ZN(new_n1141));
  NAND2_X1  g716(.A1(new_n1129), .A2(new_n1141), .ZN(G329));
  assign    G231 = 1'b0;
  AOI211_X1 g717(.A(new_n460), .B(G229), .C1(new_n939), .C2(new_n941), .ZN(new_n1144));
  NOR2_X1   g718(.A1(G401), .A2(G227), .ZN(new_n1145));
  AND3_X1   g719(.A1(new_n1144), .A2(new_n885), .A3(new_n1145), .ZN(G308));
  NAND3_X1  g720(.A1(new_n1144), .A2(new_n885), .A3(new_n1145), .ZN(G225));
endmodule


