//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 0 1 0 1 0 1 1 1 1 1 1 1 0 1 0 0 1 1 0 1 0 0 1 0 1 0 1 0 0 0 0 0 0 1 1 0 0 1 0 0 0 1 1 0 1 1 0 0 0 1 1 1 1 1 1 0 0 0 0 0 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:32:22 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n443, new_n444, new_n449, new_n453, new_n454, new_n455,
    new_n456, new_n457, new_n458, new_n461, new_n462, new_n463, new_n464,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n484, new_n485, new_n486,
    new_n487, new_n488, new_n489, new_n490, new_n491, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n533, new_n534, new_n535, new_n536, new_n537, new_n538,
    new_n539, new_n540, new_n541, new_n542, new_n543, new_n544, new_n545,
    new_n547, new_n548, new_n549, new_n550, new_n551, new_n552, new_n553,
    new_n554, new_n555, new_n556, new_n557, new_n558, new_n559, new_n560,
    new_n561, new_n562, new_n563, new_n564, new_n565, new_n566, new_n567,
    new_n568, new_n570, new_n571, new_n572, new_n573, new_n574, new_n575,
    new_n576, new_n577, new_n578, new_n579, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n590, new_n592,
    new_n593, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n611, new_n612, new_n613, new_n615, new_n616,
    new_n617, new_n619, new_n620, new_n621, new_n623, new_n624, new_n625,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n658,
    new_n661, new_n662, new_n664, new_n665, new_n667, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n687, new_n688, new_n689, new_n690, new_n691, new_n692,
    new_n693, new_n694, new_n695, new_n696, new_n697, new_n698, new_n699,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n706, new_n707,
    new_n708, new_n709, new_n710, new_n711, new_n712, new_n713, new_n714,
    new_n715, new_n716, new_n717, new_n718, new_n719, new_n720, new_n721,
    new_n723, new_n724, new_n725, new_n726, new_n727, new_n728, new_n729,
    new_n730, new_n731, new_n732, new_n733, new_n734, new_n735, new_n736,
    new_n737, new_n738, new_n739, new_n740, new_n741, new_n742, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n854, new_n855, new_n856,
    new_n857, new_n858, new_n859, new_n860, new_n861, new_n862, new_n863,
    new_n864, new_n865, new_n866, new_n867, new_n868, new_n869, new_n870,
    new_n871, new_n872, new_n873, new_n874, new_n875, new_n876, new_n877,
    new_n878, new_n879, new_n880, new_n881, new_n882, new_n883, new_n884,
    new_n885, new_n887, new_n888, new_n889, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n952, new_n953, new_n954, new_n955, new_n956, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1021, new_n1022, new_n1023, new_n1024, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1195;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  XNOR2_X1  g007(.A(KEYINPUT64), .B(G2066), .ZN(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  XNOR2_X1  g012(.A(KEYINPUT65), .B(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  INV_X1    g016(.A(G2072), .ZN(new_n442));
  INV_X1    g017(.A(G2078), .ZN(new_n443));
  NOR2_X1   g018(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  NAND3_X1  g019(.A1(new_n444), .A2(G2084), .A3(G2090), .ZN(G158));
  NAND3_X1  g020(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g021(.A(G452), .Z(G391));
  AND2_X1   g022(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g023(.A1(G7), .A2(G661), .ZN(new_n449));
  XOR2_X1   g024(.A(new_n449), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g025(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g026(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g027(.A1(G235), .A2(G237), .A3(G238), .A4(G236), .ZN(new_n453));
  XOR2_X1   g028(.A(new_n453), .B(KEYINPUT66), .Z(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR4_X1   g030(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n456));
  XNOR2_X1  g031(.A(new_n456), .B(KEYINPUT2), .ZN(new_n457));
  INV_X1    g032(.A(new_n457), .ZN(new_n458));
  NOR2_X1   g033(.A1(new_n455), .A2(new_n458), .ZN(G325));
  INV_X1    g034(.A(G325), .ZN(G261));
  AOI21_X1  g035(.A(KEYINPUT67), .B1(new_n455), .B2(G567), .ZN(new_n461));
  AOI21_X1  g036(.A(new_n461), .B1(G2106), .B2(new_n458), .ZN(new_n462));
  NAND3_X1  g037(.A1(new_n455), .A2(KEYINPUT67), .A3(G567), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  INV_X1    g039(.A(new_n464), .ZN(G319));
  NAND2_X1  g040(.A1(G101), .A2(G2104), .ZN(new_n466));
  INV_X1    g041(.A(G2104), .ZN(new_n467));
  NOR2_X1   g042(.A1(new_n467), .A2(KEYINPUT3), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n468), .A2(KEYINPUT69), .ZN(new_n469));
  INV_X1    g044(.A(KEYINPUT69), .ZN(new_n470));
  AOI21_X1  g045(.A(new_n470), .B1(KEYINPUT3), .B2(new_n467), .ZN(new_n471));
  OAI21_X1  g046(.A(new_n469), .B1(new_n468), .B2(new_n471), .ZN(new_n472));
  INV_X1    g047(.A(G137), .ZN(new_n473));
  OAI21_X1  g048(.A(new_n466), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  INV_X1    g049(.A(G2105), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n476), .A2(KEYINPUT70), .ZN(new_n477));
  INV_X1    g052(.A(KEYINPUT70), .ZN(new_n478));
  NAND3_X1  g053(.A1(new_n474), .A2(new_n478), .A3(new_n475), .ZN(new_n479));
  INV_X1    g054(.A(G125), .ZN(new_n480));
  INV_X1    g055(.A(KEYINPUT3), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n481), .A2(G2104), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n467), .A2(KEYINPUT3), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n484), .A2(KEYINPUT68), .ZN(new_n485));
  INV_X1    g060(.A(KEYINPUT68), .ZN(new_n486));
  NAND3_X1  g061(.A1(new_n482), .A2(new_n483), .A3(new_n486), .ZN(new_n487));
  AOI21_X1  g062(.A(new_n480), .B1(new_n485), .B2(new_n487), .ZN(new_n488));
  AND2_X1   g063(.A1(G113), .A2(G2104), .ZN(new_n489));
  OAI21_X1  g064(.A(G2105), .B1(new_n488), .B2(new_n489), .ZN(new_n490));
  NAND3_X1  g065(.A1(new_n477), .A2(new_n479), .A3(new_n490), .ZN(new_n491));
  INV_X1    g066(.A(new_n491), .ZN(G160));
  OR2_X1    g067(.A1(G100), .A2(G2105), .ZN(new_n493));
  OAI211_X1 g068(.A(new_n493), .B(G2104), .C1(G112), .C2(new_n475), .ZN(new_n494));
  OR2_X1    g069(.A1(new_n472), .A2(KEYINPUT71), .ZN(new_n495));
  NAND2_X1  g070(.A1(new_n472), .A2(KEYINPUT71), .ZN(new_n496));
  NAND3_X1  g071(.A1(new_n495), .A2(G2105), .A3(new_n496), .ZN(new_n497));
  INV_X1    g072(.A(G124), .ZN(new_n498));
  INV_X1    g073(.A(G136), .ZN(new_n499));
  NAND3_X1  g074(.A1(new_n495), .A2(new_n475), .A3(new_n496), .ZN(new_n500));
  OAI221_X1 g075(.A(new_n494), .B1(new_n497), .B2(new_n498), .C1(new_n499), .C2(new_n500), .ZN(new_n501));
  XNOR2_X1  g076(.A(new_n501), .B(KEYINPUT72), .ZN(new_n502));
  INV_X1    g077(.A(new_n502), .ZN(G162));
  NAND2_X1  g078(.A1(new_n475), .A2(G138), .ZN(new_n504));
  AOI21_X1  g079(.A(new_n504), .B1(new_n485), .B2(new_n487), .ZN(new_n505));
  NOR2_X1   g080(.A1(new_n505), .A2(KEYINPUT4), .ZN(new_n506));
  INV_X1    g081(.A(KEYINPUT73), .ZN(new_n507));
  OR3_X1    g082(.A1(new_n507), .A2(new_n475), .A3(G114), .ZN(new_n508));
  OAI21_X1  g083(.A(new_n507), .B1(new_n475), .B2(G114), .ZN(new_n509));
  OR2_X1    g084(.A1(G102), .A2(G2105), .ZN(new_n510));
  NAND4_X1  g085(.A1(new_n508), .A2(G2104), .A3(new_n509), .A4(new_n510), .ZN(new_n511));
  INV_X1    g086(.A(new_n504), .ZN(new_n512));
  AOI22_X1  g087(.A1(new_n512), .A2(KEYINPUT4), .B1(G126), .B2(G2105), .ZN(new_n513));
  OAI21_X1  g088(.A(new_n511), .B1(new_n472), .B2(new_n513), .ZN(new_n514));
  NOR2_X1   g089(.A1(new_n506), .A2(new_n514), .ZN(G164));
  INV_X1    g090(.A(G651), .ZN(new_n516));
  INV_X1    g091(.A(G543), .ZN(new_n517));
  OAI21_X1  g092(.A(KEYINPUT76), .B1(new_n517), .B2(KEYINPUT5), .ZN(new_n518));
  XNOR2_X1  g093(.A(KEYINPUT75), .B(G543), .ZN(new_n519));
  INV_X1    g094(.A(KEYINPUT5), .ZN(new_n520));
  OAI21_X1  g095(.A(new_n518), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  AND2_X1   g096(.A1(new_n517), .A2(KEYINPUT75), .ZN(new_n522));
  NOR2_X1   g097(.A1(new_n517), .A2(KEYINPUT75), .ZN(new_n523));
  OAI211_X1 g098(.A(KEYINPUT76), .B(KEYINPUT5), .C1(new_n522), .C2(new_n523), .ZN(new_n524));
  NAND3_X1  g099(.A1(new_n521), .A2(G62), .A3(new_n524), .ZN(new_n525));
  INV_X1    g100(.A(KEYINPUT77), .ZN(new_n526));
  AOI22_X1  g101(.A1(new_n525), .A2(new_n526), .B1(G75), .B2(G543), .ZN(new_n527));
  AND2_X1   g102(.A1(new_n521), .A2(new_n524), .ZN(new_n528));
  NAND3_X1  g103(.A1(new_n528), .A2(KEYINPUT77), .A3(G62), .ZN(new_n529));
  AOI21_X1  g104(.A(new_n516), .B1(new_n527), .B2(new_n529), .ZN(new_n530));
  INV_X1    g105(.A(KEYINPUT78), .ZN(new_n531));
  NAND2_X1  g106(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  INV_X1    g107(.A(new_n532), .ZN(new_n533));
  NAND2_X1  g108(.A1(G50), .A2(G543), .ZN(new_n534));
  NAND2_X1  g109(.A1(new_n521), .A2(new_n524), .ZN(new_n535));
  INV_X1    g110(.A(G88), .ZN(new_n536));
  OAI21_X1  g111(.A(new_n534), .B1(new_n535), .B2(new_n536), .ZN(new_n537));
  NOR2_X1   g112(.A1(new_n516), .A2(KEYINPUT6), .ZN(new_n538));
  INV_X1    g113(.A(KEYINPUT6), .ZN(new_n539));
  OAI21_X1  g114(.A(KEYINPUT74), .B1(new_n539), .B2(G651), .ZN(new_n540));
  INV_X1    g115(.A(KEYINPUT74), .ZN(new_n541));
  NAND3_X1  g116(.A1(new_n541), .A2(new_n516), .A3(KEYINPUT6), .ZN(new_n542));
  AOI21_X1  g117(.A(new_n538), .B1(new_n540), .B2(new_n542), .ZN(new_n543));
  NAND2_X1  g118(.A1(new_n537), .A2(new_n543), .ZN(new_n544));
  OAI21_X1  g119(.A(new_n544), .B1(new_n530), .B2(new_n531), .ZN(new_n545));
  NOR2_X1   g120(.A1(new_n533), .A2(new_n545), .ZN(G166));
  NAND3_X1  g121(.A1(new_n528), .A2(G89), .A3(new_n543), .ZN(new_n547));
  XOR2_X1   g122(.A(KEYINPUT81), .B(KEYINPUT7), .Z(new_n548));
  NAND3_X1  g123(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n549));
  XNOR2_X1  g124(.A(new_n548), .B(new_n549), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n547), .A2(new_n550), .ZN(new_n551));
  INV_X1    g126(.A(KEYINPUT79), .ZN(new_n552));
  OAI21_X1  g127(.A(G543), .B1(new_n543), .B2(new_n552), .ZN(new_n553));
  AOI211_X1 g128(.A(KEYINPUT79), .B(new_n538), .C1(new_n540), .C2(new_n542), .ZN(new_n554));
  INV_X1    g129(.A(G51), .ZN(new_n555));
  NOR3_X1   g130(.A1(new_n553), .A2(new_n554), .A3(new_n555), .ZN(new_n556));
  NAND4_X1  g131(.A1(new_n521), .A2(new_n524), .A3(G63), .A4(G651), .ZN(new_n557));
  INV_X1    g132(.A(new_n557), .ZN(new_n558));
  OAI21_X1  g133(.A(KEYINPUT80), .B1(new_n556), .B2(new_n558), .ZN(new_n559));
  INV_X1    g134(.A(new_n538), .ZN(new_n560));
  AOI21_X1  g135(.A(new_n541), .B1(KEYINPUT6), .B2(new_n516), .ZN(new_n561));
  NOR3_X1   g136(.A1(new_n539), .A2(KEYINPUT74), .A3(G651), .ZN(new_n562));
  OAI21_X1  g137(.A(new_n560), .B1(new_n561), .B2(new_n562), .ZN(new_n563));
  AOI21_X1  g138(.A(new_n517), .B1(new_n563), .B2(KEYINPUT79), .ZN(new_n564));
  NAND2_X1  g139(.A1(new_n543), .A2(new_n552), .ZN(new_n565));
  NAND3_X1  g140(.A1(new_n564), .A2(G51), .A3(new_n565), .ZN(new_n566));
  INV_X1    g141(.A(KEYINPUT80), .ZN(new_n567));
  NAND3_X1  g142(.A1(new_n566), .A2(new_n567), .A3(new_n557), .ZN(new_n568));
  AOI21_X1  g143(.A(new_n551), .B1(new_n559), .B2(new_n568), .ZN(G168));
  NAND2_X1  g144(.A1(new_n563), .A2(KEYINPUT79), .ZN(new_n570));
  NAND4_X1  g145(.A1(new_n570), .A2(G52), .A3(new_n565), .A4(G543), .ZN(new_n571));
  NAND4_X1  g146(.A1(new_n521), .A2(new_n524), .A3(new_n543), .A4(G90), .ZN(new_n572));
  NAND2_X1  g147(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  INV_X1    g148(.A(KEYINPUT82), .ZN(new_n574));
  NAND2_X1  g149(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  NAND3_X1  g150(.A1(new_n571), .A2(KEYINPUT82), .A3(new_n572), .ZN(new_n576));
  NAND2_X1  g151(.A1(G77), .A2(G543), .ZN(new_n577));
  INV_X1    g152(.A(G64), .ZN(new_n578));
  OAI21_X1  g153(.A(new_n577), .B1(new_n535), .B2(new_n578), .ZN(new_n579));
  AOI22_X1  g154(.A1(new_n575), .A2(new_n576), .B1(G651), .B2(new_n579), .ZN(G171));
  XOR2_X1   g155(.A(KEYINPUT83), .B(G43), .Z(new_n581));
  NOR3_X1   g156(.A1(new_n553), .A2(new_n554), .A3(new_n581), .ZN(new_n582));
  NAND3_X1  g157(.A1(new_n521), .A2(G56), .A3(new_n524), .ZN(new_n583));
  NAND2_X1  g158(.A1(G68), .A2(G543), .ZN(new_n584));
  AOI21_X1  g159(.A(new_n516), .B1(new_n583), .B2(new_n584), .ZN(new_n585));
  INV_X1    g160(.A(G81), .ZN(new_n586));
  NOR3_X1   g161(.A1(new_n535), .A2(new_n586), .A3(new_n563), .ZN(new_n587));
  NOR3_X1   g162(.A1(new_n582), .A2(new_n585), .A3(new_n587), .ZN(new_n588));
  NAND2_X1  g163(.A1(new_n588), .A2(G860), .ZN(G153));
  AND3_X1   g164(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n590));
  NAND2_X1  g165(.A1(new_n590), .A2(G36), .ZN(G176));
  NAND2_X1  g166(.A1(G1), .A2(G3), .ZN(new_n592));
  XNOR2_X1  g167(.A(new_n592), .B(KEYINPUT8), .ZN(new_n593));
  NAND2_X1  g168(.A1(new_n590), .A2(new_n593), .ZN(G188));
  INV_X1    g169(.A(KEYINPUT85), .ZN(new_n595));
  NAND3_X1  g170(.A1(new_n521), .A2(G65), .A3(new_n524), .ZN(new_n596));
  NAND2_X1  g171(.A1(G78), .A2(G543), .ZN(new_n597));
  NAND2_X1  g172(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  AOI21_X1  g173(.A(new_n595), .B1(new_n598), .B2(G651), .ZN(new_n599));
  AOI211_X1 g174(.A(KEYINPUT85), .B(new_n516), .C1(new_n596), .C2(new_n597), .ZN(new_n600));
  OR2_X1    g175(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  NAND4_X1  g176(.A1(new_n570), .A2(G53), .A3(new_n565), .A4(G543), .ZN(new_n602));
  INV_X1    g177(.A(KEYINPUT84), .ZN(new_n603));
  NAND3_X1  g178(.A1(new_n602), .A2(new_n603), .A3(KEYINPUT9), .ZN(new_n604));
  NOR2_X1   g179(.A1(new_n553), .A2(new_n554), .ZN(new_n605));
  NAND2_X1  g180(.A1(new_n603), .A2(KEYINPUT9), .ZN(new_n606));
  NAND3_X1  g181(.A1(new_n605), .A2(G53), .A3(new_n606), .ZN(new_n607));
  NOR2_X1   g182(.A1(new_n535), .A2(new_n563), .ZN(new_n608));
  AOI22_X1  g183(.A1(new_n604), .A2(new_n607), .B1(G91), .B2(new_n608), .ZN(new_n609));
  NAND2_X1  g184(.A1(new_n601), .A2(new_n609), .ZN(G299));
  NAND2_X1  g185(.A1(new_n579), .A2(G651), .ZN(new_n611));
  AND3_X1   g186(.A1(new_n571), .A2(KEYINPUT82), .A3(new_n572), .ZN(new_n612));
  AOI21_X1  g187(.A(KEYINPUT82), .B1(new_n571), .B2(new_n572), .ZN(new_n613));
  OAI21_X1  g188(.A(new_n611), .B1(new_n612), .B2(new_n613), .ZN(G301));
  INV_X1    g189(.A(new_n551), .ZN(new_n615));
  NOR3_X1   g190(.A1(new_n556), .A2(new_n558), .A3(KEYINPUT80), .ZN(new_n616));
  AOI21_X1  g191(.A(new_n567), .B1(new_n566), .B2(new_n557), .ZN(new_n617));
  OAI21_X1  g192(.A(new_n615), .B1(new_n616), .B2(new_n617), .ZN(G286));
  NAND2_X1  g193(.A1(new_n527), .A2(new_n529), .ZN(new_n619));
  NAND2_X1  g194(.A1(new_n619), .A2(G651), .ZN(new_n620));
  AOI22_X1  g195(.A1(new_n620), .A2(KEYINPUT78), .B1(new_n543), .B2(new_n537), .ZN(new_n621));
  NAND2_X1  g196(.A1(new_n621), .A2(new_n532), .ZN(G303));
  NAND2_X1  g197(.A1(new_n605), .A2(G49), .ZN(new_n623));
  NAND2_X1  g198(.A1(new_n608), .A2(G87), .ZN(new_n624));
  OAI21_X1  g199(.A(G651), .B1(new_n528), .B2(G74), .ZN(new_n625));
  NAND3_X1  g200(.A1(new_n623), .A2(new_n624), .A3(new_n625), .ZN(G288));
  NAND2_X1  g201(.A1(G48), .A2(G543), .ZN(new_n627));
  INV_X1    g202(.A(G86), .ZN(new_n628));
  OAI21_X1  g203(.A(new_n627), .B1(new_n535), .B2(new_n628), .ZN(new_n629));
  NAND2_X1  g204(.A1(new_n629), .A2(new_n543), .ZN(new_n630));
  NAND2_X1  g205(.A1(G73), .A2(G543), .ZN(new_n631));
  INV_X1    g206(.A(G61), .ZN(new_n632));
  OAI21_X1  g207(.A(new_n631), .B1(new_n535), .B2(new_n632), .ZN(new_n633));
  AND3_X1   g208(.A1(new_n633), .A2(KEYINPUT86), .A3(G651), .ZN(new_n634));
  AOI21_X1  g209(.A(KEYINPUT86), .B1(new_n633), .B2(G651), .ZN(new_n635));
  OAI21_X1  g210(.A(new_n630), .B1(new_n634), .B2(new_n635), .ZN(G305));
  NAND2_X1  g211(.A1(G72), .A2(G543), .ZN(new_n637));
  INV_X1    g212(.A(G60), .ZN(new_n638));
  OAI21_X1  g213(.A(new_n637), .B1(new_n535), .B2(new_n638), .ZN(new_n639));
  NAND2_X1  g214(.A1(new_n639), .A2(G651), .ZN(new_n640));
  NAND2_X1  g215(.A1(new_n605), .A2(G47), .ZN(new_n641));
  NAND2_X1  g216(.A1(new_n608), .A2(G85), .ZN(new_n642));
  NAND3_X1  g217(.A1(new_n640), .A2(new_n641), .A3(new_n642), .ZN(G290));
  NAND2_X1  g218(.A1(G79), .A2(G543), .ZN(new_n644));
  INV_X1    g219(.A(G66), .ZN(new_n645));
  OAI21_X1  g220(.A(new_n644), .B1(new_n535), .B2(new_n645), .ZN(new_n646));
  NAND2_X1  g221(.A1(new_n646), .A2(G651), .ZN(new_n647));
  NAND2_X1  g222(.A1(new_n605), .A2(G54), .ZN(new_n648));
  NAND4_X1  g223(.A1(new_n521), .A2(new_n524), .A3(new_n543), .A4(G92), .ZN(new_n649));
  INV_X1    g224(.A(KEYINPUT10), .ZN(new_n650));
  AND2_X1   g225(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  NOR2_X1   g226(.A1(new_n649), .A2(new_n650), .ZN(new_n652));
  OAI211_X1 g227(.A(new_n647), .B(new_n648), .C1(new_n651), .C2(new_n652), .ZN(new_n653));
  INV_X1    g228(.A(G868), .ZN(new_n654));
  NAND2_X1  g229(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  OAI21_X1  g230(.A(new_n655), .B1(G171), .B2(new_n654), .ZN(G321));
  XOR2_X1   g231(.A(G321), .B(KEYINPUT87), .Z(G284));
  NAND2_X1  g232(.A1(G299), .A2(new_n654), .ZN(new_n658));
  OAI21_X1  g233(.A(new_n658), .B1(new_n654), .B2(G168), .ZN(G297));
  OAI21_X1  g234(.A(new_n658), .B1(new_n654), .B2(G168), .ZN(G280));
  INV_X1    g235(.A(new_n653), .ZN(new_n661));
  INV_X1    g236(.A(G559), .ZN(new_n662));
  OAI21_X1  g237(.A(new_n661), .B1(new_n662), .B2(G860), .ZN(G148));
  NAND2_X1  g238(.A1(new_n661), .A2(new_n662), .ZN(new_n664));
  NAND2_X1  g239(.A1(new_n664), .A2(G868), .ZN(new_n665));
  OAI21_X1  g240(.A(new_n665), .B1(G868), .B2(new_n588), .ZN(G323));
  XNOR2_X1  g241(.A(KEYINPUT88), .B(KEYINPUT11), .ZN(new_n667));
  XNOR2_X1  g242(.A(G323), .B(new_n667), .ZN(G282));
  INV_X1    g243(.A(new_n500), .ZN(new_n669));
  NAND2_X1  g244(.A1(new_n669), .A2(G135), .ZN(new_n670));
  OR2_X1    g245(.A1(G99), .A2(G2105), .ZN(new_n671));
  OAI211_X1 g246(.A(new_n671), .B(G2104), .C1(G111), .C2(new_n475), .ZN(new_n672));
  NAND2_X1  g247(.A1(new_n670), .A2(new_n672), .ZN(new_n673));
  INV_X1    g248(.A(new_n497), .ZN(new_n674));
  AOI21_X1  g249(.A(new_n673), .B1(G123), .B2(new_n674), .ZN(new_n675));
  XNOR2_X1  g250(.A(new_n675), .B(G2096), .ZN(new_n676));
  NAND2_X1  g251(.A1(new_n485), .A2(new_n487), .ZN(new_n677));
  NOR2_X1   g252(.A1(new_n467), .A2(G2105), .ZN(new_n678));
  NAND2_X1  g253(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  XNOR2_X1  g254(.A(new_n679), .B(KEYINPUT12), .ZN(new_n680));
  INV_X1    g255(.A(KEYINPUT13), .ZN(new_n681));
  AOI22_X1  g256(.A1(new_n680), .A2(new_n681), .B1(KEYINPUT89), .B2(G2100), .ZN(new_n682));
  OAI21_X1  g257(.A(new_n682), .B1(new_n681), .B2(new_n680), .ZN(new_n683));
  NOR2_X1   g258(.A1(KEYINPUT89), .A2(G2100), .ZN(new_n684));
  XNOR2_X1  g259(.A(new_n683), .B(new_n684), .ZN(new_n685));
  NAND2_X1  g260(.A1(new_n676), .A2(new_n685), .ZN(G156));
  XNOR2_X1  g261(.A(KEYINPUT15), .B(G2435), .ZN(new_n687));
  XNOR2_X1  g262(.A(KEYINPUT91), .B(G2438), .ZN(new_n688));
  XNOR2_X1  g263(.A(new_n687), .B(new_n688), .ZN(new_n689));
  XOR2_X1   g264(.A(G2427), .B(G2430), .Z(new_n690));
  OR2_X1    g265(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  NAND2_X1  g266(.A1(new_n689), .A2(new_n690), .ZN(new_n692));
  NAND3_X1  g267(.A1(new_n691), .A2(KEYINPUT14), .A3(new_n692), .ZN(new_n693));
  XOR2_X1   g268(.A(G2443), .B(G2446), .Z(new_n694));
  XNOR2_X1  g269(.A(new_n693), .B(new_n694), .ZN(new_n695));
  XNOR2_X1  g270(.A(KEYINPUT90), .B(KEYINPUT16), .ZN(new_n696));
  XNOR2_X1  g271(.A(G2451), .B(G2454), .ZN(new_n697));
  XOR2_X1   g272(.A(new_n696), .B(new_n697), .Z(new_n698));
  XNOR2_X1  g273(.A(new_n695), .B(new_n698), .ZN(new_n699));
  XOR2_X1   g274(.A(G1341), .B(G1348), .Z(new_n700));
  INV_X1    g275(.A(new_n700), .ZN(new_n701));
  NAND2_X1  g276(.A1(new_n699), .A2(new_n701), .ZN(new_n702));
  NOR2_X1   g277(.A1(new_n699), .A2(new_n701), .ZN(new_n703));
  OAI211_X1 g278(.A(G14), .B(new_n702), .C1(new_n703), .C2(KEYINPUT92), .ZN(new_n704));
  AOI21_X1  g279(.A(new_n704), .B1(KEYINPUT92), .B2(new_n703), .ZN(G401));
  XOR2_X1   g280(.A(G2084), .B(G2090), .Z(new_n706));
  INV_X1    g281(.A(new_n706), .ZN(new_n707));
  XOR2_X1   g282(.A(G2067), .B(G2678), .Z(new_n708));
  OR2_X1    g283(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  NOR2_X1   g284(.A1(G2072), .A2(G2078), .ZN(new_n710));
  NOR2_X1   g285(.A1(new_n444), .A2(new_n710), .ZN(new_n711));
  NOR2_X1   g286(.A1(new_n709), .A2(new_n711), .ZN(new_n712));
  XNOR2_X1  g287(.A(new_n712), .B(KEYINPUT18), .ZN(new_n713));
  XNOR2_X1  g288(.A(new_n711), .B(KEYINPUT17), .ZN(new_n714));
  NAND2_X1  g289(.A1(new_n707), .A2(new_n708), .ZN(new_n715));
  NAND3_X1  g290(.A1(new_n714), .A2(new_n709), .A3(new_n715), .ZN(new_n716));
  INV_X1    g291(.A(new_n711), .ZN(new_n717));
  AOI21_X1  g292(.A(new_n715), .B1(KEYINPUT93), .B2(new_n717), .ZN(new_n718));
  OAI21_X1  g293(.A(new_n718), .B1(KEYINPUT93), .B2(new_n717), .ZN(new_n719));
  NAND3_X1  g294(.A1(new_n713), .A2(new_n716), .A3(new_n719), .ZN(new_n720));
  XOR2_X1   g295(.A(G2096), .B(G2100), .Z(new_n721));
  XNOR2_X1  g296(.A(new_n720), .B(new_n721), .ZN(G227));
  XNOR2_X1  g297(.A(G1956), .B(G2474), .ZN(new_n723));
  XNOR2_X1  g298(.A(new_n723), .B(KEYINPUT95), .ZN(new_n724));
  XOR2_X1   g299(.A(G1961), .B(G1966), .Z(new_n725));
  NAND2_X1  g300(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  XNOR2_X1  g301(.A(G1971), .B(G1976), .ZN(new_n727));
  XNOR2_X1  g302(.A(KEYINPUT94), .B(KEYINPUT19), .ZN(new_n728));
  XOR2_X1   g303(.A(new_n727), .B(new_n728), .Z(new_n729));
  NOR2_X1   g304(.A1(new_n726), .A2(new_n729), .ZN(new_n730));
  NOR2_X1   g305(.A1(new_n724), .A2(new_n725), .ZN(new_n731));
  INV_X1    g306(.A(new_n729), .ZN(new_n732));
  AOI22_X1  g307(.A1(new_n730), .A2(KEYINPUT20), .B1(new_n731), .B2(new_n732), .ZN(new_n733));
  INV_X1    g308(.A(new_n731), .ZN(new_n734));
  NAND3_X1  g309(.A1(new_n734), .A2(new_n729), .A3(new_n726), .ZN(new_n735));
  OAI211_X1 g310(.A(new_n733), .B(new_n735), .C1(KEYINPUT20), .C2(new_n730), .ZN(new_n736));
  XOR2_X1   g311(.A(G1991), .B(G1996), .Z(new_n737));
  XNOR2_X1  g312(.A(G1981), .B(G1986), .ZN(new_n738));
  XNOR2_X1  g313(.A(new_n737), .B(new_n738), .ZN(new_n739));
  XNOR2_X1  g314(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n740));
  XNOR2_X1  g315(.A(new_n740), .B(KEYINPUT96), .ZN(new_n741));
  XNOR2_X1  g316(.A(new_n739), .B(new_n741), .ZN(new_n742));
  XNOR2_X1  g317(.A(new_n736), .B(new_n742), .ZN(G229));
  INV_X1    g318(.A(G16), .ZN(new_n744));
  NAND2_X1  g319(.A1(new_n744), .A2(G4), .ZN(new_n745));
  OAI21_X1  g320(.A(new_n745), .B1(new_n661), .B2(new_n744), .ZN(new_n746));
  XOR2_X1   g321(.A(KEYINPUT100), .B(G1348), .Z(new_n747));
  XNOR2_X1  g322(.A(new_n746), .B(new_n747), .ZN(new_n748));
  INV_X1    g323(.A(G1341), .ZN(new_n749));
  NAND2_X1  g324(.A1(new_n588), .A2(G16), .ZN(new_n750));
  OAI21_X1  g325(.A(new_n750), .B1(G16), .B2(G19), .ZN(new_n751));
  INV_X1    g326(.A(G1961), .ZN(new_n752));
  NOR2_X1   g327(.A1(G5), .A2(G16), .ZN(new_n753));
  AOI21_X1  g328(.A(new_n753), .B1(G171), .B2(G16), .ZN(new_n754));
  INV_X1    g329(.A(new_n754), .ZN(new_n755));
  OAI221_X1 g330(.A(new_n748), .B1(new_n749), .B2(new_n751), .C1(new_n752), .C2(new_n755), .ZN(new_n756));
  INV_X1    g331(.A(G1966), .ZN(new_n757));
  NAND2_X1  g332(.A1(G168), .A2(G16), .ZN(new_n758));
  OAI21_X1  g333(.A(new_n758), .B1(G16), .B2(G21), .ZN(new_n759));
  AOI21_X1  g334(.A(new_n756), .B1(new_n757), .B2(new_n759), .ZN(new_n760));
  NOR2_X1   g335(.A1(new_n759), .A2(new_n757), .ZN(new_n761));
  XOR2_X1   g336(.A(new_n761), .B(KEYINPUT103), .Z(new_n762));
  NAND2_X1  g337(.A1(new_n755), .A2(new_n752), .ZN(new_n763));
  INV_X1    g338(.A(KEYINPUT24), .ZN(new_n764));
  INV_X1    g339(.A(G34), .ZN(new_n765));
  AOI21_X1  g340(.A(G29), .B1(new_n764), .B2(new_n765), .ZN(new_n766));
  OAI21_X1  g341(.A(new_n766), .B1(new_n764), .B2(new_n765), .ZN(new_n767));
  INV_X1    g342(.A(G29), .ZN(new_n768));
  OAI21_X1  g343(.A(new_n767), .B1(G160), .B2(new_n768), .ZN(new_n769));
  NAND2_X1  g344(.A1(new_n669), .A2(G141), .ZN(new_n770));
  NAND2_X1  g345(.A1(new_n674), .A2(G129), .ZN(new_n771));
  NAND3_X1  g346(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n772));
  INV_X1    g347(.A(KEYINPUT26), .ZN(new_n773));
  OR2_X1    g348(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  NAND2_X1  g349(.A1(new_n772), .A2(new_n773), .ZN(new_n775));
  AOI22_X1  g350(.A1(new_n774), .A2(new_n775), .B1(G105), .B2(new_n678), .ZN(new_n776));
  NAND3_X1  g351(.A1(new_n770), .A2(new_n771), .A3(new_n776), .ZN(new_n777));
  INV_X1    g352(.A(new_n777), .ZN(new_n778));
  NAND2_X1  g353(.A1(new_n778), .A2(G29), .ZN(new_n779));
  OAI21_X1  g354(.A(new_n779), .B1(G29), .B2(G32), .ZN(new_n780));
  XOR2_X1   g355(.A(KEYINPUT27), .B(G1996), .Z(new_n781));
  INV_X1    g356(.A(new_n781), .ZN(new_n782));
  OAI221_X1 g357(.A(new_n763), .B1(G2084), .B2(new_n769), .C1(new_n780), .C2(new_n782), .ZN(new_n783));
  INV_X1    g358(.A(KEYINPUT104), .ZN(new_n784));
  OR2_X1    g359(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  NAND2_X1  g360(.A1(new_n783), .A2(new_n784), .ZN(new_n786));
  NAND4_X1  g361(.A1(new_n760), .A2(new_n762), .A3(new_n785), .A4(new_n786), .ZN(new_n787));
  OR2_X1    g362(.A1(G29), .A2(G33), .ZN(new_n788));
  AOI22_X1  g363(.A1(new_n677), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n789));
  INV_X1    g364(.A(KEYINPUT102), .ZN(new_n790));
  AOI21_X1  g365(.A(new_n475), .B1(new_n789), .B2(new_n790), .ZN(new_n791));
  OAI21_X1  g366(.A(new_n791), .B1(new_n790), .B2(new_n789), .ZN(new_n792));
  NAND2_X1  g367(.A1(new_n669), .A2(G139), .ZN(new_n793));
  NAND2_X1  g368(.A1(new_n678), .A2(G103), .ZN(new_n794));
  XOR2_X1   g369(.A(new_n794), .B(KEYINPUT25), .Z(new_n795));
  NAND3_X1  g370(.A1(new_n792), .A2(new_n793), .A3(new_n795), .ZN(new_n796));
  OAI21_X1  g371(.A(new_n788), .B1(new_n796), .B2(new_n768), .ZN(new_n797));
  AOI22_X1  g372(.A1(new_n780), .A2(new_n782), .B1(new_n442), .B2(new_n797), .ZN(new_n798));
  OR2_X1    g373(.A1(new_n797), .A2(new_n442), .ZN(new_n799));
  NAND2_X1  g374(.A1(new_n675), .A2(G29), .ZN(new_n800));
  NAND2_X1  g375(.A1(new_n768), .A2(G27), .ZN(new_n801));
  OAI21_X1  g376(.A(new_n801), .B1(G164), .B2(new_n768), .ZN(new_n802));
  XNOR2_X1  g377(.A(new_n802), .B(new_n443), .ZN(new_n803));
  XOR2_X1   g378(.A(KEYINPUT31), .B(G11), .Z(new_n804));
  INV_X1    g379(.A(G28), .ZN(new_n805));
  OR2_X1    g380(.A1(new_n805), .A2(KEYINPUT30), .ZN(new_n806));
  AOI21_X1  g381(.A(G29), .B1(new_n805), .B2(KEYINPUT30), .ZN(new_n807));
  AOI21_X1  g382(.A(new_n804), .B1(new_n806), .B2(new_n807), .ZN(new_n808));
  AND3_X1   g383(.A1(new_n800), .A2(new_n803), .A3(new_n808), .ZN(new_n809));
  AOI22_X1  g384(.A1(new_n751), .A2(new_n749), .B1(new_n769), .B2(G2084), .ZN(new_n810));
  NAND4_X1  g385(.A1(new_n798), .A2(new_n799), .A3(new_n809), .A4(new_n810), .ZN(new_n811));
  AND2_X1   g386(.A1(new_n768), .A2(G35), .ZN(new_n812));
  AOI21_X1  g387(.A(new_n812), .B1(new_n502), .B2(G29), .ZN(new_n813));
  XOR2_X1   g388(.A(KEYINPUT29), .B(G2090), .Z(new_n814));
  INV_X1    g389(.A(new_n814), .ZN(new_n815));
  OR2_X1    g390(.A1(new_n813), .A2(new_n815), .ZN(new_n816));
  NAND2_X1  g391(.A1(new_n813), .A2(new_n815), .ZN(new_n817));
  AOI21_X1  g392(.A(new_n811), .B1(new_n816), .B2(new_n817), .ZN(new_n818));
  INV_X1    g393(.A(KEYINPUT28), .ZN(new_n819));
  INV_X1    g394(.A(G26), .ZN(new_n820));
  OAI21_X1  g395(.A(new_n819), .B1(new_n820), .B2(G29), .ZN(new_n821));
  NOR2_X1   g396(.A1(new_n820), .A2(G29), .ZN(new_n822));
  NAND2_X1  g397(.A1(new_n674), .A2(G128), .ZN(new_n823));
  NAND2_X1  g398(.A1(new_n669), .A2(G140), .ZN(new_n824));
  OR2_X1    g399(.A1(G104), .A2(G2105), .ZN(new_n825));
  OAI211_X1 g400(.A(new_n825), .B(G2104), .C1(G116), .C2(new_n475), .ZN(new_n826));
  NAND3_X1  g401(.A1(new_n823), .A2(new_n824), .A3(new_n826), .ZN(new_n827));
  INV_X1    g402(.A(KEYINPUT101), .ZN(new_n828));
  NAND2_X1  g403(.A1(new_n827), .A2(new_n828), .ZN(new_n829));
  NAND4_X1  g404(.A1(new_n823), .A2(new_n824), .A3(KEYINPUT101), .A4(new_n826), .ZN(new_n830));
  NAND2_X1  g405(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  AOI21_X1  g406(.A(new_n822), .B1(new_n831), .B2(G29), .ZN(new_n832));
  OAI21_X1  g407(.A(new_n821), .B1(new_n832), .B2(new_n819), .ZN(new_n833));
  INV_X1    g408(.A(G2067), .ZN(new_n834));
  XNOR2_X1  g409(.A(new_n833), .B(new_n834), .ZN(new_n835));
  INV_X1    g410(.A(KEYINPUT23), .ZN(new_n836));
  AND3_X1   g411(.A1(new_n836), .A2(new_n744), .A3(G20), .ZN(new_n837));
  NAND2_X1  g412(.A1(G299), .A2(G16), .ZN(new_n838));
  AOI21_X1  g413(.A(new_n836), .B1(new_n744), .B2(G20), .ZN(new_n839));
  AOI21_X1  g414(.A(new_n837), .B1(new_n838), .B2(new_n839), .ZN(new_n840));
  XNOR2_X1  g415(.A(KEYINPUT105), .B(G1956), .ZN(new_n841));
  XNOR2_X1  g416(.A(new_n840), .B(new_n841), .ZN(new_n842));
  NAND3_X1  g417(.A1(new_n818), .A2(new_n835), .A3(new_n842), .ZN(new_n843));
  NOR2_X1   g418(.A1(new_n787), .A2(new_n843), .ZN(new_n844));
  MUX2_X1   g419(.A(G23), .B(G288), .S(G16), .Z(new_n845));
  XOR2_X1   g420(.A(KEYINPUT33), .B(G1976), .Z(new_n846));
  XNOR2_X1  g421(.A(new_n845), .B(new_n846), .ZN(new_n847));
  NAND2_X1  g422(.A1(new_n744), .A2(G6), .ZN(new_n848));
  INV_X1    g423(.A(G305), .ZN(new_n849));
  OAI21_X1  g424(.A(new_n848), .B1(new_n849), .B2(new_n744), .ZN(new_n850));
  XNOR2_X1  g425(.A(KEYINPUT32), .B(G1981), .ZN(new_n851));
  NOR2_X1   g426(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  NOR2_X1   g427(.A1(new_n847), .A2(new_n852), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n850), .A2(new_n851), .ZN(new_n854));
  AND2_X1   g429(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  INV_X1    g430(.A(KEYINPUT34), .ZN(new_n856));
  NAND2_X1  g431(.A1(new_n744), .A2(G22), .ZN(new_n857));
  OAI21_X1  g432(.A(new_n857), .B1(G166), .B2(new_n744), .ZN(new_n858));
  OR2_X1    g433(.A1(new_n858), .A2(G1971), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n858), .A2(G1971), .ZN(new_n860));
  NAND4_X1  g435(.A1(new_n855), .A2(new_n856), .A3(new_n859), .A4(new_n860), .ZN(new_n861));
  NAND4_X1  g436(.A1(new_n853), .A2(new_n859), .A3(new_n860), .A4(new_n854), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n862), .A2(KEYINPUT34), .ZN(new_n863));
  MUX2_X1   g438(.A(G24), .B(G290), .S(G16), .Z(new_n864));
  XOR2_X1   g439(.A(KEYINPUT99), .B(G1986), .Z(new_n865));
  XOR2_X1   g440(.A(new_n864), .B(new_n865), .Z(new_n866));
  NAND2_X1  g441(.A1(new_n768), .A2(G25), .ZN(new_n867));
  XOR2_X1   g442(.A(new_n867), .B(KEYINPUT97), .Z(new_n868));
  NAND2_X1  g443(.A1(new_n674), .A2(G119), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n669), .A2(G131), .ZN(new_n870));
  OR2_X1    g445(.A1(G95), .A2(G2105), .ZN(new_n871));
  OAI211_X1 g446(.A(new_n871), .B(G2104), .C1(G107), .C2(new_n475), .ZN(new_n872));
  NAND3_X1  g447(.A1(new_n869), .A2(new_n870), .A3(new_n872), .ZN(new_n873));
  INV_X1    g448(.A(new_n873), .ZN(new_n874));
  OAI21_X1  g449(.A(new_n868), .B1(new_n874), .B2(new_n768), .ZN(new_n875));
  XNOR2_X1  g450(.A(KEYINPUT35), .B(G1991), .ZN(new_n876));
  XNOR2_X1  g451(.A(new_n876), .B(KEYINPUT98), .ZN(new_n877));
  INV_X1    g452(.A(new_n877), .ZN(new_n878));
  AND2_X1   g453(.A1(new_n875), .A2(new_n878), .ZN(new_n879));
  NOR2_X1   g454(.A1(new_n875), .A2(new_n878), .ZN(new_n880));
  NOR3_X1   g455(.A1(new_n866), .A2(new_n879), .A3(new_n880), .ZN(new_n881));
  NAND3_X1  g456(.A1(new_n861), .A2(new_n863), .A3(new_n881), .ZN(new_n882));
  AND2_X1   g457(.A1(new_n882), .A2(KEYINPUT36), .ZN(new_n883));
  NOR2_X1   g458(.A1(new_n882), .A2(KEYINPUT36), .ZN(new_n884));
  OAI21_X1  g459(.A(new_n844), .B1(new_n883), .B2(new_n884), .ZN(new_n885));
  INV_X1    g460(.A(new_n885), .ZN(G311));
  INV_X1    g461(.A(KEYINPUT106), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n885), .A2(new_n887), .ZN(new_n888));
  OAI211_X1 g463(.A(new_n844), .B(KEYINPUT106), .C1(new_n883), .C2(new_n884), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n888), .A2(new_n889), .ZN(G150));
  NAND3_X1  g465(.A1(new_n521), .A2(G67), .A3(new_n524), .ZN(new_n891));
  NAND2_X1  g466(.A1(G80), .A2(G543), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n893), .A2(G651), .ZN(new_n894));
  NAND3_X1  g469(.A1(new_n564), .A2(G55), .A3(new_n565), .ZN(new_n895));
  NAND3_X1  g470(.A1(new_n528), .A2(G93), .A3(new_n543), .ZN(new_n896));
  NAND3_X1  g471(.A1(new_n894), .A2(new_n895), .A3(new_n896), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n897), .A2(G860), .ZN(new_n898));
  XNOR2_X1  g473(.A(new_n898), .B(KEYINPUT109), .ZN(new_n899));
  XNOR2_X1  g474(.A(new_n899), .B(KEYINPUT37), .ZN(new_n900));
  INV_X1    g475(.A(KEYINPUT107), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n897), .A2(new_n901), .ZN(new_n902));
  OR3_X1    g477(.A1(new_n582), .A2(new_n585), .A3(new_n587), .ZN(new_n903));
  NAND4_X1  g478(.A1(new_n894), .A2(KEYINPUT107), .A3(new_n895), .A4(new_n896), .ZN(new_n904));
  NAND3_X1  g479(.A1(new_n902), .A2(new_n903), .A3(new_n904), .ZN(new_n905));
  INV_X1    g480(.A(new_n897), .ZN(new_n906));
  NAND3_X1  g481(.A1(new_n906), .A2(KEYINPUT107), .A3(new_n588), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n905), .A2(new_n907), .ZN(new_n908));
  XNOR2_X1  g483(.A(new_n908), .B(KEYINPUT38), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n661), .A2(G559), .ZN(new_n910));
  XNOR2_X1  g485(.A(new_n909), .B(new_n910), .ZN(new_n911));
  INV_X1    g486(.A(new_n911), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n912), .A2(KEYINPUT39), .ZN(new_n913));
  XOR2_X1   g488(.A(new_n913), .B(KEYINPUT108), .Z(new_n914));
  INV_X1    g489(.A(G860), .ZN(new_n915));
  OAI21_X1  g490(.A(new_n915), .B1(new_n912), .B2(KEYINPUT39), .ZN(new_n916));
  OAI21_X1  g491(.A(new_n900), .B1(new_n914), .B2(new_n916), .ZN(G145));
  XOR2_X1   g492(.A(new_n502), .B(new_n675), .Z(new_n918));
  NAND2_X1  g493(.A1(new_n674), .A2(G130), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n669), .A2(G142), .ZN(new_n920));
  OR2_X1    g495(.A1(G106), .A2(G2105), .ZN(new_n921));
  OAI211_X1 g496(.A(new_n921), .B(G2104), .C1(G118), .C2(new_n475), .ZN(new_n922));
  NAND3_X1  g497(.A1(new_n919), .A2(new_n920), .A3(new_n922), .ZN(new_n923));
  INV_X1    g498(.A(new_n680), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  NAND4_X1  g500(.A1(new_n919), .A2(new_n920), .A3(new_n680), .A4(new_n922), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n927), .A2(new_n873), .ZN(new_n928));
  NAND3_X1  g503(.A1(new_n925), .A2(new_n874), .A3(new_n926), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n930), .A2(KEYINPUT110), .ZN(new_n931));
  INV_X1    g506(.A(KEYINPUT110), .ZN(new_n932));
  NAND3_X1  g507(.A1(new_n928), .A2(new_n932), .A3(new_n929), .ZN(new_n933));
  INV_X1    g508(.A(new_n796), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n831), .A2(new_n934), .ZN(new_n935));
  XNOR2_X1  g510(.A(new_n777), .B(G164), .ZN(new_n936));
  NAND3_X1  g511(.A1(new_n829), .A2(new_n830), .A3(new_n796), .ZN(new_n937));
  NAND3_X1  g512(.A1(new_n935), .A2(new_n936), .A3(new_n937), .ZN(new_n938));
  INV_X1    g513(.A(new_n938), .ZN(new_n939));
  AOI21_X1  g514(.A(new_n936), .B1(new_n935), .B2(new_n937), .ZN(new_n940));
  OAI211_X1 g515(.A(new_n931), .B(new_n933), .C1(new_n939), .C2(new_n940), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n935), .A2(new_n937), .ZN(new_n942));
  OAI221_X1 g517(.A(new_n511), .B1(new_n472), .B2(new_n513), .C1(new_n505), .C2(KEYINPUT4), .ZN(new_n943));
  XNOR2_X1  g518(.A(new_n777), .B(new_n943), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n942), .A2(new_n944), .ZN(new_n945));
  NAND4_X1  g520(.A1(new_n945), .A2(KEYINPUT110), .A3(new_n938), .A4(new_n930), .ZN(new_n946));
  AND3_X1   g521(.A1(new_n941), .A2(new_n491), .A3(new_n946), .ZN(new_n947));
  AOI21_X1  g522(.A(new_n491), .B1(new_n941), .B2(new_n946), .ZN(new_n948));
  OAI21_X1  g523(.A(new_n918), .B1(new_n947), .B2(new_n948), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n941), .A2(new_n946), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n950), .A2(G160), .ZN(new_n951));
  INV_X1    g526(.A(new_n918), .ZN(new_n952));
  NAND3_X1  g527(.A1(new_n941), .A2(new_n491), .A3(new_n946), .ZN(new_n953));
  NAND3_X1  g528(.A1(new_n951), .A2(new_n952), .A3(new_n953), .ZN(new_n954));
  INV_X1    g529(.A(G37), .ZN(new_n955));
  NAND3_X1  g530(.A1(new_n949), .A2(new_n954), .A3(new_n955), .ZN(new_n956));
  XNOR2_X1  g531(.A(new_n956), .B(KEYINPUT40), .ZN(G395));
  XOR2_X1   g532(.A(new_n908), .B(new_n664), .Z(new_n958));
  NAND2_X1  g533(.A1(G299), .A2(new_n661), .ZN(new_n959));
  NAND3_X1  g534(.A1(new_n601), .A2(new_n609), .A3(new_n653), .ZN(new_n960));
  NAND2_X1  g535(.A1(new_n959), .A2(new_n960), .ZN(new_n961));
  INV_X1    g536(.A(new_n961), .ZN(new_n962));
  NOR2_X1   g537(.A1(new_n958), .A2(new_n962), .ZN(new_n963));
  INV_X1    g538(.A(KEYINPUT41), .ZN(new_n964));
  INV_X1    g539(.A(new_n960), .ZN(new_n965));
  AOI21_X1  g540(.A(new_n653), .B1(new_n601), .B2(new_n609), .ZN(new_n966));
  OAI21_X1  g541(.A(new_n964), .B1(new_n965), .B2(new_n966), .ZN(new_n967));
  NAND3_X1  g542(.A1(new_n959), .A2(KEYINPUT41), .A3(new_n960), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n967), .A2(new_n968), .ZN(new_n969));
  AOI21_X1  g544(.A(new_n963), .B1(new_n958), .B2(new_n969), .ZN(new_n970));
  XOR2_X1   g545(.A(KEYINPUT111), .B(KEYINPUT42), .Z(new_n971));
  INV_X1    g546(.A(new_n971), .ZN(new_n972));
  OR2_X1    g547(.A1(new_n970), .A2(new_n972), .ZN(new_n973));
  NAND2_X1  g548(.A1(G290), .A2(G288), .ZN(new_n974));
  INV_X1    g549(.A(new_n974), .ZN(new_n975));
  NOR2_X1   g550(.A1(G290), .A2(G288), .ZN(new_n976));
  OAI211_X1 g551(.A(new_n621), .B(new_n532), .C1(new_n975), .C2(new_n976), .ZN(new_n977));
  OR2_X1    g552(.A1(G290), .A2(G288), .ZN(new_n978));
  OAI211_X1 g553(.A(new_n978), .B(new_n974), .C1(new_n533), .C2(new_n545), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n977), .A2(new_n979), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n980), .A2(G305), .ZN(new_n981));
  NAND3_X1  g556(.A1(new_n977), .A2(new_n979), .A3(new_n849), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n981), .A2(new_n982), .ZN(new_n983));
  NAND2_X1  g558(.A1(new_n970), .A2(new_n972), .ZN(new_n984));
  AND3_X1   g559(.A1(new_n973), .A2(new_n983), .A3(new_n984), .ZN(new_n985));
  AOI21_X1  g560(.A(new_n983), .B1(new_n973), .B2(new_n984), .ZN(new_n986));
  OAI21_X1  g561(.A(G868), .B1(new_n985), .B2(new_n986), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n897), .A2(new_n654), .ZN(new_n988));
  NAND2_X1  g563(.A1(new_n987), .A2(new_n988), .ZN(G295));
  NAND2_X1  g564(.A1(new_n987), .A2(new_n988), .ZN(G331));
  INV_X1    g565(.A(KEYINPUT113), .ZN(new_n991));
  NAND2_X1  g566(.A1(G168), .A2(G301), .ZN(new_n992));
  NAND2_X1  g567(.A1(G171), .A2(G286), .ZN(new_n993));
  NAND3_X1  g568(.A1(new_n908), .A2(new_n992), .A3(new_n993), .ZN(new_n994));
  NOR2_X1   g569(.A1(G171), .A2(G286), .ZN(new_n995));
  NOR2_X1   g570(.A1(G168), .A2(G301), .ZN(new_n996));
  OAI211_X1 g571(.A(new_n907), .B(new_n905), .C1(new_n995), .C2(new_n996), .ZN(new_n997));
  AOI22_X1  g572(.A1(new_n994), .A2(new_n997), .B1(new_n967), .B2(new_n968), .ZN(new_n998));
  INV_X1    g573(.A(KEYINPUT112), .ZN(new_n999));
  NAND3_X1  g574(.A1(new_n997), .A2(new_n994), .A3(new_n999), .ZN(new_n1000));
  NAND4_X1  g575(.A1(new_n908), .A2(KEYINPUT112), .A3(new_n992), .A4(new_n993), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n1000), .A2(new_n1001), .ZN(new_n1002));
  AOI21_X1  g577(.A(new_n998), .B1(new_n1002), .B2(new_n961), .ZN(new_n1003));
  INV_X1    g578(.A(new_n983), .ZN(new_n1004));
  AOI21_X1  g579(.A(new_n991), .B1(new_n1003), .B2(new_n1004), .ZN(new_n1005));
  AOI21_X1  g580(.A(new_n962), .B1(new_n1000), .B2(new_n1001), .ZN(new_n1006));
  NOR4_X1   g581(.A1(new_n1006), .A2(new_n983), .A3(new_n998), .A4(KEYINPUT113), .ZN(new_n1007));
  NOR3_X1   g582(.A1(new_n1005), .A2(new_n1007), .A3(G37), .ZN(new_n1008));
  OAI21_X1  g583(.A(new_n983), .B1(new_n1006), .B2(new_n998), .ZN(new_n1009));
  AOI21_X1  g584(.A(KEYINPUT43), .B1(new_n1008), .B2(new_n1009), .ZN(new_n1010));
  NOR3_X1   g585(.A1(new_n1006), .A2(new_n983), .A3(new_n998), .ZN(new_n1011));
  OAI21_X1  g586(.A(new_n955), .B1(new_n1011), .B2(new_n991), .ZN(new_n1012));
  NAND3_X1  g587(.A1(new_n997), .A2(new_n994), .A3(new_n961), .ZN(new_n1013));
  INV_X1    g588(.A(KEYINPUT114), .ZN(new_n1014));
  XNOR2_X1  g589(.A(new_n1013), .B(new_n1014), .ZN(new_n1015));
  NAND3_X1  g590(.A1(new_n1000), .A2(new_n969), .A3(new_n1001), .ZN(new_n1016));
  AOI21_X1  g591(.A(new_n1004), .B1(new_n1015), .B2(new_n1016), .ZN(new_n1017));
  INV_X1    g592(.A(KEYINPUT43), .ZN(new_n1018));
  NOR4_X1   g593(.A1(new_n1012), .A2(new_n1017), .A3(new_n1018), .A4(new_n1007), .ZN(new_n1019));
  OAI21_X1  g594(.A(KEYINPUT44), .B1(new_n1010), .B2(new_n1019), .ZN(new_n1020));
  INV_X1    g595(.A(KEYINPUT44), .ZN(new_n1021));
  AOI21_X1  g596(.A(new_n1018), .B1(new_n1008), .B2(new_n1009), .ZN(new_n1022));
  NOR4_X1   g597(.A1(new_n1012), .A2(new_n1017), .A3(KEYINPUT43), .A4(new_n1007), .ZN(new_n1023));
  OAI21_X1  g598(.A(new_n1021), .B1(new_n1022), .B2(new_n1023), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n1020), .A2(new_n1024), .ZN(G397));
  INV_X1    g600(.A(G1384), .ZN(new_n1026));
  AOI21_X1  g601(.A(KEYINPUT45), .B1(new_n943), .B2(new_n1026), .ZN(new_n1027));
  INV_X1    g602(.A(new_n1027), .ZN(new_n1028));
  NAND4_X1  g603(.A1(new_n477), .A2(G40), .A3(new_n479), .A4(new_n490), .ZN(new_n1029));
  NOR2_X1   g604(.A1(new_n1028), .A2(new_n1029), .ZN(new_n1030));
  INV_X1    g605(.A(G1996), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n1030), .A2(new_n1031), .ZN(new_n1032));
  XOR2_X1   g607(.A(new_n1032), .B(KEYINPUT46), .Z(new_n1033));
  XNOR2_X1  g608(.A(new_n831), .B(new_n834), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n1034), .A2(new_n778), .ZN(new_n1035));
  AOI21_X1  g610(.A(new_n1033), .B1(new_n1035), .B2(new_n1030), .ZN(new_n1036));
  XNOR2_X1  g611(.A(KEYINPUT127), .B(KEYINPUT47), .ZN(new_n1037));
  XNOR2_X1  g612(.A(new_n1036), .B(new_n1037), .ZN(new_n1038));
  XNOR2_X1  g613(.A(new_n777), .B(new_n1031), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n1034), .A2(new_n1039), .ZN(new_n1040));
  OR2_X1    g615(.A1(new_n873), .A2(new_n876), .ZN(new_n1041));
  OAI22_X1  g616(.A1(new_n1040), .A2(new_n1041), .B1(G2067), .B2(new_n831), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n1042), .A2(new_n1030), .ZN(new_n1043));
  INV_X1    g618(.A(new_n1030), .ZN(new_n1044));
  NOR3_X1   g619(.A1(new_n1044), .A2(G1986), .A3(G290), .ZN(new_n1045));
  XOR2_X1   g620(.A(new_n1045), .B(KEYINPUT48), .Z(new_n1046));
  NAND2_X1  g621(.A1(new_n873), .A2(new_n876), .ZN(new_n1047));
  AND4_X1   g622(.A1(new_n1034), .A2(new_n1039), .A3(new_n1047), .A4(new_n1041), .ZN(new_n1048));
  OAI21_X1  g623(.A(new_n1046), .B1(new_n1048), .B2(new_n1044), .ZN(new_n1049));
  AND3_X1   g624(.A1(new_n1038), .A2(new_n1043), .A3(new_n1049), .ZN(new_n1050));
  INV_X1    g625(.A(KEYINPUT63), .ZN(new_n1051));
  INV_X1    g626(.A(KEYINPUT55), .ZN(new_n1052));
  INV_X1    g627(.A(G8), .ZN(new_n1053));
  OAI21_X1  g628(.A(new_n1052), .B1(G166), .B2(new_n1053), .ZN(new_n1054));
  NAND3_X1  g629(.A1(G303), .A2(KEYINPUT55), .A3(G8), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n1054), .A2(new_n1055), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n1056), .A2(KEYINPUT116), .ZN(new_n1057));
  INV_X1    g632(.A(KEYINPUT116), .ZN(new_n1058));
  NAND3_X1  g633(.A1(new_n1054), .A2(new_n1055), .A3(new_n1058), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n1057), .A2(new_n1059), .ZN(new_n1060));
  INV_X1    g635(.A(new_n1029), .ZN(new_n1061));
  INV_X1    g636(.A(G2090), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n943), .A2(new_n1026), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n1063), .A2(KEYINPUT50), .ZN(new_n1064));
  INV_X1    g639(.A(KEYINPUT50), .ZN(new_n1065));
  NAND3_X1  g640(.A1(new_n943), .A2(new_n1065), .A3(new_n1026), .ZN(new_n1066));
  NAND4_X1  g641(.A1(new_n1061), .A2(new_n1062), .A3(new_n1064), .A4(new_n1066), .ZN(new_n1067));
  INV_X1    g642(.A(KEYINPUT115), .ZN(new_n1068));
  NAND3_X1  g643(.A1(new_n943), .A2(KEYINPUT45), .A3(new_n1026), .ZN(new_n1069));
  NAND3_X1  g644(.A1(new_n1061), .A2(new_n1028), .A3(new_n1069), .ZN(new_n1070));
  INV_X1    g645(.A(G1971), .ZN(new_n1071));
  AOI22_X1  g646(.A1(new_n1067), .A2(new_n1068), .B1(new_n1070), .B2(new_n1071), .ZN(new_n1072));
  INV_X1    g647(.A(new_n1067), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n1073), .A2(KEYINPUT115), .ZN(new_n1074));
  AOI21_X1  g649(.A(new_n1053), .B1(new_n1072), .B2(new_n1074), .ZN(new_n1075));
  AOI21_X1  g650(.A(new_n1051), .B1(new_n1060), .B2(new_n1075), .ZN(new_n1076));
  NOR2_X1   g651(.A1(new_n1029), .A2(new_n1063), .ZN(new_n1077));
  NOR2_X1   g652(.A1(new_n1077), .A2(new_n1053), .ZN(new_n1078));
  XOR2_X1   g653(.A(KEYINPUT118), .B(G1981), .Z(new_n1079));
  OAI211_X1 g654(.A(new_n630), .B(new_n1079), .C1(new_n634), .C2(new_n635), .ZN(new_n1080));
  INV_X1    g655(.A(new_n630), .ZN(new_n1081));
  AND2_X1   g656(.A1(new_n633), .A2(G651), .ZN(new_n1082));
  OAI21_X1  g657(.A(G1981), .B1(new_n1081), .B2(new_n1082), .ZN(new_n1083));
  NAND3_X1  g658(.A1(new_n1080), .A2(KEYINPUT49), .A3(new_n1083), .ZN(new_n1084));
  AND2_X1   g659(.A1(new_n1078), .A2(new_n1084), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n1080), .A2(new_n1083), .ZN(new_n1086));
  INV_X1    g661(.A(KEYINPUT49), .ZN(new_n1087));
  NAND2_X1  g662(.A1(new_n1086), .A2(new_n1087), .ZN(new_n1088));
  NAND4_X1  g663(.A1(new_n623), .A2(new_n624), .A3(new_n625), .A4(G1976), .ZN(new_n1089));
  OAI211_X1 g664(.A(G8), .B(new_n1089), .C1(new_n1029), .C2(new_n1063), .ZN(new_n1090));
  NAND2_X1  g665(.A1(KEYINPUT117), .A2(KEYINPUT52), .ZN(new_n1091));
  OR2_X1    g666(.A1(new_n1090), .A2(new_n1091), .ZN(new_n1092));
  NOR2_X1   g667(.A1(KEYINPUT52), .A2(G1976), .ZN(new_n1093));
  AOI22_X1  g668(.A1(new_n1090), .A2(new_n1091), .B1(G288), .B2(new_n1093), .ZN(new_n1094));
  AOI22_X1  g669(.A1(new_n1085), .A2(new_n1088), .B1(new_n1092), .B2(new_n1094), .ZN(new_n1095));
  OAI21_X1  g670(.A(new_n1095), .B1(new_n1075), .B2(new_n1056), .ZN(new_n1096));
  INV_X1    g671(.A(KEYINPUT122), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n1096), .A2(new_n1097), .ZN(new_n1098));
  INV_X1    g673(.A(new_n1069), .ZN(new_n1099));
  NOR3_X1   g674(.A1(new_n1099), .A2(new_n1029), .A3(new_n1027), .ZN(new_n1100));
  NAND3_X1  g675(.A1(new_n1061), .A2(new_n1064), .A3(new_n1066), .ZN(new_n1101));
  OAI22_X1  g676(.A1(G1966), .A2(new_n1100), .B1(new_n1101), .B2(G2084), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n1102), .A2(G8), .ZN(new_n1103));
  NOR2_X1   g678(.A1(new_n1103), .A2(G286), .ZN(new_n1104));
  OAI211_X1 g679(.A(new_n1095), .B(KEYINPUT122), .C1(new_n1075), .C2(new_n1056), .ZN(new_n1105));
  NAND4_X1  g680(.A1(new_n1076), .A2(new_n1098), .A3(new_n1104), .A4(new_n1105), .ZN(new_n1106));
  XOR2_X1   g681(.A(KEYINPUT121), .B(KEYINPUT63), .Z(new_n1107));
  NAND2_X1  g682(.A1(new_n1106), .A2(new_n1107), .ZN(new_n1108));
  AND2_X1   g683(.A1(new_n1060), .A2(new_n1075), .ZN(new_n1109));
  XNOR2_X1  g684(.A(new_n1080), .B(KEYINPUT119), .ZN(new_n1110));
  AND2_X1   g685(.A1(new_n1085), .A2(new_n1088), .ZN(new_n1111));
  OR2_X1    g686(.A1(G288), .A2(G1976), .ZN(new_n1112));
  OAI21_X1  g687(.A(new_n1110), .B1(new_n1111), .B2(new_n1112), .ZN(new_n1113));
  AOI22_X1  g688(.A1(new_n1109), .A2(new_n1095), .B1(new_n1078), .B2(new_n1113), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n1108), .A2(new_n1114), .ZN(new_n1115));
  INV_X1    g690(.A(G1956), .ZN(new_n1116));
  NAND2_X1  g691(.A1(new_n1101), .A2(new_n1116), .ZN(new_n1117));
  NAND2_X1  g692(.A1(KEYINPUT123), .A2(KEYINPUT57), .ZN(new_n1118));
  INV_X1    g693(.A(KEYINPUT123), .ZN(new_n1119));
  INV_X1    g694(.A(KEYINPUT57), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n1119), .A2(new_n1120), .ZN(new_n1121));
  NAND3_X1  g696(.A1(G299), .A2(new_n1118), .A3(new_n1121), .ZN(new_n1122));
  NAND4_X1  g697(.A1(new_n601), .A2(new_n609), .A3(new_n1119), .A4(new_n1120), .ZN(new_n1123));
  XNOR2_X1  g698(.A(KEYINPUT56), .B(G2072), .ZN(new_n1124));
  NAND4_X1  g699(.A1(new_n1061), .A2(new_n1028), .A3(new_n1069), .A4(new_n1124), .ZN(new_n1125));
  NAND4_X1  g700(.A1(new_n1117), .A2(new_n1122), .A3(new_n1123), .A4(new_n1125), .ZN(new_n1126));
  NAND2_X1  g701(.A1(new_n1122), .A2(new_n1123), .ZN(new_n1127));
  NAND2_X1  g702(.A1(new_n1127), .A2(KEYINPUT124), .ZN(new_n1128));
  INV_X1    g703(.A(KEYINPUT124), .ZN(new_n1129));
  NAND3_X1  g704(.A1(new_n1122), .A2(new_n1129), .A3(new_n1123), .ZN(new_n1130));
  NAND2_X1  g705(.A1(new_n1117), .A2(new_n1125), .ZN(new_n1131));
  AND3_X1   g706(.A1(new_n1128), .A2(new_n1130), .A3(new_n1131), .ZN(new_n1132));
  AOI22_X1  g707(.A1(new_n1101), .A2(new_n747), .B1(new_n834), .B2(new_n1077), .ZN(new_n1133));
  NOR2_X1   g708(.A1(new_n1133), .A2(new_n653), .ZN(new_n1134));
  OAI21_X1  g709(.A(new_n1126), .B1(new_n1132), .B2(new_n1134), .ZN(new_n1135));
  AOI21_X1  g710(.A(new_n653), .B1(new_n1133), .B2(KEYINPUT60), .ZN(new_n1136));
  NAND2_X1  g711(.A1(new_n1064), .A2(new_n1066), .ZN(new_n1137));
  OAI21_X1  g712(.A(new_n747), .B1(new_n1137), .B2(new_n1029), .ZN(new_n1138));
  NAND2_X1  g713(.A1(new_n1077), .A2(new_n834), .ZN(new_n1139));
  AND4_X1   g714(.A1(KEYINPUT60), .A2(new_n1138), .A3(new_n653), .A4(new_n1139), .ZN(new_n1140));
  OAI22_X1  g715(.A1(new_n1136), .A2(new_n1140), .B1(KEYINPUT60), .B2(new_n1133), .ZN(new_n1141));
  INV_X1    g716(.A(KEYINPUT61), .ZN(new_n1142));
  INV_X1    g717(.A(new_n1126), .ZN(new_n1143));
  AOI22_X1  g718(.A1(new_n1117), .A2(new_n1125), .B1(new_n1122), .B2(new_n1123), .ZN(new_n1144));
  OAI21_X1  g719(.A(new_n1142), .B1(new_n1143), .B2(new_n1144), .ZN(new_n1145));
  XNOR2_X1  g720(.A(KEYINPUT125), .B(KEYINPUT59), .ZN(new_n1146));
  NAND4_X1  g721(.A1(new_n1061), .A2(new_n1028), .A3(new_n1031), .A4(new_n1069), .ZN(new_n1147));
  XOR2_X1   g722(.A(KEYINPUT58), .B(G1341), .Z(new_n1148));
  OAI21_X1  g723(.A(new_n1148), .B1(new_n1029), .B2(new_n1063), .ZN(new_n1149));
  AOI211_X1 g724(.A(new_n903), .B(new_n1146), .C1(new_n1147), .C2(new_n1149), .ZN(new_n1150));
  NOR2_X1   g725(.A1(KEYINPUT125), .A2(KEYINPUT59), .ZN(new_n1151));
  NAND2_X1  g726(.A1(new_n1147), .A2(new_n1149), .ZN(new_n1152));
  NAND2_X1  g727(.A1(new_n1152), .A2(new_n588), .ZN(new_n1153));
  AOI21_X1  g728(.A(new_n1150), .B1(new_n1151), .B2(new_n1153), .ZN(new_n1154));
  NAND3_X1  g729(.A1(new_n1141), .A2(new_n1145), .A3(new_n1154), .ZN(new_n1155));
  NAND2_X1  g730(.A1(new_n1126), .A2(KEYINPUT61), .ZN(new_n1156));
  NOR2_X1   g731(.A1(new_n1132), .A2(new_n1156), .ZN(new_n1157));
  OAI21_X1  g732(.A(new_n1135), .B1(new_n1155), .B2(new_n1157), .ZN(new_n1158));
  INV_X1    g733(.A(KEYINPUT54), .ZN(new_n1159));
  NAND3_X1  g734(.A1(new_n1100), .A2(KEYINPUT53), .A3(new_n443), .ZN(new_n1160));
  NAND2_X1  g735(.A1(new_n1101), .A2(new_n752), .ZN(new_n1161));
  NAND2_X1  g736(.A1(new_n1160), .A2(new_n1161), .ZN(new_n1162));
  AOI21_X1  g737(.A(KEYINPUT53), .B1(new_n1100), .B2(new_n443), .ZN(new_n1163));
  OAI21_X1  g738(.A(G171), .B1(new_n1162), .B2(new_n1163), .ZN(new_n1164));
  INV_X1    g739(.A(KEYINPUT126), .ZN(new_n1165));
  OAI21_X1  g740(.A(new_n1160), .B1(new_n1163), .B2(new_n1165), .ZN(new_n1166));
  NAND4_X1  g741(.A1(new_n1100), .A2(KEYINPUT126), .A3(KEYINPUT53), .A4(new_n443), .ZN(new_n1167));
  NAND3_X1  g742(.A1(new_n1166), .A2(new_n1167), .A3(new_n1161), .ZN(new_n1168));
  NOR2_X1   g743(.A1(new_n1163), .A2(G171), .ZN(new_n1169));
  INV_X1    g744(.A(new_n1169), .ZN(new_n1170));
  OAI211_X1 g745(.A(new_n1159), .B(new_n1164), .C1(new_n1168), .C2(new_n1170), .ZN(new_n1171));
  INV_X1    g746(.A(new_n1162), .ZN(new_n1172));
  AOI22_X1  g747(.A1(new_n1168), .A2(G171), .B1(new_n1172), .B2(new_n1169), .ZN(new_n1173));
  OAI21_X1  g748(.A(new_n1171), .B1(new_n1173), .B2(new_n1159), .ZN(new_n1174));
  OAI211_X1 g749(.A(new_n1103), .B(KEYINPUT51), .C1(new_n1053), .C2(G168), .ZN(new_n1175));
  NAND3_X1  g750(.A1(new_n1102), .A2(G8), .A3(G286), .ZN(new_n1176));
  INV_X1    g751(.A(KEYINPUT51), .ZN(new_n1177));
  OAI211_X1 g752(.A(new_n1177), .B(G8), .C1(new_n1102), .C2(G286), .ZN(new_n1178));
  NAND3_X1  g753(.A1(new_n1175), .A2(new_n1176), .A3(new_n1178), .ZN(new_n1179));
  NAND3_X1  g754(.A1(new_n1158), .A2(new_n1174), .A3(new_n1179), .ZN(new_n1180));
  NAND3_X1  g755(.A1(new_n1076), .A2(new_n1105), .A3(new_n1098), .ZN(new_n1181));
  NAND2_X1  g756(.A1(new_n1181), .A2(new_n1104), .ZN(new_n1182));
  AOI21_X1  g757(.A(new_n1164), .B1(new_n1179), .B2(KEYINPUT62), .ZN(new_n1183));
  OAI21_X1  g758(.A(new_n1183), .B1(KEYINPUT62), .B2(new_n1179), .ZN(new_n1184));
  NAND3_X1  g759(.A1(new_n1180), .A2(new_n1182), .A3(new_n1184), .ZN(new_n1185));
  XOR2_X1   g760(.A(new_n1095), .B(KEYINPUT120), .Z(new_n1186));
  OAI21_X1  g761(.A(new_n1067), .B1(new_n1100), .B2(G1971), .ZN(new_n1187));
  AOI21_X1  g762(.A(new_n1056), .B1(new_n1187), .B2(G8), .ZN(new_n1188));
  NOR3_X1   g763(.A1(new_n1186), .A2(new_n1109), .A3(new_n1188), .ZN(new_n1189));
  AOI21_X1  g764(.A(new_n1115), .B1(new_n1185), .B2(new_n1189), .ZN(new_n1190));
  XOR2_X1   g765(.A(G290), .B(G1986), .Z(new_n1191));
  AOI21_X1  g766(.A(new_n1044), .B1(new_n1048), .B2(new_n1191), .ZN(new_n1192));
  OAI21_X1  g767(.A(new_n1050), .B1(new_n1190), .B2(new_n1192), .ZN(G329));
  assign    G231 = 1'b0;
  NOR4_X1   g768(.A1(G401), .A2(new_n464), .A3(G227), .A4(G229), .ZN(new_n1195));
  OAI211_X1 g769(.A(new_n956), .B(new_n1195), .C1(new_n1022), .C2(new_n1023), .ZN(G225));
  INV_X1    g770(.A(G225), .ZN(G308));
endmodule


