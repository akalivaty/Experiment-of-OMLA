//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 1 0 0 0 0 1 1 1 1 0 0 0 0 0 0 1 0 1 1 0 0 0 1 0 1 1 0 0 0 0 0 1 0 1 0 1 1 0 1 1 0 1 0 0 1 1 0 0 0 1 1 0 0 1 0 1 0 0 0 0 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:24:09 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n699, new_n700, new_n701, new_n702, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n714, new_n715, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n730, new_n731, new_n732, new_n733, new_n734, new_n735,
    new_n736, new_n737, new_n738, new_n739, new_n740, new_n741, new_n743,
    new_n744, new_n745, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n772, new_n773,
    new_n774, new_n775, new_n776, new_n777, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n805, new_n806, new_n807, new_n808, new_n809, new_n810,
    new_n811, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n942, new_n943, new_n944, new_n945,
    new_n946, new_n947, new_n948, new_n949, new_n950, new_n951, new_n952,
    new_n953, new_n954, new_n955, new_n956, new_n957, new_n958, new_n959,
    new_n960, new_n961, new_n962, new_n963, new_n964, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n983,
    new_n984, new_n985, new_n986, new_n987, new_n988, new_n989, new_n991,
    new_n992, new_n993, new_n994, new_n995, new_n996, new_n997, new_n998,
    new_n999, new_n1000, new_n1001, new_n1002, new_n1003, new_n1005,
    new_n1006, new_n1007, new_n1008, new_n1009, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1022, new_n1023, new_n1024,
    new_n1025, new_n1026, new_n1027, new_n1028, new_n1029, new_n1030,
    new_n1031, new_n1032, new_n1033, new_n1034, new_n1035, new_n1036,
    new_n1037, new_n1038, new_n1039, new_n1040, new_n1041, new_n1042,
    new_n1043, new_n1044, new_n1045, new_n1046, new_n1047, new_n1048,
    new_n1050, new_n1051, new_n1052, new_n1053, new_n1054, new_n1055,
    new_n1056, new_n1057, new_n1058, new_n1059, new_n1060, new_n1061,
    new_n1062, new_n1063, new_n1064;
  INV_X1    g000(.A(KEYINPUT86), .ZN(new_n187));
  NOR3_X1   g001(.A1(KEYINPUT20), .A2(G475), .A3(G902), .ZN(new_n188));
  XNOR2_X1  g002(.A(G113), .B(G122), .ZN(new_n189));
  INV_X1    g003(.A(G104), .ZN(new_n190));
  XNOR2_X1  g004(.A(new_n189), .B(new_n190), .ZN(new_n191));
  INV_X1    g005(.A(KEYINPUT82), .ZN(new_n192));
  INV_X1    g006(.A(KEYINPUT19), .ZN(new_n193));
  INV_X1    g007(.A(G125), .ZN(new_n194));
  NOR2_X1   g008(.A1(new_n194), .A2(G140), .ZN(new_n195));
  INV_X1    g009(.A(G140), .ZN(new_n196));
  NOR2_X1   g010(.A1(new_n196), .A2(G125), .ZN(new_n197));
  OAI21_X1  g011(.A(new_n193), .B1(new_n195), .B2(new_n197), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n196), .A2(G125), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n194), .A2(G140), .ZN(new_n200));
  NAND3_X1  g014(.A1(new_n199), .A2(new_n200), .A3(KEYINPUT19), .ZN(new_n201));
  AOI21_X1  g015(.A(G146), .B1(new_n198), .B2(new_n201), .ZN(new_n202));
  NAND3_X1  g016(.A1(new_n199), .A2(new_n200), .A3(KEYINPUT16), .ZN(new_n203));
  INV_X1    g017(.A(KEYINPUT16), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n195), .A2(new_n204), .ZN(new_n205));
  AND3_X1   g019(.A1(new_n203), .A2(G146), .A3(new_n205), .ZN(new_n206));
  OAI21_X1  g020(.A(new_n192), .B1(new_n202), .B2(new_n206), .ZN(new_n207));
  INV_X1    g021(.A(G131), .ZN(new_n208));
  INV_X1    g022(.A(G237), .ZN(new_n209));
  INV_X1    g023(.A(G953), .ZN(new_n210));
  NAND3_X1  g024(.A1(new_n209), .A2(new_n210), .A3(G214), .ZN(new_n211));
  INV_X1    g025(.A(G143), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  NOR2_X1   g027(.A1(G237), .A2(G953), .ZN(new_n214));
  NAND3_X1  g028(.A1(new_n214), .A2(G143), .A3(G214), .ZN(new_n215));
  AOI21_X1  g029(.A(new_n208), .B1(new_n213), .B2(new_n215), .ZN(new_n216));
  INV_X1    g030(.A(new_n216), .ZN(new_n217));
  NAND3_X1  g031(.A1(new_n213), .A2(new_n208), .A3(new_n215), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  INV_X1    g033(.A(G146), .ZN(new_n220));
  AND3_X1   g034(.A1(new_n199), .A2(new_n200), .A3(KEYINPUT19), .ZN(new_n221));
  AOI21_X1  g035(.A(KEYINPUT19), .B1(new_n199), .B2(new_n200), .ZN(new_n222));
  OAI21_X1  g036(.A(new_n220), .B1(new_n221), .B2(new_n222), .ZN(new_n223));
  NAND3_X1  g037(.A1(new_n203), .A2(new_n205), .A3(G146), .ZN(new_n224));
  NAND3_X1  g038(.A1(new_n223), .A2(KEYINPUT82), .A3(new_n224), .ZN(new_n225));
  NAND3_X1  g039(.A1(new_n207), .A2(new_n219), .A3(new_n225), .ZN(new_n226));
  XNOR2_X1  g040(.A(G125), .B(G140), .ZN(new_n227));
  XNOR2_X1  g041(.A(new_n227), .B(new_n220), .ZN(new_n228));
  AND3_X1   g042(.A1(new_n214), .A2(G143), .A3(G214), .ZN(new_n229));
  AOI21_X1  g043(.A(G143), .B1(new_n214), .B2(G214), .ZN(new_n230));
  OAI211_X1 g044(.A(KEYINPUT18), .B(G131), .C1(new_n229), .C2(new_n230), .ZN(new_n231));
  NAND2_X1  g045(.A1(KEYINPUT18), .A2(G131), .ZN(new_n232));
  NAND3_X1  g046(.A1(new_n213), .A2(new_n215), .A3(new_n232), .ZN(new_n233));
  NAND3_X1  g047(.A1(new_n228), .A2(new_n231), .A3(new_n233), .ZN(new_n234));
  AOI21_X1  g048(.A(new_n191), .B1(new_n226), .B2(new_n234), .ZN(new_n235));
  NOR3_X1   g049(.A1(new_n229), .A2(new_n230), .A3(G131), .ZN(new_n236));
  NOR3_X1   g050(.A1(new_n236), .A2(new_n216), .A3(KEYINPUT17), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n203), .A2(new_n205), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n238), .A2(new_n220), .ZN(new_n239));
  OAI211_X1 g053(.A(KEYINPUT17), .B(G131), .C1(new_n229), .C2(new_n230), .ZN(new_n240));
  NAND3_X1  g054(.A1(new_n239), .A2(new_n240), .A3(new_n224), .ZN(new_n241));
  OAI211_X1 g055(.A(new_n191), .B(new_n234), .C1(new_n237), .C2(new_n241), .ZN(new_n242));
  INV_X1    g056(.A(new_n242), .ZN(new_n243));
  OAI21_X1  g057(.A(new_n188), .B1(new_n235), .B2(new_n243), .ZN(new_n244));
  INV_X1    g058(.A(KEYINPUT84), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n244), .A2(new_n245), .ZN(new_n246));
  OAI211_X1 g060(.A(KEYINPUT84), .B(new_n188), .C1(new_n235), .C2(new_n243), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n246), .A2(new_n247), .ZN(new_n248));
  INV_X1    g062(.A(new_n234), .ZN(new_n249));
  NOR2_X1   g063(.A1(new_n236), .A2(new_n216), .ZN(new_n250));
  NOR2_X1   g064(.A1(new_n202), .A2(new_n206), .ZN(new_n251));
  AOI21_X1  g065(.A(new_n250), .B1(new_n251), .B2(KEYINPUT82), .ZN(new_n252));
  AOI21_X1  g066(.A(new_n249), .B1(new_n252), .B2(new_n207), .ZN(new_n253));
  OAI211_X1 g067(.A(KEYINPUT83), .B(new_n242), .C1(new_n253), .C2(new_n191), .ZN(new_n254));
  INV_X1    g068(.A(KEYINPUT83), .ZN(new_n255));
  OAI21_X1  g069(.A(new_n255), .B1(new_n235), .B2(new_n243), .ZN(new_n256));
  NOR2_X1   g070(.A1(G475), .A2(G902), .ZN(new_n257));
  NAND3_X1  g071(.A1(new_n254), .A2(new_n256), .A3(new_n257), .ZN(new_n258));
  XOR2_X1   g072(.A(KEYINPUT81), .B(KEYINPUT20), .Z(new_n259));
  INV_X1    g073(.A(new_n259), .ZN(new_n260));
  AOI21_X1  g074(.A(new_n248), .B1(new_n258), .B2(new_n260), .ZN(new_n261));
  INV_X1    g075(.A(G475), .ZN(new_n262));
  OAI21_X1  g076(.A(new_n234), .B1(new_n237), .B2(new_n241), .ZN(new_n263));
  INV_X1    g077(.A(new_n191), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  INV_X1    g079(.A(KEYINPUT85), .ZN(new_n266));
  NOR2_X1   g080(.A1(new_n265), .A2(new_n266), .ZN(new_n267));
  NOR2_X1   g081(.A1(new_n267), .A2(G902), .ZN(new_n268));
  NAND3_X1  g082(.A1(new_n265), .A2(new_n266), .A3(new_n242), .ZN(new_n269));
  AOI21_X1  g083(.A(new_n262), .B1(new_n268), .B2(new_n269), .ZN(new_n270));
  OAI21_X1  g084(.A(new_n187), .B1(new_n261), .B2(new_n270), .ZN(new_n271));
  AND2_X1   g085(.A1(new_n246), .A2(new_n247), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n258), .A2(new_n260), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  INV_X1    g088(.A(new_n270), .ZN(new_n275));
  NAND3_X1  g089(.A1(new_n274), .A2(KEYINPUT86), .A3(new_n275), .ZN(new_n276));
  XNOR2_X1  g090(.A(KEYINPUT87), .B(G122), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n277), .A2(G116), .ZN(new_n278));
  INV_X1    g092(.A(G116), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n279), .A2(G122), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n278), .A2(new_n280), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n281), .A2(G107), .ZN(new_n282));
  INV_X1    g096(.A(G107), .ZN(new_n283));
  NAND3_X1  g097(.A1(new_n278), .A2(new_n283), .A3(new_n280), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n282), .A2(new_n284), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n212), .A2(G128), .ZN(new_n286));
  INV_X1    g100(.A(G128), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n287), .A2(G143), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n286), .A2(new_n288), .ZN(new_n289));
  INV_X1    g103(.A(new_n289), .ZN(new_n290));
  INV_X1    g104(.A(G134), .ZN(new_n291));
  INV_X1    g105(.A(KEYINPUT13), .ZN(new_n292));
  AOI21_X1  g106(.A(new_n291), .B1(new_n288), .B2(new_n292), .ZN(new_n293));
  OR2_X1    g107(.A1(new_n290), .A2(new_n293), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n290), .A2(new_n293), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n285), .A2(new_n296), .ZN(new_n297));
  XNOR2_X1  g111(.A(KEYINPUT9), .B(G234), .ZN(new_n298));
  INV_X1    g112(.A(G217), .ZN(new_n299));
  NOR3_X1   g113(.A1(new_n298), .A2(new_n299), .A3(G953), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n280), .A2(KEYINPUT14), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n301), .A2(KEYINPUT88), .ZN(new_n302));
  INV_X1    g116(.A(KEYINPUT88), .ZN(new_n303));
  NAND3_X1  g117(.A1(new_n280), .A2(new_n303), .A3(KEYINPUT14), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n302), .A2(new_n304), .ZN(new_n305));
  NOR2_X1   g119(.A1(new_n280), .A2(KEYINPUT14), .ZN(new_n306));
  AOI21_X1  g120(.A(new_n306), .B1(G116), .B2(new_n277), .ZN(new_n307));
  AOI21_X1  g121(.A(new_n283), .B1(new_n305), .B2(new_n307), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n289), .A2(new_n291), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n290), .A2(G134), .ZN(new_n310));
  NAND3_X1  g124(.A1(new_n284), .A2(new_n309), .A3(new_n310), .ZN(new_n311));
  OAI211_X1 g125(.A(new_n297), .B(new_n300), .C1(new_n308), .C2(new_n311), .ZN(new_n312));
  INV_X1    g126(.A(new_n300), .ZN(new_n313));
  NOR2_X1   g127(.A1(new_n308), .A2(new_n311), .ZN(new_n314));
  AOI22_X1  g128(.A1(new_n282), .A2(new_n284), .B1(new_n294), .B2(new_n295), .ZN(new_n315));
  OAI21_X1  g129(.A(new_n313), .B1(new_n314), .B2(new_n315), .ZN(new_n316));
  AOI21_X1  g130(.A(G902), .B1(new_n312), .B2(new_n316), .ZN(new_n317));
  INV_X1    g131(.A(G478), .ZN(new_n318));
  NOR2_X1   g132(.A1(new_n318), .A2(KEYINPUT15), .ZN(new_n319));
  XNOR2_X1  g133(.A(new_n317), .B(new_n319), .ZN(new_n320));
  INV_X1    g134(.A(new_n320), .ZN(new_n321));
  INV_X1    g135(.A(G952), .ZN(new_n322));
  NOR2_X1   g136(.A1(new_n322), .A2(G953), .ZN(new_n323));
  NAND2_X1  g137(.A1(G234), .A2(G237), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n323), .A2(new_n324), .ZN(new_n325));
  XNOR2_X1  g139(.A(KEYINPUT21), .B(G898), .ZN(new_n326));
  INV_X1    g140(.A(new_n326), .ZN(new_n327));
  NAND3_X1  g141(.A1(new_n324), .A2(G902), .A3(G953), .ZN(new_n328));
  OAI21_X1  g142(.A(new_n325), .B1(new_n327), .B2(new_n328), .ZN(new_n329));
  INV_X1    g143(.A(new_n329), .ZN(new_n330));
  NOR2_X1   g144(.A1(new_n321), .A2(new_n330), .ZN(new_n331));
  AND3_X1   g145(.A1(new_n271), .A2(new_n276), .A3(new_n331), .ZN(new_n332));
  OAI21_X1  g146(.A(G210), .B1(G237), .B2(G902), .ZN(new_n333));
  INV_X1    g147(.A(new_n333), .ZN(new_n334));
  NOR2_X1   g148(.A1(new_n220), .A2(G143), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n335), .A2(KEYINPUT1), .ZN(new_n336));
  XNOR2_X1  g150(.A(G143), .B(G146), .ZN(new_n337));
  OAI21_X1  g151(.A(new_n336), .B1(new_n337), .B2(G128), .ZN(new_n338));
  NOR2_X1   g152(.A1(new_n287), .A2(KEYINPUT1), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n220), .A2(G143), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n212), .A2(G146), .ZN(new_n341));
  AND3_X1   g155(.A1(new_n339), .A2(new_n340), .A3(new_n341), .ZN(new_n342));
  NOR3_X1   g156(.A1(new_n338), .A2(new_n342), .A3(G125), .ZN(new_n343));
  XNOR2_X1  g157(.A(KEYINPUT0), .B(G128), .ZN(new_n344));
  OAI21_X1  g158(.A(KEYINPUT64), .B1(new_n337), .B2(new_n344), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n340), .A2(new_n341), .ZN(new_n346));
  INV_X1    g160(.A(KEYINPUT64), .ZN(new_n347));
  NAND2_X1  g161(.A1(KEYINPUT0), .A2(G128), .ZN(new_n348));
  OR2_X1    g162(.A1(KEYINPUT0), .A2(G128), .ZN(new_n349));
  NAND4_X1  g163(.A1(new_n346), .A2(new_n347), .A3(new_n348), .A4(new_n349), .ZN(new_n350));
  AND2_X1   g164(.A1(KEYINPUT0), .A2(G128), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n337), .A2(new_n351), .ZN(new_n352));
  NAND3_X1  g166(.A1(new_n345), .A2(new_n350), .A3(new_n352), .ZN(new_n353));
  AOI21_X1  g167(.A(new_n343), .B1(G125), .B2(new_n353), .ZN(new_n354));
  XOR2_X1   g168(.A(KEYINPUT78), .B(G224), .Z(new_n355));
  NAND2_X1  g169(.A1(new_n355), .A2(new_n210), .ZN(new_n356));
  INV_X1    g170(.A(new_n356), .ZN(new_n357));
  XNOR2_X1  g171(.A(new_n354), .B(new_n357), .ZN(new_n358));
  OAI21_X1  g172(.A(KEYINPUT75), .B1(new_n283), .B2(G104), .ZN(new_n359));
  INV_X1    g173(.A(KEYINPUT75), .ZN(new_n360));
  NAND3_X1  g174(.A1(new_n360), .A2(new_n190), .A3(G107), .ZN(new_n361));
  INV_X1    g175(.A(G101), .ZN(new_n362));
  AND3_X1   g176(.A1(new_n359), .A2(new_n361), .A3(new_n362), .ZN(new_n363));
  NAND3_X1  g177(.A1(new_n283), .A2(KEYINPUT74), .A3(G104), .ZN(new_n364));
  INV_X1    g178(.A(KEYINPUT3), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  NAND4_X1  g180(.A1(new_n283), .A2(KEYINPUT74), .A3(KEYINPUT3), .A4(G104), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n366), .A2(new_n367), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n363), .A2(new_n368), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n359), .A2(new_n361), .ZN(new_n370));
  AOI21_X1  g184(.A(new_n370), .B1(new_n366), .B2(new_n367), .ZN(new_n371));
  OAI211_X1 g185(.A(new_n369), .B(KEYINPUT4), .C1(new_n371), .C2(new_n362), .ZN(new_n372));
  AND2_X1   g186(.A1(new_n359), .A2(new_n361), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n368), .A2(new_n373), .ZN(new_n374));
  NOR2_X1   g188(.A1(new_n362), .A2(KEYINPUT4), .ZN(new_n375));
  INV_X1    g189(.A(G119), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n376), .A2(G116), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n279), .A2(G119), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n377), .A2(new_n378), .ZN(new_n379));
  XNOR2_X1  g193(.A(KEYINPUT2), .B(G113), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n379), .A2(new_n380), .ZN(new_n381));
  XOR2_X1   g195(.A(KEYINPUT2), .B(G113), .Z(new_n382));
  XNOR2_X1  g196(.A(G116), .B(G119), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n382), .A2(new_n383), .ZN(new_n384));
  AOI22_X1  g198(.A1(new_n374), .A2(new_n375), .B1(new_n381), .B2(new_n384), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n372), .A2(new_n385), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n283), .A2(G104), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n190), .A2(G107), .ZN(new_n388));
  AOI21_X1  g202(.A(new_n362), .B1(new_n387), .B2(new_n388), .ZN(new_n389));
  AOI21_X1  g203(.A(new_n389), .B1(new_n363), .B2(new_n368), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n383), .A2(KEYINPUT5), .ZN(new_n391));
  INV_X1    g205(.A(G113), .ZN(new_n392));
  NOR2_X1   g206(.A1(new_n279), .A2(G119), .ZN(new_n393));
  INV_X1    g207(.A(KEYINPUT5), .ZN(new_n394));
  AOI21_X1  g208(.A(new_n392), .B1(new_n393), .B2(new_n394), .ZN(new_n395));
  AOI22_X1  g209(.A1(new_n391), .A2(new_n395), .B1(new_n382), .B2(new_n383), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n390), .A2(new_n396), .ZN(new_n397));
  XNOR2_X1  g211(.A(G110), .B(G122), .ZN(new_n398));
  NAND3_X1  g212(.A1(new_n386), .A2(new_n397), .A3(new_n398), .ZN(new_n399));
  INV_X1    g213(.A(KEYINPUT6), .ZN(new_n400));
  NOR2_X1   g214(.A1(new_n400), .A2(KEYINPUT77), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n399), .A2(new_n401), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n386), .A2(new_n397), .ZN(new_n403));
  INV_X1    g217(.A(new_n398), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n403), .A2(new_n404), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n402), .A2(new_n405), .ZN(new_n406));
  NAND3_X1  g220(.A1(new_n403), .A2(new_n404), .A3(new_n401), .ZN(new_n407));
  AOI21_X1  g221(.A(new_n358), .B1(new_n406), .B2(new_n407), .ZN(new_n408));
  XOR2_X1   g222(.A(new_n398), .B(KEYINPUT8), .Z(new_n409));
  NOR2_X1   g223(.A1(new_n379), .A2(new_n394), .ZN(new_n410));
  OAI21_X1  g224(.A(G113), .B1(new_n377), .B2(KEYINPUT5), .ZN(new_n411));
  OAI21_X1  g225(.A(new_n384), .B1(new_n410), .B2(new_n411), .ZN(new_n412));
  NAND3_X1  g226(.A1(new_n359), .A2(new_n361), .A3(new_n362), .ZN(new_n413));
  AOI21_X1  g227(.A(new_n413), .B1(new_n366), .B2(new_n367), .ZN(new_n414));
  OAI21_X1  g228(.A(new_n412), .B1(new_n414), .B2(new_n389), .ZN(new_n415));
  AOI21_X1  g229(.A(new_n409), .B1(new_n415), .B2(new_n397), .ZN(new_n416));
  AND2_X1   g230(.A1(new_n356), .A2(KEYINPUT7), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n353), .A2(G125), .ZN(new_n418));
  NOR2_X1   g232(.A1(new_n338), .A2(new_n342), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n419), .A2(new_n194), .ZN(new_n420));
  AOI21_X1  g234(.A(new_n417), .B1(new_n418), .B2(new_n420), .ZN(new_n421));
  NOR2_X1   g235(.A1(new_n416), .A2(new_n421), .ZN(new_n422));
  INV_X1    g236(.A(KEYINPUT79), .ZN(new_n423));
  NAND4_X1  g237(.A1(new_n354), .A2(new_n423), .A3(KEYINPUT7), .A4(new_n356), .ZN(new_n424));
  NAND4_X1  g238(.A1(new_n418), .A2(new_n420), .A3(KEYINPUT7), .A4(new_n356), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n425), .A2(KEYINPUT79), .ZN(new_n426));
  NAND4_X1  g240(.A1(new_n422), .A2(new_n399), .A3(new_n424), .A4(new_n426), .ZN(new_n427));
  INV_X1    g241(.A(G902), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n427), .A2(new_n428), .ZN(new_n429));
  OAI21_X1  g243(.A(new_n334), .B1(new_n408), .B2(new_n429), .ZN(new_n430));
  INV_X1    g244(.A(new_n401), .ZN(new_n431));
  AOI22_X1  g245(.A1(new_n372), .A2(new_n385), .B1(new_n390), .B2(new_n396), .ZN(new_n432));
  AOI21_X1  g246(.A(new_n431), .B1(new_n432), .B2(new_n398), .ZN(new_n433));
  NOR2_X1   g247(.A1(new_n432), .A2(new_n398), .ZN(new_n434));
  OAI21_X1  g248(.A(new_n407), .B1(new_n433), .B2(new_n434), .ZN(new_n435));
  INV_X1    g249(.A(new_n358), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n435), .A2(new_n436), .ZN(new_n437));
  NAND4_X1  g251(.A1(new_n437), .A2(new_n428), .A3(new_n427), .A4(new_n333), .ZN(new_n438));
  INV_X1    g252(.A(KEYINPUT80), .ZN(new_n439));
  NAND3_X1  g253(.A1(new_n430), .A2(new_n438), .A3(new_n439), .ZN(new_n440));
  OAI21_X1  g254(.A(G214), .B1(G237), .B2(G902), .ZN(new_n441));
  AND2_X1   g255(.A1(new_n427), .A2(new_n428), .ZN(new_n442));
  NAND4_X1  g256(.A1(new_n442), .A2(KEYINPUT80), .A3(new_n437), .A4(new_n333), .ZN(new_n443));
  NAND3_X1  g257(.A1(new_n440), .A2(new_n441), .A3(new_n443), .ZN(new_n444));
  INV_X1    g258(.A(G469), .ZN(new_n445));
  INV_X1    g259(.A(KEYINPUT76), .ZN(new_n446));
  AOI21_X1  g260(.A(G128), .B1(new_n340), .B2(new_n341), .ZN(new_n447));
  AND3_X1   g261(.A1(new_n212), .A2(KEYINPUT1), .A3(G146), .ZN(new_n448));
  OAI21_X1  g262(.A(new_n446), .B1(new_n447), .B2(new_n448), .ZN(new_n449));
  INV_X1    g263(.A(new_n342), .ZN(new_n450));
  OAI211_X1 g264(.A(new_n336), .B(KEYINPUT76), .C1(new_n337), .C2(G128), .ZN(new_n451));
  NAND3_X1  g265(.A1(new_n449), .A2(new_n450), .A3(new_n451), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n452), .A2(new_n390), .ZN(new_n453));
  OAI21_X1  g267(.A(new_n419), .B1(new_n414), .B2(new_n389), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  INV_X1    g269(.A(KEYINPUT11), .ZN(new_n456));
  OAI21_X1  g270(.A(new_n456), .B1(new_n291), .B2(G137), .ZN(new_n457));
  INV_X1    g271(.A(G137), .ZN(new_n458));
  NAND3_X1  g272(.A1(new_n458), .A2(KEYINPUT11), .A3(G134), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n291), .A2(G137), .ZN(new_n460));
  NAND3_X1  g274(.A1(new_n457), .A2(new_n459), .A3(new_n460), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n461), .A2(G131), .ZN(new_n462));
  NAND4_X1  g276(.A1(new_n457), .A2(new_n459), .A3(new_n208), .A4(new_n460), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  AOI21_X1  g278(.A(KEYINPUT12), .B1(new_n455), .B2(new_n464), .ZN(new_n465));
  INV_X1    g279(.A(KEYINPUT12), .ZN(new_n466));
  AND2_X1   g280(.A1(new_n462), .A2(new_n463), .ZN(new_n467));
  AOI211_X1 g281(.A(new_n466), .B(new_n467), .C1(new_n453), .C2(new_n454), .ZN(new_n468));
  NOR2_X1   g282(.A1(new_n465), .A2(new_n468), .ZN(new_n469));
  INV_X1    g283(.A(KEYINPUT10), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n453), .A2(new_n470), .ZN(new_n471));
  INV_X1    g285(.A(new_n353), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n374), .A2(new_n375), .ZN(new_n473));
  NAND3_X1  g287(.A1(new_n372), .A2(new_n472), .A3(new_n473), .ZN(new_n474));
  OAI211_X1 g288(.A(new_n390), .B(KEYINPUT10), .C1(new_n338), .C2(new_n342), .ZN(new_n475));
  NAND4_X1  g289(.A1(new_n471), .A2(new_n474), .A3(new_n467), .A4(new_n475), .ZN(new_n476));
  XNOR2_X1  g290(.A(G110), .B(G140), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n210), .A2(G227), .ZN(new_n478));
  XNOR2_X1  g292(.A(new_n477), .B(new_n478), .ZN(new_n479));
  XNOR2_X1  g293(.A(KEYINPUT72), .B(KEYINPUT73), .ZN(new_n480));
  XNOR2_X1  g294(.A(new_n479), .B(new_n480), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n476), .A2(new_n481), .ZN(new_n482));
  NOR2_X1   g296(.A1(new_n469), .A2(new_n482), .ZN(new_n483));
  NAND3_X1  g297(.A1(new_n471), .A2(new_n474), .A3(new_n475), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n484), .A2(new_n464), .ZN(new_n485));
  AOI21_X1  g299(.A(new_n481), .B1(new_n485), .B2(new_n476), .ZN(new_n486));
  OAI211_X1 g300(.A(new_n445), .B(new_n428), .C1(new_n483), .C2(new_n486), .ZN(new_n487));
  OAI21_X1  g301(.A(new_n476), .B1(new_n465), .B2(new_n468), .ZN(new_n488));
  INV_X1    g302(.A(new_n481), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  NAND3_X1  g304(.A1(new_n485), .A2(new_n476), .A3(new_n481), .ZN(new_n491));
  NAND3_X1  g305(.A1(new_n490), .A2(G469), .A3(new_n491), .ZN(new_n492));
  NAND2_X1  g306(.A1(G469), .A2(G902), .ZN(new_n493));
  NAND3_X1  g307(.A1(new_n487), .A2(new_n492), .A3(new_n493), .ZN(new_n494));
  OAI21_X1  g308(.A(G221), .B1(new_n298), .B2(G902), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  NOR2_X1   g310(.A1(new_n444), .A2(new_n496), .ZN(new_n497));
  INV_X1    g311(.A(KEYINPUT32), .ZN(new_n498));
  XOR2_X1   g312(.A(KEYINPUT26), .B(G101), .Z(new_n499));
  NAND2_X1  g313(.A1(new_n214), .A2(G210), .ZN(new_n500));
  XNOR2_X1  g314(.A(new_n499), .B(new_n500), .ZN(new_n501));
  XNOR2_X1  g315(.A(KEYINPUT65), .B(KEYINPUT27), .ZN(new_n502));
  XNOR2_X1  g316(.A(new_n501), .B(new_n502), .ZN(new_n503));
  INV_X1    g317(.A(new_n503), .ZN(new_n504));
  INV_X1    g318(.A(KEYINPUT28), .ZN(new_n505));
  INV_X1    g319(.A(new_n460), .ZN(new_n506));
  NOR2_X1   g320(.A1(new_n291), .A2(G137), .ZN(new_n507));
  OAI21_X1  g321(.A(G131), .B1(new_n506), .B2(new_n507), .ZN(new_n508));
  OAI211_X1 g322(.A(new_n463), .B(new_n508), .C1(new_n338), .C2(new_n342), .ZN(new_n509));
  OAI21_X1  g323(.A(new_n509), .B1(new_n467), .B2(new_n353), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n384), .A2(new_n381), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  INV_X1    g326(.A(new_n511), .ZN(new_n513));
  OAI211_X1 g327(.A(new_n513), .B(new_n509), .C1(new_n467), .C2(new_n353), .ZN(new_n514));
  AOI21_X1  g328(.A(new_n505), .B1(new_n512), .B2(new_n514), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n514), .A2(new_n505), .ZN(new_n516));
  INV_X1    g330(.A(new_n516), .ZN(new_n517));
  OAI21_X1  g331(.A(KEYINPUT66), .B1(new_n515), .B2(new_n517), .ZN(new_n518));
  INV_X1    g332(.A(new_n514), .ZN(new_n519));
  AND3_X1   g333(.A1(new_n340), .A2(new_n341), .A3(new_n351), .ZN(new_n520));
  NOR2_X1   g334(.A1(new_n212), .A2(G146), .ZN(new_n521));
  OAI211_X1 g335(.A(new_n348), .B(new_n349), .C1(new_n521), .C2(new_n335), .ZN(new_n522));
  AOI21_X1  g336(.A(new_n520), .B1(new_n522), .B2(KEYINPUT64), .ZN(new_n523));
  NAND3_X1  g337(.A1(new_n464), .A2(new_n523), .A3(new_n350), .ZN(new_n524));
  AOI21_X1  g338(.A(new_n513), .B1(new_n524), .B2(new_n509), .ZN(new_n525));
  OAI21_X1  g339(.A(KEYINPUT28), .B1(new_n519), .B2(new_n525), .ZN(new_n526));
  INV_X1    g340(.A(KEYINPUT66), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n518), .A2(new_n528), .ZN(new_n529));
  INV_X1    g343(.A(KEYINPUT30), .ZN(new_n530));
  OAI211_X1 g344(.A(new_n530), .B(new_n509), .C1(new_n467), .C2(new_n353), .ZN(new_n531));
  INV_X1    g345(.A(new_n531), .ZN(new_n532));
  AOI21_X1  g346(.A(new_n530), .B1(new_n524), .B2(new_n509), .ZN(new_n533));
  OAI21_X1  g347(.A(new_n511), .B1(new_n532), .B2(new_n533), .ZN(new_n534));
  NAND3_X1  g348(.A1(new_n534), .A2(new_n503), .A3(new_n514), .ZN(new_n535));
  INV_X1    g349(.A(KEYINPUT31), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  NAND4_X1  g351(.A1(new_n534), .A2(KEYINPUT31), .A3(new_n503), .A4(new_n514), .ZN(new_n538));
  AOI22_X1  g352(.A1(new_n504), .A2(new_n529), .B1(new_n537), .B2(new_n538), .ZN(new_n539));
  NOR2_X1   g353(.A1(G472), .A2(G902), .ZN(new_n540));
  INV_X1    g354(.A(new_n540), .ZN(new_n541));
  OAI21_X1  g355(.A(new_n498), .B1(new_n539), .B2(new_n541), .ZN(new_n542));
  INV_X1    g356(.A(KEYINPUT29), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n510), .A2(KEYINPUT30), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n544), .A2(new_n531), .ZN(new_n545));
  AOI21_X1  g359(.A(new_n519), .B1(new_n545), .B2(new_n511), .ZN(new_n546));
  OAI21_X1  g360(.A(new_n543), .B1(new_n546), .B2(new_n503), .ZN(new_n547));
  AOI21_X1  g361(.A(new_n527), .B1(new_n526), .B2(new_n516), .ZN(new_n548));
  NOR2_X1   g362(.A1(new_n515), .A2(KEYINPUT66), .ZN(new_n549));
  NOR2_X1   g363(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  AOI21_X1  g364(.A(new_n547), .B1(new_n550), .B2(new_n503), .ZN(new_n551));
  INV_X1    g365(.A(KEYINPUT67), .ZN(new_n552));
  NAND3_X1  g366(.A1(new_n512), .A2(new_n552), .A3(new_n514), .ZN(new_n553));
  OAI211_X1 g367(.A(new_n553), .B(KEYINPUT28), .C1(new_n552), .C2(new_n512), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n554), .A2(new_n516), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n503), .A2(KEYINPUT29), .ZN(new_n556));
  OAI21_X1  g370(.A(new_n428), .B1(new_n555), .B2(new_n556), .ZN(new_n557));
  OAI21_X1  g371(.A(G472), .B1(new_n551), .B2(new_n557), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n537), .A2(new_n538), .ZN(new_n559));
  OAI21_X1  g373(.A(new_n504), .B1(new_n548), .B2(new_n549), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  NAND3_X1  g375(.A1(new_n561), .A2(KEYINPUT32), .A3(new_n540), .ZN(new_n562));
  NAND3_X1  g376(.A1(new_n542), .A2(new_n558), .A3(new_n562), .ZN(new_n563));
  AOI21_X1  g377(.A(new_n299), .B1(G234), .B2(new_n428), .ZN(new_n564));
  NOR2_X1   g378(.A1(new_n564), .A2(G902), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n239), .A2(new_n224), .ZN(new_n566));
  OAI211_X1 g380(.A(new_n287), .B(G119), .C1(KEYINPUT68), .C2(KEYINPUT23), .ZN(new_n567));
  INV_X1    g381(.A(KEYINPUT23), .ZN(new_n568));
  AOI21_X1  g382(.A(new_n568), .B1(new_n376), .B2(G128), .ZN(new_n569));
  INV_X1    g383(.A(KEYINPUT68), .ZN(new_n570));
  OAI21_X1  g384(.A(new_n570), .B1(new_n376), .B2(G128), .ZN(new_n571));
  OAI21_X1  g385(.A(new_n567), .B1(new_n569), .B2(new_n571), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n572), .A2(G110), .ZN(new_n573));
  XOR2_X1   g387(.A(KEYINPUT24), .B(G110), .Z(new_n574));
  XNOR2_X1  g388(.A(G119), .B(G128), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  NAND3_X1  g390(.A1(new_n566), .A2(new_n573), .A3(new_n576), .ZN(new_n577));
  OAI22_X1  g391(.A1(new_n572), .A2(G110), .B1(new_n575), .B2(new_n574), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n227), .A2(new_n220), .ZN(new_n579));
  NAND3_X1  g393(.A1(new_n578), .A2(new_n224), .A3(new_n579), .ZN(new_n580));
  NAND3_X1  g394(.A1(new_n210), .A2(G221), .A3(G234), .ZN(new_n581));
  XNOR2_X1  g395(.A(new_n581), .B(KEYINPUT69), .ZN(new_n582));
  XNOR2_X1  g396(.A(KEYINPUT22), .B(G137), .ZN(new_n583));
  XNOR2_X1  g397(.A(new_n582), .B(new_n583), .ZN(new_n584));
  AND3_X1   g398(.A1(new_n577), .A2(new_n580), .A3(new_n584), .ZN(new_n585));
  AOI21_X1  g399(.A(new_n584), .B1(new_n577), .B2(new_n580), .ZN(new_n586));
  OAI21_X1  g400(.A(new_n565), .B1(new_n585), .B2(new_n586), .ZN(new_n587));
  INV_X1    g401(.A(KEYINPUT71), .ZN(new_n588));
  XNOR2_X1  g402(.A(new_n587), .B(new_n588), .ZN(new_n589));
  INV_X1    g403(.A(KEYINPUT25), .ZN(new_n590));
  AOI21_X1  g404(.A(G902), .B1(new_n590), .B2(KEYINPUT70), .ZN(new_n591));
  OAI21_X1  g405(.A(new_n591), .B1(new_n585), .B2(new_n586), .ZN(new_n592));
  NOR2_X1   g406(.A1(new_n590), .A2(KEYINPUT70), .ZN(new_n593));
  OR2_X1    g407(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  INV_X1    g408(.A(new_n564), .ZN(new_n595));
  AOI21_X1  g409(.A(new_n595), .B1(new_n592), .B2(new_n593), .ZN(new_n596));
  AOI21_X1  g410(.A(new_n589), .B1(new_n594), .B2(new_n596), .ZN(new_n597));
  NAND4_X1  g411(.A1(new_n332), .A2(new_n497), .A3(new_n563), .A4(new_n597), .ZN(new_n598));
  XNOR2_X1  g412(.A(new_n598), .B(G101), .ZN(G3));
  OAI211_X1 g413(.A(KEYINPUT91), .B(new_n313), .C1(new_n314), .C2(new_n315), .ZN(new_n600));
  NAND3_X1  g414(.A1(new_n600), .A2(new_n312), .A3(KEYINPUT33), .ZN(new_n601));
  OAI21_X1  g415(.A(new_n297), .B1(new_n308), .B2(new_n311), .ZN(new_n602));
  AOI21_X1  g416(.A(KEYINPUT91), .B1(new_n602), .B2(new_n313), .ZN(new_n603));
  OAI21_X1  g417(.A(KEYINPUT92), .B1(new_n601), .B2(new_n603), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n312), .A2(new_n316), .ZN(new_n605));
  INV_X1    g419(.A(KEYINPUT33), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  NOR2_X1   g421(.A1(new_n314), .A2(new_n315), .ZN(new_n608));
  AOI21_X1  g422(.A(new_n606), .B1(new_n608), .B2(new_n300), .ZN(new_n609));
  INV_X1    g423(.A(KEYINPUT91), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n316), .A2(new_n610), .ZN(new_n611));
  INV_X1    g425(.A(KEYINPUT92), .ZN(new_n612));
  NAND4_X1  g426(.A1(new_n609), .A2(new_n611), .A3(new_n612), .A4(new_n600), .ZN(new_n613));
  NOR2_X1   g427(.A1(new_n318), .A2(G902), .ZN(new_n614));
  NAND4_X1  g428(.A1(new_n604), .A2(new_n607), .A3(new_n613), .A4(new_n614), .ZN(new_n615));
  OR2_X1    g429(.A1(new_n317), .A2(G478), .ZN(new_n616));
  AND2_X1   g430(.A1(new_n615), .A2(new_n616), .ZN(new_n617));
  AOI21_X1  g431(.A(new_n617), .B1(new_n271), .B2(new_n276), .ZN(new_n618));
  INV_X1    g432(.A(KEYINPUT89), .ZN(new_n619));
  AND3_X1   g433(.A1(new_n430), .A2(new_n438), .A3(new_n619), .ZN(new_n620));
  OAI211_X1 g434(.A(KEYINPUT89), .B(new_n334), .C1(new_n408), .C2(new_n429), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n621), .A2(new_n441), .ZN(new_n622));
  OAI21_X1  g436(.A(KEYINPUT90), .B1(new_n620), .B2(new_n622), .ZN(new_n623));
  INV_X1    g437(.A(new_n441), .ZN(new_n624));
  AOI21_X1  g438(.A(new_n333), .B1(new_n442), .B2(new_n437), .ZN(new_n625));
  AOI21_X1  g439(.A(new_n624), .B1(new_n625), .B2(KEYINPUT89), .ZN(new_n626));
  INV_X1    g440(.A(KEYINPUT90), .ZN(new_n627));
  NAND3_X1  g441(.A1(new_n430), .A2(new_n438), .A3(new_n619), .ZN(new_n628));
  NAND3_X1  g442(.A1(new_n626), .A2(new_n627), .A3(new_n628), .ZN(new_n629));
  NAND4_X1  g443(.A1(new_n618), .A2(new_n329), .A3(new_n623), .A4(new_n629), .ZN(new_n630));
  INV_X1    g444(.A(new_n630), .ZN(new_n631));
  NAND3_X1  g445(.A1(new_n494), .A2(new_n597), .A3(new_n495), .ZN(new_n632));
  AOI21_X1  g446(.A(G902), .B1(new_n559), .B2(new_n560), .ZN(new_n633));
  INV_X1    g447(.A(G472), .ZN(new_n634));
  OAI22_X1  g448(.A1(new_n633), .A2(new_n634), .B1(new_n539), .B2(new_n541), .ZN(new_n635));
  NOR2_X1   g449(.A1(new_n632), .A2(new_n635), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n631), .A2(new_n636), .ZN(new_n637));
  XOR2_X1   g451(.A(KEYINPUT34), .B(G104), .Z(new_n638));
  XNOR2_X1  g452(.A(new_n637), .B(new_n638), .ZN(G6));
  NAND2_X1  g453(.A1(new_n321), .A2(new_n275), .ZN(new_n640));
  NAND4_X1  g454(.A1(new_n254), .A2(new_n256), .A3(new_n257), .A4(new_n259), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n273), .A2(new_n641), .ZN(new_n642));
  INV_X1    g456(.A(KEYINPUT93), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  NAND3_X1  g458(.A1(new_n273), .A2(KEYINPUT93), .A3(new_n641), .ZN(new_n645));
  AOI21_X1  g459(.A(new_n640), .B1(new_n644), .B2(new_n645), .ZN(new_n646));
  NAND4_X1  g460(.A1(new_n623), .A2(new_n629), .A3(new_n646), .A4(new_n329), .ZN(new_n647));
  AND2_X1   g461(.A1(new_n647), .A2(KEYINPUT94), .ZN(new_n648));
  NOR2_X1   g462(.A1(new_n647), .A2(KEYINPUT94), .ZN(new_n649));
  OAI21_X1  g463(.A(new_n636), .B1(new_n648), .B2(new_n649), .ZN(new_n650));
  XOR2_X1   g464(.A(KEYINPUT35), .B(G107), .Z(new_n651));
  XNOR2_X1  g465(.A(new_n650), .B(new_n651), .ZN(G9));
  INV_X1    g466(.A(new_n635), .ZN(new_n653));
  NAND2_X1  g467(.A1(new_n594), .A2(new_n596), .ZN(new_n654));
  NAND2_X1  g468(.A1(new_n577), .A2(new_n580), .ZN(new_n655));
  NOR2_X1   g469(.A1(new_n584), .A2(KEYINPUT36), .ZN(new_n656));
  XNOR2_X1  g470(.A(new_n655), .B(new_n656), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n657), .A2(new_n565), .ZN(new_n658));
  AND2_X1   g472(.A1(new_n654), .A2(new_n658), .ZN(new_n659));
  INV_X1    g473(.A(new_n659), .ZN(new_n660));
  NAND4_X1  g474(.A1(new_n332), .A2(new_n497), .A3(new_n653), .A4(new_n660), .ZN(new_n661));
  XNOR2_X1  g475(.A(KEYINPUT37), .B(G110), .ZN(new_n662));
  XNOR2_X1  g476(.A(new_n662), .B(KEYINPUT95), .ZN(new_n663));
  XNOR2_X1  g477(.A(new_n661), .B(new_n663), .ZN(G12));
  INV_X1    g478(.A(new_n496), .ZN(new_n665));
  AND3_X1   g479(.A1(new_n563), .A2(new_n665), .A3(new_n660), .ZN(new_n666));
  NOR3_X1   g480(.A1(new_n620), .A2(KEYINPUT90), .A3(new_n622), .ZN(new_n667));
  AOI21_X1  g481(.A(new_n627), .B1(new_n626), .B2(new_n628), .ZN(new_n668));
  NOR2_X1   g482(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  XOR2_X1   g483(.A(new_n325), .B(KEYINPUT96), .Z(new_n670));
  OAI21_X1  g484(.A(new_n670), .B1(G900), .B2(new_n328), .ZN(new_n671));
  NAND2_X1  g485(.A1(new_n646), .A2(new_n671), .ZN(new_n672));
  INV_X1    g486(.A(new_n672), .ZN(new_n673));
  NAND3_X1  g487(.A1(new_n666), .A2(new_n669), .A3(new_n673), .ZN(new_n674));
  XNOR2_X1  g488(.A(KEYINPUT97), .B(G128), .ZN(new_n675));
  XNOR2_X1  g489(.A(new_n674), .B(new_n675), .ZN(G30));
  NAND2_X1  g490(.A1(new_n271), .A2(new_n276), .ZN(new_n677));
  NAND2_X1  g491(.A1(new_n677), .A2(new_n321), .ZN(new_n678));
  NOR2_X1   g492(.A1(new_n678), .A2(new_n624), .ZN(new_n679));
  NAND2_X1  g493(.A1(new_n440), .A2(new_n443), .ZN(new_n680));
  INV_X1    g494(.A(KEYINPUT38), .ZN(new_n681));
  XNOR2_X1  g495(.A(new_n680), .B(new_n681), .ZN(new_n682));
  AOI21_X1  g496(.A(KEYINPUT32), .B1(new_n561), .B2(new_n540), .ZN(new_n683));
  AOI211_X1 g497(.A(new_n498), .B(new_n541), .C1(new_n559), .C2(new_n560), .ZN(new_n684));
  NOR2_X1   g498(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  OAI21_X1  g499(.A(new_n553), .B1(new_n552), .B2(new_n512), .ZN(new_n686));
  OAI211_X1 g500(.A(new_n535), .B(G472), .C1(new_n686), .C2(new_n503), .ZN(new_n687));
  NAND2_X1  g501(.A1(G472), .A2(G902), .ZN(new_n688));
  NAND2_X1  g502(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  XNOR2_X1  g503(.A(new_n689), .B(KEYINPUT98), .ZN(new_n690));
  AOI21_X1  g504(.A(new_n660), .B1(new_n685), .B2(new_n690), .ZN(new_n691));
  XNOR2_X1  g505(.A(new_n671), .B(KEYINPUT39), .ZN(new_n692));
  NAND3_X1  g506(.A1(new_n494), .A2(new_n495), .A3(new_n692), .ZN(new_n693));
  INV_X1    g507(.A(KEYINPUT40), .ZN(new_n694));
  XNOR2_X1  g508(.A(new_n693), .B(new_n694), .ZN(new_n695));
  NAND4_X1  g509(.A1(new_n679), .A2(new_n682), .A3(new_n691), .A4(new_n695), .ZN(new_n696));
  XNOR2_X1  g510(.A(new_n696), .B(KEYINPUT99), .ZN(new_n697));
  XNOR2_X1  g511(.A(new_n697), .B(G143), .ZN(G45));
  INV_X1    g512(.A(new_n671), .ZN(new_n699));
  AOI211_X1 g513(.A(new_n617), .B(new_n699), .C1(new_n271), .C2(new_n276), .ZN(new_n700));
  NAND3_X1  g514(.A1(new_n666), .A2(new_n669), .A3(new_n700), .ZN(new_n701));
  XOR2_X1   g515(.A(KEYINPUT100), .B(G146), .Z(new_n702));
  XNOR2_X1  g516(.A(new_n701), .B(new_n702), .ZN(G48));
  OAI21_X1  g517(.A(new_n428), .B1(new_n483), .B2(new_n486), .ZN(new_n704));
  NAND2_X1  g518(.A1(new_n704), .A2(G469), .ZN(new_n705));
  NAND3_X1  g519(.A1(new_n705), .A2(new_n495), .A3(new_n487), .ZN(new_n706));
  NAND2_X1  g520(.A1(new_n706), .A2(KEYINPUT101), .ZN(new_n707));
  INV_X1    g521(.A(KEYINPUT101), .ZN(new_n708));
  NAND4_X1  g522(.A1(new_n705), .A2(new_n708), .A3(new_n495), .A4(new_n487), .ZN(new_n709));
  NAND4_X1  g523(.A1(new_n563), .A2(new_n707), .A3(new_n597), .A4(new_n709), .ZN(new_n710));
  NOR2_X1   g524(.A1(new_n630), .A2(new_n710), .ZN(new_n711));
  XOR2_X1   g525(.A(KEYINPUT41), .B(G113), .Z(new_n712));
  XNOR2_X1  g526(.A(new_n711), .B(new_n712), .ZN(G15));
  INV_X1    g527(.A(new_n710), .ZN(new_n714));
  OAI21_X1  g528(.A(new_n714), .B1(new_n648), .B2(new_n649), .ZN(new_n715));
  XNOR2_X1  g529(.A(new_n715), .B(G116), .ZN(G18));
  NOR3_X1   g530(.A1(new_n667), .A2(new_n668), .A3(new_n706), .ZN(new_n717));
  INV_X1    g531(.A(KEYINPUT102), .ZN(new_n718));
  AOI21_X1  g532(.A(new_n659), .B1(new_n685), .B2(new_n558), .ZN(new_n719));
  NAND4_X1  g533(.A1(new_n717), .A2(new_n718), .A3(new_n332), .A4(new_n719), .ZN(new_n720));
  AOI211_X1 g534(.A(new_n187), .B(new_n270), .C1(new_n272), .C2(new_n273), .ZN(new_n721));
  AOI21_X1  g535(.A(KEYINPUT86), .B1(new_n274), .B2(new_n275), .ZN(new_n722));
  NOR2_X1   g536(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  NAND4_X1  g537(.A1(new_n723), .A2(new_n563), .A3(new_n331), .A4(new_n660), .ZN(new_n724));
  INV_X1    g538(.A(new_n706), .ZN(new_n725));
  NAND3_X1  g539(.A1(new_n623), .A2(new_n629), .A3(new_n725), .ZN(new_n726));
  OAI21_X1  g540(.A(KEYINPUT102), .B1(new_n724), .B2(new_n726), .ZN(new_n727));
  NAND2_X1  g541(.A1(new_n720), .A2(new_n727), .ZN(new_n728));
  XNOR2_X1  g542(.A(new_n728), .B(G119), .ZN(G21));
  NAND4_X1  g543(.A1(new_n623), .A2(new_n677), .A3(new_n321), .A4(new_n629), .ZN(new_n730));
  INV_X1    g544(.A(new_n730), .ZN(new_n731));
  NAND3_X1  g545(.A1(new_n707), .A2(new_n329), .A3(new_n709), .ZN(new_n732));
  OAI21_X1  g546(.A(G472), .B1(new_n539), .B2(G902), .ZN(new_n733));
  XOR2_X1   g547(.A(new_n540), .B(KEYINPUT103), .Z(new_n734));
  INV_X1    g548(.A(new_n734), .ZN(new_n735));
  NAND2_X1  g549(.A1(new_n555), .A2(new_n504), .ZN(new_n736));
  AOI21_X1  g550(.A(new_n735), .B1(new_n736), .B2(new_n559), .ZN(new_n737));
  INV_X1    g551(.A(new_n737), .ZN(new_n738));
  NAND3_X1  g552(.A1(new_n733), .A2(new_n738), .A3(new_n597), .ZN(new_n739));
  NOR2_X1   g553(.A1(new_n732), .A2(new_n739), .ZN(new_n740));
  NAND2_X1  g554(.A1(new_n731), .A2(new_n740), .ZN(new_n741));
  XNOR2_X1  g555(.A(new_n741), .B(G122), .ZN(G24));
  NAND3_X1  g556(.A1(new_n733), .A2(new_n660), .A3(new_n738), .ZN(new_n743));
  INV_X1    g557(.A(new_n743), .ZN(new_n744));
  NAND4_X1  g558(.A1(new_n669), .A2(new_n700), .A3(new_n725), .A4(new_n744), .ZN(new_n745));
  XNOR2_X1  g559(.A(new_n745), .B(G125), .ZN(G27));
  INV_X1    g560(.A(new_n495), .ZN(new_n747));
  NAND4_X1  g561(.A1(new_n490), .A2(KEYINPUT104), .A3(G469), .A4(new_n491), .ZN(new_n748));
  AND3_X1   g562(.A1(new_n487), .A2(new_n493), .A3(new_n748), .ZN(new_n749));
  INV_X1    g563(.A(KEYINPUT104), .ZN(new_n750));
  NAND2_X1  g564(.A1(new_n492), .A2(new_n750), .ZN(new_n751));
  AOI21_X1  g565(.A(new_n747), .B1(new_n749), .B2(new_n751), .ZN(new_n752));
  AOI21_X1  g566(.A(new_n624), .B1(new_n440), .B2(new_n443), .ZN(new_n753));
  NAND4_X1  g567(.A1(new_n752), .A2(new_n563), .A3(new_n597), .A4(new_n753), .ZN(new_n754));
  NAND2_X1  g568(.A1(new_n615), .A2(new_n616), .ZN(new_n755));
  OAI211_X1 g569(.A(new_n755), .B(new_n671), .C1(new_n721), .C2(new_n722), .ZN(new_n756));
  NOR3_X1   g570(.A1(new_n754), .A2(KEYINPUT42), .A3(new_n756), .ZN(new_n757));
  INV_X1    g571(.A(KEYINPUT106), .ZN(new_n758));
  INV_X1    g572(.A(KEYINPUT105), .ZN(new_n759));
  AOI21_X1  g573(.A(new_n759), .B1(new_n542), .B2(new_n562), .ZN(new_n760));
  NOR2_X1   g574(.A1(new_n683), .A2(KEYINPUT105), .ZN(new_n761));
  OAI21_X1  g575(.A(new_n758), .B1(new_n760), .B2(new_n761), .ZN(new_n762));
  OAI21_X1  g576(.A(KEYINPUT105), .B1(new_n683), .B2(new_n684), .ZN(new_n763));
  NAND2_X1  g577(.A1(new_n542), .A2(new_n759), .ZN(new_n764));
  NAND3_X1  g578(.A1(new_n763), .A2(KEYINPUT106), .A3(new_n764), .ZN(new_n765));
  NAND3_X1  g579(.A1(new_n762), .A2(new_n765), .A3(new_n558), .ZN(new_n766));
  NAND2_X1  g580(.A1(new_n752), .A2(new_n753), .ZN(new_n767));
  NOR2_X1   g581(.A1(new_n767), .A2(new_n756), .ZN(new_n768));
  NAND3_X1  g582(.A1(new_n766), .A2(new_n597), .A3(new_n768), .ZN(new_n769));
  AOI21_X1  g583(.A(new_n757), .B1(new_n769), .B2(KEYINPUT42), .ZN(new_n770));
  XNOR2_X1  g584(.A(new_n770), .B(G131), .ZN(G33));
  INV_X1    g585(.A(new_n589), .ZN(new_n772));
  NAND2_X1  g586(.A1(new_n772), .A2(new_n654), .ZN(new_n773));
  AOI21_X1  g587(.A(new_n773), .B1(new_n685), .B2(new_n558), .ZN(new_n774));
  NAND4_X1  g588(.A1(new_n751), .A2(new_n487), .A3(new_n493), .A4(new_n748), .ZN(new_n775));
  AND4_X1   g589(.A1(new_n441), .A2(new_n680), .A3(new_n495), .A4(new_n775), .ZN(new_n776));
  NAND3_X1  g590(.A1(new_n673), .A2(new_n774), .A3(new_n776), .ZN(new_n777));
  XNOR2_X1  g591(.A(new_n777), .B(G134), .ZN(G36));
  INV_X1    g592(.A(new_n487), .ZN(new_n779));
  AND2_X1   g593(.A1(new_n490), .A2(new_n491), .ZN(new_n780));
  OAI21_X1  g594(.A(G469), .B1(new_n780), .B2(KEYINPUT45), .ZN(new_n781));
  NAND2_X1  g595(.A1(new_n781), .A2(KEYINPUT107), .ZN(new_n782));
  INV_X1    g596(.A(KEYINPUT107), .ZN(new_n783));
  OAI211_X1 g597(.A(new_n783), .B(G469), .C1(new_n780), .C2(KEYINPUT45), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n780), .A2(KEYINPUT45), .ZN(new_n785));
  NAND3_X1  g599(.A1(new_n782), .A2(new_n784), .A3(new_n785), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n786), .A2(new_n493), .ZN(new_n787));
  INV_X1    g601(.A(KEYINPUT46), .ZN(new_n788));
  AOI21_X1  g602(.A(new_n779), .B1(new_n787), .B2(new_n788), .ZN(new_n789));
  NAND3_X1  g603(.A1(new_n786), .A2(KEYINPUT46), .A3(new_n493), .ZN(new_n790));
  AOI21_X1  g604(.A(new_n747), .B1(new_n789), .B2(new_n790), .ZN(new_n791));
  AND2_X1   g605(.A1(new_n791), .A2(new_n692), .ZN(new_n792));
  XNOR2_X1  g606(.A(new_n753), .B(KEYINPUT108), .ZN(new_n793));
  NAND3_X1  g607(.A1(new_n271), .A2(new_n276), .A3(new_n755), .ZN(new_n794));
  OR2_X1    g608(.A1(new_n794), .A2(KEYINPUT43), .ZN(new_n795));
  NAND2_X1  g609(.A1(new_n794), .A2(KEYINPUT43), .ZN(new_n796));
  NOR2_X1   g610(.A1(new_n653), .A2(new_n659), .ZN(new_n797));
  NAND3_X1  g611(.A1(new_n795), .A2(new_n796), .A3(new_n797), .ZN(new_n798));
  NAND2_X1  g612(.A1(new_n798), .A2(KEYINPUT44), .ZN(new_n799));
  INV_X1    g613(.A(KEYINPUT44), .ZN(new_n800));
  NAND4_X1  g614(.A1(new_n795), .A2(new_n800), .A3(new_n796), .A4(new_n797), .ZN(new_n801));
  AOI21_X1  g615(.A(new_n793), .B1(new_n799), .B2(new_n801), .ZN(new_n802));
  NAND2_X1  g616(.A1(new_n792), .A2(new_n802), .ZN(new_n803));
  XNOR2_X1  g617(.A(new_n803), .B(G137), .ZN(G39));
  INV_X1    g618(.A(KEYINPUT109), .ZN(new_n805));
  NAND2_X1  g619(.A1(new_n805), .A2(KEYINPUT47), .ZN(new_n806));
  NAND2_X1  g620(.A1(new_n791), .A2(new_n806), .ZN(new_n807));
  INV_X1    g621(.A(new_n753), .ZN(new_n808));
  NOR4_X1   g622(.A1(new_n756), .A2(new_n808), .A3(new_n563), .A4(new_n597), .ZN(new_n809));
  XNOR2_X1  g623(.A(KEYINPUT109), .B(KEYINPUT47), .ZN(new_n810));
  OAI211_X1 g624(.A(new_n807), .B(new_n809), .C1(new_n791), .C2(new_n810), .ZN(new_n811));
  XNOR2_X1  g625(.A(new_n811), .B(G140), .ZN(G42));
  INV_X1    g626(.A(KEYINPUT51), .ZN(new_n813));
  INV_X1    g627(.A(new_n670), .ZN(new_n814));
  AOI21_X1  g628(.A(new_n634), .B1(new_n561), .B2(new_n428), .ZN(new_n815));
  NOR3_X1   g629(.A1(new_n815), .A2(new_n773), .A3(new_n737), .ZN(new_n816));
  NAND4_X1  g630(.A1(new_n795), .A2(new_n814), .A3(new_n816), .A4(new_n796), .ZN(new_n817));
  NOR2_X1   g631(.A1(new_n817), .A2(new_n706), .ZN(new_n818));
  INV_X1    g632(.A(KEYINPUT113), .ZN(new_n819));
  OAI21_X1  g633(.A(new_n624), .B1(new_n819), .B2(KEYINPUT50), .ZN(new_n820));
  NOR2_X1   g634(.A1(new_n682), .A2(new_n820), .ZN(new_n821));
  NAND2_X1  g635(.A1(new_n818), .A2(new_n821), .ZN(new_n822));
  NAND3_X1  g636(.A1(new_n822), .A2(new_n819), .A3(KEYINPUT50), .ZN(new_n823));
  NAND3_X1  g637(.A1(new_n795), .A2(new_n814), .A3(new_n796), .ZN(new_n824));
  NAND2_X1  g638(.A1(new_n753), .A2(new_n725), .ZN(new_n825));
  NAND2_X1  g639(.A1(new_n825), .A2(KEYINPUT114), .ZN(new_n826));
  INV_X1    g640(.A(KEYINPUT114), .ZN(new_n827));
  NAND3_X1  g641(.A1(new_n753), .A2(new_n725), .A3(new_n827), .ZN(new_n828));
  AND2_X1   g642(.A1(new_n826), .A2(new_n828), .ZN(new_n829));
  NOR3_X1   g643(.A1(new_n824), .A2(new_n829), .A3(new_n743), .ZN(new_n830));
  NOR2_X1   g644(.A1(new_n773), .A2(new_n325), .ZN(new_n831));
  NAND3_X1  g645(.A1(new_n685), .A2(new_n690), .A3(new_n831), .ZN(new_n832));
  NAND2_X1  g646(.A1(new_n723), .A2(new_n617), .ZN(new_n833));
  NOR3_X1   g647(.A1(new_n829), .A2(new_n832), .A3(new_n833), .ZN(new_n834));
  NOR2_X1   g648(.A1(new_n830), .A2(new_n834), .ZN(new_n835));
  NAND2_X1  g649(.A1(new_n819), .A2(KEYINPUT50), .ZN(new_n836));
  NAND3_X1  g650(.A1(new_n818), .A2(new_n821), .A3(new_n836), .ZN(new_n837));
  NAND3_X1  g651(.A1(new_n823), .A2(new_n835), .A3(new_n837), .ZN(new_n838));
  NOR2_X1   g652(.A1(new_n817), .A2(new_n793), .ZN(new_n839));
  INV_X1    g653(.A(new_n839), .ZN(new_n840));
  OAI21_X1  g654(.A(new_n807), .B1(new_n791), .B2(new_n810), .ZN(new_n841));
  AND2_X1   g655(.A1(new_n485), .A2(new_n476), .ZN(new_n842));
  OAI22_X1  g656(.A1(new_n842), .A2(new_n481), .B1(new_n469), .B2(new_n482), .ZN(new_n843));
  AOI21_X1  g657(.A(new_n445), .B1(new_n843), .B2(new_n428), .ZN(new_n844));
  NOR2_X1   g658(.A1(new_n844), .A2(new_n779), .ZN(new_n845));
  NAND2_X1  g659(.A1(new_n845), .A2(new_n747), .ZN(new_n846));
  AOI21_X1  g660(.A(new_n840), .B1(new_n841), .B2(new_n846), .ZN(new_n847));
  OAI21_X1  g661(.A(new_n813), .B1(new_n838), .B2(new_n847), .ZN(new_n848));
  NAND2_X1  g662(.A1(new_n818), .A2(new_n669), .ZN(new_n849));
  OAI21_X1  g663(.A(new_n755), .B1(new_n721), .B2(new_n722), .ZN(new_n850));
  OR2_X1    g664(.A1(new_n829), .A2(new_n832), .ZN(new_n851));
  OAI21_X1  g665(.A(new_n849), .B1(new_n850), .B2(new_n851), .ZN(new_n852));
  NOR2_X1   g666(.A1(new_n824), .A2(new_n829), .ZN(new_n853));
  AND2_X1   g667(.A1(new_n766), .A2(new_n597), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  OR2_X1    g669(.A1(new_n855), .A2(KEYINPUT48), .ZN(new_n856));
  NAND2_X1  g670(.A1(new_n855), .A2(KEYINPUT48), .ZN(new_n857));
  AOI21_X1  g671(.A(new_n852), .B1(new_n856), .B2(new_n857), .ZN(new_n858));
  AND2_X1   g672(.A1(new_n791), .A2(new_n806), .ZN(new_n859));
  NOR2_X1   g673(.A1(new_n791), .A2(new_n810), .ZN(new_n860));
  OAI211_X1 g674(.A(KEYINPUT116), .B(new_n846), .C1(new_n859), .C2(new_n860), .ZN(new_n861));
  NAND2_X1  g675(.A1(new_n861), .A2(new_n839), .ZN(new_n862));
  AOI21_X1  g676(.A(KEYINPUT116), .B1(new_n841), .B2(new_n846), .ZN(new_n863));
  NOR2_X1   g677(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  INV_X1    g678(.A(KEYINPUT115), .ZN(new_n865));
  AOI21_X1  g679(.A(new_n813), .B1(new_n835), .B2(new_n865), .ZN(new_n866));
  OAI21_X1  g680(.A(KEYINPUT115), .B1(new_n830), .B2(new_n834), .ZN(new_n867));
  NAND4_X1  g681(.A1(new_n866), .A2(new_n823), .A3(new_n837), .A4(new_n867), .ZN(new_n868));
  OAI211_X1 g682(.A(new_n848), .B(new_n858), .C1(new_n864), .C2(new_n868), .ZN(new_n869));
  INV_X1    g683(.A(new_n869), .ZN(new_n870));
  NAND4_X1  g684(.A1(new_n816), .A2(new_n329), .A3(new_n707), .A4(new_n709), .ZN(new_n871));
  OAI22_X1  g685(.A1(new_n630), .A2(new_n710), .B1(new_n871), .B2(new_n730), .ZN(new_n872));
  AOI21_X1  g686(.A(new_n872), .B1(new_n720), .B2(new_n727), .ZN(new_n873));
  NAND3_X1  g687(.A1(new_n700), .A2(new_n776), .A3(new_n744), .ZN(new_n874));
  NAND3_X1  g688(.A1(new_n275), .A2(new_n320), .A3(new_n671), .ZN(new_n875));
  AOI21_X1  g689(.A(new_n875), .B1(new_n644), .B2(new_n645), .ZN(new_n876));
  AND2_X1   g690(.A1(new_n876), .A2(new_n753), .ZN(new_n877));
  NAND3_X1  g691(.A1(new_n719), .A2(new_n877), .A3(new_n665), .ZN(new_n878));
  NAND3_X1  g692(.A1(new_n777), .A2(new_n874), .A3(new_n878), .ZN(new_n879));
  NAND3_X1  g693(.A1(new_n271), .A2(new_n276), .A3(new_n321), .ZN(new_n880));
  NAND2_X1  g694(.A1(new_n850), .A2(new_n880), .ZN(new_n881));
  NAND4_X1  g695(.A1(new_n440), .A2(new_n329), .A3(new_n441), .A4(new_n443), .ZN(new_n882));
  NOR3_X1   g696(.A1(new_n882), .A2(new_n632), .A3(new_n635), .ZN(new_n883));
  NAND2_X1  g697(.A1(new_n881), .A2(new_n883), .ZN(new_n884));
  NAND3_X1  g698(.A1(new_n884), .A2(new_n598), .A3(new_n661), .ZN(new_n885));
  NOR2_X1   g699(.A1(new_n879), .A2(new_n885), .ZN(new_n886));
  NAND4_X1  g700(.A1(new_n770), .A2(new_n873), .A3(new_n715), .A4(new_n886), .ZN(new_n887));
  AOI21_X1  g701(.A(new_n320), .B1(new_n271), .B2(new_n276), .ZN(new_n888));
  NAND3_X1  g702(.A1(new_n775), .A2(new_n495), .A3(new_n671), .ZN(new_n889));
  INV_X1    g703(.A(new_n889), .ZN(new_n890));
  NAND4_X1  g704(.A1(new_n669), .A2(new_n691), .A3(new_n888), .A4(new_n890), .ZN(new_n891));
  NAND4_X1  g705(.A1(new_n674), .A2(new_n891), .A3(new_n701), .A4(new_n745), .ZN(new_n892));
  NAND2_X1  g706(.A1(new_n892), .A2(KEYINPUT52), .ZN(new_n893));
  NAND3_X1  g707(.A1(new_n563), .A2(new_n665), .A3(new_n660), .ZN(new_n894));
  NAND2_X1  g708(.A1(new_n623), .A2(new_n629), .ZN(new_n895));
  NOR2_X1   g709(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  NOR2_X1   g710(.A1(new_n756), .A2(new_n743), .ZN(new_n897));
  AOI22_X1  g711(.A1(new_n896), .A2(new_n673), .B1(new_n897), .B2(new_n717), .ZN(new_n898));
  INV_X1    g712(.A(KEYINPUT52), .ZN(new_n899));
  NAND4_X1  g713(.A1(new_n898), .A2(new_n899), .A3(new_n701), .A4(new_n891), .ZN(new_n900));
  NAND2_X1  g714(.A1(new_n893), .A2(new_n900), .ZN(new_n901));
  NAND2_X1  g715(.A1(new_n674), .A2(new_n745), .ZN(new_n902));
  AOI21_X1  g716(.A(KEYINPUT53), .B1(new_n902), .B2(KEYINPUT52), .ZN(new_n903));
  OR3_X1    g717(.A1(new_n887), .A2(new_n901), .A3(new_n903), .ZN(new_n904));
  INV_X1    g718(.A(KEYINPUT53), .ZN(new_n905));
  OAI21_X1  g719(.A(new_n905), .B1(new_n887), .B2(new_n901), .ZN(new_n906));
  NAND2_X1  g720(.A1(new_n904), .A2(new_n906), .ZN(new_n907));
  NAND2_X1  g721(.A1(new_n907), .A2(KEYINPUT54), .ZN(new_n908));
  NAND2_X1  g722(.A1(new_n876), .A2(new_n753), .ZN(new_n909));
  OAI22_X1  g723(.A1(new_n754), .A2(new_n672), .B1(new_n894), .B2(new_n909), .ZN(new_n910));
  NOR3_X1   g724(.A1(new_n767), .A2(new_n756), .A3(new_n743), .ZN(new_n911));
  NOR2_X1   g725(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  AND3_X1   g726(.A1(new_n884), .A2(new_n598), .A3(new_n661), .ZN(new_n913));
  INV_X1    g727(.A(KEYINPUT111), .ZN(new_n914));
  NAND3_X1  g728(.A1(new_n912), .A2(new_n913), .A3(new_n914), .ZN(new_n915));
  OAI21_X1  g729(.A(KEYINPUT111), .B1(new_n879), .B2(new_n885), .ZN(new_n916));
  AOI21_X1  g730(.A(new_n905), .B1(new_n902), .B2(KEYINPUT52), .ZN(new_n917));
  AND3_X1   g731(.A1(new_n915), .A2(new_n916), .A3(new_n917), .ZN(new_n918));
  AND2_X1   g732(.A1(new_n893), .A2(new_n900), .ZN(new_n919));
  NAND2_X1  g733(.A1(new_n769), .A2(KEYINPUT42), .ZN(new_n920));
  INV_X1    g734(.A(new_n757), .ZN(new_n921));
  NAND2_X1  g735(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  AOI22_X1  g736(.A1(new_n631), .A2(new_n714), .B1(new_n731), .B2(new_n740), .ZN(new_n923));
  NAND3_X1  g737(.A1(new_n715), .A2(new_n728), .A3(new_n923), .ZN(new_n924));
  NOR2_X1   g738(.A1(new_n922), .A2(new_n924), .ZN(new_n925));
  NAND3_X1  g739(.A1(new_n918), .A2(new_n919), .A3(new_n925), .ZN(new_n926));
  XNOR2_X1  g740(.A(KEYINPUT112), .B(KEYINPUT54), .ZN(new_n927));
  NAND3_X1  g741(.A1(new_n926), .A2(new_n906), .A3(new_n927), .ZN(new_n928));
  NAND4_X1  g742(.A1(new_n870), .A2(KEYINPUT117), .A3(new_n908), .A4(new_n928), .ZN(new_n929));
  NAND2_X1  g743(.A1(new_n929), .A2(G953), .ZN(new_n930));
  INV_X1    g744(.A(KEYINPUT117), .ZN(new_n931));
  NAND4_X1  g745(.A1(new_n870), .A2(new_n931), .A3(new_n908), .A4(new_n928), .ZN(new_n932));
  NAND2_X1  g746(.A1(new_n932), .A2(new_n323), .ZN(new_n933));
  OR4_X1    g747(.A1(new_n773), .A2(new_n794), .A3(new_n624), .A4(new_n747), .ZN(new_n934));
  NOR2_X1   g748(.A1(new_n934), .A2(KEYINPUT110), .ZN(new_n935));
  XNOR2_X1  g749(.A(new_n845), .B(KEYINPUT49), .ZN(new_n936));
  NAND3_X1  g750(.A1(new_n936), .A2(new_n685), .A3(new_n690), .ZN(new_n937));
  NOR3_X1   g751(.A1(new_n935), .A2(new_n682), .A3(new_n937), .ZN(new_n938));
  NAND2_X1  g752(.A1(new_n934), .A2(KEYINPUT110), .ZN(new_n939));
  NAND2_X1  g753(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  NAND3_X1  g754(.A1(new_n930), .A2(new_n933), .A3(new_n940), .ZN(G75));
  XNOR2_X1  g755(.A(new_n435), .B(new_n436), .ZN(new_n942));
  XNOR2_X1  g756(.A(new_n942), .B(KEYINPUT55), .ZN(new_n943));
  INV_X1    g757(.A(new_n943), .ZN(new_n944));
  NAND2_X1  g758(.A1(new_n926), .A2(new_n906), .ZN(new_n945));
  NAND2_X1  g759(.A1(G210), .A2(G902), .ZN(new_n946));
  INV_X1    g760(.A(new_n946), .ZN(new_n947));
  NAND2_X1  g761(.A1(new_n945), .A2(new_n947), .ZN(new_n948));
  AOI21_X1  g762(.A(KEYINPUT56), .B1(new_n948), .B2(KEYINPUT118), .ZN(new_n949));
  AOI21_X1  g763(.A(new_n946), .B1(new_n926), .B2(new_n906), .ZN(new_n950));
  INV_X1    g764(.A(KEYINPUT118), .ZN(new_n951));
  NAND2_X1  g765(.A1(new_n950), .A2(new_n951), .ZN(new_n952));
  AOI21_X1  g766(.A(new_n944), .B1(new_n949), .B2(new_n952), .ZN(new_n953));
  INV_X1    g767(.A(KEYINPUT56), .ZN(new_n954));
  NAND3_X1  g768(.A1(new_n948), .A2(new_n954), .A3(new_n944), .ZN(new_n955));
  NAND2_X1  g769(.A1(new_n322), .A2(G953), .ZN(new_n956));
  XNOR2_X1  g770(.A(new_n956), .B(KEYINPUT119), .ZN(new_n957));
  NAND2_X1  g771(.A1(new_n955), .A2(new_n957), .ZN(new_n958));
  OAI21_X1  g772(.A(KEYINPUT120), .B1(new_n953), .B2(new_n958), .ZN(new_n959));
  INV_X1    g773(.A(new_n952), .ZN(new_n960));
  OAI21_X1  g774(.A(new_n954), .B1(new_n950), .B2(new_n951), .ZN(new_n961));
  OAI21_X1  g775(.A(new_n943), .B1(new_n960), .B2(new_n961), .ZN(new_n962));
  INV_X1    g776(.A(KEYINPUT120), .ZN(new_n963));
  NAND4_X1  g777(.A1(new_n962), .A2(new_n963), .A3(new_n957), .A4(new_n955), .ZN(new_n964));
  NAND2_X1  g778(.A1(new_n959), .A2(new_n964), .ZN(G51));
  INV_X1    g779(.A(new_n957), .ZN(new_n966));
  XNOR2_X1  g780(.A(new_n945), .B(new_n927), .ZN(new_n967));
  XNOR2_X1  g781(.A(new_n493), .B(KEYINPUT57), .ZN(new_n968));
  OAI21_X1  g782(.A(new_n843), .B1(new_n967), .B2(new_n968), .ZN(new_n969));
  NAND2_X1  g783(.A1(new_n945), .A2(G902), .ZN(new_n970));
  OR2_X1    g784(.A1(new_n970), .A2(new_n786), .ZN(new_n971));
  AOI21_X1  g785(.A(new_n966), .B1(new_n969), .B2(new_n971), .ZN(G54));
  INV_X1    g786(.A(KEYINPUT121), .ZN(new_n973));
  NAND2_X1  g787(.A1(new_n254), .A2(new_n256), .ZN(new_n974));
  NAND2_X1  g788(.A1(KEYINPUT58), .A2(G475), .ZN(new_n975));
  OAI21_X1  g789(.A(new_n974), .B1(new_n970), .B2(new_n975), .ZN(new_n976));
  NAND2_X1  g790(.A1(new_n976), .A2(new_n957), .ZN(new_n977));
  NOR3_X1   g791(.A1(new_n970), .A2(new_n974), .A3(new_n975), .ZN(new_n978));
  OAI21_X1  g792(.A(new_n973), .B1(new_n977), .B2(new_n978), .ZN(new_n979));
  INV_X1    g793(.A(new_n978), .ZN(new_n980));
  NAND4_X1  g794(.A1(new_n980), .A2(KEYINPUT121), .A3(new_n957), .A4(new_n976), .ZN(new_n981));
  NAND2_X1  g795(.A1(new_n979), .A2(new_n981), .ZN(G60));
  AND3_X1   g796(.A1(new_n604), .A2(new_n607), .A3(new_n613), .ZN(new_n983));
  NAND2_X1  g797(.A1(G478), .A2(G902), .ZN(new_n984));
  XNOR2_X1  g798(.A(new_n984), .B(KEYINPUT59), .ZN(new_n985));
  NAND2_X1  g799(.A1(new_n983), .A2(new_n985), .ZN(new_n986));
  OAI21_X1  g800(.A(new_n957), .B1(new_n967), .B2(new_n986), .ZN(new_n987));
  NAND2_X1  g801(.A1(new_n908), .A2(new_n928), .ZN(new_n988));
  AOI21_X1  g802(.A(new_n983), .B1(new_n988), .B2(new_n985), .ZN(new_n989));
  NOR2_X1   g803(.A1(new_n987), .A2(new_n989), .ZN(G63));
  NAND2_X1  g804(.A1(G217), .A2(G902), .ZN(new_n991));
  XOR2_X1   g805(.A(new_n991), .B(KEYINPUT60), .Z(new_n992));
  NAND2_X1  g806(.A1(new_n945), .A2(new_n992), .ZN(new_n993));
  NOR2_X1   g807(.A1(new_n585), .A2(new_n586), .ZN(new_n994));
  AOI21_X1  g808(.A(new_n966), .B1(new_n993), .B2(new_n994), .ZN(new_n995));
  NAND3_X1  g809(.A1(new_n945), .A2(new_n657), .A3(new_n992), .ZN(new_n996));
  NAND2_X1  g810(.A1(new_n995), .A2(new_n996), .ZN(new_n997));
  NAND2_X1  g811(.A1(KEYINPUT122), .A2(KEYINPUT61), .ZN(new_n998));
  INV_X1    g812(.A(KEYINPUT122), .ZN(new_n999));
  INV_X1    g813(.A(KEYINPUT61), .ZN(new_n1000));
  NAND2_X1  g814(.A1(new_n999), .A2(new_n1000), .ZN(new_n1001));
  NAND3_X1  g815(.A1(new_n997), .A2(new_n998), .A3(new_n1001), .ZN(new_n1002));
  NAND4_X1  g816(.A1(new_n995), .A2(new_n999), .A3(new_n1000), .A4(new_n996), .ZN(new_n1003));
  AND2_X1   g817(.A1(new_n1002), .A2(new_n1003), .ZN(G66));
  AOI21_X1  g818(.A(new_n210), .B1(new_n327), .B2(new_n355), .ZN(new_n1005));
  NOR2_X1   g819(.A1(new_n924), .A2(new_n885), .ZN(new_n1006));
  INV_X1    g820(.A(new_n1006), .ZN(new_n1007));
  AOI21_X1  g821(.A(new_n1005), .B1(new_n1007), .B2(new_n210), .ZN(new_n1008));
  OAI211_X1 g822(.A(new_n406), .B(new_n407), .C1(G898), .C2(new_n210), .ZN(new_n1009));
  XOR2_X1   g823(.A(new_n1008), .B(new_n1009), .Z(G69));
  AOI21_X1  g824(.A(new_n210), .B1(G227), .B2(G900), .ZN(new_n1011));
  INV_X1    g825(.A(new_n1011), .ZN(new_n1012));
  INV_X1    g826(.A(KEYINPUT124), .ZN(new_n1013));
  NOR2_X1   g827(.A1(new_n221), .A2(new_n222), .ZN(new_n1014));
  XNOR2_X1  g828(.A(new_n545), .B(new_n1014), .ZN(new_n1015));
  INV_X1    g829(.A(KEYINPUT99), .ZN(new_n1016));
  OR2_X1    g830(.A1(new_n696), .A2(new_n1016), .ZN(new_n1017));
  NAND2_X1  g831(.A1(new_n696), .A2(new_n1016), .ZN(new_n1018));
  AND3_X1   g832(.A1(new_n674), .A2(new_n701), .A3(new_n745), .ZN(new_n1019));
  NAND3_X1  g833(.A1(new_n1017), .A2(new_n1018), .A3(new_n1019), .ZN(new_n1020));
  NAND2_X1  g834(.A1(new_n1020), .A2(KEYINPUT62), .ZN(new_n1021));
  NOR2_X1   g835(.A1(new_n808), .A2(new_n693), .ZN(new_n1022));
  AND3_X1   g836(.A1(new_n1022), .A2(new_n881), .A3(new_n774), .ZN(new_n1023));
  AOI21_X1  g837(.A(new_n1023), .B1(new_n792), .B2(new_n802), .ZN(new_n1024));
  NAND3_X1  g838(.A1(new_n1021), .A2(new_n811), .A3(new_n1024), .ZN(new_n1025));
  INV_X1    g839(.A(KEYINPUT123), .ZN(new_n1026));
  OAI21_X1  g840(.A(new_n1026), .B1(new_n1020), .B2(KEYINPUT62), .ZN(new_n1027));
  INV_X1    g841(.A(KEYINPUT62), .ZN(new_n1028));
  NAND4_X1  g842(.A1(new_n697), .A2(KEYINPUT123), .A3(new_n1028), .A4(new_n1019), .ZN(new_n1029));
  AOI21_X1  g843(.A(new_n1025), .B1(new_n1027), .B2(new_n1029), .ZN(new_n1030));
  OAI21_X1  g844(.A(new_n1015), .B1(new_n1030), .B2(G953), .ZN(new_n1031));
  AOI21_X1  g845(.A(new_n1015), .B1(G900), .B2(G953), .ZN(new_n1032));
  NAND2_X1  g846(.A1(new_n1019), .A2(new_n777), .ZN(new_n1033));
  AND2_X1   g847(.A1(new_n854), .A2(new_n731), .ZN(new_n1034));
  AOI21_X1  g848(.A(new_n1033), .B1(new_n1034), .B2(new_n792), .ZN(new_n1035));
  NAND4_X1  g849(.A1(new_n1035), .A2(new_n770), .A3(new_n803), .A4(new_n811), .ZN(new_n1036));
  OAI21_X1  g850(.A(new_n1032), .B1(new_n1036), .B2(G953), .ZN(new_n1037));
  AOI21_X1  g851(.A(new_n1013), .B1(new_n1031), .B2(new_n1037), .ZN(new_n1038));
  AND3_X1   g852(.A1(new_n1021), .A2(new_n811), .A3(new_n1024), .ZN(new_n1039));
  NAND2_X1  g853(.A1(new_n1027), .A2(new_n1029), .ZN(new_n1040));
  AOI21_X1  g854(.A(G953), .B1(new_n1039), .B2(new_n1040), .ZN(new_n1041));
  INV_X1    g855(.A(new_n1015), .ZN(new_n1042));
  OAI211_X1 g856(.A(new_n1013), .B(new_n1037), .C1(new_n1041), .C2(new_n1042), .ZN(new_n1043));
  INV_X1    g857(.A(new_n1043), .ZN(new_n1044));
  OAI21_X1  g858(.A(new_n1012), .B1(new_n1038), .B2(new_n1044), .ZN(new_n1045));
  OAI21_X1  g859(.A(new_n1037), .B1(new_n1041), .B2(new_n1042), .ZN(new_n1046));
  NAND2_X1  g860(.A1(new_n1046), .A2(KEYINPUT124), .ZN(new_n1047));
  NAND3_X1  g861(.A1(new_n1047), .A2(new_n1011), .A3(new_n1043), .ZN(new_n1048));
  NAND2_X1  g862(.A1(new_n1045), .A2(new_n1048), .ZN(G72));
  XNOR2_X1  g863(.A(new_n688), .B(KEYINPUT63), .ZN(new_n1050));
  INV_X1    g864(.A(new_n1050), .ZN(new_n1051));
  NOR2_X1   g865(.A1(new_n546), .A2(new_n503), .ZN(new_n1052));
  INV_X1    g866(.A(new_n535), .ZN(new_n1053));
  OAI21_X1  g867(.A(new_n1051), .B1(new_n1052), .B2(new_n1053), .ZN(new_n1054));
  AOI21_X1  g868(.A(new_n1054), .B1(new_n904), .B2(new_n906), .ZN(new_n1055));
  XOR2_X1   g869(.A(new_n1055), .B(KEYINPUT127), .Z(new_n1056));
  OAI21_X1  g870(.A(new_n1051), .B1(new_n1036), .B2(new_n1007), .ZN(new_n1057));
  XNOR2_X1  g871(.A(new_n546), .B(KEYINPUT125), .ZN(new_n1058));
  NOR2_X1   g872(.A1(new_n1058), .A2(new_n503), .ZN(new_n1059));
  XNOR2_X1  g873(.A(new_n1059), .B(KEYINPUT126), .ZN(new_n1060));
  AOI21_X1  g874(.A(new_n966), .B1(new_n1057), .B2(new_n1060), .ZN(new_n1061));
  AOI21_X1  g875(.A(new_n1050), .B1(new_n1030), .B2(new_n1006), .ZN(new_n1062));
  NAND2_X1  g876(.A1(new_n1058), .A2(new_n503), .ZN(new_n1063));
  OAI21_X1  g877(.A(new_n1061), .B1(new_n1062), .B2(new_n1063), .ZN(new_n1064));
  NOR2_X1   g878(.A1(new_n1056), .A2(new_n1064), .ZN(G57));
endmodule


