//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 0 0 0 1 0 1 1 1 0 1 1 1 1 0 1 0 0 1 1 0 0 0 1 0 1 1 0 0 1 0 1 1 0 1 1 1 0 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 0 1 0 1 1 0 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:25:04 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n595, new_n596, new_n597, new_n598, new_n599, new_n600, new_n601,
    new_n602, new_n603, new_n604, new_n605, new_n607, new_n608, new_n609,
    new_n610, new_n611, new_n612, new_n613, new_n614, new_n615, new_n616,
    new_n617, new_n619, new_n620, new_n621, new_n622, new_n623, new_n624,
    new_n625, new_n626, new_n627, new_n628, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n650, new_n651, new_n652, new_n653, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n674, new_n676, new_n677, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n691, new_n692, new_n693, new_n694,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n729, new_n730, new_n731,
    new_n732, new_n733, new_n734, new_n735, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n912, new_n913,
    new_n914, new_n915, new_n916, new_n917, new_n918, new_n919, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n966,
    new_n967, new_n968, new_n969, new_n970, new_n971, new_n972, new_n973,
    new_n974, new_n975, new_n976, new_n977, new_n978, new_n979;
  INV_X1    g000(.A(G143), .ZN(new_n187));
  NOR2_X1   g001(.A1(new_n187), .A2(G146), .ZN(new_n188));
  INV_X1    g002(.A(new_n188), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n187), .A2(KEYINPUT64), .ZN(new_n190));
  INV_X1    g004(.A(KEYINPUT64), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n191), .A2(G143), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n190), .A2(new_n192), .ZN(new_n193));
  INV_X1    g007(.A(G146), .ZN(new_n194));
  OAI21_X1  g008(.A(new_n189), .B1(new_n193), .B2(new_n194), .ZN(new_n195));
  INV_X1    g009(.A(KEYINPUT1), .ZN(new_n196));
  AOI21_X1  g010(.A(new_n196), .B1(new_n193), .B2(new_n194), .ZN(new_n197));
  INV_X1    g011(.A(G128), .ZN(new_n198));
  OAI21_X1  g012(.A(new_n195), .B1(new_n197), .B2(new_n198), .ZN(new_n199));
  INV_X1    g013(.A(KEYINPUT76), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n199), .A2(new_n200), .ZN(new_n201));
  XNOR2_X1  g015(.A(KEYINPUT68), .B(KEYINPUT1), .ZN(new_n202));
  AND2_X1   g016(.A1(new_n202), .A2(G128), .ZN(new_n203));
  XNOR2_X1  g017(.A(KEYINPUT64), .B(G143), .ZN(new_n204));
  AOI21_X1  g018(.A(new_n188), .B1(new_n204), .B2(G146), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n203), .A2(new_n205), .ZN(new_n206));
  OAI211_X1 g020(.A(KEYINPUT76), .B(new_n195), .C1(new_n197), .C2(new_n198), .ZN(new_n207));
  NAND3_X1  g021(.A1(new_n201), .A2(new_n206), .A3(new_n207), .ZN(new_n208));
  INV_X1    g022(.A(KEYINPUT3), .ZN(new_n209));
  INV_X1    g023(.A(G104), .ZN(new_n210));
  OAI21_X1  g024(.A(new_n209), .B1(new_n210), .B2(G107), .ZN(new_n211));
  INV_X1    g025(.A(G107), .ZN(new_n212));
  NAND3_X1  g026(.A1(new_n212), .A2(KEYINPUT3), .A3(G104), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n211), .A2(new_n213), .ZN(new_n214));
  NOR2_X1   g028(.A1(new_n212), .A2(G104), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n215), .A2(KEYINPUT75), .ZN(new_n216));
  INV_X1    g030(.A(G101), .ZN(new_n217));
  INV_X1    g031(.A(KEYINPUT75), .ZN(new_n218));
  OAI21_X1  g032(.A(new_n218), .B1(new_n212), .B2(G104), .ZN(new_n219));
  NAND4_X1  g033(.A1(new_n214), .A2(new_n216), .A3(new_n217), .A4(new_n219), .ZN(new_n220));
  NOR2_X1   g034(.A1(new_n210), .A2(G107), .ZN(new_n221));
  OAI21_X1  g035(.A(G101), .B1(new_n221), .B2(new_n215), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n220), .A2(new_n222), .ZN(new_n223));
  INV_X1    g037(.A(new_n223), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n208), .A2(new_n224), .ZN(new_n225));
  INV_X1    g039(.A(KEYINPUT10), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  INV_X1    g041(.A(G134), .ZN(new_n228));
  OAI21_X1  g042(.A(KEYINPUT11), .B1(new_n228), .B2(G137), .ZN(new_n229));
  INV_X1    g043(.A(KEYINPUT11), .ZN(new_n230));
  INV_X1    g044(.A(G137), .ZN(new_n231));
  NAND3_X1  g045(.A1(new_n230), .A2(new_n231), .A3(G134), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n229), .A2(new_n232), .ZN(new_n233));
  INV_X1    g047(.A(G131), .ZN(new_n234));
  OAI21_X1  g048(.A(KEYINPUT66), .B1(new_n231), .B2(G134), .ZN(new_n235));
  INV_X1    g049(.A(KEYINPUT66), .ZN(new_n236));
  NAND3_X1  g050(.A1(new_n236), .A2(new_n228), .A3(G137), .ZN(new_n237));
  NAND4_X1  g051(.A1(new_n233), .A2(new_n234), .A3(new_n235), .A4(new_n237), .ZN(new_n238));
  INV_X1    g052(.A(new_n238), .ZN(new_n239));
  AND2_X1   g053(.A1(new_n235), .A2(new_n237), .ZN(new_n240));
  AOI21_X1  g054(.A(new_n234), .B1(new_n240), .B2(new_n233), .ZN(new_n241));
  NOR2_X1   g055(.A1(new_n239), .A2(new_n241), .ZN(new_n242));
  NAND3_X1  g056(.A1(new_n214), .A2(new_n219), .A3(new_n216), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n243), .A2(G101), .ZN(new_n244));
  NAND3_X1  g058(.A1(new_n244), .A2(KEYINPUT4), .A3(new_n220), .ZN(new_n245));
  AOI21_X1  g059(.A(KEYINPUT65), .B1(new_n187), .B2(G146), .ZN(new_n246));
  OAI21_X1  g060(.A(new_n246), .B1(new_n204), .B2(G146), .ZN(new_n247));
  NAND3_X1  g061(.A1(new_n193), .A2(KEYINPUT65), .A3(new_n194), .ZN(new_n248));
  XOR2_X1   g062(.A(KEYINPUT0), .B(G128), .Z(new_n249));
  NAND3_X1  g063(.A1(new_n247), .A2(new_n248), .A3(new_n249), .ZN(new_n250));
  NAND3_X1  g064(.A1(new_n205), .A2(KEYINPUT0), .A3(G128), .ZN(new_n251));
  INV_X1    g065(.A(KEYINPUT4), .ZN(new_n252));
  NAND3_X1  g066(.A1(new_n243), .A2(new_n252), .A3(G101), .ZN(new_n253));
  NAND4_X1  g067(.A1(new_n245), .A2(new_n250), .A3(new_n251), .A4(new_n253), .ZN(new_n254));
  OAI21_X1  g068(.A(G128), .B1(new_n202), .B2(new_n188), .ZN(new_n255));
  NAND3_X1  g069(.A1(new_n255), .A2(new_n247), .A3(new_n248), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n256), .A2(new_n206), .ZN(new_n257));
  NAND3_X1  g071(.A1(new_n257), .A2(new_n224), .A3(KEYINPUT10), .ZN(new_n258));
  AND2_X1   g072(.A1(new_n254), .A2(new_n258), .ZN(new_n259));
  NAND3_X1  g073(.A1(new_n227), .A2(new_n242), .A3(new_n259), .ZN(new_n260));
  INV_X1    g074(.A(KEYINPUT77), .ZN(new_n261));
  INV_X1    g075(.A(KEYINPUT12), .ZN(new_n262));
  NOR2_X1   g076(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  NOR2_X1   g077(.A1(new_n257), .A2(new_n224), .ZN(new_n264));
  AOI21_X1  g078(.A(new_n264), .B1(new_n208), .B2(new_n224), .ZN(new_n265));
  AOI21_X1  g079(.A(new_n242), .B1(new_n261), .B2(new_n262), .ZN(new_n266));
  INV_X1    g080(.A(new_n266), .ZN(new_n267));
  OAI21_X1  g081(.A(new_n263), .B1(new_n265), .B2(new_n267), .ZN(new_n268));
  INV_X1    g082(.A(new_n263), .ZN(new_n269));
  AOI22_X1  g083(.A1(new_n199), .A2(new_n200), .B1(new_n205), .B2(new_n203), .ZN(new_n270));
  AOI21_X1  g084(.A(new_n223), .B1(new_n270), .B2(new_n207), .ZN(new_n271));
  OAI211_X1 g085(.A(new_n266), .B(new_n269), .C1(new_n271), .C2(new_n264), .ZN(new_n272));
  NAND3_X1  g086(.A1(new_n260), .A2(new_n268), .A3(new_n272), .ZN(new_n273));
  INV_X1    g087(.A(KEYINPUT78), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  NAND4_X1  g089(.A1(new_n260), .A2(new_n268), .A3(KEYINPUT78), .A4(new_n272), .ZN(new_n276));
  XNOR2_X1  g090(.A(G110), .B(G140), .ZN(new_n277));
  INV_X1    g091(.A(G953), .ZN(new_n278));
  AND2_X1   g092(.A1(new_n278), .A2(G227), .ZN(new_n279));
  XNOR2_X1  g093(.A(new_n277), .B(new_n279), .ZN(new_n280));
  XOR2_X1   g094(.A(new_n280), .B(KEYINPUT74), .Z(new_n281));
  NAND3_X1  g095(.A1(new_n275), .A2(new_n276), .A3(new_n281), .ZN(new_n282));
  INV_X1    g096(.A(KEYINPUT79), .ZN(new_n283));
  INV_X1    g097(.A(new_n242), .ZN(new_n284));
  AOI21_X1  g098(.A(KEYINPUT10), .B1(new_n208), .B2(new_n224), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n254), .A2(new_n258), .ZN(new_n286));
  OAI21_X1  g100(.A(new_n284), .B1(new_n285), .B2(new_n286), .ZN(new_n287));
  NAND3_X1  g101(.A1(new_n260), .A2(new_n283), .A3(new_n287), .ZN(new_n288));
  OAI211_X1 g102(.A(KEYINPUT79), .B(new_n284), .C1(new_n285), .C2(new_n286), .ZN(new_n289));
  AOI21_X1  g103(.A(new_n280), .B1(new_n288), .B2(new_n289), .ZN(new_n290));
  INV_X1    g104(.A(new_n290), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n282), .A2(new_n291), .ZN(new_n292));
  INV_X1    g106(.A(G902), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  INV_X1    g108(.A(KEYINPUT80), .ZN(new_n295));
  NAND3_X1  g109(.A1(new_n294), .A2(new_n295), .A3(G469), .ZN(new_n296));
  XNOR2_X1  g110(.A(KEYINPUT9), .B(G234), .ZN(new_n297));
  OAI21_X1  g111(.A(G221), .B1(new_n297), .B2(G902), .ZN(new_n298));
  AND2_X1   g112(.A1(new_n296), .A2(new_n298), .ZN(new_n299));
  NAND3_X1  g113(.A1(new_n288), .A2(new_n280), .A3(new_n289), .ZN(new_n300));
  INV_X1    g114(.A(new_n280), .ZN(new_n301));
  NAND4_X1  g115(.A1(new_n260), .A2(new_n268), .A3(new_n301), .A4(new_n272), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n300), .A2(new_n302), .ZN(new_n303));
  INV_X1    g117(.A(G469), .ZN(new_n304));
  NAND3_X1  g118(.A1(new_n303), .A2(new_n304), .A3(new_n293), .ZN(new_n305));
  AOI21_X1  g119(.A(G902), .B1(new_n282), .B2(new_n291), .ZN(new_n306));
  OAI211_X1 g120(.A(KEYINPUT80), .B(new_n305), .C1(new_n306), .C2(new_n304), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n299), .A2(new_n307), .ZN(new_n308));
  XNOR2_X1  g122(.A(G113), .B(G122), .ZN(new_n309));
  XNOR2_X1  g123(.A(new_n309), .B(new_n210), .ZN(new_n310));
  INV_X1    g124(.A(new_n310), .ZN(new_n311));
  XNOR2_X1  g125(.A(G125), .B(G140), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n312), .A2(KEYINPUT16), .ZN(new_n313));
  INV_X1    g127(.A(KEYINPUT16), .ZN(new_n314));
  INV_X1    g128(.A(G140), .ZN(new_n315));
  NAND3_X1  g129(.A1(new_n314), .A2(new_n315), .A3(G125), .ZN(new_n316));
  NAND3_X1  g130(.A1(new_n313), .A2(G146), .A3(new_n316), .ZN(new_n317));
  XOR2_X1   g131(.A(new_n312), .B(KEYINPUT19), .Z(new_n318));
  OAI21_X1  g132(.A(new_n317), .B1(new_n318), .B2(G146), .ZN(new_n319));
  INV_X1    g133(.A(G237), .ZN(new_n320));
  NAND4_X1  g134(.A1(new_n320), .A2(new_n278), .A3(G143), .A4(G214), .ZN(new_n321));
  AND3_X1   g135(.A1(new_n320), .A2(new_n278), .A3(G214), .ZN(new_n322));
  OAI21_X1  g136(.A(new_n321), .B1(new_n193), .B2(new_n322), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n323), .A2(G131), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n324), .A2(KEYINPUT86), .ZN(new_n325));
  INV_X1    g139(.A(KEYINPUT86), .ZN(new_n326));
  NAND3_X1  g140(.A1(new_n323), .A2(new_n326), .A3(G131), .ZN(new_n327));
  AND2_X1   g141(.A1(new_n325), .A2(new_n327), .ZN(new_n328));
  OR2_X1    g142(.A1(new_n323), .A2(G131), .ZN(new_n329));
  AOI21_X1  g143(.A(new_n319), .B1(new_n328), .B2(new_n329), .ZN(new_n330));
  NOR2_X1   g144(.A1(new_n323), .A2(KEYINPUT85), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n331), .A2(KEYINPUT84), .ZN(new_n332));
  AND2_X1   g146(.A1(KEYINPUT18), .A2(G131), .ZN(new_n333));
  INV_X1    g147(.A(new_n333), .ZN(new_n334));
  INV_X1    g148(.A(KEYINPUT84), .ZN(new_n335));
  AOI21_X1  g149(.A(new_n334), .B1(new_n323), .B2(new_n335), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n332), .A2(new_n336), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n331), .A2(new_n334), .ZN(new_n338));
  XNOR2_X1  g152(.A(new_n312), .B(new_n194), .ZN(new_n339));
  AND3_X1   g153(.A1(new_n337), .A2(new_n338), .A3(new_n339), .ZN(new_n340));
  OAI21_X1  g154(.A(new_n311), .B1(new_n330), .B2(new_n340), .ZN(new_n341));
  INV_X1    g155(.A(KEYINPUT17), .ZN(new_n342));
  NAND4_X1  g156(.A1(new_n325), .A2(new_n329), .A3(new_n342), .A4(new_n327), .ZN(new_n343));
  INV_X1    g157(.A(new_n317), .ZN(new_n344));
  AOI21_X1  g158(.A(G146), .B1(new_n313), .B2(new_n316), .ZN(new_n345));
  NOR2_X1   g159(.A1(new_n344), .A2(new_n345), .ZN(new_n346));
  OAI211_X1 g160(.A(new_n343), .B(new_n346), .C1(new_n328), .C2(new_n342), .ZN(new_n347));
  NAND3_X1  g161(.A1(new_n337), .A2(new_n338), .A3(new_n339), .ZN(new_n348));
  NAND3_X1  g162(.A1(new_n347), .A2(new_n348), .A3(new_n310), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n341), .A2(new_n349), .ZN(new_n350));
  INV_X1    g164(.A(KEYINPUT20), .ZN(new_n351));
  NOR2_X1   g165(.A1(G475), .A2(G902), .ZN(new_n352));
  AND3_X1   g166(.A1(new_n350), .A2(new_n351), .A3(new_n352), .ZN(new_n353));
  AOI21_X1  g167(.A(new_n351), .B1(new_n350), .B2(new_n352), .ZN(new_n354));
  INV_X1    g168(.A(G475), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n347), .A2(new_n348), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n356), .A2(new_n311), .ZN(new_n357));
  AOI21_X1  g171(.A(G902), .B1(new_n357), .B2(new_n349), .ZN(new_n358));
  OAI22_X1  g172(.A1(new_n353), .A2(new_n354), .B1(new_n355), .B2(new_n358), .ZN(new_n359));
  INV_X1    g173(.A(new_n359), .ZN(new_n360));
  NAND2_X1  g174(.A1(G234), .A2(G237), .ZN(new_n361));
  NAND3_X1  g175(.A1(new_n361), .A2(G952), .A3(new_n278), .ZN(new_n362));
  INV_X1    g176(.A(new_n362), .ZN(new_n363));
  NAND3_X1  g177(.A1(new_n361), .A2(G902), .A3(G953), .ZN(new_n364));
  INV_X1    g178(.A(new_n364), .ZN(new_n365));
  XNOR2_X1  g179(.A(KEYINPUT21), .B(G898), .ZN(new_n366));
  AOI21_X1  g180(.A(new_n363), .B1(new_n365), .B2(new_n366), .ZN(new_n367));
  INV_X1    g181(.A(new_n367), .ZN(new_n368));
  INV_X1    g182(.A(G217), .ZN(new_n369));
  NOR3_X1   g183(.A1(new_n297), .A2(new_n369), .A3(G953), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n198), .A2(G143), .ZN(new_n371));
  OAI21_X1  g185(.A(new_n371), .B1(new_n193), .B2(new_n198), .ZN(new_n372));
  XNOR2_X1  g186(.A(new_n372), .B(G134), .ZN(new_n373));
  INV_X1    g187(.A(G122), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n374), .A2(G116), .ZN(new_n375));
  AOI21_X1  g189(.A(new_n212), .B1(new_n375), .B2(KEYINPUT14), .ZN(new_n376));
  XNOR2_X1  g190(.A(G116), .B(G122), .ZN(new_n377));
  XNOR2_X1  g191(.A(new_n376), .B(new_n377), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n373), .A2(new_n378), .ZN(new_n379));
  INV_X1    g193(.A(KEYINPUT13), .ZN(new_n380));
  NAND3_X1  g194(.A1(new_n204), .A2(new_n380), .A3(G128), .ZN(new_n381));
  OAI211_X1 g195(.A(G134), .B(new_n381), .C1(new_n372), .C2(new_n380), .ZN(new_n382));
  XNOR2_X1  g196(.A(KEYINPUT87), .B(G107), .ZN(new_n383));
  XNOR2_X1  g197(.A(new_n377), .B(new_n383), .ZN(new_n384));
  OAI211_X1 g198(.A(new_n382), .B(new_n384), .C1(G134), .C2(new_n372), .ZN(new_n385));
  AOI21_X1  g199(.A(new_n370), .B1(new_n379), .B2(new_n385), .ZN(new_n386));
  INV_X1    g200(.A(new_n386), .ZN(new_n387));
  NAND3_X1  g201(.A1(new_n379), .A2(new_n385), .A3(new_n370), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n387), .A2(new_n388), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n389), .A2(new_n293), .ZN(new_n390));
  INV_X1    g204(.A(G478), .ZN(new_n391));
  INV_X1    g205(.A(KEYINPUT88), .ZN(new_n392));
  NOR2_X1   g206(.A1(new_n392), .A2(KEYINPUT15), .ZN(new_n393));
  INV_X1    g207(.A(new_n393), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n392), .A2(KEYINPUT15), .ZN(new_n395));
  AOI21_X1  g209(.A(new_n391), .B1(new_n394), .B2(new_n395), .ZN(new_n396));
  OR2_X1    g210(.A1(new_n390), .A2(new_n396), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n390), .A2(new_n396), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n397), .A2(new_n398), .ZN(new_n399));
  INV_X1    g213(.A(new_n399), .ZN(new_n400));
  NAND3_X1  g214(.A1(new_n360), .A2(new_n368), .A3(new_n400), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n250), .A2(new_n251), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n402), .A2(G125), .ZN(new_n403));
  OAI21_X1  g217(.A(new_n403), .B1(G125), .B2(new_n257), .ZN(new_n404));
  NAND3_X1  g218(.A1(new_n404), .A2(G224), .A3(new_n278), .ZN(new_n405));
  XNOR2_X1  g219(.A(G110), .B(G122), .ZN(new_n406));
  XNOR2_X1  g220(.A(new_n406), .B(KEYINPUT8), .ZN(new_n407));
  INV_X1    g221(.A(KEYINPUT5), .ZN(new_n408));
  INV_X1    g222(.A(G119), .ZN(new_n409));
  NAND3_X1  g223(.A1(new_n408), .A2(new_n409), .A3(G116), .ZN(new_n410));
  INV_X1    g224(.A(KEYINPUT82), .ZN(new_n411));
  XNOR2_X1  g225(.A(new_n410), .B(new_n411), .ZN(new_n412));
  XOR2_X1   g226(.A(G116), .B(G119), .Z(new_n413));
  OAI211_X1 g227(.A(new_n412), .B(G113), .C1(new_n408), .C2(new_n413), .ZN(new_n414));
  XNOR2_X1  g228(.A(KEYINPUT2), .B(G113), .ZN(new_n415));
  OR2_X1    g229(.A1(new_n413), .A2(new_n415), .ZN(new_n416));
  NAND3_X1  g230(.A1(new_n224), .A2(new_n414), .A3(new_n416), .ZN(new_n417));
  INV_X1    g231(.A(new_n417), .ZN(new_n418));
  AOI21_X1  g232(.A(new_n224), .B1(new_n414), .B2(new_n416), .ZN(new_n419));
  OAI21_X1  g233(.A(new_n407), .B1(new_n418), .B2(new_n419), .ZN(new_n420));
  INV_X1    g234(.A(KEYINPUT7), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n404), .A2(new_n421), .ZN(new_n422));
  AND3_X1   g236(.A1(new_n405), .A2(new_n420), .A3(new_n422), .ZN(new_n423));
  OR2_X1    g237(.A1(new_n257), .A2(G125), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n278), .A2(G224), .ZN(new_n425));
  NAND4_X1  g239(.A1(new_n424), .A2(KEYINPUT7), .A3(new_n425), .A4(new_n403), .ZN(new_n426));
  XNOR2_X1  g240(.A(new_n413), .B(new_n415), .ZN(new_n427));
  NAND3_X1  g241(.A1(new_n245), .A2(new_n427), .A3(new_n253), .ZN(new_n428));
  NAND3_X1  g242(.A1(new_n428), .A2(new_n417), .A3(new_n406), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n426), .A2(new_n429), .ZN(new_n430));
  INV_X1    g244(.A(new_n430), .ZN(new_n431));
  AOI21_X1  g245(.A(G902), .B1(new_n423), .B2(new_n431), .ZN(new_n432));
  OAI21_X1  g246(.A(G210), .B1(G237), .B2(G902), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n428), .A2(new_n417), .ZN(new_n434));
  INV_X1    g248(.A(new_n406), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  NAND3_X1  g250(.A1(new_n436), .A2(KEYINPUT6), .A3(new_n429), .ZN(new_n437));
  NAND3_X1  g251(.A1(new_n424), .A2(new_n425), .A3(new_n403), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n405), .A2(new_n438), .ZN(new_n439));
  INV_X1    g253(.A(KEYINPUT6), .ZN(new_n440));
  NAND3_X1  g254(.A1(new_n434), .A2(new_n440), .A3(new_n435), .ZN(new_n441));
  NAND3_X1  g255(.A1(new_n437), .A2(new_n439), .A3(new_n441), .ZN(new_n442));
  NAND3_X1  g256(.A1(new_n432), .A2(new_n433), .A3(new_n442), .ZN(new_n443));
  OR2_X1    g257(.A1(new_n443), .A2(KEYINPUT83), .ZN(new_n444));
  INV_X1    g258(.A(new_n433), .ZN(new_n445));
  INV_X1    g259(.A(new_n442), .ZN(new_n446));
  NAND3_X1  g260(.A1(new_n405), .A2(new_n420), .A3(new_n422), .ZN(new_n447));
  OAI21_X1  g261(.A(new_n293), .B1(new_n447), .B2(new_n430), .ZN(new_n448));
  OAI21_X1  g262(.A(new_n445), .B1(new_n446), .B2(new_n448), .ZN(new_n449));
  NAND3_X1  g263(.A1(new_n449), .A2(new_n443), .A3(KEYINPUT83), .ZN(new_n450));
  OAI21_X1  g264(.A(G214), .B1(G237), .B2(G902), .ZN(new_n451));
  XOR2_X1   g265(.A(new_n451), .B(KEYINPUT81), .Z(new_n452));
  NAND3_X1  g266(.A1(new_n444), .A2(new_n450), .A3(new_n452), .ZN(new_n453));
  NOR3_X1   g267(.A1(new_n308), .A2(new_n401), .A3(new_n453), .ZN(new_n454));
  AOI21_X1  g268(.A(new_n369), .B1(G234), .B2(new_n293), .ZN(new_n455));
  XNOR2_X1  g269(.A(KEYINPUT22), .B(G137), .ZN(new_n456));
  AND3_X1   g270(.A1(new_n278), .A2(G221), .A3(G234), .ZN(new_n457));
  XOR2_X1   g271(.A(new_n456), .B(new_n457), .Z(new_n458));
  INV_X1    g272(.A(new_n346), .ZN(new_n459));
  INV_X1    g273(.A(KEYINPUT23), .ZN(new_n460));
  OAI21_X1  g274(.A(new_n460), .B1(new_n409), .B2(G128), .ZN(new_n461));
  NAND3_X1  g275(.A1(new_n198), .A2(KEYINPUT23), .A3(G119), .ZN(new_n462));
  OAI211_X1 g276(.A(new_n461), .B(new_n462), .C1(G119), .C2(new_n198), .ZN(new_n463));
  XNOR2_X1  g277(.A(G119), .B(G128), .ZN(new_n464));
  XOR2_X1   g278(.A(KEYINPUT24), .B(G110), .Z(new_n465));
  AOI22_X1  g279(.A1(new_n463), .A2(G110), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n459), .A2(new_n466), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n467), .A2(KEYINPUT73), .ZN(new_n468));
  INV_X1    g282(.A(KEYINPUT73), .ZN(new_n469));
  NAND3_X1  g283(.A1(new_n459), .A2(new_n469), .A3(new_n466), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n468), .A2(new_n470), .ZN(new_n471));
  OAI22_X1  g285(.A1(new_n463), .A2(G110), .B1(new_n464), .B2(new_n465), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n312), .A2(new_n194), .ZN(new_n473));
  AND3_X1   g287(.A1(new_n472), .A2(new_n317), .A3(new_n473), .ZN(new_n474));
  INV_X1    g288(.A(new_n474), .ZN(new_n475));
  AOI21_X1  g289(.A(new_n458), .B1(new_n471), .B2(new_n475), .ZN(new_n476));
  INV_X1    g290(.A(new_n458), .ZN(new_n477));
  AOI211_X1 g291(.A(new_n474), .B(new_n477), .C1(new_n468), .C2(new_n470), .ZN(new_n478));
  NOR2_X1   g292(.A1(new_n476), .A2(new_n478), .ZN(new_n479));
  AOI21_X1  g293(.A(KEYINPUT25), .B1(new_n479), .B2(new_n293), .ZN(new_n480));
  INV_X1    g294(.A(KEYINPUT25), .ZN(new_n481));
  NOR4_X1   g295(.A1(new_n476), .A2(new_n478), .A3(new_n481), .A4(G902), .ZN(new_n482));
  OAI21_X1  g296(.A(new_n455), .B1(new_n480), .B2(new_n482), .ZN(new_n483));
  NOR2_X1   g297(.A1(new_n455), .A2(G902), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n479), .A2(new_n484), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n483), .A2(new_n485), .ZN(new_n486));
  NOR2_X1   g300(.A1(G472), .A2(G902), .ZN(new_n487));
  OAI21_X1  g301(.A(KEYINPUT67), .B1(new_n231), .B2(G134), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n231), .A2(G134), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  NOR3_X1   g304(.A1(new_n231), .A2(KEYINPUT67), .A3(G134), .ZN(new_n491));
  OAI21_X1  g305(.A(G131), .B1(new_n490), .B2(new_n491), .ZN(new_n492));
  AND2_X1   g306(.A1(new_n238), .A2(new_n492), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n257), .A2(new_n493), .ZN(new_n494));
  OAI211_X1 g308(.A(new_n250), .B(new_n251), .C1(new_n239), .C2(new_n241), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  NOR2_X1   g310(.A1(new_n496), .A2(new_n427), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n496), .A2(KEYINPUT30), .ZN(new_n498));
  INV_X1    g312(.A(KEYINPUT30), .ZN(new_n499));
  NAND3_X1  g313(.A1(new_n494), .A2(new_n495), .A3(new_n499), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n498), .A2(new_n500), .ZN(new_n501));
  AOI21_X1  g315(.A(new_n497), .B1(new_n501), .B2(new_n427), .ZN(new_n502));
  NAND3_X1  g316(.A1(new_n320), .A2(new_n278), .A3(G210), .ZN(new_n503));
  XNOR2_X1  g317(.A(new_n503), .B(KEYINPUT27), .ZN(new_n504));
  XNOR2_X1  g318(.A(KEYINPUT26), .B(G101), .ZN(new_n505));
  XNOR2_X1  g319(.A(new_n504), .B(new_n505), .ZN(new_n506));
  AOI21_X1  g320(.A(KEYINPUT31), .B1(new_n502), .B2(new_n506), .ZN(new_n507));
  AND3_X1   g321(.A1(new_n494), .A2(new_n499), .A3(new_n495), .ZN(new_n508));
  AOI21_X1  g322(.A(new_n499), .B1(new_n494), .B2(new_n495), .ZN(new_n509));
  OAI21_X1  g323(.A(new_n427), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  INV_X1    g324(.A(new_n496), .ZN(new_n511));
  INV_X1    g325(.A(new_n427), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  NAND3_X1  g327(.A1(new_n510), .A2(new_n513), .A3(new_n506), .ZN(new_n514));
  INV_X1    g328(.A(KEYINPUT69), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  NAND4_X1  g330(.A1(new_n510), .A2(KEYINPUT69), .A3(new_n513), .A4(new_n506), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  AOI21_X1  g332(.A(new_n507), .B1(new_n518), .B2(KEYINPUT31), .ZN(new_n519));
  NOR2_X1   g333(.A1(new_n497), .A2(KEYINPUT28), .ZN(new_n520));
  AOI21_X1  g334(.A(new_n512), .B1(new_n494), .B2(new_n495), .ZN(new_n521));
  INV_X1    g335(.A(new_n521), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n513), .A2(new_n522), .ZN(new_n523));
  AOI21_X1  g337(.A(new_n520), .B1(new_n523), .B2(KEYINPUT28), .ZN(new_n524));
  NOR2_X1   g338(.A1(new_n524), .A2(new_n506), .ZN(new_n525));
  OAI211_X1 g339(.A(KEYINPUT32), .B(new_n487), .C1(new_n519), .C2(new_n525), .ZN(new_n526));
  INV_X1    g340(.A(KEYINPUT71), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  INV_X1    g342(.A(KEYINPUT31), .ZN(new_n529));
  AOI21_X1  g343(.A(new_n529), .B1(new_n516), .B2(new_n517), .ZN(new_n530));
  OAI22_X1  g344(.A1(new_n530), .A2(new_n507), .B1(new_n524), .B2(new_n506), .ZN(new_n531));
  NAND4_X1  g345(.A1(new_n531), .A2(KEYINPUT71), .A3(KEYINPUT32), .A4(new_n487), .ZN(new_n532));
  INV_X1    g346(.A(KEYINPUT32), .ZN(new_n533));
  AOI21_X1  g347(.A(KEYINPUT69), .B1(new_n502), .B2(new_n506), .ZN(new_n534));
  INV_X1    g348(.A(new_n517), .ZN(new_n535));
  OAI21_X1  g349(.A(KEYINPUT31), .B1(new_n534), .B2(new_n535), .ZN(new_n536));
  INV_X1    g350(.A(new_n507), .ZN(new_n537));
  AOI21_X1  g351(.A(new_n525), .B1(new_n536), .B2(new_n537), .ZN(new_n538));
  INV_X1    g352(.A(new_n487), .ZN(new_n539));
  OAI21_X1  g353(.A(new_n533), .B1(new_n538), .B2(new_n539), .ZN(new_n540));
  AOI21_X1  g354(.A(KEYINPUT29), .B1(new_n524), .B2(new_n506), .ZN(new_n541));
  INV_X1    g355(.A(new_n502), .ZN(new_n542));
  INV_X1    g356(.A(new_n506), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  AOI21_X1  g358(.A(G902), .B1(new_n541), .B2(new_n544), .ZN(new_n545));
  OAI21_X1  g359(.A(KEYINPUT28), .B1(new_n497), .B2(new_n521), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n546), .A2(KEYINPUT70), .ZN(new_n547));
  INV_X1    g361(.A(new_n547), .ZN(new_n548));
  OR2_X1    g362(.A1(new_n497), .A2(KEYINPUT28), .ZN(new_n549));
  AOI21_X1  g363(.A(KEYINPUT70), .B1(new_n549), .B2(new_n546), .ZN(new_n550));
  NOR2_X1   g364(.A1(new_n548), .A2(new_n550), .ZN(new_n551));
  NAND3_X1  g365(.A1(new_n551), .A2(KEYINPUT29), .A3(new_n506), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n545), .A2(new_n552), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n553), .A2(G472), .ZN(new_n554));
  NAND4_X1  g368(.A1(new_n528), .A2(new_n532), .A3(new_n540), .A4(new_n554), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n555), .A2(KEYINPUT72), .ZN(new_n556));
  INV_X1    g370(.A(G472), .ZN(new_n557));
  AOI21_X1  g371(.A(new_n557), .B1(new_n545), .B2(new_n552), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n531), .A2(new_n487), .ZN(new_n559));
  AOI21_X1  g373(.A(new_n558), .B1(new_n559), .B2(new_n533), .ZN(new_n560));
  INV_X1    g374(.A(KEYINPUT72), .ZN(new_n561));
  NAND4_X1  g375(.A1(new_n560), .A2(new_n561), .A3(new_n528), .A4(new_n532), .ZN(new_n562));
  AOI21_X1  g376(.A(new_n486), .B1(new_n556), .B2(new_n562), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n454), .A2(new_n563), .ZN(new_n564));
  XNOR2_X1  g378(.A(new_n564), .B(G101), .ZN(G3));
  INV_X1    g379(.A(new_n486), .ZN(new_n566));
  AND4_X1   g380(.A1(new_n566), .A2(new_n307), .A3(new_n296), .A4(new_n298), .ZN(new_n567));
  AOI21_X1  g381(.A(new_n557), .B1(new_n531), .B2(new_n293), .ZN(new_n568));
  INV_X1    g382(.A(new_n568), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n569), .A2(KEYINPUT89), .ZN(new_n570));
  INV_X1    g384(.A(KEYINPUT89), .ZN(new_n571));
  AOI22_X1  g385(.A1(new_n568), .A2(new_n571), .B1(new_n487), .B2(new_n531), .ZN(new_n572));
  NAND3_X1  g386(.A1(new_n567), .A2(new_n570), .A3(new_n572), .ZN(new_n573));
  INV_X1    g387(.A(new_n573), .ZN(new_n574));
  OAI21_X1  g388(.A(KEYINPUT33), .B1(new_n370), .B2(KEYINPUT90), .ZN(new_n575));
  OR2_X1    g389(.A1(new_n389), .A2(new_n575), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n389), .A2(new_n575), .ZN(new_n577));
  AND2_X1   g391(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  NOR2_X1   g392(.A1(new_n578), .A2(new_n391), .ZN(new_n579));
  NOR2_X1   g393(.A1(new_n391), .A2(new_n293), .ZN(new_n580));
  INV_X1    g394(.A(new_n580), .ZN(new_n581));
  OAI21_X1  g395(.A(new_n581), .B1(new_n390), .B2(G478), .ZN(new_n582));
  NOR2_X1   g396(.A1(new_n579), .A2(new_n582), .ZN(new_n583));
  INV_X1    g397(.A(new_n583), .ZN(new_n584));
  NOR2_X1   g398(.A1(new_n584), .A2(new_n360), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n449), .A2(new_n443), .ZN(new_n586));
  INV_X1    g400(.A(new_n586), .ZN(new_n587));
  INV_X1    g401(.A(new_n451), .ZN(new_n588));
  NOR2_X1   g402(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  AND3_X1   g403(.A1(new_n585), .A2(new_n368), .A3(new_n589), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n574), .A2(new_n590), .ZN(new_n591));
  XNOR2_X1  g405(.A(new_n591), .B(new_n210), .ZN(new_n592));
  XNOR2_X1  g406(.A(KEYINPUT91), .B(KEYINPUT34), .ZN(new_n593));
  XNOR2_X1  g407(.A(new_n592), .B(new_n593), .ZN(G6));
  NOR2_X1   g408(.A1(new_n358), .A2(new_n355), .ZN(new_n595));
  INV_X1    g409(.A(KEYINPUT92), .ZN(new_n596));
  OR3_X1    g410(.A1(new_n353), .A2(new_n354), .A3(new_n596), .ZN(new_n597));
  OAI21_X1  g411(.A(new_n596), .B1(new_n353), .B2(new_n354), .ZN(new_n598));
  AOI21_X1  g412(.A(new_n595), .B1(new_n597), .B2(new_n598), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n599), .A2(new_n399), .ZN(new_n600));
  XNOR2_X1  g414(.A(new_n367), .B(KEYINPUT93), .ZN(new_n601));
  INV_X1    g415(.A(new_n601), .ZN(new_n602));
  NOR4_X1   g416(.A1(new_n600), .A2(new_n587), .A3(new_n588), .A4(new_n602), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n574), .A2(new_n603), .ZN(new_n604));
  XOR2_X1   g418(.A(KEYINPUT35), .B(G107), .Z(new_n605));
  XNOR2_X1  g419(.A(new_n604), .B(new_n605), .ZN(G9));
  INV_X1    g420(.A(new_n453), .ZN(new_n607));
  AND4_X1   g421(.A1(new_n607), .A2(new_n296), .A3(new_n307), .A4(new_n298), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n471), .A2(new_n475), .ZN(new_n609));
  NOR2_X1   g423(.A1(new_n477), .A2(KEYINPUT36), .ZN(new_n610));
  XNOR2_X1  g424(.A(new_n609), .B(new_n610), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n611), .A2(new_n484), .ZN(new_n612));
  AND2_X1   g426(.A1(new_n483), .A2(new_n612), .ZN(new_n613));
  NOR2_X1   g427(.A1(new_n613), .A2(new_n401), .ZN(new_n614));
  NAND4_X1  g428(.A1(new_n608), .A2(new_n570), .A3(new_n572), .A4(new_n614), .ZN(new_n615));
  XNOR2_X1  g429(.A(new_n615), .B(KEYINPUT94), .ZN(new_n616));
  XOR2_X1   g430(.A(KEYINPUT37), .B(G110), .Z(new_n617));
  XNOR2_X1  g431(.A(new_n616), .B(new_n617), .ZN(G12));
  NAND2_X1  g432(.A1(new_n556), .A2(new_n562), .ZN(new_n619));
  INV_X1    g433(.A(new_n308), .ZN(new_n620));
  INV_X1    g434(.A(new_n613), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n621), .A2(new_n589), .ZN(new_n622));
  XNOR2_X1  g436(.A(KEYINPUT95), .B(G900), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n365), .A2(new_n623), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n624), .A2(new_n362), .ZN(new_n625));
  INV_X1    g439(.A(new_n625), .ZN(new_n626));
  NOR3_X1   g440(.A1(new_n622), .A2(new_n600), .A3(new_n626), .ZN(new_n627));
  NAND3_X1  g441(.A1(new_n619), .A2(new_n620), .A3(new_n627), .ZN(new_n628));
  XNOR2_X1  g442(.A(new_n628), .B(G128), .ZN(G30));
  XNOR2_X1  g443(.A(new_n625), .B(KEYINPUT39), .ZN(new_n630));
  NAND2_X1  g444(.A1(new_n620), .A2(new_n630), .ZN(new_n631));
  OR2_X1    g445(.A1(new_n631), .A2(KEYINPUT40), .ZN(new_n632));
  AND2_X1   g446(.A1(new_n528), .A2(new_n532), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n523), .A2(new_n543), .ZN(new_n634));
  XNOR2_X1  g448(.A(new_n634), .B(KEYINPUT96), .ZN(new_n635));
  INV_X1    g449(.A(new_n518), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  AOI21_X1  g451(.A(new_n557), .B1(new_n637), .B2(new_n293), .ZN(new_n638));
  AOI21_X1  g452(.A(new_n638), .B1(new_n533), .B2(new_n559), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n633), .A2(new_n639), .ZN(new_n640));
  INV_X1    g454(.A(new_n640), .ZN(new_n641));
  NOR2_X1   g455(.A1(new_n641), .A2(new_n621), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n631), .A2(KEYINPUT40), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n444), .A2(new_n450), .ZN(new_n644));
  XOR2_X1   g458(.A(new_n644), .B(KEYINPUT38), .Z(new_n645));
  AOI21_X1  g459(.A(new_n588), .B1(new_n397), .B2(new_n398), .ZN(new_n646));
  AND3_X1   g460(.A1(new_n645), .A2(new_n359), .A3(new_n646), .ZN(new_n647));
  NAND4_X1  g461(.A1(new_n632), .A2(new_n642), .A3(new_n643), .A4(new_n647), .ZN(new_n648));
  XNOR2_X1  g462(.A(new_n648), .B(new_n193), .ZN(G45));
  NOR3_X1   g463(.A1(new_n584), .A2(new_n360), .A3(new_n626), .ZN(new_n650));
  INV_X1    g464(.A(new_n650), .ZN(new_n651));
  NOR2_X1   g465(.A1(new_n651), .A2(new_n622), .ZN(new_n652));
  NAND3_X1  g466(.A1(new_n619), .A2(new_n620), .A3(new_n652), .ZN(new_n653));
  XNOR2_X1  g467(.A(new_n653), .B(G146), .ZN(G48));
  INV_X1    g468(.A(KEYINPUT98), .ZN(new_n655));
  INV_X1    g469(.A(KEYINPUT97), .ZN(new_n656));
  AOI21_X1  g470(.A(new_n304), .B1(new_n303), .B2(new_n293), .ZN(new_n657));
  AOI211_X1 g471(.A(G469), .B(G902), .C1(new_n300), .C2(new_n302), .ZN(new_n658));
  NOR2_X1   g472(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  AOI21_X1  g473(.A(new_n656), .B1(new_n659), .B2(new_n298), .ZN(new_n660));
  INV_X1    g474(.A(new_n298), .ZN(new_n661));
  NOR4_X1   g475(.A1(new_n657), .A2(new_n658), .A3(KEYINPUT97), .A4(new_n661), .ZN(new_n662));
  OAI21_X1  g476(.A(new_n655), .B1(new_n660), .B2(new_n662), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n303), .A2(new_n293), .ZN(new_n664));
  NAND2_X1  g478(.A1(new_n664), .A2(G469), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n665), .A2(new_n305), .ZN(new_n666));
  OAI21_X1  g480(.A(KEYINPUT97), .B1(new_n666), .B2(new_n661), .ZN(new_n667));
  NAND3_X1  g481(.A1(new_n659), .A2(new_n656), .A3(new_n298), .ZN(new_n668));
  NAND3_X1  g482(.A1(new_n667), .A2(new_n668), .A3(KEYINPUT98), .ZN(new_n669));
  AND2_X1   g483(.A1(new_n663), .A2(new_n669), .ZN(new_n670));
  NAND3_X1  g484(.A1(new_n563), .A2(new_n670), .A3(new_n590), .ZN(new_n671));
  XNOR2_X1  g485(.A(KEYINPUT41), .B(G113), .ZN(new_n672));
  XNOR2_X1  g486(.A(new_n671), .B(new_n672), .ZN(G15));
  NAND3_X1  g487(.A1(new_n563), .A2(new_n670), .A3(new_n603), .ZN(new_n674));
  XNOR2_X1  g488(.A(new_n674), .B(G116), .ZN(G18));
  NAND4_X1  g489(.A1(new_n667), .A2(new_n614), .A3(new_n589), .A4(new_n668), .ZN(new_n676));
  AOI21_X1  g490(.A(new_n676), .B1(new_n556), .B2(new_n562), .ZN(new_n677));
  XNOR2_X1  g491(.A(new_n677), .B(new_n409), .ZN(G21));
  XNOR2_X1  g492(.A(new_n487), .B(KEYINPUT99), .ZN(new_n679));
  INV_X1    g493(.A(new_n679), .ZN(new_n680));
  NAND2_X1  g494(.A1(new_n536), .A2(new_n537), .ZN(new_n681));
  INV_X1    g495(.A(KEYINPUT100), .ZN(new_n682));
  OAI21_X1  g496(.A(new_n682), .B1(new_n548), .B2(new_n550), .ZN(new_n683));
  OAI211_X1 g497(.A(KEYINPUT100), .B(new_n547), .C1(new_n524), .C2(KEYINPUT70), .ZN(new_n684));
  NAND3_X1  g498(.A1(new_n683), .A2(new_n684), .A3(new_n543), .ZN(new_n685));
  AOI21_X1  g499(.A(new_n680), .B1(new_n681), .B2(new_n685), .ZN(new_n686));
  NAND4_X1  g500(.A1(new_n586), .A2(new_n646), .A3(new_n359), .A4(new_n601), .ZN(new_n687));
  NOR4_X1   g501(.A1(new_n568), .A2(new_n686), .A3(new_n486), .A4(new_n687), .ZN(new_n688));
  AND3_X1   g502(.A1(new_n663), .A2(new_n669), .A3(new_n688), .ZN(new_n689));
  XNOR2_X1  g503(.A(new_n689), .B(new_n374), .ZN(G24));
  NOR2_X1   g504(.A1(new_n568), .A2(new_n686), .ZN(new_n691));
  NAND3_X1  g505(.A1(new_n650), .A2(new_n691), .A3(new_n621), .ZN(new_n692));
  NAND3_X1  g506(.A1(new_n667), .A2(new_n668), .A3(new_n589), .ZN(new_n693));
  NOR2_X1   g507(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  XOR2_X1   g508(.A(new_n694), .B(G125), .Z(G27));
  NAND3_X1  g509(.A1(new_n644), .A2(new_n451), .A3(new_n298), .ZN(new_n696));
  INV_X1    g510(.A(KEYINPUT102), .ZN(new_n697));
  AND2_X1   g511(.A1(new_n273), .A2(new_n274), .ZN(new_n698));
  NAND2_X1  g512(.A1(new_n276), .A2(new_n281), .ZN(new_n699));
  OAI21_X1  g513(.A(KEYINPUT101), .B1(new_n698), .B2(new_n699), .ZN(new_n700));
  INV_X1    g514(.A(KEYINPUT101), .ZN(new_n701));
  NAND4_X1  g515(.A1(new_n275), .A2(new_n701), .A3(new_n276), .A4(new_n281), .ZN(new_n702));
  AOI211_X1 g516(.A(new_n304), .B(new_n290), .C1(new_n700), .C2(new_n702), .ZN(new_n703));
  NAND2_X1  g517(.A1(G469), .A2(G902), .ZN(new_n704));
  NAND2_X1  g518(.A1(new_n305), .A2(new_n704), .ZN(new_n705));
  OAI21_X1  g519(.A(new_n697), .B1(new_n703), .B2(new_n705), .ZN(new_n706));
  NAND2_X1  g520(.A1(new_n700), .A2(new_n702), .ZN(new_n707));
  NAND3_X1  g521(.A1(new_n707), .A2(G469), .A3(new_n291), .ZN(new_n708));
  INV_X1    g522(.A(new_n705), .ZN(new_n709));
  NAND3_X1  g523(.A1(new_n708), .A2(new_n709), .A3(KEYINPUT102), .ZN(new_n710));
  AOI21_X1  g524(.A(new_n696), .B1(new_n706), .B2(new_n710), .ZN(new_n711));
  NOR2_X1   g525(.A1(new_n651), .A2(KEYINPUT42), .ZN(new_n712));
  NAND3_X1  g526(.A1(new_n563), .A2(new_n711), .A3(new_n712), .ZN(new_n713));
  INV_X1    g527(.A(new_n696), .ZN(new_n714));
  NOR3_X1   g528(.A1(new_n703), .A2(new_n697), .A3(new_n705), .ZN(new_n715));
  AOI21_X1  g529(.A(KEYINPUT102), .B1(new_n708), .B2(new_n709), .ZN(new_n716));
  OAI211_X1 g530(.A(new_n650), .B(new_n714), .C1(new_n715), .C2(new_n716), .ZN(new_n717));
  INV_X1    g531(.A(KEYINPUT103), .ZN(new_n718));
  NAND3_X1  g532(.A1(new_n540), .A2(new_n718), .A3(new_n526), .ZN(new_n719));
  NAND3_X1  g533(.A1(new_n559), .A2(KEYINPUT103), .A3(new_n533), .ZN(new_n720));
  NAND2_X1  g534(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  AOI21_X1  g535(.A(new_n558), .B1(new_n721), .B2(KEYINPUT104), .ZN(new_n722));
  INV_X1    g536(.A(KEYINPUT104), .ZN(new_n723));
  NAND3_X1  g537(.A1(new_n719), .A2(new_n723), .A3(new_n720), .ZN(new_n724));
  AOI211_X1 g538(.A(new_n486), .B(new_n717), .C1(new_n722), .C2(new_n724), .ZN(new_n725));
  INV_X1    g539(.A(KEYINPUT42), .ZN(new_n726));
  OAI21_X1  g540(.A(new_n713), .B1(new_n725), .B2(new_n726), .ZN(new_n727));
  XNOR2_X1  g541(.A(new_n727), .B(new_n234), .ZN(G33));
  NOR2_X1   g542(.A1(new_n600), .A2(new_n626), .ZN(new_n729));
  NAND4_X1  g543(.A1(new_n619), .A2(new_n566), .A3(new_n729), .A4(new_n711), .ZN(new_n730));
  NAND2_X1  g544(.A1(new_n730), .A2(KEYINPUT105), .ZN(new_n731));
  INV_X1    g545(.A(KEYINPUT105), .ZN(new_n732));
  NAND4_X1  g546(.A1(new_n563), .A2(new_n732), .A3(new_n729), .A4(new_n711), .ZN(new_n733));
  NAND2_X1  g547(.A1(new_n731), .A2(new_n733), .ZN(new_n734));
  XOR2_X1   g548(.A(KEYINPUT106), .B(G134), .Z(new_n735));
  XNOR2_X1  g549(.A(new_n734), .B(new_n735), .ZN(G36));
  NAND3_X1  g550(.A1(new_n707), .A2(KEYINPUT45), .A3(new_n291), .ZN(new_n737));
  INV_X1    g551(.A(KEYINPUT45), .ZN(new_n738));
  AOI21_X1  g552(.A(new_n304), .B1(new_n292), .B2(new_n738), .ZN(new_n739));
  NAND2_X1  g553(.A1(new_n737), .A2(new_n739), .ZN(new_n740));
  AND2_X1   g554(.A1(new_n740), .A2(new_n704), .ZN(new_n741));
  OR2_X1    g555(.A1(new_n741), .A2(KEYINPUT46), .ZN(new_n742));
  NAND2_X1  g556(.A1(new_n741), .A2(KEYINPUT46), .ZN(new_n743));
  NAND3_X1  g557(.A1(new_n742), .A2(new_n305), .A3(new_n743), .ZN(new_n744));
  AND3_X1   g558(.A1(new_n744), .A2(new_n298), .A3(new_n630), .ZN(new_n745));
  NAND2_X1  g559(.A1(new_n644), .A2(new_n451), .ZN(new_n746));
  XOR2_X1   g560(.A(new_n746), .B(KEYINPUT107), .Z(new_n747));
  INV_X1    g561(.A(KEYINPUT44), .ZN(new_n748));
  NAND2_X1  g562(.A1(new_n583), .A2(new_n360), .ZN(new_n749));
  XOR2_X1   g563(.A(new_n749), .B(KEYINPUT43), .Z(new_n750));
  AND2_X1   g564(.A1(new_n750), .A2(new_n621), .ZN(new_n751));
  NAND2_X1  g565(.A1(new_n570), .A2(new_n572), .ZN(new_n752));
  AOI21_X1  g566(.A(new_n748), .B1(new_n751), .B2(new_n752), .ZN(new_n753));
  NAND2_X1  g567(.A1(new_n751), .A2(new_n752), .ZN(new_n754));
  NOR2_X1   g568(.A1(new_n754), .A2(KEYINPUT44), .ZN(new_n755));
  OAI211_X1 g569(.A(new_n745), .B(new_n747), .C1(new_n753), .C2(new_n755), .ZN(new_n756));
  XNOR2_X1  g570(.A(new_n756), .B(G137), .ZN(G39));
  NAND2_X1  g571(.A1(new_n744), .A2(new_n298), .ZN(new_n758));
  INV_X1    g572(.A(KEYINPUT47), .ZN(new_n759));
  NAND2_X1  g573(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  NAND3_X1  g574(.A1(new_n744), .A2(KEYINPUT47), .A3(new_n298), .ZN(new_n761));
  NAND2_X1  g575(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  NOR4_X1   g576(.A1(new_n619), .A2(new_n566), .A3(new_n651), .A4(new_n746), .ZN(new_n763));
  NAND2_X1  g577(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  XNOR2_X1  g578(.A(new_n764), .B(G140), .ZN(G42));
  NOR2_X1   g579(.A1(new_n677), .A2(new_n689), .ZN(new_n766));
  NAND3_X1  g580(.A1(new_n766), .A2(new_n671), .A3(new_n674), .ZN(new_n767));
  NAND2_X1  g581(.A1(new_n767), .A2(KEYINPUT110), .ZN(new_n768));
  INV_X1    g582(.A(KEYINPUT110), .ZN(new_n769));
  NAND4_X1  g583(.A1(new_n766), .A2(new_n671), .A3(new_n674), .A4(new_n769), .ZN(new_n770));
  AND2_X1   g584(.A1(new_n768), .A2(new_n770), .ZN(new_n771));
  INV_X1    g585(.A(new_n694), .ZN(new_n772));
  NAND2_X1  g586(.A1(new_n706), .A2(new_n710), .ZN(new_n773));
  AND3_X1   g587(.A1(new_n586), .A2(new_n359), .A3(new_n646), .ZN(new_n774));
  AND3_X1   g588(.A1(new_n774), .A2(new_n298), .A3(new_n625), .ZN(new_n775));
  NAND4_X1  g589(.A1(new_n640), .A2(new_n613), .A3(new_n773), .A4(new_n775), .ZN(new_n776));
  NAND4_X1  g590(.A1(new_n628), .A2(new_n653), .A3(new_n772), .A4(new_n776), .ZN(new_n777));
  INV_X1    g591(.A(KEYINPUT52), .ZN(new_n778));
  NAND2_X1  g592(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  AOI21_X1  g593(.A(new_n308), .B1(new_n556), .B2(new_n562), .ZN(new_n780));
  AOI21_X1  g594(.A(new_n694), .B1(new_n780), .B2(new_n627), .ZN(new_n781));
  NAND4_X1  g595(.A1(new_n781), .A2(KEYINPUT52), .A3(new_n653), .A4(new_n776), .ZN(new_n782));
  AOI21_X1  g596(.A(new_n727), .B1(new_n779), .B2(new_n782), .ZN(new_n783));
  NAND2_X1  g597(.A1(new_n619), .A2(new_n620), .ZN(new_n784));
  INV_X1    g598(.A(new_n746), .ZN(new_n785));
  NAND4_X1  g599(.A1(new_n785), .A2(new_n400), .A3(new_n599), .A4(new_n625), .ZN(new_n786));
  INV_X1    g600(.A(new_n691), .ZN(new_n787));
  OAI22_X1  g601(.A1(new_n784), .A2(new_n786), .B1(new_n787), .B2(new_n717), .ZN(new_n788));
  AOI22_X1  g602(.A1(new_n621), .A2(new_n788), .B1(new_n731), .B2(new_n733), .ZN(new_n789));
  NAND2_X1  g603(.A1(new_n360), .A2(new_n400), .ZN(new_n790));
  OAI21_X1  g604(.A(new_n790), .B1(new_n360), .B2(new_n583), .ZN(new_n791));
  NOR3_X1   g605(.A1(new_n791), .A2(new_n453), .A3(new_n602), .ZN(new_n792));
  NAND4_X1  g606(.A1(new_n567), .A2(new_n792), .A3(new_n570), .A4(new_n572), .ZN(new_n793));
  NAND3_X1  g607(.A1(new_n564), .A2(new_n615), .A3(new_n793), .ZN(new_n794));
  INV_X1    g608(.A(KEYINPUT53), .ZN(new_n795));
  NOR2_X1   g609(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  NAND4_X1  g610(.A1(new_n771), .A2(new_n783), .A3(new_n789), .A4(new_n796), .ZN(new_n797));
  NAND2_X1  g611(.A1(new_n779), .A2(new_n782), .ZN(new_n798));
  AOI21_X1  g612(.A(new_n486), .B1(new_n722), .B2(new_n724), .ZN(new_n799));
  NAND3_X1  g613(.A1(new_n799), .A2(new_n650), .A3(new_n711), .ZN(new_n800));
  AND2_X1   g614(.A1(new_n563), .A2(new_n711), .ZN(new_n801));
  AOI22_X1  g615(.A1(new_n800), .A2(KEYINPUT42), .B1(new_n801), .B2(new_n712), .ZN(new_n802));
  NOR2_X1   g616(.A1(new_n767), .A2(new_n794), .ZN(new_n803));
  NAND4_X1  g617(.A1(new_n798), .A2(new_n802), .A3(new_n789), .A4(new_n803), .ZN(new_n804));
  NAND2_X1  g618(.A1(new_n804), .A2(new_n795), .ZN(new_n805));
  INV_X1    g619(.A(KEYINPUT54), .ZN(new_n806));
  NAND3_X1  g620(.A1(new_n797), .A2(new_n805), .A3(new_n806), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n788), .A2(new_n621), .ZN(new_n808));
  NAND2_X1  g622(.A1(new_n808), .A2(new_n734), .ZN(new_n809));
  NAND2_X1  g623(.A1(new_n615), .A2(new_n793), .ZN(new_n810));
  AOI21_X1  g624(.A(new_n810), .B1(new_n563), .B2(new_n454), .ZN(new_n811));
  NAND4_X1  g625(.A1(new_n811), .A2(new_n671), .A3(new_n674), .A4(new_n766), .ZN(new_n812));
  NOR2_X1   g626(.A1(new_n809), .A2(new_n812), .ZN(new_n813));
  NAND3_X1  g627(.A1(new_n813), .A2(new_n783), .A3(KEYINPUT53), .ZN(new_n814));
  AOI21_X1  g628(.A(new_n806), .B1(new_n805), .B2(new_n814), .ZN(new_n815));
  INV_X1    g629(.A(KEYINPUT109), .ZN(new_n816));
  OAI21_X1  g630(.A(new_n807), .B1(new_n815), .B2(new_n816), .ZN(new_n817));
  AOI211_X1 g631(.A(KEYINPUT109), .B(new_n806), .C1(new_n805), .C2(new_n814), .ZN(new_n818));
  OAI21_X1  g632(.A(KEYINPUT111), .B1(new_n817), .B2(new_n818), .ZN(new_n819));
  NAND3_X1  g633(.A1(new_n667), .A2(new_n785), .A3(new_n668), .ZN(new_n820));
  NOR4_X1   g634(.A1(new_n640), .A2(new_n820), .A3(new_n486), .A4(new_n362), .ZN(new_n821));
  NAND3_X1  g635(.A1(new_n821), .A2(new_n360), .A3(new_n584), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n750), .A2(new_n363), .ZN(new_n823));
  NOR2_X1   g637(.A1(new_n823), .A2(new_n820), .ZN(new_n824));
  NAND3_X1  g638(.A1(new_n824), .A2(new_n621), .A3(new_n691), .ZN(new_n825));
  NAND2_X1  g639(.A1(new_n822), .A2(new_n825), .ZN(new_n826));
  NOR2_X1   g640(.A1(new_n645), .A2(new_n451), .ZN(new_n827));
  NAND3_X1  g641(.A1(new_n827), .A2(new_n668), .A3(new_n667), .ZN(new_n828));
  OR2_X1    g642(.A1(new_n828), .A2(KEYINPUT113), .ZN(new_n829));
  NOR3_X1   g643(.A1(new_n823), .A2(new_n486), .A3(new_n787), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n828), .A2(KEYINPUT113), .ZN(new_n831));
  NAND3_X1  g645(.A1(new_n829), .A2(new_n830), .A3(new_n831), .ZN(new_n832));
  INV_X1    g646(.A(KEYINPUT50), .ZN(new_n833));
  NAND2_X1  g647(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  NAND4_X1  g648(.A1(new_n829), .A2(KEYINPUT50), .A3(new_n830), .A4(new_n831), .ZN(new_n835));
  AOI21_X1  g649(.A(new_n826), .B1(new_n834), .B2(new_n835), .ZN(new_n836));
  XNOR2_X1  g650(.A(new_n666), .B(KEYINPUT108), .ZN(new_n837));
  NAND2_X1  g651(.A1(new_n837), .A2(new_n661), .ZN(new_n838));
  NAND3_X1  g652(.A1(new_n760), .A2(new_n761), .A3(new_n838), .ZN(new_n839));
  INV_X1    g653(.A(KEYINPUT114), .ZN(new_n840));
  AND2_X1   g654(.A1(new_n839), .A2(new_n840), .ZN(new_n841));
  AND2_X1   g655(.A1(new_n830), .A2(new_n747), .ZN(new_n842));
  OAI21_X1  g656(.A(new_n842), .B1(new_n839), .B2(new_n840), .ZN(new_n843));
  OAI211_X1 g657(.A(new_n836), .B(KEYINPUT51), .C1(new_n841), .C2(new_n843), .ZN(new_n844));
  NAND2_X1  g658(.A1(new_n799), .A2(new_n824), .ZN(new_n845));
  XNOR2_X1  g659(.A(new_n845), .B(KEYINPUT48), .ZN(new_n846));
  NAND2_X1  g660(.A1(new_n821), .A2(new_n585), .ZN(new_n847));
  INV_X1    g661(.A(G952), .ZN(new_n848));
  INV_X1    g662(.A(new_n693), .ZN(new_n849));
  AOI211_X1 g663(.A(new_n848), .B(G953), .C1(new_n830), .C2(new_n849), .ZN(new_n850));
  NAND3_X1  g664(.A1(new_n846), .A2(new_n847), .A3(new_n850), .ZN(new_n851));
  INV_X1    g665(.A(KEYINPUT115), .ZN(new_n852));
  AND2_X1   g666(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  NOR2_X1   g667(.A1(new_n851), .A2(new_n852), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n839), .A2(new_n842), .ZN(new_n855));
  AND2_X1   g669(.A1(new_n836), .A2(new_n855), .ZN(new_n856));
  XOR2_X1   g670(.A(KEYINPUT112), .B(KEYINPUT51), .Z(new_n857));
  OAI221_X1 g671(.A(new_n844), .B1(new_n853), .B2(new_n854), .C1(new_n856), .C2(new_n857), .ZN(new_n858));
  INV_X1    g672(.A(new_n858), .ZN(new_n859));
  NOR2_X1   g673(.A1(new_n804), .A2(new_n795), .ZN(new_n860));
  AOI21_X1  g674(.A(KEYINPUT53), .B1(new_n813), .B2(new_n783), .ZN(new_n861));
  OAI21_X1  g675(.A(KEYINPUT54), .B1(new_n860), .B2(new_n861), .ZN(new_n862));
  NAND2_X1  g676(.A1(new_n862), .A2(KEYINPUT109), .ZN(new_n863));
  NAND2_X1  g677(.A1(new_n815), .A2(new_n816), .ZN(new_n864));
  INV_X1    g678(.A(KEYINPUT111), .ZN(new_n865));
  NAND4_X1  g679(.A1(new_n863), .A2(new_n864), .A3(new_n865), .A4(new_n807), .ZN(new_n866));
  NAND3_X1  g680(.A1(new_n819), .A2(new_n859), .A3(new_n866), .ZN(new_n867));
  NAND2_X1  g681(.A1(new_n848), .A2(new_n278), .ZN(new_n868));
  NAND2_X1  g682(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  XNOR2_X1  g683(.A(new_n837), .B(KEYINPUT49), .ZN(new_n870));
  NAND3_X1  g684(.A1(new_n566), .A2(new_n452), .A3(new_n298), .ZN(new_n871));
  NOR3_X1   g685(.A1(new_n645), .A2(new_n749), .A3(new_n871), .ZN(new_n872));
  NAND3_X1  g686(.A1(new_n870), .A2(new_n872), .A3(new_n641), .ZN(new_n873));
  NAND2_X1  g687(.A1(new_n869), .A2(new_n873), .ZN(G75));
  NOR2_X1   g688(.A1(new_n278), .A2(G952), .ZN(new_n875));
  INV_X1    g689(.A(new_n875), .ZN(new_n876));
  AND4_X1   g690(.A1(new_n789), .A2(new_n768), .A3(new_n796), .A4(new_n770), .ZN(new_n877));
  AOI22_X1  g691(.A1(new_n783), .A2(new_n877), .B1(new_n804), .B2(new_n795), .ZN(new_n878));
  NOR2_X1   g692(.A1(new_n878), .A2(new_n293), .ZN(new_n879));
  AOI21_X1  g693(.A(KEYINPUT56), .B1(new_n879), .B2(G210), .ZN(new_n880));
  NAND2_X1  g694(.A1(new_n437), .A2(new_n441), .ZN(new_n881));
  XNOR2_X1  g695(.A(new_n881), .B(KEYINPUT116), .ZN(new_n882));
  XNOR2_X1  g696(.A(new_n439), .B(KEYINPUT55), .ZN(new_n883));
  XOR2_X1   g697(.A(new_n882), .B(new_n883), .Z(new_n884));
  INV_X1    g698(.A(new_n884), .ZN(new_n885));
  OAI21_X1  g699(.A(new_n876), .B1(new_n880), .B2(new_n885), .ZN(new_n886));
  AOI21_X1  g700(.A(new_n886), .B1(new_n880), .B2(new_n885), .ZN(G51));
  NOR3_X1   g701(.A1(new_n878), .A2(new_n293), .A3(new_n740), .ZN(new_n888));
  XOR2_X1   g702(.A(new_n704), .B(KEYINPUT57), .Z(new_n889));
  INV_X1    g703(.A(new_n807), .ZN(new_n890));
  AOI21_X1  g704(.A(new_n806), .B1(new_n797), .B2(new_n805), .ZN(new_n891));
  OAI21_X1  g705(.A(new_n889), .B1(new_n890), .B2(new_n891), .ZN(new_n892));
  AOI21_X1  g706(.A(new_n888), .B1(new_n892), .B2(new_n303), .ZN(new_n893));
  OAI21_X1  g707(.A(KEYINPUT117), .B1(new_n893), .B2(new_n875), .ZN(new_n894));
  INV_X1    g708(.A(KEYINPUT117), .ZN(new_n895));
  NAND2_X1  g709(.A1(new_n797), .A2(new_n805), .ZN(new_n896));
  NAND2_X1  g710(.A1(new_n896), .A2(KEYINPUT54), .ZN(new_n897));
  NAND2_X1  g711(.A1(new_n897), .A2(new_n807), .ZN(new_n898));
  AOI22_X1  g712(.A1(new_n898), .A2(new_n889), .B1(new_n300), .B2(new_n302), .ZN(new_n899));
  OAI211_X1 g713(.A(new_n895), .B(new_n876), .C1(new_n899), .C2(new_n888), .ZN(new_n900));
  NAND2_X1  g714(.A1(new_n894), .A2(new_n900), .ZN(G54));
  AND2_X1   g715(.A1(KEYINPUT58), .A2(G475), .ZN(new_n902));
  NAND3_X1  g716(.A1(new_n896), .A2(G902), .A3(new_n902), .ZN(new_n903));
  INV_X1    g717(.A(new_n350), .ZN(new_n904));
  OR3_X1    g718(.A1(new_n903), .A2(KEYINPUT118), .A3(new_n904), .ZN(new_n905));
  OAI21_X1  g719(.A(KEYINPUT118), .B1(new_n903), .B2(new_n904), .ZN(new_n906));
  NAND2_X1  g720(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  NAND2_X1  g721(.A1(new_n907), .A2(new_n876), .ZN(new_n908));
  NAND2_X1  g722(.A1(new_n903), .A2(new_n904), .ZN(new_n909));
  XNOR2_X1  g723(.A(new_n909), .B(KEYINPUT119), .ZN(new_n910));
  NOR2_X1   g724(.A1(new_n908), .A2(new_n910), .ZN(G60));
  XOR2_X1   g725(.A(new_n580), .B(KEYINPUT59), .Z(new_n912));
  NAND3_X1  g726(.A1(new_n898), .A2(new_n578), .A3(new_n912), .ZN(new_n913));
  NAND2_X1  g727(.A1(new_n913), .A2(new_n876), .ZN(new_n914));
  AOI22_X1  g728(.A1(new_n862), .A2(KEYINPUT109), .B1(new_n806), .B2(new_n878), .ZN(new_n915));
  AOI21_X1  g729(.A(new_n865), .B1(new_n915), .B2(new_n864), .ZN(new_n916));
  NOR3_X1   g730(.A1(new_n817), .A2(KEYINPUT111), .A3(new_n818), .ZN(new_n917));
  OAI21_X1  g731(.A(new_n912), .B1(new_n916), .B2(new_n917), .ZN(new_n918));
  INV_X1    g732(.A(new_n578), .ZN(new_n919));
  AOI21_X1  g733(.A(new_n914), .B1(new_n918), .B2(new_n919), .ZN(G63));
  NAND2_X1  g734(.A1(G217), .A2(G902), .ZN(new_n921));
  XOR2_X1   g735(.A(new_n921), .B(KEYINPUT60), .Z(new_n922));
  NAND3_X1  g736(.A1(new_n896), .A2(new_n611), .A3(new_n922), .ZN(new_n923));
  AND2_X1   g737(.A1(new_n896), .A2(new_n922), .ZN(new_n924));
  OAI211_X1 g738(.A(new_n876), .B(new_n923), .C1(new_n924), .C2(new_n479), .ZN(new_n925));
  XOR2_X1   g739(.A(new_n925), .B(KEYINPUT61), .Z(G66));
  INV_X1    g740(.A(G224), .ZN(new_n927));
  OAI21_X1  g741(.A(G953), .B1(new_n366), .B2(new_n927), .ZN(new_n928));
  XNOR2_X1  g742(.A(new_n928), .B(KEYINPUT120), .ZN(new_n929));
  OAI21_X1  g743(.A(new_n929), .B1(new_n803), .B2(G953), .ZN(new_n930));
  XOR2_X1   g744(.A(new_n930), .B(KEYINPUT121), .Z(new_n931));
  OAI21_X1  g745(.A(new_n882), .B1(G898), .B2(new_n278), .ZN(new_n932));
  XNOR2_X1  g746(.A(new_n931), .B(new_n932), .ZN(G69));
  XOR2_X1   g747(.A(new_n501), .B(KEYINPUT122), .Z(new_n934));
  XOR2_X1   g748(.A(new_n934), .B(new_n318), .Z(new_n935));
  INV_X1    g749(.A(new_n935), .ZN(new_n936));
  NOR3_X1   g750(.A1(new_n631), .A2(new_n746), .A3(new_n791), .ZN(new_n937));
  NAND2_X1  g751(.A1(new_n937), .A2(new_n563), .ZN(new_n938));
  AND2_X1   g752(.A1(new_n756), .A2(new_n938), .ZN(new_n939));
  AND2_X1   g753(.A1(new_n781), .A2(new_n653), .ZN(new_n940));
  NAND2_X1  g754(.A1(new_n648), .A2(new_n940), .ZN(new_n941));
  OR2_X1    g755(.A1(new_n941), .A2(KEYINPUT62), .ZN(new_n942));
  NAND2_X1  g756(.A1(new_n941), .A2(KEYINPUT62), .ZN(new_n943));
  NAND4_X1  g757(.A1(new_n939), .A2(new_n942), .A3(new_n764), .A4(new_n943), .ZN(new_n944));
  AOI21_X1  g758(.A(new_n936), .B1(new_n944), .B2(new_n278), .ZN(new_n945));
  OR2_X1    g759(.A1(new_n945), .A2(KEYINPUT123), .ZN(new_n946));
  NAND2_X1  g760(.A1(new_n945), .A2(KEYINPUT123), .ZN(new_n947));
  NOR2_X1   g761(.A1(new_n278), .A2(G900), .ZN(new_n948));
  XNOR2_X1  g762(.A(new_n948), .B(KEYINPUT124), .ZN(new_n949));
  NAND3_X1  g763(.A1(new_n764), .A2(new_n802), .A3(new_n734), .ZN(new_n950));
  NAND3_X1  g764(.A1(new_n745), .A2(new_n774), .A3(new_n799), .ZN(new_n951));
  NAND3_X1  g765(.A1(new_n756), .A2(new_n951), .A3(new_n940), .ZN(new_n952));
  NOR2_X1   g766(.A1(new_n950), .A2(new_n952), .ZN(new_n953));
  OAI21_X1  g767(.A(new_n949), .B1(new_n953), .B2(G953), .ZN(new_n954));
  NAND2_X1  g768(.A1(new_n954), .A2(new_n936), .ZN(new_n955));
  NAND3_X1  g769(.A1(new_n946), .A2(new_n947), .A3(new_n955), .ZN(new_n956));
  INV_X1    g770(.A(KEYINPUT125), .ZN(new_n957));
  NAND3_X1  g771(.A1(new_n946), .A2(new_n947), .A3(new_n957), .ZN(new_n958));
  AOI21_X1  g772(.A(new_n278), .B1(G227), .B2(G900), .ZN(new_n959));
  NAND3_X1  g773(.A1(new_n956), .A2(new_n958), .A3(new_n959), .ZN(new_n960));
  INV_X1    g774(.A(KEYINPUT123), .ZN(new_n961));
  XNOR2_X1  g775(.A(new_n945), .B(new_n961), .ZN(new_n962));
  INV_X1    g776(.A(new_n959), .ZN(new_n963));
  OAI211_X1 g777(.A(new_n962), .B(new_n955), .C1(new_n957), .C2(new_n963), .ZN(new_n964));
  NAND2_X1  g778(.A1(new_n960), .A2(new_n964), .ZN(G72));
  NAND2_X1  g779(.A1(G472), .A2(G902), .ZN(new_n966));
  XOR2_X1   g780(.A(new_n966), .B(KEYINPUT63), .Z(new_n967));
  INV_X1    g781(.A(new_n953), .ZN(new_n968));
  OAI21_X1  g782(.A(new_n967), .B1(new_n968), .B2(new_n812), .ZN(new_n969));
  NOR2_X1   g783(.A1(new_n542), .A2(new_n506), .ZN(new_n970));
  AOI21_X1  g784(.A(new_n875), .B1(new_n969), .B2(new_n970), .ZN(new_n971));
  NAND2_X1  g785(.A1(new_n636), .A2(new_n544), .ZN(new_n972));
  OAI211_X1 g786(.A(new_n967), .B(new_n972), .C1(new_n860), .C2(new_n861), .ZN(new_n973));
  OAI21_X1  g787(.A(new_n967), .B1(new_n944), .B2(new_n812), .ZN(new_n974));
  NAND3_X1  g788(.A1(new_n974), .A2(new_n506), .A3(new_n542), .ZN(new_n975));
  NAND3_X1  g789(.A1(new_n971), .A2(new_n973), .A3(new_n975), .ZN(new_n976));
  NAND2_X1  g790(.A1(new_n976), .A2(KEYINPUT126), .ZN(new_n977));
  INV_X1    g791(.A(KEYINPUT126), .ZN(new_n978));
  NAND4_X1  g792(.A1(new_n971), .A2(new_n978), .A3(new_n973), .A4(new_n975), .ZN(new_n979));
  NAND2_X1  g793(.A1(new_n977), .A2(new_n979), .ZN(G57));
endmodule


