

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585;

  NOR2_X1 U323 ( .A1(n514), .A2(n549), .ZN(n533) );
  XNOR2_X1 U324 ( .A(n428), .B(n427), .ZN(n429) );
  XNOR2_X1 U325 ( .A(n311), .B(KEYINPUT31), .ZN(n291) );
  XOR2_X1 U326 ( .A(G183GAT), .B(KEYINPUT17), .Z(n292) );
  XNOR2_X1 U327 ( .A(KEYINPUT112), .B(KEYINPUT46), .ZN(n457) );
  XNOR2_X1 U328 ( .A(n458), .B(n457), .ZN(n459) );
  INV_X1 U329 ( .A(KEYINPUT54), .ZN(n472) );
  XNOR2_X1 U330 ( .A(n469), .B(KEYINPUT48), .ZN(n470) );
  INV_X1 U331 ( .A(G190GAT), .ZN(n425) );
  XNOR2_X1 U332 ( .A(n472), .B(KEYINPUT120), .ZN(n473) );
  XNOR2_X1 U333 ( .A(n471), .B(n470), .ZN(n534) );
  XNOR2_X1 U334 ( .A(n426), .B(n425), .ZN(n427) );
  XNOR2_X1 U335 ( .A(n474), .B(n473), .ZN(n475) );
  NOR2_X1 U336 ( .A1(n582), .A2(n445), .ZN(n446) );
  NOR2_X1 U337 ( .A1(n525), .A2(n478), .ZN(n567) );
  INV_X1 U338 ( .A(G43GAT), .ZN(n453) );
  XOR2_X1 U339 ( .A(n433), .B(n432), .Z(n510) );
  XNOR2_X1 U340 ( .A(n482), .B(G176GAT), .ZN(n483) );
  XNOR2_X1 U341 ( .A(n454), .B(n453), .ZN(n455) );
  XNOR2_X1 U342 ( .A(n484), .B(n483), .ZN(G1349GAT) );
  XNOR2_X1 U343 ( .A(n456), .B(n455), .ZN(G1330GAT) );
  XOR2_X1 U344 ( .A(G141GAT), .B(G22GAT), .Z(n393) );
  XNOR2_X1 U345 ( .A(G15GAT), .B(G1GAT), .ZN(n293) );
  XNOR2_X1 U346 ( .A(n293), .B(KEYINPUT67), .ZN(n352) );
  XNOR2_X1 U347 ( .A(n393), .B(n352), .ZN(n295) );
  NAND2_X1 U348 ( .A1(G229GAT), .A2(G233GAT), .ZN(n294) );
  XNOR2_X1 U349 ( .A(n295), .B(n294), .ZN(n296) );
  XOR2_X1 U350 ( .A(G169GAT), .B(G8GAT), .Z(n424) );
  XNOR2_X1 U351 ( .A(n296), .B(n424), .ZN(n298) );
  XNOR2_X1 U352 ( .A(G197GAT), .B(G113GAT), .ZN(n297) );
  XNOR2_X1 U353 ( .A(n298), .B(n297), .ZN(n308) );
  XOR2_X1 U354 ( .A(G43GAT), .B(G29GAT), .Z(n300) );
  XNOR2_X1 U355 ( .A(KEYINPUT7), .B(G50GAT), .ZN(n299) );
  XNOR2_X1 U356 ( .A(n300), .B(n299), .ZN(n301) );
  XOR2_X1 U357 ( .A(n301), .B(KEYINPUT66), .Z(n303) );
  XNOR2_X1 U358 ( .A(G36GAT), .B(KEYINPUT8), .ZN(n302) );
  XNOR2_X1 U359 ( .A(n303), .B(n302), .ZN(n333) );
  XOR2_X1 U360 ( .A(KEYINPUT68), .B(KEYINPUT65), .Z(n305) );
  XNOR2_X1 U361 ( .A(KEYINPUT30), .B(KEYINPUT29), .ZN(n304) );
  XNOR2_X1 U362 ( .A(n305), .B(n304), .ZN(n306) );
  XOR2_X1 U363 ( .A(n333), .B(n306), .Z(n307) );
  XNOR2_X1 U364 ( .A(n308), .B(n307), .ZN(n572) );
  XNOR2_X1 U365 ( .A(KEYINPUT69), .B(n572), .ZN(n537) );
  XOR2_X1 U366 ( .A(G176GAT), .B(G64GAT), .Z(n421) );
  XNOR2_X1 U367 ( .A(KEYINPUT32), .B(KEYINPUT33), .ZN(n310) );
  AND2_X1 U368 ( .A1(G230GAT), .A2(G233GAT), .ZN(n309) );
  XNOR2_X1 U369 ( .A(n310), .B(n309), .ZN(n311) );
  XOR2_X1 U370 ( .A(G78GAT), .B(G148GAT), .Z(n313) );
  XNOR2_X1 U371 ( .A(G106GAT), .B(G204GAT), .ZN(n312) );
  XNOR2_X1 U372 ( .A(n313), .B(n312), .ZN(n383) );
  XOR2_X1 U373 ( .A(G92GAT), .B(KEYINPUT72), .Z(n315) );
  XNOR2_X1 U374 ( .A(G99GAT), .B(G85GAT), .ZN(n314) );
  XNOR2_X1 U375 ( .A(n315), .B(n314), .ZN(n325) );
  XNOR2_X1 U376 ( .A(n383), .B(n325), .ZN(n316) );
  XNOR2_X1 U377 ( .A(n291), .B(n316), .ZN(n317) );
  XNOR2_X1 U378 ( .A(n421), .B(n317), .ZN(n321) );
  XOR2_X1 U379 ( .A(G120GAT), .B(G71GAT), .Z(n355) );
  XOR2_X1 U380 ( .A(KEYINPUT13), .B(KEYINPUT70), .Z(n319) );
  XNOR2_X1 U381 ( .A(G57GAT), .B(KEYINPUT71), .ZN(n318) );
  XNOR2_X1 U382 ( .A(n319), .B(n318), .ZN(n351) );
  XNOR2_X1 U383 ( .A(n355), .B(n351), .ZN(n320) );
  XNOR2_X1 U384 ( .A(n321), .B(n320), .ZN(n576) );
  AND2_X1 U385 ( .A1(n537), .A2(n576), .ZN(n489) );
  XNOR2_X1 U386 ( .A(KEYINPUT103), .B(KEYINPUT104), .ZN(n322) );
  XNOR2_X1 U387 ( .A(n322), .B(KEYINPUT37), .ZN(n447) );
  XOR2_X1 U388 ( .A(KEYINPUT10), .B(KEYINPUT75), .Z(n324) );
  XNOR2_X1 U389 ( .A(G218GAT), .B(KEYINPUT11), .ZN(n323) );
  XNOR2_X1 U390 ( .A(n324), .B(n323), .ZN(n326) );
  XOR2_X1 U391 ( .A(n326), .B(n325), .Z(n328) );
  XOR2_X1 U392 ( .A(G190GAT), .B(G134GAT), .Z(n356) );
  XOR2_X1 U393 ( .A(KEYINPUT73), .B(G162GAT), .Z(n392) );
  XNOR2_X1 U394 ( .A(n356), .B(n392), .ZN(n327) );
  XNOR2_X1 U395 ( .A(n328), .B(n327), .ZN(n332) );
  XOR2_X1 U396 ( .A(KEYINPUT74), .B(KEYINPUT9), .Z(n330) );
  NAND2_X1 U397 ( .A1(G232GAT), .A2(G233GAT), .ZN(n329) );
  XNOR2_X1 U398 ( .A(n330), .B(n329), .ZN(n331) );
  XOR2_X1 U399 ( .A(n332), .B(n331), .Z(n335) );
  XNOR2_X1 U400 ( .A(n333), .B(G106GAT), .ZN(n334) );
  XNOR2_X1 U401 ( .A(n335), .B(n334), .ZN(n558) );
  XNOR2_X1 U402 ( .A(KEYINPUT36), .B(n558), .ZN(n582) );
  XOR2_X1 U403 ( .A(G155GAT), .B(G78GAT), .Z(n337) );
  XNOR2_X1 U404 ( .A(G22GAT), .B(G211GAT), .ZN(n336) );
  XNOR2_X1 U405 ( .A(n337), .B(n336), .ZN(n341) );
  XOR2_X1 U406 ( .A(G64GAT), .B(G127GAT), .Z(n339) );
  XNOR2_X1 U407 ( .A(G183GAT), .B(G71GAT), .ZN(n338) );
  XNOR2_X1 U408 ( .A(n339), .B(n338), .ZN(n340) );
  XOR2_X1 U409 ( .A(n341), .B(n340), .Z(n346) );
  XOR2_X1 U410 ( .A(KEYINPUT15), .B(KEYINPUT76), .Z(n343) );
  NAND2_X1 U411 ( .A1(G231GAT), .A2(G233GAT), .ZN(n342) );
  XNOR2_X1 U412 ( .A(n343), .B(n342), .ZN(n344) );
  XNOR2_X1 U413 ( .A(KEYINPUT12), .B(n344), .ZN(n345) );
  XNOR2_X1 U414 ( .A(n346), .B(n345), .ZN(n350) );
  XOR2_X1 U415 ( .A(KEYINPUT14), .B(KEYINPUT77), .Z(n348) );
  XNOR2_X1 U416 ( .A(G8GAT), .B(KEYINPUT78), .ZN(n347) );
  XNOR2_X1 U417 ( .A(n348), .B(n347), .ZN(n349) );
  XOR2_X1 U418 ( .A(n350), .B(n349), .Z(n354) );
  XNOR2_X1 U419 ( .A(n352), .B(n351), .ZN(n353) );
  XNOR2_X1 U420 ( .A(n354), .B(n353), .ZN(n579) );
  XNOR2_X1 U421 ( .A(n356), .B(n355), .ZN(n359) );
  XOR2_X1 U422 ( .A(G127GAT), .B(KEYINPUT79), .Z(n358) );
  XNOR2_X1 U423 ( .A(G113GAT), .B(KEYINPUT0), .ZN(n357) );
  XNOR2_X1 U424 ( .A(n358), .B(n357), .ZN(n405) );
  XNOR2_X1 U425 ( .A(n359), .B(n405), .ZN(n364) );
  XNOR2_X1 U426 ( .A(KEYINPUT18), .B(KEYINPUT19), .ZN(n360) );
  XNOR2_X1 U427 ( .A(n292), .B(n360), .ZN(n420) );
  XOR2_X1 U428 ( .A(G15GAT), .B(n420), .Z(n362) );
  NAND2_X1 U429 ( .A1(G227GAT), .A2(G233GAT), .ZN(n361) );
  XNOR2_X1 U430 ( .A(n362), .B(n361), .ZN(n363) );
  XOR2_X1 U431 ( .A(n364), .B(n363), .Z(n372) );
  XOR2_X1 U432 ( .A(KEYINPUT82), .B(G99GAT), .Z(n366) );
  XNOR2_X1 U433 ( .A(G169GAT), .B(G43GAT), .ZN(n365) );
  XNOR2_X1 U434 ( .A(n366), .B(n365), .ZN(n370) );
  XOR2_X1 U435 ( .A(KEYINPUT80), .B(G176GAT), .Z(n368) );
  XNOR2_X1 U436 ( .A(KEYINPUT20), .B(KEYINPUT81), .ZN(n367) );
  XNOR2_X1 U437 ( .A(n368), .B(n367), .ZN(n369) );
  XNOR2_X1 U438 ( .A(n370), .B(n369), .ZN(n371) );
  XNOR2_X1 U439 ( .A(n372), .B(n371), .ZN(n525) );
  XOR2_X1 U440 ( .A(KEYINPUT87), .B(KEYINPUT23), .Z(n374) );
  XNOR2_X1 U441 ( .A(G50GAT), .B(KEYINPUT22), .ZN(n373) );
  XNOR2_X1 U442 ( .A(n374), .B(n373), .ZN(n378) );
  XOR2_X1 U443 ( .A(KEYINPUT24), .B(KEYINPUT89), .Z(n376) );
  XNOR2_X1 U444 ( .A(KEYINPUT90), .B(KEYINPUT83), .ZN(n375) );
  XNOR2_X1 U445 ( .A(n376), .B(n375), .ZN(n377) );
  XOR2_X1 U446 ( .A(n378), .B(n377), .Z(n388) );
  XNOR2_X1 U447 ( .A(G211GAT), .B(KEYINPUT21), .ZN(n379) );
  XNOR2_X1 U448 ( .A(n379), .B(KEYINPUT84), .ZN(n380) );
  XOR2_X1 U449 ( .A(n380), .B(KEYINPUT85), .Z(n382) );
  XNOR2_X1 U450 ( .A(G197GAT), .B(G218GAT), .ZN(n381) );
  XNOR2_X1 U451 ( .A(n382), .B(n381), .ZN(n431) );
  XOR2_X1 U452 ( .A(KEYINPUT88), .B(n383), .Z(n385) );
  NAND2_X1 U453 ( .A1(G228GAT), .A2(G233GAT), .ZN(n384) );
  XNOR2_X1 U454 ( .A(n385), .B(n384), .ZN(n386) );
  XNOR2_X1 U455 ( .A(n431), .B(n386), .ZN(n387) );
  XNOR2_X1 U456 ( .A(n388), .B(n387), .ZN(n391) );
  XOR2_X1 U457 ( .A(G155GAT), .B(KEYINPUT2), .Z(n390) );
  XNOR2_X1 U458 ( .A(KEYINPUT3), .B(KEYINPUT86), .ZN(n389) );
  XNOR2_X1 U459 ( .A(n390), .B(n389), .ZN(n404) );
  XOR2_X1 U460 ( .A(n391), .B(n404), .Z(n395) );
  XNOR2_X1 U461 ( .A(n393), .B(n392), .ZN(n394) );
  XNOR2_X1 U462 ( .A(n395), .B(n394), .ZN(n476) );
  XOR2_X1 U463 ( .A(n476), .B(KEYINPUT28), .Z(n514) );
  XOR2_X1 U464 ( .A(KEYINPUT95), .B(KEYINPUT6), .Z(n397) );
  XNOR2_X1 U465 ( .A(KEYINPUT5), .B(G57GAT), .ZN(n396) );
  XNOR2_X1 U466 ( .A(n397), .B(n396), .ZN(n409) );
  XOR2_X1 U467 ( .A(KEYINPUT1), .B(KEYINPUT4), .Z(n399) );
  XNOR2_X1 U468 ( .A(G1GAT), .B(G120GAT), .ZN(n398) );
  XNOR2_X1 U469 ( .A(n399), .B(n398), .ZN(n403) );
  XOR2_X1 U470 ( .A(KEYINPUT91), .B(KEYINPUT94), .Z(n401) );
  XNOR2_X1 U471 ( .A(KEYINPUT92), .B(KEYINPUT93), .ZN(n400) );
  XNOR2_X1 U472 ( .A(n401), .B(n400), .ZN(n402) );
  XOR2_X1 U473 ( .A(n403), .B(n402), .Z(n407) );
  XNOR2_X1 U474 ( .A(n405), .B(n404), .ZN(n406) );
  XNOR2_X1 U475 ( .A(n407), .B(n406), .ZN(n408) );
  XNOR2_X1 U476 ( .A(n409), .B(n408), .ZN(n417) );
  NAND2_X1 U477 ( .A1(G225GAT), .A2(G233GAT), .ZN(n415) );
  XOR2_X1 U478 ( .A(G85GAT), .B(G148GAT), .Z(n411) );
  XNOR2_X1 U479 ( .A(G29GAT), .B(G141GAT), .ZN(n410) );
  XNOR2_X1 U480 ( .A(n411), .B(n410), .ZN(n413) );
  XOR2_X1 U481 ( .A(G134GAT), .B(G162GAT), .Z(n412) );
  XNOR2_X1 U482 ( .A(n413), .B(n412), .ZN(n414) );
  XNOR2_X1 U483 ( .A(n415), .B(n414), .ZN(n416) );
  XNOR2_X1 U484 ( .A(n417), .B(n416), .ZN(n507) );
  XOR2_X1 U485 ( .A(KEYINPUT96), .B(KEYINPUT76), .Z(n419) );
  XNOR2_X1 U486 ( .A(G204GAT), .B(G92GAT), .ZN(n418) );
  XNOR2_X1 U487 ( .A(n419), .B(n418), .ZN(n430) );
  XOR2_X1 U488 ( .A(n421), .B(n420), .Z(n423) );
  NAND2_X1 U489 ( .A1(G226GAT), .A2(G233GAT), .ZN(n422) );
  XNOR2_X1 U490 ( .A(n423), .B(n422), .ZN(n428) );
  XNOR2_X1 U491 ( .A(G36GAT), .B(n424), .ZN(n426) );
  XNOR2_X1 U492 ( .A(n430), .B(n429), .ZN(n433) );
  INV_X1 U493 ( .A(n431), .ZN(n432) );
  INV_X1 U494 ( .A(n510), .ZN(n522) );
  XOR2_X1 U495 ( .A(KEYINPUT27), .B(n522), .Z(n436) );
  NAND2_X1 U496 ( .A1(n507), .A2(n436), .ZN(n549) );
  NAND2_X1 U497 ( .A1(n525), .A2(n533), .ZN(n434) );
  XOR2_X1 U498 ( .A(KEYINPUT97), .B(n434), .Z(n444) );
  INV_X1 U499 ( .A(n525), .ZN(n532) );
  NOR2_X1 U500 ( .A1(n532), .A2(n476), .ZN(n435) );
  XNOR2_X1 U501 ( .A(n435), .B(KEYINPUT26), .ZN(n570) );
  NAND2_X1 U502 ( .A1(n436), .A2(n570), .ZN(n441) );
  NAND2_X1 U503 ( .A1(n532), .A2(n510), .ZN(n437) );
  NAND2_X1 U504 ( .A1(n437), .A2(n476), .ZN(n438) );
  XNOR2_X1 U505 ( .A(n438), .B(KEYINPUT25), .ZN(n439) );
  XOR2_X1 U506 ( .A(KEYINPUT98), .B(n439), .Z(n440) );
  NAND2_X1 U507 ( .A1(n441), .A2(n440), .ZN(n442) );
  INV_X1 U508 ( .A(n507), .ZN(n519) );
  NAND2_X1 U509 ( .A1(n442), .A2(n519), .ZN(n443) );
  NAND2_X1 U510 ( .A1(n444), .A2(n443), .ZN(n486) );
  NAND2_X1 U511 ( .A1(n579), .A2(n486), .ZN(n445) );
  XNOR2_X1 U512 ( .A(n447), .B(n446), .ZN(n517) );
  AND2_X1 U513 ( .A1(n489), .A2(n517), .ZN(n448) );
  XNOR2_X1 U514 ( .A(n448), .B(KEYINPUT38), .ZN(n501) );
  NAND2_X1 U515 ( .A1(n501), .A2(n507), .ZN(n452) );
  XOR2_X1 U516 ( .A(KEYINPUT39), .B(KEYINPUT105), .Z(n450) );
  INV_X1 U517 ( .A(G29GAT), .ZN(n449) );
  XNOR2_X1 U518 ( .A(n450), .B(n449), .ZN(n451) );
  XNOR2_X1 U519 ( .A(n452), .B(n451), .ZN(G1328GAT) );
  NAND2_X1 U520 ( .A1(n501), .A2(n532), .ZN(n456) );
  XOR2_X1 U521 ( .A(KEYINPUT40), .B(KEYINPUT106), .Z(n454) );
  XNOR2_X1 U522 ( .A(n576), .B(KEYINPUT41), .ZN(n539) );
  INV_X1 U523 ( .A(n572), .ZN(n504) );
  NAND2_X1 U524 ( .A1(n539), .A2(n504), .ZN(n458) );
  NAND2_X1 U525 ( .A1(n459), .A2(n579), .ZN(n460) );
  XNOR2_X1 U526 ( .A(n460), .B(KEYINPUT113), .ZN(n461) );
  NAND2_X1 U527 ( .A1(n461), .A2(n558), .ZN(n462) );
  XNOR2_X1 U528 ( .A(n462), .B(KEYINPUT47), .ZN(n468) );
  NOR2_X1 U529 ( .A1(n579), .A2(n582), .ZN(n464) );
  XNOR2_X1 U530 ( .A(KEYINPUT45), .B(KEYINPUT114), .ZN(n463) );
  XNOR2_X1 U531 ( .A(n464), .B(n463), .ZN(n465) );
  NAND2_X1 U532 ( .A1(n576), .A2(n465), .ZN(n466) );
  NOR2_X1 U533 ( .A1(n466), .A2(n537), .ZN(n467) );
  NOR2_X1 U534 ( .A1(n468), .A2(n467), .ZN(n471) );
  XOR2_X1 U535 ( .A(KEYINPUT64), .B(KEYINPUT115), .Z(n469) );
  NOR2_X1 U536 ( .A1(n534), .A2(n522), .ZN(n474) );
  NOR2_X1 U537 ( .A1(n507), .A2(n475), .ZN(n571) );
  AND2_X1 U538 ( .A1(n476), .A2(n571), .ZN(n477) );
  XNOR2_X1 U539 ( .A(n477), .B(KEYINPUT55), .ZN(n478) );
  NAND2_X1 U540 ( .A1(n567), .A2(n537), .ZN(n481) );
  XOR2_X1 U541 ( .A(G169GAT), .B(KEYINPUT121), .Z(n479) );
  XNOR2_X1 U542 ( .A(n479), .B(KEYINPUT122), .ZN(n480) );
  XNOR2_X1 U543 ( .A(n481), .B(n480), .ZN(G1348GAT) );
  NAND2_X1 U544 ( .A1(n567), .A2(n539), .ZN(n484) );
  XOR2_X1 U545 ( .A(KEYINPUT56), .B(KEYINPUT57), .Z(n482) );
  INV_X1 U546 ( .A(n558), .ZN(n566) );
  NOR2_X1 U547 ( .A1(n579), .A2(n566), .ZN(n485) );
  XNOR2_X1 U548 ( .A(KEYINPUT16), .B(n485), .ZN(n487) );
  NAND2_X1 U549 ( .A1(n487), .A2(n486), .ZN(n488) );
  XNOR2_X1 U550 ( .A(n488), .B(KEYINPUT99), .ZN(n505) );
  NAND2_X1 U551 ( .A1(n489), .A2(n505), .ZN(n497) );
  NOR2_X1 U552 ( .A1(n519), .A2(n497), .ZN(n491) );
  XNOR2_X1 U553 ( .A(KEYINPUT34), .B(KEYINPUT100), .ZN(n490) );
  XNOR2_X1 U554 ( .A(n491), .B(n490), .ZN(n492) );
  XOR2_X1 U555 ( .A(G1GAT), .B(n492), .Z(G1324GAT) );
  NOR2_X1 U556 ( .A1(n522), .A2(n497), .ZN(n493) );
  XOR2_X1 U557 ( .A(G8GAT), .B(n493), .Z(G1325GAT) );
  NOR2_X1 U558 ( .A1(n525), .A2(n497), .ZN(n495) );
  XNOR2_X1 U559 ( .A(KEYINPUT101), .B(KEYINPUT35), .ZN(n494) );
  XNOR2_X1 U560 ( .A(n495), .B(n494), .ZN(n496) );
  XOR2_X1 U561 ( .A(G15GAT), .B(n496), .Z(G1326GAT) );
  INV_X1 U562 ( .A(n514), .ZN(n529) );
  NOR2_X1 U563 ( .A1(n529), .A2(n497), .ZN(n498) );
  XOR2_X1 U564 ( .A(KEYINPUT102), .B(n498), .Z(n499) );
  XNOR2_X1 U565 ( .A(G22GAT), .B(n499), .ZN(G1327GAT) );
  NAND2_X1 U566 ( .A1(n501), .A2(n510), .ZN(n500) );
  XNOR2_X1 U567 ( .A(n500), .B(G36GAT), .ZN(G1329GAT) );
  XOR2_X1 U568 ( .A(G50GAT), .B(KEYINPUT107), .Z(n503) );
  NAND2_X1 U569 ( .A1(n514), .A2(n501), .ZN(n502) );
  XNOR2_X1 U570 ( .A(n503), .B(n502), .ZN(G1331GAT) );
  INV_X1 U571 ( .A(n539), .ZN(n552) );
  NOR2_X1 U572 ( .A1(n504), .A2(n552), .ZN(n518) );
  NAND2_X1 U573 ( .A1(n505), .A2(n518), .ZN(n506) );
  XOR2_X1 U574 ( .A(KEYINPUT108), .B(n506), .Z(n513) );
  NAND2_X1 U575 ( .A1(n513), .A2(n507), .ZN(n508) );
  XNOR2_X1 U576 ( .A(n508), .B(KEYINPUT42), .ZN(n509) );
  XNOR2_X1 U577 ( .A(G57GAT), .B(n509), .ZN(G1332GAT) );
  NAND2_X1 U578 ( .A1(n513), .A2(n510), .ZN(n511) );
  XNOR2_X1 U579 ( .A(n511), .B(G64GAT), .ZN(G1333GAT) );
  NAND2_X1 U580 ( .A1(n513), .A2(n532), .ZN(n512) );
  XNOR2_X1 U581 ( .A(n512), .B(G71GAT), .ZN(G1334GAT) );
  XOR2_X1 U582 ( .A(G78GAT), .B(KEYINPUT43), .Z(n516) );
  NAND2_X1 U583 ( .A1(n514), .A2(n513), .ZN(n515) );
  XNOR2_X1 U584 ( .A(n516), .B(n515), .ZN(G1335GAT) );
  NAND2_X1 U585 ( .A1(n518), .A2(n517), .ZN(n528) );
  NOR2_X1 U586 ( .A1(n519), .A2(n528), .ZN(n521) );
  XNOR2_X1 U587 ( .A(G85GAT), .B(KEYINPUT109), .ZN(n520) );
  XNOR2_X1 U588 ( .A(n521), .B(n520), .ZN(G1336GAT) );
  NOR2_X1 U589 ( .A1(n522), .A2(n528), .ZN(n523) );
  XOR2_X1 U590 ( .A(KEYINPUT110), .B(n523), .Z(n524) );
  XNOR2_X1 U591 ( .A(G92GAT), .B(n524), .ZN(G1337GAT) );
  NOR2_X1 U592 ( .A1(n525), .A2(n528), .ZN(n527) );
  XNOR2_X1 U593 ( .A(G99GAT), .B(KEYINPUT111), .ZN(n526) );
  XNOR2_X1 U594 ( .A(n527), .B(n526), .ZN(G1338GAT) );
  NOR2_X1 U595 ( .A1(n529), .A2(n528), .ZN(n530) );
  XOR2_X1 U596 ( .A(KEYINPUT44), .B(n530), .Z(n531) );
  XNOR2_X1 U597 ( .A(G106GAT), .B(n531), .ZN(G1339GAT) );
  NAND2_X1 U598 ( .A1(n533), .A2(n532), .ZN(n535) );
  NOR2_X1 U599 ( .A1(n535), .A2(n534), .ZN(n536) );
  XNOR2_X1 U600 ( .A(n536), .B(KEYINPUT116), .ZN(n545) );
  NAND2_X1 U601 ( .A1(n537), .A2(n545), .ZN(n538) );
  XNOR2_X1 U602 ( .A(G113GAT), .B(n538), .ZN(G1340GAT) );
  XOR2_X1 U603 ( .A(KEYINPUT49), .B(KEYINPUT117), .Z(n541) );
  NAND2_X1 U604 ( .A1(n545), .A2(n539), .ZN(n540) );
  XNOR2_X1 U605 ( .A(n541), .B(n540), .ZN(n542) );
  XOR2_X1 U606 ( .A(G120GAT), .B(n542), .Z(G1341GAT) );
  INV_X1 U607 ( .A(n579), .ZN(n561) );
  NAND2_X1 U608 ( .A1(n545), .A2(n561), .ZN(n543) );
  XNOR2_X1 U609 ( .A(n543), .B(KEYINPUT50), .ZN(n544) );
  XNOR2_X1 U610 ( .A(G127GAT), .B(n544), .ZN(G1342GAT) );
  XOR2_X1 U611 ( .A(KEYINPUT118), .B(KEYINPUT51), .Z(n547) );
  NAND2_X1 U612 ( .A1(n545), .A2(n566), .ZN(n546) );
  XNOR2_X1 U613 ( .A(n547), .B(n546), .ZN(n548) );
  XNOR2_X1 U614 ( .A(G134GAT), .B(n548), .ZN(G1343GAT) );
  NOR2_X1 U615 ( .A1(n534), .A2(n549), .ZN(n550) );
  NAND2_X1 U616 ( .A1(n550), .A2(n570), .ZN(n557) );
  NOR2_X1 U617 ( .A1(n572), .A2(n557), .ZN(n551) );
  XOR2_X1 U618 ( .A(G141GAT), .B(n551), .Z(G1344GAT) );
  NOR2_X1 U619 ( .A1(n552), .A2(n557), .ZN(n554) );
  XNOR2_X1 U620 ( .A(KEYINPUT53), .B(KEYINPUT52), .ZN(n553) );
  XNOR2_X1 U621 ( .A(n554), .B(n553), .ZN(n555) );
  XNOR2_X1 U622 ( .A(G148GAT), .B(n555), .ZN(G1345GAT) );
  NOR2_X1 U623 ( .A1(n579), .A2(n557), .ZN(n556) );
  XOR2_X1 U624 ( .A(G155GAT), .B(n556), .Z(G1346GAT) );
  NOR2_X1 U625 ( .A1(n558), .A2(n557), .ZN(n560) );
  XNOR2_X1 U626 ( .A(G162GAT), .B(KEYINPUT119), .ZN(n559) );
  XNOR2_X1 U627 ( .A(n560), .B(n559), .ZN(G1347GAT) );
  XOR2_X1 U628 ( .A(G183GAT), .B(KEYINPUT123), .Z(n563) );
  NAND2_X1 U629 ( .A1(n567), .A2(n561), .ZN(n562) );
  XNOR2_X1 U630 ( .A(n563), .B(n562), .ZN(G1350GAT) );
  XNOR2_X1 U631 ( .A(G190GAT), .B(KEYINPUT125), .ZN(n564) );
  XNOR2_X1 U632 ( .A(n564), .B(KEYINPUT124), .ZN(n565) );
  XOR2_X1 U633 ( .A(KEYINPUT58), .B(n565), .Z(n569) );
  NAND2_X1 U634 ( .A1(n567), .A2(n566), .ZN(n568) );
  XNOR2_X1 U635 ( .A(n569), .B(n568), .ZN(G1351GAT) );
  NAND2_X1 U636 ( .A1(n571), .A2(n570), .ZN(n581) );
  NOR2_X1 U637 ( .A1(n572), .A2(n581), .ZN(n574) );
  XNOR2_X1 U638 ( .A(KEYINPUT60), .B(KEYINPUT59), .ZN(n573) );
  XNOR2_X1 U639 ( .A(n574), .B(n573), .ZN(n575) );
  XNOR2_X1 U640 ( .A(G197GAT), .B(n575), .ZN(G1352GAT) );
  NOR2_X1 U641 ( .A1(n576), .A2(n581), .ZN(n578) );
  XNOR2_X1 U642 ( .A(G204GAT), .B(KEYINPUT61), .ZN(n577) );
  XNOR2_X1 U643 ( .A(n578), .B(n577), .ZN(G1353GAT) );
  NOR2_X1 U644 ( .A1(n579), .A2(n581), .ZN(n580) );
  XOR2_X1 U645 ( .A(G211GAT), .B(n580), .Z(G1354GAT) );
  NOR2_X1 U646 ( .A1(n582), .A2(n581), .ZN(n584) );
  XNOR2_X1 U647 ( .A(KEYINPUT126), .B(KEYINPUT62), .ZN(n583) );
  XNOR2_X1 U648 ( .A(n584), .B(n583), .ZN(n585) );
  XOR2_X1 U649 ( .A(G218GAT), .B(n585), .Z(G1355GAT) );
endmodule

