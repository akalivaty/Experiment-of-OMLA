//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 0 1 0 0 0 0 1 1 0 0 1 0 0 1 0 0 1 0 1 0 1 0 1 0 1 1 0 0 0 1 1 1 1 1 0 1 0 1 0 1 0 1 1 1 1 0 1 1 1 1 1 1 1 1 0 1 0 0 1 0 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:29:26 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n437, new_n444, new_n449, new_n452, new_n454, new_n455,
    new_n456, new_n459, new_n460, new_n461, new_n462, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n523, new_n524, new_n525,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n531, new_n532,
    new_n533, new_n534, new_n535, new_n537, new_n538, new_n539, new_n540,
    new_n541, new_n544, new_n545, new_n546, new_n547, new_n548, new_n549,
    new_n550, new_n551, new_n552, new_n555, new_n556, new_n558, new_n559,
    new_n560, new_n561, new_n562, new_n563, new_n564, new_n565, new_n566,
    new_n567, new_n568, new_n569, new_n570, new_n571, new_n572, new_n573,
    new_n574, new_n575, new_n576, new_n577, new_n579, new_n580, new_n581,
    new_n582, new_n583, new_n586, new_n587, new_n588, new_n589, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n619, new_n621, new_n622, new_n623, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1217, new_n1218,
    new_n1219, new_n1220, new_n1221, new_n1222, new_n1223, new_n1224,
    new_n1225, new_n1226, new_n1227, new_n1228, new_n1229, new_n1230,
    new_n1231, new_n1232, new_n1233, new_n1234, new_n1235, new_n1236,
    new_n1237, new_n1238, new_n1241;
  XOR2_X1   g000(.A(KEYINPUT64), .B(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  XOR2_X1   g002(.A(KEYINPUT65), .B(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(new_n436));
  INV_X1    g011(.A(KEYINPUT66), .ZN(new_n437));
  XNOR2_X1  g012(.A(new_n436), .B(new_n437), .ZN(G220));
  INV_X1    g013(.A(G96), .ZN(G221));
  INV_X1    g014(.A(G69), .ZN(G235));
  INV_X1    g015(.A(G120), .ZN(G236));
  INV_X1    g016(.A(G57), .ZN(G237));
  INV_X1    g017(.A(G108), .ZN(G238));
  AND2_X1   g018(.A1(G2072), .A2(G2078), .ZN(new_n444));
  NAND3_X1  g019(.A1(new_n444), .A2(G2084), .A3(G2090), .ZN(G158));
  NAND3_X1  g020(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g021(.A(G452), .Z(G391));
  AND2_X1   g022(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g023(.A1(G7), .A2(G661), .ZN(new_n449));
  XOR2_X1   g024(.A(new_n449), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g025(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g026(.A1(G7), .A2(G661), .A3(G2106), .ZN(new_n452));
  XNOR2_X1  g027(.A(new_n452), .B(KEYINPUT67), .ZN(G217));
  NOR4_X1   g028(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n454));
  XOR2_X1   g029(.A(new_n454), .B(KEYINPUT2), .Z(new_n455));
  NAND4_X1  g030(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n456));
  NOR2_X1   g031(.A1(new_n455), .A2(new_n456), .ZN(G325));
  INV_X1    g032(.A(G325), .ZN(G261));
  NAND2_X1  g033(.A1(new_n455), .A2(G2106), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n456), .A2(G567), .ZN(new_n460));
  XOR2_X1   g035(.A(new_n460), .B(KEYINPUT68), .Z(new_n461));
  NAND2_X1  g036(.A1(new_n459), .A2(new_n461), .ZN(new_n462));
  INV_X1    g037(.A(new_n462), .ZN(G319));
  XNOR2_X1  g038(.A(KEYINPUT3), .B(G2104), .ZN(new_n464));
  INV_X1    g039(.A(G2105), .ZN(new_n465));
  NAND3_X1  g040(.A1(new_n464), .A2(G137), .A3(new_n465), .ZN(new_n466));
  AND2_X1   g041(.A1(new_n465), .A2(G2104), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n467), .A2(G101), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n466), .A2(new_n468), .ZN(new_n469));
  AND2_X1   g044(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n470));
  NOR2_X1   g045(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n471));
  OAI21_X1  g046(.A(G125), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  NAND2_X1  g047(.A1(G113), .A2(G2104), .ZN(new_n473));
  AOI21_X1  g048(.A(new_n465), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  NOR2_X1   g049(.A1(new_n469), .A2(new_n474), .ZN(G160));
  NOR2_X1   g050(.A1(new_n470), .A2(new_n471), .ZN(new_n476));
  NOR2_X1   g051(.A1(new_n476), .A2(KEYINPUT69), .ZN(new_n477));
  INV_X1    g052(.A(KEYINPUT69), .ZN(new_n478));
  NOR2_X1   g053(.A1(new_n464), .A2(new_n478), .ZN(new_n479));
  OAI21_X1  g054(.A(new_n465), .B1(new_n477), .B2(new_n479), .ZN(new_n480));
  INV_X1    g055(.A(new_n480), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n481), .A2(G136), .ZN(new_n482));
  OAI21_X1  g057(.A(G2105), .B1(new_n477), .B2(new_n479), .ZN(new_n483));
  INV_X1    g058(.A(new_n483), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n484), .A2(G124), .ZN(new_n485));
  OR2_X1    g060(.A1(G100), .A2(G2105), .ZN(new_n486));
  OAI211_X1 g061(.A(new_n486), .B(G2104), .C1(G112), .C2(new_n465), .ZN(new_n487));
  NAND3_X1  g062(.A1(new_n482), .A2(new_n485), .A3(new_n487), .ZN(new_n488));
  INV_X1    g063(.A(new_n488), .ZN(G162));
  NAND2_X1  g064(.A1(G126), .A2(G2105), .ZN(new_n490));
  NOR2_X1   g065(.A1(new_n465), .A2(G114), .ZN(new_n491));
  OAI21_X1  g066(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n492));
  OAI22_X1  g067(.A1(new_n476), .A2(new_n490), .B1(new_n491), .B2(new_n492), .ZN(new_n493));
  OAI21_X1  g068(.A(new_n465), .B1(new_n470), .B2(new_n471), .ZN(new_n494));
  INV_X1    g069(.A(G138), .ZN(new_n495));
  NOR2_X1   g070(.A1(new_n495), .A2(KEYINPUT70), .ZN(new_n496));
  INV_X1    g071(.A(new_n496), .ZN(new_n497));
  OAI21_X1  g072(.A(KEYINPUT4), .B1(new_n494), .B2(new_n497), .ZN(new_n498));
  INV_X1    g073(.A(KEYINPUT4), .ZN(new_n499));
  NAND4_X1  g074(.A1(new_n464), .A2(new_n499), .A3(new_n465), .A4(new_n496), .ZN(new_n500));
  AOI21_X1  g075(.A(new_n493), .B1(new_n498), .B2(new_n500), .ZN(G164));
  INV_X1    g076(.A(KEYINPUT5), .ZN(new_n502));
  INV_X1    g077(.A(G543), .ZN(new_n503));
  NAND2_X1  g078(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  NAND2_X1  g079(.A1(KEYINPUT5), .A2(G543), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  AOI22_X1  g081(.A1(new_n506), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n507));
  INV_X1    g082(.A(G651), .ZN(new_n508));
  NOR2_X1   g083(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  INV_X1    g084(.A(KEYINPUT6), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n510), .A2(new_n508), .ZN(new_n511));
  NAND2_X1  g086(.A1(KEYINPUT6), .A2(G651), .ZN(new_n512));
  AOI21_X1  g087(.A(new_n503), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n513), .A2(G50), .ZN(new_n514));
  INV_X1    g089(.A(G88), .ZN(new_n515));
  NOR2_X1   g090(.A1(KEYINPUT5), .A2(G543), .ZN(new_n516));
  AND2_X1   g091(.A1(KEYINPUT5), .A2(G543), .ZN(new_n517));
  AND2_X1   g092(.A1(KEYINPUT6), .A2(G651), .ZN(new_n518));
  NOR2_X1   g093(.A1(KEYINPUT6), .A2(G651), .ZN(new_n519));
  OAI22_X1  g094(.A1(new_n516), .A2(new_n517), .B1(new_n518), .B2(new_n519), .ZN(new_n520));
  OAI21_X1  g095(.A(new_n514), .B1(new_n515), .B2(new_n520), .ZN(new_n521));
  NOR2_X1   g096(.A1(new_n509), .A2(new_n521), .ZN(G166));
  NAND3_X1  g097(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n523), .A2(KEYINPUT7), .ZN(new_n524));
  INV_X1    g099(.A(KEYINPUT7), .ZN(new_n525));
  NAND4_X1  g100(.A1(new_n525), .A2(G76), .A3(G543), .A4(G651), .ZN(new_n526));
  NAND2_X1  g101(.A1(new_n524), .A2(new_n526), .ZN(new_n527));
  OAI211_X1 g102(.A(G51), .B(G543), .C1(new_n518), .C2(new_n519), .ZN(new_n528));
  NAND2_X1  g103(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  INV_X1    g104(.A(new_n529), .ZN(new_n530));
  OAI21_X1  g105(.A(G89), .B1(new_n518), .B2(new_n519), .ZN(new_n531));
  NAND2_X1  g106(.A1(G63), .A2(G651), .ZN(new_n532));
  NAND2_X1  g107(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  NAND2_X1  g108(.A1(new_n533), .A2(new_n506), .ZN(new_n534));
  NAND2_X1  g109(.A1(new_n530), .A2(new_n534), .ZN(new_n535));
  INV_X1    g110(.A(new_n535), .ZN(G168));
  AND2_X1   g111(.A1(new_n506), .A2(G64), .ZN(new_n537));
  AND2_X1   g112(.A1(G77), .A2(G543), .ZN(new_n538));
  OAI21_X1  g113(.A(G651), .B1(new_n537), .B2(new_n538), .ZN(new_n539));
  AOI22_X1  g114(.A1(new_n504), .A2(new_n505), .B1(new_n511), .B2(new_n512), .ZN(new_n540));
  AOI22_X1  g115(.A1(new_n540), .A2(G90), .B1(new_n513), .B2(G52), .ZN(new_n541));
  NAND2_X1  g116(.A1(new_n539), .A2(new_n541), .ZN(G301));
  INV_X1    g117(.A(G301), .ZN(G171));
  AOI22_X1  g118(.A1(new_n540), .A2(G81), .B1(new_n513), .B2(G43), .ZN(new_n544));
  OAI21_X1  g119(.A(G56), .B1(new_n517), .B2(new_n516), .ZN(new_n545));
  NAND2_X1  g120(.A1(G68), .A2(G543), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  AOI21_X1  g122(.A(KEYINPUT71), .B1(new_n547), .B2(G651), .ZN(new_n548));
  INV_X1    g123(.A(KEYINPUT71), .ZN(new_n549));
  AOI211_X1 g124(.A(new_n549), .B(new_n508), .C1(new_n545), .C2(new_n546), .ZN(new_n550));
  OAI21_X1  g125(.A(new_n544), .B1(new_n548), .B2(new_n550), .ZN(new_n551));
  INV_X1    g126(.A(new_n551), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n552), .A2(G860), .ZN(G153));
  NAND4_X1  g128(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g129(.A1(G1), .A2(G3), .ZN(new_n555));
  XNOR2_X1  g130(.A(new_n555), .B(KEYINPUT8), .ZN(new_n556));
  NAND4_X1  g131(.A1(G319), .A2(G483), .A3(G661), .A4(new_n556), .ZN(G188));
  NAND2_X1  g132(.A1(G78), .A2(G543), .ZN(new_n558));
  NOR2_X1   g133(.A1(new_n517), .A2(new_n516), .ZN(new_n559));
  INV_X1    g134(.A(G65), .ZN(new_n560));
  OAI21_X1  g135(.A(new_n558), .B1(new_n559), .B2(new_n560), .ZN(new_n561));
  AOI22_X1  g136(.A1(new_n561), .A2(G651), .B1(new_n540), .B2(G91), .ZN(new_n562));
  AND2_X1   g137(.A1(G53), .A2(G543), .ZN(new_n563));
  NAND2_X1  g138(.A1(KEYINPUT72), .A2(KEYINPUT9), .ZN(new_n564));
  OAI211_X1 g139(.A(new_n563), .B(new_n564), .C1(new_n518), .C2(new_n519), .ZN(new_n565));
  INV_X1    g140(.A(KEYINPUT73), .ZN(new_n566));
  NAND2_X1  g141(.A1(G53), .A2(G543), .ZN(new_n567));
  AOI21_X1  g142(.A(new_n567), .B1(new_n511), .B2(new_n512), .ZN(new_n568));
  INV_X1    g143(.A(new_n564), .ZN(new_n569));
  NOR2_X1   g144(.A1(KEYINPUT72), .A2(KEYINPUT9), .ZN(new_n570));
  NOR2_X1   g145(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  OAI211_X1 g146(.A(new_n565), .B(new_n566), .C1(new_n568), .C2(new_n571), .ZN(new_n572));
  INV_X1    g147(.A(new_n572), .ZN(new_n573));
  OAI21_X1  g148(.A(new_n563), .B1(new_n518), .B2(new_n519), .ZN(new_n574));
  XNOR2_X1  g149(.A(KEYINPUT72), .B(KEYINPUT9), .ZN(new_n575));
  NAND2_X1  g150(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  AOI21_X1  g151(.A(new_n566), .B1(new_n576), .B2(new_n565), .ZN(new_n577));
  OAI21_X1  g152(.A(new_n562), .B1(new_n573), .B2(new_n577), .ZN(G299));
  INV_X1    g153(.A(KEYINPUT74), .ZN(new_n579));
  NAND3_X1  g154(.A1(new_n530), .A2(new_n534), .A3(new_n579), .ZN(new_n580));
  AOI21_X1  g155(.A(new_n559), .B1(new_n531), .B2(new_n532), .ZN(new_n581));
  OAI21_X1  g156(.A(KEYINPUT74), .B1(new_n581), .B2(new_n529), .ZN(new_n582));
  NAND2_X1  g157(.A1(new_n580), .A2(new_n582), .ZN(new_n583));
  INV_X1    g158(.A(new_n583), .ZN(G286));
  INV_X1    g159(.A(G166), .ZN(G303));
  OAI21_X1  g160(.A(G651), .B1(new_n506), .B2(G74), .ZN(new_n586));
  NAND2_X1  g161(.A1(new_n511), .A2(new_n512), .ZN(new_n587));
  NAND3_X1  g162(.A1(new_n506), .A2(new_n587), .A3(G87), .ZN(new_n588));
  NAND3_X1  g163(.A1(new_n587), .A2(G49), .A3(G543), .ZN(new_n589));
  NAND3_X1  g164(.A1(new_n586), .A2(new_n588), .A3(new_n589), .ZN(G288));
  AOI22_X1  g165(.A1(new_n540), .A2(G86), .B1(new_n513), .B2(G48), .ZN(new_n591));
  OAI21_X1  g166(.A(G61), .B1(new_n517), .B2(new_n516), .ZN(new_n592));
  NAND2_X1  g167(.A1(G73), .A2(G543), .ZN(new_n593));
  AOI21_X1  g168(.A(new_n508), .B1(new_n592), .B2(new_n593), .ZN(new_n594));
  INV_X1    g169(.A(new_n594), .ZN(new_n595));
  NAND2_X1  g170(.A1(new_n591), .A2(new_n595), .ZN(G305));
  AOI22_X1  g171(.A1(new_n506), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n597));
  NOR2_X1   g172(.A1(new_n597), .A2(new_n508), .ZN(new_n598));
  NAND2_X1  g173(.A1(new_n513), .A2(G47), .ZN(new_n599));
  INV_X1    g174(.A(G85), .ZN(new_n600));
  OAI21_X1  g175(.A(new_n599), .B1(new_n600), .B2(new_n520), .ZN(new_n601));
  NOR2_X1   g176(.A1(new_n598), .A2(new_n601), .ZN(new_n602));
  INV_X1    g177(.A(new_n602), .ZN(G290));
  NAND2_X1  g178(.A1(G301), .A2(G868), .ZN(new_n604));
  NAND2_X1  g179(.A1(new_n513), .A2(G54), .ZN(new_n605));
  INV_X1    g180(.A(G79), .ZN(new_n606));
  NOR2_X1   g181(.A1(new_n606), .A2(new_n503), .ZN(new_n607));
  AOI21_X1  g182(.A(new_n607), .B1(new_n506), .B2(G66), .ZN(new_n608));
  OAI21_X1  g183(.A(new_n605), .B1(new_n608), .B2(new_n508), .ZN(new_n609));
  INV_X1    g184(.A(KEYINPUT10), .ZN(new_n610));
  INV_X1    g185(.A(G92), .ZN(new_n611));
  OAI21_X1  g186(.A(new_n610), .B1(new_n520), .B2(new_n611), .ZN(new_n612));
  NAND3_X1  g187(.A1(new_n540), .A2(KEYINPUT10), .A3(G92), .ZN(new_n613));
  AOI21_X1  g188(.A(new_n609), .B1(new_n612), .B2(new_n613), .ZN(new_n614));
  OAI21_X1  g189(.A(new_n604), .B1(new_n614), .B2(G868), .ZN(G284));
  OAI21_X1  g190(.A(new_n604), .B1(new_n614), .B2(G868), .ZN(G321));
  MUX2_X1   g191(.A(G299), .B(G286), .S(G868), .Z(G280));
  XOR2_X1   g192(.A(G280), .B(KEYINPUT75), .Z(G297));
  XOR2_X1   g193(.A(KEYINPUT76), .B(G559), .Z(new_n619));
  OAI21_X1  g194(.A(new_n614), .B1(G860), .B2(new_n619), .ZN(G148));
  INV_X1    g195(.A(G868), .ZN(new_n621));
  NAND2_X1  g196(.A1(new_n551), .A2(new_n621), .ZN(new_n622));
  AND2_X1   g197(.A1(new_n614), .A2(new_n619), .ZN(new_n623));
  OAI21_X1  g198(.A(new_n622), .B1(new_n623), .B2(new_n621), .ZN(G323));
  XNOR2_X1  g199(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g200(.A1(new_n464), .A2(new_n467), .ZN(new_n626));
  XNOR2_X1  g201(.A(new_n626), .B(KEYINPUT12), .ZN(new_n627));
  XNOR2_X1  g202(.A(new_n627), .B(KEYINPUT13), .ZN(new_n628));
  XNOR2_X1  g203(.A(new_n628), .B(G2100), .ZN(new_n629));
  NAND2_X1  g204(.A1(new_n481), .A2(G135), .ZN(new_n630));
  NAND2_X1  g205(.A1(new_n484), .A2(G123), .ZN(new_n631));
  OAI21_X1  g206(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n632));
  INV_X1    g207(.A(KEYINPUT78), .ZN(new_n633));
  OR2_X1    g208(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  NAND2_X1  g209(.A1(new_n632), .A2(new_n633), .ZN(new_n635));
  OR3_X1    g210(.A1(new_n465), .A2(KEYINPUT77), .A3(G111), .ZN(new_n636));
  OAI21_X1  g211(.A(KEYINPUT77), .B1(new_n465), .B2(G111), .ZN(new_n637));
  NAND4_X1  g212(.A1(new_n634), .A2(new_n635), .A3(new_n636), .A4(new_n637), .ZN(new_n638));
  NAND3_X1  g213(.A1(new_n630), .A2(new_n631), .A3(new_n638), .ZN(new_n639));
  OR2_X1    g214(.A1(new_n639), .A2(G2096), .ZN(new_n640));
  NAND2_X1  g215(.A1(new_n639), .A2(G2096), .ZN(new_n641));
  NAND3_X1  g216(.A1(new_n629), .A2(new_n640), .A3(new_n641), .ZN(G156));
  XNOR2_X1  g217(.A(G2427), .B(G2438), .ZN(new_n643));
  XNOR2_X1  g218(.A(new_n643), .B(G2430), .ZN(new_n644));
  XNOR2_X1  g219(.A(KEYINPUT15), .B(G2435), .ZN(new_n645));
  OR2_X1    g220(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  NAND2_X1  g221(.A1(new_n644), .A2(new_n645), .ZN(new_n647));
  NAND3_X1  g222(.A1(new_n646), .A2(KEYINPUT14), .A3(new_n647), .ZN(new_n648));
  XNOR2_X1  g223(.A(new_n648), .B(KEYINPUT79), .ZN(new_n649));
  XNOR2_X1  g224(.A(G2451), .B(G2454), .ZN(new_n650));
  XNOR2_X1  g225(.A(new_n650), .B(KEYINPUT16), .ZN(new_n651));
  XNOR2_X1  g226(.A(G2443), .B(G2446), .ZN(new_n652));
  XNOR2_X1  g227(.A(new_n651), .B(new_n652), .ZN(new_n653));
  XNOR2_X1  g228(.A(new_n649), .B(new_n653), .ZN(new_n654));
  XNOR2_X1  g229(.A(G1341), .B(G1348), .ZN(new_n655));
  OR2_X1    g230(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  NAND2_X1  g231(.A1(new_n654), .A2(new_n655), .ZN(new_n657));
  NAND3_X1  g232(.A1(new_n656), .A2(new_n657), .A3(G14), .ZN(new_n658));
  INV_X1    g233(.A(new_n658), .ZN(G401));
  XNOR2_X1  g234(.A(G2084), .B(G2090), .ZN(new_n660));
  XNOR2_X1  g235(.A(new_n660), .B(KEYINPUT80), .ZN(new_n661));
  XNOR2_X1  g236(.A(G2067), .B(G2678), .ZN(new_n662));
  NAND2_X1  g237(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  AND2_X1   g238(.A1(new_n663), .A2(KEYINPUT17), .ZN(new_n664));
  OR2_X1    g239(.A1(new_n661), .A2(new_n662), .ZN(new_n665));
  AOI21_X1  g240(.A(KEYINPUT18), .B1(new_n664), .B2(new_n665), .ZN(new_n666));
  XNOR2_X1  g241(.A(new_n666), .B(G2100), .ZN(new_n667));
  NOR2_X1   g242(.A1(G2072), .A2(G2078), .ZN(new_n668));
  NOR2_X1   g243(.A1(new_n444), .A2(new_n668), .ZN(new_n669));
  AOI21_X1  g244(.A(new_n669), .B1(new_n663), .B2(KEYINPUT18), .ZN(new_n670));
  XOR2_X1   g245(.A(new_n670), .B(G2096), .Z(new_n671));
  XNOR2_X1  g246(.A(new_n667), .B(new_n671), .ZN(G227));
  XOR2_X1   g247(.A(G1971), .B(G1976), .Z(new_n673));
  XNOR2_X1  g248(.A(new_n673), .B(KEYINPUT19), .ZN(new_n674));
  XOR2_X1   g249(.A(G1956), .B(G2474), .Z(new_n675));
  XOR2_X1   g250(.A(G1961), .B(G1966), .Z(new_n676));
  AND2_X1   g251(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  NAND2_X1  g252(.A1(new_n674), .A2(new_n677), .ZN(new_n678));
  XNOR2_X1  g253(.A(new_n678), .B(KEYINPUT20), .ZN(new_n679));
  NOR2_X1   g254(.A1(new_n675), .A2(new_n676), .ZN(new_n680));
  NOR3_X1   g255(.A1(new_n674), .A2(new_n677), .A3(new_n680), .ZN(new_n681));
  AOI21_X1  g256(.A(new_n681), .B1(new_n674), .B2(new_n680), .ZN(new_n682));
  NAND2_X1  g257(.A1(new_n679), .A2(new_n682), .ZN(new_n683));
  XNOR2_X1  g258(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n684));
  XOR2_X1   g259(.A(new_n684), .B(KEYINPUT81), .Z(new_n685));
  XNOR2_X1  g260(.A(new_n683), .B(new_n685), .ZN(new_n686));
  XNOR2_X1  g261(.A(G1991), .B(G1996), .ZN(new_n687));
  XNOR2_X1  g262(.A(new_n686), .B(new_n687), .ZN(new_n688));
  XNOR2_X1  g263(.A(G1981), .B(G1986), .ZN(new_n689));
  XNOR2_X1  g264(.A(new_n688), .B(new_n689), .ZN(G229));
  NOR2_X1   g265(.A1(G6), .A2(G16), .ZN(new_n691));
  INV_X1    g266(.A(G305), .ZN(new_n692));
  AOI21_X1  g267(.A(new_n691), .B1(new_n692), .B2(G16), .ZN(new_n693));
  XOR2_X1   g268(.A(KEYINPUT32), .B(G1981), .Z(new_n694));
  XNOR2_X1  g269(.A(new_n693), .B(new_n694), .ZN(new_n695));
  INV_X1    g270(.A(G16), .ZN(new_n696));
  NAND2_X1  g271(.A1(new_n696), .A2(G22), .ZN(new_n697));
  OAI21_X1  g272(.A(new_n697), .B1(G166), .B2(new_n696), .ZN(new_n698));
  INV_X1    g273(.A(G1971), .ZN(new_n699));
  XNOR2_X1  g274(.A(new_n698), .B(new_n699), .ZN(new_n700));
  NAND2_X1  g275(.A1(new_n696), .A2(G23), .ZN(new_n701));
  INV_X1    g276(.A(G288), .ZN(new_n702));
  OAI21_X1  g277(.A(new_n701), .B1(new_n702), .B2(new_n696), .ZN(new_n703));
  XNOR2_X1  g278(.A(KEYINPUT33), .B(G1976), .ZN(new_n704));
  XNOR2_X1  g279(.A(new_n703), .B(new_n704), .ZN(new_n705));
  NAND3_X1  g280(.A1(new_n695), .A2(new_n700), .A3(new_n705), .ZN(new_n706));
  XOR2_X1   g281(.A(new_n706), .B(KEYINPUT82), .Z(new_n707));
  INV_X1    g282(.A(KEYINPUT34), .ZN(new_n708));
  OR2_X1    g283(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  NAND2_X1  g284(.A1(new_n707), .A2(new_n708), .ZN(new_n710));
  NAND2_X1  g285(.A1(new_n481), .A2(G131), .ZN(new_n711));
  NAND2_X1  g286(.A1(new_n484), .A2(G119), .ZN(new_n712));
  OR2_X1    g287(.A1(G95), .A2(G2105), .ZN(new_n713));
  OAI211_X1 g288(.A(new_n713), .B(G2104), .C1(G107), .C2(new_n465), .ZN(new_n714));
  NAND3_X1  g289(.A1(new_n711), .A2(new_n712), .A3(new_n714), .ZN(new_n715));
  INV_X1    g290(.A(new_n715), .ZN(new_n716));
  NAND2_X1  g291(.A1(new_n716), .A2(G29), .ZN(new_n717));
  OAI21_X1  g292(.A(new_n717), .B1(G25), .B2(G29), .ZN(new_n718));
  XOR2_X1   g293(.A(KEYINPUT35), .B(G1991), .Z(new_n719));
  AND2_X1   g294(.A1(new_n718), .A2(new_n719), .ZN(new_n720));
  NOR2_X1   g295(.A1(new_n718), .A2(new_n719), .ZN(new_n721));
  NAND2_X1  g296(.A1(new_n696), .A2(G24), .ZN(new_n722));
  OAI21_X1  g297(.A(new_n722), .B1(new_n602), .B2(new_n696), .ZN(new_n723));
  XNOR2_X1  g298(.A(new_n723), .B(G1986), .ZN(new_n724));
  NOR3_X1   g299(.A1(new_n720), .A2(new_n721), .A3(new_n724), .ZN(new_n725));
  NAND3_X1  g300(.A1(new_n709), .A2(new_n710), .A3(new_n725), .ZN(new_n726));
  XNOR2_X1  g301(.A(new_n726), .B(KEYINPUT36), .ZN(new_n727));
  NAND2_X1  g302(.A1(new_n696), .A2(G4), .ZN(new_n728));
  OAI21_X1  g303(.A(new_n728), .B1(new_n614), .B2(new_n696), .ZN(new_n729));
  XNOR2_X1  g304(.A(new_n729), .B(KEYINPUT83), .ZN(new_n730));
  INV_X1    g305(.A(G1348), .ZN(new_n731));
  XNOR2_X1  g306(.A(new_n730), .B(new_n731), .ZN(new_n732));
  INV_X1    g307(.A(G29), .ZN(new_n733));
  INV_X1    g308(.A(KEYINPUT24), .ZN(new_n734));
  OAI21_X1  g309(.A(new_n733), .B1(new_n734), .B2(G34), .ZN(new_n735));
  OR2_X1    g310(.A1(new_n735), .A2(KEYINPUT88), .ZN(new_n736));
  NAND2_X1  g311(.A1(new_n735), .A2(KEYINPUT88), .ZN(new_n737));
  NAND2_X1  g312(.A1(new_n734), .A2(G34), .ZN(new_n738));
  NAND3_X1  g313(.A1(new_n736), .A2(new_n737), .A3(new_n738), .ZN(new_n739));
  XNOR2_X1  g314(.A(new_n739), .B(KEYINPUT89), .ZN(new_n740));
  AOI21_X1  g315(.A(new_n740), .B1(G29), .B2(G160), .ZN(new_n741));
  NAND2_X1  g316(.A1(new_n741), .A2(G2084), .ZN(new_n742));
  XOR2_X1   g317(.A(new_n742), .B(KEYINPUT90), .Z(new_n743));
  INV_X1    g318(.A(G1961), .ZN(new_n744));
  NAND2_X1  g319(.A1(new_n744), .A2(KEYINPUT93), .ZN(new_n745));
  NOR2_X1   g320(.A1(G171), .A2(new_n696), .ZN(new_n746));
  AND2_X1   g321(.A1(new_n696), .A2(G5), .ZN(new_n747));
  OAI21_X1  g322(.A(new_n745), .B1(new_n746), .B2(new_n747), .ZN(new_n748));
  NOR2_X1   g323(.A1(new_n744), .A2(KEYINPUT93), .ZN(new_n749));
  XOR2_X1   g324(.A(new_n748), .B(new_n749), .Z(new_n750));
  NAND2_X1  g325(.A1(new_n696), .A2(G21), .ZN(new_n751));
  OAI21_X1  g326(.A(new_n751), .B1(G168), .B2(new_n696), .ZN(new_n752));
  NAND2_X1  g327(.A1(new_n752), .A2(G1966), .ZN(new_n753));
  OAI221_X1 g328(.A(new_n753), .B1(new_n639), .B2(new_n733), .C1(new_n741), .C2(G2084), .ZN(new_n754));
  NOR4_X1   g329(.A1(new_n732), .A2(new_n743), .A3(new_n750), .A4(new_n754), .ZN(new_n755));
  NAND2_X1  g330(.A1(new_n696), .A2(G20), .ZN(new_n756));
  XOR2_X1   g331(.A(new_n756), .B(KEYINPUT23), .Z(new_n757));
  AOI21_X1  g332(.A(new_n757), .B1(G299), .B2(G16), .ZN(new_n758));
  XNOR2_X1  g333(.A(new_n758), .B(G1956), .ZN(new_n759));
  NAND2_X1  g334(.A1(new_n696), .A2(G19), .ZN(new_n760));
  OAI21_X1  g335(.A(new_n760), .B1(new_n552), .B2(new_n696), .ZN(new_n761));
  XOR2_X1   g336(.A(new_n761), .B(G1341), .Z(new_n762));
  INV_X1    g337(.A(G28), .ZN(new_n763));
  OR2_X1    g338(.A1(new_n763), .A2(KEYINPUT30), .ZN(new_n764));
  AOI21_X1  g339(.A(G29), .B1(new_n763), .B2(KEYINPUT30), .ZN(new_n765));
  OR2_X1    g340(.A1(KEYINPUT31), .A2(G11), .ZN(new_n766));
  NAND2_X1  g341(.A1(KEYINPUT31), .A2(G11), .ZN(new_n767));
  AOI22_X1  g342(.A1(new_n764), .A2(new_n765), .B1(new_n766), .B2(new_n767), .ZN(new_n768));
  OAI21_X1  g343(.A(new_n768), .B1(new_n752), .B2(G1966), .ZN(new_n769));
  NOR2_X1   g344(.A1(G27), .A2(G29), .ZN(new_n770));
  AOI21_X1  g345(.A(new_n770), .B1(G164), .B2(G29), .ZN(new_n771));
  XOR2_X1   g346(.A(KEYINPUT94), .B(G2078), .Z(new_n772));
  AND2_X1   g347(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  NOR2_X1   g348(.A1(new_n771), .A2(new_n772), .ZN(new_n774));
  NOR3_X1   g349(.A1(new_n769), .A2(new_n773), .A3(new_n774), .ZN(new_n775));
  NAND4_X1  g350(.A1(new_n755), .A2(new_n759), .A3(new_n762), .A4(new_n775), .ZN(new_n776));
  NAND2_X1  g351(.A1(new_n733), .A2(G35), .ZN(new_n777));
  OAI21_X1  g352(.A(new_n777), .B1(G162), .B2(new_n733), .ZN(new_n778));
  XOR2_X1   g353(.A(new_n778), .B(KEYINPUT29), .Z(new_n779));
  INV_X1    g354(.A(G2090), .ZN(new_n780));
  OR2_X1    g355(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  XOR2_X1   g356(.A(KEYINPUT85), .B(KEYINPUT28), .Z(new_n782));
  NAND2_X1  g357(.A1(new_n733), .A2(G26), .ZN(new_n783));
  XNOR2_X1  g358(.A(new_n782), .B(new_n783), .ZN(new_n784));
  OAI21_X1  g359(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n785));
  INV_X1    g360(.A(G116), .ZN(new_n786));
  AOI21_X1  g361(.A(new_n785), .B1(new_n786), .B2(G2105), .ZN(new_n787));
  AOI21_X1  g362(.A(new_n787), .B1(new_n484), .B2(G128), .ZN(new_n788));
  NAND2_X1  g363(.A1(new_n481), .A2(G140), .ZN(new_n789));
  AND2_X1   g364(.A1(new_n789), .A2(KEYINPUT84), .ZN(new_n790));
  NOR2_X1   g365(.A1(new_n789), .A2(KEYINPUT84), .ZN(new_n791));
  OAI21_X1  g366(.A(new_n788), .B1(new_n790), .B2(new_n791), .ZN(new_n792));
  INV_X1    g367(.A(new_n792), .ZN(new_n793));
  OAI21_X1  g368(.A(new_n784), .B1(new_n793), .B2(new_n733), .ZN(new_n794));
  INV_X1    g369(.A(G2067), .ZN(new_n795));
  XNOR2_X1  g370(.A(new_n794), .B(new_n795), .ZN(new_n796));
  NOR2_X1   g371(.A1(G29), .A2(G33), .ZN(new_n797));
  XOR2_X1   g372(.A(new_n797), .B(KEYINPUT86), .Z(new_n798));
  NAND3_X1  g373(.A1(new_n465), .A2(G103), .A3(G2104), .ZN(new_n799));
  XOR2_X1   g374(.A(new_n799), .B(KEYINPUT25), .Z(new_n800));
  AOI22_X1  g375(.A1(new_n464), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n801));
  INV_X1    g376(.A(G139), .ZN(new_n802));
  OAI221_X1 g377(.A(new_n800), .B1(new_n465), .B2(new_n801), .C1(new_n480), .C2(new_n802), .ZN(new_n803));
  INV_X1    g378(.A(KEYINPUT87), .ZN(new_n804));
  XNOR2_X1  g379(.A(new_n803), .B(new_n804), .ZN(new_n805));
  OAI21_X1  g380(.A(new_n798), .B1(new_n805), .B2(new_n733), .ZN(new_n806));
  XNOR2_X1  g381(.A(new_n806), .B(G2072), .ZN(new_n807));
  NAND2_X1  g382(.A1(new_n779), .A2(new_n780), .ZN(new_n808));
  NAND4_X1  g383(.A1(new_n781), .A2(new_n796), .A3(new_n807), .A4(new_n808), .ZN(new_n809));
  NAND3_X1  g384(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n810));
  INV_X1    g385(.A(KEYINPUT26), .ZN(new_n811));
  OR2_X1    g386(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  NAND2_X1  g387(.A1(new_n810), .A2(new_n811), .ZN(new_n813));
  AOI22_X1  g388(.A1(new_n812), .A2(new_n813), .B1(G105), .B2(new_n467), .ZN(new_n814));
  INV_X1    g389(.A(G141), .ZN(new_n815));
  INV_X1    g390(.A(G129), .ZN(new_n816));
  OAI221_X1 g391(.A(new_n814), .B1(new_n480), .B2(new_n815), .C1(new_n816), .C2(new_n483), .ZN(new_n817));
  NAND2_X1  g392(.A1(new_n817), .A2(KEYINPUT91), .ZN(new_n818));
  INV_X1    g393(.A(new_n818), .ZN(new_n819));
  NOR2_X1   g394(.A1(new_n817), .A2(KEYINPUT91), .ZN(new_n820));
  NOR2_X1   g395(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  NAND2_X1  g396(.A1(new_n821), .A2(G29), .ZN(new_n822));
  INV_X1    g397(.A(KEYINPUT92), .ZN(new_n823));
  OAI21_X1  g398(.A(new_n823), .B1(G29), .B2(G32), .ZN(new_n824));
  NAND2_X1  g399(.A1(new_n822), .A2(new_n824), .ZN(new_n825));
  OAI21_X1  g400(.A(new_n825), .B1(KEYINPUT92), .B2(new_n822), .ZN(new_n826));
  XNOR2_X1  g401(.A(KEYINPUT27), .B(G1996), .ZN(new_n827));
  XNOR2_X1  g402(.A(new_n826), .B(new_n827), .ZN(new_n828));
  NOR3_X1   g403(.A1(new_n776), .A2(new_n809), .A3(new_n828), .ZN(new_n829));
  NAND2_X1  g404(.A1(new_n727), .A2(new_n829), .ZN(G150));
  INV_X1    g405(.A(G150), .ZN(G311));
  NAND3_X1  g406(.A1(new_n506), .A2(new_n587), .A3(G93), .ZN(new_n832));
  NAND3_X1  g407(.A1(new_n587), .A2(G55), .A3(G543), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  OAI21_X1  g409(.A(G67), .B1(new_n517), .B2(new_n516), .ZN(new_n835));
  NAND2_X1  g410(.A1(G80), .A2(G543), .ZN(new_n836));
  AOI21_X1  g411(.A(new_n508), .B1(new_n835), .B2(new_n836), .ZN(new_n837));
  OAI21_X1  g412(.A(KEYINPUT95), .B1(new_n834), .B2(new_n837), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n835), .A2(new_n836), .ZN(new_n839));
  NAND2_X1  g414(.A1(new_n839), .A2(G651), .ZN(new_n840));
  INV_X1    g415(.A(KEYINPUT95), .ZN(new_n841));
  NAND4_X1  g416(.A1(new_n840), .A2(new_n841), .A3(new_n833), .A4(new_n832), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n838), .A2(new_n842), .ZN(new_n843));
  NAND2_X1  g418(.A1(new_n843), .A2(new_n551), .ZN(new_n844));
  AOI21_X1  g419(.A(new_n508), .B1(new_n545), .B2(new_n546), .ZN(new_n845));
  XNOR2_X1  g420(.A(new_n845), .B(KEYINPUT71), .ZN(new_n846));
  NAND4_X1  g421(.A1(new_n846), .A2(new_n544), .A3(new_n838), .A4(new_n842), .ZN(new_n847));
  NAND2_X1  g422(.A1(new_n844), .A2(new_n847), .ZN(new_n848));
  XOR2_X1   g423(.A(new_n848), .B(KEYINPUT38), .Z(new_n849));
  NAND2_X1  g424(.A1(new_n614), .A2(G559), .ZN(new_n850));
  XNOR2_X1  g425(.A(new_n849), .B(new_n850), .ZN(new_n851));
  OR2_X1    g426(.A1(new_n851), .A2(KEYINPUT39), .ZN(new_n852));
  INV_X1    g427(.A(G860), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n851), .A2(KEYINPUT39), .ZN(new_n854));
  NAND3_X1  g429(.A1(new_n852), .A2(new_n853), .A3(new_n854), .ZN(new_n855));
  NOR2_X1   g430(.A1(new_n834), .A2(new_n837), .ZN(new_n856));
  NOR2_X1   g431(.A1(new_n856), .A2(new_n853), .ZN(new_n857));
  XNOR2_X1  g432(.A(new_n857), .B(KEYINPUT37), .ZN(new_n858));
  NAND2_X1  g433(.A1(new_n855), .A2(new_n858), .ZN(G145));
  NAND2_X1  g434(.A1(new_n805), .A2(new_n792), .ZN(new_n860));
  INV_X1    g435(.A(new_n860), .ZN(new_n861));
  NOR2_X1   g436(.A1(new_n805), .A2(new_n792), .ZN(new_n862));
  OR2_X1    g437(.A1(G106), .A2(G2105), .ZN(new_n863));
  OAI211_X1 g438(.A(new_n863), .B(G2104), .C1(G118), .C2(new_n465), .ZN(new_n864));
  INV_X1    g439(.A(G142), .ZN(new_n865));
  INV_X1    g440(.A(G130), .ZN(new_n866));
  OAI221_X1 g441(.A(new_n864), .B1(new_n480), .B2(new_n865), .C1(new_n866), .C2(new_n483), .ZN(new_n867));
  XNOR2_X1  g442(.A(new_n867), .B(new_n627), .ZN(new_n868));
  NOR3_X1   g443(.A1(new_n861), .A2(new_n862), .A3(new_n868), .ZN(new_n869));
  INV_X1    g444(.A(new_n868), .ZN(new_n870));
  OR2_X1    g445(.A1(new_n805), .A2(new_n792), .ZN(new_n871));
  AOI21_X1  g446(.A(new_n870), .B1(new_n871), .B2(new_n860), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n498), .A2(new_n500), .ZN(new_n873));
  INV_X1    g448(.A(new_n493), .ZN(new_n874));
  NAND2_X1  g449(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  OAI21_X1  g450(.A(new_n875), .B1(new_n819), .B2(new_n820), .ZN(new_n876));
  INV_X1    g451(.A(new_n820), .ZN(new_n877));
  NAND3_X1  g452(.A1(new_n877), .A2(G164), .A3(new_n818), .ZN(new_n878));
  NAND3_X1  g453(.A1(new_n876), .A2(new_n878), .A3(new_n715), .ZN(new_n879));
  INV_X1    g454(.A(new_n879), .ZN(new_n880));
  AOI21_X1  g455(.A(new_n715), .B1(new_n876), .B2(new_n878), .ZN(new_n881));
  OAI22_X1  g456(.A1(new_n869), .A2(new_n872), .B1(new_n880), .B2(new_n881), .ZN(new_n882));
  INV_X1    g457(.A(new_n881), .ZN(new_n883));
  OAI21_X1  g458(.A(new_n868), .B1(new_n861), .B2(new_n862), .ZN(new_n884));
  NAND3_X1  g459(.A1(new_n871), .A2(new_n860), .A3(new_n870), .ZN(new_n885));
  NAND4_X1  g460(.A1(new_n883), .A2(new_n879), .A3(new_n884), .A4(new_n885), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n882), .A2(new_n886), .ZN(new_n887));
  INV_X1    g462(.A(new_n887), .ZN(new_n888));
  OAI21_X1  g463(.A(new_n488), .B1(new_n474), .B2(new_n469), .ZN(new_n889));
  INV_X1    g464(.A(KEYINPUT96), .ZN(new_n890));
  NAND4_X1  g465(.A1(new_n482), .A2(new_n485), .A3(G160), .A4(new_n487), .ZN(new_n891));
  AND3_X1   g466(.A1(new_n889), .A2(new_n890), .A3(new_n891), .ZN(new_n892));
  AOI21_X1  g467(.A(new_n890), .B1(new_n889), .B2(new_n891), .ZN(new_n893));
  OAI21_X1  g468(.A(new_n639), .B1(new_n892), .B2(new_n893), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n889), .A2(new_n891), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n895), .A2(KEYINPUT96), .ZN(new_n896));
  INV_X1    g471(.A(new_n639), .ZN(new_n897));
  NAND3_X1  g472(.A1(new_n889), .A2(new_n890), .A3(new_n891), .ZN(new_n898));
  NAND3_X1  g473(.A1(new_n896), .A2(new_n897), .A3(new_n898), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n894), .A2(new_n899), .ZN(new_n900));
  AOI21_X1  g475(.A(G37), .B1(new_n888), .B2(new_n900), .ZN(new_n901));
  INV_X1    g476(.A(KEYINPUT97), .ZN(new_n902));
  XNOR2_X1  g477(.A(new_n900), .B(new_n902), .ZN(new_n903));
  INV_X1    g478(.A(KEYINPUT98), .ZN(new_n904));
  AND3_X1   g479(.A1(new_n903), .A2(new_n904), .A3(new_n887), .ZN(new_n905));
  AOI21_X1  g480(.A(new_n904), .B1(new_n903), .B2(new_n887), .ZN(new_n906));
  OAI21_X1  g481(.A(new_n901), .B1(new_n905), .B2(new_n906), .ZN(new_n907));
  XNOR2_X1  g482(.A(KEYINPUT99), .B(KEYINPUT40), .ZN(new_n908));
  XNOR2_X1  g483(.A(new_n907), .B(new_n908), .ZN(G395));
  OAI21_X1  g484(.A(KEYINPUT100), .B1(new_n614), .B2(G299), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n614), .A2(G299), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n613), .A2(new_n612), .ZN(new_n912));
  INV_X1    g487(.A(G66), .ZN(new_n913));
  OAI22_X1  g488(.A1(new_n559), .A2(new_n913), .B1(new_n606), .B2(new_n503), .ZN(new_n914));
  AOI22_X1  g489(.A1(new_n914), .A2(G651), .B1(G54), .B2(new_n513), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n912), .A2(new_n915), .ZN(new_n916));
  INV_X1    g491(.A(KEYINPUT100), .ZN(new_n917));
  OAI21_X1  g492(.A(new_n565), .B1(new_n568), .B2(new_n571), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n918), .A2(KEYINPUT73), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n919), .A2(new_n572), .ZN(new_n920));
  NAND4_X1  g495(.A1(new_n916), .A2(new_n917), .A3(new_n562), .A4(new_n920), .ZN(new_n921));
  NAND3_X1  g496(.A1(new_n910), .A2(new_n911), .A3(new_n921), .ZN(new_n922));
  INV_X1    g497(.A(KEYINPUT41), .ZN(new_n923));
  AND3_X1   g498(.A1(new_n922), .A2(KEYINPUT101), .A3(new_n923), .ZN(new_n924));
  AOI21_X1  g499(.A(KEYINPUT101), .B1(new_n922), .B2(new_n923), .ZN(new_n925));
  AOI21_X1  g500(.A(new_n923), .B1(new_n614), .B2(G299), .ZN(new_n926));
  NAND3_X1  g501(.A1(new_n916), .A2(new_n562), .A3(new_n920), .ZN(new_n927));
  AND2_X1   g502(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  NOR3_X1   g503(.A1(new_n924), .A2(new_n925), .A3(new_n928), .ZN(new_n929));
  XOR2_X1   g504(.A(new_n848), .B(new_n623), .Z(new_n930));
  NOR2_X1   g505(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  INV_X1    g506(.A(KEYINPUT42), .ZN(new_n932));
  NOR2_X1   g507(.A1(new_n932), .A2(KEYINPUT102), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n911), .A2(new_n927), .ZN(new_n934));
  AND2_X1   g509(.A1(new_n930), .A2(new_n934), .ZN(new_n935));
  OR3_X1    g510(.A1(new_n931), .A2(new_n933), .A3(new_n935), .ZN(new_n936));
  NAND2_X1  g511(.A1(G303), .A2(new_n702), .ZN(new_n937));
  NAND2_X1  g512(.A1(G166), .A2(G288), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  NAND2_X1  g514(.A1(G290), .A2(new_n692), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n602), .A2(G305), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n939), .A2(new_n942), .ZN(new_n943));
  NAND4_X1  g518(.A1(new_n937), .A2(new_n940), .A3(new_n938), .A4(new_n941), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  INV_X1    g520(.A(new_n945), .ZN(new_n946));
  AOI21_X1  g521(.A(new_n946), .B1(KEYINPUT102), .B2(new_n932), .ZN(new_n947));
  OAI21_X1  g522(.A(new_n933), .B1(new_n931), .B2(new_n935), .ZN(new_n948));
  AND3_X1   g523(.A1(new_n936), .A2(new_n947), .A3(new_n948), .ZN(new_n949));
  AOI21_X1  g524(.A(new_n947), .B1(new_n936), .B2(new_n948), .ZN(new_n950));
  OAI21_X1  g525(.A(G868), .B1(new_n949), .B2(new_n950), .ZN(new_n951));
  OAI21_X1  g526(.A(new_n951), .B1(G868), .B2(new_n856), .ZN(G295));
  OAI21_X1  g527(.A(new_n951), .B1(G868), .B2(new_n856), .ZN(G331));
  AOI22_X1  g528(.A1(new_n539), .A2(new_n541), .B1(new_n534), .B2(new_n530), .ZN(new_n954));
  AOI21_X1  g529(.A(new_n954), .B1(G171), .B2(new_n583), .ZN(new_n955));
  NOR2_X1   g530(.A1(new_n843), .A2(new_n551), .ZN(new_n956));
  AOI22_X1  g531(.A1(new_n846), .A2(new_n544), .B1(new_n838), .B2(new_n842), .ZN(new_n957));
  OAI21_X1  g532(.A(new_n955), .B1(new_n956), .B2(new_n957), .ZN(new_n958));
  AOI21_X1  g533(.A(G301), .B1(new_n582), .B2(new_n580), .ZN(new_n959));
  OAI211_X1 g534(.A(new_n844), .B(new_n847), .C1(new_n959), .C2(new_n954), .ZN(new_n960));
  NAND2_X1  g535(.A1(new_n958), .A2(new_n960), .ZN(new_n961));
  NAND2_X1  g536(.A1(new_n961), .A2(new_n934), .ZN(new_n962));
  OAI211_X1 g537(.A(new_n945), .B(new_n962), .C1(new_n929), .C2(new_n961), .ZN(new_n963));
  AND3_X1   g538(.A1(new_n910), .A2(new_n926), .A3(new_n921), .ZN(new_n964));
  AOI21_X1  g539(.A(KEYINPUT41), .B1(new_n911), .B2(new_n927), .ZN(new_n965));
  OAI211_X1 g540(.A(new_n960), .B(new_n958), .C1(new_n964), .C2(new_n965), .ZN(new_n966));
  NAND3_X1  g541(.A1(new_n966), .A2(new_n962), .A3(KEYINPUT103), .ZN(new_n967));
  AOI22_X1  g542(.A1(new_n958), .A2(new_n960), .B1(new_n911), .B2(new_n927), .ZN(new_n968));
  INV_X1    g543(.A(KEYINPUT103), .ZN(new_n969));
  AOI21_X1  g544(.A(new_n945), .B1(new_n968), .B2(new_n969), .ZN(new_n970));
  AOI21_X1  g545(.A(G37), .B1(new_n967), .B2(new_n970), .ZN(new_n971));
  INV_X1    g546(.A(KEYINPUT43), .ZN(new_n972));
  AND3_X1   g547(.A1(new_n963), .A2(new_n971), .A3(new_n972), .ZN(new_n973));
  INV_X1    g548(.A(KEYINPUT104), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n922), .A2(new_n923), .ZN(new_n975));
  INV_X1    g550(.A(KEYINPUT101), .ZN(new_n976));
  AOI21_X1  g551(.A(new_n928), .B1(new_n975), .B2(new_n976), .ZN(new_n977));
  NAND3_X1  g552(.A1(new_n922), .A2(KEYINPUT101), .A3(new_n923), .ZN(new_n978));
  AOI21_X1  g553(.A(new_n961), .B1(new_n977), .B2(new_n978), .ZN(new_n979));
  OAI21_X1  g554(.A(new_n946), .B1(new_n979), .B2(new_n968), .ZN(new_n980));
  INV_X1    g555(.A(G37), .ZN(new_n981));
  NAND3_X1  g556(.A1(new_n980), .A2(new_n963), .A3(new_n981), .ZN(new_n982));
  AOI22_X1  g557(.A1(new_n973), .A2(new_n974), .B1(new_n982), .B2(KEYINPUT43), .ZN(new_n983));
  NAND3_X1  g558(.A1(new_n963), .A2(new_n971), .A3(new_n972), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n984), .A2(KEYINPUT104), .ZN(new_n985));
  AOI21_X1  g560(.A(KEYINPUT44), .B1(new_n983), .B2(new_n985), .ZN(new_n986));
  INV_X1    g561(.A(KEYINPUT44), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n982), .A2(new_n972), .ZN(new_n988));
  NAND3_X1  g563(.A1(new_n963), .A2(new_n971), .A3(KEYINPUT43), .ZN(new_n989));
  AOI21_X1  g564(.A(new_n987), .B1(new_n988), .B2(new_n989), .ZN(new_n990));
  OAI21_X1  g565(.A(KEYINPUT105), .B1(new_n986), .B2(new_n990), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n982), .A2(KEYINPUT43), .ZN(new_n992));
  NAND4_X1  g567(.A1(new_n963), .A2(new_n971), .A3(new_n974), .A4(new_n972), .ZN(new_n993));
  NAND3_X1  g568(.A1(new_n992), .A2(new_n985), .A3(new_n993), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n994), .A2(new_n987), .ZN(new_n995));
  INV_X1    g570(.A(new_n990), .ZN(new_n996));
  INV_X1    g571(.A(KEYINPUT105), .ZN(new_n997));
  NAND3_X1  g572(.A1(new_n995), .A2(new_n996), .A3(new_n997), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n991), .A2(new_n998), .ZN(G397));
  INV_X1    g574(.A(KEYINPUT119), .ZN(new_n1000));
  NOR2_X1   g575(.A1(new_n1000), .A2(KEYINPUT59), .ZN(new_n1001));
  AOI21_X1  g576(.A(G1384), .B1(new_n873), .B2(new_n874), .ZN(new_n1002));
  INV_X1    g577(.A(G40), .ZN(new_n1003));
  NOR3_X1   g578(.A1(new_n469), .A2(new_n474), .A3(new_n1003), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n1002), .A2(new_n1004), .ZN(new_n1005));
  XOR2_X1   g580(.A(KEYINPUT58), .B(G1341), .Z(new_n1006));
  NAND2_X1  g581(.A1(new_n1005), .A2(new_n1006), .ZN(new_n1007));
  INV_X1    g582(.A(new_n1007), .ZN(new_n1008));
  INV_X1    g583(.A(G1996), .ZN(new_n1009));
  INV_X1    g584(.A(new_n474), .ZN(new_n1010));
  NAND4_X1  g585(.A1(new_n1010), .A2(G40), .A3(new_n468), .A4(new_n466), .ZN(new_n1011));
  AOI21_X1  g586(.A(new_n1011), .B1(new_n1002), .B2(KEYINPUT45), .ZN(new_n1012));
  INV_X1    g587(.A(KEYINPUT107), .ZN(new_n1013));
  INV_X1    g588(.A(G1384), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n875), .A2(new_n1014), .ZN(new_n1015));
  INV_X1    g590(.A(KEYINPUT45), .ZN(new_n1016));
  AOI21_X1  g591(.A(new_n1013), .B1(new_n1015), .B2(new_n1016), .ZN(new_n1017));
  OAI211_X1 g592(.A(new_n1013), .B(new_n1016), .C1(G164), .C2(G1384), .ZN(new_n1018));
  INV_X1    g593(.A(new_n1018), .ZN(new_n1019));
  OAI211_X1 g594(.A(new_n1009), .B(new_n1012), .C1(new_n1017), .C2(new_n1019), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n1020), .A2(KEYINPUT117), .ZN(new_n1021));
  OAI21_X1  g596(.A(new_n1016), .B1(G164), .B2(G1384), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n1022), .A2(KEYINPUT107), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n1023), .A2(new_n1018), .ZN(new_n1024));
  INV_X1    g599(.A(KEYINPUT117), .ZN(new_n1025));
  NAND4_X1  g600(.A1(new_n1024), .A2(new_n1025), .A3(new_n1009), .A4(new_n1012), .ZN(new_n1026));
  AOI21_X1  g601(.A(new_n1008), .B1(new_n1021), .B2(new_n1026), .ZN(new_n1027));
  OAI21_X1  g602(.A(new_n552), .B1(new_n1027), .B2(KEYINPUT118), .ZN(new_n1028));
  INV_X1    g603(.A(KEYINPUT118), .ZN(new_n1029));
  AOI211_X1 g604(.A(new_n1029), .B(new_n1008), .C1(new_n1021), .C2(new_n1026), .ZN(new_n1030));
  OAI21_X1  g605(.A(new_n1001), .B1(new_n1028), .B2(new_n1030), .ZN(new_n1031));
  XNOR2_X1  g606(.A(KEYINPUT56), .B(G2072), .ZN(new_n1032));
  OAI211_X1 g607(.A(new_n1012), .B(new_n1032), .C1(new_n1017), .C2(new_n1019), .ZN(new_n1033));
  OAI211_X1 g608(.A(new_n562), .B(KEYINPUT57), .C1(new_n573), .C2(new_n577), .ZN(new_n1034));
  NOR2_X1   g609(.A1(new_n1034), .A2(KEYINPUT116), .ZN(new_n1035));
  AND2_X1   g610(.A1(new_n1034), .A2(KEYINPUT116), .ZN(new_n1036));
  INV_X1    g611(.A(KEYINPUT115), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n918), .A2(new_n1037), .ZN(new_n1038));
  NAND3_X1  g613(.A1(new_n576), .A2(KEYINPUT115), .A3(new_n565), .ZN(new_n1039));
  NAND3_X1  g614(.A1(new_n562), .A2(new_n1038), .A3(new_n1039), .ZN(new_n1040));
  INV_X1    g615(.A(KEYINPUT57), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n1040), .A2(new_n1041), .ZN(new_n1042));
  AOI21_X1  g617(.A(new_n1035), .B1(new_n1036), .B2(new_n1042), .ZN(new_n1043));
  INV_X1    g618(.A(KEYINPUT50), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n1002), .A2(new_n1044), .ZN(new_n1045));
  XOR2_X1   g620(.A(KEYINPUT108), .B(KEYINPUT50), .Z(new_n1046));
  INV_X1    g621(.A(new_n1046), .ZN(new_n1047));
  OAI21_X1  g622(.A(new_n1047), .B1(G164), .B2(G1384), .ZN(new_n1048));
  NAND3_X1  g623(.A1(new_n1045), .A2(new_n1004), .A3(new_n1048), .ZN(new_n1049));
  INV_X1    g624(.A(G1956), .ZN(new_n1050));
  NAND2_X1  g625(.A1(new_n1049), .A2(new_n1050), .ZN(new_n1051));
  NAND3_X1  g626(.A1(new_n1033), .A2(new_n1043), .A3(new_n1051), .ZN(new_n1052));
  INV_X1    g627(.A(KEYINPUT120), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n1053), .A2(KEYINPUT61), .ZN(new_n1054));
  NAND2_X1  g629(.A1(new_n1052), .A2(new_n1054), .ZN(new_n1055));
  NAND4_X1  g630(.A1(new_n1033), .A2(new_n1043), .A3(new_n1053), .A4(new_n1051), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n1033), .A2(new_n1051), .ZN(new_n1057));
  INV_X1    g632(.A(new_n1043), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n1057), .A2(new_n1058), .ZN(new_n1059));
  NAND3_X1  g634(.A1(new_n1055), .A2(new_n1056), .A3(new_n1059), .ZN(new_n1060));
  AOI21_X1  g635(.A(new_n1011), .B1(new_n1002), .B2(new_n1046), .ZN(new_n1061));
  OAI21_X1  g636(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n1062));
  AOI21_X1  g637(.A(G1348), .B1(new_n1061), .B2(new_n1062), .ZN(new_n1063));
  NAND3_X1  g638(.A1(new_n1002), .A2(new_n795), .A3(new_n1004), .ZN(new_n1064));
  INV_X1    g639(.A(new_n1064), .ZN(new_n1065));
  OAI21_X1  g640(.A(new_n614), .B1(new_n1063), .B2(new_n1065), .ZN(new_n1066));
  NAND3_X1  g641(.A1(new_n875), .A2(new_n1014), .A3(new_n1046), .ZN(new_n1067));
  NAND3_X1  g642(.A1(new_n1067), .A2(new_n1062), .A3(new_n1004), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n1068), .A2(new_n731), .ZN(new_n1069));
  NAND3_X1  g644(.A1(new_n1069), .A2(new_n916), .A3(new_n1064), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n1066), .A2(new_n1070), .ZN(new_n1071));
  NOR2_X1   g646(.A1(new_n1063), .A2(new_n1065), .ZN(new_n1072));
  NOR2_X1   g647(.A1(new_n916), .A2(KEYINPUT60), .ZN(new_n1073));
  AOI22_X1  g648(.A1(new_n1071), .A2(KEYINPUT60), .B1(new_n1072), .B2(new_n1073), .ZN(new_n1074));
  INV_X1    g649(.A(KEYINPUT61), .ZN(new_n1075));
  AND3_X1   g650(.A1(new_n1033), .A2(new_n1043), .A3(new_n1051), .ZN(new_n1076));
  AOI21_X1  g651(.A(new_n1043), .B1(new_n1033), .B2(new_n1051), .ZN(new_n1077));
  OAI21_X1  g652(.A(new_n1075), .B1(new_n1076), .B2(new_n1077), .ZN(new_n1078));
  AND3_X1   g653(.A1(new_n1060), .A2(new_n1074), .A3(new_n1078), .ZN(new_n1079));
  NAND3_X1  g654(.A1(new_n875), .A2(KEYINPUT45), .A3(new_n1014), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1080), .A2(new_n1004), .ZN(new_n1081));
  AOI21_X1  g656(.A(new_n1081), .B1(new_n1023), .B2(new_n1018), .ZN(new_n1082));
  AOI21_X1  g657(.A(new_n1025), .B1(new_n1082), .B2(new_n1009), .ZN(new_n1083));
  INV_X1    g658(.A(new_n1026), .ZN(new_n1084));
  OAI21_X1  g659(.A(new_n1007), .B1(new_n1083), .B2(new_n1084), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n1085), .A2(new_n1029), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n1027), .A2(KEYINPUT118), .ZN(new_n1087));
  XNOR2_X1  g662(.A(KEYINPUT119), .B(KEYINPUT59), .ZN(new_n1088));
  NAND4_X1  g663(.A1(new_n1086), .A2(new_n552), .A3(new_n1087), .A4(new_n1088), .ZN(new_n1089));
  NAND3_X1  g664(.A1(new_n1031), .A2(new_n1079), .A3(new_n1089), .ZN(new_n1090));
  INV_X1    g665(.A(new_n1066), .ZN(new_n1091));
  OAI21_X1  g666(.A(new_n1052), .B1(new_n1077), .B2(new_n1091), .ZN(new_n1092));
  NAND2_X1  g667(.A1(new_n1090), .A2(new_n1092), .ZN(new_n1093));
  INV_X1    g668(.A(new_n1022), .ZN(new_n1094));
  NOR2_X1   g669(.A1(new_n1081), .A2(new_n1094), .ZN(new_n1095));
  INV_X1    g670(.A(KEYINPUT53), .ZN(new_n1096));
  NOR2_X1   g671(.A1(new_n1096), .A2(G2078), .ZN(new_n1097));
  MUX2_X1   g672(.A(G2078), .B(new_n1097), .S(KEYINPUT124), .Z(new_n1098));
  NAND2_X1  g673(.A1(new_n1095), .A2(new_n1098), .ZN(new_n1099));
  AND3_X1   g674(.A1(new_n1068), .A2(KEYINPUT123), .A3(new_n744), .ZN(new_n1100));
  AOI21_X1  g675(.A(KEYINPUT123), .B1(new_n1068), .B2(new_n744), .ZN(new_n1101));
  OAI21_X1  g676(.A(new_n1099), .B1(new_n1100), .B2(new_n1101), .ZN(new_n1102));
  INV_X1    g677(.A(G2078), .ZN(new_n1103));
  AOI21_X1  g678(.A(KEYINPUT53), .B1(new_n1082), .B2(new_n1103), .ZN(new_n1104));
  OAI21_X1  g679(.A(G171), .B1(new_n1102), .B2(new_n1104), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n1024), .A2(new_n1012), .ZN(new_n1106));
  OAI21_X1  g681(.A(new_n1096), .B1(new_n1106), .B2(G2078), .ZN(new_n1107));
  AOI22_X1  g682(.A1(new_n1095), .A2(new_n1097), .B1(new_n744), .B2(new_n1068), .ZN(new_n1108));
  NAND3_X1  g683(.A1(new_n1107), .A2(G301), .A3(new_n1108), .ZN(new_n1109));
  NAND3_X1  g684(.A1(new_n1105), .A2(KEYINPUT54), .A3(new_n1109), .ZN(new_n1110));
  INV_X1    g685(.A(G8), .ZN(new_n1111));
  NOR2_X1   g686(.A1(G166), .A2(new_n1111), .ZN(new_n1112));
  XNOR2_X1  g687(.A(KEYINPUT109), .B(KEYINPUT55), .ZN(new_n1113));
  OR2_X1    g688(.A1(new_n1112), .A2(new_n1113), .ZN(new_n1114));
  INV_X1    g689(.A(KEYINPUT109), .ZN(new_n1115));
  OAI21_X1  g690(.A(new_n1112), .B1(new_n1115), .B2(KEYINPUT55), .ZN(new_n1116));
  NAND2_X1  g691(.A1(new_n1114), .A2(new_n1116), .ZN(new_n1117));
  INV_X1    g692(.A(new_n1117), .ZN(new_n1118));
  AND4_X1   g693(.A1(new_n780), .A2(new_n1045), .A3(new_n1004), .A4(new_n1048), .ZN(new_n1119));
  AOI21_X1  g694(.A(new_n1119), .B1(new_n1106), .B2(new_n699), .ZN(new_n1120));
  OAI21_X1  g695(.A(new_n1118), .B1(new_n1120), .B2(new_n1111), .ZN(new_n1121));
  INV_X1    g696(.A(KEYINPUT112), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n1121), .A2(new_n1122), .ZN(new_n1123));
  AOI21_X1  g698(.A(G1971), .B1(new_n1024), .B2(new_n1012), .ZN(new_n1124));
  NOR2_X1   g699(.A1(new_n1068), .A2(G2090), .ZN(new_n1125));
  OAI211_X1 g700(.A(G8), .B(new_n1117), .C1(new_n1124), .C2(new_n1125), .ZN(new_n1126));
  AND4_X1   g701(.A1(G1976), .A2(new_n586), .A3(new_n588), .A4(new_n589), .ZN(new_n1127));
  INV_X1    g702(.A(new_n1127), .ZN(new_n1128));
  INV_X1    g703(.A(G1976), .ZN(new_n1129));
  AOI21_X1  g704(.A(KEYINPUT52), .B1(G288), .B2(new_n1129), .ZN(new_n1130));
  NAND4_X1  g705(.A1(new_n1005), .A2(G8), .A3(new_n1128), .A4(new_n1130), .ZN(new_n1131));
  AOI211_X1 g706(.A(new_n1111), .B(new_n1127), .C1(new_n1002), .C2(new_n1004), .ZN(new_n1132));
  INV_X1    g707(.A(KEYINPUT52), .ZN(new_n1133));
  OAI21_X1  g708(.A(new_n1131), .B1(new_n1132), .B2(new_n1133), .ZN(new_n1134));
  INV_X1    g709(.A(G1981), .ZN(new_n1135));
  AOI21_X1  g710(.A(new_n1135), .B1(new_n591), .B2(new_n595), .ZN(new_n1136));
  INV_X1    g711(.A(new_n1136), .ZN(new_n1137));
  NAND3_X1  g712(.A1(new_n591), .A2(new_n595), .A3(new_n1135), .ZN(new_n1138));
  NAND3_X1  g713(.A1(new_n1137), .A2(new_n1138), .A3(KEYINPUT49), .ZN(new_n1139));
  INV_X1    g714(.A(KEYINPUT49), .ZN(new_n1140));
  AND3_X1   g715(.A1(new_n591), .A2(new_n595), .A3(new_n1135), .ZN(new_n1141));
  OAI21_X1  g716(.A(new_n1140), .B1(new_n1141), .B2(new_n1136), .ZN(new_n1142));
  AOI21_X1  g717(.A(new_n1111), .B1(new_n1002), .B2(new_n1004), .ZN(new_n1143));
  NAND3_X1  g718(.A1(new_n1139), .A2(new_n1142), .A3(new_n1143), .ZN(new_n1144));
  NAND2_X1  g719(.A1(new_n1144), .A2(KEYINPUT110), .ZN(new_n1145));
  INV_X1    g720(.A(KEYINPUT110), .ZN(new_n1146));
  NAND4_X1  g721(.A1(new_n1139), .A2(new_n1142), .A3(new_n1143), .A4(new_n1146), .ZN(new_n1147));
  AOI21_X1  g722(.A(new_n1134), .B1(new_n1145), .B2(new_n1147), .ZN(new_n1148));
  AND2_X1   g723(.A1(new_n1126), .A2(new_n1148), .ZN(new_n1149));
  OAI211_X1 g724(.A(KEYINPUT112), .B(new_n1118), .C1(new_n1120), .C2(new_n1111), .ZN(new_n1150));
  NAND4_X1  g725(.A1(new_n1110), .A2(new_n1123), .A3(new_n1149), .A4(new_n1150), .ZN(new_n1151));
  INV_X1    g726(.A(KEYINPUT113), .ZN(new_n1152));
  OAI21_X1  g727(.A(new_n1152), .B1(new_n1068), .B2(G2084), .ZN(new_n1153));
  INV_X1    g728(.A(G1966), .ZN(new_n1154));
  OAI21_X1  g729(.A(new_n1154), .B1(new_n1081), .B2(new_n1094), .ZN(new_n1155));
  INV_X1    g730(.A(G2084), .ZN(new_n1156));
  NAND4_X1  g731(.A1(new_n1061), .A2(KEYINPUT113), .A3(new_n1156), .A4(new_n1062), .ZN(new_n1157));
  NAND4_X1  g732(.A1(new_n1153), .A2(new_n1155), .A3(G168), .A4(new_n1157), .ZN(new_n1158));
  NAND2_X1  g733(.A1(KEYINPUT121), .A2(KEYINPUT51), .ZN(new_n1159));
  OR2_X1    g734(.A1(KEYINPUT121), .A2(KEYINPUT51), .ZN(new_n1160));
  AND4_X1   g735(.A1(G8), .A2(new_n1158), .A3(new_n1159), .A4(new_n1160), .ZN(new_n1161));
  NAND3_X1  g736(.A1(new_n1153), .A2(new_n1155), .A3(new_n1157), .ZN(new_n1162));
  AND3_X1   g737(.A1(new_n1162), .A2(G8), .A3(new_n535), .ZN(new_n1163));
  AOI21_X1  g738(.A(new_n1159), .B1(new_n1158), .B2(G8), .ZN(new_n1164));
  NOR3_X1   g739(.A1(new_n1161), .A2(new_n1163), .A3(new_n1164), .ZN(new_n1165));
  XOR2_X1   g740(.A(KEYINPUT122), .B(KEYINPUT54), .Z(new_n1166));
  OR3_X1    g741(.A1(new_n1102), .A2(new_n1104), .A3(G171), .ZN(new_n1167));
  NAND2_X1  g742(.A1(new_n1107), .A2(new_n1108), .ZN(new_n1168));
  NAND2_X1  g743(.A1(new_n1168), .A2(G171), .ZN(new_n1169));
  AOI21_X1  g744(.A(new_n1166), .B1(new_n1167), .B2(new_n1169), .ZN(new_n1170));
  NOR3_X1   g745(.A1(new_n1151), .A2(new_n1165), .A3(new_n1170), .ZN(new_n1171));
  NAND2_X1  g746(.A1(new_n1093), .A2(new_n1171), .ZN(new_n1172));
  AND3_X1   g747(.A1(new_n1162), .A2(G8), .A3(new_n583), .ZN(new_n1173));
  NAND4_X1  g748(.A1(new_n1123), .A2(new_n1149), .A3(new_n1150), .A4(new_n1173), .ZN(new_n1174));
  INV_X1    g749(.A(KEYINPUT63), .ZN(new_n1175));
  NAND2_X1  g750(.A1(new_n1174), .A2(new_n1175), .ZN(new_n1176));
  NAND2_X1  g751(.A1(new_n1126), .A2(new_n1148), .ZN(new_n1177));
  OAI22_X1  g752(.A1(new_n1082), .A2(G1971), .B1(G2090), .B2(new_n1068), .ZN(new_n1178));
  AOI21_X1  g753(.A(new_n1117), .B1(new_n1178), .B2(G8), .ZN(new_n1179));
  NOR3_X1   g754(.A1(new_n1177), .A2(new_n1179), .A3(new_n1175), .ZN(new_n1180));
  NAND2_X1  g755(.A1(new_n1180), .A2(new_n1173), .ZN(new_n1181));
  NAND2_X1  g756(.A1(new_n1176), .A2(new_n1181), .ZN(new_n1182));
  INV_X1    g757(.A(KEYINPUT114), .ZN(new_n1183));
  XNOR2_X1  g758(.A(new_n1143), .B(KEYINPUT111), .ZN(new_n1184));
  NAND2_X1  g759(.A1(new_n1145), .A2(new_n1147), .ZN(new_n1185));
  NOR2_X1   g760(.A1(G288), .A2(G1976), .ZN(new_n1186));
  NAND2_X1  g761(.A1(new_n1185), .A2(new_n1186), .ZN(new_n1187));
  AOI21_X1  g762(.A(new_n1184), .B1(new_n1187), .B2(new_n1138), .ZN(new_n1188));
  INV_X1    g763(.A(new_n1148), .ZN(new_n1189));
  NOR2_X1   g764(.A1(new_n1189), .A2(new_n1126), .ZN(new_n1190));
  NOR2_X1   g765(.A1(new_n1188), .A2(new_n1190), .ZN(new_n1191));
  NAND3_X1  g766(.A1(new_n1182), .A2(new_n1183), .A3(new_n1191), .ZN(new_n1192));
  AOI22_X1  g767(.A1(new_n1174), .A2(new_n1175), .B1(new_n1180), .B2(new_n1173), .ZN(new_n1193));
  INV_X1    g768(.A(new_n1191), .ZN(new_n1194));
  OAI21_X1  g769(.A(KEYINPUT114), .B1(new_n1193), .B2(new_n1194), .ZN(new_n1195));
  INV_X1    g770(.A(KEYINPUT62), .ZN(new_n1196));
  OR2_X1    g771(.A1(new_n1165), .A2(new_n1196), .ZN(new_n1197));
  NAND2_X1  g772(.A1(new_n1165), .A2(new_n1196), .ZN(new_n1198));
  INV_X1    g773(.A(new_n1169), .ZN(new_n1199));
  AND3_X1   g774(.A1(new_n1123), .A2(new_n1149), .A3(new_n1150), .ZN(new_n1200));
  NAND4_X1  g775(.A1(new_n1197), .A2(new_n1198), .A3(new_n1199), .A4(new_n1200), .ZN(new_n1201));
  NAND4_X1  g776(.A1(new_n1172), .A2(new_n1192), .A3(new_n1195), .A4(new_n1201), .ZN(new_n1202));
  NAND2_X1  g777(.A1(new_n1094), .A2(new_n1004), .ZN(new_n1203));
  INV_X1    g778(.A(new_n1203), .ZN(new_n1204));
  XNOR2_X1  g779(.A(new_n792), .B(new_n795), .ZN(new_n1205));
  NAND2_X1  g780(.A1(new_n821), .A2(new_n1009), .ZN(new_n1206));
  OAI21_X1  g781(.A(G1996), .B1(new_n819), .B2(new_n820), .ZN(new_n1207));
  XNOR2_X1  g782(.A(new_n715), .B(new_n719), .ZN(new_n1208));
  NAND4_X1  g783(.A1(new_n1205), .A2(new_n1206), .A3(new_n1207), .A4(new_n1208), .ZN(new_n1209));
  OR2_X1    g784(.A1(G290), .A2(G1986), .ZN(new_n1210));
  INV_X1    g785(.A(KEYINPUT106), .ZN(new_n1211));
  NAND2_X1  g786(.A1(new_n1210), .A2(new_n1211), .ZN(new_n1212));
  NAND2_X1  g787(.A1(G290), .A2(G1986), .ZN(new_n1213));
  XNOR2_X1  g788(.A(new_n1212), .B(new_n1213), .ZN(new_n1214));
  OAI21_X1  g789(.A(new_n1204), .B1(new_n1209), .B2(new_n1214), .ZN(new_n1215));
  NAND2_X1  g790(.A1(new_n1202), .A2(new_n1215), .ZN(new_n1216));
  NOR2_X1   g791(.A1(new_n1210), .A2(new_n1203), .ZN(new_n1217));
  XNOR2_X1  g792(.A(new_n1217), .B(KEYINPUT127), .ZN(new_n1218));
  XOR2_X1   g793(.A(new_n1218), .B(KEYINPUT48), .Z(new_n1219));
  NAND3_X1  g794(.A1(new_n1209), .A2(KEYINPUT126), .A3(new_n1204), .ZN(new_n1220));
  NAND2_X1  g795(.A1(new_n1219), .A2(new_n1220), .ZN(new_n1221));
  AOI21_X1  g796(.A(KEYINPUT126), .B1(new_n1209), .B2(new_n1204), .ZN(new_n1222));
  INV_X1    g797(.A(KEYINPUT47), .ZN(new_n1223));
  NAND2_X1  g798(.A1(new_n1205), .A2(new_n821), .ZN(new_n1224));
  NAND2_X1  g799(.A1(new_n1224), .A2(new_n1204), .ZN(new_n1225));
  NAND2_X1  g800(.A1(new_n1204), .A2(new_n1009), .ZN(new_n1226));
  XNOR2_X1  g801(.A(new_n1226), .B(KEYINPUT46), .ZN(new_n1227));
  AOI21_X1  g802(.A(new_n1223), .B1(new_n1225), .B2(new_n1227), .ZN(new_n1228));
  AND3_X1   g803(.A1(new_n1225), .A2(new_n1223), .A3(new_n1227), .ZN(new_n1229));
  OAI22_X1  g804(.A1(new_n1221), .A2(new_n1222), .B1(new_n1228), .B2(new_n1229), .ZN(new_n1230));
  NAND3_X1  g805(.A1(new_n1205), .A2(new_n1206), .A3(new_n1207), .ZN(new_n1231));
  NAND2_X1  g806(.A1(new_n1231), .A2(new_n1204), .ZN(new_n1232));
  AND2_X1   g807(.A1(new_n716), .A2(new_n719), .ZN(new_n1233));
  AOI22_X1  g808(.A1(new_n1232), .A2(new_n1233), .B1(new_n795), .B2(new_n793), .ZN(new_n1234));
  INV_X1    g809(.A(KEYINPUT125), .ZN(new_n1235));
  OR2_X1    g810(.A1(new_n1234), .A2(new_n1235), .ZN(new_n1236));
  AOI21_X1  g811(.A(new_n1203), .B1(new_n1234), .B2(new_n1235), .ZN(new_n1237));
  AOI21_X1  g812(.A(new_n1230), .B1(new_n1236), .B2(new_n1237), .ZN(new_n1238));
  NAND2_X1  g813(.A1(new_n1216), .A2(new_n1238), .ZN(G329));
  assign    G231 = 1'b0;
  NOR4_X1   g814(.A1(G229), .A2(new_n462), .A3(G401), .A4(G227), .ZN(new_n1241));
  NAND3_X1  g815(.A1(new_n907), .A2(new_n1241), .A3(new_n994), .ZN(G225));
  INV_X1    g816(.A(G225), .ZN(G308));
endmodule


