//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 0 1 0 0 0 0 0 0 1 0 1 1 0 1 0 1 1 0 1 1 0 1 1 1 0 1 1 0 1 0 1 0 1 1 1 1 0 1 1 0 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 0 1 0 0 0 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:21:32 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n705,
    new_n707, new_n708, new_n710, new_n711, new_n712, new_n713, new_n714,
    new_n715, new_n716, new_n717, new_n718, new_n720, new_n721, new_n722,
    new_n723, new_n724, new_n725, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n756, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n783, new_n784, new_n785, new_n786, new_n787, new_n788, new_n789,
    new_n790, new_n791, new_n792, new_n793, new_n794, new_n795, new_n796,
    new_n797, new_n798, new_n799, new_n800, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n912, new_n913, new_n914, new_n915, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n932, new_n933, new_n934,
    new_n935, new_n936, new_n937, new_n938, new_n939, new_n940, new_n941,
    new_n942, new_n943, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n951, new_n952, new_n953, new_n954, new_n955, new_n956,
    new_n958, new_n959, new_n960, new_n961, new_n962, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n989, new_n990, new_n991, new_n992, new_n993, new_n994,
    new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003;
  INV_X1    g000(.A(KEYINPUT32), .ZN(new_n187));
  OR2_X1    g001(.A1(KEYINPUT72), .A2(G953), .ZN(new_n188));
  NAND2_X1  g002(.A1(KEYINPUT72), .A2(G953), .ZN(new_n189));
  AOI21_X1  g003(.A(G237), .B1(new_n188), .B2(new_n189), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n190), .A2(G210), .ZN(new_n191));
  XOR2_X1   g005(.A(KEYINPUT26), .B(G101), .Z(new_n192));
  XNOR2_X1  g006(.A(new_n191), .B(new_n192), .ZN(new_n193));
  XNOR2_X1  g007(.A(KEYINPUT73), .B(KEYINPUT27), .ZN(new_n194));
  XNOR2_X1  g008(.A(new_n193), .B(new_n194), .ZN(new_n195));
  INV_X1    g009(.A(G128), .ZN(new_n196));
  NOR2_X1   g010(.A1(new_n196), .A2(KEYINPUT1), .ZN(new_n197));
  INV_X1    g011(.A(G146), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n198), .A2(G143), .ZN(new_n199));
  INV_X1    g013(.A(G143), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n200), .A2(G146), .ZN(new_n201));
  NAND3_X1  g015(.A1(new_n197), .A2(new_n199), .A3(new_n201), .ZN(new_n202));
  NAND3_X1  g016(.A1(new_n196), .A2(new_n198), .A3(G143), .ZN(new_n203));
  OAI211_X1 g017(.A(new_n200), .B(G146), .C1(new_n196), .C2(KEYINPUT1), .ZN(new_n204));
  NAND3_X1  g018(.A1(new_n202), .A2(new_n203), .A3(new_n204), .ZN(new_n205));
  INV_X1    g019(.A(G134), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n206), .A2(G137), .ZN(new_n207));
  INV_X1    g021(.A(new_n207), .ZN(new_n208));
  NOR2_X1   g022(.A1(new_n206), .A2(G137), .ZN(new_n209));
  OAI21_X1  g023(.A(G131), .B1(new_n208), .B2(new_n209), .ZN(new_n210));
  INV_X1    g024(.A(KEYINPUT11), .ZN(new_n211));
  OAI21_X1  g025(.A(new_n211), .B1(new_n206), .B2(G137), .ZN(new_n212));
  INV_X1    g026(.A(G137), .ZN(new_n213));
  NAND3_X1  g027(.A1(new_n213), .A2(KEYINPUT11), .A3(G134), .ZN(new_n214));
  INV_X1    g028(.A(G131), .ZN(new_n215));
  NAND4_X1  g029(.A1(new_n212), .A2(new_n214), .A3(new_n215), .A4(new_n207), .ZN(new_n216));
  NAND3_X1  g030(.A1(new_n205), .A2(new_n210), .A3(new_n216), .ZN(new_n217));
  INV_X1    g031(.A(KEYINPUT71), .ZN(new_n218));
  XNOR2_X1  g032(.A(new_n217), .B(new_n218), .ZN(new_n219));
  NAND2_X1  g033(.A1(KEYINPUT2), .A2(G113), .ZN(new_n220));
  INV_X1    g034(.A(KEYINPUT66), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  NAND3_X1  g036(.A1(KEYINPUT66), .A2(KEYINPUT2), .A3(G113), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  OR2_X1    g038(.A1(KEYINPUT2), .A2(G113), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  INV_X1    g040(.A(new_n226), .ZN(new_n227));
  INV_X1    g041(.A(KEYINPUT69), .ZN(new_n228));
  INV_X1    g042(.A(G119), .ZN(new_n229));
  OR2_X1    g043(.A1(KEYINPUT68), .A2(G116), .ZN(new_n230));
  NAND2_X1  g044(.A1(KEYINPUT68), .A2(G116), .ZN(new_n231));
  AOI21_X1  g045(.A(new_n229), .B1(new_n230), .B2(new_n231), .ZN(new_n232));
  INV_X1    g046(.A(G116), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n229), .A2(KEYINPUT67), .ZN(new_n234));
  INV_X1    g048(.A(KEYINPUT67), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n235), .A2(G119), .ZN(new_n236));
  AOI21_X1  g050(.A(new_n233), .B1(new_n234), .B2(new_n236), .ZN(new_n237));
  OAI21_X1  g051(.A(new_n228), .B1(new_n232), .B2(new_n237), .ZN(new_n238));
  AND2_X1   g052(.A1(KEYINPUT68), .A2(G116), .ZN(new_n239));
  NOR2_X1   g053(.A1(KEYINPUT68), .A2(G116), .ZN(new_n240));
  OAI21_X1  g054(.A(G119), .B1(new_n239), .B2(new_n240), .ZN(new_n241));
  XNOR2_X1  g055(.A(KEYINPUT67), .B(G119), .ZN(new_n242));
  OAI211_X1 g056(.A(new_n241), .B(KEYINPUT69), .C1(new_n233), .C2(new_n242), .ZN(new_n243));
  AOI21_X1  g057(.A(new_n227), .B1(new_n238), .B2(new_n243), .ZN(new_n244));
  NOR3_X1   g058(.A1(new_n226), .A2(new_n237), .A3(new_n232), .ZN(new_n245));
  NOR2_X1   g059(.A1(new_n244), .A2(new_n245), .ZN(new_n246));
  NAND3_X1  g060(.A1(new_n212), .A2(new_n207), .A3(new_n214), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n247), .A2(G131), .ZN(new_n248));
  NAND3_X1  g062(.A1(new_n248), .A2(KEYINPUT64), .A3(new_n216), .ZN(new_n249));
  INV_X1    g063(.A(KEYINPUT64), .ZN(new_n250));
  NAND3_X1  g064(.A1(new_n247), .A2(new_n250), .A3(G131), .ZN(new_n251));
  XNOR2_X1  g065(.A(G143), .B(G146), .ZN(new_n252));
  INV_X1    g066(.A(KEYINPUT0), .ZN(new_n253));
  OAI21_X1  g067(.A(new_n252), .B1(new_n253), .B2(new_n196), .ZN(new_n254));
  XOR2_X1   g068(.A(KEYINPUT0), .B(G128), .Z(new_n255));
  OAI21_X1  g069(.A(new_n254), .B1(new_n252), .B2(new_n255), .ZN(new_n256));
  NAND3_X1  g070(.A1(new_n249), .A2(new_n251), .A3(new_n256), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n257), .A2(KEYINPUT70), .ZN(new_n258));
  INV_X1    g072(.A(KEYINPUT70), .ZN(new_n259));
  NAND4_X1  g073(.A1(new_n249), .A2(new_n256), .A3(new_n259), .A4(new_n251), .ZN(new_n260));
  NAND4_X1  g074(.A1(new_n219), .A2(new_n246), .A3(new_n258), .A4(new_n260), .ZN(new_n261));
  INV_X1    g075(.A(new_n217), .ZN(new_n262));
  INV_X1    g076(.A(KEYINPUT65), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n257), .A2(new_n263), .ZN(new_n264));
  NAND4_X1  g078(.A1(new_n249), .A2(new_n256), .A3(KEYINPUT65), .A4(new_n251), .ZN(new_n265));
  AOI21_X1  g079(.A(new_n262), .B1(new_n264), .B2(new_n265), .ZN(new_n266));
  OAI21_X1  g080(.A(new_n261), .B1(new_n266), .B2(new_n246), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n267), .A2(KEYINPUT28), .ZN(new_n268));
  AND3_X1   g082(.A1(new_n246), .A2(new_n217), .A3(new_n257), .ZN(new_n269));
  NOR2_X1   g083(.A1(new_n269), .A2(KEYINPUT28), .ZN(new_n270));
  INV_X1    g084(.A(new_n270), .ZN(new_n271));
  AOI21_X1  g085(.A(new_n195), .B1(new_n268), .B2(new_n271), .ZN(new_n272));
  INV_X1    g086(.A(KEYINPUT31), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n261), .A2(new_n195), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n274), .A2(KEYINPUT74), .ZN(new_n275));
  INV_X1    g089(.A(KEYINPUT74), .ZN(new_n276));
  NAND3_X1  g090(.A1(new_n261), .A2(new_n276), .A3(new_n195), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n275), .A2(new_n277), .ZN(new_n278));
  NAND3_X1  g092(.A1(new_n219), .A2(new_n258), .A3(new_n260), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n279), .A2(KEYINPUT30), .ZN(new_n280));
  INV_X1    g094(.A(KEYINPUT30), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n266), .A2(new_n281), .ZN(new_n282));
  AOI21_X1  g096(.A(new_n246), .B1(new_n280), .B2(new_n282), .ZN(new_n283));
  OAI21_X1  g097(.A(new_n273), .B1(new_n278), .B2(new_n283), .ZN(new_n284));
  AND3_X1   g098(.A1(new_n261), .A2(new_n276), .A3(new_n195), .ZN(new_n285));
  AOI21_X1  g099(.A(new_n276), .B1(new_n261), .B2(new_n195), .ZN(new_n286));
  NOR2_X1   g100(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n280), .A2(new_n282), .ZN(new_n288));
  INV_X1    g102(.A(new_n246), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  NAND3_X1  g104(.A1(new_n287), .A2(KEYINPUT31), .A3(new_n290), .ZN(new_n291));
  AOI21_X1  g105(.A(new_n272), .B1(new_n284), .B2(new_n291), .ZN(new_n292));
  NOR2_X1   g106(.A1(G472), .A2(G902), .ZN(new_n293));
  INV_X1    g107(.A(new_n293), .ZN(new_n294));
  OAI21_X1  g108(.A(new_n187), .B1(new_n292), .B2(new_n294), .ZN(new_n295));
  INV_X1    g109(.A(new_n272), .ZN(new_n296));
  AOI21_X1  g110(.A(KEYINPUT31), .B1(new_n287), .B2(new_n290), .ZN(new_n297));
  NOR4_X1   g111(.A1(new_n283), .A2(new_n285), .A3(new_n286), .A4(new_n273), .ZN(new_n298));
  OAI21_X1  g112(.A(new_n296), .B1(new_n297), .B2(new_n298), .ZN(new_n299));
  NAND3_X1  g113(.A1(new_n299), .A2(KEYINPUT32), .A3(new_n293), .ZN(new_n300));
  INV_X1    g114(.A(KEYINPUT75), .ZN(new_n301));
  NAND3_X1  g115(.A1(new_n295), .A2(new_n300), .A3(new_n301), .ZN(new_n302));
  NOR2_X1   g116(.A1(new_n292), .A2(new_n294), .ZN(new_n303));
  NAND3_X1  g117(.A1(new_n303), .A2(KEYINPUT75), .A3(KEYINPUT32), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n302), .A2(new_n304), .ZN(new_n305));
  INV_X1    g119(.A(G472), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n290), .A2(new_n261), .ZN(new_n307));
  INV_X1    g121(.A(new_n195), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  INV_X1    g123(.A(KEYINPUT29), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n268), .A2(new_n271), .ZN(new_n311));
  OAI211_X1 g125(.A(new_n309), .B(new_n310), .C1(new_n308), .C2(new_n311), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n279), .A2(new_n289), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n313), .A2(new_n261), .ZN(new_n314));
  AOI21_X1  g128(.A(new_n270), .B1(new_n314), .B2(KEYINPUT28), .ZN(new_n315));
  NOR2_X1   g129(.A1(new_n308), .A2(new_n310), .ZN(new_n316));
  AOI21_X1  g130(.A(G902), .B1(new_n315), .B2(new_n316), .ZN(new_n317));
  AOI21_X1  g131(.A(new_n306), .B1(new_n312), .B2(new_n317), .ZN(new_n318));
  INV_X1    g132(.A(new_n318), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n305), .A2(new_n319), .ZN(new_n320));
  INV_X1    g134(.A(G125), .ZN(new_n321));
  NOR3_X1   g135(.A1(new_n321), .A2(KEYINPUT16), .A3(G140), .ZN(new_n322));
  NAND2_X1  g136(.A1(KEYINPUT76), .A2(G125), .ZN(new_n323));
  INV_X1    g137(.A(G140), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n323), .A2(new_n324), .ZN(new_n325));
  NAND3_X1  g139(.A1(KEYINPUT76), .A2(G125), .A3(G140), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  AOI211_X1 g141(.A(new_n198), .B(new_n322), .C1(new_n327), .C2(KEYINPUT16), .ZN(new_n328));
  INV_X1    g142(.A(G110), .ZN(new_n329));
  INV_X1    g143(.A(KEYINPUT23), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n234), .A2(new_n236), .ZN(new_n331));
  OAI21_X1  g145(.A(new_n330), .B1(new_n331), .B2(G128), .ZN(new_n332));
  NOR2_X1   g146(.A1(new_n229), .A2(G128), .ZN(new_n333));
  AOI21_X1  g147(.A(new_n333), .B1(new_n331), .B2(G128), .ZN(new_n334));
  OAI211_X1 g148(.A(new_n329), .B(new_n332), .C1(new_n334), .C2(new_n330), .ZN(new_n335));
  INV_X1    g149(.A(new_n333), .ZN(new_n336));
  OAI21_X1  g150(.A(new_n336), .B1(new_n242), .B2(new_n196), .ZN(new_n337));
  XNOR2_X1  g151(.A(KEYINPUT24), .B(G110), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n337), .A2(new_n338), .ZN(new_n339));
  AOI21_X1  g153(.A(new_n328), .B1(new_n335), .B2(new_n339), .ZN(new_n340));
  XNOR2_X1  g154(.A(G125), .B(G140), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n341), .A2(new_n198), .ZN(new_n342));
  NAND3_X1  g156(.A1(new_n340), .A2(KEYINPUT77), .A3(new_n342), .ZN(new_n343));
  INV_X1    g157(.A(new_n343), .ZN(new_n344));
  AOI21_X1  g158(.A(KEYINPUT77), .B1(new_n340), .B2(new_n342), .ZN(new_n345));
  NOR2_X1   g159(.A1(new_n344), .A2(new_n345), .ZN(new_n346));
  INV_X1    g160(.A(KEYINPUT79), .ZN(new_n347));
  OR2_X1    g161(.A1(new_n337), .A2(new_n338), .ZN(new_n348));
  AOI21_X1  g162(.A(new_n322), .B1(new_n327), .B2(KEYINPUT16), .ZN(new_n349));
  NOR2_X1   g163(.A1(new_n349), .A2(G146), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n337), .A2(KEYINPUT23), .ZN(new_n351));
  AND2_X1   g165(.A1(new_n351), .A2(new_n332), .ZN(new_n352));
  OAI221_X1 g166(.A(new_n348), .B1(new_n328), .B2(new_n350), .C1(new_n352), .C2(new_n329), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n188), .A2(new_n189), .ZN(new_n354));
  NAND3_X1  g168(.A1(new_n354), .A2(G221), .A3(G234), .ZN(new_n355));
  OR2_X1    g169(.A1(new_n355), .A2(KEYINPUT22), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n355), .A2(KEYINPUT22), .ZN(new_n357));
  AND3_X1   g171(.A1(new_n356), .A2(G137), .A3(new_n357), .ZN(new_n358));
  AOI21_X1  g172(.A(G137), .B1(new_n356), .B2(new_n357), .ZN(new_n359));
  NOR2_X1   g173(.A1(new_n358), .A2(new_n359), .ZN(new_n360));
  NAND4_X1  g174(.A1(new_n346), .A2(new_n347), .A3(new_n353), .A4(new_n360), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n335), .A2(new_n339), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n349), .A2(G146), .ZN(new_n363));
  NAND3_X1  g177(.A1(new_n362), .A2(new_n363), .A3(new_n342), .ZN(new_n364));
  INV_X1    g178(.A(KEYINPUT77), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  NAND3_X1  g180(.A1(new_n366), .A2(new_n353), .A3(new_n343), .ZN(new_n367));
  INV_X1    g181(.A(new_n360), .ZN(new_n368));
  OAI21_X1  g182(.A(KEYINPUT79), .B1(new_n367), .B2(new_n368), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n361), .A2(new_n369), .ZN(new_n370));
  INV_X1    g184(.A(G902), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n367), .A2(new_n368), .ZN(new_n372));
  INV_X1    g186(.A(KEYINPUT78), .ZN(new_n373));
  NOR2_X1   g187(.A1(new_n372), .A2(new_n373), .ZN(new_n374));
  AOI21_X1  g188(.A(KEYINPUT78), .B1(new_n367), .B2(new_n368), .ZN(new_n375));
  OAI211_X1 g189(.A(new_n370), .B(new_n371), .C1(new_n374), .C2(new_n375), .ZN(new_n376));
  NOR2_X1   g190(.A1(KEYINPUT80), .A2(KEYINPUT25), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n376), .A2(new_n377), .ZN(new_n378));
  XNOR2_X1  g192(.A(new_n372), .B(new_n373), .ZN(new_n379));
  INV_X1    g193(.A(new_n377), .ZN(new_n380));
  NAND4_X1  g194(.A1(new_n379), .A2(new_n371), .A3(new_n370), .A4(new_n380), .ZN(new_n381));
  NAND2_X1  g195(.A1(KEYINPUT80), .A2(KEYINPUT25), .ZN(new_n382));
  NAND3_X1  g196(.A1(new_n378), .A2(new_n381), .A3(new_n382), .ZN(new_n383));
  INV_X1    g197(.A(G217), .ZN(new_n384));
  AOI21_X1  g198(.A(new_n384), .B1(G234), .B2(new_n371), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n383), .A2(new_n385), .ZN(new_n386));
  AND2_X1   g200(.A1(new_n379), .A2(new_n370), .ZN(new_n387));
  NOR2_X1   g201(.A1(new_n385), .A2(G902), .ZN(new_n388));
  XNOR2_X1  g202(.A(new_n388), .B(KEYINPUT81), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n387), .A2(new_n389), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n386), .A2(new_n390), .ZN(new_n391));
  INV_X1    g205(.A(new_n391), .ZN(new_n392));
  NAND2_X1  g206(.A1(G469), .A2(G902), .ZN(new_n393));
  INV_X1    g207(.A(KEYINPUT84), .ZN(new_n394));
  XNOR2_X1  g208(.A(G104), .B(G107), .ZN(new_n395));
  INV_X1    g209(.A(G101), .ZN(new_n396));
  OAI21_X1  g210(.A(new_n394), .B1(new_n395), .B2(new_n396), .ZN(new_n397));
  XNOR2_X1  g211(.A(KEYINPUT83), .B(G101), .ZN(new_n398));
  INV_X1    g212(.A(G104), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n399), .A2(G107), .ZN(new_n400));
  INV_X1    g214(.A(KEYINPUT3), .ZN(new_n401));
  INV_X1    g215(.A(G107), .ZN(new_n402));
  NAND3_X1  g216(.A1(new_n401), .A2(new_n402), .A3(G104), .ZN(new_n403));
  OAI21_X1  g217(.A(KEYINPUT3), .B1(new_n399), .B2(G107), .ZN(new_n404));
  NAND4_X1  g218(.A1(new_n398), .A2(new_n400), .A3(new_n403), .A4(new_n404), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n402), .A2(G104), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n400), .A2(new_n406), .ZN(new_n407));
  NAND3_X1  g221(.A1(new_n407), .A2(KEYINPUT84), .A3(G101), .ZN(new_n408));
  NAND3_X1  g222(.A1(new_n397), .A2(new_n405), .A3(new_n408), .ZN(new_n409));
  INV_X1    g223(.A(new_n205), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n409), .A2(new_n410), .ZN(new_n411));
  NAND4_X1  g225(.A1(new_n205), .A2(new_n397), .A3(new_n405), .A4(new_n408), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n411), .A2(new_n412), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n249), .A2(new_n251), .ZN(new_n414));
  INV_X1    g228(.A(new_n414), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n413), .A2(new_n415), .ZN(new_n416));
  INV_X1    g230(.A(KEYINPUT12), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  NAND3_X1  g232(.A1(new_n413), .A2(new_n415), .A3(KEYINPUT12), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n418), .A2(new_n419), .ZN(new_n420));
  AND2_X1   g234(.A1(new_n397), .A2(new_n408), .ZN(new_n421));
  NAND4_X1  g235(.A1(new_n421), .A2(KEYINPUT10), .A3(new_n205), .A4(new_n405), .ZN(new_n422));
  NAND3_X1  g236(.A1(new_n404), .A2(new_n403), .A3(new_n400), .ZN(new_n423));
  INV_X1    g237(.A(KEYINPUT4), .ZN(new_n424));
  NAND3_X1  g238(.A1(new_n423), .A2(new_n424), .A3(G101), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n405), .A2(KEYINPUT4), .ZN(new_n426));
  AND2_X1   g240(.A1(new_n423), .A2(G101), .ZN(new_n427));
  OAI211_X1 g241(.A(new_n256), .B(new_n425), .C1(new_n426), .C2(new_n427), .ZN(new_n428));
  INV_X1    g242(.A(KEYINPUT10), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n412), .A2(new_n429), .ZN(new_n430));
  NAND4_X1  g244(.A1(new_n422), .A2(new_n428), .A3(new_n430), .A4(new_n414), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n354), .A2(G227), .ZN(new_n432));
  XNOR2_X1  g246(.A(G110), .B(G140), .ZN(new_n433));
  XNOR2_X1  g247(.A(new_n432), .B(new_n433), .ZN(new_n434));
  AND2_X1   g248(.A1(new_n431), .A2(new_n434), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n420), .A2(new_n435), .ZN(new_n436));
  NAND3_X1  g250(.A1(new_n422), .A2(new_n428), .A3(new_n430), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n437), .A2(new_n415), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n438), .A2(new_n431), .ZN(new_n439));
  INV_X1    g253(.A(new_n434), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n439), .A2(new_n440), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n436), .A2(new_n441), .ZN(new_n442));
  INV_X1    g256(.A(G469), .ZN(new_n443));
  NAND3_X1  g257(.A1(new_n442), .A2(new_n443), .A3(new_n371), .ZN(new_n444));
  INV_X1    g258(.A(KEYINPUT85), .ZN(new_n445));
  AOI21_X1  g259(.A(new_n434), .B1(new_n420), .B2(new_n431), .ZN(new_n446));
  AND3_X1   g260(.A1(new_n438), .A2(new_n431), .A3(new_n434), .ZN(new_n447));
  OAI21_X1  g261(.A(new_n445), .B1(new_n446), .B2(new_n447), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n435), .A2(new_n438), .ZN(new_n449));
  INV_X1    g263(.A(new_n437), .ZN(new_n450));
  AOI22_X1  g264(.A1(new_n418), .A2(new_n419), .B1(new_n450), .B2(new_n414), .ZN(new_n451));
  OAI211_X1 g265(.A(new_n449), .B(KEYINPUT85), .C1(new_n451), .C2(new_n434), .ZN(new_n452));
  AND2_X1   g266(.A1(new_n448), .A2(new_n452), .ZN(new_n453));
  OAI211_X1 g267(.A(new_n393), .B(new_n444), .C1(new_n453), .C2(new_n443), .ZN(new_n454));
  XNOR2_X1  g268(.A(KEYINPUT9), .B(G234), .ZN(new_n455));
  OAI21_X1  g269(.A(G221), .B1(new_n455), .B2(G902), .ZN(new_n456));
  XNOR2_X1  g270(.A(new_n456), .B(KEYINPUT82), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n454), .A2(new_n457), .ZN(new_n458));
  INV_X1    g272(.A(new_n458), .ZN(new_n459));
  XOR2_X1   g273(.A(G110), .B(G122), .Z(new_n460));
  OAI21_X1  g274(.A(new_n425), .B1(new_n426), .B2(new_n427), .ZN(new_n461));
  NOR2_X1   g275(.A1(new_n246), .A2(new_n461), .ZN(new_n462));
  NAND3_X1  g276(.A1(new_n238), .A2(KEYINPUT5), .A3(new_n243), .ZN(new_n463));
  INV_X1    g277(.A(G113), .ZN(new_n464));
  INV_X1    g278(.A(KEYINPUT5), .ZN(new_n465));
  AOI21_X1  g279(.A(new_n464), .B1(new_n237), .B2(new_n465), .ZN(new_n466));
  AOI211_X1 g280(.A(new_n409), .B(new_n245), .C1(new_n463), .C2(new_n466), .ZN(new_n467));
  OAI21_X1  g281(.A(new_n460), .B1(new_n462), .B2(new_n467), .ZN(new_n468));
  OAI221_X1 g282(.A(new_n425), .B1(new_n427), .B2(new_n426), .C1(new_n244), .C2(new_n245), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n463), .A2(new_n466), .ZN(new_n470));
  INV_X1    g284(.A(new_n245), .ZN(new_n471));
  NAND4_X1  g285(.A1(new_n470), .A2(new_n471), .A3(new_n405), .A4(new_n421), .ZN(new_n472));
  INV_X1    g286(.A(new_n460), .ZN(new_n473));
  NAND3_X1  g287(.A1(new_n469), .A2(new_n472), .A3(new_n473), .ZN(new_n474));
  NAND3_X1  g288(.A1(new_n468), .A2(new_n474), .A3(KEYINPUT6), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n256), .A2(G125), .ZN(new_n476));
  OAI21_X1  g290(.A(new_n476), .B1(G125), .B2(new_n410), .ZN(new_n477));
  XNOR2_X1  g291(.A(KEYINPUT87), .B(G224), .ZN(new_n478));
  INV_X1    g292(.A(G953), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  XNOR2_X1  g294(.A(new_n477), .B(new_n480), .ZN(new_n481));
  INV_X1    g295(.A(KEYINPUT6), .ZN(new_n482));
  OAI211_X1 g296(.A(new_n482), .B(new_n460), .C1(new_n462), .C2(new_n467), .ZN(new_n483));
  NAND3_X1  g297(.A1(new_n475), .A2(new_n481), .A3(new_n483), .ZN(new_n484));
  NAND3_X1  g298(.A1(new_n470), .A2(new_n471), .A3(new_n409), .ZN(new_n485));
  XOR2_X1   g299(.A(new_n460), .B(KEYINPUT8), .Z(new_n486));
  XNOR2_X1  g300(.A(new_n466), .B(KEYINPUT88), .ZN(new_n487));
  OAI211_X1 g301(.A(new_n241), .B(KEYINPUT5), .C1(new_n233), .C2(new_n242), .ZN(new_n488));
  AOI21_X1  g302(.A(new_n245), .B1(new_n487), .B2(new_n488), .ZN(new_n489));
  OAI211_X1 g303(.A(new_n485), .B(new_n486), .C1(new_n489), .C2(new_n409), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n480), .A2(KEYINPUT7), .ZN(new_n491));
  XNOR2_X1  g305(.A(new_n477), .B(new_n491), .ZN(new_n492));
  NAND3_X1  g306(.A1(new_n490), .A2(new_n474), .A3(new_n492), .ZN(new_n493));
  NAND3_X1  g307(.A1(new_n484), .A2(new_n371), .A3(new_n493), .ZN(new_n494));
  OAI21_X1  g308(.A(G210), .B1(G237), .B2(G902), .ZN(new_n495));
  INV_X1    g309(.A(new_n495), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n494), .A2(new_n496), .ZN(new_n497));
  NAND4_X1  g311(.A1(new_n484), .A2(new_n371), .A3(new_n495), .A4(new_n493), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  OAI21_X1  g313(.A(G214), .B1(G237), .B2(G902), .ZN(new_n500));
  XOR2_X1   g314(.A(new_n500), .B(KEYINPUT86), .Z(new_n501));
  INV_X1    g315(.A(G952), .ZN(new_n502));
  AOI211_X1 g316(.A(G953), .B(new_n502), .C1(G234), .C2(G237), .ZN(new_n503));
  AOI211_X1 g317(.A(new_n371), .B(new_n354), .C1(G234), .C2(G237), .ZN(new_n504));
  XOR2_X1   g318(.A(KEYINPUT21), .B(G898), .Z(new_n505));
  INV_X1    g319(.A(new_n505), .ZN(new_n506));
  AOI21_X1  g320(.A(new_n503), .B1(new_n504), .B2(new_n506), .ZN(new_n507));
  INV_X1    g321(.A(new_n507), .ZN(new_n508));
  NAND3_X1  g322(.A1(new_n499), .A2(new_n501), .A3(new_n508), .ZN(new_n509));
  INV_X1    g323(.A(new_n509), .ZN(new_n510));
  INV_X1    g324(.A(KEYINPUT92), .ZN(new_n511));
  XNOR2_X1  g325(.A(G113), .B(G122), .ZN(new_n512));
  XNOR2_X1  g326(.A(new_n512), .B(new_n399), .ZN(new_n513));
  INV_X1    g327(.A(new_n513), .ZN(new_n514));
  AOI21_X1  g328(.A(G143), .B1(new_n190), .B2(G214), .ZN(new_n515));
  INV_X1    g329(.A(G237), .ZN(new_n516));
  AND2_X1   g330(.A1(KEYINPUT72), .A2(G953), .ZN(new_n517));
  NOR2_X1   g331(.A1(KEYINPUT72), .A2(G953), .ZN(new_n518));
  OAI211_X1 g332(.A(G214), .B(new_n516), .C1(new_n517), .C2(new_n518), .ZN(new_n519));
  NOR2_X1   g333(.A1(new_n519), .A2(new_n200), .ZN(new_n520));
  OAI21_X1  g334(.A(G131), .B1(new_n515), .B2(new_n520), .ZN(new_n521));
  INV_X1    g335(.A(KEYINPUT18), .ZN(new_n522));
  NOR2_X1   g336(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  OAI21_X1  g337(.A(new_n342), .B1(new_n327), .B2(new_n198), .ZN(new_n524));
  NAND3_X1  g338(.A1(new_n190), .A2(G143), .A3(G214), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n519), .A2(new_n200), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  NOR2_X1   g341(.A1(new_n522), .A2(new_n215), .ZN(new_n528));
  OAI21_X1  g342(.A(new_n524), .B1(new_n527), .B2(new_n528), .ZN(new_n529));
  NOR2_X1   g343(.A1(new_n523), .A2(new_n529), .ZN(new_n530));
  NOR2_X1   g344(.A1(new_n341), .A2(KEYINPUT19), .ZN(new_n531));
  INV_X1    g345(.A(KEYINPUT19), .ZN(new_n532));
  AOI21_X1  g346(.A(new_n532), .B1(new_n325), .B2(new_n326), .ZN(new_n533));
  NOR2_X1   g347(.A1(new_n531), .A2(new_n533), .ZN(new_n534));
  OAI21_X1  g348(.A(new_n363), .B1(new_n534), .B2(G146), .ZN(new_n535));
  NAND3_X1  g349(.A1(new_n525), .A2(new_n215), .A3(new_n526), .ZN(new_n536));
  AOI21_X1  g350(.A(new_n535), .B1(new_n521), .B2(new_n536), .ZN(new_n537));
  OAI21_X1  g351(.A(new_n514), .B1(new_n530), .B2(new_n537), .ZN(new_n538));
  NOR2_X1   g352(.A1(new_n350), .A2(new_n328), .ZN(new_n539));
  NAND3_X1  g353(.A1(new_n527), .A2(KEYINPUT17), .A3(G131), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n521), .A2(new_n536), .ZN(new_n541));
  OAI211_X1 g355(.A(new_n539), .B(new_n540), .C1(new_n541), .C2(KEYINPUT17), .ZN(new_n542));
  OAI221_X1 g356(.A(new_n524), .B1(new_n527), .B2(new_n528), .C1(new_n521), .C2(new_n522), .ZN(new_n543));
  NAND3_X1  g357(.A1(new_n542), .A2(new_n543), .A3(new_n513), .ZN(new_n544));
  AOI21_X1  g358(.A(G475), .B1(new_n538), .B2(new_n544), .ZN(new_n545));
  NAND3_X1  g359(.A1(new_n545), .A2(KEYINPUT20), .A3(new_n371), .ZN(new_n546));
  INV_X1    g360(.A(new_n546), .ZN(new_n547));
  AOI21_X1  g361(.A(KEYINPUT20), .B1(new_n545), .B2(new_n371), .ZN(new_n548));
  NOR2_X1   g362(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  INV_X1    g363(.A(new_n544), .ZN(new_n550));
  AOI21_X1  g364(.A(new_n513), .B1(new_n542), .B2(new_n543), .ZN(new_n551));
  OAI21_X1  g365(.A(new_n371), .B1(new_n550), .B2(new_n551), .ZN(new_n552));
  INV_X1    g366(.A(KEYINPUT89), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  OAI211_X1 g368(.A(KEYINPUT89), .B(new_n371), .C1(new_n550), .C2(new_n551), .ZN(new_n555));
  NAND3_X1  g369(.A1(new_n554), .A2(G475), .A3(new_n555), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n549), .A2(new_n556), .ZN(new_n557));
  INV_X1    g371(.A(G122), .ZN(new_n558));
  AOI21_X1  g372(.A(new_n558), .B1(new_n230), .B2(new_n231), .ZN(new_n559));
  NOR2_X1   g373(.A1(new_n233), .A2(G122), .ZN(new_n560));
  OAI21_X1  g374(.A(G107), .B1(new_n559), .B2(new_n560), .ZN(new_n561));
  OAI21_X1  g375(.A(G122), .B1(new_n239), .B2(new_n240), .ZN(new_n562));
  INV_X1    g376(.A(new_n560), .ZN(new_n563));
  NAND3_X1  g377(.A1(new_n562), .A2(new_n402), .A3(new_n563), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n561), .A2(new_n564), .ZN(new_n565));
  XNOR2_X1  g379(.A(G128), .B(G143), .ZN(new_n566));
  AOI21_X1  g380(.A(new_n206), .B1(new_n566), .B2(KEYINPUT13), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n200), .A2(G128), .ZN(new_n568));
  OAI21_X1  g382(.A(new_n567), .B1(KEYINPUT13), .B2(new_n568), .ZN(new_n569));
  INV_X1    g383(.A(KEYINPUT90), .ZN(new_n570));
  AOI21_X1  g384(.A(new_n570), .B1(new_n566), .B2(new_n206), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n196), .A2(G143), .ZN(new_n572));
  AND4_X1   g386(.A1(new_n570), .A2(new_n572), .A3(new_n568), .A4(new_n206), .ZN(new_n573));
  NOR2_X1   g387(.A1(new_n571), .A2(new_n573), .ZN(new_n574));
  NAND3_X1  g388(.A1(new_n565), .A2(new_n569), .A3(new_n574), .ZN(new_n575));
  INV_X1    g389(.A(KEYINPUT14), .ZN(new_n576));
  NAND3_X1  g390(.A1(new_n562), .A2(new_n576), .A3(new_n563), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n559), .A2(KEYINPUT14), .ZN(new_n578));
  NAND3_X1  g392(.A1(new_n577), .A2(new_n578), .A3(G107), .ZN(new_n579));
  XNOR2_X1  g393(.A(new_n566), .B(new_n206), .ZN(new_n580));
  NAND3_X1  g394(.A1(new_n579), .A2(new_n580), .A3(new_n564), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n575), .A2(new_n581), .ZN(new_n582));
  NOR3_X1   g396(.A1(new_n455), .A2(new_n384), .A3(G953), .ZN(new_n583));
  INV_X1    g397(.A(new_n583), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n582), .A2(new_n584), .ZN(new_n585));
  NAND3_X1  g399(.A1(new_n575), .A2(new_n581), .A3(new_n583), .ZN(new_n586));
  NAND3_X1  g400(.A1(new_n585), .A2(KEYINPUT91), .A3(new_n586), .ZN(new_n587));
  INV_X1    g401(.A(KEYINPUT91), .ZN(new_n588));
  NAND3_X1  g402(.A1(new_n582), .A2(new_n588), .A3(new_n584), .ZN(new_n589));
  NAND3_X1  g403(.A1(new_n587), .A2(new_n371), .A3(new_n589), .ZN(new_n590));
  INV_X1    g404(.A(G478), .ZN(new_n591));
  NOR2_X1   g405(.A1(new_n591), .A2(KEYINPUT15), .ZN(new_n592));
  XOR2_X1   g406(.A(new_n590), .B(new_n592), .Z(new_n593));
  INV_X1    g407(.A(new_n593), .ZN(new_n594));
  NOR2_X1   g408(.A1(new_n557), .A2(new_n594), .ZN(new_n595));
  NAND4_X1  g409(.A1(new_n459), .A2(new_n510), .A3(new_n511), .A4(new_n595), .ZN(new_n596));
  NAND3_X1  g410(.A1(new_n595), .A2(new_n457), .A3(new_n454), .ZN(new_n597));
  OAI21_X1  g411(.A(KEYINPUT92), .B1(new_n597), .B2(new_n509), .ZN(new_n598));
  NAND4_X1  g412(.A1(new_n320), .A2(new_n392), .A3(new_n596), .A4(new_n598), .ZN(new_n599));
  XOR2_X1   g413(.A(new_n599), .B(new_n398), .Z(G3));
  NAND2_X1  g414(.A1(new_n299), .A2(new_n371), .ZN(new_n601));
  AOI21_X1  g415(.A(new_n303), .B1(G472), .B2(new_n601), .ZN(new_n602));
  AND4_X1   g416(.A1(new_n390), .A2(new_n602), .A3(new_n459), .A4(new_n386), .ZN(new_n603));
  XOR2_X1   g417(.A(new_n603), .B(KEYINPUT93), .Z(new_n604));
  INV_X1    g418(.A(KEYINPUT33), .ZN(new_n605));
  NAND3_X1  g419(.A1(new_n587), .A2(new_n605), .A3(new_n589), .ZN(new_n606));
  INV_X1    g420(.A(KEYINPUT95), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  AND2_X1   g422(.A1(new_n585), .A2(new_n586), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n609), .A2(KEYINPUT33), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n608), .A2(new_n610), .ZN(new_n611));
  NAND3_X1  g425(.A1(new_n609), .A2(new_n607), .A3(KEYINPUT33), .ZN(new_n612));
  NAND4_X1  g426(.A1(new_n611), .A2(G478), .A3(new_n371), .A4(new_n612), .ZN(new_n613));
  INV_X1    g427(.A(KEYINPUT96), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  INV_X1    g429(.A(new_n612), .ZN(new_n616));
  AOI21_X1  g430(.A(new_n616), .B1(new_n608), .B2(new_n610), .ZN(new_n617));
  NAND4_X1  g431(.A1(new_n617), .A2(KEYINPUT96), .A3(G478), .A4(new_n371), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n590), .A2(new_n591), .ZN(new_n619));
  NAND3_X1  g433(.A1(new_n615), .A2(new_n618), .A3(new_n619), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n620), .A2(new_n557), .ZN(new_n621));
  INV_X1    g435(.A(new_n500), .ZN(new_n622));
  INV_X1    g436(.A(new_n498), .ZN(new_n623));
  INV_X1    g437(.A(KEYINPUT94), .ZN(new_n624));
  AOI21_X1  g438(.A(new_n622), .B1(new_n623), .B2(new_n624), .ZN(new_n625));
  NAND3_X1  g439(.A1(new_n497), .A2(KEYINPUT94), .A3(new_n498), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  NOR3_X1   g441(.A1(new_n621), .A2(new_n507), .A3(new_n627), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n604), .A2(new_n628), .ZN(new_n629));
  XOR2_X1   g443(.A(KEYINPUT34), .B(G104), .Z(new_n630));
  XNOR2_X1  g444(.A(new_n629), .B(new_n630), .ZN(G6));
  AND2_X1   g445(.A1(new_n625), .A2(new_n626), .ZN(new_n632));
  INV_X1    g446(.A(KEYINPUT97), .ZN(new_n633));
  AND3_X1   g447(.A1(new_n554), .A2(G475), .A3(new_n555), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n545), .A2(new_n371), .ZN(new_n635));
  INV_X1    g449(.A(KEYINPUT20), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n637), .A2(new_n546), .ZN(new_n638));
  NOR3_X1   g452(.A1(new_n634), .A2(new_n638), .A3(new_n593), .ZN(new_n639));
  NAND4_X1  g453(.A1(new_n632), .A2(new_n633), .A3(new_n508), .A4(new_n639), .ZN(new_n640));
  NAND4_X1  g454(.A1(new_n639), .A2(new_n625), .A3(new_n508), .A4(new_n626), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n641), .A2(KEYINPUT97), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n640), .A2(new_n642), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n604), .A2(new_n643), .ZN(new_n644));
  XOR2_X1   g458(.A(KEYINPUT35), .B(G107), .Z(new_n645));
  XNOR2_X1  g459(.A(new_n644), .B(new_n645), .ZN(G9));
  NOR2_X1   g460(.A1(new_n368), .A2(KEYINPUT36), .ZN(new_n647));
  XNOR2_X1  g461(.A(new_n647), .B(new_n367), .ZN(new_n648));
  NAND2_X1  g462(.A1(new_n648), .A2(new_n389), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n386), .A2(new_n649), .ZN(new_n650));
  NAND4_X1  g464(.A1(new_n598), .A2(new_n596), .A3(new_n602), .A4(new_n650), .ZN(new_n651));
  XNOR2_X1  g465(.A(new_n651), .B(KEYINPUT98), .ZN(new_n652));
  XOR2_X1   g466(.A(KEYINPUT37), .B(G110), .Z(new_n653));
  XNOR2_X1  g467(.A(new_n652), .B(new_n653), .ZN(G12));
  AOI21_X1  g468(.A(new_n318), .B1(new_n302), .B2(new_n304), .ZN(new_n655));
  NOR2_X1   g469(.A1(new_n655), .A2(new_n458), .ZN(new_n656));
  AOI22_X1  g470(.A1(new_n383), .A2(new_n385), .B1(new_n389), .B2(new_n648), .ZN(new_n657));
  INV_X1    g471(.A(G900), .ZN(new_n658));
  AOI21_X1  g472(.A(new_n503), .B1(new_n504), .B2(new_n658), .ZN(new_n659));
  NOR3_X1   g473(.A1(new_n557), .A2(new_n593), .A3(new_n659), .ZN(new_n660));
  NAND3_X1  g474(.A1(new_n632), .A2(KEYINPUT99), .A3(new_n660), .ZN(new_n661));
  INV_X1    g475(.A(KEYINPUT99), .ZN(new_n662));
  INV_X1    g476(.A(new_n659), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n639), .A2(new_n663), .ZN(new_n664));
  OAI21_X1  g478(.A(new_n662), .B1(new_n664), .B2(new_n627), .ZN(new_n665));
  AOI21_X1  g479(.A(new_n657), .B1(new_n661), .B2(new_n665), .ZN(new_n666));
  NAND2_X1  g480(.A1(new_n656), .A2(new_n666), .ZN(new_n667));
  XNOR2_X1  g481(.A(new_n667), .B(G128), .ZN(G30));
  NAND2_X1  g482(.A1(new_n557), .A2(new_n594), .ZN(new_n669));
  XNOR2_X1  g483(.A(new_n659), .B(KEYINPUT39), .ZN(new_n670));
  NOR2_X1   g484(.A1(new_n458), .A2(new_n670), .ZN(new_n671));
  OR2_X1    g485(.A1(new_n671), .A2(KEYINPUT40), .ZN(new_n672));
  NAND2_X1  g486(.A1(new_n671), .A2(KEYINPUT40), .ZN(new_n673));
  AOI21_X1  g487(.A(new_n669), .B1(new_n672), .B2(new_n673), .ZN(new_n674));
  NAND2_X1  g488(.A1(new_n314), .A2(new_n308), .ZN(new_n675));
  OAI21_X1  g489(.A(new_n675), .B1(new_n278), .B2(new_n283), .ZN(new_n676));
  AOI21_X1  g490(.A(new_n306), .B1(new_n676), .B2(new_n371), .ZN(new_n677));
  AOI21_X1  g491(.A(new_n677), .B1(new_n302), .B2(new_n304), .ZN(new_n678));
  AND3_X1   g492(.A1(new_n497), .A2(KEYINPUT38), .A3(new_n498), .ZN(new_n679));
  AOI21_X1  g493(.A(KEYINPUT38), .B1(new_n497), .B2(new_n498), .ZN(new_n680));
  OR2_X1    g494(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  NOR3_X1   g495(.A1(new_n678), .A2(new_n650), .A3(new_n681), .ZN(new_n682));
  NAND3_X1  g496(.A1(new_n674), .A2(new_n682), .A3(new_n500), .ZN(new_n683));
  XNOR2_X1  g497(.A(new_n683), .B(KEYINPUT100), .ZN(new_n684));
  XNOR2_X1  g498(.A(new_n684), .B(G143), .ZN(G45));
  NAND3_X1  g499(.A1(new_n620), .A2(new_n557), .A3(new_n663), .ZN(new_n686));
  NAND2_X1  g500(.A1(new_n686), .A2(KEYINPUT101), .ZN(new_n687));
  INV_X1    g501(.A(KEYINPUT101), .ZN(new_n688));
  NAND4_X1  g502(.A1(new_n620), .A2(new_n688), .A3(new_n557), .A4(new_n663), .ZN(new_n689));
  AND2_X1   g503(.A1(new_n687), .A2(new_n689), .ZN(new_n690));
  NOR2_X1   g504(.A1(new_n657), .A2(new_n627), .ZN(new_n691));
  NAND4_X1  g505(.A1(new_n690), .A2(new_n320), .A3(new_n459), .A4(new_n691), .ZN(new_n692));
  XNOR2_X1  g506(.A(new_n692), .B(G146), .ZN(G48));
  INV_X1    g507(.A(new_n456), .ZN(new_n694));
  AOI22_X1  g508(.A1(new_n420), .A2(new_n435), .B1(new_n439), .B2(new_n440), .ZN(new_n695));
  OAI21_X1  g509(.A(G469), .B1(new_n695), .B2(G902), .ZN(new_n696));
  INV_X1    g510(.A(KEYINPUT102), .ZN(new_n697));
  NAND3_X1  g511(.A1(new_n696), .A2(new_n444), .A3(new_n697), .ZN(new_n698));
  OAI211_X1 g512(.A(KEYINPUT102), .B(G469), .C1(new_n695), .C2(G902), .ZN(new_n699));
  AOI21_X1  g513(.A(new_n694), .B1(new_n698), .B2(new_n699), .ZN(new_n700));
  XNOR2_X1  g514(.A(new_n700), .B(KEYINPUT103), .ZN(new_n701));
  NAND4_X1  g515(.A1(new_n320), .A2(new_n392), .A3(new_n628), .A4(new_n701), .ZN(new_n702));
  XNOR2_X1  g516(.A(new_n702), .B(KEYINPUT41), .ZN(new_n703));
  XNOR2_X1  g517(.A(new_n703), .B(G113), .ZN(G15));
  NAND4_X1  g518(.A1(new_n643), .A2(new_n320), .A3(new_n392), .A4(new_n701), .ZN(new_n705));
  XNOR2_X1  g519(.A(new_n705), .B(G116), .ZN(G18));
  AND3_X1   g520(.A1(new_n595), .A2(new_n700), .A3(new_n508), .ZN(new_n707));
  NAND3_X1  g521(.A1(new_n320), .A2(new_n691), .A3(new_n707), .ZN(new_n708));
  XNOR2_X1  g522(.A(new_n708), .B(G119), .ZN(G21));
  OAI21_X1  g523(.A(G472), .B1(new_n292), .B2(G902), .ZN(new_n710));
  INV_X1    g524(.A(KEYINPUT105), .ZN(new_n711));
  NAND2_X1  g525(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  NAND3_X1  g526(.A1(new_n601), .A2(KEYINPUT105), .A3(G472), .ZN(new_n713));
  OAI22_X1  g527(.A1(new_n297), .A2(new_n298), .B1(new_n195), .B2(new_n315), .ZN(new_n714));
  XNOR2_X1  g528(.A(new_n293), .B(KEYINPUT104), .ZN(new_n715));
  AOI22_X1  g529(.A1(new_n712), .A2(new_n713), .B1(new_n714), .B2(new_n715), .ZN(new_n716));
  NOR3_X1   g530(.A1(new_n627), .A2(new_n507), .A3(new_n669), .ZN(new_n717));
  NAND4_X1  g531(.A1(new_n716), .A2(new_n392), .A3(new_n701), .A4(new_n717), .ZN(new_n718));
  XNOR2_X1  g532(.A(new_n718), .B(G122), .ZN(G24));
  NAND2_X1  g533(.A1(new_n712), .A2(new_n713), .ZN(new_n720));
  NAND2_X1  g534(.A1(new_n714), .A2(new_n715), .ZN(new_n721));
  AND3_X1   g535(.A1(new_n720), .A2(new_n650), .A3(new_n721), .ZN(new_n722));
  INV_X1    g536(.A(new_n700), .ZN(new_n723));
  NOR2_X1   g537(.A1(new_n627), .A2(new_n723), .ZN(new_n724));
  NAND3_X1  g538(.A1(new_n690), .A2(new_n722), .A3(new_n724), .ZN(new_n725));
  XNOR2_X1  g539(.A(new_n725), .B(G125), .ZN(G27));
  NAND3_X1  g540(.A1(new_n497), .A2(new_n500), .A3(new_n498), .ZN(new_n727));
  INV_X1    g541(.A(KEYINPUT107), .ZN(new_n728));
  NAND2_X1  g542(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  NAND4_X1  g543(.A1(new_n497), .A2(KEYINPUT107), .A3(new_n500), .A4(new_n498), .ZN(new_n730));
  NAND2_X1  g544(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  NOR3_X1   g545(.A1(new_n655), .A2(new_n391), .A3(new_n731), .ZN(new_n732));
  XNOR2_X1  g546(.A(new_n393), .B(KEYINPUT106), .ZN(new_n733));
  OAI21_X1  g547(.A(new_n449), .B1(new_n451), .B2(new_n434), .ZN(new_n734));
  OAI211_X1 g548(.A(new_n444), .B(new_n733), .C1(new_n443), .C2(new_n734), .ZN(new_n735));
  NAND2_X1  g549(.A1(new_n735), .A2(new_n456), .ZN(new_n736));
  INV_X1    g550(.A(new_n736), .ZN(new_n737));
  NAND3_X1  g551(.A1(new_n732), .A2(new_n690), .A3(new_n737), .ZN(new_n738));
  INV_X1    g552(.A(KEYINPUT42), .ZN(new_n739));
  NAND2_X1  g553(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  INV_X1    g554(.A(KEYINPUT108), .ZN(new_n741));
  INV_X1    g555(.A(KEYINPUT109), .ZN(new_n742));
  AND3_X1   g556(.A1(new_n295), .A2(new_n741), .A3(new_n742), .ZN(new_n743));
  AOI21_X1  g557(.A(new_n742), .B1(new_n295), .B2(new_n741), .ZN(new_n744));
  NOR2_X1   g558(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  INV_X1    g559(.A(new_n300), .ZN(new_n746));
  NAND2_X1  g560(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  OAI21_X1  g561(.A(new_n300), .B1(new_n743), .B2(new_n744), .ZN(new_n748));
  NAND3_X1  g562(.A1(new_n747), .A2(new_n748), .A3(new_n319), .ZN(new_n749));
  NAND2_X1  g563(.A1(new_n687), .A2(new_n689), .ZN(new_n750));
  NOR2_X1   g564(.A1(new_n750), .A2(new_n731), .ZN(new_n751));
  NOR2_X1   g565(.A1(new_n736), .A2(new_n739), .ZN(new_n752));
  NAND4_X1  g566(.A1(new_n749), .A2(new_n392), .A3(new_n751), .A4(new_n752), .ZN(new_n753));
  NAND2_X1  g567(.A1(new_n740), .A2(new_n753), .ZN(new_n754));
  XNOR2_X1  g568(.A(new_n754), .B(G131), .ZN(G33));
  NAND3_X1  g569(.A1(new_n732), .A2(new_n660), .A3(new_n737), .ZN(new_n756));
  XNOR2_X1  g570(.A(new_n756), .B(G134), .ZN(G36));
  INV_X1    g571(.A(KEYINPUT43), .ZN(new_n758));
  OAI21_X1  g572(.A(KEYINPUT111), .B1(new_n634), .B2(new_n638), .ZN(new_n759));
  INV_X1    g573(.A(KEYINPUT111), .ZN(new_n760));
  NAND3_X1  g574(.A1(new_n549), .A2(new_n760), .A3(new_n556), .ZN(new_n761));
  NAND2_X1  g575(.A1(new_n759), .A2(new_n761), .ZN(new_n762));
  AOI21_X1  g576(.A(new_n758), .B1(new_n762), .B2(new_n620), .ZN(new_n763));
  INV_X1    g577(.A(new_n557), .ZN(new_n764));
  AND3_X1   g578(.A1(new_n620), .A2(new_n758), .A3(new_n764), .ZN(new_n765));
  NOR4_X1   g579(.A1(new_n763), .A2(new_n765), .A3(new_n602), .A4(new_n657), .ZN(new_n766));
  OR2_X1    g580(.A1(new_n766), .A2(KEYINPUT44), .ZN(new_n767));
  INV_X1    g581(.A(KEYINPUT45), .ZN(new_n768));
  NAND3_X1  g582(.A1(new_n448), .A2(new_n768), .A3(new_n452), .ZN(new_n769));
  OR2_X1    g583(.A1(new_n734), .A2(new_n768), .ZN(new_n770));
  NAND3_X1  g584(.A1(new_n769), .A2(G469), .A3(new_n770), .ZN(new_n771));
  NAND3_X1  g585(.A1(new_n771), .A2(KEYINPUT46), .A3(new_n733), .ZN(new_n772));
  AND3_X1   g586(.A1(new_n772), .A2(KEYINPUT110), .A3(new_n444), .ZN(new_n773));
  AOI21_X1  g587(.A(KEYINPUT110), .B1(new_n772), .B2(new_n444), .ZN(new_n774));
  AOI21_X1  g588(.A(KEYINPUT46), .B1(new_n771), .B2(new_n733), .ZN(new_n775));
  NOR3_X1   g589(.A1(new_n773), .A2(new_n774), .A3(new_n775), .ZN(new_n776));
  NOR3_X1   g590(.A1(new_n776), .A2(new_n694), .A3(new_n670), .ZN(new_n777));
  NAND2_X1  g591(.A1(new_n766), .A2(KEYINPUT44), .ZN(new_n778));
  XNOR2_X1  g592(.A(new_n731), .B(KEYINPUT112), .ZN(new_n779));
  INV_X1    g593(.A(new_n779), .ZN(new_n780));
  NAND4_X1  g594(.A1(new_n767), .A2(new_n777), .A3(new_n778), .A4(new_n780), .ZN(new_n781));
  XNOR2_X1  g595(.A(new_n781), .B(G137), .ZN(G39));
  NAND2_X1  g596(.A1(new_n772), .A2(new_n444), .ZN(new_n783));
  INV_X1    g597(.A(KEYINPUT110), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  INV_X1    g599(.A(new_n775), .ZN(new_n786));
  NAND3_X1  g600(.A1(new_n772), .A2(KEYINPUT110), .A3(new_n444), .ZN(new_n787));
  NAND3_X1  g601(.A1(new_n785), .A2(new_n786), .A3(new_n787), .ZN(new_n788));
  XOR2_X1   g602(.A(KEYINPUT113), .B(KEYINPUT47), .Z(new_n789));
  INV_X1    g603(.A(new_n789), .ZN(new_n790));
  AND3_X1   g604(.A1(new_n788), .A2(new_n456), .A3(new_n790), .ZN(new_n791));
  NOR2_X1   g605(.A1(KEYINPUT113), .A2(KEYINPUT47), .ZN(new_n792));
  AOI21_X1  g606(.A(new_n792), .B1(new_n788), .B2(new_n456), .ZN(new_n793));
  NOR2_X1   g607(.A1(new_n791), .A2(new_n793), .ZN(new_n794));
  NOR3_X1   g608(.A1(new_n750), .A2(new_n320), .A3(new_n731), .ZN(new_n795));
  NAND3_X1  g609(.A1(new_n794), .A2(new_n391), .A3(new_n795), .ZN(new_n796));
  INV_X1    g610(.A(KEYINPUT114), .ZN(new_n797));
  OR2_X1    g611(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  NAND2_X1  g612(.A1(new_n796), .A2(new_n797), .ZN(new_n799));
  NAND2_X1  g613(.A1(new_n798), .A2(new_n799), .ZN(new_n800));
  XNOR2_X1  g614(.A(new_n800), .B(G140), .ZN(G42));
  INV_X1    g615(.A(KEYINPUT54), .ZN(new_n802));
  INV_X1    g616(.A(KEYINPUT53), .ZN(new_n803));
  NAND4_X1  g617(.A1(new_n705), .A2(new_n702), .A3(new_n708), .A4(new_n718), .ZN(new_n804));
  XNOR2_X1  g618(.A(new_n593), .B(KEYINPUT115), .ZN(new_n805));
  OAI21_X1  g619(.A(new_n621), .B1(new_n557), .B2(new_n805), .ZN(new_n806));
  NAND3_X1  g620(.A1(new_n603), .A2(new_n510), .A3(new_n806), .ZN(new_n807));
  NAND3_X1  g621(.A1(new_n807), .A2(new_n599), .A3(new_n651), .ZN(new_n808));
  NOR2_X1   g622(.A1(new_n804), .A2(new_n808), .ZN(new_n809));
  INV_X1    g623(.A(new_n731), .ZN(new_n810));
  NOR2_X1   g624(.A1(new_n557), .A2(new_n659), .ZN(new_n811));
  AND3_X1   g625(.A1(new_n656), .A2(new_n805), .A3(new_n811), .ZN(new_n812));
  AND4_X1   g626(.A1(new_n689), .A2(new_n716), .A3(new_n687), .A4(new_n737), .ZN(new_n813));
  OAI211_X1 g627(.A(new_n650), .B(new_n810), .C1(new_n812), .C2(new_n813), .ZN(new_n814));
  AND4_X1   g628(.A1(new_n754), .A2(new_n809), .A3(new_n814), .A4(new_n756), .ZN(new_n815));
  INV_X1    g629(.A(KEYINPUT52), .ZN(new_n816));
  INV_X1    g630(.A(new_n677), .ZN(new_n817));
  AOI21_X1  g631(.A(new_n736), .B1(new_n305), .B2(new_n817), .ZN(new_n818));
  NOR2_X1   g632(.A1(new_n627), .A2(new_n669), .ZN(new_n819));
  AND3_X1   g633(.A1(new_n819), .A2(new_n657), .A3(new_n663), .ZN(new_n820));
  AOI21_X1  g634(.A(new_n816), .B1(new_n818), .B2(new_n820), .ZN(new_n821));
  NAND4_X1  g635(.A1(new_n692), .A2(new_n821), .A3(new_n725), .A4(new_n667), .ZN(new_n822));
  INV_X1    g636(.A(KEYINPUT116), .ZN(new_n823));
  NAND2_X1  g637(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  NAND2_X1  g638(.A1(new_n818), .A2(new_n820), .ZN(new_n825));
  NAND4_X1  g639(.A1(new_n692), .A2(new_n725), .A3(new_n667), .A4(new_n825), .ZN(new_n826));
  XOR2_X1   g640(.A(KEYINPUT117), .B(KEYINPUT52), .Z(new_n827));
  NAND2_X1  g641(.A1(new_n826), .A2(new_n827), .ZN(new_n828));
  NAND3_X1  g642(.A1(new_n720), .A2(new_n650), .A3(new_n721), .ZN(new_n829));
  NOR2_X1   g643(.A1(new_n750), .A2(new_n829), .ZN(new_n830));
  AOI22_X1  g644(.A1(new_n830), .A2(new_n724), .B1(new_n656), .B2(new_n666), .ZN(new_n831));
  NAND4_X1  g645(.A1(new_n831), .A2(KEYINPUT116), .A3(new_n692), .A4(new_n821), .ZN(new_n832));
  NAND3_X1  g646(.A1(new_n824), .A2(new_n828), .A3(new_n832), .ZN(new_n833));
  AOI21_X1  g647(.A(new_n803), .B1(new_n815), .B2(new_n833), .ZN(new_n834));
  NAND4_X1  g648(.A1(new_n754), .A2(new_n809), .A3(new_n814), .A4(new_n756), .ZN(new_n835));
  AND3_X1   g649(.A1(new_n692), .A2(new_n725), .A3(new_n667), .ZN(new_n836));
  AOI22_X1  g650(.A1(new_n836), .A2(new_n821), .B1(new_n826), .B2(new_n816), .ZN(new_n837));
  NOR3_X1   g651(.A1(new_n835), .A2(new_n837), .A3(KEYINPUT53), .ZN(new_n838));
  OAI21_X1  g652(.A(new_n802), .B1(new_n834), .B2(new_n838), .ZN(new_n839));
  AND3_X1   g653(.A1(new_n824), .A2(new_n828), .A3(new_n832), .ZN(new_n840));
  OAI21_X1  g654(.A(new_n803), .B1(new_n840), .B2(new_n835), .ZN(new_n841));
  INV_X1    g655(.A(new_n837), .ZN(new_n842));
  NAND3_X1  g656(.A1(new_n815), .A2(new_n842), .A3(KEYINPUT53), .ZN(new_n843));
  AOI21_X1  g657(.A(new_n802), .B1(new_n841), .B2(new_n843), .ZN(new_n844));
  INV_X1    g658(.A(KEYINPUT118), .ZN(new_n845));
  OAI21_X1  g659(.A(new_n839), .B1(new_n844), .B2(new_n845), .ZN(new_n846));
  NOR2_X1   g660(.A1(KEYINPUT121), .A2(KEYINPUT51), .ZN(new_n847));
  INV_X1    g661(.A(new_n847), .ZN(new_n848));
  NOR2_X1   g662(.A1(new_n763), .A2(new_n765), .ZN(new_n849));
  AND4_X1   g663(.A1(new_n503), .A2(new_n729), .A3(new_n700), .A4(new_n730), .ZN(new_n850));
  AOI21_X1  g664(.A(KEYINPUT120), .B1(new_n849), .B2(new_n850), .ZN(new_n851));
  NAND2_X1  g665(.A1(new_n762), .A2(new_n620), .ZN(new_n852));
  NAND2_X1  g666(.A1(new_n852), .A2(KEYINPUT43), .ZN(new_n853));
  NAND3_X1  g667(.A1(new_n620), .A2(new_n758), .A3(new_n764), .ZN(new_n854));
  AND4_X1   g668(.A1(KEYINPUT120), .A2(new_n853), .A3(new_n850), .A4(new_n854), .ZN(new_n855));
  OAI21_X1  g669(.A(new_n722), .B1(new_n851), .B2(new_n855), .ZN(new_n856));
  NAND4_X1  g670(.A1(new_n849), .A2(new_n392), .A3(new_n503), .A4(new_n716), .ZN(new_n857));
  OAI211_X1 g671(.A(new_n622), .B(new_n700), .C1(new_n679), .C2(new_n680), .ZN(new_n858));
  XNOR2_X1  g672(.A(new_n858), .B(KEYINPUT119), .ZN(new_n859));
  OAI21_X1  g673(.A(KEYINPUT50), .B1(new_n857), .B2(new_n859), .ZN(new_n860));
  AND2_X1   g674(.A1(new_n678), .A2(new_n392), .ZN(new_n861));
  INV_X1    g675(.A(new_n620), .ZN(new_n862));
  NAND4_X1  g676(.A1(new_n861), .A2(new_n764), .A3(new_n862), .A4(new_n850), .ZN(new_n863));
  NAND3_X1  g677(.A1(new_n856), .A2(new_n860), .A3(new_n863), .ZN(new_n864));
  NOR2_X1   g678(.A1(new_n859), .A2(KEYINPUT50), .ZN(new_n865));
  INV_X1    g679(.A(new_n865), .ZN(new_n866));
  NAND2_X1  g680(.A1(new_n698), .A2(new_n699), .ZN(new_n867));
  INV_X1    g681(.A(new_n867), .ZN(new_n868));
  NOR2_X1   g682(.A1(new_n868), .A2(new_n457), .ZN(new_n869));
  INV_X1    g683(.A(new_n792), .ZN(new_n870));
  OAI21_X1  g684(.A(new_n870), .B1(new_n776), .B2(new_n694), .ZN(new_n871));
  NAND3_X1  g685(.A1(new_n788), .A2(new_n456), .A3(new_n790), .ZN(new_n872));
  AOI21_X1  g686(.A(new_n869), .B1(new_n871), .B2(new_n872), .ZN(new_n873));
  OAI21_X1  g687(.A(new_n866), .B1(new_n873), .B2(new_n779), .ZN(new_n874));
  INV_X1    g688(.A(new_n857), .ZN(new_n875));
  AOI21_X1  g689(.A(new_n864), .B1(new_n874), .B2(new_n875), .ZN(new_n876));
  AND2_X1   g690(.A1(KEYINPUT121), .A2(KEYINPUT51), .ZN(new_n877));
  OAI21_X1  g691(.A(new_n848), .B1(new_n876), .B2(new_n877), .ZN(new_n878));
  NOR2_X1   g692(.A1(new_n502), .A2(G953), .ZN(new_n879));
  NAND4_X1  g693(.A1(new_n861), .A2(new_n557), .A3(new_n620), .A4(new_n850), .ZN(new_n880));
  AND3_X1   g694(.A1(new_n856), .A2(new_n860), .A3(new_n863), .ZN(new_n881));
  INV_X1    g695(.A(new_n869), .ZN(new_n882));
  OAI21_X1  g696(.A(new_n882), .B1(new_n791), .B2(new_n793), .ZN(new_n883));
  AOI21_X1  g697(.A(new_n865), .B1(new_n883), .B2(new_n780), .ZN(new_n884));
  OAI21_X1  g698(.A(new_n881), .B1(new_n884), .B2(new_n857), .ZN(new_n885));
  NAND2_X1  g699(.A1(new_n885), .A2(new_n847), .ZN(new_n886));
  NAND4_X1  g700(.A1(new_n878), .A2(new_n879), .A3(new_n880), .A4(new_n886), .ZN(new_n887));
  NOR2_X1   g701(.A1(new_n851), .A2(new_n855), .ZN(new_n888));
  NAND2_X1  g702(.A1(new_n749), .A2(new_n392), .ZN(new_n889));
  NOR2_X1   g703(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  XNOR2_X1  g704(.A(new_n890), .B(KEYINPUT48), .ZN(new_n891));
  NOR3_X1   g705(.A1(new_n857), .A2(new_n627), .A3(new_n723), .ZN(new_n892));
  NOR3_X1   g706(.A1(new_n887), .A2(new_n891), .A3(new_n892), .ZN(new_n893));
  OAI21_X1  g707(.A(KEYINPUT53), .B1(new_n840), .B2(new_n835), .ZN(new_n894));
  NAND3_X1  g708(.A1(new_n815), .A2(new_n842), .A3(new_n803), .ZN(new_n895));
  AOI21_X1  g709(.A(KEYINPUT54), .B1(new_n894), .B2(new_n895), .ZN(new_n896));
  NAND2_X1  g710(.A1(new_n896), .A2(KEYINPUT118), .ZN(new_n897));
  NAND3_X1  g711(.A1(new_n846), .A2(new_n893), .A3(new_n897), .ZN(new_n898));
  NAND2_X1  g712(.A1(new_n502), .A2(new_n479), .ZN(new_n899));
  NAND2_X1  g713(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  INV_X1    g714(.A(new_n681), .ZN(new_n901));
  OAI21_X1  g715(.A(new_n457), .B1(new_n868), .B2(KEYINPUT49), .ZN(new_n902));
  NOR3_X1   g716(.A1(new_n901), .A2(new_n852), .A3(new_n902), .ZN(new_n903));
  NAND2_X1  g717(.A1(new_n868), .A2(KEYINPUT49), .ZN(new_n904));
  NAND4_X1  g718(.A1(new_n861), .A2(new_n903), .A3(new_n501), .A4(new_n904), .ZN(new_n905));
  NAND2_X1  g719(.A1(new_n900), .A2(new_n905), .ZN(G75));
  NAND4_X1  g720(.A1(new_n894), .A2(new_n895), .A3(G210), .A4(G902), .ZN(new_n907));
  INV_X1    g721(.A(KEYINPUT56), .ZN(new_n908));
  NAND3_X1  g722(.A1(new_n907), .A2(KEYINPUT122), .A3(new_n908), .ZN(new_n909));
  NAND2_X1  g723(.A1(new_n475), .A2(new_n483), .ZN(new_n910));
  XNOR2_X1  g724(.A(new_n910), .B(new_n481), .ZN(new_n911));
  XOR2_X1   g725(.A(new_n911), .B(KEYINPUT55), .Z(new_n912));
  AND2_X1   g726(.A1(new_n909), .A2(new_n912), .ZN(new_n913));
  NOR2_X1   g727(.A1(new_n909), .A2(new_n912), .ZN(new_n914));
  NOR2_X1   g728(.A1(new_n354), .A2(G952), .ZN(new_n915));
  NOR3_X1   g729(.A1(new_n913), .A2(new_n914), .A3(new_n915), .ZN(G51));
  NAND2_X1  g730(.A1(new_n733), .A2(KEYINPUT57), .ZN(new_n917));
  OR2_X1    g731(.A1(new_n733), .A2(KEYINPUT57), .ZN(new_n918));
  NOR3_X1   g732(.A1(new_n834), .A2(new_n838), .A3(new_n802), .ZN(new_n919));
  OAI211_X1 g733(.A(new_n917), .B(new_n918), .C1(new_n919), .C2(new_n896), .ZN(new_n920));
  NAND2_X1  g734(.A1(new_n920), .A2(new_n442), .ZN(new_n921));
  NOR3_X1   g735(.A1(new_n834), .A2(new_n838), .A3(new_n371), .ZN(new_n922));
  INV_X1    g736(.A(new_n771), .ZN(new_n923));
  NAND2_X1  g737(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  AOI21_X1  g738(.A(new_n915), .B1(new_n921), .B2(new_n924), .ZN(G54));
  NAND3_X1  g739(.A1(new_n922), .A2(KEYINPUT58), .A3(G475), .ZN(new_n926));
  NAND3_X1  g740(.A1(new_n926), .A2(new_n544), .A3(new_n538), .ZN(new_n927));
  INV_X1    g741(.A(new_n915), .ZN(new_n928));
  NAND2_X1  g742(.A1(new_n538), .A2(new_n544), .ZN(new_n929));
  NAND4_X1  g743(.A1(new_n922), .A2(KEYINPUT58), .A3(G475), .A4(new_n929), .ZN(new_n930));
  AND3_X1   g744(.A1(new_n927), .A2(new_n928), .A3(new_n930), .ZN(G60));
  NAND2_X1  g745(.A1(G478), .A2(G902), .ZN(new_n932));
  XOR2_X1   g746(.A(new_n932), .B(KEYINPUT59), .Z(new_n933));
  INV_X1    g747(.A(new_n933), .ZN(new_n934));
  OAI211_X1 g748(.A(new_n617), .B(new_n934), .C1(new_n919), .C2(new_n896), .ZN(new_n935));
  NAND2_X1  g749(.A1(new_n935), .A2(new_n928), .ZN(new_n936));
  AOI21_X1  g750(.A(KEYINPUT53), .B1(new_n815), .B2(new_n833), .ZN(new_n937));
  NOR3_X1   g751(.A1(new_n835), .A2(new_n837), .A3(new_n803), .ZN(new_n938));
  OAI21_X1  g752(.A(KEYINPUT54), .B1(new_n937), .B2(new_n938), .ZN(new_n939));
  AOI21_X1  g753(.A(new_n896), .B1(KEYINPUT118), .B2(new_n939), .ZN(new_n940));
  NOR2_X1   g754(.A1(new_n839), .A2(new_n845), .ZN(new_n941));
  OAI21_X1  g755(.A(new_n934), .B1(new_n940), .B2(new_n941), .ZN(new_n942));
  INV_X1    g756(.A(new_n617), .ZN(new_n943));
  AOI21_X1  g757(.A(new_n936), .B1(new_n942), .B2(new_n943), .ZN(G63));
  XNOR2_X1  g758(.A(new_n387), .B(KEYINPUT124), .ZN(new_n945));
  INV_X1    g759(.A(new_n945), .ZN(new_n946));
  NOR2_X1   g760(.A1(new_n834), .A2(new_n838), .ZN(new_n947));
  NAND2_X1  g761(.A1(G217), .A2(G902), .ZN(new_n948));
  XNOR2_X1  g762(.A(new_n948), .B(KEYINPUT123), .ZN(new_n949));
  XNOR2_X1  g763(.A(new_n949), .B(KEYINPUT60), .ZN(new_n950));
  AOI21_X1  g764(.A(new_n946), .B1(new_n947), .B2(new_n950), .ZN(new_n951));
  NAND4_X1  g765(.A1(new_n894), .A2(new_n895), .A3(new_n648), .A4(new_n950), .ZN(new_n952));
  NAND2_X1  g766(.A1(new_n952), .A2(new_n928), .ZN(new_n953));
  INV_X1    g767(.A(KEYINPUT61), .ZN(new_n954));
  OR3_X1    g768(.A1(new_n951), .A2(new_n953), .A3(new_n954), .ZN(new_n955));
  OAI21_X1  g769(.A(new_n954), .B1(new_n951), .B2(new_n953), .ZN(new_n956));
  NAND2_X1  g770(.A1(new_n955), .A2(new_n956), .ZN(G66));
  INV_X1    g771(.A(new_n478), .ZN(new_n958));
  OAI21_X1  g772(.A(G953), .B1(new_n506), .B2(new_n958), .ZN(new_n959));
  INV_X1    g773(.A(new_n354), .ZN(new_n960));
  OAI21_X1  g774(.A(new_n959), .B1(new_n809), .B2(new_n960), .ZN(new_n961));
  OAI21_X1  g775(.A(new_n910), .B1(G898), .B2(new_n354), .ZN(new_n962));
  XNOR2_X1  g776(.A(new_n961), .B(new_n962), .ZN(G69));
  XNOR2_X1  g777(.A(new_n288), .B(new_n534), .ZN(new_n964));
  NAND2_X1  g778(.A1(new_n836), .A2(new_n683), .ZN(new_n965));
  INV_X1    g779(.A(KEYINPUT62), .ZN(new_n966));
  NAND2_X1  g780(.A1(new_n965), .A2(new_n966), .ZN(new_n967));
  NAND3_X1  g781(.A1(new_n836), .A2(KEYINPUT62), .A3(new_n683), .ZN(new_n968));
  NAND2_X1  g782(.A1(new_n967), .A2(new_n968), .ZN(new_n969));
  NAND3_X1  g783(.A1(new_n732), .A2(new_n671), .A3(new_n806), .ZN(new_n970));
  NAND4_X1  g784(.A1(new_n800), .A2(new_n969), .A3(new_n781), .A4(new_n970), .ZN(new_n971));
  INV_X1    g785(.A(new_n971), .ZN(new_n972));
  OAI21_X1  g786(.A(new_n964), .B1(new_n972), .B2(new_n960), .ZN(new_n973));
  NOR2_X1   g787(.A1(new_n354), .A2(G900), .ZN(new_n974));
  XNOR2_X1  g788(.A(new_n974), .B(KEYINPUT125), .ZN(new_n975));
  INV_X1    g789(.A(new_n975), .ZN(new_n976));
  INV_X1    g790(.A(new_n781), .ZN(new_n977));
  AOI21_X1  g791(.A(new_n977), .B1(new_n798), .B2(new_n799), .ZN(new_n978));
  NAND4_X1  g792(.A1(new_n777), .A2(new_n749), .A3(new_n392), .A4(new_n819), .ZN(new_n979));
  AND3_X1   g793(.A1(new_n754), .A2(new_n756), .A3(new_n836), .ZN(new_n980));
  NAND3_X1  g794(.A1(new_n978), .A2(new_n979), .A3(new_n980), .ZN(new_n981));
  AOI21_X1  g795(.A(new_n976), .B1(new_n981), .B2(new_n354), .ZN(new_n982));
  OAI21_X1  g796(.A(new_n973), .B1(new_n964), .B2(new_n982), .ZN(new_n983));
  AOI21_X1  g797(.A(new_n354), .B1(G227), .B2(G900), .ZN(new_n984));
  NAND2_X1  g798(.A1(new_n983), .A2(new_n984), .ZN(new_n985));
  INV_X1    g799(.A(new_n984), .ZN(new_n986));
  OAI211_X1 g800(.A(new_n973), .B(new_n986), .C1(new_n964), .C2(new_n982), .ZN(new_n987));
  NAND2_X1  g801(.A1(new_n985), .A2(new_n987), .ZN(G72));
  NAND4_X1  g802(.A1(new_n978), .A2(new_n809), .A3(new_n969), .A4(new_n970), .ZN(new_n989));
  XNOR2_X1  g803(.A(KEYINPUT126), .B(KEYINPUT63), .ZN(new_n990));
  NAND2_X1  g804(.A1(G472), .A2(G902), .ZN(new_n991));
  XNOR2_X1  g805(.A(new_n990), .B(new_n991), .ZN(new_n992));
  NAND3_X1  g806(.A1(new_n989), .A2(KEYINPUT127), .A3(new_n992), .ZN(new_n993));
  NAND2_X1  g807(.A1(new_n993), .A2(new_n195), .ZN(new_n994));
  INV_X1    g808(.A(new_n307), .ZN(new_n995));
  AOI21_X1  g809(.A(KEYINPUT127), .B1(new_n989), .B2(new_n992), .ZN(new_n996));
  NOR3_X1   g810(.A1(new_n994), .A2(new_n995), .A3(new_n996), .ZN(new_n997));
  INV_X1    g811(.A(new_n809), .ZN(new_n998));
  OAI21_X1  g812(.A(new_n992), .B1(new_n981), .B2(new_n998), .ZN(new_n999));
  NAND3_X1  g813(.A1(new_n999), .A2(new_n995), .A3(new_n308), .ZN(new_n1000));
  OAI21_X1  g814(.A(new_n309), .B1(new_n283), .B2(new_n278), .ZN(new_n1001));
  OAI211_X1 g815(.A(new_n992), .B(new_n1001), .C1(new_n937), .C2(new_n938), .ZN(new_n1002));
  NAND3_X1  g816(.A1(new_n1000), .A2(new_n928), .A3(new_n1002), .ZN(new_n1003));
  NOR2_X1   g817(.A1(new_n997), .A2(new_n1003), .ZN(G57));
endmodule


