//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 1 0 1 0 0 0 1 0 0 0 1 0 1 1 1 1 0 0 0 0 1 1 1 0 1 1 0 1 0 0 1 0 0 1 0 1 0 0 0 1 1 1 1 0 0 0 1 1 1 0 0 0 1 0 1 0 1 1 1 1 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:25:14 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n611, new_n612, new_n613, new_n614, new_n615,
    new_n617, new_n618, new_n619, new_n620, new_n621, new_n622, new_n623,
    new_n624, new_n625, new_n627, new_n628, new_n629, new_n630, new_n631,
    new_n632, new_n633, new_n634, new_n635, new_n636, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n655, new_n656, new_n657, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n669, new_n670,
    new_n671, new_n673, new_n674, new_n675, new_n676, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n719, new_n720, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n870,
    new_n871, new_n872, new_n873, new_n874, new_n875, new_n876, new_n877,
    new_n878, new_n880, new_n881, new_n882, new_n883, new_n884, new_n885,
    new_n886, new_n887, new_n888, new_n889, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n906, new_n907, new_n908,
    new_n909, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n935, new_n936, new_n937, new_n938,
    new_n939, new_n940, new_n941, new_n942, new_n943, new_n944, new_n945,
    new_n946, new_n947, new_n948, new_n949, new_n950, new_n951, new_n952,
    new_n953, new_n954;
  INV_X1    g000(.A(G104), .ZN(new_n187));
  NOR2_X1   g001(.A1(new_n187), .A2(KEYINPUT3), .ZN(new_n188));
  INV_X1    g002(.A(KEYINPUT78), .ZN(new_n189));
  NOR2_X1   g003(.A1(new_n189), .A2(G107), .ZN(new_n190));
  INV_X1    g004(.A(G107), .ZN(new_n191));
  NOR2_X1   g005(.A1(new_n191), .A2(KEYINPUT78), .ZN(new_n192));
  OAI21_X1  g006(.A(new_n188), .B1(new_n190), .B2(new_n192), .ZN(new_n193));
  NOR2_X1   g007(.A1(new_n191), .A2(G104), .ZN(new_n194));
  INV_X1    g008(.A(new_n194), .ZN(new_n195));
  OAI21_X1  g009(.A(KEYINPUT3), .B1(new_n187), .B2(G107), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n196), .A2(KEYINPUT77), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n191), .A2(G104), .ZN(new_n198));
  INV_X1    g012(.A(KEYINPUT77), .ZN(new_n199));
  NAND3_X1  g013(.A1(new_n198), .A2(new_n199), .A3(KEYINPUT3), .ZN(new_n200));
  NAND4_X1  g014(.A1(new_n193), .A2(new_n195), .A3(new_n197), .A4(new_n200), .ZN(new_n201));
  INV_X1    g015(.A(KEYINPUT4), .ZN(new_n202));
  NAND3_X1  g016(.A1(new_n201), .A2(new_n202), .A3(G101), .ZN(new_n203));
  NOR2_X1   g017(.A1(KEYINPUT2), .A2(G113), .ZN(new_n204));
  NAND2_X1  g018(.A1(KEYINPUT2), .A2(G113), .ZN(new_n205));
  INV_X1    g019(.A(KEYINPUT67), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  NAND3_X1  g021(.A1(KEYINPUT67), .A2(KEYINPUT2), .A3(G113), .ZN(new_n208));
  AOI21_X1  g022(.A(new_n204), .B1(new_n207), .B2(new_n208), .ZN(new_n209));
  XNOR2_X1  g023(.A(G116), .B(G119), .ZN(new_n210));
  XNOR2_X1  g024(.A(new_n209), .B(new_n210), .ZN(new_n211));
  XNOR2_X1  g025(.A(KEYINPUT79), .B(G101), .ZN(new_n212));
  OAI21_X1  g026(.A(KEYINPUT4), .B1(new_n201), .B2(new_n212), .ZN(new_n213));
  INV_X1    g027(.A(G101), .ZN(new_n214));
  AND2_X1   g028(.A1(new_n197), .A2(new_n200), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n191), .A2(KEYINPUT78), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n189), .A2(G107), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  AOI21_X1  g032(.A(new_n194), .B1(new_n218), .B2(new_n188), .ZN(new_n219));
  AOI21_X1  g033(.A(new_n214), .B1(new_n215), .B2(new_n219), .ZN(new_n220));
  OAI211_X1 g034(.A(new_n203), .B(new_n211), .C1(new_n213), .C2(new_n220), .ZN(new_n221));
  XNOR2_X1  g035(.A(KEYINPUT78), .B(G107), .ZN(new_n222));
  INV_X1    g036(.A(new_n188), .ZN(new_n223));
  OAI21_X1  g037(.A(new_n195), .B1(new_n222), .B2(new_n223), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n197), .A2(new_n200), .ZN(new_n225));
  NOR2_X1   g039(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  INV_X1    g040(.A(new_n212), .ZN(new_n227));
  OAI21_X1  g041(.A(new_n198), .B1(new_n218), .B2(G104), .ZN(new_n228));
  AOI22_X1  g042(.A1(new_n226), .A2(new_n227), .B1(G101), .B2(new_n228), .ZN(new_n229));
  AND2_X1   g043(.A1(new_n209), .A2(new_n210), .ZN(new_n230));
  INV_X1    g044(.A(G116), .ZN(new_n231));
  NOR3_X1   g045(.A1(new_n231), .A2(KEYINPUT5), .A3(G119), .ZN(new_n232));
  AOI21_X1  g046(.A(new_n232), .B1(new_n210), .B2(KEYINPUT5), .ZN(new_n233));
  AOI21_X1  g047(.A(new_n230), .B1(G113), .B2(new_n233), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n229), .A2(new_n234), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n221), .A2(new_n235), .ZN(new_n236));
  XOR2_X1   g050(.A(G110), .B(G122), .Z(new_n237));
  NAND2_X1  g051(.A1(new_n236), .A2(new_n237), .ZN(new_n238));
  INV_X1    g052(.A(new_n237), .ZN(new_n239));
  NAND3_X1  g053(.A1(new_n221), .A2(new_n235), .A3(new_n239), .ZN(new_n240));
  NAND3_X1  g054(.A1(new_n238), .A2(KEYINPUT6), .A3(new_n240), .ZN(new_n241));
  INV_X1    g055(.A(G146), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n242), .A2(G143), .ZN(new_n243));
  INV_X1    g057(.A(G143), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n244), .A2(G146), .ZN(new_n245));
  NAND4_X1  g059(.A1(new_n243), .A2(new_n245), .A3(KEYINPUT0), .A4(G128), .ZN(new_n246));
  INV_X1    g060(.A(KEYINPUT64), .ZN(new_n247));
  OAI21_X1  g061(.A(new_n247), .B1(new_n242), .B2(G143), .ZN(new_n248));
  NAND3_X1  g062(.A1(new_n244), .A2(KEYINPUT64), .A3(G146), .ZN(new_n249));
  AOI22_X1  g063(.A1(new_n248), .A2(new_n249), .B1(G143), .B2(new_n242), .ZN(new_n250));
  XNOR2_X1  g064(.A(KEYINPUT0), .B(G128), .ZN(new_n251));
  OAI21_X1  g065(.A(new_n246), .B1(new_n250), .B2(new_n251), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n252), .A2(G125), .ZN(new_n253));
  INV_X1    g067(.A(KEYINPUT1), .ZN(new_n254));
  NAND4_X1  g068(.A1(new_n243), .A2(new_n245), .A3(new_n254), .A4(G128), .ZN(new_n255));
  INV_X1    g069(.A(G128), .ZN(new_n256));
  AOI21_X1  g070(.A(new_n256), .B1(new_n243), .B2(KEYINPUT1), .ZN(new_n257));
  OAI21_X1  g071(.A(new_n255), .B1(new_n250), .B2(new_n257), .ZN(new_n258));
  OAI21_X1  g072(.A(new_n253), .B1(G125), .B2(new_n258), .ZN(new_n259));
  INV_X1    g073(.A(G953), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n260), .A2(G224), .ZN(new_n261));
  XOR2_X1   g075(.A(new_n259), .B(new_n261), .Z(new_n262));
  INV_X1    g076(.A(KEYINPUT6), .ZN(new_n263));
  NAND3_X1  g077(.A1(new_n236), .A2(new_n263), .A3(new_n237), .ZN(new_n264));
  NAND3_X1  g078(.A1(new_n241), .A2(new_n262), .A3(new_n264), .ZN(new_n265));
  INV_X1    g079(.A(G902), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n261), .A2(KEYINPUT7), .ZN(new_n267));
  XOR2_X1   g081(.A(new_n259), .B(new_n267), .Z(new_n268));
  NAND2_X1  g082(.A1(new_n228), .A2(G101), .ZN(new_n269));
  OAI21_X1  g083(.A(new_n269), .B1(new_n201), .B2(new_n212), .ZN(new_n270));
  XNOR2_X1  g084(.A(new_n234), .B(new_n270), .ZN(new_n271));
  XNOR2_X1  g085(.A(new_n237), .B(KEYINPUT8), .ZN(new_n272));
  OAI211_X1 g086(.A(new_n268), .B(new_n240), .C1(new_n271), .C2(new_n272), .ZN(new_n273));
  NAND3_X1  g087(.A1(new_n265), .A2(new_n266), .A3(new_n273), .ZN(new_n274));
  OAI21_X1  g088(.A(G210), .B1(G237), .B2(G902), .ZN(new_n275));
  INV_X1    g089(.A(new_n275), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n274), .A2(new_n276), .ZN(new_n277));
  INV_X1    g091(.A(KEYINPUT84), .ZN(new_n278));
  NAND4_X1  g092(.A1(new_n265), .A2(new_n266), .A3(new_n275), .A4(new_n273), .ZN(new_n279));
  NAND3_X1  g093(.A1(new_n277), .A2(new_n278), .A3(new_n279), .ZN(new_n280));
  OR2_X1    g094(.A1(new_n279), .A2(new_n278), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  XOR2_X1   g096(.A(KEYINPUT21), .B(G898), .Z(new_n283));
  INV_X1    g097(.A(new_n283), .ZN(new_n284));
  NAND2_X1  g098(.A1(G234), .A2(G237), .ZN(new_n285));
  AND3_X1   g099(.A1(new_n285), .A2(G902), .A3(G953), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n284), .A2(new_n286), .ZN(new_n287));
  XNOR2_X1  g101(.A(KEYINPUT95), .B(G952), .ZN(new_n288));
  NOR2_X1   g102(.A1(new_n288), .A2(G953), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n289), .A2(new_n285), .ZN(new_n290));
  AND2_X1   g104(.A1(new_n287), .A2(new_n290), .ZN(new_n291));
  OAI21_X1  g105(.A(G214), .B1(G237), .B2(G902), .ZN(new_n292));
  INV_X1    g106(.A(new_n292), .ZN(new_n293));
  OR2_X1    g107(.A1(new_n291), .A2(new_n293), .ZN(new_n294));
  XOR2_X1   g108(.A(G113), .B(G122), .Z(new_n295));
  XNOR2_X1  g109(.A(new_n295), .B(KEYINPUT90), .ZN(new_n296));
  XNOR2_X1  g110(.A(new_n296), .B(G104), .ZN(new_n297));
  INV_X1    g111(.A(G140), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n298), .A2(G125), .ZN(new_n299));
  INV_X1    g113(.A(G125), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n300), .A2(G140), .ZN(new_n301));
  NAND3_X1  g115(.A1(new_n299), .A2(new_n301), .A3(KEYINPUT72), .ZN(new_n302));
  OR3_X1    g116(.A1(new_n300), .A2(KEYINPUT72), .A3(G140), .ZN(new_n303));
  NAND3_X1  g117(.A1(new_n302), .A2(new_n303), .A3(G146), .ZN(new_n304));
  XNOR2_X1  g118(.A(G125), .B(G140), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n305), .A2(new_n242), .ZN(new_n306));
  AND3_X1   g120(.A1(new_n304), .A2(KEYINPUT86), .A3(new_n306), .ZN(new_n307));
  NOR2_X1   g121(.A1(new_n304), .A2(KEYINPUT86), .ZN(new_n308));
  OAI21_X1  g122(.A(KEYINPUT87), .B1(new_n307), .B2(new_n308), .ZN(new_n309));
  INV_X1    g123(.A(G237), .ZN(new_n310));
  NAND3_X1  g124(.A1(new_n310), .A2(new_n260), .A3(G214), .ZN(new_n311));
  XNOR2_X1  g125(.A(new_n311), .B(new_n244), .ZN(new_n312));
  NAND2_X1  g126(.A1(KEYINPUT18), .A2(G131), .ZN(new_n313));
  OAI21_X1  g127(.A(KEYINPUT88), .B1(new_n313), .B2(KEYINPUT85), .ZN(new_n314));
  OR2_X1    g128(.A1(new_n312), .A2(new_n314), .ZN(new_n315));
  NAND3_X1  g129(.A1(new_n304), .A2(KEYINPUT86), .A3(new_n306), .ZN(new_n316));
  INV_X1    g130(.A(KEYINPUT87), .ZN(new_n317));
  OAI211_X1 g131(.A(new_n316), .B(new_n317), .C1(KEYINPUT86), .C2(new_n304), .ZN(new_n318));
  NOR2_X1   g132(.A1(new_n313), .A2(KEYINPUT88), .ZN(new_n319));
  OAI21_X1  g133(.A(new_n314), .B1(new_n312), .B2(new_n319), .ZN(new_n320));
  NAND4_X1  g134(.A1(new_n309), .A2(new_n315), .A3(new_n318), .A4(new_n320), .ZN(new_n321));
  NOR2_X1   g135(.A1(new_n299), .A2(KEYINPUT16), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n302), .A2(new_n303), .ZN(new_n323));
  AOI21_X1  g137(.A(new_n322), .B1(new_n323), .B2(KEYINPUT16), .ZN(new_n324));
  NOR2_X1   g138(.A1(new_n324), .A2(G146), .ZN(new_n325));
  INV_X1    g139(.A(new_n325), .ZN(new_n326));
  INV_X1    g140(.A(G131), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n327), .A2(KEYINPUT66), .ZN(new_n328));
  INV_X1    g142(.A(KEYINPUT66), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n329), .A2(G131), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n328), .A2(new_n330), .ZN(new_n331));
  INV_X1    g145(.A(new_n331), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n312), .A2(new_n332), .ZN(new_n333));
  XNOR2_X1  g147(.A(new_n311), .B(G143), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n334), .A2(new_n331), .ZN(new_n335));
  INV_X1    g149(.A(KEYINPUT17), .ZN(new_n336));
  NAND3_X1  g150(.A1(new_n333), .A2(new_n335), .A3(new_n336), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n324), .A2(G146), .ZN(new_n338));
  NAND3_X1  g152(.A1(new_n312), .A2(KEYINPUT17), .A3(new_n332), .ZN(new_n339));
  NAND4_X1  g153(.A1(new_n326), .A2(new_n337), .A3(new_n338), .A4(new_n339), .ZN(new_n340));
  AOI21_X1  g154(.A(new_n297), .B1(new_n321), .B2(new_n340), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n341), .A2(KEYINPUT92), .ZN(new_n342));
  NAND3_X1  g156(.A1(new_n321), .A2(new_n340), .A3(new_n297), .ZN(new_n343));
  INV_X1    g157(.A(KEYINPUT92), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  OAI211_X1 g159(.A(new_n342), .B(new_n266), .C1(new_n345), .C2(new_n341), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n346), .A2(G475), .ZN(new_n347));
  INV_X1    g161(.A(KEYINPUT89), .ZN(new_n348));
  AOI211_X1 g162(.A(new_n242), .B(new_n322), .C1(new_n323), .C2(KEYINPUT16), .ZN(new_n349));
  NAND3_X1  g163(.A1(new_n302), .A2(new_n303), .A3(KEYINPUT19), .ZN(new_n350));
  INV_X1    g164(.A(KEYINPUT19), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n305), .A2(new_n351), .ZN(new_n352));
  AND3_X1   g166(.A1(new_n350), .A2(new_n242), .A3(new_n352), .ZN(new_n353));
  OAI21_X1  g167(.A(new_n348), .B1(new_n349), .B2(new_n353), .ZN(new_n354));
  NAND3_X1  g168(.A1(new_n350), .A2(new_n242), .A3(new_n352), .ZN(new_n355));
  NAND3_X1  g169(.A1(new_n338), .A2(KEYINPUT89), .A3(new_n355), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n333), .A2(new_n335), .ZN(new_n357));
  NAND3_X1  g171(.A1(new_n354), .A2(new_n356), .A3(new_n357), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n358), .A2(new_n321), .ZN(new_n359));
  INV_X1    g173(.A(new_n297), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n359), .A2(new_n360), .ZN(new_n361));
  AOI21_X1  g175(.A(G475), .B1(new_n361), .B2(new_n343), .ZN(new_n362));
  INV_X1    g176(.A(KEYINPUT91), .ZN(new_n363));
  AND3_X1   g177(.A1(new_n321), .A2(new_n340), .A3(new_n297), .ZN(new_n364));
  AOI21_X1  g178(.A(new_n297), .B1(new_n358), .B2(new_n321), .ZN(new_n365));
  OAI21_X1  g179(.A(new_n363), .B1(new_n364), .B2(new_n365), .ZN(new_n366));
  INV_X1    g180(.A(KEYINPUT20), .ZN(new_n367));
  NAND4_X1  g181(.A1(new_n362), .A2(new_n366), .A3(new_n367), .A4(new_n266), .ZN(new_n368));
  INV_X1    g182(.A(new_n368), .ZN(new_n369));
  AOI22_X1  g183(.A1(new_n266), .A2(new_n362), .B1(new_n366), .B2(new_n367), .ZN(new_n370));
  OAI21_X1  g184(.A(new_n347), .B1(new_n369), .B2(new_n370), .ZN(new_n371));
  XNOR2_X1  g185(.A(KEYINPUT9), .B(G234), .ZN(new_n372));
  INV_X1    g186(.A(G217), .ZN(new_n373));
  NOR3_X1   g187(.A1(new_n372), .A2(new_n373), .A3(G953), .ZN(new_n374));
  XNOR2_X1  g188(.A(G128), .B(G143), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n375), .A2(KEYINPUT13), .ZN(new_n376));
  OR3_X1    g190(.A1(new_n256), .A2(KEYINPUT13), .A3(G143), .ZN(new_n377));
  NAND3_X1  g191(.A1(new_n376), .A2(G134), .A3(new_n377), .ZN(new_n378));
  INV_X1    g192(.A(G134), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n375), .A2(new_n379), .ZN(new_n380));
  XNOR2_X1  g194(.A(G116), .B(G122), .ZN(new_n381));
  NOR2_X1   g195(.A1(new_n218), .A2(new_n381), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n218), .A2(new_n381), .ZN(new_n383));
  INV_X1    g197(.A(new_n383), .ZN(new_n384));
  OAI211_X1 g198(.A(new_n378), .B(new_n380), .C1(new_n382), .C2(new_n384), .ZN(new_n385));
  XNOR2_X1  g199(.A(new_n375), .B(new_n379), .ZN(new_n386));
  INV_X1    g200(.A(KEYINPUT14), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n381), .A2(new_n387), .ZN(new_n388));
  NAND3_X1  g202(.A1(new_n231), .A2(KEYINPUT14), .A3(G122), .ZN(new_n389));
  NAND3_X1  g203(.A1(new_n388), .A2(G107), .A3(new_n389), .ZN(new_n390));
  NAND3_X1  g204(.A1(new_n386), .A2(new_n383), .A3(new_n390), .ZN(new_n391));
  AOI21_X1  g205(.A(new_n374), .B1(new_n385), .B2(new_n391), .ZN(new_n392));
  INV_X1    g206(.A(new_n392), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n393), .A2(KEYINPUT94), .ZN(new_n394));
  NAND3_X1  g208(.A1(new_n385), .A2(new_n391), .A3(new_n374), .ZN(new_n395));
  INV_X1    g209(.A(KEYINPUT93), .ZN(new_n396));
  OR2_X1    g210(.A1(new_n395), .A2(new_n396), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n395), .A2(new_n396), .ZN(new_n398));
  INV_X1    g212(.A(KEYINPUT94), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n392), .A2(new_n399), .ZN(new_n400));
  NAND4_X1  g214(.A1(new_n394), .A2(new_n397), .A3(new_n398), .A4(new_n400), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n401), .A2(new_n266), .ZN(new_n402));
  INV_X1    g216(.A(KEYINPUT15), .ZN(new_n403));
  NAND3_X1  g217(.A1(new_n402), .A2(new_n403), .A3(G478), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n403), .A2(G478), .ZN(new_n405));
  NAND3_X1  g219(.A1(new_n401), .A2(new_n266), .A3(new_n405), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n404), .A2(new_n406), .ZN(new_n407));
  NOR4_X1   g221(.A1(new_n282), .A2(new_n294), .A3(new_n371), .A4(new_n407), .ZN(new_n408));
  INV_X1    g222(.A(G221), .ZN(new_n409));
  INV_X1    g223(.A(new_n372), .ZN(new_n410));
  AOI21_X1  g224(.A(new_n409), .B1(new_n410), .B2(new_n266), .ZN(new_n411));
  INV_X1    g225(.A(G469), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n248), .A2(new_n249), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n413), .A2(new_n243), .ZN(new_n414));
  INV_X1    g228(.A(new_n251), .ZN(new_n415));
  AND3_X1   g229(.A1(new_n243), .A2(new_n245), .A3(G128), .ZN(new_n416));
  AOI22_X1  g230(.A1(new_n414), .A2(new_n415), .B1(new_n416), .B2(KEYINPUT0), .ZN(new_n417));
  OAI211_X1 g231(.A(new_n417), .B(new_n203), .C1(new_n213), .C2(new_n220), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n243), .A2(new_n245), .ZN(new_n419));
  OAI211_X1 g233(.A(KEYINPUT80), .B(KEYINPUT1), .C1(new_n244), .C2(G146), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n420), .A2(G128), .ZN(new_n421));
  AOI21_X1  g235(.A(KEYINPUT80), .B1(new_n243), .B2(KEYINPUT1), .ZN(new_n422));
  OAI21_X1  g236(.A(new_n419), .B1(new_n421), .B2(new_n422), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n423), .A2(new_n255), .ZN(new_n424));
  NAND4_X1  g238(.A1(new_n219), .A2(new_n227), .A3(new_n197), .A4(new_n200), .ZN(new_n425));
  NAND3_X1  g239(.A1(new_n424), .A2(new_n425), .A3(new_n269), .ZN(new_n426));
  INV_X1    g240(.A(KEYINPUT10), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n426), .A2(new_n427), .ZN(new_n428));
  INV_X1    g242(.A(KEYINPUT11), .ZN(new_n429));
  OAI21_X1  g243(.A(new_n429), .B1(new_n379), .B2(G137), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n379), .A2(G137), .ZN(new_n431));
  INV_X1    g245(.A(G137), .ZN(new_n432));
  NAND3_X1  g246(.A1(new_n432), .A2(KEYINPUT11), .A3(G134), .ZN(new_n433));
  NAND3_X1  g247(.A1(new_n430), .A2(new_n431), .A3(new_n433), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n434), .A2(G131), .ZN(new_n435));
  NAND4_X1  g249(.A1(new_n331), .A2(new_n431), .A3(new_n433), .A4(new_n430), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n435), .A2(new_n436), .ZN(new_n437));
  INV_X1    g251(.A(new_n437), .ZN(new_n438));
  NAND4_X1  g252(.A1(new_n425), .A2(KEYINPUT10), .A3(new_n269), .A4(new_n258), .ZN(new_n439));
  NAND4_X1  g253(.A1(new_n418), .A2(new_n428), .A3(new_n438), .A4(new_n439), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n440), .A2(KEYINPUT81), .ZN(new_n441));
  INV_X1    g255(.A(new_n258), .ZN(new_n442));
  NOR2_X1   g256(.A1(new_n442), .A2(new_n427), .ZN(new_n443));
  AOI22_X1  g257(.A1(new_n229), .A2(new_n443), .B1(new_n426), .B2(new_n427), .ZN(new_n444));
  INV_X1    g258(.A(KEYINPUT81), .ZN(new_n445));
  NAND4_X1  g259(.A1(new_n444), .A2(new_n445), .A3(new_n438), .A4(new_n418), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n441), .A2(new_n446), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n270), .A2(new_n442), .ZN(new_n448));
  AOI21_X1  g262(.A(new_n438), .B1(new_n448), .B2(new_n426), .ZN(new_n449));
  XNOR2_X1  g263(.A(new_n449), .B(KEYINPUT12), .ZN(new_n450));
  XNOR2_X1  g264(.A(G110), .B(G140), .ZN(new_n451));
  XNOR2_X1  g265(.A(new_n451), .B(KEYINPUT76), .ZN(new_n452));
  AND2_X1   g266(.A1(new_n260), .A2(G227), .ZN(new_n453));
  XNOR2_X1  g267(.A(new_n452), .B(new_n453), .ZN(new_n454));
  INV_X1    g268(.A(new_n454), .ZN(new_n455));
  AND3_X1   g269(.A1(new_n447), .A2(new_n450), .A3(new_n455), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n444), .A2(new_n418), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n457), .A2(new_n437), .ZN(new_n458));
  AOI21_X1  g272(.A(new_n455), .B1(new_n447), .B2(new_n458), .ZN(new_n459));
  OAI211_X1 g273(.A(new_n412), .B(new_n266), .C1(new_n456), .C2(new_n459), .ZN(new_n460));
  NOR2_X1   g274(.A1(new_n412), .A2(new_n266), .ZN(new_n461));
  INV_X1    g275(.A(new_n461), .ZN(new_n462));
  AND2_X1   g276(.A1(new_n460), .A2(new_n462), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n447), .A2(new_n450), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n464), .A2(KEYINPUT82), .ZN(new_n465));
  INV_X1    g279(.A(KEYINPUT82), .ZN(new_n466));
  NAND3_X1  g280(.A1(new_n447), .A2(new_n450), .A3(new_n466), .ZN(new_n467));
  NAND3_X1  g281(.A1(new_n465), .A2(new_n454), .A3(new_n467), .ZN(new_n468));
  AOI21_X1  g282(.A(new_n454), .B1(new_n441), .B2(new_n446), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n469), .A2(new_n458), .ZN(new_n470));
  NAND3_X1  g284(.A1(new_n468), .A2(G469), .A3(new_n470), .ZN(new_n471));
  AOI211_X1 g285(.A(KEYINPUT83), .B(new_n411), .C1(new_n463), .C2(new_n471), .ZN(new_n472));
  INV_X1    g286(.A(KEYINPUT83), .ZN(new_n473));
  NAND3_X1  g287(.A1(new_n471), .A2(new_n460), .A3(new_n462), .ZN(new_n474));
  INV_X1    g288(.A(new_n411), .ZN(new_n475));
  AOI21_X1  g289(.A(new_n473), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  OAI21_X1  g290(.A(new_n408), .B1(new_n472), .B2(new_n476), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n477), .A2(KEYINPUT96), .ZN(new_n478));
  INV_X1    g292(.A(KEYINPUT96), .ZN(new_n479));
  OAI211_X1 g293(.A(new_n408), .B(new_n479), .C1(new_n472), .C2(new_n476), .ZN(new_n480));
  INV_X1    g294(.A(KEYINPUT25), .ZN(new_n481));
  INV_X1    g295(.A(G119), .ZN(new_n482));
  OAI21_X1  g296(.A(KEYINPUT23), .B1(new_n482), .B2(G128), .ZN(new_n483));
  INV_X1    g297(.A(KEYINPUT23), .ZN(new_n484));
  NAND3_X1  g298(.A1(new_n484), .A2(new_n256), .A3(G119), .ZN(new_n485));
  AOI22_X1  g299(.A1(new_n483), .A2(new_n485), .B1(new_n482), .B2(G128), .ZN(new_n486));
  INV_X1    g300(.A(new_n486), .ZN(new_n487));
  NAND3_X1  g301(.A1(new_n487), .A2(KEYINPUT71), .A3(G110), .ZN(new_n488));
  INV_X1    g302(.A(KEYINPUT71), .ZN(new_n489));
  INV_X1    g303(.A(G110), .ZN(new_n490));
  OAI21_X1  g304(.A(new_n489), .B1(new_n486), .B2(new_n490), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n488), .A2(new_n491), .ZN(new_n492));
  XOR2_X1   g306(.A(G119), .B(G128), .Z(new_n493));
  INV_X1    g307(.A(KEYINPUT70), .ZN(new_n494));
  XNOR2_X1  g308(.A(KEYINPUT24), .B(G110), .ZN(new_n495));
  OR3_X1    g309(.A1(new_n493), .A2(new_n494), .A3(new_n495), .ZN(new_n496));
  OAI21_X1  g310(.A(new_n494), .B1(new_n493), .B2(new_n495), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  OAI211_X1 g312(.A(new_n492), .B(new_n498), .C1(new_n325), .C2(new_n349), .ZN(new_n499));
  NOR2_X1   g313(.A1(new_n487), .A2(G110), .ZN(new_n500));
  AND2_X1   g314(.A1(new_n493), .A2(new_n495), .ZN(new_n501));
  OAI211_X1 g315(.A(new_n338), .B(new_n306), .C1(new_n500), .C2(new_n501), .ZN(new_n502));
  XNOR2_X1  g316(.A(KEYINPUT22), .B(G137), .ZN(new_n503));
  XNOR2_X1  g317(.A(new_n503), .B(KEYINPUT73), .ZN(new_n504));
  AND3_X1   g318(.A1(new_n260), .A2(G221), .A3(G234), .ZN(new_n505));
  XNOR2_X1  g319(.A(new_n504), .B(new_n505), .ZN(new_n506));
  AND3_X1   g320(.A1(new_n499), .A2(new_n502), .A3(new_n506), .ZN(new_n507));
  AOI21_X1  g321(.A(new_n506), .B1(new_n499), .B2(new_n502), .ZN(new_n508));
  NOR3_X1   g322(.A1(new_n507), .A2(new_n508), .A3(G902), .ZN(new_n509));
  OAI21_X1  g323(.A(new_n481), .B1(new_n509), .B2(KEYINPUT74), .ZN(new_n510));
  AOI21_X1  g324(.A(new_n373), .B1(G234), .B2(new_n266), .ZN(new_n511));
  INV_X1    g325(.A(new_n508), .ZN(new_n512));
  NAND3_X1  g326(.A1(new_n499), .A2(new_n502), .A3(new_n506), .ZN(new_n513));
  NAND3_X1  g327(.A1(new_n512), .A2(new_n266), .A3(new_n513), .ZN(new_n514));
  INV_X1    g328(.A(KEYINPUT74), .ZN(new_n515));
  NAND3_X1  g329(.A1(new_n514), .A2(new_n515), .A3(KEYINPUT25), .ZN(new_n516));
  NAND3_X1  g330(.A1(new_n510), .A2(new_n511), .A3(new_n516), .ZN(new_n517));
  NOR2_X1   g331(.A1(new_n511), .A2(G902), .ZN(new_n518));
  XOR2_X1   g332(.A(new_n518), .B(KEYINPUT75), .Z(new_n519));
  NAND3_X1  g333(.A1(new_n512), .A2(new_n519), .A3(new_n513), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n517), .A2(new_n520), .ZN(new_n521));
  XNOR2_X1  g335(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n522));
  XNOR2_X1  g336(.A(new_n522), .B(G101), .ZN(new_n523));
  NAND3_X1  g337(.A1(new_n310), .A2(new_n260), .A3(G210), .ZN(new_n524));
  XNOR2_X1  g338(.A(new_n523), .B(new_n524), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n417), .A2(new_n437), .ZN(new_n526));
  NOR2_X1   g340(.A1(new_n209), .A2(new_n210), .ZN(new_n527));
  NOR2_X1   g341(.A1(new_n230), .A2(new_n527), .ZN(new_n528));
  INV_X1    g342(.A(new_n431), .ZN(new_n529));
  NOR2_X1   g343(.A1(new_n379), .A2(G137), .ZN(new_n530));
  OAI21_X1  g344(.A(G131), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  NAND3_X1  g345(.A1(new_n258), .A2(new_n436), .A3(new_n531), .ZN(new_n532));
  AND3_X1   g346(.A1(new_n526), .A2(new_n528), .A3(new_n532), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n252), .A2(KEYINPUT65), .ZN(new_n534));
  INV_X1    g348(.A(KEYINPUT65), .ZN(new_n535));
  OAI211_X1 g349(.A(new_n535), .B(new_n246), .C1(new_n250), .C2(new_n251), .ZN(new_n536));
  NAND3_X1  g350(.A1(new_n534), .A2(new_n437), .A3(new_n536), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n537), .A2(new_n532), .ZN(new_n538));
  AOI22_X1  g352(.A1(KEYINPUT28), .A2(new_n533), .B1(new_n538), .B2(new_n211), .ZN(new_n539));
  NAND3_X1  g353(.A1(new_n526), .A2(new_n528), .A3(new_n532), .ZN(new_n540));
  INV_X1    g354(.A(KEYINPUT28), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  AOI21_X1  g356(.A(new_n525), .B1(new_n539), .B2(new_n542), .ZN(new_n543));
  INV_X1    g357(.A(new_n543), .ZN(new_n544));
  AND3_X1   g358(.A1(new_n540), .A2(KEYINPUT68), .A3(new_n525), .ZN(new_n545));
  AOI21_X1  g359(.A(KEYINPUT68), .B1(new_n540), .B2(new_n525), .ZN(new_n546));
  NOR2_X1   g360(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  AOI21_X1  g361(.A(KEYINPUT30), .B1(new_n537), .B2(new_n532), .ZN(new_n548));
  AND3_X1   g362(.A1(new_n526), .A2(KEYINPUT30), .A3(new_n532), .ZN(new_n549));
  NOR3_X1   g363(.A1(new_n548), .A2(new_n549), .A3(new_n528), .ZN(new_n550));
  INV_X1    g364(.A(KEYINPUT31), .ZN(new_n551));
  NOR3_X1   g365(.A1(new_n547), .A2(new_n550), .A3(new_n551), .ZN(new_n552));
  NOR2_X1   g366(.A1(new_n548), .A2(new_n549), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n553), .A2(new_n211), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n540), .A2(new_n525), .ZN(new_n555));
  INV_X1    g369(.A(KEYINPUT68), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  NAND3_X1  g371(.A1(new_n540), .A2(new_n525), .A3(KEYINPUT68), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  AOI21_X1  g373(.A(KEYINPUT31), .B1(new_n554), .B2(new_n559), .ZN(new_n560));
  OAI21_X1  g374(.A(new_n544), .B1(new_n552), .B2(new_n560), .ZN(new_n561));
  INV_X1    g375(.A(KEYINPUT32), .ZN(new_n562));
  NOR2_X1   g376(.A1(G472), .A2(G902), .ZN(new_n563));
  NAND3_X1  g377(.A1(new_n561), .A2(new_n562), .A3(new_n563), .ZN(new_n564));
  OAI21_X1  g378(.A(new_n551), .B1(new_n547), .B2(new_n550), .ZN(new_n565));
  NAND3_X1  g379(.A1(new_n554), .A2(new_n559), .A3(KEYINPUT31), .ZN(new_n566));
  AOI21_X1  g380(.A(new_n543), .B1(new_n565), .B2(new_n566), .ZN(new_n567));
  INV_X1    g381(.A(new_n563), .ZN(new_n568));
  OAI21_X1  g382(.A(KEYINPUT32), .B1(new_n567), .B2(new_n568), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n564), .A2(new_n569), .ZN(new_n570));
  AOI21_X1  g384(.A(new_n525), .B1(new_n554), .B2(new_n540), .ZN(new_n571));
  AND3_X1   g385(.A1(new_n539), .A2(new_n525), .A3(new_n542), .ZN(new_n572));
  NOR3_X1   g386(.A1(new_n571), .A2(new_n572), .A3(KEYINPUT29), .ZN(new_n573));
  AOI21_X1  g387(.A(new_n528), .B1(new_n526), .B2(new_n532), .ZN(new_n574));
  OAI21_X1  g388(.A(KEYINPUT28), .B1(new_n533), .B2(new_n574), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n575), .A2(KEYINPUT69), .ZN(new_n576));
  INV_X1    g390(.A(KEYINPUT69), .ZN(new_n577));
  OAI211_X1 g391(.A(new_n577), .B(KEYINPUT28), .C1(new_n533), .C2(new_n574), .ZN(new_n578));
  NAND4_X1  g392(.A1(new_n576), .A2(KEYINPUT29), .A3(new_n542), .A4(new_n578), .ZN(new_n579));
  INV_X1    g393(.A(new_n525), .ZN(new_n580));
  OAI21_X1  g394(.A(new_n266), .B1(new_n579), .B2(new_n580), .ZN(new_n581));
  OAI21_X1  g395(.A(G472), .B1(new_n573), .B2(new_n581), .ZN(new_n582));
  AOI21_X1  g396(.A(new_n521), .B1(new_n570), .B2(new_n582), .ZN(new_n583));
  NAND3_X1  g397(.A1(new_n478), .A2(new_n480), .A3(new_n583), .ZN(new_n584));
  XNOR2_X1  g398(.A(new_n584), .B(KEYINPUT97), .ZN(new_n585));
  XNOR2_X1  g399(.A(new_n585), .B(new_n227), .ZN(G3));
  OR2_X1    g400(.A1(new_n472), .A2(new_n476), .ZN(new_n587));
  INV_X1    g401(.A(new_n521), .ZN(new_n588));
  OAI21_X1  g402(.A(G472), .B1(new_n567), .B2(G902), .ZN(new_n589));
  OAI21_X1  g403(.A(new_n589), .B1(new_n567), .B2(new_n568), .ZN(new_n590));
  INV_X1    g404(.A(new_n590), .ZN(new_n591));
  NAND3_X1  g405(.A1(new_n587), .A2(new_n588), .A3(new_n591), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n277), .A2(new_n279), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n593), .A2(new_n292), .ZN(new_n594));
  NOR2_X1   g408(.A1(new_n594), .A2(new_n291), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n366), .A2(new_n367), .ZN(new_n596));
  INV_X1    g410(.A(G475), .ZN(new_n597));
  OAI211_X1 g411(.A(new_n597), .B(new_n266), .C1(new_n364), .C2(new_n365), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n596), .A2(new_n598), .ZN(new_n599));
  AOI22_X1  g413(.A1(new_n599), .A2(new_n368), .B1(G475), .B2(new_n346), .ZN(new_n600));
  AOI21_X1  g414(.A(G478), .B1(new_n401), .B2(new_n266), .ZN(new_n601));
  AND3_X1   g415(.A1(new_n393), .A2(KEYINPUT33), .A3(new_n395), .ZN(new_n602));
  INV_X1    g416(.A(KEYINPUT33), .ZN(new_n603));
  AOI211_X1 g417(.A(G902), .B(new_n602), .C1(new_n401), .C2(new_n603), .ZN(new_n604));
  AOI21_X1  g418(.A(new_n601), .B1(new_n604), .B2(G478), .ZN(new_n605));
  NOR2_X1   g419(.A1(new_n600), .A2(new_n605), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n595), .A2(new_n606), .ZN(new_n607));
  NOR2_X1   g421(.A1(new_n592), .A2(new_n607), .ZN(new_n608));
  XNOR2_X1  g422(.A(KEYINPUT34), .B(G104), .ZN(new_n609));
  XNOR2_X1  g423(.A(new_n608), .B(new_n609), .ZN(G6));
  NAND2_X1  g424(.A1(new_n598), .A2(new_n367), .ZN(new_n611));
  NAND3_X1  g425(.A1(new_n362), .A2(KEYINPUT20), .A3(new_n266), .ZN(new_n612));
  NAND4_X1  g426(.A1(new_n407), .A2(new_n347), .A3(new_n611), .A4(new_n612), .ZN(new_n613));
  NOR4_X1   g427(.A1(new_n592), .A2(new_n291), .A3(new_n594), .A4(new_n613), .ZN(new_n614));
  XNOR2_X1  g428(.A(KEYINPUT35), .B(G107), .ZN(new_n615));
  XNOR2_X1  g429(.A(new_n614), .B(new_n615), .ZN(G9));
  INV_X1    g430(.A(new_n506), .ZN(new_n617));
  NOR2_X1   g431(.A1(new_n617), .A2(KEYINPUT36), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n499), .A2(new_n502), .ZN(new_n619));
  XNOR2_X1  g433(.A(new_n618), .B(new_n619), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n620), .A2(new_n519), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n517), .A2(new_n621), .ZN(new_n622));
  NAND4_X1  g436(.A1(new_n478), .A2(new_n480), .A3(new_n591), .A4(new_n622), .ZN(new_n623));
  XNOR2_X1  g437(.A(KEYINPUT98), .B(KEYINPUT37), .ZN(new_n624));
  XNOR2_X1  g438(.A(new_n624), .B(G110), .ZN(new_n625));
  XNOR2_X1  g439(.A(new_n623), .B(new_n625), .ZN(G12));
  AOI21_X1  g440(.A(new_n562), .B1(new_n561), .B2(new_n563), .ZN(new_n627));
  NOR3_X1   g441(.A1(new_n567), .A2(KEYINPUT32), .A3(new_n568), .ZN(new_n628));
  OAI21_X1  g442(.A(new_n582), .B1(new_n627), .B2(new_n628), .ZN(new_n629));
  INV_X1    g443(.A(G900), .ZN(new_n630));
  NAND2_X1  g444(.A1(new_n286), .A2(new_n630), .ZN(new_n631));
  AND2_X1   g445(.A1(new_n290), .A2(new_n631), .ZN(new_n632));
  NOR2_X1   g446(.A1(new_n613), .A2(new_n632), .ZN(new_n633));
  AOI21_X1  g447(.A(new_n293), .B1(new_n277), .B2(new_n279), .ZN(new_n634));
  AND4_X1   g448(.A1(new_n629), .A2(new_n633), .A3(new_n634), .A4(new_n622), .ZN(new_n635));
  NAND2_X1  g449(.A1(new_n587), .A2(new_n635), .ZN(new_n636));
  XNOR2_X1  g450(.A(new_n636), .B(G128), .ZN(G30));
  XNOR2_X1  g451(.A(new_n282), .B(KEYINPUT38), .ZN(new_n638));
  INV_X1    g452(.A(new_n638), .ZN(new_n639));
  INV_X1    g453(.A(new_n407), .ZN(new_n640));
  NOR3_X1   g454(.A1(new_n600), .A2(new_n293), .A3(new_n640), .ZN(new_n641));
  OAI21_X1  g455(.A(new_n580), .B1(new_n533), .B2(new_n574), .ZN(new_n642));
  XOR2_X1   g456(.A(new_n642), .B(KEYINPUT99), .Z(new_n643));
  NOR2_X1   g457(.A1(new_n547), .A2(new_n550), .ZN(new_n644));
  OAI21_X1  g458(.A(new_n266), .B1(new_n643), .B2(new_n644), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n645), .A2(G472), .ZN(new_n646));
  AOI21_X1  g460(.A(new_n622), .B1(new_n570), .B2(new_n646), .ZN(new_n647));
  NAND3_X1  g461(.A1(new_n639), .A2(new_n641), .A3(new_n647), .ZN(new_n648));
  XOR2_X1   g462(.A(new_n632), .B(KEYINPUT39), .Z(new_n649));
  AOI21_X1  g463(.A(KEYINPUT40), .B1(new_n587), .B2(new_n649), .ZN(new_n650));
  INV_X1    g464(.A(new_n650), .ZN(new_n651));
  NAND3_X1  g465(.A1(new_n587), .A2(KEYINPUT40), .A3(new_n649), .ZN(new_n652));
  AOI21_X1  g466(.A(new_n648), .B1(new_n651), .B2(new_n652), .ZN(new_n653));
  XNOR2_X1  g467(.A(new_n653), .B(new_n244), .ZN(G45));
  NOR3_X1   g468(.A1(new_n600), .A2(new_n605), .A3(new_n632), .ZN(new_n655));
  AND4_X1   g469(.A1(new_n629), .A2(new_n655), .A3(new_n634), .A4(new_n622), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n587), .A2(new_n656), .ZN(new_n657));
  XNOR2_X1  g471(.A(new_n657), .B(G146), .ZN(G48));
  NOR2_X1   g472(.A1(new_n412), .A2(KEYINPUT100), .ZN(new_n659));
  NAND2_X1  g473(.A1(new_n447), .A2(new_n458), .ZN(new_n660));
  AOI22_X1  g474(.A1(new_n660), .A2(new_n454), .B1(new_n469), .B2(new_n450), .ZN(new_n661));
  OAI21_X1  g475(.A(new_n659), .B1(new_n661), .B2(G902), .ZN(new_n662));
  INV_X1    g476(.A(new_n659), .ZN(new_n663));
  OAI211_X1 g477(.A(new_n266), .B(new_n663), .C1(new_n456), .C2(new_n459), .ZN(new_n664));
  AND3_X1   g478(.A1(new_n662), .A2(new_n664), .A3(new_n475), .ZN(new_n665));
  NAND4_X1  g479(.A1(new_n595), .A2(new_n583), .A3(new_n606), .A4(new_n665), .ZN(new_n666));
  XNOR2_X1  g480(.A(KEYINPUT41), .B(G113), .ZN(new_n667));
  XNOR2_X1  g481(.A(new_n666), .B(new_n667), .ZN(G15));
  INV_X1    g482(.A(new_n613), .ZN(new_n669));
  NAND4_X1  g483(.A1(new_n595), .A2(new_n583), .A3(new_n669), .A4(new_n665), .ZN(new_n670));
  XNOR2_X1  g484(.A(KEYINPUT101), .B(G116), .ZN(new_n671));
  XNOR2_X1  g485(.A(new_n670), .B(new_n671), .ZN(G18));
  AND3_X1   g486(.A1(new_n629), .A2(new_n634), .A3(new_n622), .ZN(new_n673));
  NAND3_X1  g487(.A1(new_n662), .A2(new_n664), .A3(new_n475), .ZN(new_n674));
  NOR2_X1   g488(.A1(new_n674), .A2(new_n291), .ZN(new_n675));
  NAND4_X1  g489(.A1(new_n673), .A2(new_n640), .A3(new_n600), .A4(new_n675), .ZN(new_n676));
  XNOR2_X1  g490(.A(new_n676), .B(G119), .ZN(G21));
  INV_X1    g491(.A(KEYINPUT102), .ZN(new_n678));
  NAND3_X1  g492(.A1(new_n641), .A2(new_n678), .A3(new_n593), .ZN(new_n679));
  NAND4_X1  g493(.A1(new_n371), .A2(new_n593), .A3(new_n292), .A4(new_n407), .ZN(new_n680));
  NAND2_X1  g494(.A1(new_n680), .A2(KEYINPUT102), .ZN(new_n681));
  NAND2_X1  g495(.A1(new_n679), .A2(new_n681), .ZN(new_n682));
  NAND3_X1  g496(.A1(new_n576), .A2(new_n542), .A3(new_n578), .ZN(new_n683));
  NAND2_X1  g497(.A1(new_n683), .A2(new_n580), .ZN(new_n684));
  OAI21_X1  g498(.A(new_n684), .B1(new_n560), .B2(new_n552), .ZN(new_n685));
  NAND2_X1  g499(.A1(new_n685), .A2(new_n563), .ZN(new_n686));
  NAND2_X1  g500(.A1(new_n686), .A2(new_n589), .ZN(new_n687));
  NOR4_X1   g501(.A1(new_n674), .A2(new_n687), .A3(new_n291), .A4(new_n521), .ZN(new_n688));
  NAND2_X1  g502(.A1(new_n682), .A2(new_n688), .ZN(new_n689));
  XOR2_X1   g503(.A(new_n689), .B(KEYINPUT103), .Z(new_n690));
  XNOR2_X1  g504(.A(new_n690), .B(G122), .ZN(G24));
  AND3_X1   g505(.A1(new_n622), .A2(new_n686), .A3(new_n589), .ZN(new_n692));
  NAND4_X1  g506(.A1(new_n655), .A2(new_n665), .A3(new_n692), .A4(new_n634), .ZN(new_n693));
  INV_X1    g507(.A(KEYINPUT104), .ZN(new_n694));
  NAND2_X1  g508(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  NOR2_X1   g509(.A1(new_n674), .A2(new_n594), .ZN(new_n696));
  NAND4_X1  g510(.A1(new_n696), .A2(KEYINPUT104), .A3(new_n655), .A4(new_n692), .ZN(new_n697));
  NAND2_X1  g511(.A1(new_n695), .A2(new_n697), .ZN(new_n698));
  XNOR2_X1  g512(.A(new_n698), .B(G125), .ZN(G27));
  INV_X1    g513(.A(KEYINPUT42), .ZN(new_n700));
  INV_X1    g514(.A(KEYINPUT105), .ZN(new_n701));
  NAND2_X1  g515(.A1(new_n471), .A2(new_n701), .ZN(new_n702));
  NAND4_X1  g516(.A1(new_n468), .A2(KEYINPUT105), .A3(G469), .A4(new_n470), .ZN(new_n703));
  NAND3_X1  g517(.A1(new_n702), .A2(new_n463), .A3(new_n703), .ZN(new_n704));
  NAND3_X1  g518(.A1(new_n704), .A2(new_n475), .A3(new_n583), .ZN(new_n705));
  AOI21_X1  g519(.A(new_n293), .B1(new_n280), .B2(new_n281), .ZN(new_n706));
  NAND2_X1  g520(.A1(new_n706), .A2(new_n655), .ZN(new_n707));
  OAI21_X1  g521(.A(new_n700), .B1(new_n705), .B2(new_n707), .ZN(new_n708));
  INV_X1    g522(.A(KEYINPUT106), .ZN(new_n709));
  NAND2_X1  g523(.A1(new_n460), .A2(new_n462), .ZN(new_n710));
  AOI21_X1  g524(.A(new_n710), .B1(new_n701), .B2(new_n471), .ZN(new_n711));
  AOI21_X1  g525(.A(new_n411), .B1(new_n711), .B2(new_n703), .ZN(new_n712));
  AND2_X1   g526(.A1(new_n706), .A2(new_n655), .ZN(new_n713));
  NAND4_X1  g527(.A1(new_n712), .A2(new_n713), .A3(KEYINPUT42), .A4(new_n583), .ZN(new_n714));
  AND3_X1   g528(.A1(new_n708), .A2(new_n709), .A3(new_n714), .ZN(new_n715));
  AOI21_X1  g529(.A(new_n709), .B1(new_n708), .B2(new_n714), .ZN(new_n716));
  NOR2_X1   g530(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  XNOR2_X1  g531(.A(new_n717), .B(new_n327), .ZN(G33));
  INV_X1    g532(.A(new_n706), .ZN(new_n719));
  NOR4_X1   g533(.A1(new_n705), .A2(new_n613), .A3(new_n632), .A4(new_n719), .ZN(new_n720));
  XNOR2_X1  g534(.A(new_n720), .B(new_n379), .ZN(G36));
  INV_X1    g535(.A(KEYINPUT107), .ZN(new_n722));
  AND3_X1   g536(.A1(new_n447), .A2(new_n450), .A3(new_n466), .ZN(new_n723));
  AOI21_X1  g537(.A(new_n466), .B1(new_n447), .B2(new_n450), .ZN(new_n724));
  NOR2_X1   g538(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  AOI22_X1  g539(.A1(new_n725), .A2(new_n454), .B1(new_n469), .B2(new_n458), .ZN(new_n726));
  OAI211_X1 g540(.A(new_n722), .B(G469), .C1(new_n726), .C2(KEYINPUT45), .ZN(new_n727));
  NAND2_X1  g541(.A1(KEYINPUT45), .A2(G469), .ZN(new_n728));
  NAND3_X1  g542(.A1(new_n471), .A2(KEYINPUT107), .A3(new_n728), .ZN(new_n729));
  NAND2_X1  g543(.A1(new_n726), .A2(KEYINPUT45), .ZN(new_n730));
  NAND3_X1  g544(.A1(new_n727), .A2(new_n729), .A3(new_n730), .ZN(new_n731));
  NAND2_X1  g545(.A1(new_n731), .A2(new_n462), .ZN(new_n732));
  INV_X1    g546(.A(KEYINPUT46), .ZN(new_n733));
  NAND2_X1  g547(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  NAND3_X1  g548(.A1(new_n731), .A2(KEYINPUT46), .A3(new_n462), .ZN(new_n735));
  NAND3_X1  g549(.A1(new_n734), .A2(new_n460), .A3(new_n735), .ZN(new_n736));
  AND2_X1   g550(.A1(new_n736), .A2(new_n475), .ZN(new_n737));
  AND2_X1   g551(.A1(new_n737), .A2(new_n649), .ZN(new_n738));
  INV_X1    g552(.A(KEYINPUT43), .ZN(new_n739));
  OAI21_X1  g553(.A(new_n739), .B1(new_n371), .B2(KEYINPUT108), .ZN(new_n740));
  NOR2_X1   g554(.A1(new_n371), .A2(new_n605), .ZN(new_n741));
  XNOR2_X1  g555(.A(new_n740), .B(new_n741), .ZN(new_n742));
  NAND3_X1  g556(.A1(new_n742), .A2(new_n590), .A3(new_n622), .ZN(new_n743));
  INV_X1    g557(.A(KEYINPUT44), .ZN(new_n744));
  NAND2_X1  g558(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  INV_X1    g559(.A(KEYINPUT109), .ZN(new_n746));
  XNOR2_X1  g560(.A(new_n745), .B(new_n746), .ZN(new_n747));
  OR2_X1    g561(.A1(new_n743), .A2(new_n744), .ZN(new_n748));
  NAND4_X1  g562(.A1(new_n738), .A2(new_n706), .A3(new_n747), .A4(new_n748), .ZN(new_n749));
  XNOR2_X1  g563(.A(new_n749), .B(G137), .ZN(G39));
  OR2_X1    g564(.A1(new_n573), .A2(new_n581), .ZN(new_n751));
  AOI22_X1  g565(.A1(new_n751), .A2(G472), .B1(new_n564), .B2(new_n569), .ZN(new_n752));
  NOR2_X1   g566(.A1(new_n707), .A2(new_n588), .ZN(new_n753));
  AND3_X1   g567(.A1(new_n736), .A2(KEYINPUT47), .A3(new_n475), .ZN(new_n754));
  AOI21_X1  g568(.A(KEYINPUT47), .B1(new_n736), .B2(new_n475), .ZN(new_n755));
  OAI211_X1 g569(.A(new_n752), .B(new_n753), .C1(new_n754), .C2(new_n755), .ZN(new_n756));
  XNOR2_X1  g570(.A(new_n756), .B(G140), .ZN(G42));
  OR2_X1    g571(.A1(G952), .A2(G953), .ZN(new_n758));
  INV_X1    g572(.A(new_n290), .ZN(new_n759));
  NOR2_X1   g573(.A1(new_n687), .A2(new_n521), .ZN(new_n760));
  AND3_X1   g574(.A1(new_n742), .A2(new_n759), .A3(new_n760), .ZN(new_n761));
  NAND2_X1  g575(.A1(new_n665), .A2(new_n293), .ZN(new_n762));
  OR2_X1    g576(.A1(new_n762), .A2(KEYINPUT114), .ZN(new_n763));
  NAND2_X1  g577(.A1(new_n762), .A2(KEYINPUT114), .ZN(new_n764));
  NAND2_X1  g578(.A1(new_n638), .A2(new_n764), .ZN(new_n765));
  INV_X1    g579(.A(new_n765), .ZN(new_n766));
  NAND4_X1  g580(.A1(new_n761), .A2(KEYINPUT50), .A3(new_n763), .A4(new_n766), .ZN(new_n767));
  INV_X1    g581(.A(KEYINPUT50), .ZN(new_n768));
  NAND4_X1  g582(.A1(new_n742), .A2(new_n763), .A3(new_n759), .A4(new_n760), .ZN(new_n769));
  OAI21_X1  g583(.A(new_n768), .B1(new_n769), .B2(new_n765), .ZN(new_n770));
  NAND2_X1  g584(.A1(new_n767), .A2(new_n770), .ZN(new_n771));
  NOR3_X1   g585(.A1(new_n719), .A2(new_n290), .A3(new_n674), .ZN(new_n772));
  NAND3_X1  g586(.A1(new_n742), .A2(new_n772), .A3(new_n692), .ZN(new_n773));
  AND3_X1   g587(.A1(new_n570), .A2(new_n588), .A3(new_n646), .ZN(new_n774));
  NAND4_X1  g588(.A1(new_n772), .A2(new_n600), .A3(new_n605), .A4(new_n774), .ZN(new_n775));
  AND2_X1   g589(.A1(new_n773), .A2(new_n775), .ZN(new_n776));
  AND2_X1   g590(.A1(new_n771), .A2(new_n776), .ZN(new_n777));
  NAND2_X1  g591(.A1(new_n662), .A2(new_n664), .ZN(new_n778));
  XOR2_X1   g592(.A(new_n778), .B(KEYINPUT110), .Z(new_n779));
  NOR2_X1   g593(.A1(new_n779), .A2(new_n475), .ZN(new_n780));
  NOR3_X1   g594(.A1(new_n754), .A2(new_n755), .A3(new_n780), .ZN(new_n781));
  NAND2_X1  g595(.A1(new_n761), .A2(new_n706), .ZN(new_n782));
  OAI211_X1 g596(.A(new_n777), .B(KEYINPUT51), .C1(new_n781), .C2(new_n782), .ZN(new_n783));
  NAND2_X1  g597(.A1(new_n761), .A2(new_n696), .ZN(new_n784));
  NAND3_X1  g598(.A1(new_n772), .A2(new_n606), .A3(new_n774), .ZN(new_n785));
  NAND4_X1  g599(.A1(new_n783), .A2(new_n289), .A3(new_n784), .A4(new_n785), .ZN(new_n786));
  NAND3_X1  g600(.A1(new_n742), .A2(new_n772), .A3(new_n583), .ZN(new_n787));
  XOR2_X1   g601(.A(new_n787), .B(KEYINPUT48), .Z(new_n788));
  NOR2_X1   g602(.A1(new_n786), .A2(new_n788), .ZN(new_n789));
  OAI22_X1  g603(.A1(new_n656), .A2(new_n635), .B1(new_n472), .B2(new_n476), .ZN(new_n790));
  INV_X1    g604(.A(new_n632), .ZN(new_n791));
  AND2_X1   g605(.A1(new_n647), .A2(new_n791), .ZN(new_n792));
  NAND3_X1  g606(.A1(new_n682), .A2(new_n712), .A3(new_n792), .ZN(new_n793));
  NAND3_X1  g607(.A1(new_n790), .A2(new_n698), .A3(new_n793), .ZN(new_n794));
  NAND2_X1  g608(.A1(new_n794), .A2(KEYINPUT52), .ZN(new_n795));
  INV_X1    g609(.A(KEYINPUT52), .ZN(new_n796));
  NAND4_X1  g610(.A1(new_n790), .A2(new_n698), .A3(new_n793), .A4(new_n796), .ZN(new_n797));
  AND3_X1   g611(.A1(new_n347), .A2(new_n611), .A3(new_n612), .ZN(new_n798));
  NOR2_X1   g612(.A1(new_n752), .A2(new_n407), .ZN(new_n799));
  OAI211_X1 g613(.A(new_n798), .B(new_n799), .C1(new_n472), .C2(new_n476), .ZN(new_n800));
  INV_X1    g614(.A(new_n687), .ZN(new_n801));
  NAND3_X1  g615(.A1(new_n712), .A2(new_n606), .A3(new_n801), .ZN(new_n802));
  NAND2_X1  g616(.A1(new_n800), .A2(new_n802), .ZN(new_n803));
  NAND4_X1  g617(.A1(new_n803), .A2(new_n622), .A3(new_n791), .A4(new_n706), .ZN(new_n804));
  NAND3_X1  g618(.A1(new_n795), .A2(new_n797), .A3(new_n804), .ZN(new_n805));
  INV_X1    g619(.A(new_n720), .ZN(new_n806));
  OAI21_X1  g620(.A(new_n806), .B1(new_n715), .B2(new_n716), .ZN(new_n807));
  NOR2_X1   g621(.A1(new_n805), .A2(new_n807), .ZN(new_n808));
  AND4_X1   g622(.A1(new_n666), .A2(new_n689), .A3(new_n670), .A4(new_n676), .ZN(new_n809));
  OAI21_X1  g623(.A(KEYINPUT111), .B1(new_n371), .B2(new_n640), .ZN(new_n810));
  INV_X1    g624(.A(KEYINPUT111), .ZN(new_n811));
  NAND3_X1  g625(.A1(new_n600), .A2(new_n811), .A3(new_n407), .ZN(new_n812));
  OAI211_X1 g626(.A(new_n810), .B(new_n812), .C1(new_n600), .C2(new_n605), .ZN(new_n813));
  NOR2_X1   g627(.A1(new_n282), .A2(new_n294), .ZN(new_n814));
  AND2_X1   g628(.A1(new_n813), .A2(new_n814), .ZN(new_n815));
  NAND4_X1  g629(.A1(new_n815), .A2(new_n587), .A3(new_n588), .A4(new_n591), .ZN(new_n816));
  NAND4_X1  g630(.A1(new_n623), .A2(new_n809), .A3(new_n584), .A4(new_n816), .ZN(new_n817));
  INV_X1    g631(.A(new_n817), .ZN(new_n818));
  AOI21_X1  g632(.A(KEYINPUT53), .B1(new_n808), .B2(new_n818), .ZN(new_n819));
  AND2_X1   g633(.A1(new_n708), .A2(new_n714), .ZN(new_n820));
  NAND2_X1  g634(.A1(new_n806), .A2(KEYINPUT53), .ZN(new_n821));
  NOR4_X1   g635(.A1(new_n805), .A2(new_n817), .A3(new_n820), .A4(new_n821), .ZN(new_n822));
  NOR2_X1   g636(.A1(new_n819), .A2(new_n822), .ZN(new_n823));
  XNOR2_X1  g637(.A(KEYINPUT113), .B(KEYINPUT54), .ZN(new_n824));
  INV_X1    g638(.A(new_n824), .ZN(new_n825));
  NAND2_X1  g639(.A1(new_n823), .A2(new_n825), .ZN(new_n826));
  INV_X1    g640(.A(KEYINPUT53), .ZN(new_n827));
  NOR4_X1   g641(.A1(new_n805), .A2(new_n817), .A3(new_n807), .A4(new_n827), .ZN(new_n828));
  OAI21_X1  g642(.A(KEYINPUT54), .B1(new_n819), .B2(new_n828), .ZN(new_n829));
  INV_X1    g643(.A(KEYINPUT112), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  OAI211_X1 g645(.A(KEYINPUT112), .B(KEYINPUT54), .C1(new_n819), .C2(new_n828), .ZN(new_n832));
  NAND4_X1  g646(.A1(new_n789), .A2(new_n826), .A3(new_n831), .A4(new_n832), .ZN(new_n833));
  INV_X1    g647(.A(KEYINPUT51), .ZN(new_n834));
  OR2_X1    g648(.A1(new_n771), .A2(KEYINPUT115), .ZN(new_n835));
  NAND2_X1  g649(.A1(new_n771), .A2(KEYINPUT115), .ZN(new_n836));
  NAND3_X1  g650(.A1(new_n835), .A2(new_n776), .A3(new_n836), .ZN(new_n837));
  NOR2_X1   g651(.A1(new_n781), .A2(new_n782), .ZN(new_n838));
  OAI21_X1  g652(.A(new_n834), .B1(new_n837), .B2(new_n838), .ZN(new_n839));
  XNOR2_X1  g653(.A(new_n839), .B(KEYINPUT116), .ZN(new_n840));
  OAI21_X1  g654(.A(new_n758), .B1(new_n833), .B2(new_n840), .ZN(new_n841));
  OR2_X1    g655(.A1(new_n779), .A2(KEYINPUT49), .ZN(new_n842));
  NAND2_X1  g656(.A1(new_n779), .A2(KEYINPUT49), .ZN(new_n843));
  AND4_X1   g657(.A1(new_n741), .A2(new_n842), .A3(new_n843), .A4(new_n774), .ZN(new_n844));
  NAND4_X1  g658(.A1(new_n844), .A2(new_n475), .A3(new_n292), .A4(new_n638), .ZN(new_n845));
  NAND2_X1  g659(.A1(new_n841), .A2(new_n845), .ZN(G75));
  INV_X1    g660(.A(new_n823), .ZN(new_n847));
  NAND3_X1  g661(.A1(new_n847), .A2(G210), .A3(G902), .ZN(new_n848));
  INV_X1    g662(.A(KEYINPUT56), .ZN(new_n849));
  AND2_X1   g663(.A1(new_n241), .A2(new_n264), .ZN(new_n850));
  XNOR2_X1  g664(.A(new_n850), .B(new_n262), .ZN(new_n851));
  NOR2_X1   g665(.A1(new_n851), .A2(KEYINPUT55), .ZN(new_n852));
  AND2_X1   g666(.A1(new_n851), .A2(KEYINPUT55), .ZN(new_n853));
  AOI211_X1 g667(.A(new_n852), .B(new_n853), .C1(KEYINPUT117), .C2(new_n849), .ZN(new_n854));
  AND3_X1   g668(.A1(new_n848), .A2(new_n849), .A3(new_n854), .ZN(new_n855));
  AOI21_X1  g669(.A(new_n854), .B1(new_n848), .B2(new_n849), .ZN(new_n856));
  NOR2_X1   g670(.A1(new_n260), .A2(G952), .ZN(new_n857));
  NOR3_X1   g671(.A1(new_n855), .A2(new_n856), .A3(new_n857), .ZN(G51));
  NAND2_X1  g672(.A1(new_n462), .A2(KEYINPUT57), .ZN(new_n859));
  OAI21_X1  g673(.A(new_n824), .B1(new_n819), .B2(new_n822), .ZN(new_n860));
  INV_X1    g674(.A(new_n860), .ZN(new_n861));
  NOR3_X1   g675(.A1(new_n819), .A2(new_n822), .A3(new_n824), .ZN(new_n862));
  OAI21_X1  g676(.A(new_n859), .B1(new_n861), .B2(new_n862), .ZN(new_n863));
  NOR2_X1   g677(.A1(new_n462), .A2(KEYINPUT57), .ZN(new_n864));
  OAI22_X1  g678(.A1(new_n863), .A2(new_n864), .B1(new_n459), .B2(new_n456), .ZN(new_n865));
  NOR2_X1   g679(.A1(new_n823), .A2(new_n266), .ZN(new_n866));
  XOR2_X1   g680(.A(new_n731), .B(KEYINPUT118), .Z(new_n867));
  NAND2_X1  g681(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  AOI21_X1  g682(.A(new_n857), .B1(new_n865), .B2(new_n868), .ZN(G54));
  INV_X1    g683(.A(KEYINPUT119), .ZN(new_n870));
  INV_X1    g684(.A(KEYINPUT58), .ZN(new_n871));
  OAI21_X1  g685(.A(new_n870), .B1(new_n871), .B2(new_n597), .ZN(new_n872));
  NAND3_X1  g686(.A1(KEYINPUT119), .A2(KEYINPUT58), .A3(G475), .ZN(new_n873));
  NAND3_X1  g687(.A1(new_n866), .A2(new_n872), .A3(new_n873), .ZN(new_n874));
  NAND3_X1  g688(.A1(new_n874), .A2(new_n343), .A3(new_n361), .ZN(new_n875));
  INV_X1    g689(.A(new_n857), .ZN(new_n876));
  NAND2_X1  g690(.A1(new_n361), .A2(new_n343), .ZN(new_n877));
  NAND4_X1  g691(.A1(new_n866), .A2(new_n877), .A3(new_n872), .A4(new_n873), .ZN(new_n878));
  AND3_X1   g692(.A1(new_n875), .A2(new_n876), .A3(new_n878), .ZN(G60));
  AND2_X1   g693(.A1(new_n401), .A2(new_n603), .ZN(new_n880));
  OR2_X1    g694(.A1(new_n880), .A2(new_n602), .ZN(new_n881));
  XNOR2_X1  g695(.A(new_n881), .B(KEYINPUT120), .ZN(new_n882));
  INV_X1    g696(.A(new_n882), .ZN(new_n883));
  NAND3_X1  g697(.A1(new_n831), .A2(new_n826), .A3(new_n832), .ZN(new_n884));
  NAND2_X1  g698(.A1(G478), .A2(G902), .ZN(new_n885));
  XOR2_X1   g699(.A(new_n885), .B(KEYINPUT59), .Z(new_n886));
  INV_X1    g700(.A(new_n886), .ZN(new_n887));
  AOI21_X1  g701(.A(new_n883), .B1(new_n884), .B2(new_n887), .ZN(new_n888));
  AOI211_X1 g702(.A(new_n882), .B(new_n886), .C1(new_n826), .C2(new_n860), .ZN(new_n889));
  NOR3_X1   g703(.A1(new_n888), .A2(new_n857), .A3(new_n889), .ZN(G63));
  NAND2_X1  g704(.A1(G217), .A2(G902), .ZN(new_n891));
  XOR2_X1   g705(.A(new_n891), .B(KEYINPUT121), .Z(new_n892));
  XOR2_X1   g706(.A(new_n892), .B(KEYINPUT60), .Z(new_n893));
  INV_X1    g707(.A(new_n893), .ZN(new_n894));
  OAI22_X1  g708(.A1(new_n823), .A2(new_n894), .B1(new_n507), .B2(new_n508), .ZN(new_n895));
  AND2_X1   g709(.A1(new_n895), .A2(new_n876), .ZN(new_n896));
  NAND2_X1  g710(.A1(KEYINPUT122), .A2(KEYINPUT61), .ZN(new_n897));
  XOR2_X1   g711(.A(new_n897), .B(KEYINPUT123), .Z(new_n898));
  NAND3_X1  g712(.A1(new_n847), .A2(new_n620), .A3(new_n893), .ZN(new_n899));
  OR2_X1    g713(.A1(KEYINPUT122), .A2(KEYINPUT61), .ZN(new_n900));
  NAND4_X1  g714(.A1(new_n896), .A2(new_n898), .A3(new_n899), .A4(new_n900), .ZN(new_n901));
  NAND4_X1  g715(.A1(new_n899), .A2(new_n895), .A3(new_n876), .A4(new_n900), .ZN(new_n902));
  INV_X1    g716(.A(new_n898), .ZN(new_n903));
  NAND2_X1  g717(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  NAND2_X1  g718(.A1(new_n901), .A2(new_n904), .ZN(G66));
  AOI21_X1  g719(.A(new_n260), .B1(new_n283), .B2(G224), .ZN(new_n906));
  AOI21_X1  g720(.A(new_n906), .B1(new_n817), .B2(new_n260), .ZN(new_n907));
  INV_X1    g721(.A(G898), .ZN(new_n908));
  AOI21_X1  g722(.A(new_n850), .B1(new_n908), .B2(G953), .ZN(new_n909));
  XNOR2_X1  g723(.A(new_n907), .B(new_n909), .ZN(G69));
  NAND2_X1  g724(.A1(new_n350), .A2(new_n352), .ZN(new_n911));
  XNOR2_X1  g725(.A(new_n553), .B(new_n911), .ZN(new_n912));
  AND2_X1   g726(.A1(new_n813), .A2(new_n583), .ZN(new_n913));
  AND4_X1   g727(.A1(new_n587), .A2(new_n913), .A3(new_n649), .A4(new_n706), .ZN(new_n914));
  INV_X1    g728(.A(KEYINPUT62), .ZN(new_n915));
  NAND2_X1  g729(.A1(new_n790), .A2(new_n698), .ZN(new_n916));
  OAI21_X1  g730(.A(new_n915), .B1(new_n653), .B2(new_n916), .ZN(new_n917));
  INV_X1    g731(.A(new_n916), .ZN(new_n918));
  INV_X1    g732(.A(new_n652), .ZN(new_n919));
  NOR2_X1   g733(.A1(new_n919), .A2(new_n650), .ZN(new_n920));
  OAI211_X1 g734(.A(KEYINPUT62), .B(new_n918), .C1(new_n920), .C2(new_n648), .ZN(new_n921));
  AOI21_X1  g735(.A(new_n914), .B1(new_n917), .B2(new_n921), .ZN(new_n922));
  AND3_X1   g736(.A1(new_n922), .A2(new_n749), .A3(new_n756), .ZN(new_n923));
  OAI21_X1  g737(.A(new_n912), .B1(new_n923), .B2(G953), .ZN(new_n924));
  AOI21_X1  g738(.A(new_n912), .B1(G900), .B2(G953), .ZN(new_n925));
  OR2_X1    g739(.A1(new_n807), .A2(new_n916), .ZN(new_n926));
  INV_X1    g740(.A(new_n926), .ZN(new_n927));
  NAND3_X1  g741(.A1(new_n738), .A2(new_n583), .A3(new_n682), .ZN(new_n928));
  NAND4_X1  g742(.A1(new_n749), .A2(new_n927), .A3(new_n928), .A4(new_n756), .ZN(new_n929));
  OAI21_X1  g743(.A(new_n925), .B1(new_n929), .B2(G953), .ZN(new_n930));
  NAND2_X1  g744(.A1(new_n924), .A2(new_n930), .ZN(new_n931));
  AOI21_X1  g745(.A(new_n260), .B1(G227), .B2(G900), .ZN(new_n932));
  XNOR2_X1  g746(.A(new_n932), .B(KEYINPUT124), .ZN(new_n933));
  XNOR2_X1  g747(.A(new_n931), .B(new_n933), .ZN(G72));
  NAND4_X1  g748(.A1(new_n922), .A2(new_n749), .A3(new_n756), .A4(new_n818), .ZN(new_n935));
  XOR2_X1   g749(.A(KEYINPUT125), .B(KEYINPUT63), .Z(new_n936));
  NAND2_X1  g750(.A1(G472), .A2(G902), .ZN(new_n937));
  XNOR2_X1  g751(.A(new_n936), .B(new_n937), .ZN(new_n938));
  NAND2_X1  g752(.A1(new_n935), .A2(new_n938), .ZN(new_n939));
  INV_X1    g753(.A(KEYINPUT126), .ZN(new_n940));
  NAND2_X1  g754(.A1(new_n939), .A2(new_n940), .ZN(new_n941));
  NAND2_X1  g755(.A1(new_n554), .A2(new_n540), .ZN(new_n942));
  NAND3_X1  g756(.A1(new_n935), .A2(KEYINPUT126), .A3(new_n938), .ZN(new_n943));
  NAND4_X1  g757(.A1(new_n941), .A2(new_n525), .A3(new_n942), .A4(new_n943), .ZN(new_n944));
  OAI21_X1  g758(.A(new_n938), .B1(new_n929), .B2(new_n817), .ZN(new_n945));
  NAND2_X1  g759(.A1(new_n945), .A2(KEYINPUT127), .ZN(new_n946));
  NOR2_X1   g760(.A1(new_n942), .A2(new_n525), .ZN(new_n947));
  INV_X1    g761(.A(KEYINPUT127), .ZN(new_n948));
  OAI211_X1 g762(.A(new_n948), .B(new_n938), .C1(new_n929), .C2(new_n817), .ZN(new_n949));
  NAND3_X1  g763(.A1(new_n946), .A2(new_n947), .A3(new_n949), .ZN(new_n950));
  NOR2_X1   g764(.A1(new_n819), .A2(new_n828), .ZN(new_n951));
  NOR2_X1   g765(.A1(new_n571), .A2(new_n644), .ZN(new_n952));
  NOR2_X1   g766(.A1(new_n951), .A2(new_n952), .ZN(new_n953));
  AOI21_X1  g767(.A(new_n857), .B1(new_n953), .B2(new_n938), .ZN(new_n954));
  AND3_X1   g768(.A1(new_n944), .A2(new_n950), .A3(new_n954), .ZN(G57));
endmodule


