

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304,
         n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315,
         n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326,
         n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, n337,
         n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, n348,
         n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359,
         n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370,
         n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381,
         n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392,
         n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403,
         n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414,
         n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425,
         n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436,
         n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447,
         n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458,
         n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469,
         n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480,
         n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491,
         n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502,
         n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513,
         n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592;

  NOR2_X1 U326 ( .A1(n524), .A2(n454), .ZN(n568) );
  XNOR2_X1 U327 ( .A(n383), .B(n382), .ZN(n384) );
  XOR2_X1 U328 ( .A(KEYINPUT116), .B(n407), .Z(n294) );
  XOR2_X1 U329 ( .A(n400), .B(KEYINPUT14), .Z(n295) );
  NOR2_X1 U330 ( .A1(n588), .A2(n559), .ZN(n405) );
  NOR2_X1 U331 ( .A1(n533), .A2(n431), .ZN(n432) );
  XNOR2_X1 U332 ( .A(KEYINPUT64), .B(KEYINPUT48), .ZN(n418) );
  XNOR2_X1 U333 ( .A(n419), .B(n418), .ZN(n533) );
  XNOR2_X1 U334 ( .A(n385), .B(n384), .ZN(n386) );
  AND2_X1 U335 ( .A1(n470), .A2(n574), .ZN(n453) );
  XOR2_X1 U336 ( .A(n404), .B(n403), .Z(n584) );
  XOR2_X1 U337 ( .A(n389), .B(n388), .Z(n567) );
  XNOR2_X1 U338 ( .A(n456), .B(n455), .ZN(n457) );
  XNOR2_X1 U339 ( .A(n458), .B(n457), .ZN(G1349GAT) );
  XOR2_X1 U340 ( .A(KEYINPUT20), .B(G71GAT), .Z(n297) );
  XNOR2_X1 U341 ( .A(G99GAT), .B(G190GAT), .ZN(n296) );
  XNOR2_X1 U342 ( .A(n297), .B(n296), .ZN(n298) );
  XOR2_X1 U343 ( .A(n298), .B(G120GAT), .Z(n300) );
  XOR2_X1 U344 ( .A(G15GAT), .B(G127GAT), .Z(n401) );
  XNOR2_X1 U345 ( .A(G43GAT), .B(n401), .ZN(n299) );
  XNOR2_X1 U346 ( .A(n300), .B(n299), .ZN(n313) );
  XOR2_X1 U347 ( .A(KEYINPUT83), .B(G183GAT), .Z(n302) );
  NAND2_X1 U348 ( .A1(G227GAT), .A2(G233GAT), .ZN(n301) );
  XNOR2_X1 U349 ( .A(n302), .B(n301), .ZN(n303) );
  XOR2_X1 U350 ( .A(n303), .B(KEYINPUT84), .Z(n311) );
  XOR2_X1 U351 ( .A(KEYINPUT82), .B(G134GAT), .Z(n305) );
  XNOR2_X1 U352 ( .A(KEYINPUT81), .B(KEYINPUT0), .ZN(n304) );
  XNOR2_X1 U353 ( .A(n305), .B(n304), .ZN(n306) );
  XOR2_X1 U354 ( .A(G113GAT), .B(n306), .Z(n448) );
  XOR2_X1 U355 ( .A(KEYINPUT17), .B(KEYINPUT19), .Z(n308) );
  XNOR2_X1 U356 ( .A(KEYINPUT18), .B(G176GAT), .ZN(n307) );
  XNOR2_X1 U357 ( .A(n308), .B(n307), .ZN(n309) );
  XNOR2_X1 U358 ( .A(G169GAT), .B(n309), .ZN(n429) );
  XOR2_X1 U359 ( .A(n448), .B(n429), .Z(n310) );
  XNOR2_X1 U360 ( .A(n311), .B(n310), .ZN(n312) );
  XNOR2_X1 U361 ( .A(n313), .B(n312), .ZN(n536) );
  INV_X1 U362 ( .A(n536), .ZN(n524) );
  XOR2_X1 U363 ( .A(KEYINPUT89), .B(KEYINPUT23), .Z(n315) );
  XNOR2_X1 U364 ( .A(G22GAT), .B(KEYINPUT24), .ZN(n314) );
  XNOR2_X1 U365 ( .A(n315), .B(n314), .ZN(n321) );
  XOR2_X1 U366 ( .A(KEYINPUT87), .B(KEYINPUT21), .Z(n317) );
  XNOR2_X1 U367 ( .A(G197GAT), .B(G218GAT), .ZN(n316) );
  XNOR2_X1 U368 ( .A(n317), .B(n316), .ZN(n426) );
  XOR2_X1 U369 ( .A(G50GAT), .B(G162GAT), .Z(n383) );
  XOR2_X1 U370 ( .A(n426), .B(n383), .Z(n319) );
  NAND2_X1 U371 ( .A1(G228GAT), .A2(G233GAT), .ZN(n318) );
  XNOR2_X1 U372 ( .A(n319), .B(n318), .ZN(n320) );
  XNOR2_X1 U373 ( .A(n321), .B(n320), .ZN(n333) );
  XOR2_X1 U374 ( .A(G148GAT), .B(G155GAT), .Z(n323) );
  XNOR2_X1 U375 ( .A(G211GAT), .B(G204GAT), .ZN(n322) );
  XNOR2_X1 U376 ( .A(n323), .B(n322), .ZN(n324) );
  XOR2_X1 U377 ( .A(n324), .B(KEYINPUT90), .Z(n326) );
  XOR2_X1 U378 ( .A(G106GAT), .B(KEYINPUT72), .Z(n368) );
  XNOR2_X1 U379 ( .A(n368), .B(KEYINPUT22), .ZN(n325) );
  XNOR2_X1 U380 ( .A(n326), .B(n325), .ZN(n327) );
  XOR2_X1 U381 ( .A(n327), .B(G78GAT), .Z(n331) );
  XOR2_X1 U382 ( .A(KEYINPUT2), .B(KEYINPUT88), .Z(n329) );
  XNOR2_X1 U383 ( .A(G141GAT), .B(KEYINPUT3), .ZN(n328) );
  XNOR2_X1 U384 ( .A(n329), .B(n328), .ZN(n438) );
  XNOR2_X1 U385 ( .A(n438), .B(KEYINPUT86), .ZN(n330) );
  XNOR2_X1 U386 ( .A(n331), .B(n330), .ZN(n332) );
  XNOR2_X1 U387 ( .A(n333), .B(n332), .ZN(n470) );
  XOR2_X1 U388 ( .A(KEYINPUT30), .B(KEYINPUT66), .Z(n335) );
  XNOR2_X1 U389 ( .A(G1GAT), .B(KEYINPUT67), .ZN(n334) );
  XNOR2_X1 U390 ( .A(n335), .B(n334), .ZN(n352) );
  XOR2_X1 U391 ( .A(G197GAT), .B(G141GAT), .Z(n337) );
  XNOR2_X1 U392 ( .A(G36GAT), .B(G50GAT), .ZN(n336) );
  XNOR2_X1 U393 ( .A(n337), .B(n336), .ZN(n341) );
  XOR2_X1 U394 ( .A(G8GAT), .B(G113GAT), .Z(n339) );
  XNOR2_X1 U395 ( .A(G169GAT), .B(G15GAT), .ZN(n338) );
  XNOR2_X1 U396 ( .A(n339), .B(n338), .ZN(n340) );
  XOR2_X1 U397 ( .A(n341), .B(n340), .Z(n350) );
  XOR2_X1 U398 ( .A(KEYINPUT8), .B(KEYINPUT68), .Z(n343) );
  XNOR2_X1 U399 ( .A(G43GAT), .B(G29GAT), .ZN(n342) );
  XNOR2_X1 U400 ( .A(n343), .B(n342), .ZN(n344) );
  XOR2_X1 U401 ( .A(KEYINPUT7), .B(n344), .Z(n374) );
  XNOR2_X1 U402 ( .A(G22GAT), .B(KEYINPUT70), .ZN(n345) );
  XNOR2_X1 U403 ( .A(n345), .B(KEYINPUT69), .ZN(n391) );
  XOR2_X1 U404 ( .A(n391), .B(KEYINPUT29), .Z(n347) );
  NAND2_X1 U405 ( .A1(G229GAT), .A2(G233GAT), .ZN(n346) );
  XNOR2_X1 U406 ( .A(n347), .B(n346), .ZN(n348) );
  XNOR2_X1 U407 ( .A(n374), .B(n348), .ZN(n349) );
  XNOR2_X1 U408 ( .A(n350), .B(n349), .ZN(n351) );
  XOR2_X1 U409 ( .A(n352), .B(n351), .Z(n553) );
  INV_X1 U410 ( .A(n553), .ZN(n578) );
  XNOR2_X1 U411 ( .A(G204GAT), .B(G92GAT), .ZN(n353) );
  XNOR2_X1 U412 ( .A(n353), .B(G64GAT), .ZN(n425) );
  XOR2_X1 U413 ( .A(G99GAT), .B(G85GAT), .Z(n381) );
  XNOR2_X1 U414 ( .A(n425), .B(n381), .ZN(n355) );
  AND2_X1 U415 ( .A1(G230GAT), .A2(G233GAT), .ZN(n354) );
  XNOR2_X1 U416 ( .A(n355), .B(n354), .ZN(n358) );
  INV_X1 U417 ( .A(n358), .ZN(n357) );
  INV_X1 U418 ( .A(KEYINPUT32), .ZN(n356) );
  NAND2_X1 U419 ( .A1(n357), .A2(n356), .ZN(n360) );
  NAND2_X1 U420 ( .A1(n358), .A2(KEYINPUT32), .ZN(n359) );
  NAND2_X1 U421 ( .A1(n360), .A2(n359), .ZN(n363) );
  XNOR2_X1 U422 ( .A(G71GAT), .B(G78GAT), .ZN(n361) );
  XOR2_X1 U423 ( .A(n361), .B(KEYINPUT13), .Z(n390) );
  XNOR2_X1 U424 ( .A(n390), .B(KEYINPUT31), .ZN(n362) );
  XNOR2_X1 U425 ( .A(n363), .B(n362), .ZN(n367) );
  XOR2_X1 U426 ( .A(KEYINPUT71), .B(KEYINPUT33), .Z(n365) );
  XNOR2_X1 U427 ( .A(G176GAT), .B(G57GAT), .ZN(n364) );
  XOR2_X1 U428 ( .A(n365), .B(n364), .Z(n366) );
  XNOR2_X1 U429 ( .A(n367), .B(n366), .ZN(n370) );
  XOR2_X1 U430 ( .A(G120GAT), .B(G148GAT), .Z(n433) );
  XNOR2_X1 U431 ( .A(n368), .B(n433), .ZN(n369) );
  XNOR2_X1 U432 ( .A(n370), .B(n369), .ZN(n409) );
  XOR2_X1 U433 ( .A(KEYINPUT73), .B(KEYINPUT75), .Z(n372) );
  XNOR2_X1 U434 ( .A(KEYINPUT10), .B(KEYINPUT9), .ZN(n371) );
  XNOR2_X1 U435 ( .A(n372), .B(n371), .ZN(n373) );
  XNOR2_X1 U436 ( .A(n374), .B(n373), .ZN(n389) );
  XOR2_X1 U437 ( .A(KEYINPUT76), .B(KEYINPUT77), .Z(n376) );
  XNOR2_X1 U438 ( .A(G218GAT), .B(G92GAT), .ZN(n375) );
  XNOR2_X1 U439 ( .A(n376), .B(n375), .ZN(n380) );
  XOR2_X1 U440 ( .A(KEYINPUT74), .B(KEYINPUT11), .Z(n378) );
  XNOR2_X1 U441 ( .A(G134GAT), .B(G106GAT), .ZN(n377) );
  XNOR2_X1 U442 ( .A(n378), .B(n377), .ZN(n379) );
  XOR2_X1 U443 ( .A(n380), .B(n379), .Z(n387) );
  XOR2_X1 U444 ( .A(G36GAT), .B(G190GAT), .Z(n420) );
  XOR2_X1 U445 ( .A(n381), .B(n420), .Z(n385) );
  NAND2_X1 U446 ( .A1(G232GAT), .A2(G233GAT), .ZN(n382) );
  XNOR2_X1 U447 ( .A(n387), .B(n386), .ZN(n388) );
  XOR2_X1 U448 ( .A(KEYINPUT36), .B(n567), .Z(n588) );
  XNOR2_X1 U449 ( .A(n391), .B(n390), .ZN(n404) );
  XOR2_X1 U450 ( .A(KEYINPUT12), .B(KEYINPUT79), .Z(n393) );
  NAND2_X1 U451 ( .A1(G231GAT), .A2(G233GAT), .ZN(n392) );
  XNOR2_X1 U452 ( .A(n393), .B(n392), .ZN(n394) );
  XOR2_X1 U453 ( .A(n394), .B(KEYINPUT15), .Z(n399) );
  XNOR2_X1 U454 ( .A(G1GAT), .B(G155GAT), .ZN(n395) );
  XNOR2_X1 U455 ( .A(n395), .B(G57GAT), .ZN(n434) );
  XOR2_X1 U456 ( .A(KEYINPUT78), .B(G211GAT), .Z(n397) );
  XNOR2_X1 U457 ( .A(G8GAT), .B(G183GAT), .ZN(n396) );
  XNOR2_X1 U458 ( .A(n397), .B(n396), .ZN(n424) );
  XNOR2_X1 U459 ( .A(n434), .B(n424), .ZN(n398) );
  XNOR2_X1 U460 ( .A(n399), .B(n398), .ZN(n400) );
  XNOR2_X1 U461 ( .A(n401), .B(G64GAT), .ZN(n402) );
  XNOR2_X1 U462 ( .A(n295), .B(n402), .ZN(n403) );
  INV_X1 U463 ( .A(n584), .ZN(n559) );
  XOR2_X1 U464 ( .A(KEYINPUT45), .B(n405), .Z(n406) );
  NOR2_X1 U465 ( .A1(n409), .A2(n406), .ZN(n407) );
  NOR2_X1 U466 ( .A1(n578), .A2(n294), .ZN(n417) );
  XOR2_X1 U467 ( .A(KEYINPUT113), .B(n584), .Z(n565) );
  INV_X1 U468 ( .A(KEYINPUT41), .ZN(n408) );
  XNOR2_X1 U469 ( .A(n409), .B(n408), .ZN(n539) );
  AND2_X1 U470 ( .A1(n578), .A2(n539), .ZN(n410) );
  XNOR2_X1 U471 ( .A(n410), .B(KEYINPUT46), .ZN(n411) );
  NOR2_X1 U472 ( .A1(n565), .A2(n411), .ZN(n412) );
  INV_X1 U473 ( .A(n567), .ZN(n562) );
  NAND2_X1 U474 ( .A1(n412), .A2(n562), .ZN(n414) );
  XOR2_X1 U475 ( .A(KEYINPUT114), .B(KEYINPUT115), .Z(n413) );
  XNOR2_X1 U476 ( .A(n414), .B(n413), .ZN(n415) );
  XNOR2_X1 U477 ( .A(n415), .B(KEYINPUT47), .ZN(n416) );
  NOR2_X1 U478 ( .A1(n417), .A2(n416), .ZN(n419) );
  XOR2_X1 U479 ( .A(KEYINPUT94), .B(n420), .Z(n422) );
  NAND2_X1 U480 ( .A1(G226GAT), .A2(G233GAT), .ZN(n421) );
  XNOR2_X1 U481 ( .A(n422), .B(n421), .ZN(n423) );
  XOR2_X1 U482 ( .A(n424), .B(n423), .Z(n428) );
  XNOR2_X1 U483 ( .A(n426), .B(n425), .ZN(n427) );
  XNOR2_X1 U484 ( .A(n428), .B(n427), .ZN(n430) );
  XOR2_X1 U485 ( .A(n430), .B(n429), .Z(n508) );
  XNOR2_X1 U486 ( .A(KEYINPUT121), .B(n508), .ZN(n431) );
  XNOR2_X1 U487 ( .A(n432), .B(KEYINPUT54), .ZN(n451) );
  XOR2_X1 U488 ( .A(n434), .B(n433), .Z(n436) );
  NAND2_X1 U489 ( .A1(G225GAT), .A2(G233GAT), .ZN(n435) );
  XNOR2_X1 U490 ( .A(n436), .B(n435), .ZN(n437) );
  XOR2_X1 U491 ( .A(n437), .B(KEYINPUT92), .Z(n440) );
  XNOR2_X1 U492 ( .A(n438), .B(KEYINPUT6), .ZN(n439) );
  XNOR2_X1 U493 ( .A(n440), .B(n439), .ZN(n444) );
  XOR2_X1 U494 ( .A(G85GAT), .B(G162GAT), .Z(n442) );
  XNOR2_X1 U495 ( .A(G29GAT), .B(G127GAT), .ZN(n441) );
  XNOR2_X1 U496 ( .A(n442), .B(n441), .ZN(n443) );
  XOR2_X1 U497 ( .A(n444), .B(n443), .Z(n450) );
  XOR2_X1 U498 ( .A(KEYINPUT5), .B(KEYINPUT1), .Z(n446) );
  XNOR2_X1 U499 ( .A(KEYINPUT91), .B(KEYINPUT4), .ZN(n445) );
  XNOR2_X1 U500 ( .A(n446), .B(n445), .ZN(n447) );
  XNOR2_X1 U501 ( .A(n448), .B(n447), .ZN(n449) );
  XNOR2_X1 U502 ( .A(n450), .B(n449), .ZN(n468) );
  XNOR2_X1 U503 ( .A(KEYINPUT93), .B(n468), .ZN(n551) );
  INV_X1 U504 ( .A(n551), .ZN(n519) );
  NAND2_X1 U505 ( .A1(n451), .A2(n519), .ZN(n452) );
  XNOR2_X1 U506 ( .A(n452), .B(KEYINPUT65), .ZN(n574) );
  XNOR2_X1 U507 ( .A(KEYINPUT55), .B(n453), .ZN(n454) );
  NAND2_X1 U508 ( .A1(n568), .A2(n539), .ZN(n458) );
  XOR2_X1 U509 ( .A(G176GAT), .B(KEYINPUT122), .Z(n456) );
  XNOR2_X1 U510 ( .A(KEYINPUT56), .B(KEYINPUT57), .ZN(n455) );
  XOR2_X1 U511 ( .A(KEYINPUT97), .B(KEYINPUT98), .Z(n460) );
  XNOR2_X1 U512 ( .A(G1GAT), .B(KEYINPUT34), .ZN(n459) );
  XNOR2_X1 U513 ( .A(n460), .B(n459), .ZN(n479) );
  NOR2_X1 U514 ( .A1(n553), .A2(n409), .ZN(n490) );
  XOR2_X1 U515 ( .A(KEYINPUT80), .B(KEYINPUT16), .Z(n462) );
  NAND2_X1 U516 ( .A1(n584), .A2(n562), .ZN(n461) );
  XNOR2_X1 U517 ( .A(n462), .B(n461), .ZN(n477) );
  NAND2_X1 U518 ( .A1(n536), .A2(n508), .ZN(n463) );
  NAND2_X1 U519 ( .A1(n470), .A2(n463), .ZN(n464) );
  XOR2_X1 U520 ( .A(KEYINPUT25), .B(n464), .Z(n467) );
  NOR2_X1 U521 ( .A1(n470), .A2(n536), .ZN(n466) );
  XNOR2_X1 U522 ( .A(KEYINPUT26), .B(KEYINPUT96), .ZN(n465) );
  XNOR2_X1 U523 ( .A(n466), .B(n465), .ZN(n575) );
  XNOR2_X1 U524 ( .A(n508), .B(KEYINPUT27), .ZN(n472) );
  NAND2_X1 U525 ( .A1(n575), .A2(n472), .ZN(n550) );
  NAND2_X1 U526 ( .A1(n467), .A2(n550), .ZN(n469) );
  NAND2_X1 U527 ( .A1(n469), .A2(n468), .ZN(n476) );
  XNOR2_X1 U528 ( .A(n470), .B(KEYINPUT28), .ZN(n529) );
  INV_X1 U529 ( .A(n529), .ZN(n513) );
  NOR2_X1 U530 ( .A1(n519), .A2(n513), .ZN(n471) );
  NAND2_X1 U531 ( .A1(n472), .A2(n471), .ZN(n534) );
  XOR2_X1 U532 ( .A(KEYINPUT85), .B(n536), .Z(n473) );
  NOR2_X1 U533 ( .A1(n534), .A2(n473), .ZN(n474) );
  XNOR2_X1 U534 ( .A(KEYINPUT95), .B(n474), .ZN(n475) );
  NAND2_X1 U535 ( .A1(n476), .A2(n475), .ZN(n486) );
  AND2_X1 U536 ( .A1(n477), .A2(n486), .ZN(n503) );
  NAND2_X1 U537 ( .A1(n490), .A2(n503), .ZN(n484) );
  NOR2_X1 U538 ( .A1(n519), .A2(n484), .ZN(n478) );
  XOR2_X1 U539 ( .A(n479), .B(n478), .Z(G1324GAT) );
  INV_X1 U540 ( .A(n508), .ZN(n522) );
  NOR2_X1 U541 ( .A1(n522), .A2(n484), .ZN(n481) );
  XNOR2_X1 U542 ( .A(G8GAT), .B(KEYINPUT99), .ZN(n480) );
  XNOR2_X1 U543 ( .A(n481), .B(n480), .ZN(G1325GAT) );
  NOR2_X1 U544 ( .A1(n524), .A2(n484), .ZN(n483) );
  XNOR2_X1 U545 ( .A(G15GAT), .B(KEYINPUT35), .ZN(n482) );
  XNOR2_X1 U546 ( .A(n483), .B(n482), .ZN(G1326GAT) );
  NOR2_X1 U547 ( .A1(n529), .A2(n484), .ZN(n485) );
  XOR2_X1 U548 ( .A(G22GAT), .B(n485), .Z(G1327GAT) );
  XNOR2_X1 U549 ( .A(KEYINPUT100), .B(KEYINPUT39), .ZN(n493) );
  NAND2_X1 U550 ( .A1(n559), .A2(n486), .ZN(n487) );
  XOR2_X1 U551 ( .A(KEYINPUT101), .B(n487), .Z(n488) );
  NOR2_X1 U552 ( .A1(n588), .A2(n488), .ZN(n489) );
  XOR2_X1 U553 ( .A(KEYINPUT37), .B(n489), .Z(n518) );
  NAND2_X1 U554 ( .A1(n518), .A2(n490), .ZN(n491) );
  XNOR2_X1 U555 ( .A(KEYINPUT38), .B(n491), .ZN(n501) );
  NOR2_X1 U556 ( .A1(n519), .A2(n501), .ZN(n492) );
  XNOR2_X1 U557 ( .A(n493), .B(n492), .ZN(n494) );
  XNOR2_X1 U558 ( .A(G29GAT), .B(n494), .ZN(G1328GAT) );
  NOR2_X1 U559 ( .A1(n522), .A2(n501), .ZN(n495) );
  XOR2_X1 U560 ( .A(KEYINPUT102), .B(n495), .Z(n496) );
  XNOR2_X1 U561 ( .A(G36GAT), .B(n496), .ZN(G1329GAT) );
  XOR2_X1 U562 ( .A(KEYINPUT40), .B(KEYINPUT104), .Z(n498) );
  XNOR2_X1 U563 ( .A(G43GAT), .B(KEYINPUT103), .ZN(n497) );
  XNOR2_X1 U564 ( .A(n498), .B(n497), .ZN(n500) );
  NOR2_X1 U565 ( .A1(n524), .A2(n501), .ZN(n499) );
  XOR2_X1 U566 ( .A(n500), .B(n499), .Z(G1330GAT) );
  NOR2_X1 U567 ( .A1(n501), .A2(n529), .ZN(n502) );
  XOR2_X1 U568 ( .A(G50GAT), .B(n502), .Z(G1331GAT) );
  INV_X1 U569 ( .A(n539), .ZN(n555) );
  NOR2_X1 U570 ( .A1(n578), .A2(n555), .ZN(n517) );
  NAND2_X1 U571 ( .A1(n517), .A2(n503), .ZN(n504) );
  XOR2_X1 U572 ( .A(KEYINPUT106), .B(n504), .Z(n512) );
  NAND2_X1 U573 ( .A1(n512), .A2(n551), .ZN(n507) );
  XOR2_X1 U574 ( .A(G57GAT), .B(KEYINPUT105), .Z(n505) );
  XNOR2_X1 U575 ( .A(KEYINPUT42), .B(n505), .ZN(n506) );
  XNOR2_X1 U576 ( .A(n507), .B(n506), .ZN(G1332GAT) );
  XOR2_X1 U577 ( .A(G64GAT), .B(KEYINPUT107), .Z(n510) );
  NAND2_X1 U578 ( .A1(n512), .A2(n508), .ZN(n509) );
  XNOR2_X1 U579 ( .A(n510), .B(n509), .ZN(G1333GAT) );
  NAND2_X1 U580 ( .A1(n512), .A2(n536), .ZN(n511) );
  XNOR2_X1 U581 ( .A(n511), .B(G71GAT), .ZN(G1334GAT) );
  XOR2_X1 U582 ( .A(KEYINPUT108), .B(KEYINPUT43), .Z(n515) );
  NAND2_X1 U583 ( .A1(n513), .A2(n512), .ZN(n514) );
  XNOR2_X1 U584 ( .A(n515), .B(n514), .ZN(n516) );
  XNOR2_X1 U585 ( .A(G78GAT), .B(n516), .ZN(G1335GAT) );
  NAND2_X1 U586 ( .A1(n518), .A2(n517), .ZN(n528) );
  NOR2_X1 U587 ( .A1(n519), .A2(n528), .ZN(n521) );
  XNOR2_X1 U588 ( .A(G85GAT), .B(KEYINPUT109), .ZN(n520) );
  XNOR2_X1 U589 ( .A(n521), .B(n520), .ZN(G1336GAT) );
  NOR2_X1 U590 ( .A1(n522), .A2(n528), .ZN(n523) );
  XOR2_X1 U591 ( .A(G92GAT), .B(n523), .Z(G1337GAT) );
  NOR2_X1 U592 ( .A1(n524), .A2(n528), .ZN(n526) );
  XNOR2_X1 U593 ( .A(KEYINPUT110), .B(KEYINPUT111), .ZN(n525) );
  XNOR2_X1 U594 ( .A(n526), .B(n525), .ZN(n527) );
  XNOR2_X1 U595 ( .A(G99GAT), .B(n527), .ZN(G1338GAT) );
  NOR2_X1 U596 ( .A1(n529), .A2(n528), .ZN(n531) );
  XNOR2_X1 U597 ( .A(KEYINPUT44), .B(KEYINPUT112), .ZN(n530) );
  XNOR2_X1 U598 ( .A(n531), .B(n530), .ZN(n532) );
  XOR2_X1 U599 ( .A(G106GAT), .B(n532), .Z(G1339GAT) );
  NOR2_X1 U600 ( .A1(n533), .A2(n534), .ZN(n535) );
  NAND2_X1 U601 ( .A1(n536), .A2(n535), .ZN(n537) );
  XNOR2_X1 U602 ( .A(n537), .B(KEYINPUT117), .ZN(n546) );
  NAND2_X1 U603 ( .A1(n578), .A2(n546), .ZN(n538) );
  XNOR2_X1 U604 ( .A(n538), .B(G113GAT), .ZN(G1340GAT) );
  XOR2_X1 U605 ( .A(KEYINPUT118), .B(KEYINPUT49), .Z(n541) );
  NAND2_X1 U606 ( .A1(n546), .A2(n539), .ZN(n540) );
  XNOR2_X1 U607 ( .A(n541), .B(n540), .ZN(n542) );
  XNOR2_X1 U608 ( .A(G120GAT), .B(n542), .ZN(G1341GAT) );
  XOR2_X1 U609 ( .A(KEYINPUT50), .B(KEYINPUT119), .Z(n544) );
  NAND2_X1 U610 ( .A1(n546), .A2(n565), .ZN(n543) );
  XNOR2_X1 U611 ( .A(n544), .B(n543), .ZN(n545) );
  XNOR2_X1 U612 ( .A(G127GAT), .B(n545), .ZN(G1342GAT) );
  XOR2_X1 U613 ( .A(KEYINPUT120), .B(KEYINPUT51), .Z(n548) );
  NAND2_X1 U614 ( .A1(n546), .A2(n567), .ZN(n547) );
  XNOR2_X1 U615 ( .A(n548), .B(n547), .ZN(n549) );
  XNOR2_X1 U616 ( .A(G134GAT), .B(n549), .ZN(G1343GAT) );
  NOR2_X1 U617 ( .A1(n533), .A2(n550), .ZN(n552) );
  NAND2_X1 U618 ( .A1(n552), .A2(n551), .ZN(n561) );
  NOR2_X1 U619 ( .A1(n553), .A2(n561), .ZN(n554) );
  XOR2_X1 U620 ( .A(G141GAT), .B(n554), .Z(G1344GAT) );
  NOR2_X1 U621 ( .A1(n555), .A2(n561), .ZN(n557) );
  XNOR2_X1 U622 ( .A(KEYINPUT53), .B(KEYINPUT52), .ZN(n556) );
  XNOR2_X1 U623 ( .A(n557), .B(n556), .ZN(n558) );
  XNOR2_X1 U624 ( .A(G148GAT), .B(n558), .ZN(G1345GAT) );
  NOR2_X1 U625 ( .A1(n559), .A2(n561), .ZN(n560) );
  XOR2_X1 U626 ( .A(G155GAT), .B(n560), .Z(G1346GAT) );
  NOR2_X1 U627 ( .A1(n562), .A2(n561), .ZN(n563) );
  XOR2_X1 U628 ( .A(G162GAT), .B(n563), .Z(G1347GAT) );
  NAND2_X1 U629 ( .A1(n578), .A2(n568), .ZN(n564) );
  XNOR2_X1 U630 ( .A(n564), .B(G169GAT), .ZN(G1348GAT) );
  NAND2_X1 U631 ( .A1(n568), .A2(n565), .ZN(n566) );
  XNOR2_X1 U632 ( .A(n566), .B(G183GAT), .ZN(G1350GAT) );
  XNOR2_X1 U633 ( .A(G190GAT), .B(KEYINPUT58), .ZN(n570) );
  NAND2_X1 U634 ( .A1(n568), .A2(n567), .ZN(n569) );
  XNOR2_X1 U635 ( .A(n570), .B(n569), .ZN(G1351GAT) );
  XOR2_X1 U636 ( .A(KEYINPUT60), .B(KEYINPUT125), .Z(n572) );
  XNOR2_X1 U637 ( .A(G197GAT), .B(KEYINPUT124), .ZN(n571) );
  XNOR2_X1 U638 ( .A(n572), .B(n571), .ZN(n573) );
  XOR2_X1 U639 ( .A(KEYINPUT59), .B(n573), .Z(n580) );
  NAND2_X1 U640 ( .A1(n575), .A2(n574), .ZN(n577) );
  INV_X1 U641 ( .A(KEYINPUT123), .ZN(n576) );
  XNOR2_X1 U642 ( .A(n577), .B(n576), .ZN(n589) );
  INV_X1 U643 ( .A(n589), .ZN(n585) );
  NAND2_X1 U644 ( .A1(n585), .A2(n578), .ZN(n579) );
  XNOR2_X1 U645 ( .A(n580), .B(n579), .ZN(G1352GAT) );
  XOR2_X1 U646 ( .A(KEYINPUT126), .B(KEYINPUT61), .Z(n582) );
  NAND2_X1 U647 ( .A1(n585), .A2(n409), .ZN(n581) );
  XNOR2_X1 U648 ( .A(n582), .B(n581), .ZN(n583) );
  XNOR2_X1 U649 ( .A(G204GAT), .B(n583), .ZN(G1353GAT) );
  XOR2_X1 U650 ( .A(G211GAT), .B(KEYINPUT127), .Z(n587) );
  NAND2_X1 U651 ( .A1(n585), .A2(n584), .ZN(n586) );
  XNOR2_X1 U652 ( .A(n587), .B(n586), .ZN(G1354GAT) );
  INV_X1 U653 ( .A(KEYINPUT62), .ZN(n591) );
  NOR2_X1 U654 ( .A1(n589), .A2(n588), .ZN(n590) );
  XNOR2_X1 U655 ( .A(n591), .B(n590), .ZN(n592) );
  XNOR2_X1 U656 ( .A(G218GAT), .B(n592), .ZN(G1355GAT) );
endmodule

