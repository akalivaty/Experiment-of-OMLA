//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 0 1 0 1 1 0 1 1 1 0 1 1 1 1 1 0 1 1 0 0 0 0 0 0 1 0 0 0 0 0 1 1 0 1 0 1 1 0 1 1 1 1 0 0 0 0 0 1 1 0 0 1 1 1 0 0 1 1 0 1 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:36:58 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n245, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1193,
    new_n1194, new_n1195, new_n1196, new_n1197, new_n1198, new_n1199,
    new_n1200, new_n1201, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1216, new_n1217, new_n1218,
    new_n1219, new_n1221, new_n1222, new_n1223, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1285, new_n1286, new_n1287,
    new_n1288, new_n1289;
  INV_X1    g0000(.A(G50), .ZN(new_n201));
  INV_X1    g0001(.A(G58), .ZN(new_n202));
  INV_X1    g0002(.A(G68), .ZN(new_n203));
  NAND3_X1  g0003(.A1(new_n201), .A2(new_n202), .A3(new_n203), .ZN(new_n204));
  NOR2_X1   g0004(.A1(new_n204), .A2(G77), .ZN(G353));
  OAI21_X1  g0005(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0006(.A(G1), .ZN(new_n207));
  INV_X1    g0007(.A(G20), .ZN(new_n208));
  NOR2_X1   g0008(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  INV_X1    g0009(.A(new_n209), .ZN(new_n210));
  NOR2_X1   g0010(.A1(new_n210), .A2(G13), .ZN(new_n211));
  OAI211_X1 g0011(.A(new_n211), .B(G250), .C1(G257), .C2(G264), .ZN(new_n212));
  XNOR2_X1  g0012(.A(new_n212), .B(KEYINPUT0), .ZN(new_n213));
  NAND2_X1  g0013(.A1(G1), .A2(G13), .ZN(new_n214));
  INV_X1    g0014(.A(new_n214), .ZN(new_n215));
  NAND2_X1  g0015(.A1(new_n215), .A2(G20), .ZN(new_n216));
  OAI21_X1  g0016(.A(G50), .B1(G58), .B2(G68), .ZN(new_n217));
  AOI22_X1  g0017(.A1(G107), .A2(G264), .B1(G116), .B2(G270), .ZN(new_n218));
  INV_X1    g0018(.A(G77), .ZN(new_n219));
  INV_X1    g0019(.A(G244), .ZN(new_n220));
  INV_X1    g0020(.A(G87), .ZN(new_n221));
  INV_X1    g0021(.A(G250), .ZN(new_n222));
  OAI221_X1 g0022(.A(new_n218), .B1(new_n219), .B2(new_n220), .C1(new_n221), .C2(new_n222), .ZN(new_n223));
  AOI22_X1  g0023(.A1(G50), .A2(G226), .B1(G97), .B2(G257), .ZN(new_n224));
  INV_X1    g0024(.A(G232), .ZN(new_n225));
  INV_X1    g0025(.A(G238), .ZN(new_n226));
  OAI221_X1 g0026(.A(new_n224), .B1(new_n202), .B2(new_n225), .C1(new_n203), .C2(new_n226), .ZN(new_n227));
  OAI21_X1  g0027(.A(new_n210), .B1(new_n223), .B2(new_n227), .ZN(new_n228));
  OAI221_X1 g0028(.A(new_n213), .B1(new_n216), .B2(new_n217), .C1(KEYINPUT1), .C2(new_n228), .ZN(new_n229));
  AOI21_X1  g0029(.A(new_n229), .B1(KEYINPUT1), .B2(new_n228), .ZN(G361));
  XNOR2_X1  g0030(.A(G238), .B(G244), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n231), .B(KEYINPUT2), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n232), .B(G226), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n233), .B(new_n225), .ZN(new_n234));
  XNOR2_X1  g0034(.A(G250), .B(G257), .ZN(new_n235));
  XNOR2_X1  g0035(.A(G264), .B(G270), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n234), .B(new_n237), .ZN(G358));
  XOR2_X1   g0038(.A(G50), .B(G58), .Z(new_n239));
  XNOR2_X1  g0039(.A(new_n239), .B(KEYINPUT64), .ZN(new_n240));
  XNOR2_X1  g0040(.A(G68), .B(G77), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XOR2_X1   g0042(.A(G87), .B(G97), .Z(new_n243));
  XNOR2_X1  g0043(.A(G107), .B(G116), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XOR2_X1   g0045(.A(new_n242), .B(new_n245), .Z(G351));
  NAND3_X1  g0046(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n247));
  NAND2_X1  g0047(.A1(new_n247), .A2(new_n214), .ZN(new_n248));
  INV_X1    g0048(.A(new_n248), .ZN(new_n249));
  INV_X1    g0049(.A(KEYINPUT68), .ZN(new_n250));
  INV_X1    g0050(.A(G33), .ZN(new_n251));
  NAND3_X1  g0051(.A1(new_n250), .A2(new_n208), .A3(new_n251), .ZN(new_n252));
  OAI21_X1  g0052(.A(KEYINPUT68), .B1(G20), .B2(G33), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n252), .A2(new_n253), .ZN(new_n254));
  NAND2_X1  g0054(.A1(new_n254), .A2(G50), .ZN(new_n255));
  XOR2_X1   g0055(.A(new_n255), .B(KEYINPUT71), .Z(new_n256));
  OAI21_X1  g0056(.A(KEYINPUT67), .B1(new_n251), .B2(G20), .ZN(new_n257));
  INV_X1    g0057(.A(KEYINPUT67), .ZN(new_n258));
  NAND3_X1  g0058(.A1(new_n258), .A2(new_n208), .A3(G33), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n257), .A2(new_n259), .ZN(new_n260));
  INV_X1    g0060(.A(new_n260), .ZN(new_n261));
  AOI22_X1  g0061(.A1(new_n261), .A2(G77), .B1(G20), .B2(new_n203), .ZN(new_n262));
  AOI21_X1  g0062(.A(new_n249), .B1(new_n256), .B2(new_n262), .ZN(new_n263));
  OR2_X1    g0063(.A1(new_n263), .A2(KEYINPUT11), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n263), .A2(KEYINPUT11), .ZN(new_n265));
  NAND3_X1  g0065(.A1(new_n207), .A2(G13), .A3(G20), .ZN(new_n266));
  INV_X1    g0066(.A(new_n266), .ZN(new_n267));
  AOI21_X1  g0067(.A(KEYINPUT12), .B1(new_n267), .B2(new_n203), .ZN(new_n268));
  AND3_X1   g0068(.A1(new_n267), .A2(KEYINPUT12), .A3(new_n203), .ZN(new_n269));
  AOI21_X1  g0069(.A(new_n248), .B1(new_n207), .B2(G20), .ZN(new_n270));
  AOI211_X1 g0070(.A(new_n268), .B(new_n269), .C1(G68), .C2(new_n270), .ZN(new_n271));
  NAND3_X1  g0071(.A1(new_n264), .A2(new_n265), .A3(new_n271), .ZN(new_n272));
  INV_X1    g0072(.A(new_n272), .ZN(new_n273));
  INV_X1    g0073(.A(KEYINPUT72), .ZN(new_n274));
  INV_X1    g0074(.A(KEYINPUT70), .ZN(new_n275));
  INV_X1    g0075(.A(KEYINPUT3), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n276), .A2(new_n251), .ZN(new_n277));
  NAND2_X1  g0077(.A1(KEYINPUT3), .A2(G33), .ZN(new_n278));
  INV_X1    g0078(.A(G1698), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n279), .A2(G226), .ZN(new_n280));
  NAND2_X1  g0080(.A1(G232), .A2(G1698), .ZN(new_n281));
  AOI22_X1  g0081(.A1(new_n277), .A2(new_n278), .B1(new_n280), .B2(new_n281), .ZN(new_n282));
  NAND2_X1  g0082(.A1(G33), .A2(G97), .ZN(new_n283));
  INV_X1    g0083(.A(new_n283), .ZN(new_n284));
  OAI21_X1  g0084(.A(new_n275), .B1(new_n282), .B2(new_n284), .ZN(new_n285));
  AND2_X1   g0085(.A1(new_n280), .A2(new_n281), .ZN(new_n286));
  AND2_X1   g0086(.A1(KEYINPUT3), .A2(G33), .ZN(new_n287));
  NOR2_X1   g0087(.A1(KEYINPUT3), .A2(G33), .ZN(new_n288));
  NOR2_X1   g0088(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  OAI211_X1 g0089(.A(KEYINPUT70), .B(new_n283), .C1(new_n286), .C2(new_n289), .ZN(new_n290));
  NAND2_X1  g0090(.A1(G33), .A2(G41), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n215), .A2(new_n291), .ZN(new_n292));
  INV_X1    g0092(.A(new_n292), .ZN(new_n293));
  NAND3_X1  g0093(.A1(new_n285), .A2(new_n290), .A3(new_n293), .ZN(new_n294));
  INV_X1    g0094(.A(KEYINPUT13), .ZN(new_n295));
  AND2_X1   g0095(.A1(G33), .A2(G41), .ZN(new_n296));
  OAI21_X1  g0096(.A(KEYINPUT65), .B1(new_n296), .B2(new_n214), .ZN(new_n297));
  INV_X1    g0097(.A(KEYINPUT65), .ZN(new_n298));
  NAND4_X1  g0098(.A1(new_n291), .A2(new_n298), .A3(G1), .A4(G13), .ZN(new_n299));
  OAI21_X1  g0099(.A(new_n207), .B1(G41), .B2(G45), .ZN(new_n300));
  NAND4_X1  g0100(.A1(new_n297), .A2(G238), .A3(new_n299), .A4(new_n300), .ZN(new_n301));
  INV_X1    g0101(.A(new_n300), .ZN(new_n302));
  NAND4_X1  g0102(.A1(new_n297), .A2(new_n302), .A3(G274), .A4(new_n299), .ZN(new_n303));
  AND2_X1   g0103(.A1(new_n301), .A2(new_n303), .ZN(new_n304));
  AND3_X1   g0104(.A1(new_n294), .A2(new_n295), .A3(new_n304), .ZN(new_n305));
  AOI21_X1  g0105(.A(new_n295), .B1(new_n294), .B2(new_n304), .ZN(new_n306));
  NOR2_X1   g0106(.A1(new_n305), .A2(new_n306), .ZN(new_n307));
  AOI21_X1  g0107(.A(new_n274), .B1(new_n307), .B2(G179), .ZN(new_n308));
  INV_X1    g0108(.A(G179), .ZN(new_n309));
  NOR4_X1   g0109(.A1(new_n305), .A2(new_n306), .A3(KEYINPUT72), .A4(new_n309), .ZN(new_n310));
  NOR2_X1   g0110(.A1(new_n308), .A2(new_n310), .ZN(new_n311));
  OAI21_X1  g0111(.A(G169), .B1(new_n305), .B2(new_n306), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n312), .A2(KEYINPUT14), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n294), .A2(new_n304), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n314), .A2(KEYINPUT13), .ZN(new_n315));
  NAND3_X1  g0115(.A1(new_n294), .A2(new_n295), .A3(new_n304), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n315), .A2(new_n316), .ZN(new_n317));
  INV_X1    g0117(.A(KEYINPUT14), .ZN(new_n318));
  NAND3_X1  g0118(.A1(new_n317), .A2(new_n318), .A3(G169), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n313), .A2(new_n319), .ZN(new_n320));
  OAI21_X1  g0120(.A(KEYINPUT73), .B1(new_n311), .B2(new_n320), .ZN(new_n321));
  OAI21_X1  g0121(.A(KEYINPUT72), .B1(new_n317), .B2(new_n309), .ZN(new_n322));
  NAND3_X1  g0122(.A1(new_n307), .A2(new_n274), .A3(G179), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  INV_X1    g0124(.A(KEYINPUT73), .ZN(new_n325));
  NAND4_X1  g0125(.A1(new_n324), .A2(new_n325), .A3(new_n313), .A4(new_n319), .ZN(new_n326));
  AOI21_X1  g0126(.A(new_n273), .B1(new_n321), .B2(new_n326), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n307), .A2(G190), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n317), .A2(G200), .ZN(new_n329));
  NAND3_X1  g0129(.A1(new_n273), .A2(new_n328), .A3(new_n329), .ZN(new_n330));
  INV_X1    g0130(.A(new_n330), .ZN(new_n331));
  NOR2_X1   g0131(.A1(new_n327), .A2(new_n331), .ZN(new_n332));
  AND2_X1   g0132(.A1(new_n297), .A2(new_n299), .ZN(new_n333));
  NAND3_X1  g0133(.A1(new_n333), .A2(G226), .A3(new_n300), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n277), .A2(new_n278), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n279), .A2(G222), .ZN(new_n336));
  NAND2_X1  g0136(.A1(G223), .A2(G1698), .ZN(new_n337));
  NAND3_X1  g0137(.A1(new_n335), .A2(new_n336), .A3(new_n337), .ZN(new_n338));
  OAI211_X1 g0138(.A(new_n338), .B(new_n293), .C1(G77), .C2(new_n335), .ZN(new_n339));
  NAND3_X1  g0139(.A1(new_n334), .A2(new_n339), .A3(new_n303), .ZN(new_n340));
  AND2_X1   g0140(.A1(new_n340), .A2(G200), .ZN(new_n341));
  INV_X1    g0141(.A(G190), .ZN(new_n342));
  NOR2_X1   g0142(.A1(new_n340), .A2(new_n342), .ZN(new_n343));
  NOR2_X1   g0143(.A1(new_n341), .A2(new_n343), .ZN(new_n344));
  XNOR2_X1  g0144(.A(KEYINPUT8), .B(G58), .ZN(new_n345));
  INV_X1    g0145(.A(KEYINPUT66), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n345), .A2(new_n346), .ZN(new_n347));
  NAND3_X1  g0147(.A1(new_n202), .A2(KEYINPUT66), .A3(KEYINPUT8), .ZN(new_n348));
  NAND3_X1  g0148(.A1(new_n261), .A2(new_n347), .A3(new_n348), .ZN(new_n349));
  AOI22_X1  g0149(.A1(new_n254), .A2(G150), .B1(G20), .B2(new_n204), .ZN(new_n350));
  AOI21_X1  g0150(.A(new_n249), .B1(new_n349), .B2(new_n350), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n267), .A2(new_n201), .ZN(new_n352));
  INV_X1    g0152(.A(new_n270), .ZN(new_n353));
  OAI21_X1  g0153(.A(new_n352), .B1(new_n353), .B2(new_n201), .ZN(new_n354));
  NOR2_X1   g0154(.A1(new_n351), .A2(new_n354), .ZN(new_n355));
  INV_X1    g0155(.A(KEYINPUT9), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n355), .A2(new_n356), .ZN(new_n357));
  OAI21_X1  g0157(.A(KEYINPUT9), .B1(new_n351), .B2(new_n354), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n357), .A2(new_n358), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n344), .A2(new_n359), .ZN(new_n360));
  OAI211_X1 g0160(.A(new_n360), .B(KEYINPUT10), .C1(KEYINPUT69), .C2(new_n341), .ZN(new_n361));
  OAI21_X1  g0161(.A(KEYINPUT10), .B1(new_n341), .B2(KEYINPUT69), .ZN(new_n362));
  NAND3_X1  g0162(.A1(new_n362), .A2(new_n359), .A3(new_n344), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n361), .A2(new_n363), .ZN(new_n364));
  NOR2_X1   g0164(.A1(new_n340), .A2(G179), .ZN(new_n365));
  INV_X1    g0165(.A(G169), .ZN(new_n366));
  AOI211_X1 g0166(.A(new_n355), .B(new_n365), .C1(new_n366), .C2(new_n340), .ZN(new_n367));
  INV_X1    g0167(.A(new_n367), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n364), .A2(new_n368), .ZN(new_n369));
  INV_X1    g0169(.A(KEYINPUT17), .ZN(new_n370));
  NAND4_X1  g0170(.A1(new_n297), .A2(G232), .A3(new_n299), .A4(new_n300), .ZN(new_n371));
  NOR2_X1   g0171(.A1(new_n251), .A2(new_n221), .ZN(new_n372));
  NOR2_X1   g0172(.A1(G223), .A2(G1698), .ZN(new_n373));
  INV_X1    g0173(.A(G226), .ZN(new_n374));
  AOI21_X1  g0174(.A(new_n373), .B1(new_n374), .B2(G1698), .ZN(new_n375));
  AOI21_X1  g0175(.A(new_n372), .B1(new_n375), .B2(new_n335), .ZN(new_n376));
  OAI211_X1 g0176(.A(new_n303), .B(new_n371), .C1(new_n376), .C2(new_n292), .ZN(new_n377));
  INV_X1    g0177(.A(G200), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n377), .A2(new_n378), .ZN(new_n379));
  OAI21_X1  g0179(.A(KEYINPUT75), .B1(new_n376), .B2(new_n292), .ZN(new_n380));
  OR2_X1    g0180(.A1(G223), .A2(G1698), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n374), .A2(G1698), .ZN(new_n382));
  OAI211_X1 g0182(.A(new_n381), .B(new_n382), .C1(new_n287), .C2(new_n288), .ZN(new_n383));
  INV_X1    g0183(.A(new_n372), .ZN(new_n384));
  AOI21_X1  g0184(.A(new_n292), .B1(new_n383), .B2(new_n384), .ZN(new_n385));
  INV_X1    g0185(.A(KEYINPUT75), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n385), .A2(new_n386), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n380), .A2(new_n387), .ZN(new_n388));
  NAND3_X1  g0188(.A1(new_n303), .A2(new_n371), .A3(new_n342), .ZN(new_n389));
  OAI21_X1  g0189(.A(new_n379), .B1(new_n388), .B2(new_n389), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n347), .A2(new_n348), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n391), .A2(new_n267), .ZN(new_n392));
  OAI21_X1  g0192(.A(new_n392), .B1(new_n353), .B2(new_n391), .ZN(new_n393));
  INV_X1    g0193(.A(new_n393), .ZN(new_n394));
  INV_X1    g0194(.A(KEYINPUT74), .ZN(new_n395));
  NAND3_X1  g0195(.A1(new_n277), .A2(new_n208), .A3(new_n278), .ZN(new_n396));
  INV_X1    g0196(.A(KEYINPUT7), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n396), .A2(new_n397), .ZN(new_n398));
  NAND4_X1  g0198(.A1(new_n277), .A2(KEYINPUT7), .A3(new_n208), .A4(new_n278), .ZN(new_n399));
  AOI21_X1  g0199(.A(new_n395), .B1(new_n398), .B2(new_n399), .ZN(new_n400));
  AOI21_X1  g0200(.A(KEYINPUT74), .B1(new_n396), .B2(new_n397), .ZN(new_n401));
  OAI21_X1  g0201(.A(G68), .B1(new_n400), .B2(new_n401), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n254), .A2(G159), .ZN(new_n403));
  XNOR2_X1  g0203(.A(G58), .B(G68), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n404), .A2(G20), .ZN(new_n405));
  AND2_X1   g0205(.A1(new_n403), .A2(new_n405), .ZN(new_n406));
  AOI21_X1  g0206(.A(KEYINPUT16), .B1(new_n402), .B2(new_n406), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n398), .A2(new_n399), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n408), .A2(G68), .ZN(new_n409));
  NAND3_X1  g0209(.A1(new_n409), .A2(KEYINPUT16), .A3(new_n406), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n410), .A2(new_n248), .ZN(new_n411));
  OAI211_X1 g0211(.A(new_n390), .B(new_n394), .C1(new_n407), .C2(new_n411), .ZN(new_n412));
  INV_X1    g0212(.A(KEYINPUT76), .ZN(new_n413));
  OAI21_X1  g0213(.A(new_n370), .B1(new_n412), .B2(new_n413), .ZN(new_n414));
  INV_X1    g0214(.A(KEYINPUT16), .ZN(new_n415));
  AOI21_X1  g0215(.A(KEYINPUT7), .B1(new_n289), .B2(new_n208), .ZN(new_n416));
  INV_X1    g0216(.A(new_n399), .ZN(new_n417));
  OAI21_X1  g0217(.A(KEYINPUT74), .B1(new_n416), .B2(new_n417), .ZN(new_n418));
  INV_X1    g0218(.A(new_n401), .ZN(new_n419));
  AOI21_X1  g0219(.A(new_n203), .B1(new_n418), .B2(new_n419), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n403), .A2(new_n405), .ZN(new_n421));
  OAI21_X1  g0221(.A(new_n415), .B1(new_n420), .B2(new_n421), .ZN(new_n422));
  AOI21_X1  g0222(.A(new_n421), .B1(G68), .B2(new_n408), .ZN(new_n423));
  AOI21_X1  g0223(.A(new_n249), .B1(new_n423), .B2(KEYINPUT16), .ZN(new_n424));
  AOI21_X1  g0224(.A(new_n393), .B1(new_n422), .B2(new_n424), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n377), .A2(new_n366), .ZN(new_n426));
  NAND3_X1  g0226(.A1(new_n303), .A2(new_n371), .A3(new_n309), .ZN(new_n427));
  OAI21_X1  g0227(.A(new_n426), .B1(new_n388), .B2(new_n427), .ZN(new_n428));
  OAI21_X1  g0228(.A(KEYINPUT18), .B1(new_n425), .B2(new_n428), .ZN(new_n429));
  NAND4_X1  g0229(.A1(new_n425), .A2(KEYINPUT76), .A3(KEYINPUT17), .A4(new_n390), .ZN(new_n430));
  OAI21_X1  g0230(.A(new_n394), .B1(new_n407), .B2(new_n411), .ZN(new_n431));
  INV_X1    g0231(.A(KEYINPUT18), .ZN(new_n432));
  INV_X1    g0232(.A(new_n428), .ZN(new_n433));
  NAND3_X1  g0233(.A1(new_n431), .A2(new_n432), .A3(new_n433), .ZN(new_n434));
  NAND4_X1  g0234(.A1(new_n414), .A2(new_n429), .A3(new_n430), .A4(new_n434), .ZN(new_n435));
  INV_X1    g0235(.A(new_n345), .ZN(new_n436));
  AOI22_X1  g0236(.A1(new_n436), .A2(new_n254), .B1(G20), .B2(G77), .ZN(new_n437));
  XNOR2_X1  g0237(.A(KEYINPUT15), .B(G87), .ZN(new_n438));
  OAI21_X1  g0238(.A(new_n437), .B1(new_n260), .B2(new_n438), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n439), .A2(new_n248), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n270), .A2(G77), .ZN(new_n441));
  OAI211_X1 g0241(.A(new_n440), .B(new_n441), .C1(G77), .C2(new_n266), .ZN(new_n442));
  NAND2_X1  g0242(.A1(G238), .A2(G1698), .ZN(new_n443));
  OAI211_X1 g0243(.A(new_n335), .B(new_n443), .C1(new_n225), .C2(G1698), .ZN(new_n444));
  OAI211_X1 g0244(.A(new_n444), .B(new_n293), .C1(G107), .C2(new_n335), .ZN(new_n445));
  NAND3_X1  g0245(.A1(new_n333), .A2(G244), .A3(new_n300), .ZN(new_n446));
  NAND3_X1  g0246(.A1(new_n445), .A2(new_n303), .A3(new_n446), .ZN(new_n447));
  AND2_X1   g0247(.A1(new_n447), .A2(G200), .ZN(new_n448));
  NOR2_X1   g0248(.A1(new_n442), .A2(new_n448), .ZN(new_n449));
  OAI21_X1  g0249(.A(new_n449), .B1(new_n342), .B2(new_n447), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n447), .A2(new_n366), .ZN(new_n451));
  NAND4_X1  g0251(.A1(new_n445), .A2(new_n446), .A3(new_n309), .A4(new_n303), .ZN(new_n452));
  NAND3_X1  g0252(.A1(new_n442), .A2(new_n451), .A3(new_n452), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n450), .A2(new_n453), .ZN(new_n454));
  NOR3_X1   g0254(.A1(new_n369), .A2(new_n435), .A3(new_n454), .ZN(new_n455));
  AND2_X1   g0255(.A1(new_n332), .A2(new_n455), .ZN(new_n456));
  INV_X1    g0256(.A(KEYINPUT19), .ZN(new_n457));
  INV_X1    g0257(.A(G97), .ZN(new_n458));
  OAI21_X1  g0258(.A(new_n457), .B1(new_n260), .B2(new_n458), .ZN(new_n459));
  NAND3_X1  g0259(.A1(new_n335), .A2(new_n208), .A3(G68), .ZN(new_n460));
  OAI21_X1  g0260(.A(new_n208), .B1(new_n283), .B2(new_n457), .ZN(new_n461));
  INV_X1    g0261(.A(KEYINPUT82), .ZN(new_n462));
  INV_X1    g0262(.A(G107), .ZN(new_n463));
  NAND3_X1  g0263(.A1(new_n221), .A2(new_n458), .A3(new_n463), .ZN(new_n464));
  NAND3_X1  g0264(.A1(new_n461), .A2(new_n462), .A3(new_n464), .ZN(new_n465));
  INV_X1    g0265(.A(new_n465), .ZN(new_n466));
  AOI21_X1  g0266(.A(new_n462), .B1(new_n461), .B2(new_n464), .ZN(new_n467));
  OAI211_X1 g0267(.A(new_n459), .B(new_n460), .C1(new_n466), .C2(new_n467), .ZN(new_n468));
  INV_X1    g0268(.A(KEYINPUT83), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  INV_X1    g0270(.A(new_n467), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n471), .A2(new_n465), .ZN(new_n472));
  NAND4_X1  g0272(.A1(new_n472), .A2(KEYINPUT83), .A3(new_n460), .A4(new_n459), .ZN(new_n473));
  NAND3_X1  g0273(.A1(new_n470), .A2(new_n473), .A3(new_n248), .ZN(new_n474));
  INV_X1    g0274(.A(new_n438), .ZN(new_n475));
  NOR2_X1   g0275(.A1(new_n475), .A2(new_n266), .ZN(new_n476));
  INV_X1    g0276(.A(new_n476), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n207), .A2(G33), .ZN(new_n478));
  NAND4_X1  g0278(.A1(new_n266), .A2(new_n478), .A3(new_n214), .A4(new_n247), .ZN(new_n479));
  OR2_X1    g0279(.A1(new_n479), .A2(new_n221), .ZN(new_n480));
  AND3_X1   g0280(.A1(new_n474), .A2(new_n477), .A3(new_n480), .ZN(new_n481));
  INV_X1    g0281(.A(KEYINPUT81), .ZN(new_n482));
  INV_X1    g0282(.A(G45), .ZN(new_n483));
  OR3_X1    g0283(.A1(new_n483), .A2(G1), .A3(G274), .ZN(new_n484));
  OAI21_X1  g0284(.A(new_n222), .B1(new_n483), .B2(G1), .ZN(new_n485));
  NAND4_X1  g0285(.A1(new_n297), .A2(new_n484), .A3(new_n299), .A4(new_n485), .ZN(new_n486));
  INV_X1    g0286(.A(new_n486), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n226), .A2(new_n279), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n220), .A2(G1698), .ZN(new_n489));
  OAI211_X1 g0289(.A(new_n488), .B(new_n489), .C1(new_n287), .C2(new_n288), .ZN(new_n490));
  NAND2_X1  g0290(.A1(G33), .A2(G116), .ZN(new_n491));
  AOI21_X1  g0291(.A(new_n292), .B1(new_n490), .B2(new_n491), .ZN(new_n492));
  OAI21_X1  g0292(.A(new_n482), .B1(new_n487), .B2(new_n492), .ZN(new_n493));
  AND2_X1   g0293(.A1(new_n490), .A2(new_n491), .ZN(new_n494));
  OAI211_X1 g0294(.A(KEYINPUT81), .B(new_n486), .C1(new_n494), .C2(new_n292), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n493), .A2(new_n495), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n496), .A2(G200), .ZN(new_n497));
  NAND3_X1  g0297(.A1(new_n493), .A2(new_n495), .A3(G190), .ZN(new_n498));
  AND2_X1   g0298(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  AOI21_X1  g0299(.A(G169), .B1(new_n493), .B2(new_n495), .ZN(new_n500));
  AND2_X1   g0300(.A1(new_n493), .A2(new_n495), .ZN(new_n501));
  AOI21_X1  g0301(.A(new_n500), .B1(new_n309), .B2(new_n501), .ZN(new_n502));
  NOR2_X1   g0302(.A1(new_n479), .A2(new_n438), .ZN(new_n503));
  XNOR2_X1  g0303(.A(new_n503), .B(KEYINPUT84), .ZN(new_n504));
  NAND3_X1  g0304(.A1(new_n474), .A2(new_n477), .A3(new_n504), .ZN(new_n505));
  AOI22_X1  g0305(.A1(new_n481), .A2(new_n499), .B1(new_n502), .B2(new_n505), .ZN(new_n506));
  INV_X1    g0306(.A(G41), .ZN(new_n507));
  OAI211_X1 g0307(.A(new_n207), .B(G45), .C1(new_n507), .C2(KEYINPUT5), .ZN(new_n508));
  AND2_X1   g0308(.A1(new_n507), .A2(KEYINPUT5), .ZN(new_n509));
  OR2_X1    g0309(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  NAND4_X1  g0310(.A1(new_n510), .A2(new_n297), .A3(G257), .A4(new_n299), .ZN(new_n511));
  NOR2_X1   g0311(.A1(new_n508), .A2(new_n509), .ZN(new_n512));
  NAND4_X1  g0312(.A1(new_n512), .A2(G274), .A3(new_n297), .A4(new_n299), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n511), .A2(new_n513), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n279), .A2(G244), .ZN(new_n515));
  AOI21_X1  g0315(.A(new_n515), .B1(new_n277), .B2(new_n278), .ZN(new_n516));
  AOI22_X1  g0316(.A1(new_n516), .A2(KEYINPUT4), .B1(G33), .B2(G283), .ZN(new_n517));
  INV_X1    g0317(.A(KEYINPUT78), .ZN(new_n518));
  OAI21_X1  g0318(.A(new_n518), .B1(new_n516), .B2(KEYINPUT4), .ZN(new_n519));
  NAND3_X1  g0319(.A1(new_n335), .A2(G250), .A3(G1698), .ZN(new_n520));
  OAI211_X1 g0320(.A(G244), .B(new_n279), .C1(new_n287), .C2(new_n288), .ZN(new_n521));
  INV_X1    g0321(.A(KEYINPUT4), .ZN(new_n522));
  NAND3_X1  g0322(.A1(new_n521), .A2(KEYINPUT78), .A3(new_n522), .ZN(new_n523));
  NAND4_X1  g0323(.A1(new_n517), .A2(new_n519), .A3(new_n520), .A4(new_n523), .ZN(new_n524));
  AOI21_X1  g0324(.A(new_n514), .B1(new_n524), .B2(new_n293), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n525), .A2(G190), .ZN(new_n526));
  OAI21_X1  g0326(.A(G107), .B1(new_n400), .B2(new_n401), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n254), .A2(G77), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n528), .A2(KEYINPUT77), .ZN(new_n529));
  INV_X1    g0329(.A(KEYINPUT77), .ZN(new_n530));
  NAND3_X1  g0330(.A1(new_n254), .A2(new_n530), .A3(G77), .ZN(new_n531));
  NAND3_X1  g0331(.A1(new_n463), .A2(KEYINPUT6), .A3(G97), .ZN(new_n532));
  XOR2_X1   g0332(.A(G97), .B(G107), .Z(new_n533));
  OAI21_X1  g0333(.A(new_n532), .B1(new_n533), .B2(KEYINPUT6), .ZN(new_n534));
  AOI22_X1  g0334(.A1(new_n529), .A2(new_n531), .B1(new_n534), .B2(G20), .ZN(new_n535));
  AOI21_X1  g0335(.A(new_n249), .B1(new_n527), .B2(new_n535), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n267), .A2(new_n458), .ZN(new_n537));
  OAI21_X1  g0337(.A(new_n537), .B1(new_n479), .B2(new_n458), .ZN(new_n538));
  NOR2_X1   g0338(.A1(new_n536), .A2(new_n538), .ZN(new_n539));
  OAI21_X1  g0339(.A(G200), .B1(new_n525), .B2(KEYINPUT79), .ZN(new_n540));
  INV_X1    g0340(.A(KEYINPUT79), .ZN(new_n541));
  AOI211_X1 g0341(.A(new_n541), .B(new_n514), .C1(new_n293), .C2(new_n524), .ZN(new_n542));
  OAI211_X1 g0342(.A(new_n526), .B(new_n539), .C1(new_n540), .C2(new_n542), .ZN(new_n543));
  INV_X1    g0343(.A(new_n536), .ZN(new_n544));
  INV_X1    g0344(.A(new_n538), .ZN(new_n545));
  NAND3_X1  g0345(.A1(new_n544), .A2(KEYINPUT80), .A3(new_n545), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n524), .A2(new_n293), .ZN(new_n547));
  NAND4_X1  g0347(.A1(new_n547), .A2(G179), .A3(new_n513), .A4(new_n511), .ZN(new_n548));
  OAI21_X1  g0348(.A(new_n548), .B1(new_n366), .B2(new_n525), .ZN(new_n549));
  INV_X1    g0349(.A(KEYINPUT80), .ZN(new_n550));
  OAI21_X1  g0350(.A(new_n550), .B1(new_n536), .B2(new_n538), .ZN(new_n551));
  NAND3_X1  g0351(.A1(new_n546), .A2(new_n549), .A3(new_n551), .ZN(new_n552));
  NAND4_X1  g0352(.A1(new_n506), .A2(KEYINPUT85), .A3(new_n543), .A4(new_n552), .ZN(new_n553));
  INV_X1    g0353(.A(KEYINPUT85), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n552), .A2(new_n543), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n502), .A2(new_n505), .ZN(new_n556));
  AOI21_X1  g0356(.A(new_n249), .B1(new_n468), .B2(new_n469), .ZN(new_n557));
  AOI21_X1  g0357(.A(new_n476), .B1(new_n557), .B2(new_n473), .ZN(new_n558));
  NAND4_X1  g0358(.A1(new_n558), .A2(new_n480), .A3(new_n497), .A4(new_n498), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n556), .A2(new_n559), .ZN(new_n560));
  OAI21_X1  g0360(.A(new_n554), .B1(new_n555), .B2(new_n560), .ZN(new_n561));
  NAND3_X1  g0361(.A1(new_n333), .A2(G270), .A3(new_n510), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n279), .A2(G257), .ZN(new_n563));
  NAND2_X1  g0363(.A1(G264), .A2(G1698), .ZN(new_n564));
  NAND3_X1  g0364(.A1(new_n335), .A2(new_n563), .A3(new_n564), .ZN(new_n565));
  INV_X1    g0365(.A(G303), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n289), .A2(new_n566), .ZN(new_n567));
  NAND3_X1  g0367(.A1(new_n565), .A2(new_n293), .A3(new_n567), .ZN(new_n568));
  NAND3_X1  g0368(.A1(new_n562), .A2(new_n513), .A3(new_n568), .ZN(new_n569));
  INV_X1    g0369(.A(G116), .ZN(new_n570));
  OR2_X1    g0370(.A1(new_n479), .A2(new_n570), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n267), .A2(new_n570), .ZN(new_n572));
  AOI22_X1  g0372(.A1(new_n247), .A2(new_n214), .B1(G20), .B2(new_n570), .ZN(new_n573));
  NAND2_X1  g0373(.A1(G33), .A2(G283), .ZN(new_n574));
  OAI211_X1 g0374(.A(new_n574), .B(new_n208), .C1(G33), .C2(new_n458), .ZN(new_n575));
  AND3_X1   g0375(.A1(new_n573), .A2(KEYINPUT20), .A3(new_n575), .ZN(new_n576));
  AOI21_X1  g0376(.A(KEYINPUT20), .B1(new_n573), .B2(new_n575), .ZN(new_n577));
  OAI211_X1 g0377(.A(new_n571), .B(new_n572), .C1(new_n576), .C2(new_n577), .ZN(new_n578));
  NAND3_X1  g0378(.A1(new_n569), .A2(new_n578), .A3(G169), .ZN(new_n579));
  INV_X1    g0379(.A(KEYINPUT21), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  NOR2_X1   g0381(.A1(new_n569), .A2(new_n309), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n582), .A2(new_n578), .ZN(new_n583));
  NAND4_X1  g0383(.A1(new_n569), .A2(new_n578), .A3(KEYINPUT21), .A4(G169), .ZN(new_n584));
  AND3_X1   g0384(.A1(new_n581), .A2(new_n583), .A3(new_n584), .ZN(new_n585));
  AOI21_X1  g0385(.A(new_n578), .B1(new_n569), .B2(G200), .ZN(new_n586));
  OAI21_X1  g0386(.A(new_n586), .B1(new_n342), .B2(new_n569), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n585), .A2(new_n587), .ZN(new_n588));
  NOR2_X1   g0388(.A1(new_n491), .A2(G20), .ZN(new_n589));
  INV_X1    g0389(.A(KEYINPUT23), .ZN(new_n590));
  OAI21_X1  g0390(.A(new_n590), .B1(new_n208), .B2(G107), .ZN(new_n591));
  NAND3_X1  g0391(.A1(new_n463), .A2(KEYINPUT23), .A3(G20), .ZN(new_n592));
  AOI21_X1  g0392(.A(new_n589), .B1(new_n591), .B2(new_n592), .ZN(new_n593));
  OAI211_X1 g0393(.A(new_n208), .B(G87), .C1(new_n287), .C2(new_n288), .ZN(new_n594));
  INV_X1    g0394(.A(KEYINPUT22), .ZN(new_n595));
  NOR2_X1   g0395(.A1(new_n595), .A2(KEYINPUT86), .ZN(new_n596));
  AND2_X1   g0396(.A1(new_n594), .A2(new_n596), .ZN(new_n597));
  NOR2_X1   g0397(.A1(new_n594), .A2(new_n596), .ZN(new_n598));
  OAI21_X1  g0398(.A(new_n593), .B1(new_n597), .B2(new_n598), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n599), .A2(KEYINPUT24), .ZN(new_n600));
  INV_X1    g0400(.A(KEYINPUT24), .ZN(new_n601));
  OAI211_X1 g0401(.A(new_n601), .B(new_n593), .C1(new_n597), .C2(new_n598), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n600), .A2(new_n602), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n603), .A2(new_n248), .ZN(new_n604));
  NAND3_X1  g0404(.A1(new_n267), .A2(KEYINPUT25), .A3(new_n463), .ZN(new_n605));
  INV_X1    g0405(.A(new_n605), .ZN(new_n606));
  AOI21_X1  g0406(.A(KEYINPUT25), .B1(new_n267), .B2(new_n463), .ZN(new_n607));
  OAI22_X1  g0407(.A1(new_n606), .A2(new_n607), .B1(new_n463), .B2(new_n479), .ZN(new_n608));
  INV_X1    g0408(.A(new_n608), .ZN(new_n609));
  OAI211_X1 g0409(.A(G250), .B(new_n279), .C1(new_n287), .C2(new_n288), .ZN(new_n610));
  OAI211_X1 g0410(.A(G257), .B(G1698), .C1(new_n287), .C2(new_n288), .ZN(new_n611));
  INV_X1    g0411(.A(G294), .ZN(new_n612));
  OAI211_X1 g0412(.A(new_n610), .B(new_n611), .C1(new_n251), .C2(new_n612), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n613), .A2(new_n293), .ZN(new_n614));
  NAND3_X1  g0414(.A1(new_n333), .A2(G264), .A3(new_n510), .ZN(new_n615));
  NAND3_X1  g0415(.A1(new_n614), .A2(new_n615), .A3(new_n513), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n616), .A2(G200), .ZN(new_n617));
  AND2_X1   g0417(.A1(new_n614), .A2(new_n615), .ZN(new_n618));
  NAND3_X1  g0418(.A1(new_n618), .A2(G190), .A3(new_n513), .ZN(new_n619));
  NAND4_X1  g0419(.A1(new_n604), .A2(new_n609), .A3(new_n617), .A4(new_n619), .ZN(new_n620));
  NAND4_X1  g0420(.A1(new_n614), .A2(new_n615), .A3(new_n309), .A4(new_n513), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n616), .A2(new_n366), .ZN(new_n622));
  AOI21_X1  g0422(.A(new_n249), .B1(new_n600), .B2(new_n602), .ZN(new_n623));
  OAI211_X1 g0423(.A(new_n621), .B(new_n622), .C1(new_n623), .C2(new_n608), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n620), .A2(new_n624), .ZN(new_n625));
  NOR2_X1   g0425(.A1(new_n588), .A2(new_n625), .ZN(new_n626));
  AND4_X1   g0426(.A1(new_n456), .A2(new_n553), .A3(new_n561), .A4(new_n626), .ZN(G372));
  NAND2_X1  g0427(.A1(new_n414), .A2(new_n430), .ZN(new_n628));
  INV_X1    g0428(.A(new_n326), .ZN(new_n629));
  AND2_X1   g0429(.A1(new_n313), .A2(new_n319), .ZN(new_n630));
  AOI21_X1  g0430(.A(new_n325), .B1(new_n630), .B2(new_n324), .ZN(new_n631));
  OAI21_X1  g0431(.A(new_n272), .B1(new_n629), .B2(new_n631), .ZN(new_n632));
  INV_X1    g0432(.A(new_n453), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n330), .A2(new_n633), .ZN(new_n634));
  AOI21_X1  g0434(.A(new_n628), .B1(new_n632), .B2(new_n634), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n429), .A2(new_n434), .ZN(new_n636));
  OAI21_X1  g0436(.A(new_n364), .B1(new_n635), .B2(new_n636), .ZN(new_n637));
  AND2_X1   g0437(.A1(new_n637), .A2(new_n368), .ZN(new_n638));
  INV_X1    g0438(.A(new_n456), .ZN(new_n639));
  INV_X1    g0439(.A(KEYINPUT87), .ZN(new_n640));
  NAND3_X1  g0440(.A1(new_n585), .A2(new_n624), .A3(new_n640), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n622), .A2(new_n621), .ZN(new_n642));
  AOI21_X1  g0442(.A(new_n642), .B1(new_n604), .B2(new_n609), .ZN(new_n643));
  NAND3_X1  g0443(.A1(new_n581), .A2(new_n583), .A3(new_n584), .ZN(new_n644));
  OAI21_X1  g0444(.A(KEYINPUT87), .B1(new_n643), .B2(new_n644), .ZN(new_n645));
  OAI21_X1  g0445(.A(new_n486), .B1(new_n494), .B2(new_n292), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n646), .A2(G200), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n498), .A2(new_n647), .ZN(new_n648));
  INV_X1    g0448(.A(new_n648), .ZN(new_n649));
  NAND3_X1  g0449(.A1(new_n493), .A2(new_n495), .A3(new_n309), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n646), .A2(new_n366), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  INV_X1    g0452(.A(new_n652), .ZN(new_n653));
  AOI22_X1  g0453(.A1(new_n481), .A2(new_n649), .B1(new_n653), .B2(new_n505), .ZN(new_n654));
  NAND3_X1  g0454(.A1(new_n641), .A2(new_n645), .A3(new_n654), .ZN(new_n655));
  NAND3_X1  g0455(.A1(new_n552), .A2(new_n543), .A3(new_n620), .ZN(new_n656));
  NOR2_X1   g0456(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  OAI21_X1  g0457(.A(KEYINPUT26), .B1(new_n560), .B2(new_n552), .ZN(new_n658));
  INV_X1    g0458(.A(KEYINPUT26), .ZN(new_n659));
  INV_X1    g0459(.A(new_n539), .ZN(new_n660));
  NAND4_X1  g0460(.A1(new_n654), .A2(new_n659), .A3(new_n660), .A4(new_n549), .ZN(new_n661));
  AND3_X1   g0461(.A1(new_n474), .A2(new_n477), .A3(new_n504), .ZN(new_n662));
  NOR3_X1   g0462(.A1(new_n662), .A2(KEYINPUT88), .A3(new_n652), .ZN(new_n663));
  INV_X1    g0463(.A(KEYINPUT88), .ZN(new_n664));
  AOI21_X1  g0464(.A(new_n664), .B1(new_n653), .B2(new_n505), .ZN(new_n665));
  NOR2_X1   g0465(.A1(new_n663), .A2(new_n665), .ZN(new_n666));
  NAND3_X1  g0466(.A1(new_n658), .A2(new_n661), .A3(new_n666), .ZN(new_n667));
  NOR2_X1   g0467(.A1(new_n657), .A2(new_n667), .ZN(new_n668));
  OAI21_X1  g0468(.A(new_n638), .B1(new_n639), .B2(new_n668), .ZN(G369));
  NAND3_X1  g0469(.A1(new_n207), .A2(new_n208), .A3(G13), .ZN(new_n670));
  OR2_X1    g0470(.A1(new_n670), .A2(KEYINPUT27), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n670), .A2(KEYINPUT27), .ZN(new_n672));
  NAND3_X1  g0472(.A1(new_n671), .A2(G213), .A3(new_n672), .ZN(new_n673));
  INV_X1    g0473(.A(G343), .ZN(new_n674));
  NOR2_X1   g0474(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  AND2_X1   g0475(.A1(new_n578), .A2(new_n675), .ZN(new_n676));
  OR2_X1    g0476(.A1(new_n588), .A2(new_n676), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n644), .A2(new_n676), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  INV_X1    g0479(.A(new_n679), .ZN(new_n680));
  INV_X1    g0480(.A(G330), .ZN(new_n681));
  NOR2_X1   g0481(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  OAI21_X1  g0482(.A(new_n675), .B1(new_n623), .B2(new_n608), .ZN(new_n683));
  NAND3_X1  g0483(.A1(new_n620), .A2(new_n624), .A3(new_n683), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n643), .A2(new_n675), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n682), .A2(new_n686), .ZN(new_n687));
  INV_X1    g0487(.A(new_n675), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n644), .A2(new_n688), .ZN(new_n689));
  NOR2_X1   g0489(.A1(new_n625), .A2(new_n689), .ZN(new_n690));
  AOI21_X1  g0490(.A(new_n690), .B1(new_n643), .B2(new_n688), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n687), .A2(new_n691), .ZN(G399));
  OR2_X1    g0492(.A1(new_n464), .A2(G116), .ZN(new_n693));
  XOR2_X1   g0493(.A(new_n693), .B(KEYINPUT89), .Z(new_n694));
  NAND2_X1  g0494(.A1(new_n211), .A2(new_n507), .ZN(new_n695));
  INV_X1    g0495(.A(new_n695), .ZN(new_n696));
  NOR3_X1   g0496(.A1(new_n694), .A2(new_n207), .A3(new_n696), .ZN(new_n697));
  INV_X1    g0497(.A(new_n217), .ZN(new_n698));
  AOI21_X1  g0498(.A(new_n697), .B1(new_n698), .B2(new_n696), .ZN(new_n699));
  XOR2_X1   g0499(.A(new_n699), .B(KEYINPUT28), .Z(new_n700));
  NAND4_X1  g0500(.A1(new_n561), .A2(new_n553), .A3(new_n626), .A4(new_n688), .ZN(new_n701));
  INV_X1    g0501(.A(KEYINPUT30), .ZN(new_n702));
  NAND3_X1  g0502(.A1(new_n501), .A2(new_n582), .A3(new_n618), .ZN(new_n703));
  INV_X1    g0503(.A(new_n525), .ZN(new_n704));
  OAI21_X1  g0504(.A(new_n702), .B1(new_n703), .B2(new_n704), .ZN(new_n705));
  AND3_X1   g0505(.A1(new_n618), .A2(new_n493), .A3(new_n495), .ZN(new_n706));
  NAND4_X1  g0506(.A1(new_n706), .A2(KEYINPUT30), .A3(new_n525), .A4(new_n582), .ZN(new_n707));
  AND2_X1   g0507(.A1(new_n646), .A2(new_n309), .ZN(new_n708));
  NAND4_X1  g0508(.A1(new_n704), .A2(new_n616), .A3(new_n569), .A4(new_n708), .ZN(new_n709));
  NAND3_X1  g0509(.A1(new_n705), .A2(new_n707), .A3(new_n709), .ZN(new_n710));
  AND3_X1   g0510(.A1(new_n710), .A2(KEYINPUT31), .A3(new_n675), .ZN(new_n711));
  AOI21_X1  g0511(.A(KEYINPUT31), .B1(new_n710), .B2(new_n675), .ZN(new_n712));
  NOR2_X1   g0512(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  AOI21_X1  g0513(.A(new_n681), .B1(new_n701), .B2(new_n713), .ZN(new_n714));
  INV_X1    g0514(.A(KEYINPUT29), .ZN(new_n715));
  OAI21_X1  g0515(.A(new_n715), .B1(new_n668), .B2(new_n675), .ZN(new_n716));
  INV_X1    g0516(.A(new_n552), .ZN(new_n717));
  NAND3_X1  g0517(.A1(new_n717), .A2(new_n506), .A3(new_n659), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n558), .A2(new_n480), .ZN(new_n719));
  OAI22_X1  g0519(.A1(new_n662), .A2(new_n652), .B1(new_n719), .B2(new_n648), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n660), .A2(new_n549), .ZN(new_n721));
  OAI21_X1  g0521(.A(KEYINPUT26), .B1(new_n720), .B2(new_n721), .ZN(new_n722));
  NAND3_X1  g0522(.A1(new_n718), .A2(new_n722), .A3(new_n666), .ZN(new_n723));
  OAI21_X1  g0523(.A(new_n654), .B1(new_n643), .B2(new_n644), .ZN(new_n724));
  NOR2_X1   g0524(.A1(new_n724), .A2(new_n656), .ZN(new_n725));
  OAI211_X1 g0525(.A(KEYINPUT29), .B(new_n688), .C1(new_n723), .C2(new_n725), .ZN(new_n726));
  AOI21_X1  g0526(.A(new_n714), .B1(new_n716), .B2(new_n726), .ZN(new_n727));
  OAI21_X1  g0527(.A(new_n700), .B1(new_n727), .B2(G1), .ZN(G364));
  INV_X1    g0528(.A(G13), .ZN(new_n729));
  NOR2_X1   g0529(.A1(new_n729), .A2(G20), .ZN(new_n730));
  AOI21_X1  g0530(.A(new_n207), .B1(new_n730), .B2(G45), .ZN(new_n731));
  INV_X1    g0531(.A(new_n731), .ZN(new_n732));
  NOR2_X1   g0532(.A1(new_n696), .A2(new_n732), .ZN(new_n733));
  NOR2_X1   g0533(.A1(new_n682), .A2(new_n733), .ZN(new_n734));
  OAI21_X1  g0534(.A(new_n734), .B1(G330), .B2(new_n679), .ZN(new_n735));
  NAND2_X1  g0535(.A1(new_n211), .A2(new_n335), .ZN(new_n736));
  INV_X1    g0536(.A(G355), .ZN(new_n737));
  OAI22_X1  g0537(.A1(new_n736), .A2(new_n737), .B1(G116), .B2(new_n211), .ZN(new_n738));
  NAND2_X1  g0538(.A1(new_n242), .A2(G45), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n211), .A2(new_n289), .ZN(new_n740));
  AOI21_X1  g0540(.A(new_n740), .B1(new_n483), .B2(new_n698), .ZN(new_n741));
  AOI21_X1  g0541(.A(new_n738), .B1(new_n739), .B2(new_n741), .ZN(new_n742));
  AOI21_X1  g0542(.A(new_n214), .B1(G20), .B2(new_n366), .ZN(new_n743));
  OR2_X1    g0543(.A1(new_n743), .A2(KEYINPUT90), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n743), .A2(KEYINPUT90), .ZN(new_n745));
  NAND2_X1  g0545(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  NOR2_X1   g0546(.A1(G13), .A2(G33), .ZN(new_n747));
  INV_X1    g0547(.A(new_n747), .ZN(new_n748));
  NOR2_X1   g0548(.A1(new_n748), .A2(G20), .ZN(new_n749));
  NOR2_X1   g0549(.A1(new_n746), .A2(new_n749), .ZN(new_n750));
  INV_X1    g0550(.A(new_n750), .ZN(new_n751));
  OAI21_X1  g0551(.A(new_n733), .B1(new_n742), .B2(new_n751), .ZN(new_n752));
  NOR2_X1   g0552(.A1(new_n342), .A2(new_n378), .ZN(new_n753));
  NOR2_X1   g0553(.A1(new_n208), .A2(new_n309), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  INV_X1    g0555(.A(new_n755), .ZN(new_n756));
  AOI21_X1  g0556(.A(new_n335), .B1(new_n756), .B2(G326), .ZN(new_n757));
  INV_X1    g0557(.A(G311), .ZN(new_n758));
  NOR2_X1   g0558(.A1(G190), .A2(G200), .ZN(new_n759));
  NAND2_X1  g0559(.A1(new_n754), .A2(new_n759), .ZN(new_n760));
  INV_X1    g0560(.A(G322), .ZN(new_n761));
  NAND3_X1  g0561(.A1(new_n754), .A2(G190), .A3(new_n378), .ZN(new_n762));
  OAI221_X1 g0562(.A(new_n757), .B1(new_n758), .B2(new_n760), .C1(new_n761), .C2(new_n762), .ZN(new_n763));
  NOR2_X1   g0563(.A1(new_n208), .A2(G190), .ZN(new_n764));
  NAND3_X1  g0564(.A1(new_n764), .A2(new_n309), .A3(G200), .ZN(new_n765));
  INV_X1    g0565(.A(G283), .ZN(new_n766));
  INV_X1    g0566(.A(G329), .ZN(new_n767));
  NAND3_X1  g0567(.A1(new_n759), .A2(G20), .A3(new_n309), .ZN(new_n768));
  OAI22_X1  g0568(.A1(new_n765), .A2(new_n766), .B1(new_n767), .B2(new_n768), .ZN(new_n769));
  NAND3_X1  g0569(.A1(new_n764), .A2(G179), .A3(G200), .ZN(new_n770));
  XOR2_X1   g0570(.A(KEYINPUT33), .B(G317), .Z(new_n771));
  NAND3_X1  g0571(.A1(new_n753), .A2(G20), .A3(new_n309), .ZN(new_n772));
  OAI22_X1  g0572(.A1(new_n770), .A2(new_n771), .B1(new_n772), .B2(new_n566), .ZN(new_n773));
  NOR3_X1   g0573(.A1(new_n342), .A2(G179), .A3(G200), .ZN(new_n774));
  NOR2_X1   g0574(.A1(new_n774), .A2(new_n208), .ZN(new_n775));
  NOR2_X1   g0575(.A1(new_n775), .A2(new_n612), .ZN(new_n776));
  NOR4_X1   g0576(.A1(new_n763), .A2(new_n769), .A3(new_n773), .A4(new_n776), .ZN(new_n777));
  XNOR2_X1  g0577(.A(new_n777), .B(KEYINPUT92), .ZN(new_n778));
  AOI21_X1  g0578(.A(new_n289), .B1(new_n756), .B2(G50), .ZN(new_n779));
  INV_X1    g0579(.A(new_n775), .ZN(new_n780));
  NAND2_X1  g0580(.A1(new_n780), .A2(G97), .ZN(new_n781));
  INV_X1    g0581(.A(G159), .ZN(new_n782));
  OAI21_X1  g0582(.A(KEYINPUT32), .B1(new_n768), .B2(new_n782), .ZN(new_n783));
  OR3_X1    g0583(.A1(new_n768), .A2(KEYINPUT32), .A3(new_n782), .ZN(new_n784));
  NAND4_X1  g0584(.A1(new_n779), .A2(new_n781), .A3(new_n783), .A4(new_n784), .ZN(new_n785));
  INV_X1    g0585(.A(new_n772), .ZN(new_n786));
  INV_X1    g0586(.A(new_n765), .ZN(new_n787));
  AOI22_X1  g0587(.A1(G87), .A2(new_n786), .B1(new_n787), .B2(G107), .ZN(new_n788));
  OAI21_X1  g0588(.A(new_n788), .B1(new_n203), .B2(new_n770), .ZN(new_n789));
  INV_X1    g0589(.A(new_n762), .ZN(new_n790));
  INV_X1    g0590(.A(new_n760), .ZN(new_n791));
  AOI22_X1  g0591(.A1(new_n790), .A2(G58), .B1(new_n791), .B2(G77), .ZN(new_n792));
  AOI21_X1  g0592(.A(new_n789), .B1(KEYINPUT91), .B2(new_n792), .ZN(new_n793));
  OAI21_X1  g0593(.A(new_n793), .B1(KEYINPUT91), .B2(new_n792), .ZN(new_n794));
  OAI21_X1  g0594(.A(new_n778), .B1(new_n785), .B2(new_n794), .ZN(new_n795));
  OR2_X1    g0595(.A1(new_n795), .A2(KEYINPUT93), .ZN(new_n796));
  INV_X1    g0596(.A(new_n746), .ZN(new_n797));
  AOI21_X1  g0597(.A(new_n797), .B1(new_n795), .B2(KEYINPUT93), .ZN(new_n798));
  AOI21_X1  g0598(.A(new_n752), .B1(new_n796), .B2(new_n798), .ZN(new_n799));
  XNOR2_X1  g0599(.A(new_n749), .B(KEYINPUT94), .ZN(new_n800));
  OAI21_X1  g0600(.A(new_n799), .B1(new_n679), .B2(new_n800), .ZN(new_n801));
  AND2_X1   g0601(.A1(new_n735), .A2(new_n801), .ZN(new_n802));
  INV_X1    g0602(.A(new_n802), .ZN(G396));
  NOR2_X1   g0603(.A1(new_n453), .A2(new_n688), .ZN(new_n804));
  INV_X1    g0604(.A(KEYINPUT97), .ZN(new_n805));
  XNOR2_X1  g0605(.A(new_n804), .B(new_n805), .ZN(new_n806));
  NAND2_X1  g0606(.A1(new_n633), .A2(KEYINPUT96), .ZN(new_n807));
  INV_X1    g0607(.A(KEYINPUT96), .ZN(new_n808));
  NAND2_X1  g0608(.A1(new_n453), .A2(new_n808), .ZN(new_n809));
  NAND2_X1  g0609(.A1(new_n442), .A2(new_n675), .ZN(new_n810));
  NAND4_X1  g0610(.A1(new_n807), .A2(new_n450), .A3(new_n809), .A4(new_n810), .ZN(new_n811));
  NAND2_X1  g0611(.A1(new_n806), .A2(new_n811), .ZN(new_n812));
  INV_X1    g0612(.A(new_n812), .ZN(new_n813));
  OAI21_X1  g0613(.A(new_n813), .B1(new_n668), .B2(new_n675), .ZN(new_n814));
  OAI211_X1 g0614(.A(new_n688), .B(new_n812), .C1(new_n657), .C2(new_n667), .ZN(new_n815));
  AOI21_X1  g0615(.A(new_n714), .B1(new_n814), .B2(new_n815), .ZN(new_n816));
  NOR2_X1   g0616(.A1(new_n816), .A2(new_n733), .ZN(new_n817));
  NAND3_X1  g0617(.A1(new_n814), .A2(new_n714), .A3(new_n815), .ZN(new_n818));
  NAND2_X1  g0618(.A1(new_n817), .A2(new_n818), .ZN(new_n819));
  NOR2_X1   g0619(.A1(new_n746), .A2(new_n747), .ZN(new_n820));
  INV_X1    g0620(.A(new_n820), .ZN(new_n821));
  OAI21_X1  g0621(.A(new_n733), .B1(new_n821), .B2(G77), .ZN(new_n822));
  OAI22_X1  g0622(.A1(new_n765), .A2(new_n221), .B1(new_n758), .B2(new_n768), .ZN(new_n823));
  AOI211_X1 g0623(.A(new_n335), .B(new_n823), .C1(G107), .C2(new_n786), .ZN(new_n824));
  AOI22_X1  g0624(.A1(new_n790), .A2(G294), .B1(new_n791), .B2(G116), .ZN(new_n825));
  INV_X1    g0625(.A(new_n770), .ZN(new_n826));
  AOI22_X1  g0626(.A1(G303), .A2(new_n756), .B1(new_n826), .B2(G283), .ZN(new_n827));
  NAND4_X1  g0627(.A1(new_n824), .A2(new_n781), .A3(new_n825), .A4(new_n827), .ZN(new_n828));
  AOI22_X1  g0628(.A1(G137), .A2(new_n756), .B1(new_n791), .B2(G159), .ZN(new_n829));
  INV_X1    g0629(.A(G150), .ZN(new_n830));
  XNOR2_X1  g0630(.A(KEYINPUT95), .B(G143), .ZN(new_n831));
  OAI221_X1 g0631(.A(new_n829), .B1(new_n830), .B2(new_n770), .C1(new_n762), .C2(new_n831), .ZN(new_n832));
  XOR2_X1   g0632(.A(new_n832), .B(KEYINPUT34), .Z(new_n833));
  INV_X1    g0633(.A(new_n768), .ZN(new_n834));
  AOI22_X1  g0634(.A1(new_n786), .A2(G50), .B1(G132), .B2(new_n834), .ZN(new_n835));
  AOI21_X1  g0635(.A(new_n289), .B1(new_n787), .B2(G68), .ZN(new_n836));
  OAI211_X1 g0636(.A(new_n835), .B(new_n836), .C1(new_n202), .C2(new_n775), .ZN(new_n837));
  OAI21_X1  g0637(.A(new_n828), .B1(new_n833), .B2(new_n837), .ZN(new_n838));
  AOI21_X1  g0638(.A(new_n822), .B1(new_n838), .B2(new_n746), .ZN(new_n839));
  OAI21_X1  g0639(.A(new_n839), .B1(new_n812), .B2(new_n748), .ZN(new_n840));
  NAND2_X1  g0640(.A1(new_n819), .A2(new_n840), .ZN(G384));
  OAI21_X1  g0641(.A(G77), .B1(new_n202), .B2(new_n203), .ZN(new_n842));
  OAI22_X1  g0642(.A1(new_n842), .A2(new_n217), .B1(G50), .B2(new_n203), .ZN(new_n843));
  NAND3_X1  g0643(.A1(new_n843), .A2(G1), .A3(new_n729), .ZN(new_n844));
  XOR2_X1   g0644(.A(new_n844), .B(KEYINPUT98), .Z(new_n845));
  AOI211_X1 g0645(.A(new_n570), .B(new_n216), .C1(new_n534), .C2(KEYINPUT35), .ZN(new_n846));
  OAI21_X1  g0646(.A(new_n846), .B1(KEYINPUT35), .B2(new_n534), .ZN(new_n847));
  INV_X1    g0647(.A(KEYINPUT36), .ZN(new_n848));
  OAI21_X1  g0648(.A(new_n845), .B1(new_n847), .B2(new_n848), .ZN(new_n849));
  AOI21_X1  g0649(.A(new_n849), .B1(new_n848), .B2(new_n847), .ZN(new_n850));
  NAND2_X1  g0650(.A1(new_n701), .A2(new_n713), .ZN(new_n851));
  NOR2_X1   g0651(.A1(new_n273), .A2(new_n688), .ZN(new_n852));
  NOR3_X1   g0652(.A1(new_n327), .A2(new_n331), .A3(new_n852), .ZN(new_n853));
  INV_X1    g0653(.A(new_n852), .ZN(new_n854));
  AOI21_X1  g0654(.A(new_n854), .B1(new_n321), .B2(new_n326), .ZN(new_n855));
  OAI211_X1 g0655(.A(new_n851), .B(new_n812), .C1(new_n853), .C2(new_n855), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n856), .A2(KEYINPUT102), .ZN(new_n857));
  NAND3_X1  g0657(.A1(new_n632), .A2(new_n330), .A3(new_n854), .ZN(new_n858));
  OAI21_X1  g0658(.A(new_n852), .B1(new_n629), .B2(new_n631), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  INV_X1    g0660(.A(KEYINPUT102), .ZN(new_n861));
  NAND4_X1  g0661(.A1(new_n860), .A2(new_n861), .A3(new_n851), .A4(new_n812), .ZN(new_n862));
  INV_X1    g0662(.A(KEYINPUT100), .ZN(new_n863));
  XOR2_X1   g0663(.A(new_n673), .B(KEYINPUT99), .Z(new_n864));
  INV_X1    g0664(.A(new_n864), .ZN(new_n865));
  OAI21_X1  g0665(.A(new_n863), .B1(new_n425), .B2(new_n865), .ZN(new_n866));
  NAND3_X1  g0666(.A1(new_n431), .A2(KEYINPUT100), .A3(new_n864), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  OAI21_X1  g0668(.A(new_n412), .B1(new_n425), .B2(new_n428), .ZN(new_n869));
  INV_X1    g0669(.A(new_n869), .ZN(new_n870));
  INV_X1    g0670(.A(KEYINPUT37), .ZN(new_n871));
  NAND3_X1  g0671(.A1(new_n868), .A2(new_n870), .A3(new_n871), .ZN(new_n872));
  OAI21_X1  g0672(.A(new_n424), .B1(KEYINPUT16), .B2(new_n423), .ZN(new_n873));
  AOI22_X1  g0673(.A1(new_n873), .A2(new_n394), .B1(new_n428), .B2(new_n673), .ZN(new_n874));
  INV_X1    g0674(.A(new_n412), .ZN(new_n875));
  OAI21_X1  g0675(.A(KEYINPUT37), .B1(new_n874), .B2(new_n875), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n872), .A2(new_n876), .ZN(new_n877));
  AOI21_X1  g0677(.A(new_n673), .B1(new_n873), .B2(new_n394), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n435), .A2(new_n878), .ZN(new_n879));
  AND3_X1   g0679(.A1(new_n877), .A2(KEYINPUT38), .A3(new_n879), .ZN(new_n880));
  AOI21_X1  g0680(.A(KEYINPUT38), .B1(new_n877), .B2(new_n879), .ZN(new_n881));
  NOR2_X1   g0681(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  INV_X1    g0682(.A(new_n882), .ZN(new_n883));
  NAND3_X1  g0683(.A1(new_n857), .A2(new_n862), .A3(new_n883), .ZN(new_n884));
  XNOR2_X1  g0684(.A(KEYINPUT101), .B(KEYINPUT40), .ZN(new_n885));
  INV_X1    g0685(.A(new_n885), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n884), .A2(new_n886), .ZN(new_n887));
  NAND3_X1  g0687(.A1(new_n877), .A2(KEYINPUT38), .A3(new_n879), .ZN(new_n888));
  AND3_X1   g0688(.A1(new_n431), .A2(KEYINPUT100), .A3(new_n864), .ZN(new_n889));
  AOI21_X1  g0689(.A(KEYINPUT100), .B1(new_n431), .B2(new_n864), .ZN(new_n890));
  NOR2_X1   g0690(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  OAI21_X1  g0691(.A(KEYINPUT37), .B1(new_n891), .B2(new_n869), .ZN(new_n892));
  AOI22_X1  g0692(.A1(new_n892), .A2(new_n872), .B1(new_n435), .B2(new_n891), .ZN(new_n893));
  OAI211_X1 g0693(.A(new_n888), .B(KEYINPUT103), .C1(new_n893), .C2(KEYINPUT38), .ZN(new_n894));
  INV_X1    g0694(.A(new_n894), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n435), .A2(new_n891), .ZN(new_n896));
  AND3_X1   g0696(.A1(new_n868), .A2(new_n871), .A3(new_n870), .ZN(new_n897));
  AOI21_X1  g0697(.A(new_n871), .B1(new_n868), .B2(new_n870), .ZN(new_n898));
  OAI21_X1  g0698(.A(new_n896), .B1(new_n897), .B2(new_n898), .ZN(new_n899));
  INV_X1    g0699(.A(KEYINPUT38), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  AOI21_X1  g0701(.A(KEYINPUT103), .B1(new_n901), .B2(new_n888), .ZN(new_n902));
  NOR2_X1   g0702(.A1(new_n895), .A2(new_n902), .ZN(new_n903));
  NAND4_X1  g0703(.A1(new_n860), .A2(KEYINPUT40), .A3(new_n851), .A4(new_n812), .ZN(new_n904));
  OAI21_X1  g0704(.A(new_n887), .B1(new_n903), .B2(new_n904), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n456), .A2(new_n851), .ZN(new_n906));
  OR2_X1    g0706(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n905), .A2(new_n906), .ZN(new_n908));
  NAND3_X1  g0708(.A1(new_n907), .A2(G330), .A3(new_n908), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n807), .A2(new_n809), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n910), .A2(new_n688), .ZN(new_n911));
  AOI22_X1  g0711(.A1(new_n815), .A2(new_n911), .B1(new_n858), .B2(new_n859), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n912), .A2(new_n883), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n636), .A2(new_n865), .ZN(new_n914));
  OAI21_X1  g0714(.A(KEYINPUT39), .B1(new_n880), .B2(new_n881), .ZN(new_n915));
  INV_X1    g0715(.A(KEYINPUT39), .ZN(new_n916));
  OAI211_X1 g0716(.A(new_n888), .B(new_n916), .C1(new_n893), .C2(KEYINPUT38), .ZN(new_n917));
  AND2_X1   g0717(.A1(new_n915), .A2(new_n917), .ZN(new_n918));
  NOR2_X1   g0718(.A1(new_n632), .A2(new_n675), .ZN(new_n919));
  INV_X1    g0719(.A(new_n919), .ZN(new_n920));
  OAI211_X1 g0720(.A(new_n913), .B(new_n914), .C1(new_n918), .C2(new_n920), .ZN(new_n921));
  NAND3_X1  g0721(.A1(new_n456), .A2(new_n716), .A3(new_n726), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n638), .A2(new_n922), .ZN(new_n923));
  XNOR2_X1  g0723(.A(new_n921), .B(new_n923), .ZN(new_n924));
  OAI22_X1  g0724(.A1(new_n909), .A2(new_n924), .B1(new_n207), .B2(new_n730), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n925), .A2(KEYINPUT104), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n909), .A2(new_n924), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  NOR2_X1   g0728(.A1(new_n925), .A2(KEYINPUT104), .ZN(new_n929));
  OAI21_X1  g0729(.A(new_n850), .B1(new_n928), .B2(new_n929), .ZN(G367));
  OAI21_X1  g0730(.A(new_n750), .B1(new_n211), .B2(new_n438), .ZN(new_n931));
  AND3_X1   g0731(.A1(new_n237), .A2(new_n211), .A3(new_n289), .ZN(new_n932));
  OAI21_X1  g0732(.A(new_n733), .B1(new_n931), .B2(new_n932), .ZN(new_n933));
  INV_X1    g0733(.A(G137), .ZN(new_n934));
  OAI22_X1  g0734(.A1(new_n772), .A2(new_n202), .B1(new_n934), .B2(new_n768), .ZN(new_n935));
  AOI211_X1 g0735(.A(new_n289), .B(new_n935), .C1(G50), .C2(new_n791), .ZN(new_n936));
  NOR2_X1   g0736(.A1(new_n765), .A2(new_n219), .ZN(new_n937));
  AOI21_X1  g0737(.A(new_n937), .B1(G150), .B2(new_n790), .ZN(new_n938));
  INV_X1    g0738(.A(new_n831), .ZN(new_n939));
  AOI22_X1  g0739(.A1(new_n756), .A2(new_n939), .B1(new_n826), .B2(G159), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n780), .A2(G68), .ZN(new_n941));
  NAND4_X1  g0741(.A1(new_n936), .A2(new_n938), .A3(new_n940), .A4(new_n941), .ZN(new_n942));
  INV_X1    g0742(.A(KEYINPUT46), .ZN(new_n943));
  NOR3_X1   g0743(.A1(new_n772), .A2(new_n943), .A3(new_n570), .ZN(new_n944));
  AOI211_X1 g0744(.A(new_n335), .B(new_n944), .C1(G311), .C2(new_n756), .ZN(new_n945));
  AOI22_X1  g0745(.A1(G303), .A2(new_n790), .B1(new_n787), .B2(G97), .ZN(new_n946));
  AOI22_X1  g0746(.A1(new_n826), .A2(G294), .B1(new_n834), .B2(G317), .ZN(new_n947));
  OAI21_X1  g0747(.A(new_n943), .B1(new_n772), .B2(new_n570), .ZN(new_n948));
  NAND4_X1  g0748(.A1(new_n945), .A2(new_n946), .A3(new_n947), .A4(new_n948), .ZN(new_n949));
  OAI22_X1  g0749(.A1(new_n775), .A2(new_n463), .B1(new_n760), .B2(new_n766), .ZN(new_n950));
  XNOR2_X1  g0750(.A(new_n950), .B(KEYINPUT107), .ZN(new_n951));
  OAI21_X1  g0751(.A(new_n942), .B1(new_n949), .B2(new_n951), .ZN(new_n952));
  INV_X1    g0752(.A(KEYINPUT47), .ZN(new_n953));
  OR2_X1    g0753(.A1(new_n952), .A2(new_n953), .ZN(new_n954));
  AOI21_X1  g0754(.A(new_n797), .B1(new_n952), .B2(new_n953), .ZN(new_n955));
  AOI21_X1  g0755(.A(new_n933), .B1(new_n954), .B2(new_n955), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n719), .A2(new_n675), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n654), .A2(new_n957), .ZN(new_n958));
  OAI21_X1  g0758(.A(new_n958), .B1(new_n666), .B2(new_n957), .ZN(new_n959));
  OAI21_X1  g0759(.A(new_n956), .B1(new_n959), .B2(new_n800), .ZN(new_n960));
  NOR2_X1   g0760(.A1(new_n539), .A2(new_n688), .ZN(new_n961));
  OAI22_X1  g0761(.A1(new_n555), .A2(new_n961), .B1(new_n721), .B2(new_n688), .ZN(new_n962));
  NOR2_X1   g0762(.A1(new_n691), .A2(new_n962), .ZN(new_n963));
  XOR2_X1   g0763(.A(new_n963), .B(KEYINPUT44), .Z(new_n964));
  NAND2_X1  g0764(.A1(new_n691), .A2(new_n962), .ZN(new_n965));
  XNOR2_X1  g0765(.A(new_n965), .B(KEYINPUT45), .ZN(new_n966));
  NOR2_X1   g0766(.A1(new_n964), .A2(new_n966), .ZN(new_n967));
  INV_X1    g0767(.A(new_n687), .ZN(new_n968));
  AND2_X1   g0768(.A1(new_n968), .A2(KEYINPUT106), .ZN(new_n969));
  XNOR2_X1  g0769(.A(new_n967), .B(new_n969), .ZN(new_n970));
  NAND3_X1  g0770(.A1(new_n684), .A2(new_n685), .A3(new_n689), .ZN(new_n971));
  OAI21_X1  g0771(.A(new_n971), .B1(new_n625), .B2(new_n689), .ZN(new_n972));
  XNOR2_X1  g0772(.A(new_n682), .B(new_n972), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n973), .A2(new_n727), .ZN(new_n974));
  INV_X1    g0774(.A(new_n974), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n970), .A2(new_n975), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n976), .A2(new_n727), .ZN(new_n977));
  XOR2_X1   g0777(.A(new_n695), .B(KEYINPUT41), .Z(new_n978));
  AOI21_X1  g0778(.A(new_n732), .B1(new_n977), .B2(new_n978), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n962), .A2(new_n690), .ZN(new_n980));
  XNOR2_X1  g0780(.A(new_n980), .B(KEYINPUT42), .ZN(new_n981));
  AND2_X1   g0781(.A1(new_n962), .A2(new_n643), .ZN(new_n982));
  OR2_X1    g0782(.A1(new_n982), .A2(new_n717), .ZN(new_n983));
  AOI21_X1  g0783(.A(new_n981), .B1(new_n688), .B2(new_n983), .ZN(new_n984));
  NOR2_X1   g0784(.A1(new_n959), .A2(KEYINPUT43), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n984), .A2(new_n985), .ZN(new_n986));
  XNOR2_X1  g0786(.A(new_n986), .B(KEYINPUT105), .ZN(new_n987));
  AND2_X1   g0787(.A1(new_n959), .A2(KEYINPUT43), .ZN(new_n988));
  OR3_X1    g0788(.A1(new_n984), .A2(new_n988), .A3(new_n985), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n987), .A2(new_n989), .ZN(new_n990));
  NAND2_X1  g0790(.A1(new_n968), .A2(new_n962), .ZN(new_n991));
  NAND2_X1  g0791(.A1(new_n990), .A2(new_n991), .ZN(new_n992));
  NAND4_X1  g0792(.A1(new_n987), .A2(new_n968), .A3(new_n962), .A4(new_n989), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n992), .A2(new_n993), .ZN(new_n994));
  OAI21_X1  g0794(.A(new_n960), .B1(new_n979), .B2(new_n994), .ZN(G387));
  NOR2_X1   g0795(.A1(new_n973), .A2(new_n727), .ZN(new_n996));
  INV_X1    g0796(.A(new_n996), .ZN(new_n997));
  NAND4_X1  g0797(.A1(new_n997), .A2(new_n507), .A3(new_n211), .A4(new_n974), .ZN(new_n998));
  NOR2_X1   g0798(.A1(new_n686), .A2(new_n800), .ZN(new_n999));
  INV_X1    g0799(.A(new_n694), .ZN(new_n1000));
  OAI22_X1  g0800(.A1(new_n1000), .A2(new_n736), .B1(G107), .B2(new_n211), .ZN(new_n1001));
  NAND2_X1  g0801(.A1(new_n234), .A2(G45), .ZN(new_n1002));
  XNOR2_X1  g0802(.A(KEYINPUT108), .B(KEYINPUT50), .ZN(new_n1003));
  NAND3_X1  g0803(.A1(new_n436), .A2(new_n1003), .A3(new_n201), .ZN(new_n1004));
  OAI211_X1 g0804(.A(new_n1004), .B(new_n483), .C1(new_n203), .C2(new_n219), .ZN(new_n1005));
  AOI21_X1  g0805(.A(new_n1003), .B1(new_n436), .B2(new_n201), .ZN(new_n1006));
  NOR2_X1   g0806(.A1(new_n1005), .A2(new_n1006), .ZN(new_n1007));
  AOI21_X1  g0807(.A(new_n740), .B1(new_n1000), .B2(new_n1007), .ZN(new_n1008));
  AOI21_X1  g0808(.A(new_n1001), .B1(new_n1002), .B2(new_n1008), .ZN(new_n1009));
  OAI21_X1  g0809(.A(new_n733), .B1(new_n1009), .B2(new_n751), .ZN(new_n1010));
  OAI22_X1  g0810(.A1(new_n755), .A2(new_n782), .B1(new_n830), .B2(new_n768), .ZN(new_n1011));
  AOI211_X1 g0811(.A(new_n289), .B(new_n1011), .C1(G97), .C2(new_n787), .ZN(new_n1012));
  OAI22_X1  g0812(.A1(new_n762), .A2(new_n201), .B1(new_n760), .B2(new_n203), .ZN(new_n1013));
  AOI21_X1  g0813(.A(new_n1013), .B1(G77), .B2(new_n786), .ZN(new_n1014));
  NAND2_X1  g0814(.A1(new_n780), .A2(new_n475), .ZN(new_n1015));
  NAND3_X1  g0815(.A1(new_n826), .A2(new_n347), .A3(new_n348), .ZN(new_n1016));
  NAND4_X1  g0816(.A1(new_n1012), .A2(new_n1014), .A3(new_n1015), .A4(new_n1016), .ZN(new_n1017));
  AOI21_X1  g0817(.A(new_n335), .B1(new_n834), .B2(G326), .ZN(new_n1018));
  AOI22_X1  g0818(.A1(G322), .A2(new_n756), .B1(new_n791), .B2(G303), .ZN(new_n1019));
  INV_X1    g0819(.A(G317), .ZN(new_n1020));
  OAI221_X1 g0820(.A(new_n1019), .B1(new_n758), .B2(new_n770), .C1(new_n1020), .C2(new_n762), .ZN(new_n1021));
  INV_X1    g0821(.A(KEYINPUT48), .ZN(new_n1022));
  OR2_X1    g0822(.A1(new_n1021), .A2(new_n1022), .ZN(new_n1023));
  NAND2_X1  g0823(.A1(new_n1021), .A2(new_n1022), .ZN(new_n1024));
  AOI22_X1  g0824(.A1(G283), .A2(new_n780), .B1(new_n786), .B2(G294), .ZN(new_n1025));
  NAND3_X1  g0825(.A1(new_n1023), .A2(new_n1024), .A3(new_n1025), .ZN(new_n1026));
  XOR2_X1   g0826(.A(new_n1026), .B(KEYINPUT49), .Z(new_n1027));
  INV_X1    g0827(.A(KEYINPUT109), .ZN(new_n1028));
  OAI221_X1 g0828(.A(new_n1018), .B1(new_n570), .B2(new_n765), .C1(new_n1027), .C2(new_n1028), .ZN(new_n1029));
  AND2_X1   g0829(.A1(new_n1027), .A2(new_n1028), .ZN(new_n1030));
  OAI21_X1  g0830(.A(new_n1017), .B1(new_n1029), .B2(new_n1030), .ZN(new_n1031));
  AOI211_X1 g0831(.A(new_n999), .B(new_n1010), .C1(new_n1031), .C2(new_n746), .ZN(new_n1032));
  AOI21_X1  g0832(.A(new_n1032), .B1(new_n973), .B2(new_n732), .ZN(new_n1033));
  NAND2_X1  g0833(.A1(new_n998), .A2(new_n1033), .ZN(new_n1034));
  INV_X1    g0834(.A(KEYINPUT110), .ZN(new_n1035));
  NAND2_X1  g0835(.A1(new_n1034), .A2(new_n1035), .ZN(new_n1036));
  NAND3_X1  g0836(.A1(new_n998), .A2(KEYINPUT110), .A3(new_n1033), .ZN(new_n1037));
  NAND2_X1  g0837(.A1(new_n1036), .A2(new_n1037), .ZN(G393));
  XNOR2_X1  g0838(.A(new_n967), .B(new_n687), .ZN(new_n1039));
  NAND2_X1  g0839(.A1(new_n1039), .A2(new_n974), .ZN(new_n1040));
  NAND3_X1  g0840(.A1(new_n976), .A2(new_n1040), .A3(new_n696), .ZN(new_n1041));
  OR2_X1    g0841(.A1(new_n1039), .A2(new_n731), .ZN(new_n1042));
  INV_X1    g0842(.A(new_n733), .ZN(new_n1043));
  OAI221_X1 g0843(.A(new_n750), .B1(new_n458), .B2(new_n211), .C1(new_n245), .C2(new_n740), .ZN(new_n1044));
  AOI21_X1  g0844(.A(new_n1043), .B1(new_n1044), .B2(KEYINPUT111), .ZN(new_n1045));
  OAI21_X1  g0845(.A(new_n1045), .B1(KEYINPUT111), .B2(new_n1044), .ZN(new_n1046));
  OAI22_X1  g0846(.A1(new_n762), .A2(new_n782), .B1(new_n755), .B2(new_n830), .ZN(new_n1047));
  XOR2_X1   g0847(.A(new_n1047), .B(KEYINPUT51), .Z(new_n1048));
  OAI22_X1  g0848(.A1(new_n770), .A2(new_n201), .B1(new_n831), .B2(new_n768), .ZN(new_n1049));
  OAI22_X1  g0849(.A1(new_n772), .A2(new_n203), .B1(new_n760), .B2(new_n345), .ZN(new_n1050));
  NAND2_X1  g0850(.A1(new_n780), .A2(G77), .ZN(new_n1051));
  OAI211_X1 g0851(.A(new_n1051), .B(new_n335), .C1(new_n221), .C2(new_n765), .ZN(new_n1052));
  OR4_X1    g0852(.A1(new_n1048), .A2(new_n1049), .A3(new_n1050), .A4(new_n1052), .ZN(new_n1053));
  OAI22_X1  g0853(.A1(new_n772), .A2(new_n766), .B1(new_n761), .B2(new_n768), .ZN(new_n1054));
  AOI211_X1 g0854(.A(new_n335), .B(new_n1054), .C1(G107), .C2(new_n787), .ZN(new_n1055));
  OR2_X1    g0855(.A1(new_n1055), .A2(KEYINPUT112), .ZN(new_n1056));
  NAND2_X1  g0856(.A1(new_n1055), .A2(KEYINPUT112), .ZN(new_n1057));
  OAI22_X1  g0857(.A1(new_n762), .A2(new_n758), .B1(new_n755), .B2(new_n1020), .ZN(new_n1058));
  XNOR2_X1  g0858(.A(new_n1058), .B(KEYINPUT52), .ZN(new_n1059));
  NAND3_X1  g0859(.A1(new_n1056), .A2(new_n1057), .A3(new_n1059), .ZN(new_n1060));
  AOI22_X1  g0860(.A1(G303), .A2(new_n826), .B1(new_n791), .B2(G294), .ZN(new_n1061));
  OAI21_X1  g0861(.A(new_n1061), .B1(new_n570), .B2(new_n775), .ZN(new_n1062));
  XNOR2_X1  g0862(.A(new_n1062), .B(KEYINPUT113), .ZN(new_n1063));
  OAI21_X1  g0863(.A(new_n1053), .B1(new_n1060), .B2(new_n1063), .ZN(new_n1064));
  AOI21_X1  g0864(.A(new_n1046), .B1(new_n1064), .B2(new_n746), .ZN(new_n1065));
  INV_X1    g0865(.A(new_n749), .ZN(new_n1066));
  OAI21_X1  g0866(.A(new_n1065), .B1(new_n962), .B2(new_n1066), .ZN(new_n1067));
  NAND3_X1  g0867(.A1(new_n1041), .A2(new_n1042), .A3(new_n1067), .ZN(G390));
  NAND2_X1  g0868(.A1(new_n918), .A2(new_n747), .ZN(new_n1069));
  AOI22_X1  g0869(.A1(new_n787), .A2(G50), .B1(new_n834), .B2(G125), .ZN(new_n1070));
  INV_X1    g0870(.A(G132), .ZN(new_n1071));
  OAI21_X1  g0871(.A(new_n1070), .B1(new_n1071), .B2(new_n762), .ZN(new_n1072));
  XNOR2_X1  g0872(.A(KEYINPUT54), .B(G143), .ZN(new_n1073));
  OAI21_X1  g0873(.A(new_n335), .B1(new_n760), .B2(new_n1073), .ZN(new_n1074));
  INV_X1    g0874(.A(G128), .ZN(new_n1075));
  OAI22_X1  g0875(.A1(new_n1075), .A2(new_n755), .B1(new_n770), .B2(new_n934), .ZN(new_n1076));
  NOR3_X1   g0876(.A1(new_n1072), .A2(new_n1074), .A3(new_n1076), .ZN(new_n1077));
  NOR2_X1   g0877(.A1(new_n772), .A2(new_n830), .ZN(new_n1078));
  XNOR2_X1  g0878(.A(KEYINPUT115), .B(KEYINPUT53), .ZN(new_n1079));
  AOI22_X1  g0879(.A1(new_n1078), .A2(new_n1079), .B1(new_n780), .B2(G159), .ZN(new_n1080));
  OAI211_X1 g0880(.A(new_n1077), .B(new_n1080), .C1(new_n1078), .C2(new_n1079), .ZN(new_n1081));
  OAI22_X1  g0881(.A1(new_n203), .A2(new_n765), .B1(new_n760), .B2(new_n458), .ZN(new_n1082));
  AOI211_X1 g0882(.A(new_n335), .B(new_n1082), .C1(G87), .C2(new_n786), .ZN(new_n1083));
  AOI22_X1  g0883(.A1(new_n790), .A2(G116), .B1(G294), .B2(new_n834), .ZN(new_n1084));
  AOI22_X1  g0884(.A1(G283), .A2(new_n756), .B1(new_n826), .B2(G107), .ZN(new_n1085));
  NAND4_X1  g0885(.A1(new_n1083), .A2(new_n1051), .A3(new_n1084), .A4(new_n1085), .ZN(new_n1086));
  AOI21_X1  g0886(.A(new_n797), .B1(new_n1081), .B2(new_n1086), .ZN(new_n1087));
  AOI211_X1 g0887(.A(new_n1043), .B(new_n1087), .C1(new_n391), .C2(new_n820), .ZN(new_n1088));
  XOR2_X1   g0888(.A(new_n1088), .B(KEYINPUT116), .Z(new_n1089));
  NAND2_X1  g0889(.A1(new_n1069), .A2(new_n1089), .ZN(new_n1090));
  OAI211_X1 g0890(.A(new_n915), .B(new_n917), .C1(new_n912), .C2(new_n919), .ZN(new_n1091));
  OAI211_X1 g0891(.A(new_n688), .B(new_n812), .C1(new_n723), .C2(new_n725), .ZN(new_n1092));
  NAND2_X1  g0892(.A1(new_n1092), .A2(new_n911), .ZN(new_n1093));
  NAND2_X1  g0893(.A1(new_n860), .A2(new_n1093), .ZN(new_n1094));
  OAI211_X1 g0894(.A(new_n1094), .B(new_n920), .C1(new_n895), .C2(new_n902), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n1091), .A2(new_n1095), .ZN(new_n1096));
  OAI211_X1 g0896(.A(new_n714), .B(new_n812), .C1(new_n853), .C2(new_n855), .ZN(new_n1097));
  INV_X1    g0897(.A(new_n1097), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n1096), .A2(new_n1098), .ZN(new_n1099));
  NAND3_X1  g0899(.A1(new_n1091), .A2(new_n1095), .A3(new_n1097), .ZN(new_n1100));
  NAND2_X1  g0900(.A1(new_n1099), .A2(new_n1100), .ZN(new_n1101));
  OAI21_X1  g0901(.A(new_n1090), .B1(new_n1101), .B2(new_n731), .ZN(new_n1102));
  NAND2_X1  g0902(.A1(new_n456), .A2(new_n714), .ZN(new_n1103));
  NAND4_X1  g0903(.A1(new_n922), .A2(new_n1103), .A3(new_n368), .A4(new_n637), .ZN(new_n1104));
  NAND3_X1  g0904(.A1(new_n851), .A2(G330), .A3(new_n812), .ZN(new_n1105));
  AOI21_X1  g0905(.A(new_n855), .B1(new_n332), .B2(new_n854), .ZN(new_n1106));
  NAND2_X1  g0906(.A1(new_n1105), .A2(new_n1106), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n1107), .A2(new_n1097), .ZN(new_n1108));
  AND2_X1   g0908(.A1(new_n815), .A2(new_n911), .ZN(new_n1109));
  INV_X1    g0909(.A(new_n1109), .ZN(new_n1110));
  NAND2_X1  g0910(.A1(new_n1108), .A2(new_n1110), .ZN(new_n1111));
  NAND4_X1  g0911(.A1(new_n1107), .A2(new_n1097), .A3(new_n911), .A4(new_n1092), .ZN(new_n1112));
  AOI21_X1  g0912(.A(new_n1104), .B1(new_n1111), .B2(new_n1112), .ZN(new_n1113));
  NAND3_X1  g0913(.A1(new_n1099), .A2(new_n1113), .A3(new_n1100), .ZN(new_n1114));
  AND2_X1   g0914(.A1(new_n1114), .A2(new_n696), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n1111), .A2(new_n1112), .ZN(new_n1116));
  INV_X1    g0916(.A(new_n1104), .ZN(new_n1117));
  NAND2_X1  g0917(.A1(new_n1116), .A2(new_n1117), .ZN(new_n1118));
  INV_X1    g0918(.A(KEYINPUT114), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n1118), .A2(new_n1119), .ZN(new_n1120));
  NAND2_X1  g0920(.A1(new_n1113), .A2(KEYINPUT114), .ZN(new_n1121));
  NAND3_X1  g0921(.A1(new_n1120), .A2(new_n1101), .A3(new_n1121), .ZN(new_n1122));
  AOI21_X1  g0922(.A(new_n1102), .B1(new_n1115), .B2(new_n1122), .ZN(new_n1123));
  INV_X1    g0923(.A(new_n1123), .ZN(G378));
  XNOR2_X1  g0924(.A(KEYINPUT118), .B(KEYINPUT56), .ZN(new_n1125));
  XNOR2_X1  g0925(.A(new_n369), .B(new_n1125), .ZN(new_n1126));
  NOR2_X1   g0926(.A1(new_n355), .A2(new_n673), .ZN(new_n1127));
  INV_X1    g0927(.A(new_n1127), .ZN(new_n1128));
  OR2_X1    g0928(.A1(new_n1126), .A2(new_n1128), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n1126), .A2(new_n1128), .ZN(new_n1130));
  XNOR2_X1  g0930(.A(KEYINPUT119), .B(KEYINPUT55), .ZN(new_n1131));
  AND3_X1   g0931(.A1(new_n1129), .A2(new_n1130), .A3(new_n1131), .ZN(new_n1132));
  AOI21_X1  g0932(.A(new_n1131), .B1(new_n1129), .B2(new_n1130), .ZN(new_n1133));
  NOR2_X1   g0933(.A1(new_n1132), .A2(new_n1133), .ZN(new_n1134));
  INV_X1    g0934(.A(new_n1134), .ZN(new_n1135));
  NOR3_X1   g0935(.A1(new_n1109), .A2(new_n882), .A3(new_n1106), .ZN(new_n1136));
  AOI21_X1  g0936(.A(new_n920), .B1(new_n915), .B2(new_n917), .ZN(new_n1137));
  INV_X1    g0937(.A(new_n914), .ZN(new_n1138));
  NOR3_X1   g0938(.A1(new_n1136), .A2(new_n1137), .A3(new_n1138), .ZN(new_n1139));
  AOI21_X1  g0939(.A(new_n882), .B1(new_n856), .B2(KEYINPUT102), .ZN(new_n1140));
  AOI21_X1  g0940(.A(new_n885), .B1(new_n1140), .B2(new_n862), .ZN(new_n1141));
  OAI21_X1  g0941(.A(G330), .B1(new_n903), .B2(new_n904), .ZN(new_n1142));
  NOR3_X1   g0942(.A1(new_n1139), .A2(new_n1141), .A3(new_n1142), .ZN(new_n1143));
  INV_X1    g0943(.A(new_n904), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n901), .A2(new_n888), .ZN(new_n1145));
  INV_X1    g0945(.A(KEYINPUT103), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n1145), .A2(new_n1146), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n1147), .A2(new_n894), .ZN(new_n1148));
  AOI21_X1  g0948(.A(new_n681), .B1(new_n1144), .B2(new_n1148), .ZN(new_n1149));
  AOI21_X1  g0949(.A(new_n921), .B1(new_n887), .B2(new_n1149), .ZN(new_n1150));
  OAI21_X1  g0950(.A(new_n1135), .B1(new_n1143), .B2(new_n1150), .ZN(new_n1151));
  NAND2_X1  g0951(.A1(new_n1114), .A2(new_n1117), .ZN(new_n1152));
  OAI21_X1  g0952(.A(new_n1139), .B1(new_n1141), .B2(new_n1142), .ZN(new_n1153));
  NAND3_X1  g0953(.A1(new_n887), .A2(new_n1149), .A3(new_n921), .ZN(new_n1154));
  NAND3_X1  g0954(.A1(new_n1153), .A2(new_n1154), .A3(new_n1134), .ZN(new_n1155));
  NAND3_X1  g0955(.A1(new_n1151), .A2(new_n1152), .A3(new_n1155), .ZN(new_n1156));
  INV_X1    g0956(.A(KEYINPUT57), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n1156), .A2(new_n1157), .ZN(new_n1158));
  NAND4_X1  g0958(.A1(new_n1151), .A2(new_n1152), .A3(KEYINPUT57), .A4(new_n1155), .ZN(new_n1159));
  NAND3_X1  g0959(.A1(new_n1158), .A2(new_n696), .A3(new_n1159), .ZN(new_n1160));
  NAND3_X1  g0960(.A1(new_n1151), .A2(new_n732), .A3(new_n1155), .ZN(new_n1161));
  NOR2_X1   g0961(.A1(new_n821), .A2(G50), .ZN(new_n1162));
  NAND2_X1  g0962(.A1(new_n790), .A2(G128), .ZN(new_n1163));
  OAI21_X1  g0963(.A(new_n1163), .B1(new_n772), .B2(new_n1073), .ZN(new_n1164));
  AOI22_X1  g0964(.A1(G125), .A2(new_n756), .B1(new_n791), .B2(G137), .ZN(new_n1165));
  OAI21_X1  g0965(.A(new_n1165), .B1(new_n1071), .B2(new_n770), .ZN(new_n1166));
  AOI211_X1 g0966(.A(new_n1164), .B(new_n1166), .C1(G150), .C2(new_n780), .ZN(new_n1167));
  INV_X1    g0967(.A(new_n1167), .ZN(new_n1168));
  OR2_X1    g0968(.A1(new_n1168), .A2(KEYINPUT59), .ZN(new_n1169));
  NAND2_X1  g0969(.A1(new_n1168), .A2(KEYINPUT59), .ZN(new_n1170));
  INV_X1    g0970(.A(KEYINPUT117), .ZN(new_n1171));
  OR2_X1    g0971(.A1(new_n1171), .A2(G124), .ZN(new_n1172));
  NAND2_X1  g0972(.A1(new_n1171), .A2(G124), .ZN(new_n1173));
  NAND3_X1  g0973(.A1(new_n834), .A2(new_n1172), .A3(new_n1173), .ZN(new_n1174));
  NAND3_X1  g0974(.A1(new_n1174), .A2(new_n251), .A3(new_n507), .ZN(new_n1175));
  AOI21_X1  g0975(.A(new_n1175), .B1(G159), .B2(new_n787), .ZN(new_n1176));
  NAND3_X1  g0976(.A1(new_n1169), .A2(new_n1170), .A3(new_n1176), .ZN(new_n1177));
  NAND2_X1  g0977(.A1(new_n289), .A2(new_n507), .ZN(new_n1178));
  OAI22_X1  g0978(.A1(new_n760), .A2(new_n438), .B1(new_n768), .B2(new_n766), .ZN(new_n1179));
  AOI211_X1 g0979(.A(new_n1178), .B(new_n1179), .C1(G77), .C2(new_n786), .ZN(new_n1180));
  AOI22_X1  g0980(.A1(G107), .A2(new_n790), .B1(new_n787), .B2(G58), .ZN(new_n1181));
  AOI22_X1  g0981(.A1(G116), .A2(new_n756), .B1(new_n826), .B2(G97), .ZN(new_n1182));
  AND4_X1   g0982(.A1(new_n941), .A2(new_n1180), .A3(new_n1181), .A4(new_n1182), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n1183), .A2(KEYINPUT58), .ZN(new_n1184));
  OR2_X1    g0984(.A1(new_n1183), .A2(KEYINPUT58), .ZN(new_n1185));
  OAI211_X1 g0985(.A(new_n1178), .B(new_n201), .C1(G33), .C2(G41), .ZN(new_n1186));
  NAND4_X1  g0986(.A1(new_n1177), .A2(new_n1184), .A3(new_n1185), .A4(new_n1186), .ZN(new_n1187));
  AOI211_X1 g0987(.A(new_n1043), .B(new_n1162), .C1(new_n1187), .C2(new_n746), .ZN(new_n1188));
  OAI21_X1  g0988(.A(new_n1188), .B1(new_n1134), .B2(new_n748), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n1161), .A2(new_n1189), .ZN(new_n1190));
  INV_X1    g0990(.A(new_n1190), .ZN(new_n1191));
  NAND2_X1  g0991(.A1(new_n1160), .A2(new_n1191), .ZN(G375));
  NAND3_X1  g0992(.A1(new_n1111), .A2(new_n1104), .A3(new_n1112), .ZN(new_n1193));
  XOR2_X1   g0993(.A(new_n978), .B(KEYINPUT120), .Z(new_n1194));
  NAND4_X1  g0994(.A1(new_n1120), .A2(new_n1121), .A3(new_n1193), .A4(new_n1194), .ZN(new_n1195));
  AOI22_X1  g0995(.A1(G294), .A2(new_n756), .B1(new_n791), .B2(G107), .ZN(new_n1196));
  OAI21_X1  g0996(.A(new_n1196), .B1(new_n570), .B2(new_n770), .ZN(new_n1197));
  XOR2_X1   g0997(.A(new_n1197), .B(KEYINPUT121), .Z(new_n1198));
  OAI22_X1  g0998(.A1(new_n772), .A2(new_n458), .B1(new_n566), .B2(new_n768), .ZN(new_n1199));
  NOR4_X1   g0999(.A1(new_n1198), .A2(new_n335), .A3(new_n937), .A4(new_n1199), .ZN(new_n1200));
  OAI21_X1  g1000(.A(new_n1015), .B1(new_n766), .B2(new_n762), .ZN(new_n1201));
  XOR2_X1   g1001(.A(new_n1201), .B(KEYINPUT122), .Z(new_n1202));
  OAI22_X1  g1002(.A1(new_n775), .A2(new_n201), .B1(new_n760), .B2(new_n830), .ZN(new_n1203));
  XOR2_X1   g1003(.A(new_n1203), .B(KEYINPUT123), .Z(new_n1204));
  OAI22_X1  g1004(.A1(new_n772), .A2(new_n782), .B1(new_n770), .B2(new_n1073), .ZN(new_n1205));
  OAI22_X1  g1005(.A1(new_n762), .A2(new_n934), .B1(new_n1075), .B2(new_n768), .ZN(new_n1206));
  OAI21_X1  g1006(.A(new_n335), .B1(new_n765), .B2(new_n202), .ZN(new_n1207));
  NOR2_X1   g1007(.A1(new_n755), .A2(new_n1071), .ZN(new_n1208));
  NOR4_X1   g1008(.A1(new_n1205), .A2(new_n1206), .A3(new_n1207), .A4(new_n1208), .ZN(new_n1209));
  AOI22_X1  g1009(.A1(new_n1200), .A2(new_n1202), .B1(new_n1204), .B2(new_n1209), .ZN(new_n1210));
  OAI221_X1 g1010(.A(new_n733), .B1(G68), .B2(new_n821), .C1(new_n1210), .C2(new_n797), .ZN(new_n1211));
  AOI21_X1  g1011(.A(new_n1211), .B1(new_n1106), .B2(new_n747), .ZN(new_n1212));
  AOI21_X1  g1012(.A(new_n1212), .B1(new_n1116), .B2(new_n732), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(new_n1195), .A2(new_n1213), .ZN(new_n1214));
  XOR2_X1   g1014(.A(new_n1214), .B(KEYINPUT124), .Z(G381));
  NOR2_X1   g1015(.A1(G387), .A2(G390), .ZN(new_n1216));
  INV_X1    g1016(.A(G384), .ZN(new_n1217));
  NOR2_X1   g1017(.A1(G393), .A2(G396), .ZN(new_n1218));
  NAND3_X1  g1018(.A1(new_n1216), .A2(new_n1217), .A3(new_n1218), .ZN(new_n1219));
  OR4_X1    g1019(.A1(G378), .A2(new_n1219), .A3(G375), .A4(G381), .ZN(G407));
  NAND2_X1  g1020(.A1(new_n674), .A2(G213), .ZN(new_n1221));
  INV_X1    g1021(.A(new_n1221), .ZN(new_n1222));
  NAND2_X1  g1022(.A1(new_n1123), .A2(new_n1222), .ZN(new_n1223));
  OAI211_X1 g1023(.A(G407), .B(G213), .C1(G375), .C2(new_n1223), .ZN(G409));
  INV_X1    g1024(.A(KEYINPUT61), .ZN(new_n1225));
  NAND3_X1  g1025(.A1(new_n1160), .A2(G378), .A3(new_n1191), .ZN(new_n1226));
  AND3_X1   g1026(.A1(new_n1153), .A2(new_n1154), .A3(new_n1134), .ZN(new_n1227));
  AOI21_X1  g1027(.A(new_n1134), .B1(new_n1153), .B2(new_n1154), .ZN(new_n1228));
  OAI21_X1  g1028(.A(KEYINPUT125), .B1(new_n1227), .B2(new_n1228), .ZN(new_n1229));
  INV_X1    g1029(.A(KEYINPUT125), .ZN(new_n1230));
  NAND3_X1  g1030(.A1(new_n1151), .A2(new_n1230), .A3(new_n1155), .ZN(new_n1231));
  AND3_X1   g1031(.A1(new_n1229), .A2(new_n732), .A3(new_n1231), .ZN(new_n1232));
  NAND4_X1  g1032(.A1(new_n1151), .A2(new_n1152), .A3(new_n1155), .A4(new_n1194), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(new_n1233), .A2(new_n1189), .ZN(new_n1234));
  OAI21_X1  g1034(.A(new_n1123), .B1(new_n1232), .B2(new_n1234), .ZN(new_n1235));
  AOI21_X1  g1035(.A(new_n1222), .B1(new_n1226), .B2(new_n1235), .ZN(new_n1236));
  INV_X1    g1036(.A(KEYINPUT60), .ZN(new_n1237));
  OAI211_X1 g1037(.A(new_n1118), .B(new_n696), .C1(new_n1237), .C2(new_n1193), .ZN(new_n1238));
  AND2_X1   g1038(.A1(new_n1193), .A2(new_n1237), .ZN(new_n1239));
  OAI21_X1  g1039(.A(new_n1213), .B1(new_n1238), .B2(new_n1239), .ZN(new_n1240));
  OR2_X1    g1040(.A1(new_n1240), .A2(new_n1217), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(new_n1240), .A2(new_n1217), .ZN(new_n1242));
  AND2_X1   g1042(.A1(new_n1222), .A2(G2897), .ZN(new_n1243));
  AND3_X1   g1043(.A1(new_n1241), .A2(new_n1242), .A3(new_n1243), .ZN(new_n1244));
  AOI21_X1  g1044(.A(new_n1243), .B1(new_n1241), .B2(new_n1242), .ZN(new_n1245));
  NOR2_X1   g1045(.A1(new_n1244), .A2(new_n1245), .ZN(new_n1246));
  OAI21_X1  g1046(.A(new_n1225), .B1(new_n1236), .B2(new_n1246), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n1241), .A2(new_n1242), .ZN(new_n1248));
  INV_X1    g1048(.A(new_n1248), .ZN(new_n1249));
  AOI21_X1  g1049(.A(new_n695), .B1(new_n1156), .B2(new_n1157), .ZN(new_n1250));
  AOI211_X1 g1050(.A(new_n1123), .B(new_n1190), .C1(new_n1250), .C2(new_n1159), .ZN(new_n1251));
  INV_X1    g1051(.A(new_n1234), .ZN(new_n1252));
  NAND3_X1  g1052(.A1(new_n1229), .A2(new_n1231), .A3(new_n732), .ZN(new_n1253));
  AOI21_X1  g1053(.A(G378), .B1(new_n1252), .B2(new_n1253), .ZN(new_n1254));
  OAI211_X1 g1054(.A(new_n1221), .B(new_n1249), .C1(new_n1251), .C2(new_n1254), .ZN(new_n1255));
  INV_X1    g1055(.A(KEYINPUT62), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(new_n1255), .A2(new_n1256), .ZN(new_n1257));
  NAND3_X1  g1057(.A1(new_n1236), .A2(KEYINPUT62), .A3(new_n1249), .ZN(new_n1258));
  AOI21_X1  g1058(.A(new_n1247), .B1(new_n1257), .B2(new_n1258), .ZN(new_n1259));
  INV_X1    g1059(.A(G390), .ZN(new_n1260));
  OAI211_X1 g1060(.A(new_n1260), .B(new_n960), .C1(new_n979), .C2(new_n994), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(G387), .A2(G390), .ZN(new_n1262));
  NAND2_X1  g1062(.A1(new_n1261), .A2(new_n1262), .ZN(new_n1263));
  AOI21_X1  g1063(.A(new_n802), .B1(new_n1036), .B2(new_n1037), .ZN(new_n1264));
  NOR2_X1   g1064(.A1(new_n1218), .A2(new_n1264), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(new_n1263), .A2(new_n1265), .ZN(new_n1266));
  INV_X1    g1066(.A(new_n1265), .ZN(new_n1267));
  NAND3_X1  g1067(.A1(new_n1267), .A2(new_n1261), .A3(new_n1262), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1266), .A2(new_n1268), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n1269), .A2(KEYINPUT127), .ZN(new_n1270));
  INV_X1    g1070(.A(KEYINPUT127), .ZN(new_n1271));
  NAND3_X1  g1071(.A1(new_n1266), .A2(new_n1271), .A3(new_n1268), .ZN(new_n1272));
  NAND2_X1  g1072(.A1(new_n1270), .A2(new_n1272), .ZN(new_n1273));
  INV_X1    g1073(.A(KEYINPUT63), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n1255), .A2(new_n1274), .ZN(new_n1275));
  AND3_X1   g1075(.A1(new_n1266), .A2(new_n1225), .A3(new_n1268), .ZN(new_n1276));
  NAND3_X1  g1076(.A1(new_n1236), .A2(KEYINPUT63), .A3(new_n1249), .ZN(new_n1277));
  NAND3_X1  g1077(.A1(new_n1275), .A2(new_n1276), .A3(new_n1277), .ZN(new_n1278));
  OAI211_X1 g1078(.A(KEYINPUT126), .B(new_n1221), .C1(new_n1251), .C2(new_n1254), .ZN(new_n1279));
  INV_X1    g1079(.A(new_n1246), .ZN(new_n1280));
  NAND2_X1  g1080(.A1(new_n1279), .A2(new_n1280), .ZN(new_n1281));
  NOR2_X1   g1081(.A1(new_n1236), .A2(KEYINPUT126), .ZN(new_n1282));
  NOR2_X1   g1082(.A1(new_n1281), .A2(new_n1282), .ZN(new_n1283));
  OAI22_X1  g1083(.A1(new_n1259), .A2(new_n1273), .B1(new_n1278), .B2(new_n1283), .ZN(G405));
  NAND2_X1  g1084(.A1(G375), .A2(new_n1123), .ZN(new_n1285));
  NAND2_X1  g1085(.A1(new_n1285), .A2(new_n1226), .ZN(new_n1286));
  NAND2_X1  g1086(.A1(new_n1286), .A2(new_n1249), .ZN(new_n1287));
  NAND3_X1  g1087(.A1(new_n1285), .A2(new_n1226), .A3(new_n1248), .ZN(new_n1288));
  NAND2_X1  g1088(.A1(new_n1287), .A2(new_n1288), .ZN(new_n1289));
  XNOR2_X1  g1089(.A(new_n1289), .B(new_n1269), .ZN(G402));
endmodule


