//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 0 1 1 0 0 0 1 0 0 1 0 1 1 1 1 1 0 0 0 1 0 1 1 0 1 0 1 1 0 1 0 0 0 1 0 0 0 1 0 0 0 0 1 1 1 1 0 0 1 0 1 0 1 0 1 1 0 1 1 0 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:23:33 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n702, new_n703,
    new_n704, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n716, new_n717, new_n719, new_n720,
    new_n722, new_n723, new_n724, new_n725, new_n726, new_n727, new_n728,
    new_n730, new_n731, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n761, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n790, new_n791, new_n792, new_n793, new_n794, new_n795, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n913, new_n914, new_n915, new_n916, new_n918, new_n919, new_n920,
    new_n921, new_n922, new_n923, new_n924, new_n925, new_n926, new_n927,
    new_n928, new_n929, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n951, new_n952, new_n953, new_n954, new_n955, new_n957,
    new_n958, new_n959, new_n960, new_n961, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015;
  OAI21_X1  g000(.A(G214), .B1(G237), .B2(G902), .ZN(new_n187));
  INV_X1    g001(.A(KEYINPUT79), .ZN(new_n188));
  INV_X1    g002(.A(G107), .ZN(new_n189));
  OAI21_X1  g003(.A(new_n188), .B1(new_n189), .B2(G104), .ZN(new_n190));
  INV_X1    g004(.A(G104), .ZN(new_n191));
  NAND3_X1  g005(.A1(new_n191), .A2(KEYINPUT79), .A3(G107), .ZN(new_n192));
  AND3_X1   g006(.A1(new_n189), .A2(KEYINPUT3), .A3(G104), .ZN(new_n193));
  AOI21_X1  g007(.A(KEYINPUT3), .B1(new_n189), .B2(G104), .ZN(new_n194));
  OAI211_X1 g008(.A(new_n190), .B(new_n192), .C1(new_n193), .C2(new_n194), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n195), .A2(G101), .ZN(new_n196));
  INV_X1    g010(.A(KEYINPUT3), .ZN(new_n197));
  OAI21_X1  g011(.A(new_n197), .B1(new_n191), .B2(G107), .ZN(new_n198));
  NAND3_X1  g012(.A1(new_n189), .A2(KEYINPUT3), .A3(G104), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n198), .A2(new_n199), .ZN(new_n200));
  INV_X1    g014(.A(G101), .ZN(new_n201));
  NAND4_X1  g015(.A1(new_n200), .A2(new_n201), .A3(new_n190), .A4(new_n192), .ZN(new_n202));
  NAND3_X1  g016(.A1(new_n196), .A2(KEYINPUT4), .A3(new_n202), .ZN(new_n203));
  XOR2_X1   g017(.A(KEYINPUT2), .B(G113), .Z(new_n204));
  XNOR2_X1  g018(.A(G116), .B(G119), .ZN(new_n205));
  OR2_X1    g019(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n204), .A2(new_n205), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  INV_X1    g022(.A(KEYINPUT4), .ZN(new_n209));
  NAND3_X1  g023(.A1(new_n195), .A2(new_n209), .A3(G101), .ZN(new_n210));
  NAND3_X1  g024(.A1(new_n203), .A2(new_n208), .A3(new_n210), .ZN(new_n211));
  XNOR2_X1  g025(.A(G110), .B(G122), .ZN(new_n212));
  NOR2_X1   g026(.A1(new_n191), .A2(G107), .ZN(new_n213));
  NOR2_X1   g027(.A1(new_n189), .A2(G104), .ZN(new_n214));
  OAI21_X1  g028(.A(G101), .B1(new_n213), .B2(new_n214), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n202), .A2(new_n215), .ZN(new_n216));
  INV_X1    g030(.A(G119), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n217), .A2(G116), .ZN(new_n218));
  INV_X1    g032(.A(G116), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n219), .A2(G119), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n218), .A2(new_n220), .ZN(new_n221));
  INV_X1    g035(.A(KEYINPUT5), .ZN(new_n222));
  NOR2_X1   g036(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  OAI21_X1  g037(.A(G113), .B1(new_n218), .B2(KEYINPUT5), .ZN(new_n224));
  OAI21_X1  g038(.A(new_n207), .B1(new_n223), .B2(new_n224), .ZN(new_n225));
  OR2_X1    g039(.A1(new_n216), .A2(new_n225), .ZN(new_n226));
  NAND3_X1  g040(.A1(new_n211), .A2(new_n212), .A3(new_n226), .ZN(new_n227));
  XNOR2_X1  g041(.A(KEYINPUT69), .B(KEYINPUT1), .ZN(new_n228));
  INV_X1    g042(.A(G146), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n229), .A2(G143), .ZN(new_n230));
  INV_X1    g044(.A(new_n230), .ZN(new_n231));
  OAI21_X1  g045(.A(G128), .B1(new_n228), .B2(new_n231), .ZN(new_n232));
  INV_X1    g046(.A(G143), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n233), .A2(G146), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n230), .A2(new_n234), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n232), .A2(new_n235), .ZN(new_n236));
  INV_X1    g050(.A(KEYINPUT64), .ZN(new_n237));
  OAI21_X1  g051(.A(new_n237), .B1(new_n233), .B2(G146), .ZN(new_n238));
  NAND3_X1  g052(.A1(new_n229), .A2(KEYINPUT64), .A3(G143), .ZN(new_n239));
  AND3_X1   g053(.A1(new_n238), .A2(new_n239), .A3(new_n234), .ZN(new_n240));
  INV_X1    g054(.A(KEYINPUT1), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n241), .A2(KEYINPUT69), .ZN(new_n242));
  INV_X1    g056(.A(KEYINPUT69), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n243), .A2(KEYINPUT1), .ZN(new_n244));
  NAND3_X1  g058(.A1(new_n242), .A2(new_n244), .A3(G128), .ZN(new_n245));
  INV_X1    g059(.A(new_n245), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n240), .A2(new_n246), .ZN(new_n247));
  INV_X1    g061(.A(G125), .ZN(new_n248));
  NAND3_X1  g062(.A1(new_n236), .A2(new_n247), .A3(new_n248), .ZN(new_n249));
  NAND2_X1  g063(.A1(KEYINPUT0), .A2(G128), .ZN(new_n250));
  OR2_X1    g064(.A1(KEYINPUT0), .A2(G128), .ZN(new_n251));
  AND3_X1   g065(.A1(new_n235), .A2(new_n250), .A3(new_n251), .ZN(new_n252));
  AND2_X1   g066(.A1(new_n239), .A2(new_n234), .ZN(new_n253));
  INV_X1    g067(.A(KEYINPUT65), .ZN(new_n254));
  INV_X1    g068(.A(new_n250), .ZN(new_n255));
  NAND4_X1  g069(.A1(new_n253), .A2(new_n254), .A3(new_n255), .A4(new_n238), .ZN(new_n256));
  NAND4_X1  g070(.A1(new_n238), .A2(new_n239), .A3(new_n255), .A4(new_n234), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n257), .A2(KEYINPUT65), .ZN(new_n258));
  AOI21_X1  g072(.A(new_n252), .B1(new_n256), .B2(new_n258), .ZN(new_n259));
  OAI21_X1  g073(.A(new_n249), .B1(new_n259), .B2(new_n248), .ZN(new_n260));
  INV_X1    g074(.A(G953), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n261), .A2(G224), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n262), .A2(KEYINPUT7), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n260), .A2(new_n263), .ZN(new_n264));
  INV_X1    g078(.A(KEYINPUT85), .ZN(new_n265));
  OAI21_X1  g079(.A(KEYINPUT7), .B1(new_n262), .B2(new_n265), .ZN(new_n266));
  AOI21_X1  g080(.A(new_n266), .B1(new_n265), .B2(new_n262), .ZN(new_n267));
  OAI211_X1 g081(.A(new_n249), .B(new_n267), .C1(new_n259), .C2(new_n248), .ZN(new_n268));
  AND3_X1   g082(.A1(new_n227), .A2(new_n264), .A3(new_n268), .ZN(new_n269));
  XNOR2_X1  g083(.A(new_n212), .B(KEYINPUT8), .ZN(new_n270));
  AND2_X1   g084(.A1(new_n202), .A2(new_n215), .ZN(new_n271));
  OAI21_X1  g085(.A(KEYINPUT83), .B1(new_n221), .B2(new_n222), .ZN(new_n272));
  INV_X1    g086(.A(new_n224), .ZN(new_n273));
  INV_X1    g087(.A(KEYINPUT83), .ZN(new_n274));
  NAND3_X1  g088(.A1(new_n205), .A2(new_n274), .A3(KEYINPUT5), .ZN(new_n275));
  NAND3_X1  g089(.A1(new_n272), .A2(new_n273), .A3(new_n275), .ZN(new_n276));
  NAND3_X1  g090(.A1(new_n271), .A2(new_n207), .A3(new_n276), .ZN(new_n277));
  AND2_X1   g091(.A1(new_n277), .A2(KEYINPUT84), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n216), .A2(new_n225), .ZN(new_n279));
  OAI21_X1  g093(.A(new_n279), .B1(new_n277), .B2(KEYINPUT84), .ZN(new_n280));
  OAI21_X1  g094(.A(new_n270), .B1(new_n278), .B2(new_n280), .ZN(new_n281));
  AOI21_X1  g095(.A(G902), .B1(new_n269), .B2(new_n281), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n211), .A2(new_n226), .ZN(new_n283));
  INV_X1    g097(.A(new_n212), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  NAND3_X1  g099(.A1(new_n285), .A2(KEYINPUT6), .A3(new_n227), .ZN(new_n286));
  XOR2_X1   g100(.A(new_n262), .B(KEYINPUT82), .Z(new_n287));
  INV_X1    g101(.A(new_n287), .ZN(new_n288));
  XNOR2_X1  g102(.A(new_n260), .B(new_n288), .ZN(new_n289));
  INV_X1    g103(.A(KEYINPUT6), .ZN(new_n290));
  NAND3_X1  g104(.A1(new_n283), .A2(new_n290), .A3(new_n284), .ZN(new_n291));
  NAND3_X1  g105(.A1(new_n286), .A2(new_n289), .A3(new_n291), .ZN(new_n292));
  OAI21_X1  g106(.A(G210), .B1(G237), .B2(G902), .ZN(new_n293));
  AND3_X1   g107(.A1(new_n282), .A2(new_n292), .A3(new_n293), .ZN(new_n294));
  AOI21_X1  g108(.A(new_n293), .B1(new_n282), .B2(new_n292), .ZN(new_n295));
  OAI21_X1  g109(.A(new_n187), .B1(new_n294), .B2(new_n295), .ZN(new_n296));
  INV_X1    g110(.A(G902), .ZN(new_n297));
  XNOR2_X1  g111(.A(G116), .B(G122), .ZN(new_n298));
  INV_X1    g112(.A(KEYINPUT89), .ZN(new_n299));
  AND3_X1   g113(.A1(new_n298), .A2(new_n299), .A3(new_n189), .ZN(new_n300));
  AOI21_X1  g114(.A(new_n299), .B1(new_n298), .B2(new_n189), .ZN(new_n301));
  NOR2_X1   g115(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  INV_X1    g116(.A(G122), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n303), .A2(G116), .ZN(new_n304));
  INV_X1    g118(.A(KEYINPUT14), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  INV_X1    g120(.A(KEYINPUT90), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n219), .A2(G122), .ZN(new_n308));
  NAND3_X1  g122(.A1(new_n306), .A2(new_n307), .A3(new_n308), .ZN(new_n309));
  NOR2_X1   g123(.A1(new_n303), .A2(G116), .ZN(new_n310));
  AOI21_X1  g124(.A(new_n310), .B1(new_n305), .B2(new_n304), .ZN(new_n311));
  OAI21_X1  g125(.A(KEYINPUT90), .B1(new_n308), .B2(KEYINPUT14), .ZN(new_n312));
  OAI211_X1 g126(.A(new_n309), .B(G107), .C1(new_n311), .C2(new_n312), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n233), .A2(G128), .ZN(new_n314));
  INV_X1    g128(.A(G128), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n315), .A2(G143), .ZN(new_n316));
  AOI21_X1  g130(.A(KEYINPUT88), .B1(new_n314), .B2(new_n316), .ZN(new_n317));
  INV_X1    g131(.A(new_n317), .ZN(new_n318));
  XNOR2_X1  g132(.A(G128), .B(G143), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n319), .A2(KEYINPUT88), .ZN(new_n320));
  AOI21_X1  g134(.A(G134), .B1(new_n318), .B2(new_n320), .ZN(new_n321));
  AND3_X1   g135(.A1(new_n314), .A2(new_n316), .A3(KEYINPUT88), .ZN(new_n322));
  INV_X1    g136(.A(G134), .ZN(new_n323));
  NOR3_X1   g137(.A1(new_n322), .A2(new_n317), .A3(new_n323), .ZN(new_n324));
  OAI211_X1 g138(.A(new_n302), .B(new_n313), .C1(new_n321), .C2(new_n324), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n319), .A2(KEYINPUT13), .ZN(new_n326));
  OAI211_X1 g140(.A(new_n326), .B(G134), .C1(KEYINPUT13), .C2(new_n314), .ZN(new_n327));
  XNOR2_X1  g141(.A(new_n298), .B(new_n189), .ZN(new_n328));
  OAI21_X1  g142(.A(new_n323), .B1(new_n322), .B2(new_n317), .ZN(new_n329));
  NAND3_X1  g143(.A1(new_n327), .A2(new_n328), .A3(new_n329), .ZN(new_n330));
  XNOR2_X1  g144(.A(KEYINPUT9), .B(G234), .ZN(new_n331));
  INV_X1    g145(.A(G217), .ZN(new_n332));
  NOR3_X1   g146(.A1(new_n331), .A2(new_n332), .A3(G953), .ZN(new_n333));
  AND3_X1   g147(.A1(new_n325), .A2(new_n330), .A3(new_n333), .ZN(new_n334));
  AOI21_X1  g148(.A(new_n333), .B1(new_n325), .B2(new_n330), .ZN(new_n335));
  OAI21_X1  g149(.A(new_n297), .B1(new_n334), .B2(new_n335), .ZN(new_n336));
  INV_X1    g150(.A(G478), .ZN(new_n337));
  NOR2_X1   g151(.A1(new_n337), .A2(KEYINPUT15), .ZN(new_n338));
  OR2_X1    g152(.A1(new_n336), .A2(new_n338), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n336), .A2(new_n338), .ZN(new_n340));
  AND2_X1   g154(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  NOR2_X1   g155(.A1(G475), .A2(G902), .ZN(new_n342));
  XNOR2_X1  g156(.A(G113), .B(G122), .ZN(new_n343));
  XNOR2_X1  g157(.A(new_n343), .B(new_n191), .ZN(new_n344));
  INV_X1    g158(.A(G140), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n345), .A2(G125), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n248), .A2(G140), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n346), .A2(new_n347), .ZN(new_n348));
  INV_X1    g162(.A(KEYINPUT19), .ZN(new_n349));
  NOR2_X1   g163(.A1(new_n348), .A2(new_n349), .ZN(new_n350));
  XNOR2_X1  g164(.A(G125), .B(G140), .ZN(new_n351));
  NOR2_X1   g165(.A1(new_n351), .A2(KEYINPUT19), .ZN(new_n352));
  OAI21_X1  g166(.A(new_n229), .B1(new_n350), .B2(new_n352), .ZN(new_n353));
  NAND3_X1  g167(.A1(new_n346), .A2(new_n347), .A3(KEYINPUT16), .ZN(new_n354));
  OR3_X1    g168(.A1(new_n248), .A2(KEYINPUT16), .A3(G140), .ZN(new_n355));
  NAND3_X1  g169(.A1(new_n354), .A2(new_n355), .A3(G146), .ZN(new_n356));
  NAND3_X1  g170(.A1(new_n353), .A2(KEYINPUT86), .A3(new_n356), .ZN(new_n357));
  INV_X1    g171(.A(KEYINPUT86), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n348), .A2(new_n349), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n351), .A2(KEYINPUT19), .ZN(new_n360));
  AOI21_X1  g174(.A(G146), .B1(new_n359), .B2(new_n360), .ZN(new_n361));
  INV_X1    g175(.A(new_n356), .ZN(new_n362));
  OAI21_X1  g176(.A(new_n358), .B1(new_n361), .B2(new_n362), .ZN(new_n363));
  NOR2_X1   g177(.A1(G237), .A2(G953), .ZN(new_n364));
  NAND3_X1  g178(.A1(new_n364), .A2(G143), .A3(G214), .ZN(new_n365));
  INV_X1    g179(.A(new_n365), .ZN(new_n366));
  AOI21_X1  g180(.A(G143), .B1(new_n364), .B2(G214), .ZN(new_n367));
  OAI21_X1  g181(.A(G131), .B1(new_n366), .B2(new_n367), .ZN(new_n368));
  INV_X1    g182(.A(new_n367), .ZN(new_n369));
  INV_X1    g183(.A(G131), .ZN(new_n370));
  NAND3_X1  g184(.A1(new_n369), .A2(new_n370), .A3(new_n365), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n368), .A2(new_n371), .ZN(new_n372));
  NAND3_X1  g186(.A1(new_n357), .A2(new_n363), .A3(new_n372), .ZN(new_n373));
  XNOR2_X1  g187(.A(new_n351), .B(new_n229), .ZN(new_n374));
  OAI211_X1 g188(.A(KEYINPUT18), .B(G131), .C1(new_n366), .C2(new_n367), .ZN(new_n375));
  NAND2_X1  g189(.A1(KEYINPUT18), .A2(G131), .ZN(new_n376));
  NAND3_X1  g190(.A1(new_n369), .A2(new_n365), .A3(new_n376), .ZN(new_n377));
  NAND3_X1  g191(.A1(new_n374), .A2(new_n375), .A3(new_n377), .ZN(new_n378));
  AOI21_X1  g192(.A(new_n344), .B1(new_n373), .B2(new_n378), .ZN(new_n379));
  INV_X1    g193(.A(KEYINPUT17), .ZN(new_n380));
  NAND3_X1  g194(.A1(new_n368), .A2(new_n371), .A3(new_n380), .ZN(new_n381));
  INV_X1    g195(.A(new_n381), .ZN(new_n382));
  OAI211_X1 g196(.A(KEYINPUT17), .B(G131), .C1(new_n366), .C2(new_n367), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n354), .A2(new_n355), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n384), .A2(new_n229), .ZN(new_n385));
  NAND3_X1  g199(.A1(new_n383), .A2(new_n385), .A3(new_n356), .ZN(new_n386));
  OAI211_X1 g200(.A(new_n344), .B(new_n378), .C1(new_n382), .C2(new_n386), .ZN(new_n387));
  INV_X1    g201(.A(new_n387), .ZN(new_n388));
  OAI21_X1  g202(.A(new_n342), .B1(new_n379), .B2(new_n388), .ZN(new_n389));
  XOR2_X1   g203(.A(KEYINPUT87), .B(KEYINPUT20), .Z(new_n390));
  INV_X1    g204(.A(new_n390), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n389), .A2(new_n391), .ZN(new_n392));
  NAND2_X1  g206(.A1(KEYINPUT87), .A2(KEYINPUT20), .ZN(new_n393));
  OAI211_X1 g207(.A(new_n342), .B(new_n393), .C1(new_n379), .C2(new_n388), .ZN(new_n394));
  NAND4_X1  g208(.A1(new_n381), .A2(new_n385), .A3(new_n356), .A4(new_n383), .ZN(new_n395));
  AOI21_X1  g209(.A(new_n344), .B1(new_n395), .B2(new_n378), .ZN(new_n396));
  OAI21_X1  g210(.A(new_n297), .B1(new_n388), .B2(new_n396), .ZN(new_n397));
  AOI22_X1  g211(.A1(new_n392), .A2(new_n394), .B1(G475), .B2(new_n397), .ZN(new_n398));
  INV_X1    g212(.A(G234), .ZN(new_n399));
  INV_X1    g213(.A(G237), .ZN(new_n400));
  OAI211_X1 g214(.A(G952), .B(new_n261), .C1(new_n399), .C2(new_n400), .ZN(new_n401));
  XNOR2_X1  g215(.A(new_n401), .B(KEYINPUT91), .ZN(new_n402));
  OAI211_X1 g216(.A(G902), .B(G953), .C1(new_n399), .C2(new_n400), .ZN(new_n403));
  XOR2_X1   g217(.A(new_n403), .B(KEYINPUT92), .Z(new_n404));
  XNOR2_X1  g218(.A(KEYINPUT21), .B(G898), .ZN(new_n405));
  AOI21_X1  g219(.A(new_n402), .B1(new_n404), .B2(new_n405), .ZN(new_n406));
  INV_X1    g220(.A(new_n406), .ZN(new_n407));
  NAND3_X1  g221(.A1(new_n341), .A2(new_n398), .A3(new_n407), .ZN(new_n408));
  NOR2_X1   g222(.A1(new_n296), .A2(new_n408), .ZN(new_n409));
  INV_X1    g223(.A(G221), .ZN(new_n410));
  INV_X1    g224(.A(new_n331), .ZN(new_n411));
  AOI21_X1  g225(.A(new_n410), .B1(new_n411), .B2(new_n297), .ZN(new_n412));
  INV_X1    g226(.A(new_n412), .ZN(new_n413));
  NAND3_X1  g227(.A1(new_n216), .A2(new_n247), .A3(new_n236), .ZN(new_n414));
  AOI21_X1  g228(.A(new_n315), .B1(new_n230), .B2(KEYINPUT1), .ZN(new_n415));
  AOI21_X1  g229(.A(new_n415), .B1(new_n253), .B2(new_n238), .ZN(new_n416));
  NAND3_X1  g230(.A1(new_n238), .A2(new_n239), .A3(new_n234), .ZN(new_n417));
  NOR2_X1   g231(.A1(new_n417), .A2(new_n245), .ZN(new_n418));
  OAI211_X1 g232(.A(new_n202), .B(new_n215), .C1(new_n416), .C2(new_n418), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n414), .A2(new_n419), .ZN(new_n420));
  NAND2_X1  g234(.A1(KEYINPUT11), .A2(G134), .ZN(new_n421));
  OAI21_X1  g235(.A(KEYINPUT67), .B1(new_n421), .B2(G137), .ZN(new_n422));
  INV_X1    g236(.A(KEYINPUT67), .ZN(new_n423));
  INV_X1    g237(.A(G137), .ZN(new_n424));
  NAND4_X1  g238(.A1(new_n423), .A2(new_n424), .A3(KEYINPUT11), .A4(G134), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n422), .A2(new_n425), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n323), .A2(G137), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n424), .A2(G134), .ZN(new_n428));
  INV_X1    g242(.A(KEYINPUT11), .ZN(new_n429));
  AOI21_X1  g243(.A(KEYINPUT66), .B1(new_n428), .B2(new_n429), .ZN(new_n430));
  OAI211_X1 g244(.A(KEYINPUT66), .B(new_n429), .C1(new_n323), .C2(G137), .ZN(new_n431));
  INV_X1    g245(.A(new_n431), .ZN(new_n432));
  OAI211_X1 g246(.A(new_n426), .B(new_n427), .C1(new_n430), .C2(new_n432), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n433), .A2(G131), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n427), .A2(new_n370), .ZN(new_n435));
  INV_X1    g249(.A(new_n435), .ZN(new_n436));
  OAI211_X1 g250(.A(new_n426), .B(new_n436), .C1(new_n430), .C2(new_n432), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n434), .A2(new_n437), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n420), .A2(new_n438), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n439), .A2(KEYINPUT12), .ZN(new_n440));
  NAND3_X1  g254(.A1(new_n203), .A2(new_n259), .A3(new_n210), .ZN(new_n441));
  INV_X1    g255(.A(KEYINPUT10), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n419), .A2(new_n442), .ZN(new_n443));
  AOI21_X1  g257(.A(new_n442), .B1(new_n236), .B2(new_n247), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n444), .A2(new_n271), .ZN(new_n445));
  OAI21_X1  g259(.A(new_n429), .B1(new_n323), .B2(G137), .ZN(new_n446));
  INV_X1    g260(.A(KEYINPUT66), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n446), .A2(new_n447), .ZN(new_n448));
  AOI22_X1  g262(.A1(new_n448), .A2(new_n431), .B1(new_n422), .B2(new_n425), .ZN(new_n449));
  AOI22_X1  g263(.A1(new_n433), .A2(G131), .B1(new_n449), .B2(new_n436), .ZN(new_n450));
  NAND4_X1  g264(.A1(new_n441), .A2(new_n443), .A3(new_n445), .A4(new_n450), .ZN(new_n451));
  INV_X1    g265(.A(KEYINPUT12), .ZN(new_n452));
  NAND3_X1  g266(.A1(new_n420), .A2(new_n452), .A3(new_n438), .ZN(new_n453));
  NAND3_X1  g267(.A1(new_n440), .A2(new_n451), .A3(new_n453), .ZN(new_n454));
  XNOR2_X1  g268(.A(G110), .B(G140), .ZN(new_n455));
  AND2_X1   g269(.A1(new_n261), .A2(G227), .ZN(new_n456));
  XNOR2_X1  g270(.A(new_n455), .B(new_n456), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n454), .A2(new_n457), .ZN(new_n458));
  NAND3_X1  g272(.A1(new_n441), .A2(new_n443), .A3(new_n445), .ZN(new_n459));
  AOI21_X1  g273(.A(new_n370), .B1(new_n449), .B2(new_n427), .ZN(new_n460));
  INV_X1    g274(.A(new_n437), .ZN(new_n461));
  OAI21_X1  g275(.A(KEYINPUT80), .B1(new_n460), .B2(new_n461), .ZN(new_n462));
  INV_X1    g276(.A(new_n462), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n459), .A2(new_n463), .ZN(new_n464));
  AOI22_X1  g278(.A1(new_n442), .A2(new_n419), .B1(new_n444), .B2(new_n271), .ZN(new_n465));
  NAND3_X1  g279(.A1(new_n465), .A2(new_n441), .A3(new_n462), .ZN(new_n466));
  INV_X1    g280(.A(new_n457), .ZN(new_n467));
  NAND3_X1  g281(.A1(new_n464), .A2(new_n466), .A3(new_n467), .ZN(new_n468));
  NAND3_X1  g282(.A1(new_n458), .A2(G469), .A3(new_n468), .ZN(new_n469));
  NAND2_X1  g283(.A1(G469), .A2(G902), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  AOI21_X1  g285(.A(new_n462), .B1(new_n465), .B2(new_n441), .ZN(new_n472));
  AND4_X1   g286(.A1(new_n441), .A2(new_n462), .A3(new_n443), .A4(new_n445), .ZN(new_n473));
  OAI21_X1  g287(.A(new_n457), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  NAND4_X1  g288(.A1(new_n440), .A2(new_n467), .A3(new_n451), .A4(new_n453), .ZN(new_n475));
  AOI211_X1 g289(.A(G469), .B(G902), .C1(new_n474), .C2(new_n475), .ZN(new_n476));
  OAI211_X1 g290(.A(KEYINPUT81), .B(new_n413), .C1(new_n471), .C2(new_n476), .ZN(new_n477));
  INV_X1    g291(.A(new_n477), .ZN(new_n478));
  INV_X1    g292(.A(G469), .ZN(new_n479));
  INV_X1    g293(.A(new_n475), .ZN(new_n480));
  AOI21_X1  g294(.A(new_n467), .B1(new_n464), .B2(new_n466), .ZN(new_n481));
  OAI211_X1 g295(.A(new_n479), .B(new_n297), .C1(new_n480), .C2(new_n481), .ZN(new_n482));
  NAND3_X1  g296(.A1(new_n482), .A2(new_n470), .A3(new_n469), .ZN(new_n483));
  AOI21_X1  g297(.A(KEYINPUT81), .B1(new_n483), .B2(new_n413), .ZN(new_n484));
  OAI21_X1  g298(.A(new_n409), .B1(new_n478), .B2(new_n484), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n485), .A2(KEYINPUT93), .ZN(new_n486));
  OAI21_X1  g300(.A(new_n413), .B1(new_n471), .B2(new_n476), .ZN(new_n487));
  INV_X1    g301(.A(KEYINPUT81), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n489), .A2(new_n477), .ZN(new_n490));
  INV_X1    g304(.A(KEYINPUT93), .ZN(new_n491));
  NAND3_X1  g305(.A1(new_n490), .A2(new_n491), .A3(new_n409), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n486), .A2(new_n492), .ZN(new_n493));
  AOI21_X1  g307(.A(new_n332), .B1(G234), .B2(new_n297), .ZN(new_n494));
  XNOR2_X1  g308(.A(KEYINPUT22), .B(G137), .ZN(new_n495));
  NOR3_X1   g309(.A1(new_n410), .A2(new_n399), .A3(G953), .ZN(new_n496));
  XOR2_X1   g310(.A(new_n495), .B(new_n496), .Z(new_n497));
  XNOR2_X1  g311(.A(G119), .B(G128), .ZN(new_n498));
  XOR2_X1   g312(.A(KEYINPUT24), .B(G110), .Z(new_n499));
  AOI22_X1  g313(.A1(new_n385), .A2(new_n356), .B1(new_n498), .B2(new_n499), .ZN(new_n500));
  INV_X1    g314(.A(KEYINPUT23), .ZN(new_n501));
  OAI21_X1  g315(.A(new_n501), .B1(new_n217), .B2(G128), .ZN(new_n502));
  NAND3_X1  g316(.A1(new_n315), .A2(KEYINPUT23), .A3(G119), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n217), .A2(G128), .ZN(new_n504));
  NAND3_X1  g318(.A1(new_n502), .A2(new_n503), .A3(new_n504), .ZN(new_n505));
  INV_X1    g319(.A(KEYINPUT75), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  NAND4_X1  g321(.A1(new_n502), .A2(new_n503), .A3(KEYINPUT75), .A4(new_n504), .ZN(new_n508));
  NAND3_X1  g322(.A1(new_n507), .A2(G110), .A3(new_n508), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n509), .A2(KEYINPUT76), .ZN(new_n510));
  INV_X1    g324(.A(KEYINPUT76), .ZN(new_n511));
  NAND4_X1  g325(.A1(new_n507), .A2(new_n511), .A3(G110), .A4(new_n508), .ZN(new_n512));
  NAND3_X1  g326(.A1(new_n500), .A2(new_n510), .A3(new_n512), .ZN(new_n513));
  OAI22_X1  g327(.A1(new_n505), .A2(G110), .B1(new_n499), .B2(new_n498), .ZN(new_n514));
  OAI211_X1 g328(.A(new_n514), .B(new_n356), .C1(G146), .C2(new_n348), .ZN(new_n515));
  AND3_X1   g329(.A1(new_n513), .A2(KEYINPUT77), .A3(new_n515), .ZN(new_n516));
  AOI21_X1  g330(.A(KEYINPUT77), .B1(new_n513), .B2(new_n515), .ZN(new_n517));
  OAI21_X1  g331(.A(new_n497), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  INV_X1    g332(.A(new_n497), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n513), .A2(new_n515), .ZN(new_n520));
  INV_X1    g334(.A(KEYINPUT77), .ZN(new_n521));
  OAI21_X1  g335(.A(new_n519), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  NAND3_X1  g336(.A1(new_n518), .A2(new_n297), .A3(new_n522), .ZN(new_n523));
  INV_X1    g337(.A(KEYINPUT78), .ZN(new_n524));
  NOR2_X1   g338(.A1(new_n524), .A2(KEYINPUT25), .ZN(new_n525));
  AND2_X1   g339(.A1(new_n523), .A2(new_n525), .ZN(new_n526));
  NOR2_X1   g340(.A1(new_n523), .A2(new_n525), .ZN(new_n527));
  OAI21_X1  g341(.A(new_n494), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  AND2_X1   g342(.A1(new_n518), .A2(new_n522), .ZN(new_n529));
  NOR2_X1   g343(.A1(new_n494), .A2(G902), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n528), .A2(new_n531), .ZN(new_n532));
  XNOR2_X1  g346(.A(KEYINPUT72), .B(KEYINPUT32), .ZN(new_n533));
  INV_X1    g347(.A(new_n252), .ZN(new_n534));
  AND2_X1   g348(.A1(new_n257), .A2(KEYINPUT65), .ZN(new_n535));
  NOR2_X1   g349(.A1(new_n257), .A2(KEYINPUT65), .ZN(new_n536));
  OAI21_X1  g350(.A(new_n534), .B1(new_n535), .B2(new_n536), .ZN(new_n537));
  NOR2_X1   g351(.A1(new_n450), .A2(new_n537), .ZN(new_n538));
  AND2_X1   g352(.A1(new_n206), .A2(new_n207), .ZN(new_n539));
  XNOR2_X1  g353(.A(G134), .B(G137), .ZN(new_n540));
  OAI21_X1  g354(.A(KEYINPUT68), .B1(new_n540), .B2(new_n370), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n428), .A2(new_n427), .ZN(new_n542));
  INV_X1    g356(.A(KEYINPUT68), .ZN(new_n543));
  NAND3_X1  g357(.A1(new_n542), .A2(new_n543), .A3(G131), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n541), .A2(new_n544), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n545), .A2(new_n437), .ZN(new_n546));
  AOI22_X1  g360(.A1(new_n235), .A2(new_n232), .B1(new_n240), .B2(new_n246), .ZN(new_n547));
  OAI21_X1  g361(.A(new_n539), .B1(new_n546), .B2(new_n547), .ZN(new_n548));
  OAI21_X1  g362(.A(KEYINPUT70), .B1(new_n538), .B2(new_n548), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n242), .A2(new_n244), .ZN(new_n550));
  AOI21_X1  g364(.A(new_n315), .B1(new_n550), .B2(new_n230), .ZN(new_n551));
  INV_X1    g365(.A(new_n235), .ZN(new_n552));
  NOR2_X1   g366(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  OAI211_X1 g367(.A(new_n437), .B(new_n545), .C1(new_n553), .C2(new_n418), .ZN(new_n554));
  OAI21_X1  g368(.A(new_n554), .B1(new_n450), .B2(new_n537), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n555), .A2(new_n208), .ZN(new_n556));
  OAI21_X1  g370(.A(new_n259), .B1(new_n460), .B2(new_n461), .ZN(new_n557));
  INV_X1    g371(.A(KEYINPUT70), .ZN(new_n558));
  NAND4_X1  g372(.A1(new_n557), .A2(new_n558), .A3(new_n539), .A4(new_n554), .ZN(new_n559));
  NAND3_X1  g373(.A1(new_n549), .A2(new_n556), .A3(new_n559), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n560), .A2(KEYINPUT28), .ZN(new_n561));
  INV_X1    g375(.A(KEYINPUT28), .ZN(new_n562));
  OAI21_X1  g376(.A(new_n562), .B1(new_n538), .B2(new_n548), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n561), .A2(new_n563), .ZN(new_n564));
  XOR2_X1   g378(.A(KEYINPUT71), .B(KEYINPUT27), .Z(new_n565));
  NAND2_X1  g379(.A1(new_n364), .A2(G210), .ZN(new_n566));
  XNOR2_X1  g380(.A(new_n565), .B(new_n566), .ZN(new_n567));
  XNOR2_X1  g381(.A(KEYINPUT26), .B(G101), .ZN(new_n568));
  XNOR2_X1  g382(.A(new_n567), .B(new_n568), .ZN(new_n569));
  INV_X1    g383(.A(new_n569), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n564), .A2(new_n570), .ZN(new_n571));
  INV_X1    g385(.A(KEYINPUT31), .ZN(new_n572));
  OAI21_X1  g386(.A(KEYINPUT30), .B1(new_n546), .B2(new_n547), .ZN(new_n573));
  OAI21_X1  g387(.A(new_n208), .B1(new_n538), .B2(new_n573), .ZN(new_n574));
  AOI21_X1  g388(.A(KEYINPUT30), .B1(new_n557), .B2(new_n554), .ZN(new_n575));
  OAI211_X1 g389(.A(new_n549), .B(new_n559), .C1(new_n574), .C2(new_n575), .ZN(new_n576));
  OAI21_X1  g390(.A(new_n572), .B1(new_n576), .B2(new_n570), .ZN(new_n577));
  AND2_X1   g391(.A1(new_n549), .A2(new_n559), .ZN(new_n578));
  INV_X1    g392(.A(KEYINPUT30), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n555), .A2(new_n579), .ZN(new_n580));
  NAND3_X1  g394(.A1(new_n557), .A2(KEYINPUT30), .A3(new_n554), .ZN(new_n581));
  NAND3_X1  g395(.A1(new_n580), .A2(new_n208), .A3(new_n581), .ZN(new_n582));
  NAND4_X1  g396(.A1(new_n578), .A2(KEYINPUT31), .A3(new_n569), .A4(new_n582), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n577), .A2(new_n583), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n571), .A2(new_n584), .ZN(new_n585));
  NOR2_X1   g399(.A1(G472), .A2(G902), .ZN(new_n586));
  AOI21_X1  g400(.A(new_n533), .B1(new_n585), .B2(new_n586), .ZN(new_n587));
  INV_X1    g401(.A(KEYINPUT32), .ZN(new_n588));
  INV_X1    g402(.A(new_n586), .ZN(new_n589));
  AOI211_X1 g403(.A(new_n588), .B(new_n589), .C1(new_n571), .C2(new_n584), .ZN(new_n590));
  NOR2_X1   g404(.A1(new_n587), .A2(new_n590), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n576), .A2(new_n570), .ZN(new_n592));
  INV_X1    g406(.A(KEYINPUT29), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n563), .A2(new_n569), .ZN(new_n595));
  AOI21_X1  g409(.A(new_n595), .B1(new_n560), .B2(KEYINPUT28), .ZN(new_n596));
  OAI21_X1  g410(.A(KEYINPUT73), .B1(new_n594), .B2(new_n596), .ZN(new_n597));
  INV_X1    g411(.A(new_n596), .ZN(new_n598));
  INV_X1    g412(.A(KEYINPUT73), .ZN(new_n599));
  AOI21_X1  g413(.A(KEYINPUT29), .B1(new_n576), .B2(new_n570), .ZN(new_n600));
  NAND3_X1  g414(.A1(new_n598), .A2(new_n599), .A3(new_n600), .ZN(new_n601));
  INV_X1    g415(.A(KEYINPUT74), .ZN(new_n602));
  NAND3_X1  g416(.A1(new_n563), .A2(KEYINPUT29), .A3(new_n569), .ZN(new_n603));
  AOI21_X1  g417(.A(new_n603), .B1(KEYINPUT28), .B2(new_n560), .ZN(new_n604));
  OAI21_X1  g418(.A(new_n602), .B1(new_n604), .B2(G902), .ZN(new_n605));
  INV_X1    g419(.A(new_n603), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n561), .A2(new_n606), .ZN(new_n607));
  NAND3_X1  g421(.A1(new_n607), .A2(KEYINPUT74), .A3(new_n297), .ZN(new_n608));
  NAND4_X1  g422(.A1(new_n597), .A2(new_n601), .A3(new_n605), .A4(new_n608), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n609), .A2(G472), .ZN(new_n610));
  AOI21_X1  g424(.A(new_n532), .B1(new_n591), .B2(new_n610), .ZN(new_n611));
  INV_X1    g425(.A(new_n611), .ZN(new_n612));
  NOR2_X1   g426(.A1(new_n493), .A2(new_n612), .ZN(new_n613));
  XNOR2_X1  g427(.A(new_n613), .B(new_n201), .ZN(G3));
  AOI21_X1  g428(.A(G902), .B1(new_n571), .B2(new_n584), .ZN(new_n615));
  INV_X1    g429(.A(G472), .ZN(new_n616));
  AOI22_X1  g430(.A1(new_n564), .A2(new_n570), .B1(new_n577), .B2(new_n583), .ZN(new_n617));
  OAI22_X1  g431(.A1(new_n615), .A2(new_n616), .B1(new_n617), .B2(new_n589), .ZN(new_n618));
  NOR2_X1   g432(.A1(new_n618), .A2(new_n532), .ZN(new_n619));
  AND2_X1   g433(.A1(new_n619), .A2(new_n490), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n282), .A2(new_n292), .ZN(new_n621));
  INV_X1    g435(.A(new_n293), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  INV_X1    g437(.A(KEYINPUT94), .ZN(new_n624));
  NAND3_X1  g438(.A1(new_n282), .A2(new_n292), .A3(new_n293), .ZN(new_n625));
  NAND3_X1  g439(.A1(new_n623), .A2(new_n624), .A3(new_n625), .ZN(new_n626));
  NAND4_X1  g440(.A1(new_n282), .A2(new_n292), .A3(KEYINPUT94), .A4(new_n293), .ZN(new_n627));
  AND2_X1   g441(.A1(new_n627), .A2(new_n187), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n626), .A2(new_n628), .ZN(new_n629));
  INV_X1    g443(.A(new_n398), .ZN(new_n630));
  NAND2_X1  g444(.A1(G478), .A2(G902), .ZN(new_n631));
  OAI21_X1  g445(.A(new_n631), .B1(new_n336), .B2(G478), .ZN(new_n632));
  INV_X1    g446(.A(new_n335), .ZN(new_n633));
  INV_X1    g447(.A(KEYINPUT33), .ZN(new_n634));
  NAND3_X1  g448(.A1(new_n325), .A2(new_n330), .A3(new_n333), .ZN(new_n635));
  NAND3_X1  g449(.A1(new_n633), .A2(new_n634), .A3(new_n635), .ZN(new_n636));
  OAI21_X1  g450(.A(KEYINPUT33), .B1(new_n334), .B2(new_n335), .ZN(new_n637));
  AND2_X1   g451(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  AOI21_X1  g452(.A(new_n632), .B1(new_n638), .B2(G478), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n630), .A2(new_n639), .ZN(new_n640));
  NOR3_X1   g454(.A1(new_n629), .A2(new_n406), .A3(new_n640), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n620), .A2(new_n641), .ZN(new_n642));
  XOR2_X1   g456(.A(KEYINPUT34), .B(G104), .Z(new_n643));
  XNOR2_X1  g457(.A(new_n642), .B(new_n643), .ZN(G6));
  NAND2_X1  g458(.A1(new_n392), .A2(new_n394), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n397), .A2(G475), .ZN(new_n646));
  INV_X1    g460(.A(KEYINPUT95), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  NAND3_X1  g462(.A1(new_n397), .A2(KEYINPUT95), .A3(G475), .ZN(new_n649));
  NAND3_X1  g463(.A1(new_n645), .A2(new_n648), .A3(new_n649), .ZN(new_n650));
  NOR4_X1   g464(.A1(new_n629), .A2(new_n650), .A3(new_n406), .A4(new_n341), .ZN(new_n651));
  NAND2_X1  g465(.A1(new_n620), .A2(new_n651), .ZN(new_n652));
  XOR2_X1   g466(.A(KEYINPUT35), .B(G107), .Z(new_n653));
  XNOR2_X1  g467(.A(new_n652), .B(new_n653), .ZN(G9));
  NOR2_X1   g468(.A1(new_n519), .A2(KEYINPUT36), .ZN(new_n655));
  XNOR2_X1  g469(.A(new_n520), .B(new_n655), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n656), .A2(new_n530), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n528), .A2(new_n657), .ZN(new_n658));
  INV_X1    g472(.A(new_n658), .ZN(new_n659));
  NOR2_X1   g473(.A1(new_n659), .A2(new_n618), .ZN(new_n660));
  INV_X1    g474(.A(new_n660), .ZN(new_n661));
  NOR2_X1   g475(.A1(new_n493), .A2(new_n661), .ZN(new_n662));
  XNOR2_X1  g476(.A(new_n662), .B(KEYINPUT96), .ZN(new_n663));
  XOR2_X1   g477(.A(KEYINPUT37), .B(G110), .Z(new_n664));
  XNOR2_X1  g478(.A(new_n663), .B(new_n664), .ZN(G12));
  NAND3_X1  g479(.A1(new_n585), .A2(KEYINPUT32), .A3(new_n586), .ZN(new_n666));
  INV_X1    g480(.A(new_n533), .ZN(new_n667));
  OAI21_X1  g481(.A(new_n667), .B1(new_n617), .B2(new_n589), .ZN(new_n668));
  NAND3_X1  g482(.A1(new_n610), .A2(new_n666), .A3(new_n668), .ZN(new_n669));
  AOI21_X1  g483(.A(new_n629), .B1(new_n489), .B2(new_n477), .ZN(new_n670));
  INV_X1    g484(.A(G900), .ZN(new_n671));
  NAND2_X1  g485(.A1(new_n404), .A2(new_n671), .ZN(new_n672));
  INV_X1    g486(.A(new_n402), .ZN(new_n673));
  NAND2_X1  g487(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  XOR2_X1   g488(.A(new_n674), .B(KEYINPUT97), .Z(new_n675));
  INV_X1    g489(.A(new_n675), .ZN(new_n676));
  NOR3_X1   g490(.A1(new_n650), .A2(new_n341), .A3(new_n676), .ZN(new_n677));
  NAND4_X1  g491(.A1(new_n669), .A2(new_n670), .A3(new_n658), .A4(new_n677), .ZN(new_n678));
  XNOR2_X1  g492(.A(new_n678), .B(G128), .ZN(G30));
  XNOR2_X1  g493(.A(new_n675), .B(KEYINPUT39), .ZN(new_n680));
  NAND2_X1  g494(.A1(new_n490), .A2(new_n680), .ZN(new_n681));
  INV_X1    g495(.A(KEYINPUT40), .ZN(new_n682));
  XNOR2_X1  g496(.A(new_n681), .B(new_n682), .ZN(new_n683));
  INV_X1    g497(.A(new_n576), .ZN(new_n684));
  NOR2_X1   g498(.A1(new_n684), .A2(new_n570), .ZN(new_n685));
  OAI21_X1  g499(.A(new_n297), .B1(new_n560), .B2(new_n569), .ZN(new_n686));
  OAI21_X1  g500(.A(G472), .B1(new_n685), .B2(new_n686), .ZN(new_n687));
  NAND3_X1  g501(.A1(new_n668), .A2(new_n666), .A3(new_n687), .ZN(new_n688));
  INV_X1    g502(.A(new_n688), .ZN(new_n689));
  NAND2_X1  g503(.A1(new_n623), .A2(new_n625), .ZN(new_n690));
  INV_X1    g504(.A(KEYINPUT38), .ZN(new_n691));
  XNOR2_X1  g505(.A(new_n690), .B(new_n691), .ZN(new_n692));
  NAND2_X1  g506(.A1(new_n339), .A2(new_n340), .ZN(new_n693));
  NAND3_X1  g507(.A1(new_n630), .A2(new_n187), .A3(new_n693), .ZN(new_n694));
  NOR4_X1   g508(.A1(new_n689), .A2(new_n692), .A3(new_n658), .A4(new_n694), .ZN(new_n695));
  NAND2_X1  g509(.A1(new_n683), .A2(new_n695), .ZN(new_n696));
  NAND2_X1  g510(.A1(new_n696), .A2(KEYINPUT98), .ZN(new_n697));
  INV_X1    g511(.A(KEYINPUT98), .ZN(new_n698));
  NAND3_X1  g512(.A1(new_n683), .A2(new_n698), .A3(new_n695), .ZN(new_n699));
  NAND2_X1  g513(.A1(new_n697), .A2(new_n699), .ZN(new_n700));
  XNOR2_X1  g514(.A(new_n700), .B(new_n233), .ZN(G45));
  NOR2_X1   g515(.A1(new_n640), .A2(new_n676), .ZN(new_n702));
  NAND4_X1  g516(.A1(new_n669), .A2(new_n670), .A3(new_n658), .A4(new_n702), .ZN(new_n703));
  XNOR2_X1  g517(.A(KEYINPUT99), .B(G146), .ZN(new_n704));
  XNOR2_X1  g518(.A(new_n703), .B(new_n704), .ZN(G48));
  NAND2_X1  g519(.A1(new_n474), .A2(new_n475), .ZN(new_n706));
  NAND2_X1  g520(.A1(new_n706), .A2(new_n297), .ZN(new_n707));
  NAND2_X1  g521(.A1(new_n707), .A2(G469), .ZN(new_n708));
  NAND3_X1  g522(.A1(new_n708), .A2(new_n413), .A3(new_n482), .ZN(new_n709));
  INV_X1    g523(.A(new_n709), .ZN(new_n710));
  NAND2_X1  g524(.A1(new_n611), .A2(new_n710), .ZN(new_n711));
  INV_X1    g525(.A(new_n711), .ZN(new_n712));
  NAND2_X1  g526(.A1(new_n712), .A2(new_n641), .ZN(new_n713));
  XNOR2_X1  g527(.A(KEYINPUT41), .B(G113), .ZN(new_n714));
  XNOR2_X1  g528(.A(new_n713), .B(new_n714), .ZN(G15));
  NAND2_X1  g529(.A1(new_n712), .A2(new_n651), .ZN(new_n716));
  XOR2_X1   g530(.A(KEYINPUT100), .B(G116), .Z(new_n717));
  XNOR2_X1  g531(.A(new_n716), .B(new_n717), .ZN(G18));
  NOR3_X1   g532(.A1(new_n629), .A2(new_n408), .A3(new_n709), .ZN(new_n719));
  NAND3_X1  g533(.A1(new_n669), .A2(new_n658), .A3(new_n719), .ZN(new_n720));
  XNOR2_X1  g534(.A(new_n720), .B(G119), .ZN(G21));
  NAND4_X1  g535(.A1(new_n708), .A2(new_n413), .A3(new_n482), .A4(new_n407), .ZN(new_n722));
  NOR3_X1   g536(.A1(new_n618), .A2(new_n532), .A3(new_n722), .ZN(new_n723));
  NAND3_X1  g537(.A1(new_n630), .A2(KEYINPUT101), .A3(new_n693), .ZN(new_n724));
  INV_X1    g538(.A(KEYINPUT101), .ZN(new_n725));
  OAI21_X1  g539(.A(new_n725), .B1(new_n341), .B2(new_n398), .ZN(new_n726));
  AND4_X1   g540(.A1(new_n626), .A2(new_n724), .A3(new_n628), .A4(new_n726), .ZN(new_n727));
  NAND2_X1  g541(.A1(new_n723), .A2(new_n727), .ZN(new_n728));
  XNOR2_X1  g542(.A(new_n728), .B(G122), .ZN(G24));
  NOR2_X1   g543(.A1(new_n629), .A2(new_n709), .ZN(new_n730));
  NAND3_X1  g544(.A1(new_n660), .A2(new_n702), .A3(new_n730), .ZN(new_n731));
  XNOR2_X1  g545(.A(new_n731), .B(G125), .ZN(G27));
  INV_X1    g546(.A(KEYINPUT105), .ZN(new_n733));
  OAI21_X1  g547(.A(new_n588), .B1(new_n617), .B2(new_n589), .ZN(new_n734));
  NAND3_X1  g548(.A1(new_n610), .A2(new_n666), .A3(new_n734), .ZN(new_n735));
  INV_X1    g549(.A(new_n532), .ZN(new_n736));
  NAND2_X1  g550(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  INV_X1    g551(.A(new_n187), .ZN(new_n738));
  NOR2_X1   g552(.A1(new_n412), .A2(new_n738), .ZN(new_n739));
  NAND3_X1  g553(.A1(new_n623), .A2(new_n625), .A3(new_n739), .ZN(new_n740));
  NAND2_X1  g554(.A1(new_n458), .A2(new_n468), .ZN(new_n741));
  NAND2_X1  g555(.A1(new_n741), .A2(KEYINPUT103), .ZN(new_n742));
  INV_X1    g556(.A(KEYINPUT103), .ZN(new_n743));
  NAND2_X1  g557(.A1(new_n468), .A2(new_n743), .ZN(new_n744));
  NAND3_X1  g558(.A1(new_n742), .A2(new_n744), .A3(G469), .ZN(new_n745));
  XOR2_X1   g559(.A(new_n470), .B(KEYINPUT102), .Z(new_n746));
  INV_X1    g560(.A(new_n746), .ZN(new_n747));
  NOR2_X1   g561(.A1(new_n476), .A2(new_n747), .ZN(new_n748));
  AOI21_X1  g562(.A(new_n740), .B1(new_n745), .B2(new_n748), .ZN(new_n749));
  NAND3_X1  g563(.A1(new_n749), .A2(KEYINPUT42), .A3(new_n702), .ZN(new_n750));
  OAI21_X1  g564(.A(new_n733), .B1(new_n737), .B2(new_n750), .ZN(new_n751));
  INV_X1    g565(.A(new_n750), .ZN(new_n752));
  NAND4_X1  g566(.A1(new_n752), .A2(KEYINPUT105), .A3(new_n736), .A4(new_n735), .ZN(new_n753));
  NAND2_X1  g567(.A1(new_n751), .A2(new_n753), .ZN(new_n754));
  NAND4_X1  g568(.A1(new_n669), .A2(new_n736), .A3(new_n702), .A4(new_n749), .ZN(new_n755));
  INV_X1    g569(.A(KEYINPUT42), .ZN(new_n756));
  AND3_X1   g570(.A1(new_n755), .A2(KEYINPUT104), .A3(new_n756), .ZN(new_n757));
  AOI21_X1  g571(.A(KEYINPUT104), .B1(new_n755), .B2(new_n756), .ZN(new_n758));
  OAI21_X1  g572(.A(new_n754), .B1(new_n757), .B2(new_n758), .ZN(new_n759));
  XNOR2_X1  g573(.A(new_n759), .B(G131), .ZN(G33));
  NAND4_X1  g574(.A1(new_n669), .A2(new_n736), .A3(new_n677), .A4(new_n749), .ZN(new_n761));
  XNOR2_X1  g575(.A(new_n761), .B(G134), .ZN(G36));
  NAND3_X1  g576(.A1(new_n742), .A2(new_n744), .A3(KEYINPUT45), .ZN(new_n763));
  INV_X1    g577(.A(KEYINPUT106), .ZN(new_n764));
  OR2_X1    g578(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  NAND2_X1  g579(.A1(new_n763), .A2(new_n764), .ZN(new_n766));
  AND2_X1   g580(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  INV_X1    g581(.A(KEYINPUT45), .ZN(new_n768));
  AOI21_X1  g582(.A(new_n479), .B1(new_n741), .B2(new_n768), .ZN(new_n769));
  INV_X1    g583(.A(new_n769), .ZN(new_n770));
  OAI211_X1 g584(.A(KEYINPUT46), .B(new_n746), .C1(new_n767), .C2(new_n770), .ZN(new_n771));
  INV_X1    g585(.A(KEYINPUT46), .ZN(new_n772));
  AOI21_X1  g586(.A(new_n770), .B1(new_n765), .B2(new_n766), .ZN(new_n773));
  OAI21_X1  g587(.A(new_n772), .B1(new_n773), .B2(new_n747), .ZN(new_n774));
  NAND3_X1  g588(.A1(new_n771), .A2(new_n774), .A3(new_n482), .ZN(new_n775));
  AND3_X1   g589(.A1(new_n775), .A2(new_n413), .A3(new_n680), .ZN(new_n776));
  NAND2_X1  g590(.A1(new_n639), .A2(new_n398), .ZN(new_n777));
  XOR2_X1   g591(.A(new_n777), .B(KEYINPUT43), .Z(new_n778));
  NAND3_X1  g592(.A1(new_n778), .A2(new_n618), .A3(new_n658), .ZN(new_n779));
  INV_X1    g593(.A(KEYINPUT44), .ZN(new_n780));
  NAND2_X1  g594(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  NAND4_X1  g595(.A1(new_n778), .A2(KEYINPUT44), .A3(new_n618), .A4(new_n658), .ZN(new_n782));
  NOR2_X1   g596(.A1(new_n690), .A2(new_n738), .ZN(new_n783));
  NAND3_X1  g597(.A1(new_n781), .A2(new_n782), .A3(new_n783), .ZN(new_n784));
  INV_X1    g598(.A(KEYINPUT107), .ZN(new_n785));
  OR2_X1    g599(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n784), .A2(new_n785), .ZN(new_n787));
  NAND3_X1  g601(.A1(new_n776), .A2(new_n786), .A3(new_n787), .ZN(new_n788));
  XNOR2_X1  g602(.A(new_n788), .B(G137), .ZN(G39));
  NAND3_X1  g603(.A1(new_n702), .A2(new_n532), .A3(new_n783), .ZN(new_n790));
  NOR2_X1   g604(.A1(new_n669), .A2(new_n790), .ZN(new_n791));
  NAND3_X1  g605(.A1(new_n775), .A2(KEYINPUT47), .A3(new_n413), .ZN(new_n792));
  INV_X1    g606(.A(new_n792), .ZN(new_n793));
  AOI21_X1  g607(.A(KEYINPUT47), .B1(new_n775), .B2(new_n413), .ZN(new_n794));
  OAI21_X1  g608(.A(new_n791), .B1(new_n793), .B2(new_n794), .ZN(new_n795));
  XNOR2_X1  g609(.A(new_n795), .B(G140), .ZN(G42));
  NAND3_X1  g610(.A1(new_n619), .A2(new_n402), .A3(new_n778), .ZN(new_n797));
  INV_X1    g611(.A(new_n730), .ZN(new_n798));
  OAI211_X1 g612(.A(G952), .B(new_n261), .C1(new_n797), .C2(new_n798), .ZN(new_n799));
  INV_X1    g613(.A(new_n783), .ZN(new_n800));
  NOR3_X1   g614(.A1(new_n800), .A2(new_n673), .A3(new_n709), .ZN(new_n801));
  AND3_X1   g615(.A1(new_n801), .A2(new_n736), .A3(new_n689), .ZN(new_n802));
  INV_X1    g616(.A(new_n640), .ZN(new_n803));
  AOI21_X1  g617(.A(new_n799), .B1(new_n802), .B2(new_n803), .ZN(new_n804));
  NAND2_X1  g618(.A1(new_n801), .A2(new_n778), .ZN(new_n805));
  NOR2_X1   g619(.A1(new_n805), .A2(new_n737), .ZN(new_n806));
  XOR2_X1   g620(.A(new_n806), .B(KEYINPUT114), .Z(new_n807));
  XNOR2_X1  g621(.A(KEYINPUT115), .B(KEYINPUT48), .ZN(new_n808));
  OAI21_X1  g622(.A(new_n804), .B1(new_n807), .B2(new_n808), .ZN(new_n809));
  NOR2_X1   g623(.A1(KEYINPUT115), .A2(KEYINPUT48), .ZN(new_n810));
  AOI21_X1  g624(.A(new_n809), .B1(new_n807), .B2(new_n810), .ZN(new_n811));
  NAND3_X1  g625(.A1(new_n692), .A2(new_n710), .A3(new_n738), .ZN(new_n812));
  NOR2_X1   g626(.A1(new_n797), .A2(new_n812), .ZN(new_n813));
  XNOR2_X1  g627(.A(new_n813), .B(KEYINPUT50), .ZN(new_n814));
  INV_X1    g628(.A(KEYINPUT51), .ZN(new_n815));
  NOR2_X1   g629(.A1(new_n805), .A2(new_n661), .ZN(new_n816));
  NOR2_X1   g630(.A1(new_n630), .A2(new_n639), .ZN(new_n817));
  AOI21_X1  g631(.A(new_n816), .B1(new_n802), .B2(new_n817), .ZN(new_n818));
  NAND3_X1  g632(.A1(new_n814), .A2(new_n815), .A3(new_n818), .ZN(new_n819));
  NOR2_X1   g633(.A1(new_n793), .A2(new_n794), .ZN(new_n820));
  NAND2_X1  g634(.A1(new_n820), .A2(KEYINPUT112), .ZN(new_n821));
  NAND2_X1  g635(.A1(new_n775), .A2(new_n413), .ZN(new_n822));
  INV_X1    g636(.A(KEYINPUT47), .ZN(new_n823));
  NAND2_X1  g637(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  NAND2_X1  g638(.A1(new_n824), .A2(new_n792), .ZN(new_n825));
  INV_X1    g639(.A(KEYINPUT112), .ZN(new_n826));
  NAND2_X1  g640(.A1(new_n825), .A2(new_n826), .ZN(new_n827));
  AND2_X1   g641(.A1(new_n708), .A2(new_n482), .ZN(new_n828));
  NAND2_X1  g642(.A1(new_n828), .A2(new_n412), .ZN(new_n829));
  NAND3_X1  g643(.A1(new_n821), .A2(new_n827), .A3(new_n829), .ZN(new_n830));
  NOR2_X1   g644(.A1(new_n797), .A2(new_n800), .ZN(new_n831));
  XNOR2_X1  g645(.A(new_n831), .B(KEYINPUT111), .ZN(new_n832));
  AOI21_X1  g646(.A(new_n819), .B1(new_n830), .B2(new_n832), .ZN(new_n833));
  NAND2_X1  g647(.A1(new_n814), .A2(new_n818), .ZN(new_n834));
  XNOR2_X1  g648(.A(new_n834), .B(KEYINPUT113), .ZN(new_n835));
  NAND2_X1  g649(.A1(new_n820), .A2(new_n829), .ZN(new_n836));
  NAND2_X1  g650(.A1(new_n836), .A2(new_n832), .ZN(new_n837));
  AOI21_X1  g651(.A(new_n815), .B1(new_n835), .B2(new_n837), .ZN(new_n838));
  OAI21_X1  g652(.A(new_n811), .B1(new_n833), .B2(new_n838), .ZN(new_n839));
  AOI211_X1 g653(.A(new_n412), .B(new_n676), .C1(new_n745), .C2(new_n748), .ZN(new_n840));
  NAND4_X1  g654(.A1(new_n727), .A2(new_n840), .A3(new_n659), .A4(new_n688), .ZN(new_n841));
  NAND4_X1  g655(.A1(new_n678), .A2(new_n703), .A3(new_n731), .A4(new_n841), .ZN(new_n842));
  INV_X1    g656(.A(KEYINPUT52), .ZN(new_n843));
  XNOR2_X1  g657(.A(new_n842), .B(new_n843), .ZN(new_n844));
  NOR3_X1   g658(.A1(new_n650), .A2(new_n693), .A3(new_n676), .ZN(new_n845));
  AND2_X1   g659(.A1(new_n783), .A2(new_n845), .ZN(new_n846));
  NAND4_X1  g660(.A1(new_n669), .A2(new_n490), .A3(new_n658), .A4(new_n846), .ZN(new_n847));
  NAND3_X1  g661(.A1(new_n660), .A2(new_n702), .A3(new_n749), .ZN(new_n848));
  AND3_X1   g662(.A1(new_n761), .A2(new_n847), .A3(new_n848), .ZN(new_n849));
  NAND2_X1  g663(.A1(new_n341), .A2(new_n398), .ZN(new_n850));
  OAI21_X1  g664(.A(new_n850), .B1(new_n639), .B2(new_n398), .ZN(new_n851));
  NOR3_X1   g665(.A1(new_n851), .A2(new_n296), .A3(new_n406), .ZN(new_n852));
  NAND3_X1  g666(.A1(new_n619), .A2(new_n490), .A3(new_n852), .ZN(new_n853));
  AND3_X1   g667(.A1(new_n720), .A2(new_n728), .A3(new_n853), .ZN(new_n854));
  OAI211_X1 g668(.A(new_n492), .B(new_n486), .C1(new_n611), .C2(new_n660), .ZN(new_n855));
  OAI211_X1 g669(.A(new_n611), .B(new_n710), .C1(new_n641), .C2(new_n651), .ZN(new_n856));
  NAND4_X1  g670(.A1(new_n849), .A2(new_n854), .A3(new_n855), .A4(new_n856), .ZN(new_n857));
  INV_X1    g671(.A(new_n857), .ZN(new_n858));
  NAND3_X1  g672(.A1(new_n844), .A2(new_n858), .A3(new_n759), .ZN(new_n859));
  NAND2_X1  g673(.A1(new_n859), .A2(KEYINPUT53), .ZN(new_n860));
  AND3_X1   g674(.A1(new_n842), .A2(KEYINPUT110), .A3(new_n843), .ZN(new_n861));
  AOI21_X1  g675(.A(new_n843), .B1(new_n842), .B2(KEYINPUT110), .ZN(new_n862));
  OR2_X1    g676(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  INV_X1    g677(.A(KEYINPUT53), .ZN(new_n864));
  AOI21_X1  g678(.A(new_n659), .B1(new_n591), .B2(new_n610), .ZN(new_n865));
  AOI22_X1  g679(.A1(new_n865), .A2(new_n719), .B1(new_n723), .B2(new_n727), .ZN(new_n866));
  AND4_X1   g680(.A1(new_n853), .A2(new_n855), .A3(new_n856), .A4(new_n866), .ZN(new_n867));
  INV_X1    g681(.A(KEYINPUT109), .ZN(new_n868));
  NAND4_X1  g682(.A1(new_n759), .A2(new_n867), .A3(new_n868), .A4(new_n849), .ZN(new_n869));
  NAND3_X1  g683(.A1(new_n863), .A2(new_n864), .A3(new_n869), .ZN(new_n870));
  NAND2_X1  g684(.A1(new_n755), .A2(new_n756), .ZN(new_n871));
  INV_X1    g685(.A(KEYINPUT104), .ZN(new_n872));
  NAND2_X1  g686(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  NAND3_X1  g687(.A1(new_n755), .A2(KEYINPUT104), .A3(new_n756), .ZN(new_n874));
  AOI22_X1  g688(.A1(new_n873), .A2(new_n874), .B1(new_n751), .B2(new_n753), .ZN(new_n875));
  NOR2_X1   g689(.A1(new_n875), .A2(new_n857), .ZN(new_n876));
  NOR2_X1   g690(.A1(new_n876), .A2(new_n868), .ZN(new_n877));
  OAI211_X1 g691(.A(new_n860), .B(KEYINPUT54), .C1(new_n870), .C2(new_n877), .ZN(new_n878));
  NAND2_X1  g692(.A1(new_n859), .A2(new_n864), .ZN(new_n879));
  NAND3_X1  g693(.A1(new_n863), .A2(new_n876), .A3(KEYINPUT53), .ZN(new_n880));
  INV_X1    g694(.A(KEYINPUT54), .ZN(new_n881));
  NAND3_X1  g695(.A1(new_n879), .A2(new_n880), .A3(new_n881), .ZN(new_n882));
  NAND2_X1  g696(.A1(new_n878), .A2(new_n882), .ZN(new_n883));
  OAI22_X1  g697(.A1(new_n839), .A2(new_n883), .B1(G952), .B2(G953), .ZN(new_n884));
  INV_X1    g698(.A(new_n777), .ZN(new_n885));
  INV_X1    g699(.A(KEYINPUT49), .ZN(new_n886));
  OAI211_X1 g700(.A(new_n739), .B(new_n885), .C1(new_n828), .C2(new_n886), .ZN(new_n887));
  AOI21_X1  g701(.A(KEYINPUT108), .B1(new_n828), .B2(new_n886), .ZN(new_n888));
  NOR2_X1   g702(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  NAND3_X1  g703(.A1(new_n828), .A2(KEYINPUT108), .A3(new_n886), .ZN(new_n890));
  NAND4_X1  g704(.A1(new_n889), .A2(new_n692), .A3(new_n736), .A4(new_n890), .ZN(new_n891));
  OAI21_X1  g705(.A(new_n884), .B1(new_n688), .B2(new_n891), .ZN(G75));
  AOI21_X1  g706(.A(new_n297), .B1(new_n879), .B2(new_n880), .ZN(new_n893));
  NAND2_X1  g707(.A1(new_n893), .A2(G210), .ZN(new_n894));
  XNOR2_X1  g708(.A(new_n289), .B(KEYINPUT117), .ZN(new_n895));
  XNOR2_X1  g709(.A(new_n895), .B(KEYINPUT55), .ZN(new_n896));
  NAND2_X1  g710(.A1(new_n286), .A2(new_n291), .ZN(new_n897));
  XNOR2_X1  g711(.A(new_n897), .B(KEYINPUT116), .ZN(new_n898));
  XOR2_X1   g712(.A(new_n896), .B(new_n898), .Z(new_n899));
  INV_X1    g713(.A(KEYINPUT118), .ZN(new_n900));
  NOR2_X1   g714(.A1(new_n900), .A2(KEYINPUT56), .ZN(new_n901));
  AND3_X1   g715(.A1(new_n894), .A2(new_n899), .A3(new_n901), .ZN(new_n902));
  AOI21_X1  g716(.A(new_n899), .B1(new_n894), .B2(new_n901), .ZN(new_n903));
  NOR2_X1   g717(.A1(new_n261), .A2(G952), .ZN(new_n904));
  NOR3_X1   g718(.A1(new_n902), .A2(new_n903), .A3(new_n904), .ZN(G51));
  INV_X1    g719(.A(new_n882), .ZN(new_n906));
  AOI21_X1  g720(.A(new_n881), .B1(new_n879), .B2(new_n880), .ZN(new_n907));
  NOR2_X1   g721(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  XNOR2_X1  g722(.A(new_n746), .B(KEYINPUT57), .ZN(new_n909));
  OAI21_X1  g723(.A(new_n706), .B1(new_n908), .B2(new_n909), .ZN(new_n910));
  NAND2_X1  g724(.A1(new_n893), .A2(new_n773), .ZN(new_n911));
  AOI21_X1  g725(.A(new_n904), .B1(new_n910), .B2(new_n911), .ZN(G54));
  NAND3_X1  g726(.A1(new_n893), .A2(KEYINPUT58), .A3(G475), .ZN(new_n913));
  NOR2_X1   g727(.A1(new_n379), .A2(new_n388), .ZN(new_n914));
  AND2_X1   g728(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  NOR2_X1   g729(.A1(new_n913), .A2(new_n914), .ZN(new_n916));
  NOR3_X1   g730(.A1(new_n915), .A2(new_n916), .A3(new_n904), .ZN(G60));
  INV_X1    g731(.A(new_n904), .ZN(new_n918));
  XOR2_X1   g732(.A(new_n631), .B(KEYINPUT59), .Z(new_n919));
  AOI21_X1  g733(.A(new_n919), .B1(new_n878), .B2(new_n882), .ZN(new_n920));
  INV_X1    g734(.A(new_n638), .ZN(new_n921));
  OAI21_X1  g735(.A(new_n918), .B1(new_n920), .B2(new_n921), .ZN(new_n922));
  INV_X1    g736(.A(new_n907), .ZN(new_n923));
  NAND2_X1  g737(.A1(new_n923), .A2(new_n882), .ZN(new_n924));
  NOR2_X1   g738(.A1(new_n638), .A2(new_n919), .ZN(new_n925));
  NAND2_X1  g739(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  INV_X1    g740(.A(KEYINPUT119), .ZN(new_n927));
  NAND2_X1  g741(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  NAND3_X1  g742(.A1(new_n924), .A2(KEYINPUT119), .A3(new_n925), .ZN(new_n929));
  AOI21_X1  g743(.A(new_n922), .B1(new_n928), .B2(new_n929), .ZN(G63));
  INV_X1    g744(.A(KEYINPUT61), .ZN(new_n931));
  XNOR2_X1  g745(.A(KEYINPUT120), .B(KEYINPUT60), .ZN(new_n932));
  NOR2_X1   g746(.A1(new_n332), .A2(new_n297), .ZN(new_n933));
  XNOR2_X1  g747(.A(new_n932), .B(new_n933), .ZN(new_n934));
  AOI21_X1  g748(.A(KEYINPUT53), .B1(new_n876), .B2(new_n844), .ZN(new_n935));
  NAND4_X1  g749(.A1(new_n759), .A2(new_n867), .A3(KEYINPUT53), .A4(new_n849), .ZN(new_n936));
  NOR2_X1   g750(.A1(new_n861), .A2(new_n862), .ZN(new_n937));
  NOR2_X1   g751(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  OAI211_X1 g752(.A(new_n656), .B(new_n934), .C1(new_n935), .C2(new_n938), .ZN(new_n939));
  OAI21_X1  g753(.A(new_n934), .B1(new_n935), .B2(new_n938), .ZN(new_n940));
  INV_X1    g754(.A(new_n529), .ZN(new_n941));
  AOI21_X1  g755(.A(new_n904), .B1(new_n940), .B2(new_n941), .ZN(new_n942));
  INV_X1    g756(.A(KEYINPUT121), .ZN(new_n943));
  OAI21_X1  g757(.A(new_n939), .B1(new_n942), .B2(new_n943), .ZN(new_n944));
  INV_X1    g758(.A(new_n934), .ZN(new_n945));
  AOI21_X1  g759(.A(new_n945), .B1(new_n879), .B2(new_n880), .ZN(new_n946));
  OAI211_X1 g760(.A(new_n943), .B(new_n918), .C1(new_n946), .C2(new_n529), .ZN(new_n947));
  INV_X1    g761(.A(new_n947), .ZN(new_n948));
  OAI21_X1  g762(.A(new_n931), .B1(new_n944), .B2(new_n948), .ZN(new_n949));
  INV_X1    g763(.A(KEYINPUT122), .ZN(new_n950));
  OAI21_X1  g764(.A(new_n918), .B1(new_n946), .B2(new_n529), .ZN(new_n951));
  NAND2_X1  g765(.A1(new_n939), .A2(KEYINPUT61), .ZN(new_n952));
  OAI21_X1  g766(.A(new_n950), .B1(new_n951), .B2(new_n952), .ZN(new_n953));
  NAND4_X1  g767(.A1(new_n942), .A2(KEYINPUT122), .A3(KEYINPUT61), .A4(new_n939), .ZN(new_n954));
  NAND2_X1  g768(.A1(new_n953), .A2(new_n954), .ZN(new_n955));
  NAND2_X1  g769(.A1(new_n949), .A2(new_n955), .ZN(G66));
  INV_X1    g770(.A(new_n405), .ZN(new_n957));
  AOI21_X1  g771(.A(new_n261), .B1(new_n957), .B2(G224), .ZN(new_n958));
  NAND3_X1  g772(.A1(new_n854), .A2(new_n855), .A3(new_n856), .ZN(new_n959));
  AOI21_X1  g773(.A(new_n958), .B1(new_n959), .B2(new_n261), .ZN(new_n960));
  OAI21_X1  g774(.A(new_n898), .B1(G898), .B2(new_n261), .ZN(new_n961));
  XOR2_X1   g775(.A(new_n960), .B(new_n961), .Z(G69));
  NAND2_X1  g776(.A1(new_n580), .A2(new_n581), .ZN(new_n963));
  NAND2_X1  g777(.A1(new_n359), .A2(new_n360), .ZN(new_n964));
  XNOR2_X1  g778(.A(new_n963), .B(new_n964), .ZN(new_n965));
  INV_X1    g779(.A(new_n965), .ZN(new_n966));
  NAND3_X1  g780(.A1(new_n775), .A2(new_n413), .A3(new_n680), .ZN(new_n967));
  NOR2_X1   g781(.A1(new_n784), .A2(new_n785), .ZN(new_n968));
  NOR2_X1   g782(.A1(new_n967), .A2(new_n968), .ZN(new_n969));
  AOI22_X1  g783(.A1(new_n825), .A2(new_n791), .B1(new_n969), .B2(new_n787), .ZN(new_n970));
  NOR4_X1   g784(.A1(new_n612), .A2(new_n681), .A3(new_n800), .A4(new_n851), .ZN(new_n971));
  AND3_X1   g785(.A1(new_n678), .A2(new_n703), .A3(new_n731), .ZN(new_n972));
  NAND3_X1  g786(.A1(new_n697), .A2(new_n699), .A3(new_n972), .ZN(new_n973));
  AOI21_X1  g787(.A(new_n971), .B1(new_n973), .B2(KEYINPUT62), .ZN(new_n974));
  OAI211_X1 g788(.A(new_n970), .B(new_n974), .C1(KEYINPUT62), .C2(new_n973), .ZN(new_n975));
  AOI21_X1  g789(.A(new_n966), .B1(new_n975), .B2(new_n261), .ZN(new_n976));
  NOR2_X1   g790(.A1(new_n261), .A2(G900), .ZN(new_n977));
  XNOR2_X1  g791(.A(new_n977), .B(KEYINPUT124), .ZN(new_n978));
  NAND2_X1  g792(.A1(new_n972), .A2(new_n761), .ZN(new_n979));
  NAND3_X1  g793(.A1(new_n735), .A2(new_n736), .A3(new_n727), .ZN(new_n980));
  INV_X1    g794(.A(new_n980), .ZN(new_n981));
  AOI21_X1  g795(.A(new_n979), .B1(new_n776), .B2(new_n981), .ZN(new_n982));
  NAND4_X1  g796(.A1(new_n795), .A2(new_n982), .A3(new_n759), .A4(new_n788), .ZN(new_n983));
  AOI21_X1  g797(.A(new_n978), .B1(new_n983), .B2(new_n261), .ZN(new_n984));
  NOR2_X1   g798(.A1(new_n984), .A2(new_n965), .ZN(new_n985));
  NOR2_X1   g799(.A1(new_n976), .A2(new_n985), .ZN(new_n986));
  INV_X1    g800(.A(KEYINPUT123), .ZN(new_n987));
  OAI21_X1  g801(.A(new_n987), .B1(new_n984), .B2(new_n965), .ZN(new_n988));
  AOI21_X1  g802(.A(new_n261), .B1(G227), .B2(G900), .ZN(new_n989));
  INV_X1    g803(.A(new_n989), .ZN(new_n990));
  NAND2_X1  g804(.A1(new_n988), .A2(new_n990), .ZN(new_n991));
  NAND2_X1  g805(.A1(new_n986), .A2(new_n991), .ZN(new_n992));
  OAI211_X1 g806(.A(new_n990), .B(new_n988), .C1(new_n976), .C2(new_n985), .ZN(new_n993));
  AND2_X1   g807(.A1(new_n992), .A2(new_n993), .ZN(G72));
  NAND2_X1  g808(.A1(G472), .A2(G902), .ZN(new_n995));
  XOR2_X1   g809(.A(new_n995), .B(KEYINPUT63), .Z(new_n996));
  OAI21_X1  g810(.A(new_n996), .B1(new_n975), .B2(new_n959), .ZN(new_n997));
  NAND2_X1  g811(.A1(new_n997), .A2(new_n685), .ZN(new_n998));
  AOI21_X1  g812(.A(KEYINPUT127), .B1(new_n684), .B2(new_n569), .ZN(new_n999));
  XOR2_X1   g813(.A(new_n999), .B(new_n592), .Z(new_n1000));
  AND2_X1   g814(.A1(new_n1000), .A2(new_n996), .ZN(new_n1001));
  OAI211_X1 g815(.A(new_n860), .B(new_n1001), .C1(new_n870), .C2(new_n877), .ZN(new_n1002));
  NAND2_X1  g816(.A1(new_n998), .A2(new_n1002), .ZN(new_n1003));
  INV_X1    g817(.A(KEYINPUT125), .ZN(new_n1004));
  OAI211_X1 g818(.A(new_n1004), .B(new_n996), .C1(new_n983), .C2(new_n959), .ZN(new_n1005));
  NOR2_X1   g819(.A1(new_n576), .A2(new_n569), .ZN(new_n1006));
  NAND2_X1  g820(.A1(new_n1005), .A2(new_n1006), .ZN(new_n1007));
  NOR2_X1   g821(.A1(new_n967), .A2(new_n980), .ZN(new_n1008));
  NOR3_X1   g822(.A1(new_n1008), .A2(new_n875), .A3(new_n979), .ZN(new_n1009));
  NAND3_X1  g823(.A1(new_n970), .A2(new_n867), .A3(new_n1009), .ZN(new_n1010));
  AOI21_X1  g824(.A(new_n1004), .B1(new_n1010), .B2(new_n996), .ZN(new_n1011));
  OAI21_X1  g825(.A(new_n918), .B1(new_n1007), .B2(new_n1011), .ZN(new_n1012));
  INV_X1    g826(.A(KEYINPUT126), .ZN(new_n1013));
  NAND2_X1  g827(.A1(new_n1012), .A2(new_n1013), .ZN(new_n1014));
  OAI211_X1 g828(.A(KEYINPUT126), .B(new_n918), .C1(new_n1007), .C2(new_n1011), .ZN(new_n1015));
  AOI21_X1  g829(.A(new_n1003), .B1(new_n1014), .B2(new_n1015), .ZN(G57));
endmodule


