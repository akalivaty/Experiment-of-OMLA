//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 0 0 1 0 0 0 1 1 0 1 1 1 0 1 1 0 1 0 1 0 1 0 1 0 1 1 1 1 1 0 1 1 0 0 1 1 0 1 0 0 0 0 0 1 1 0 1 0 1 0 1 1 1 1 0 0 0 1 0 1 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:35:15 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n205, new_n206, new_n207, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n252, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1113, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1261, new_n1262, new_n1263, new_n1264, new_n1265,
    new_n1266, new_n1267, new_n1268, new_n1269, new_n1270, new_n1271,
    new_n1273, new_n1274, new_n1275, new_n1276, new_n1277, new_n1278,
    new_n1279, new_n1281, new_n1282, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1350, new_n1351, new_n1352, new_n1353,
    new_n1354, new_n1355, new_n1356;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  INV_X1    g0004(.A(G97), .ZN(new_n205));
  INV_X1    g0005(.A(G107), .ZN(new_n206));
  NAND2_X1  g0006(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  NAND2_X1  g0007(.A1(new_n207), .A2(G87), .ZN(G355));
  INV_X1    g0008(.A(G1), .ZN(new_n209));
  INV_X1    g0009(.A(G20), .ZN(new_n210));
  NOR2_X1   g0010(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  INV_X1    g0011(.A(new_n211), .ZN(new_n212));
  NOR2_X1   g0012(.A1(new_n212), .A2(G13), .ZN(new_n213));
  OAI211_X1 g0013(.A(new_n213), .B(G250), .C1(G257), .C2(G264), .ZN(new_n214));
  XNOR2_X1  g0014(.A(new_n214), .B(KEYINPUT0), .ZN(new_n215));
  INV_X1    g0015(.A(new_n201), .ZN(new_n216));
  NAND2_X1  g0016(.A1(new_n216), .A2(G50), .ZN(new_n217));
  INV_X1    g0017(.A(new_n217), .ZN(new_n218));
  NAND2_X1  g0018(.A1(G1), .A2(G13), .ZN(new_n219));
  NOR2_X1   g0019(.A1(new_n219), .A2(new_n210), .ZN(new_n220));
  NAND2_X1  g0020(.A1(new_n218), .A2(new_n220), .ZN(new_n221));
  AOI22_X1  g0021(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n222));
  INV_X1    g0022(.A(G68), .ZN(new_n223));
  INV_X1    g0023(.A(G238), .ZN(new_n224));
  INV_X1    g0024(.A(G87), .ZN(new_n225));
  INV_X1    g0025(.A(G250), .ZN(new_n226));
  OAI221_X1 g0026(.A(new_n222), .B1(new_n223), .B2(new_n224), .C1(new_n225), .C2(new_n226), .ZN(new_n227));
  AOI22_X1  g0027(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n228));
  INV_X1    g0028(.A(G77), .ZN(new_n229));
  INV_X1    g0029(.A(G244), .ZN(new_n230));
  INV_X1    g0030(.A(G264), .ZN(new_n231));
  OAI221_X1 g0031(.A(new_n228), .B1(new_n229), .B2(new_n230), .C1(new_n206), .C2(new_n231), .ZN(new_n232));
  OAI21_X1  g0032(.A(new_n212), .B1(new_n227), .B2(new_n232), .ZN(new_n233));
  OAI211_X1 g0033(.A(new_n215), .B(new_n221), .C1(KEYINPUT1), .C2(new_n233), .ZN(new_n234));
  AOI21_X1  g0034(.A(new_n234), .B1(KEYINPUT1), .B2(new_n233), .ZN(G361));
  XNOR2_X1  g0035(.A(G238), .B(G244), .ZN(new_n236));
  INV_X1    g0036(.A(G232), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XOR2_X1   g0038(.A(KEYINPUT2), .B(G226), .Z(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XOR2_X1   g0040(.A(G264), .B(G270), .Z(new_n241));
  XNOR2_X1  g0041(.A(G250), .B(G257), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n240), .B(new_n243), .ZN(G358));
  XOR2_X1   g0044(.A(G87), .B(G97), .Z(new_n245));
  XNOR2_X1  g0045(.A(new_n245), .B(KEYINPUT64), .ZN(new_n246));
  XNOR2_X1  g0046(.A(G107), .B(G116), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n246), .B(new_n247), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n248), .B(KEYINPUT65), .ZN(new_n249));
  XNOR2_X1  g0049(.A(G50), .B(G68), .ZN(new_n250));
  XNOR2_X1  g0050(.A(G58), .B(G77), .ZN(new_n251));
  XNOR2_X1  g0051(.A(new_n250), .B(new_n251), .ZN(new_n252));
  XNOR2_X1  g0052(.A(new_n249), .B(new_n252), .ZN(G351));
  NAND3_X1  g0053(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n254));
  NAND2_X1  g0054(.A1(new_n254), .A2(new_n219), .ZN(new_n255));
  INV_X1    g0055(.A(new_n255), .ZN(new_n256));
  XNOR2_X1  g0056(.A(KEYINPUT8), .B(G58), .ZN(new_n257));
  INV_X1    g0057(.A(new_n257), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n210), .A2(G33), .ZN(new_n259));
  INV_X1    g0059(.A(new_n259), .ZN(new_n260));
  NOR2_X1   g0060(.A1(G20), .A2(G33), .ZN(new_n261));
  AOI22_X1  g0061(.A1(new_n258), .A2(new_n260), .B1(G150), .B2(new_n261), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n203), .A2(G20), .ZN(new_n263));
  AOI21_X1  g0063(.A(new_n256), .B1(new_n262), .B2(new_n263), .ZN(new_n264));
  NAND3_X1  g0064(.A1(new_n209), .A2(G13), .A3(G20), .ZN(new_n265));
  INV_X1    g0065(.A(new_n265), .ZN(new_n266));
  NOR2_X1   g0066(.A1(new_n266), .A2(new_n255), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n209), .A2(G20), .ZN(new_n268));
  NAND3_X1  g0068(.A1(new_n267), .A2(G50), .A3(new_n268), .ZN(new_n269));
  OAI21_X1  g0069(.A(new_n269), .B1(G50), .B2(new_n265), .ZN(new_n270));
  NOR2_X1   g0070(.A1(new_n264), .A2(new_n270), .ZN(new_n271));
  XOR2_X1   g0071(.A(new_n271), .B(KEYINPUT9), .Z(new_n272));
  INV_X1    g0072(.A(G33), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n273), .A2(KEYINPUT3), .ZN(new_n274));
  INV_X1    g0074(.A(KEYINPUT3), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n275), .A2(G33), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n274), .A2(new_n276), .ZN(new_n277));
  INV_X1    g0077(.A(G1698), .ZN(new_n278));
  NOR2_X1   g0078(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  AOI22_X1  g0079(.A1(new_n279), .A2(G223), .B1(G77), .B2(new_n277), .ZN(new_n280));
  NOR2_X1   g0080(.A1(new_n277), .A2(G1698), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n281), .A2(G222), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n280), .A2(new_n282), .ZN(new_n283));
  AOI21_X1  g0083(.A(new_n219), .B1(G33), .B2(G41), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  INV_X1    g0085(.A(new_n284), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n286), .A2(G274), .ZN(new_n287));
  INV_X1    g0087(.A(G41), .ZN(new_n288));
  INV_X1    g0088(.A(G45), .ZN(new_n289));
  AOI21_X1  g0089(.A(G1), .B1(new_n288), .B2(new_n289), .ZN(new_n290));
  INV_X1    g0090(.A(new_n290), .ZN(new_n291));
  NOR2_X1   g0091(.A1(new_n287), .A2(new_n291), .ZN(new_n292));
  NOR2_X1   g0092(.A1(new_n284), .A2(new_n290), .ZN(new_n293));
  AOI21_X1  g0093(.A(new_n292), .B1(G226), .B2(new_n293), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n285), .A2(new_n294), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n295), .A2(G200), .ZN(new_n296));
  INV_X1    g0096(.A(G190), .ZN(new_n297));
  OAI211_X1 g0097(.A(new_n272), .B(new_n296), .C1(new_n297), .C2(new_n295), .ZN(new_n298));
  XNOR2_X1  g0098(.A(new_n298), .B(KEYINPUT10), .ZN(new_n299));
  INV_X1    g0099(.A(G169), .ZN(new_n300));
  AOI21_X1  g0100(.A(new_n271), .B1(new_n295), .B2(new_n300), .ZN(new_n301));
  OR2_X1    g0101(.A1(new_n301), .A2(KEYINPUT66), .ZN(new_n302));
  INV_X1    g0102(.A(G179), .ZN(new_n303));
  NAND3_X1  g0103(.A1(new_n285), .A2(new_n294), .A3(new_n303), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n301), .A2(KEYINPUT66), .ZN(new_n305));
  NAND3_X1  g0105(.A1(new_n302), .A2(new_n304), .A3(new_n305), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n299), .A2(new_n306), .ZN(new_n307));
  INV_X1    g0107(.A(new_n307), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n266), .A2(new_n223), .ZN(new_n309));
  XNOR2_X1  g0109(.A(new_n309), .B(KEYINPUT12), .ZN(new_n310));
  AOI22_X1  g0110(.A1(new_n261), .A2(G50), .B1(G20), .B2(new_n223), .ZN(new_n311));
  OAI21_X1  g0111(.A(new_n311), .B1(new_n229), .B2(new_n259), .ZN(new_n312));
  NAND3_X1  g0112(.A1(new_n312), .A2(KEYINPUT11), .A3(new_n255), .ZN(new_n313));
  NAND3_X1  g0113(.A1(new_n267), .A2(G68), .A3(new_n268), .ZN(new_n314));
  NAND3_X1  g0114(.A1(new_n310), .A2(new_n313), .A3(new_n314), .ZN(new_n315));
  AOI21_X1  g0115(.A(KEYINPUT11), .B1(new_n312), .B2(new_n255), .ZN(new_n316));
  NOR2_X1   g0116(.A1(new_n315), .A2(new_n316), .ZN(new_n317));
  INV_X1    g0117(.A(new_n317), .ZN(new_n318));
  AND2_X1   g0118(.A1(new_n286), .A2(G274), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n319), .A2(new_n290), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n286), .A2(new_n291), .ZN(new_n321));
  OAI21_X1  g0121(.A(new_n320), .B1(new_n224), .B2(new_n321), .ZN(new_n322));
  NAND4_X1  g0122(.A1(new_n274), .A2(new_n276), .A3(G232), .A4(G1698), .ZN(new_n323));
  XNOR2_X1  g0123(.A(new_n323), .B(KEYINPUT68), .ZN(new_n324));
  NOR2_X1   g0124(.A1(new_n273), .A2(new_n205), .ZN(new_n325));
  AOI21_X1  g0125(.A(new_n325), .B1(new_n281), .B2(G226), .ZN(new_n326));
  AOI21_X1  g0126(.A(new_n286), .B1(new_n324), .B2(new_n326), .ZN(new_n327));
  OR3_X1    g0127(.A1(new_n322), .A2(new_n327), .A3(KEYINPUT13), .ZN(new_n328));
  OAI21_X1  g0128(.A(KEYINPUT13), .B1(new_n322), .B2(new_n327), .ZN(new_n329));
  NAND3_X1  g0129(.A1(new_n328), .A2(G179), .A3(new_n329), .ZN(new_n330));
  NOR2_X1   g0130(.A1(new_n300), .A2(KEYINPUT69), .ZN(new_n331));
  INV_X1    g0131(.A(new_n331), .ZN(new_n332));
  AOI21_X1  g0132(.A(new_n332), .B1(new_n328), .B2(new_n329), .ZN(new_n333));
  INV_X1    g0133(.A(KEYINPUT14), .ZN(new_n334));
  OAI21_X1  g0134(.A(new_n330), .B1(new_n333), .B2(new_n334), .ZN(new_n335));
  AOI211_X1 g0135(.A(KEYINPUT14), .B(new_n332), .C1(new_n328), .C2(new_n329), .ZN(new_n336));
  OAI21_X1  g0136(.A(new_n318), .B1(new_n335), .B2(new_n336), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n328), .A2(new_n329), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n338), .A2(G200), .ZN(new_n339));
  OAI211_X1 g0139(.A(new_n339), .B(new_n317), .C1(new_n297), .C2(new_n338), .ZN(new_n340));
  AOI22_X1  g0140(.A1(new_n258), .A2(new_n261), .B1(G20), .B2(G77), .ZN(new_n341));
  XNOR2_X1  g0141(.A(KEYINPUT15), .B(G87), .ZN(new_n342));
  INV_X1    g0142(.A(new_n342), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n343), .A2(new_n260), .ZN(new_n344));
  AOI21_X1  g0144(.A(new_n256), .B1(new_n341), .B2(new_n344), .ZN(new_n345));
  NAND3_X1  g0145(.A1(new_n267), .A2(G77), .A3(new_n268), .ZN(new_n346));
  OAI21_X1  g0146(.A(new_n346), .B1(G77), .B2(new_n265), .ZN(new_n347));
  NOR2_X1   g0147(.A1(new_n345), .A2(new_n347), .ZN(new_n348));
  INV_X1    g0148(.A(new_n348), .ZN(new_n349));
  OAI21_X1  g0149(.A(new_n320), .B1(new_n230), .B2(new_n321), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n281), .A2(G232), .ZN(new_n351));
  INV_X1    g0151(.A(new_n277), .ZN(new_n352));
  NAND3_X1  g0152(.A1(new_n352), .A2(G238), .A3(G1698), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n277), .A2(G107), .ZN(new_n354));
  NAND3_X1  g0154(.A1(new_n351), .A2(new_n353), .A3(new_n354), .ZN(new_n355));
  AOI21_X1  g0155(.A(new_n286), .B1(new_n355), .B2(KEYINPUT67), .ZN(new_n356));
  INV_X1    g0156(.A(KEYINPUT67), .ZN(new_n357));
  NAND4_X1  g0157(.A1(new_n351), .A2(new_n353), .A3(new_n357), .A4(new_n354), .ZN(new_n358));
  AOI21_X1  g0158(.A(new_n350), .B1(new_n356), .B2(new_n358), .ZN(new_n359));
  OAI21_X1  g0159(.A(new_n349), .B1(new_n359), .B2(G169), .ZN(new_n360));
  AOI21_X1  g0160(.A(new_n360), .B1(new_n303), .B2(new_n359), .ZN(new_n361));
  AND2_X1   g0161(.A1(new_n356), .A2(new_n358), .ZN(new_n362));
  OAI21_X1  g0162(.A(G200), .B1(new_n362), .B2(new_n350), .ZN(new_n363));
  AOI21_X1  g0163(.A(new_n349), .B1(new_n359), .B2(G190), .ZN(new_n364));
  AOI21_X1  g0164(.A(new_n361), .B1(new_n363), .B2(new_n364), .ZN(new_n365));
  NAND4_X1  g0165(.A1(new_n308), .A2(new_n337), .A3(new_n340), .A4(new_n365), .ZN(new_n366));
  NAND3_X1  g0166(.A1(new_n267), .A2(new_n258), .A3(new_n268), .ZN(new_n367));
  OAI21_X1  g0167(.A(new_n367), .B1(new_n265), .B2(new_n258), .ZN(new_n368));
  INV_X1    g0168(.A(new_n368), .ZN(new_n369));
  INV_X1    g0169(.A(new_n276), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n275), .A2(KEYINPUT70), .ZN(new_n371));
  INV_X1    g0171(.A(KEYINPUT70), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n372), .A2(KEYINPUT3), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n371), .A2(new_n373), .ZN(new_n374));
  AOI21_X1  g0174(.A(new_n370), .B1(new_n374), .B2(new_n273), .ZN(new_n375));
  INV_X1    g0175(.A(KEYINPUT7), .ZN(new_n376));
  NOR2_X1   g0176(.A1(new_n376), .A2(G20), .ZN(new_n377));
  INV_X1    g0177(.A(new_n377), .ZN(new_n378));
  OAI21_X1  g0178(.A(KEYINPUT72), .B1(new_n375), .B2(new_n378), .ZN(new_n379));
  XNOR2_X1  g0179(.A(KEYINPUT70), .B(KEYINPUT3), .ZN(new_n380));
  OAI21_X1  g0180(.A(new_n276), .B1(new_n380), .B2(G33), .ZN(new_n381));
  INV_X1    g0181(.A(KEYINPUT72), .ZN(new_n382));
  NAND3_X1  g0182(.A1(new_n381), .A2(new_n382), .A3(new_n377), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n379), .A2(new_n383), .ZN(new_n384));
  AOI21_X1  g0184(.A(KEYINPUT7), .B1(new_n277), .B2(new_n210), .ZN(new_n385));
  INV_X1    g0185(.A(new_n385), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n384), .A2(new_n386), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n387), .A2(G68), .ZN(new_n388));
  NAND2_X1  g0188(.A1(G58), .A2(G68), .ZN(new_n389));
  AOI21_X1  g0189(.A(new_n210), .B1(new_n216), .B2(new_n389), .ZN(new_n390));
  AOI21_X1  g0190(.A(new_n390), .B1(G159), .B2(new_n261), .ZN(new_n391));
  AOI21_X1  g0191(.A(KEYINPUT16), .B1(new_n388), .B2(new_n391), .ZN(new_n392));
  NAND3_X1  g0192(.A1(new_n371), .A2(new_n373), .A3(G33), .ZN(new_n393));
  INV_X1    g0193(.A(KEYINPUT71), .ZN(new_n394));
  OAI21_X1  g0194(.A(new_n394), .B1(new_n275), .B2(G33), .ZN(new_n395));
  INV_X1    g0195(.A(new_n395), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n393), .A2(new_n396), .ZN(new_n397));
  NAND4_X1  g0197(.A1(new_n371), .A2(new_n373), .A3(KEYINPUT71), .A4(G33), .ZN(new_n398));
  NAND3_X1  g0198(.A1(new_n397), .A2(new_n210), .A3(new_n398), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n399), .A2(KEYINPUT7), .ZN(new_n400));
  NAND4_X1  g0200(.A1(new_n397), .A2(new_n376), .A3(new_n210), .A4(new_n398), .ZN(new_n401));
  NAND3_X1  g0201(.A1(new_n400), .A2(G68), .A3(new_n401), .ZN(new_n402));
  NAND3_X1  g0202(.A1(new_n402), .A2(KEYINPUT16), .A3(new_n391), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n403), .A2(new_n255), .ZN(new_n404));
  OAI21_X1  g0204(.A(new_n369), .B1(new_n392), .B2(new_n404), .ZN(new_n405));
  OAI21_X1  g0205(.A(KEYINPUT73), .B1(new_n321), .B2(new_n237), .ZN(new_n406));
  INV_X1    g0206(.A(KEYINPUT73), .ZN(new_n407));
  NAND3_X1  g0207(.A1(new_n293), .A2(new_n407), .A3(G232), .ZN(new_n408));
  AOI21_X1  g0208(.A(new_n292), .B1(new_n406), .B2(new_n408), .ZN(new_n409));
  OR2_X1    g0209(.A1(G223), .A2(G1698), .ZN(new_n410));
  OAI21_X1  g0210(.A(new_n410), .B1(G226), .B2(new_n278), .ZN(new_n411));
  AOI21_X1  g0211(.A(new_n411), .B1(new_n397), .B2(new_n398), .ZN(new_n412));
  NOR2_X1   g0212(.A1(new_n273), .A2(new_n225), .ZN(new_n413));
  OAI21_X1  g0213(.A(new_n284), .B1(new_n412), .B2(new_n413), .ZN(new_n414));
  AOI21_X1  g0214(.A(new_n300), .B1(new_n409), .B2(new_n414), .ZN(new_n415));
  AND2_X1   g0215(.A1(new_n409), .A2(new_n414), .ZN(new_n416));
  AOI21_X1  g0216(.A(new_n415), .B1(G179), .B2(new_n416), .ZN(new_n417));
  INV_X1    g0217(.A(new_n417), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n405), .A2(new_n418), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n419), .A2(KEYINPUT18), .ZN(new_n420));
  AOI21_X1  g0220(.A(new_n385), .B1(new_n379), .B2(new_n383), .ZN(new_n421));
  OAI21_X1  g0221(.A(new_n391), .B1(new_n421), .B2(new_n223), .ZN(new_n422));
  INV_X1    g0222(.A(KEYINPUT16), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  NAND3_X1  g0224(.A1(new_n424), .A2(new_n255), .A3(new_n403), .ZN(new_n425));
  AOI21_X1  g0225(.A(new_n417), .B1(new_n425), .B2(new_n369), .ZN(new_n426));
  INV_X1    g0226(.A(KEYINPUT18), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n426), .A2(new_n427), .ZN(new_n428));
  INV_X1    g0228(.A(G200), .ZN(new_n429));
  AOI21_X1  g0229(.A(new_n429), .B1(new_n409), .B2(new_n414), .ZN(new_n430));
  AND2_X1   g0230(.A1(new_n297), .A2(KEYINPUT74), .ZN(new_n431));
  NOR2_X1   g0231(.A1(new_n297), .A2(KEYINPUT74), .ZN(new_n432));
  NOR2_X1   g0232(.A1(new_n431), .A2(new_n432), .ZN(new_n433));
  INV_X1    g0233(.A(new_n433), .ZN(new_n434));
  AOI21_X1  g0234(.A(new_n430), .B1(new_n416), .B2(new_n434), .ZN(new_n435));
  NAND3_X1  g0235(.A1(new_n425), .A2(new_n435), .A3(new_n369), .ZN(new_n436));
  INV_X1    g0236(.A(KEYINPUT17), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n436), .A2(new_n437), .ZN(new_n438));
  NAND4_X1  g0238(.A1(new_n425), .A2(new_n435), .A3(KEYINPUT17), .A4(new_n369), .ZN(new_n439));
  NAND4_X1  g0239(.A1(new_n420), .A2(new_n428), .A3(new_n438), .A4(new_n439), .ZN(new_n440));
  NOR2_X1   g0240(.A1(new_n366), .A2(new_n440), .ZN(new_n441));
  INV_X1    g0241(.A(new_n441), .ZN(new_n442));
  NOR4_X1   g0242(.A1(new_n277), .A2(KEYINPUT22), .A3(G20), .A4(new_n225), .ZN(new_n443));
  INV_X1    g0243(.A(new_n443), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n397), .A2(new_n398), .ZN(new_n445));
  NAND4_X1  g0245(.A1(new_n445), .A2(KEYINPUT79), .A3(new_n210), .A4(G87), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n446), .A2(KEYINPUT22), .ZN(new_n447));
  AOI21_X1  g0247(.A(G20), .B1(new_n397), .B2(new_n398), .ZN(new_n448));
  AOI21_X1  g0248(.A(KEYINPUT79), .B1(new_n448), .B2(G87), .ZN(new_n449));
  OAI21_X1  g0249(.A(new_n444), .B1(new_n447), .B2(new_n449), .ZN(new_n450));
  INV_X1    g0250(.A(KEYINPUT24), .ZN(new_n451));
  OR3_X1    g0251(.A1(new_n210), .A2(KEYINPUT23), .A3(G107), .ZN(new_n452));
  NAND2_X1  g0252(.A1(G33), .A2(G116), .ZN(new_n453));
  OAI21_X1  g0253(.A(KEYINPUT23), .B1(new_n210), .B2(G107), .ZN(new_n454));
  INV_X1    g0254(.A(KEYINPUT80), .ZN(new_n455));
  OAI221_X1 g0255(.A(new_n452), .B1(G20), .B2(new_n453), .C1(new_n454), .C2(new_n455), .ZN(new_n456));
  AND2_X1   g0256(.A1(new_n454), .A2(new_n455), .ZN(new_n457));
  NOR2_X1   g0257(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  AND3_X1   g0258(.A1(new_n450), .A2(new_n451), .A3(new_n458), .ZN(new_n459));
  AOI21_X1  g0259(.A(new_n451), .B1(new_n450), .B2(new_n458), .ZN(new_n460));
  OAI21_X1  g0260(.A(new_n255), .B1(new_n459), .B2(new_n460), .ZN(new_n461));
  INV_X1    g0261(.A(KEYINPUT81), .ZN(new_n462));
  OAI21_X1  g0262(.A(new_n206), .B1(new_n462), .B2(KEYINPUT25), .ZN(new_n463));
  NOR2_X1   g0263(.A1(new_n463), .A2(new_n265), .ZN(new_n464));
  AOI21_X1  g0264(.A(new_n464), .B1(new_n462), .B2(KEYINPUT25), .ZN(new_n465));
  INV_X1    g0265(.A(new_n465), .ZN(new_n466));
  NAND3_X1  g0266(.A1(new_n464), .A2(new_n462), .A3(KEYINPUT25), .ZN(new_n467));
  NOR2_X1   g0267(.A1(new_n273), .A2(G1), .ZN(new_n468));
  NOR3_X1   g0268(.A1(new_n266), .A2(new_n255), .A3(new_n468), .ZN(new_n469));
  AOI22_X1  g0269(.A1(new_n466), .A2(new_n467), .B1(G107), .B2(new_n469), .ZN(new_n470));
  AOI21_X1  g0270(.A(new_n395), .B1(new_n380), .B2(G33), .ZN(new_n471));
  AND4_X1   g0271(.A1(KEYINPUT71), .A2(new_n371), .A3(new_n373), .A4(G33), .ZN(new_n472));
  OAI211_X1 g0272(.A(G257), .B(G1698), .C1(new_n471), .C2(new_n472), .ZN(new_n473));
  NAND2_X1  g0273(.A1(G33), .A2(G294), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n278), .A2(G250), .ZN(new_n475));
  AOI21_X1  g0275(.A(new_n475), .B1(new_n397), .B2(new_n398), .ZN(new_n476));
  OAI211_X1 g0276(.A(new_n473), .B(new_n474), .C1(KEYINPUT82), .C2(new_n476), .ZN(new_n477));
  AND2_X1   g0277(.A1(new_n476), .A2(KEYINPUT82), .ZN(new_n478));
  OAI21_X1  g0278(.A(new_n284), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  XNOR2_X1  g0279(.A(KEYINPUT5), .B(G41), .ZN(new_n480));
  NOR2_X1   g0280(.A1(new_n289), .A2(G1), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  OR2_X1    g0282(.A1(new_n287), .A2(new_n482), .ZN(new_n483));
  INV_X1    g0283(.A(KEYINPUT83), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n482), .A2(new_n286), .ZN(new_n485));
  OAI21_X1  g0285(.A(new_n484), .B1(new_n485), .B2(new_n231), .ZN(new_n486));
  AOI21_X1  g0286(.A(new_n284), .B1(new_n481), .B2(new_n480), .ZN(new_n487));
  NAND3_X1  g0287(.A1(new_n487), .A2(KEYINPUT83), .A3(G264), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n486), .A2(new_n488), .ZN(new_n489));
  NAND4_X1  g0289(.A1(new_n479), .A2(new_n297), .A3(new_n483), .A4(new_n489), .ZN(new_n490));
  NOR2_X1   g0290(.A1(new_n287), .A2(new_n482), .ZN(new_n491));
  AOI21_X1  g0291(.A(KEYINPUT83), .B1(new_n487), .B2(G264), .ZN(new_n492));
  AND4_X1   g0292(.A1(KEYINPUT83), .A2(new_n482), .A3(G264), .A4(new_n286), .ZN(new_n493));
  OAI21_X1  g0293(.A(KEYINPUT84), .B1(new_n492), .B2(new_n493), .ZN(new_n494));
  INV_X1    g0294(.A(KEYINPUT84), .ZN(new_n495));
  NAND3_X1  g0295(.A1(new_n486), .A2(new_n495), .A3(new_n488), .ZN(new_n496));
  AOI21_X1  g0296(.A(new_n491), .B1(new_n494), .B2(new_n496), .ZN(new_n497));
  AOI21_X1  g0297(.A(G200), .B1(new_n497), .B2(new_n479), .ZN(new_n498));
  INV_X1    g0298(.A(KEYINPUT85), .ZN(new_n499));
  OAI21_X1  g0299(.A(new_n490), .B1(new_n498), .B2(new_n499), .ZN(new_n500));
  AOI211_X1 g0300(.A(KEYINPUT85), .B(G200), .C1(new_n497), .C2(new_n479), .ZN(new_n501));
  OAI211_X1 g0301(.A(new_n461), .B(new_n470), .C1(new_n500), .C2(new_n501), .ZN(new_n502));
  NAND3_X1  g0302(.A1(new_n479), .A2(new_n483), .A3(new_n489), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n503), .A2(G169), .ZN(new_n504));
  NAND3_X1  g0304(.A1(new_n497), .A2(new_n479), .A3(G179), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  INV_X1    g0306(.A(KEYINPUT22), .ZN(new_n507));
  AOI211_X1 g0307(.A(G20), .B(new_n225), .C1(new_n397), .C2(new_n398), .ZN(new_n508));
  AOI21_X1  g0308(.A(new_n507), .B1(new_n508), .B2(KEYINPUT79), .ZN(new_n509));
  INV_X1    g0309(.A(new_n449), .ZN(new_n510));
  AOI21_X1  g0310(.A(new_n443), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  INV_X1    g0311(.A(new_n458), .ZN(new_n512));
  OAI21_X1  g0312(.A(KEYINPUT24), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  NAND3_X1  g0313(.A1(new_n450), .A2(new_n451), .A3(new_n458), .ZN(new_n514));
  AOI21_X1  g0314(.A(new_n256), .B1(new_n513), .B2(new_n514), .ZN(new_n515));
  INV_X1    g0315(.A(new_n470), .ZN(new_n516));
  OAI21_X1  g0316(.A(new_n506), .B1(new_n515), .B2(new_n516), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n502), .A2(new_n517), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n487), .A2(G257), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n483), .A2(new_n519), .ZN(new_n520));
  NAND4_X1  g0320(.A1(new_n274), .A2(new_n276), .A3(G250), .A4(G1698), .ZN(new_n521));
  NAND2_X1  g0321(.A1(G33), .A2(G283), .ZN(new_n522));
  AND2_X1   g0322(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  INV_X1    g0323(.A(KEYINPUT4), .ZN(new_n524));
  NOR2_X1   g0324(.A1(new_n524), .A2(new_n230), .ZN(new_n525));
  NAND3_X1  g0325(.A1(new_n352), .A2(new_n278), .A3(new_n525), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n278), .A2(G244), .ZN(new_n527));
  AOI21_X1  g0327(.A(new_n527), .B1(new_n397), .B2(new_n398), .ZN(new_n528));
  OAI211_X1 g0328(.A(new_n523), .B(new_n526), .C1(new_n528), .C2(KEYINPUT4), .ZN(new_n529));
  AOI21_X1  g0329(.A(new_n520), .B1(new_n529), .B2(new_n284), .ZN(new_n530));
  INV_X1    g0330(.A(KEYINPUT77), .ZN(new_n531));
  NAND3_X1  g0331(.A1(new_n530), .A2(new_n531), .A3(new_n303), .ZN(new_n532));
  AOI21_X1  g0332(.A(new_n491), .B1(G257), .B2(new_n487), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n523), .A2(new_n526), .ZN(new_n534));
  OAI211_X1 g0334(.A(G244), .B(new_n278), .C1(new_n471), .C2(new_n472), .ZN(new_n535));
  AOI21_X1  g0335(.A(new_n534), .B1(new_n535), .B2(new_n524), .ZN(new_n536));
  OAI21_X1  g0336(.A(new_n533), .B1(new_n536), .B2(new_n286), .ZN(new_n537));
  OAI21_X1  g0337(.A(KEYINPUT77), .B1(new_n537), .B2(G179), .ZN(new_n538));
  NOR2_X1   g0338(.A1(new_n530), .A2(G169), .ZN(new_n539));
  OAI21_X1  g0339(.A(new_n532), .B1(new_n538), .B2(new_n539), .ZN(new_n540));
  AOI21_X1  g0340(.A(new_n206), .B1(new_n384), .B2(new_n386), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n261), .A2(G77), .ZN(new_n542));
  INV_X1    g0342(.A(KEYINPUT6), .ZN(new_n543));
  NOR3_X1   g0343(.A1(new_n543), .A2(new_n205), .A3(G107), .ZN(new_n544));
  XNOR2_X1  g0344(.A(G97), .B(G107), .ZN(new_n545));
  AOI21_X1  g0345(.A(new_n544), .B1(new_n545), .B2(new_n543), .ZN(new_n546));
  OAI21_X1  g0346(.A(new_n542), .B1(new_n546), .B2(new_n210), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n547), .A2(KEYINPUT75), .ZN(new_n548));
  INV_X1    g0348(.A(KEYINPUT75), .ZN(new_n549));
  OAI211_X1 g0349(.A(new_n549), .B(new_n542), .C1(new_n546), .C2(new_n210), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n548), .A2(new_n550), .ZN(new_n551));
  OAI21_X1  g0351(.A(new_n255), .B1(new_n541), .B2(new_n551), .ZN(new_n552));
  NOR2_X1   g0352(.A1(new_n265), .A2(G97), .ZN(new_n553));
  AOI21_X1  g0353(.A(new_n553), .B1(new_n469), .B2(G97), .ZN(new_n554));
  AOI21_X1  g0354(.A(KEYINPUT76), .B1(new_n552), .B2(new_n554), .ZN(new_n555));
  INV_X1    g0355(.A(new_n555), .ZN(new_n556));
  INV_X1    g0356(.A(new_n554), .ZN(new_n557));
  OAI211_X1 g0357(.A(new_n550), .B(new_n548), .C1(new_n421), .C2(new_n206), .ZN(new_n558));
  AOI21_X1  g0358(.A(new_n557), .B1(new_n558), .B2(new_n255), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n559), .A2(KEYINPUT76), .ZN(new_n560));
  NAND3_X1  g0360(.A1(new_n540), .A2(new_n556), .A3(new_n560), .ZN(new_n561));
  OAI211_X1 g0361(.A(new_n522), .B(new_n210), .C1(G33), .C2(new_n205), .ZN(new_n562));
  OAI211_X1 g0362(.A(new_n562), .B(new_n255), .C1(new_n210), .C2(G116), .ZN(new_n563));
  INV_X1    g0363(.A(KEYINPUT20), .ZN(new_n564));
  XNOR2_X1  g0364(.A(new_n563), .B(new_n564), .ZN(new_n565));
  NOR2_X1   g0365(.A1(new_n265), .A2(G116), .ZN(new_n566));
  AOI21_X1  g0366(.A(new_n566), .B1(new_n469), .B2(G116), .ZN(new_n567));
  AND2_X1   g0367(.A1(new_n565), .A2(new_n567), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n231), .A2(G1698), .ZN(new_n569));
  OAI21_X1  g0369(.A(new_n569), .B1(G257), .B2(G1698), .ZN(new_n570));
  AOI21_X1  g0370(.A(new_n570), .B1(new_n397), .B2(new_n398), .ZN(new_n571));
  INV_X1    g0371(.A(G303), .ZN(new_n572));
  NOR2_X1   g0372(.A1(new_n352), .A2(new_n572), .ZN(new_n573));
  OAI21_X1  g0373(.A(new_n284), .B1(new_n571), .B2(new_n573), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n487), .A2(G270), .ZN(new_n575));
  NAND3_X1  g0375(.A1(new_n574), .A2(new_n483), .A3(new_n575), .ZN(new_n576));
  OAI21_X1  g0376(.A(new_n568), .B1(new_n576), .B2(new_n433), .ZN(new_n577));
  AOI21_X1  g0377(.A(new_n577), .B1(G200), .B2(new_n576), .ZN(new_n578));
  AND2_X1   g0378(.A1(new_n574), .A2(new_n575), .ZN(new_n579));
  AOI21_X1  g0379(.A(new_n303), .B1(new_n565), .B2(new_n567), .ZN(new_n580));
  NAND3_X1  g0380(.A1(new_n579), .A2(new_n580), .A3(new_n483), .ZN(new_n581));
  AOI21_X1  g0381(.A(new_n300), .B1(new_n565), .B2(new_n567), .ZN(new_n582));
  NAND3_X1  g0382(.A1(new_n582), .A2(new_n576), .A3(KEYINPUT21), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n581), .A2(new_n583), .ZN(new_n584));
  AOI21_X1  g0384(.A(KEYINPUT21), .B1(new_n582), .B2(new_n576), .ZN(new_n585));
  NOR3_X1   g0385(.A1(new_n578), .A2(new_n584), .A3(new_n585), .ZN(new_n586));
  NOR2_X1   g0386(.A1(new_n343), .A2(new_n265), .ZN(new_n587));
  OAI211_X1 g0387(.A(new_n210), .B(G68), .C1(new_n471), .C2(new_n472), .ZN(new_n588));
  OAI22_X1  g0388(.A1(new_n325), .A2(G20), .B1(new_n207), .B2(G87), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n589), .A2(KEYINPUT19), .ZN(new_n590));
  NOR3_X1   g0390(.A1(new_n259), .A2(KEYINPUT19), .A3(new_n205), .ZN(new_n591));
  INV_X1    g0391(.A(new_n591), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n590), .A2(new_n592), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n588), .A2(new_n593), .ZN(new_n594));
  AOI21_X1  g0394(.A(new_n587), .B1(new_n594), .B2(new_n255), .ZN(new_n595));
  INV_X1    g0395(.A(new_n469), .ZN(new_n596));
  OAI21_X1  g0396(.A(new_n595), .B1(new_n342), .B2(new_n596), .ZN(new_n597));
  NOR2_X1   g0397(.A1(G238), .A2(G1698), .ZN(new_n598));
  AOI21_X1  g0398(.A(new_n598), .B1(new_n230), .B2(G1698), .ZN(new_n599));
  OAI21_X1  g0399(.A(new_n599), .B1(new_n471), .B2(new_n472), .ZN(new_n600));
  AOI21_X1  g0400(.A(new_n286), .B1(new_n600), .B2(new_n453), .ZN(new_n601));
  NOR2_X1   g0401(.A1(new_n481), .A2(new_n226), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n286), .A2(new_n602), .ZN(new_n603));
  INV_X1    g0403(.A(new_n481), .ZN(new_n604));
  OAI21_X1  g0404(.A(new_n603), .B1(new_n287), .B2(new_n604), .ZN(new_n605));
  NOR2_X1   g0405(.A1(new_n601), .A2(new_n605), .ZN(new_n606));
  INV_X1    g0406(.A(KEYINPUT78), .ZN(new_n607));
  NAND3_X1  g0407(.A1(new_n606), .A2(new_n607), .A3(new_n303), .ZN(new_n608));
  INV_X1    g0408(.A(new_n599), .ZN(new_n609));
  AOI21_X1  g0409(.A(new_n609), .B1(new_n397), .B2(new_n398), .ZN(new_n610));
  INV_X1    g0410(.A(new_n453), .ZN(new_n611));
  OAI21_X1  g0411(.A(new_n284), .B1(new_n610), .B2(new_n611), .ZN(new_n612));
  INV_X1    g0412(.A(new_n605), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  OAI21_X1  g0414(.A(KEYINPUT78), .B1(new_n614), .B2(G179), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n614), .A2(new_n300), .ZN(new_n616));
  NAND4_X1  g0416(.A1(new_n597), .A2(new_n608), .A3(new_n615), .A4(new_n616), .ZN(new_n617));
  INV_X1    g0417(.A(new_n587), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n469), .A2(G87), .ZN(new_n619));
  AOI21_X1  g0419(.A(new_n591), .B1(new_n589), .B2(KEYINPUT19), .ZN(new_n620));
  AOI21_X1  g0420(.A(new_n620), .B1(new_n448), .B2(G68), .ZN(new_n621));
  OAI211_X1 g0421(.A(new_n618), .B(new_n619), .C1(new_n621), .C2(new_n256), .ZN(new_n622));
  INV_X1    g0422(.A(new_n622), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n606), .A2(G190), .ZN(new_n624));
  OAI21_X1  g0424(.A(G200), .B1(new_n601), .B2(new_n605), .ZN(new_n625));
  NAND3_X1  g0425(.A1(new_n623), .A2(new_n624), .A3(new_n625), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n617), .A2(new_n626), .ZN(new_n627));
  INV_X1    g0427(.A(new_n627), .ZN(new_n628));
  OAI211_X1 g0428(.A(G190), .B(new_n533), .C1(new_n536), .C2(new_n286), .ZN(new_n629));
  OAI21_X1  g0429(.A(new_n629), .B1(new_n530), .B2(new_n429), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n552), .A2(new_n554), .ZN(new_n631));
  NOR2_X1   g0431(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  INV_X1    g0432(.A(new_n632), .ZN(new_n633));
  NAND4_X1  g0433(.A1(new_n561), .A2(new_n586), .A3(new_n628), .A4(new_n633), .ZN(new_n634));
  NOR3_X1   g0434(.A1(new_n442), .A2(new_n518), .A3(new_n634), .ZN(G372));
  INV_X1    g0435(.A(new_n306), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n340), .A2(new_n361), .ZN(new_n637));
  AND2_X1   g0437(.A1(new_n637), .A2(new_n337), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n438), .A2(new_n439), .ZN(new_n639));
  OAI211_X1 g0439(.A(new_n420), .B(new_n428), .C1(new_n638), .C2(new_n639), .ZN(new_n640));
  AOI21_X1  g0440(.A(new_n636), .B1(new_n640), .B2(new_n299), .ZN(new_n641));
  OAI211_X1 g0441(.A(new_n597), .B(new_n616), .C1(G179), .C2(new_n614), .ZN(new_n642));
  INV_X1    g0442(.A(KEYINPUT76), .ZN(new_n643));
  AOI211_X1 g0443(.A(new_n643), .B(new_n557), .C1(new_n558), .C2(new_n255), .ZN(new_n644));
  NOR2_X1   g0444(.A1(new_n644), .A2(new_n555), .ZN(new_n645));
  AOI21_X1  g0445(.A(new_n632), .B1(new_n645), .B2(new_n540), .ZN(new_n646));
  AOI22_X1  g0446(.A1(new_n461), .A2(new_n470), .B1(new_n504), .B2(new_n505), .ZN(new_n647));
  NOR2_X1   g0447(.A1(new_n584), .A2(new_n585), .ZN(new_n648));
  INV_X1    g0448(.A(new_n648), .ZN(new_n649));
  OAI211_X1 g0449(.A(new_n646), .B(new_n502), .C1(new_n647), .C2(new_n649), .ZN(new_n650));
  AOI21_X1  g0450(.A(new_n429), .B1(new_n612), .B2(new_n613), .ZN(new_n651));
  OAI21_X1  g0451(.A(KEYINPUT86), .B1(new_n622), .B2(new_n651), .ZN(new_n652));
  INV_X1    g0452(.A(KEYINPUT86), .ZN(new_n653));
  NAND4_X1  g0453(.A1(new_n625), .A2(new_n595), .A3(new_n653), .A4(new_n619), .ZN(new_n654));
  NAND3_X1  g0454(.A1(new_n652), .A2(new_n654), .A3(new_n624), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n655), .A2(new_n642), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n656), .A2(KEYINPUT87), .ZN(new_n657));
  INV_X1    g0457(.A(KEYINPUT87), .ZN(new_n658));
  NAND3_X1  g0458(.A1(new_n655), .A2(new_n642), .A3(new_n658), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n657), .A2(new_n659), .ZN(new_n660));
  INV_X1    g0460(.A(new_n660), .ZN(new_n661));
  OAI21_X1  g0461(.A(new_n642), .B1(new_n650), .B2(new_n661), .ZN(new_n662));
  INV_X1    g0462(.A(KEYINPUT26), .ZN(new_n663));
  NOR3_X1   g0463(.A1(new_n561), .A2(new_n663), .A3(new_n627), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n540), .A2(new_n631), .ZN(new_n665));
  INV_X1    g0465(.A(new_n665), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n660), .A2(new_n666), .ZN(new_n667));
  AOI21_X1  g0467(.A(new_n664), .B1(new_n667), .B2(new_n663), .ZN(new_n668));
  NOR2_X1   g0468(.A1(new_n662), .A2(new_n668), .ZN(new_n669));
  OAI21_X1  g0469(.A(new_n641), .B1(new_n442), .B2(new_n669), .ZN(G369));
  NAND3_X1  g0470(.A1(new_n209), .A2(new_n210), .A3(G13), .ZN(new_n671));
  XNOR2_X1  g0471(.A(new_n671), .B(KEYINPUT88), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n672), .A2(KEYINPUT27), .ZN(new_n673));
  OR2_X1    g0473(.A1(new_n671), .A2(KEYINPUT88), .ZN(new_n674));
  INV_X1    g0474(.A(KEYINPUT27), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n671), .A2(KEYINPUT88), .ZN(new_n676));
  NAND3_X1  g0476(.A1(new_n674), .A2(new_n675), .A3(new_n676), .ZN(new_n677));
  NAND3_X1  g0477(.A1(new_n673), .A2(new_n677), .A3(G213), .ZN(new_n678));
  INV_X1    g0478(.A(G343), .ZN(new_n679));
  NOR2_X1   g0479(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  INV_X1    g0480(.A(KEYINPUT89), .ZN(new_n681));
  XNOR2_X1  g0481(.A(new_n680), .B(new_n681), .ZN(new_n682));
  NOR2_X1   g0482(.A1(new_n517), .A2(new_n682), .ZN(new_n683));
  OAI21_X1  g0483(.A(new_n682), .B1(new_n515), .B2(new_n516), .ZN(new_n684));
  NAND3_X1  g0484(.A1(new_n502), .A2(new_n517), .A3(new_n684), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n647), .A2(new_n682), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n687), .A2(KEYINPUT90), .ZN(new_n688));
  INV_X1    g0488(.A(KEYINPUT90), .ZN(new_n689));
  NAND3_X1  g0489(.A1(new_n685), .A2(new_n689), .A3(new_n686), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n688), .A2(new_n690), .ZN(new_n691));
  NOR2_X1   g0491(.A1(new_n648), .A2(new_n682), .ZN(new_n692));
  AOI21_X1  g0492(.A(new_n683), .B1(new_n691), .B2(new_n692), .ZN(new_n693));
  XNOR2_X1  g0493(.A(new_n680), .B(KEYINPUT89), .ZN(new_n694));
  NOR2_X1   g0494(.A1(new_n694), .A2(new_n568), .ZN(new_n695));
  MUX2_X1   g0495(.A(new_n586), .B(new_n649), .S(new_n695), .Z(new_n696));
  NAND2_X1  g0496(.A1(new_n696), .A2(G330), .ZN(new_n697));
  INV_X1    g0497(.A(new_n697), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n691), .A2(new_n698), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n693), .A2(new_n699), .ZN(new_n700));
  XNOR2_X1  g0500(.A(new_n700), .B(KEYINPUT91), .ZN(G399));
  INV_X1    g0501(.A(new_n213), .ZN(new_n702));
  NOR2_X1   g0502(.A1(new_n702), .A2(G41), .ZN(new_n703));
  INV_X1    g0503(.A(new_n703), .ZN(new_n704));
  NOR3_X1   g0504(.A1(new_n207), .A2(G87), .A3(G116), .ZN(new_n705));
  NAND3_X1  g0505(.A1(new_n704), .A2(G1), .A3(new_n705), .ZN(new_n706));
  OAI21_X1  g0506(.A(new_n706), .B1(new_n217), .B2(new_n704), .ZN(new_n707));
  XNOR2_X1  g0507(.A(new_n707), .B(KEYINPUT28), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n667), .A2(KEYINPUT26), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n517), .A2(new_n648), .ZN(new_n710));
  NAND4_X1  g0510(.A1(new_n710), .A2(new_n502), .A3(new_n660), .A4(new_n646), .ZN(new_n711));
  AND3_X1   g0511(.A1(new_n540), .A2(new_n556), .A3(new_n560), .ZN(new_n712));
  NAND3_X1  g0512(.A1(new_n712), .A2(new_n663), .A3(new_n628), .ZN(new_n713));
  NAND4_X1  g0513(.A1(new_n709), .A2(new_n711), .A3(new_n642), .A4(new_n713), .ZN(new_n714));
  NAND3_X1  g0514(.A1(new_n714), .A2(KEYINPUT29), .A3(new_n694), .ZN(new_n715));
  INV_X1    g0515(.A(new_n715), .ZN(new_n716));
  INV_X1    g0516(.A(KEYINPUT29), .ZN(new_n717));
  NAND3_X1  g0517(.A1(new_n712), .A2(KEYINPUT26), .A3(new_n628), .ZN(new_n718));
  AOI21_X1  g0518(.A(new_n665), .B1(new_n657), .B2(new_n659), .ZN(new_n719));
  OAI21_X1  g0519(.A(new_n718), .B1(new_n719), .B2(KEYINPUT26), .ZN(new_n720));
  NAND3_X1  g0520(.A1(new_n720), .A2(new_n711), .A3(new_n642), .ZN(new_n721));
  INV_X1    g0521(.A(KEYINPUT92), .ZN(new_n722));
  AND3_X1   g0522(.A1(new_n721), .A2(new_n722), .A3(new_n694), .ZN(new_n723));
  AOI21_X1  g0523(.A(new_n722), .B1(new_n721), .B2(new_n694), .ZN(new_n724));
  OAI21_X1  g0524(.A(new_n717), .B1(new_n723), .B2(new_n724), .ZN(new_n725));
  NAND2_X1  g0525(.A1(new_n725), .A2(KEYINPUT93), .ZN(new_n726));
  INV_X1    g0526(.A(KEYINPUT93), .ZN(new_n727));
  OAI211_X1 g0527(.A(new_n727), .B(new_n717), .C1(new_n723), .C2(new_n724), .ZN(new_n728));
  AOI21_X1  g0528(.A(new_n716), .B1(new_n726), .B2(new_n728), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n497), .A2(new_n479), .ZN(new_n730));
  INV_X1    g0530(.A(new_n730), .ZN(new_n731));
  NAND4_X1  g0531(.A1(new_n612), .A2(new_n574), .A3(new_n613), .A4(new_n575), .ZN(new_n732));
  NOR2_X1   g0532(.A1(new_n537), .A2(new_n732), .ZN(new_n733));
  NAND4_X1  g0533(.A1(new_n731), .A2(KEYINPUT30), .A3(G179), .A4(new_n733), .ZN(new_n734));
  INV_X1    g0534(.A(KEYINPUT30), .ZN(new_n735));
  NAND3_X1  g0535(.A1(new_n530), .A2(new_n606), .A3(new_n579), .ZN(new_n736));
  OAI21_X1  g0536(.A(new_n735), .B1(new_n505), .B2(new_n736), .ZN(new_n737));
  NOR3_X1   g0537(.A1(new_n530), .A2(G179), .A3(new_n606), .ZN(new_n738));
  NAND3_X1  g0538(.A1(new_n738), .A2(new_n730), .A3(new_n576), .ZN(new_n739));
  NAND3_X1  g0539(.A1(new_n734), .A2(new_n737), .A3(new_n739), .ZN(new_n740));
  NAND3_X1  g0540(.A1(new_n740), .A2(KEYINPUT31), .A3(new_n682), .ZN(new_n741));
  INV_X1    g0541(.A(new_n741), .ZN(new_n742));
  AOI21_X1  g0542(.A(KEYINPUT31), .B1(new_n740), .B2(new_n682), .ZN(new_n743));
  NOR2_X1   g0543(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  AND4_X1   g0544(.A1(new_n561), .A2(new_n586), .A3(new_n633), .A4(new_n628), .ZN(new_n745));
  NAND4_X1  g0545(.A1(new_n745), .A2(new_n517), .A3(new_n502), .A4(new_n694), .ZN(new_n746));
  NAND2_X1  g0546(.A1(new_n744), .A2(new_n746), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n747), .A2(G330), .ZN(new_n748));
  INV_X1    g0548(.A(new_n748), .ZN(new_n749));
  NOR2_X1   g0549(.A1(new_n729), .A2(new_n749), .ZN(new_n750));
  OAI21_X1  g0550(.A(new_n708), .B1(new_n750), .B2(G1), .ZN(G364));
  INV_X1    g0551(.A(G13), .ZN(new_n752));
  NOR3_X1   g0552(.A1(new_n752), .A2(new_n289), .A3(G20), .ZN(new_n753));
  OR2_X1    g0553(.A1(new_n753), .A2(KEYINPUT94), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n753), .A2(KEYINPUT94), .ZN(new_n755));
  NAND3_X1  g0555(.A1(new_n754), .A2(G1), .A3(new_n755), .ZN(new_n756));
  NOR2_X1   g0556(.A1(new_n703), .A2(new_n756), .ZN(new_n757));
  NOR2_X1   g0557(.A1(new_n696), .A2(G330), .ZN(new_n758));
  NOR3_X1   g0558(.A1(new_n698), .A2(new_n757), .A3(new_n758), .ZN(new_n759));
  XOR2_X1   g0559(.A(new_n759), .B(KEYINPUT95), .Z(new_n760));
  NAND2_X1  g0560(.A1(new_n213), .A2(new_n352), .ZN(new_n761));
  INV_X1    g0561(.A(G355), .ZN(new_n762));
  OAI22_X1  g0562(.A1(new_n761), .A2(new_n762), .B1(G116), .B2(new_n213), .ZN(new_n763));
  NOR2_X1   g0563(.A1(new_n217), .A2(G45), .ZN(new_n764));
  AOI21_X1  g0564(.A(new_n764), .B1(new_n252), .B2(G45), .ZN(new_n765));
  NOR2_X1   g0565(.A1(new_n445), .A2(new_n702), .ZN(new_n766));
  AOI21_X1  g0566(.A(new_n763), .B1(new_n765), .B2(new_n766), .ZN(new_n767));
  NOR2_X1   g0567(.A1(G13), .A2(G33), .ZN(new_n768));
  INV_X1    g0568(.A(new_n768), .ZN(new_n769));
  NOR2_X1   g0569(.A1(new_n769), .A2(G20), .ZN(new_n770));
  AOI21_X1  g0570(.A(new_n219), .B1(G20), .B2(new_n300), .ZN(new_n771));
  NOR2_X1   g0571(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  INV_X1    g0572(.A(new_n772), .ZN(new_n773));
  OAI21_X1  g0573(.A(new_n757), .B1(new_n767), .B2(new_n773), .ZN(new_n774));
  INV_X1    g0574(.A(new_n770), .ZN(new_n775));
  NOR2_X1   g0575(.A1(new_n696), .A2(new_n775), .ZN(new_n776));
  NOR3_X1   g0576(.A1(new_n210), .A2(new_n303), .A3(G200), .ZN(new_n777));
  NAND2_X1  g0577(.A1(new_n434), .A2(new_n777), .ZN(new_n778));
  INV_X1    g0578(.A(new_n778), .ZN(new_n779));
  AOI21_X1  g0579(.A(new_n352), .B1(new_n779), .B2(G322), .ZN(new_n780));
  NOR3_X1   g0580(.A1(new_n210), .A2(new_n303), .A3(new_n429), .ZN(new_n781));
  INV_X1    g0581(.A(new_n781), .ZN(new_n782));
  NOR2_X1   g0582(.A1(new_n782), .A2(G190), .ZN(new_n783));
  INV_X1    g0583(.A(new_n783), .ZN(new_n784));
  XOR2_X1   g0584(.A(KEYINPUT33), .B(G317), .Z(new_n785));
  OAI21_X1  g0585(.A(new_n780), .B1(new_n784), .B2(new_n785), .ZN(new_n786));
  NOR4_X1   g0586(.A1(new_n210), .A2(G179), .A3(G190), .A4(G200), .ZN(new_n787));
  INV_X1    g0587(.A(new_n787), .ZN(new_n788));
  OR2_X1    g0588(.A1(new_n788), .A2(KEYINPUT96), .ZN(new_n789));
  NAND2_X1  g0589(.A1(new_n788), .A2(KEYINPUT96), .ZN(new_n790));
  NAND2_X1  g0590(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  INV_X1    g0591(.A(new_n791), .ZN(new_n792));
  AOI21_X1  g0592(.A(new_n786), .B1(G329), .B2(new_n792), .ZN(new_n793));
  NAND2_X1  g0593(.A1(new_n777), .A2(new_n297), .ZN(new_n794));
  INV_X1    g0594(.A(G311), .ZN(new_n795));
  NOR3_X1   g0595(.A1(new_n297), .A2(G179), .A3(G200), .ZN(new_n796));
  NOR2_X1   g0596(.A1(new_n796), .A2(new_n210), .ZN(new_n797));
  INV_X1    g0597(.A(G294), .ZN(new_n798));
  OAI22_X1  g0598(.A1(new_n794), .A2(new_n795), .B1(new_n797), .B2(new_n798), .ZN(new_n799));
  NOR2_X1   g0599(.A1(new_n782), .A2(new_n433), .ZN(new_n800));
  AOI21_X1  g0600(.A(new_n799), .B1(G326), .B2(new_n800), .ZN(new_n801));
  XNOR2_X1  g0601(.A(new_n801), .B(KEYINPUT100), .ZN(new_n802));
  AOI21_X1  g0602(.A(KEYINPUT98), .B1(new_n303), .B2(G200), .ZN(new_n803));
  NOR2_X1   g0603(.A1(new_n803), .A2(new_n210), .ZN(new_n804));
  NAND3_X1  g0604(.A1(new_n303), .A2(KEYINPUT98), .A3(G200), .ZN(new_n805));
  NAND2_X1  g0605(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  NOR2_X1   g0606(.A1(new_n806), .A2(G190), .ZN(new_n807));
  NOR2_X1   g0607(.A1(new_n806), .A2(new_n297), .ZN(new_n808));
  AOI22_X1  g0608(.A1(G283), .A2(new_n807), .B1(new_n808), .B2(G303), .ZN(new_n809));
  NAND3_X1  g0609(.A1(new_n793), .A2(new_n802), .A3(new_n809), .ZN(new_n810));
  XNOR2_X1  g0610(.A(KEYINPUT97), .B(G159), .ZN(new_n811));
  NAND2_X1  g0611(.A1(new_n792), .A2(new_n811), .ZN(new_n812));
  XOR2_X1   g0612(.A(new_n812), .B(KEYINPUT32), .Z(new_n813));
  INV_X1    g0613(.A(new_n794), .ZN(new_n814));
  AOI22_X1  g0614(.A1(new_n779), .A2(G58), .B1(G77), .B2(new_n814), .ZN(new_n815));
  INV_X1    g0615(.A(new_n797), .ZN(new_n816));
  NAND2_X1  g0616(.A1(new_n816), .A2(G97), .ZN(new_n817));
  AOI22_X1  g0617(.A1(G50), .A2(new_n800), .B1(new_n783), .B2(G68), .ZN(new_n818));
  NAND4_X1  g0618(.A1(new_n813), .A2(new_n815), .A3(new_n817), .A4(new_n818), .ZN(new_n819));
  NAND2_X1  g0619(.A1(new_n808), .A2(G87), .ZN(new_n820));
  INV_X1    g0620(.A(new_n807), .ZN(new_n821));
  OAI211_X1 g0621(.A(new_n820), .B(new_n352), .C1(new_n821), .C2(new_n206), .ZN(new_n822));
  XOR2_X1   g0622(.A(new_n822), .B(KEYINPUT99), .Z(new_n823));
  OAI21_X1  g0623(.A(new_n810), .B1(new_n819), .B2(new_n823), .ZN(new_n824));
  AOI211_X1 g0624(.A(new_n774), .B(new_n776), .C1(new_n771), .C2(new_n824), .ZN(new_n825));
  NOR2_X1   g0625(.A1(new_n760), .A2(new_n825), .ZN(new_n826));
  INV_X1    g0626(.A(new_n826), .ZN(G396));
  INV_X1    g0627(.A(new_n724), .ZN(new_n828));
  NAND3_X1  g0628(.A1(new_n721), .A2(new_n722), .A3(new_n694), .ZN(new_n829));
  NAND2_X1  g0629(.A1(new_n828), .A2(new_n829), .ZN(new_n830));
  INV_X1    g0630(.A(KEYINPUT103), .ZN(new_n831));
  NAND2_X1  g0631(.A1(new_n363), .A2(new_n364), .ZN(new_n832));
  NAND2_X1  g0632(.A1(new_n682), .A2(new_n349), .ZN(new_n833));
  INV_X1    g0633(.A(new_n360), .ZN(new_n834));
  NAND2_X1  g0634(.A1(new_n359), .A2(new_n303), .ZN(new_n835));
  AOI22_X1  g0635(.A1(new_n832), .A2(new_n833), .B1(new_n834), .B2(new_n835), .ZN(new_n836));
  AND3_X1   g0636(.A1(new_n834), .A2(new_n835), .A3(new_n694), .ZN(new_n837));
  OAI21_X1  g0637(.A(new_n831), .B1(new_n836), .B2(new_n837), .ZN(new_n838));
  NAND3_X1  g0638(.A1(new_n834), .A2(new_n835), .A3(new_n694), .ZN(new_n839));
  AOI22_X1  g0639(.A1(new_n363), .A2(new_n364), .B1(new_n682), .B2(new_n349), .ZN(new_n840));
  OAI211_X1 g0640(.A(KEYINPUT103), .B(new_n839), .C1(new_n840), .C2(new_n361), .ZN(new_n841));
  AND2_X1   g0641(.A1(new_n838), .A2(new_n841), .ZN(new_n842));
  NAND2_X1  g0642(.A1(new_n830), .A2(new_n842), .ZN(new_n843));
  AOI21_X1  g0643(.A(new_n682), .B1(new_n838), .B2(new_n841), .ZN(new_n844));
  OAI21_X1  g0644(.A(new_n844), .B1(new_n662), .B2(new_n668), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n843), .A2(new_n845), .ZN(new_n846));
  AOI21_X1  g0646(.A(new_n757), .B1(new_n846), .B2(new_n748), .ZN(new_n847));
  NAND3_X1  g0647(.A1(new_n843), .A2(new_n749), .A3(new_n845), .ZN(new_n848));
  NAND2_X1  g0648(.A1(new_n847), .A2(new_n848), .ZN(new_n849));
  OR2_X1    g0649(.A1(new_n771), .A2(new_n768), .ZN(new_n850));
  OAI21_X1  g0650(.A(new_n757), .B1(G77), .B2(new_n850), .ZN(new_n851));
  INV_X1    g0651(.A(G116), .ZN(new_n852));
  OAI22_X1  g0652(.A1(new_n778), .A2(new_n798), .B1(new_n852), .B2(new_n794), .ZN(new_n853));
  INV_X1    g0653(.A(new_n800), .ZN(new_n854));
  OAI221_X1 g0654(.A(new_n817), .B1(new_n572), .B2(new_n854), .C1(new_n791), .C2(new_n795), .ZN(new_n855));
  AOI211_X1 g0655(.A(new_n853), .B(new_n855), .C1(G283), .C2(new_n783), .ZN(new_n856));
  AOI21_X1  g0656(.A(new_n352), .B1(new_n808), .B2(G107), .ZN(new_n857));
  XNOR2_X1  g0657(.A(new_n857), .B(KEYINPUT101), .ZN(new_n858));
  OAI211_X1 g0658(.A(new_n856), .B(new_n858), .C1(new_n225), .C2(new_n821), .ZN(new_n859));
  NOR2_X1   g0659(.A1(new_n821), .A2(new_n223), .ZN(new_n860));
  INV_X1    g0660(.A(G58), .ZN(new_n861));
  INV_X1    g0661(.A(G132), .ZN(new_n862));
  OAI221_X1 g0662(.A(new_n445), .B1(new_n861), .B2(new_n797), .C1(new_n791), .C2(new_n862), .ZN(new_n863));
  AOI211_X1 g0663(.A(new_n860), .B(new_n863), .C1(G50), .C2(new_n808), .ZN(new_n864));
  XNOR2_X1  g0664(.A(new_n864), .B(KEYINPUT102), .ZN(new_n865));
  AOI22_X1  g0665(.A1(new_n779), .A2(G143), .B1(G150), .B2(new_n783), .ZN(new_n866));
  AOI22_X1  g0666(.A1(new_n800), .A2(G137), .B1(new_n814), .B2(new_n811), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  XOR2_X1   g0668(.A(new_n868), .B(KEYINPUT34), .Z(new_n869));
  OAI21_X1  g0669(.A(new_n859), .B1(new_n865), .B2(new_n869), .ZN(new_n870));
  AOI21_X1  g0670(.A(new_n851), .B1(new_n870), .B2(new_n771), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n838), .A2(new_n841), .ZN(new_n872));
  OAI21_X1  g0672(.A(new_n871), .B1(new_n872), .B2(new_n769), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n849), .A2(new_n873), .ZN(G384));
  INV_X1    g0674(.A(new_n546), .ZN(new_n875));
  OR2_X1    g0675(.A1(new_n875), .A2(KEYINPUT35), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n875), .A2(KEYINPUT35), .ZN(new_n877));
  NAND4_X1  g0677(.A1(new_n876), .A2(new_n877), .A3(G116), .A4(new_n220), .ZN(new_n878));
  XNOR2_X1  g0678(.A(KEYINPUT104), .B(KEYINPUT36), .ZN(new_n879));
  XNOR2_X1  g0679(.A(new_n878), .B(new_n879), .ZN(new_n880));
  NAND3_X1  g0680(.A1(new_n218), .A2(G77), .A3(new_n389), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n202), .A2(G68), .ZN(new_n882));
  AOI211_X1 g0682(.A(new_n209), .B(G13), .C1(new_n881), .C2(new_n882), .ZN(new_n883));
  NOR2_X1   g0683(.A1(new_n880), .A2(new_n883), .ZN(new_n884));
  INV_X1    g0684(.A(new_n641), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n726), .A2(new_n728), .ZN(new_n886));
  NOR2_X1   g0686(.A1(new_n442), .A2(new_n716), .ZN(new_n887));
  AOI21_X1  g0687(.A(new_n885), .B1(new_n886), .B2(new_n887), .ZN(new_n888));
  INV_X1    g0688(.A(new_n678), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n405), .A2(new_n889), .ZN(new_n890));
  OAI211_X1 g0690(.A(new_n436), .B(new_n890), .C1(new_n419), .C2(KEYINPUT107), .ZN(new_n891));
  INV_X1    g0691(.A(KEYINPUT37), .ZN(new_n892));
  INV_X1    g0692(.A(KEYINPUT107), .ZN(new_n893));
  OAI21_X1  g0693(.A(new_n892), .B1(new_n426), .B2(new_n893), .ZN(new_n894));
  AOI21_X1  g0694(.A(KEYINPUT16), .B1(new_n402), .B2(new_n391), .ZN(new_n895));
  OAI21_X1  g0695(.A(new_n369), .B1(new_n404), .B2(new_n895), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n418), .A2(new_n896), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n896), .A2(new_n889), .ZN(new_n898));
  AND3_X1   g0698(.A1(new_n897), .A2(new_n898), .A3(new_n436), .ZN(new_n899));
  OAI22_X1  g0699(.A1(new_n891), .A2(new_n894), .B1(new_n899), .B2(new_n892), .ZN(new_n900));
  INV_X1    g0700(.A(new_n898), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n440), .A2(new_n901), .ZN(new_n902));
  AND3_X1   g0702(.A1(new_n900), .A2(new_n902), .A3(KEYINPUT38), .ZN(new_n903));
  AOI21_X1  g0703(.A(KEYINPUT38), .B1(new_n900), .B2(new_n902), .ZN(new_n904));
  NOR2_X1   g0704(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  INV_X1    g0705(.A(new_n905), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n337), .A2(KEYINPUT106), .ZN(new_n907));
  NOR2_X1   g0707(.A1(new_n694), .A2(new_n317), .ZN(new_n908));
  INV_X1    g0708(.A(new_n908), .ZN(new_n909));
  AND2_X1   g0709(.A1(new_n340), .A2(new_n909), .ZN(new_n910));
  INV_X1    g0710(.A(KEYINPUT106), .ZN(new_n911));
  OAI211_X1 g0711(.A(new_n911), .B(new_n318), .C1(new_n335), .C2(new_n336), .ZN(new_n912));
  NAND3_X1  g0712(.A1(new_n907), .A2(new_n910), .A3(new_n912), .ZN(new_n913));
  NOR2_X1   g0713(.A1(new_n335), .A2(new_n336), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n914), .A2(new_n340), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n915), .A2(new_n908), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n913), .A2(new_n916), .ZN(new_n917));
  AOI21_X1  g0717(.A(KEYINPUT105), .B1(new_n845), .B2(new_n839), .ZN(new_n918));
  INV_X1    g0718(.A(KEYINPUT105), .ZN(new_n919));
  AOI211_X1 g0719(.A(new_n919), .B(new_n837), .C1(new_n721), .C2(new_n844), .ZN(new_n920));
  OAI211_X1 g0720(.A(new_n906), .B(new_n917), .C1(new_n918), .C2(new_n920), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n420), .A2(new_n428), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n922), .A2(new_n678), .ZN(new_n923));
  NAND3_X1  g0723(.A1(new_n900), .A2(new_n902), .A3(KEYINPUT38), .ZN(new_n924));
  AOI21_X1  g0724(.A(new_n678), .B1(new_n425), .B2(new_n369), .ZN(new_n925));
  AND2_X1   g0725(.A1(new_n440), .A2(new_n925), .ZN(new_n926));
  AOI21_X1  g0726(.A(KEYINPUT37), .B1(new_n419), .B2(KEYINPUT107), .ZN(new_n927));
  AND3_X1   g0727(.A1(new_n425), .A2(new_n369), .A3(new_n435), .ZN(new_n928));
  NOR2_X1   g0728(.A1(new_n928), .A2(new_n925), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n426), .A2(new_n893), .ZN(new_n930));
  NAND3_X1  g0730(.A1(new_n927), .A2(new_n929), .A3(new_n930), .ZN(new_n931));
  NAND3_X1  g0731(.A1(new_n419), .A2(new_n890), .A3(new_n436), .ZN(new_n932));
  AOI22_X1  g0732(.A1(new_n931), .A2(KEYINPUT108), .B1(KEYINPUT37), .B2(new_n932), .ZN(new_n933));
  OR3_X1    g0733(.A1(new_n891), .A2(new_n894), .A3(KEYINPUT108), .ZN(new_n934));
  AOI21_X1  g0734(.A(new_n926), .B1(new_n933), .B2(new_n934), .ZN(new_n935));
  OAI21_X1  g0735(.A(new_n924), .B1(new_n935), .B2(KEYINPUT38), .ZN(new_n936));
  INV_X1    g0736(.A(KEYINPUT39), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  NOR3_X1   g0738(.A1(new_n903), .A2(new_n904), .A3(new_n937), .ZN(new_n939));
  INV_X1    g0739(.A(new_n939), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n938), .A2(new_n940), .ZN(new_n941));
  AOI21_X1  g0741(.A(new_n682), .B1(new_n907), .B2(new_n912), .ZN(new_n942));
  INV_X1    g0742(.A(new_n942), .ZN(new_n943));
  OAI211_X1 g0743(.A(new_n921), .B(new_n923), .C1(new_n941), .C2(new_n943), .ZN(new_n944));
  XOR2_X1   g0744(.A(new_n888), .B(new_n944), .Z(new_n945));
  AOI21_X1  g0745(.A(new_n842), .B1(new_n916), .B2(new_n913), .ZN(new_n946));
  NAND3_X1  g0746(.A1(new_n946), .A2(KEYINPUT40), .A3(new_n747), .ZN(new_n947));
  INV_X1    g0747(.A(new_n947), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n948), .A2(new_n936), .ZN(new_n949));
  OAI211_X1 g0749(.A(new_n946), .B(new_n747), .C1(new_n903), .C2(new_n904), .ZN(new_n950));
  INV_X1    g0750(.A(KEYINPUT40), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n950), .A2(new_n951), .ZN(new_n952));
  NAND3_X1  g0752(.A1(new_n949), .A2(G330), .A3(new_n952), .ZN(new_n953));
  NOR2_X1   g0753(.A1(new_n442), .A2(new_n748), .ZN(new_n954));
  INV_X1    g0754(.A(new_n954), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n953), .A2(new_n955), .ZN(new_n956));
  XNOR2_X1  g0756(.A(new_n956), .B(KEYINPUT109), .ZN(new_n957));
  AOI22_X1  g0757(.A1(new_n948), .A2(new_n936), .B1(new_n950), .B2(new_n951), .ZN(new_n958));
  NAND3_X1  g0758(.A1(new_n958), .A2(new_n441), .A3(new_n747), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n957), .A2(new_n959), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n945), .A2(new_n960), .ZN(new_n961));
  OAI21_X1  g0761(.A(G1), .B1(new_n752), .B2(G20), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n961), .A2(new_n962), .ZN(new_n963));
  NOR2_X1   g0763(.A1(new_n945), .A2(new_n960), .ZN(new_n964));
  OAI21_X1  g0764(.A(new_n884), .B1(new_n963), .B2(new_n964), .ZN(G367));
  NOR2_X1   g0765(.A1(new_n694), .A2(new_n623), .ZN(new_n966));
  MUX2_X1   g0766(.A(new_n661), .B(new_n642), .S(new_n966), .Z(new_n967));
  NAND2_X1  g0767(.A1(new_n967), .A2(new_n770), .ZN(new_n968));
  XNOR2_X1  g0768(.A(KEYINPUT113), .B(G317), .ZN(new_n969));
  NOR2_X1   g0769(.A1(new_n791), .A2(new_n969), .ZN(new_n970));
  OAI22_X1  g0770(.A1(new_n854), .A2(new_n795), .B1(new_n784), .B2(new_n798), .ZN(new_n971));
  NOR3_X1   g0771(.A1(new_n970), .A2(new_n971), .A3(new_n445), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n808), .A2(G116), .ZN(new_n973));
  XNOR2_X1  g0773(.A(new_n973), .B(KEYINPUT46), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n807), .A2(G97), .ZN(new_n975));
  OAI22_X1  g0775(.A1(new_n778), .A2(new_n572), .B1(new_n206), .B2(new_n797), .ZN(new_n976));
  AOI21_X1  g0776(.A(new_n976), .B1(G283), .B2(new_n814), .ZN(new_n977));
  NAND4_X1  g0777(.A1(new_n972), .A2(new_n974), .A3(new_n975), .A4(new_n977), .ZN(new_n978));
  NOR2_X1   g0778(.A1(new_n797), .A2(new_n223), .ZN(new_n979));
  AOI211_X1 g0779(.A(new_n277), .B(new_n979), .C1(new_n792), .C2(G137), .ZN(new_n980));
  AOI22_X1  g0780(.A1(new_n783), .A2(new_n811), .B1(new_n814), .B2(G50), .ZN(new_n981));
  AOI22_X1  g0781(.A1(new_n779), .A2(G150), .B1(G143), .B2(new_n800), .ZN(new_n982));
  NAND3_X1  g0782(.A1(new_n980), .A2(new_n981), .A3(new_n982), .ZN(new_n983));
  INV_X1    g0783(.A(new_n808), .ZN(new_n984));
  OAI22_X1  g0784(.A1(new_n861), .A2(new_n984), .B1(new_n821), .B2(new_n229), .ZN(new_n985));
  OAI21_X1  g0785(.A(new_n978), .B1(new_n983), .B2(new_n985), .ZN(new_n986));
  XNOR2_X1  g0786(.A(new_n986), .B(KEYINPUT47), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n987), .A2(new_n771), .ZN(new_n988));
  INV_X1    g0788(.A(new_n766), .ZN(new_n989));
  OAI221_X1 g0789(.A(new_n772), .B1(new_n213), .B2(new_n342), .C1(new_n989), .C2(new_n243), .ZN(new_n990));
  NAND4_X1  g0790(.A1(new_n968), .A2(new_n757), .A3(new_n988), .A4(new_n990), .ZN(new_n991));
  INV_X1    g0791(.A(new_n699), .ZN(new_n992));
  AND3_X1   g0792(.A1(new_n685), .A2(new_n689), .A3(new_n686), .ZN(new_n993));
  AOI21_X1  g0793(.A(new_n689), .B1(new_n685), .B2(new_n686), .ZN(new_n994));
  OAI21_X1  g0794(.A(new_n692), .B1(new_n993), .B2(new_n994), .ZN(new_n995));
  INV_X1    g0795(.A(new_n683), .ZN(new_n996));
  NAND2_X1  g0796(.A1(new_n995), .A2(new_n996), .ZN(new_n997));
  OAI21_X1  g0797(.A(new_n646), .B1(new_n559), .B2(new_n694), .ZN(new_n998));
  NAND2_X1  g0798(.A1(new_n666), .A2(new_n682), .ZN(new_n999));
  AND2_X1   g0799(.A1(new_n998), .A2(new_n999), .ZN(new_n1000));
  AOI21_X1  g0800(.A(KEYINPUT44), .B1(new_n997), .B2(new_n1000), .ZN(new_n1001));
  INV_X1    g0801(.A(KEYINPUT44), .ZN(new_n1002));
  INV_X1    g0802(.A(new_n1000), .ZN(new_n1003));
  AOI211_X1 g0803(.A(new_n1002), .B(new_n1003), .C1(new_n995), .C2(new_n996), .ZN(new_n1004));
  NOR2_X1   g0804(.A1(new_n1001), .A2(new_n1004), .ZN(new_n1005));
  XOR2_X1   g0805(.A(KEYINPUT112), .B(KEYINPUT45), .Z(new_n1006));
  NAND3_X1  g0806(.A1(new_n693), .A2(new_n1003), .A3(new_n1006), .ZN(new_n1007));
  NAND3_X1  g0807(.A1(new_n995), .A2(new_n996), .A3(new_n1003), .ZN(new_n1008));
  INV_X1    g0808(.A(new_n1006), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n1008), .A2(new_n1009), .ZN(new_n1010));
  NAND2_X1  g0810(.A1(new_n1007), .A2(new_n1010), .ZN(new_n1011));
  OAI21_X1  g0811(.A(new_n992), .B1(new_n1005), .B2(new_n1011), .ZN(new_n1012));
  OAI21_X1  g0812(.A(new_n1002), .B1(new_n693), .B2(new_n1003), .ZN(new_n1013));
  NAND3_X1  g0813(.A1(new_n997), .A2(KEYINPUT44), .A3(new_n1000), .ZN(new_n1014));
  NAND2_X1  g0814(.A1(new_n1013), .A2(new_n1014), .ZN(new_n1015));
  NAND4_X1  g0815(.A1(new_n1015), .A2(new_n699), .A3(new_n1007), .A4(new_n1010), .ZN(new_n1016));
  NAND2_X1  g0816(.A1(new_n1012), .A2(new_n1016), .ZN(new_n1017));
  NOR2_X1   g0817(.A1(new_n691), .A2(new_n692), .ZN(new_n1018));
  INV_X1    g0818(.A(new_n995), .ZN(new_n1019));
  NOR2_X1   g0819(.A1(new_n1018), .A2(new_n1019), .ZN(new_n1020));
  XNOR2_X1  g0820(.A(new_n1020), .B(new_n698), .ZN(new_n1021));
  OAI21_X1  g0821(.A(new_n750), .B1(new_n1017), .B2(new_n1021), .ZN(new_n1022));
  XOR2_X1   g0822(.A(new_n703), .B(KEYINPUT41), .Z(new_n1023));
  INV_X1    g0823(.A(new_n1023), .ZN(new_n1024));
  AOI21_X1  g0824(.A(new_n756), .B1(new_n1022), .B2(new_n1024), .ZN(new_n1025));
  INV_X1    g0825(.A(KEYINPUT42), .ZN(new_n1026));
  OAI21_X1  g0826(.A(new_n1026), .B1(new_n995), .B2(new_n1000), .ZN(new_n1027));
  NAND3_X1  g0827(.A1(new_n1019), .A2(KEYINPUT42), .A3(new_n1003), .ZN(new_n1028));
  INV_X1    g0828(.A(KEYINPUT111), .ZN(new_n1029));
  OAI211_X1 g0829(.A(new_n1029), .B(new_n561), .C1(new_n1000), .C2(new_n517), .ZN(new_n1030));
  OAI21_X1  g0830(.A(new_n561), .B1(new_n1000), .B2(new_n517), .ZN(new_n1031));
  AOI21_X1  g0831(.A(new_n682), .B1(new_n1031), .B2(KEYINPUT111), .ZN(new_n1032));
  AOI22_X1  g0832(.A1(new_n1027), .A2(new_n1028), .B1(new_n1030), .B2(new_n1032), .ZN(new_n1033));
  XOR2_X1   g0833(.A(KEYINPUT110), .B(KEYINPUT43), .Z(new_n1034));
  NAND3_X1  g0834(.A1(new_n1033), .A2(new_n967), .A3(new_n1034), .ZN(new_n1035));
  MUX2_X1   g0835(.A(KEYINPUT43), .B(new_n1034), .S(new_n967), .Z(new_n1036));
  OAI21_X1  g0836(.A(new_n1035), .B1(new_n1033), .B2(new_n1036), .ZN(new_n1037));
  NAND2_X1  g0837(.A1(new_n992), .A2(new_n1003), .ZN(new_n1038));
  XNOR2_X1  g0838(.A(new_n1037), .B(new_n1038), .ZN(new_n1039));
  OAI21_X1  g0839(.A(new_n991), .B1(new_n1025), .B2(new_n1039), .ZN(G387));
  INV_X1    g0840(.A(new_n1021), .ZN(new_n1041));
  NAND2_X1  g0841(.A1(new_n750), .A2(new_n1041), .ZN(new_n1042));
  OAI21_X1  g0842(.A(new_n1021), .B1(new_n729), .B2(new_n749), .ZN(new_n1043));
  NAND3_X1  g0843(.A1(new_n1042), .A2(new_n703), .A3(new_n1043), .ZN(new_n1044));
  NAND3_X1  g0844(.A1(new_n688), .A2(new_n690), .A3(new_n770), .ZN(new_n1045));
  OAI22_X1  g0845(.A1(new_n761), .A2(new_n705), .B1(G107), .B2(new_n213), .ZN(new_n1046));
  OR2_X1    g0846(.A1(new_n240), .A2(new_n289), .ZN(new_n1047));
  INV_X1    g0847(.A(new_n705), .ZN(new_n1048));
  AOI211_X1 g0848(.A(G45), .B(new_n1048), .C1(G68), .C2(G77), .ZN(new_n1049));
  NOR2_X1   g0849(.A1(new_n257), .A2(G50), .ZN(new_n1050));
  XNOR2_X1  g0850(.A(new_n1050), .B(KEYINPUT50), .ZN(new_n1051));
  AOI21_X1  g0851(.A(new_n989), .B1(new_n1049), .B2(new_n1051), .ZN(new_n1052));
  AOI21_X1  g0852(.A(new_n1046), .B1(new_n1047), .B2(new_n1052), .ZN(new_n1053));
  OAI21_X1  g0853(.A(new_n757), .B1(new_n1053), .B2(new_n773), .ZN(new_n1054));
  AOI22_X1  g0854(.A1(G322), .A2(new_n800), .B1(new_n783), .B2(G311), .ZN(new_n1055));
  OAI221_X1 g0855(.A(new_n1055), .B1(new_n572), .B2(new_n794), .C1(new_n778), .C2(new_n969), .ZN(new_n1056));
  XNOR2_X1  g0856(.A(new_n1056), .B(KEYINPUT114), .ZN(new_n1057));
  INV_X1    g0857(.A(KEYINPUT48), .ZN(new_n1058));
  OR2_X1    g0858(.A1(new_n1057), .A2(new_n1058), .ZN(new_n1059));
  NAND2_X1  g0859(.A1(new_n1057), .A2(new_n1058), .ZN(new_n1060));
  AOI22_X1  g0860(.A1(new_n808), .A2(G294), .B1(G283), .B2(new_n816), .ZN(new_n1061));
  AND3_X1   g0861(.A1(new_n1059), .A2(new_n1060), .A3(new_n1061), .ZN(new_n1062));
  NAND2_X1  g0862(.A1(new_n1062), .A2(KEYINPUT49), .ZN(new_n1063));
  AOI21_X1  g0863(.A(new_n445), .B1(new_n792), .B2(G326), .ZN(new_n1064));
  OAI211_X1 g0864(.A(new_n1063), .B(new_n1064), .C1(new_n852), .C2(new_n821), .ZN(new_n1065));
  NOR2_X1   g0865(.A1(new_n1062), .A2(KEYINPUT49), .ZN(new_n1066));
  AOI22_X1  g0866(.A1(new_n800), .A2(G159), .B1(new_n814), .B2(G68), .ZN(new_n1067));
  INV_X1    g0867(.A(G150), .ZN(new_n1068));
  OAI211_X1 g0868(.A(new_n445), .B(new_n1067), .C1(new_n791), .C2(new_n1068), .ZN(new_n1069));
  NAND2_X1  g0869(.A1(new_n779), .A2(G50), .ZN(new_n1070));
  NAND2_X1  g0870(.A1(new_n808), .A2(G77), .ZN(new_n1071));
  AOI22_X1  g0871(.A1(new_n783), .A2(new_n258), .B1(new_n816), .B2(new_n343), .ZN(new_n1072));
  NAND4_X1  g0872(.A1(new_n1070), .A2(new_n975), .A3(new_n1071), .A4(new_n1072), .ZN(new_n1073));
  OAI22_X1  g0873(.A1(new_n1065), .A2(new_n1066), .B1(new_n1069), .B2(new_n1073), .ZN(new_n1074));
  AOI21_X1  g0874(.A(new_n1054), .B1(new_n1074), .B2(new_n771), .ZN(new_n1075));
  AOI22_X1  g0875(.A1(new_n1041), .A2(new_n756), .B1(new_n1045), .B2(new_n1075), .ZN(new_n1076));
  NAND2_X1  g0876(.A1(new_n1044), .A2(new_n1076), .ZN(G393));
  AND2_X1   g0877(.A1(new_n1012), .A2(new_n1016), .ZN(new_n1078));
  NOR3_X1   g0878(.A1(new_n729), .A2(new_n1021), .A3(new_n749), .ZN(new_n1079));
  AOI21_X1  g0879(.A(new_n704), .B1(new_n1078), .B2(new_n1079), .ZN(new_n1080));
  NAND2_X1  g0880(.A1(new_n1042), .A2(new_n1017), .ZN(new_n1081));
  NAND2_X1  g0881(.A1(new_n1080), .A2(new_n1081), .ZN(new_n1082));
  NAND3_X1  g0882(.A1(new_n1012), .A2(new_n1016), .A3(new_n756), .ZN(new_n1083));
  AND2_X1   g0883(.A1(new_n248), .A2(new_n766), .ZN(new_n1084));
  OAI21_X1  g0884(.A(new_n772), .B1(new_n205), .B2(new_n213), .ZN(new_n1085));
  OAI21_X1  g0885(.A(new_n757), .B1(new_n1084), .B2(new_n1085), .ZN(new_n1086));
  INV_X1    g0886(.A(G159), .ZN(new_n1087));
  OAI22_X1  g0887(.A1(new_n854), .A2(new_n1068), .B1(new_n778), .B2(new_n1087), .ZN(new_n1088));
  INV_X1    g0888(.A(KEYINPUT51), .ZN(new_n1089));
  AOI22_X1  g0889(.A1(new_n1088), .A2(new_n1089), .B1(G87), .B2(new_n807), .ZN(new_n1090));
  OAI221_X1 g0890(.A(new_n1090), .B1(new_n1089), .B2(new_n1088), .C1(new_n223), .C2(new_n984), .ZN(new_n1091));
  INV_X1    g0891(.A(new_n445), .ZN(new_n1092));
  AOI21_X1  g0892(.A(new_n1092), .B1(new_n792), .B2(G143), .ZN(new_n1093));
  NOR2_X1   g0893(.A1(new_n797), .A2(new_n229), .ZN(new_n1094));
  AOI21_X1  g0894(.A(new_n1094), .B1(new_n258), .B2(new_n814), .ZN(new_n1095));
  OAI211_X1 g0895(.A(new_n1093), .B(new_n1095), .C1(new_n202), .C2(new_n784), .ZN(new_n1096));
  NOR2_X1   g0896(.A1(new_n1091), .A2(new_n1096), .ZN(new_n1097));
  INV_X1    g0897(.A(new_n1097), .ZN(new_n1098));
  OR2_X1    g0898(.A1(new_n1098), .A2(KEYINPUT115), .ZN(new_n1099));
  AOI22_X1  g0899(.A1(new_n779), .A2(G311), .B1(G317), .B2(new_n800), .ZN(new_n1100));
  NOR2_X1   g0900(.A1(new_n1100), .A2(KEYINPUT52), .ZN(new_n1101));
  AOI21_X1  g0901(.A(new_n1101), .B1(G107), .B2(new_n807), .ZN(new_n1102));
  OAI21_X1  g0902(.A(new_n277), .B1(new_n794), .B2(new_n798), .ZN(new_n1103));
  OAI22_X1  g0903(.A1(new_n784), .A2(new_n572), .B1(new_n797), .B2(new_n852), .ZN(new_n1104));
  AOI211_X1 g0904(.A(new_n1103), .B(new_n1104), .C1(G322), .C2(new_n792), .ZN(new_n1105));
  AOI22_X1  g0905(.A1(new_n1100), .A2(KEYINPUT52), .B1(G283), .B2(new_n808), .ZN(new_n1106));
  NAND3_X1  g0906(.A1(new_n1102), .A2(new_n1105), .A3(new_n1106), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n1098), .A2(KEYINPUT115), .ZN(new_n1108));
  NAND3_X1  g0908(.A1(new_n1099), .A2(new_n1107), .A3(new_n1108), .ZN(new_n1109));
  AOI21_X1  g0909(.A(new_n1086), .B1(new_n1109), .B2(new_n771), .ZN(new_n1110));
  OAI21_X1  g0910(.A(new_n1110), .B1(new_n1003), .B2(new_n775), .ZN(new_n1111));
  NAND2_X1  g0911(.A1(new_n1083), .A2(new_n1111), .ZN(new_n1112));
  INV_X1    g0912(.A(new_n1112), .ZN(new_n1113));
  NAND2_X1  g0913(.A1(new_n1082), .A2(new_n1113), .ZN(G390));
  INV_X1    g0914(.A(new_n917), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n845), .A2(new_n839), .ZN(new_n1116));
  NAND2_X1  g0916(.A1(new_n1116), .A2(new_n919), .ZN(new_n1117));
  NAND3_X1  g0917(.A1(new_n845), .A2(KEYINPUT105), .A3(new_n839), .ZN(new_n1118));
  AOI21_X1  g0918(.A(new_n1115), .B1(new_n1117), .B2(new_n1118), .ZN(new_n1119));
  OAI21_X1  g0919(.A(new_n941), .B1(new_n1119), .B2(new_n942), .ZN(new_n1120));
  NAND2_X1  g0920(.A1(new_n936), .A2(new_n943), .ZN(new_n1121));
  NAND3_X1  g0921(.A1(new_n714), .A2(new_n694), .A3(new_n872), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n1122), .A2(new_n839), .ZN(new_n1123));
  AOI21_X1  g0923(.A(new_n1121), .B1(new_n917), .B2(new_n1123), .ZN(new_n1124));
  INV_X1    g0924(.A(new_n1124), .ZN(new_n1125));
  NAND4_X1  g0925(.A1(new_n747), .A2(G330), .A3(new_n872), .A4(new_n917), .ZN(new_n1126));
  NAND3_X1  g0926(.A1(new_n1120), .A2(new_n1125), .A3(new_n1126), .ZN(new_n1127));
  INV_X1    g0927(.A(new_n1126), .ZN(new_n1128));
  AOI21_X1  g0928(.A(new_n939), .B1(new_n936), .B2(new_n937), .ZN(new_n1129));
  OAI21_X1  g0929(.A(new_n917), .B1(new_n918), .B2(new_n920), .ZN(new_n1130));
  AOI21_X1  g0930(.A(new_n1129), .B1(new_n1130), .B2(new_n943), .ZN(new_n1131));
  OAI21_X1  g0931(.A(new_n1128), .B1(new_n1131), .B2(new_n1124), .ZN(new_n1132));
  NAND2_X1  g0932(.A1(new_n1127), .A2(new_n1132), .ZN(new_n1133));
  INV_X1    g0933(.A(new_n743), .ZN(new_n1134));
  NAND2_X1  g0934(.A1(new_n1134), .A2(new_n741), .ZN(new_n1135));
  NOR3_X1   g0935(.A1(new_n518), .A2(new_n634), .A3(new_n682), .ZN(new_n1136));
  OAI211_X1 g0936(.A(G330), .B(new_n872), .C1(new_n1135), .C2(new_n1136), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n1137), .A2(new_n1115), .ZN(new_n1138));
  NAND2_X1  g0938(.A1(new_n1138), .A2(new_n1126), .ZN(new_n1139));
  OAI21_X1  g0939(.A(new_n1139), .B1(new_n918), .B2(new_n920), .ZN(new_n1140));
  OAI21_X1  g0940(.A(new_n1140), .B1(new_n1123), .B2(new_n1139), .ZN(new_n1141));
  NAND3_X1  g0941(.A1(new_n888), .A2(new_n955), .A3(new_n1141), .ZN(new_n1142));
  AOI21_X1  g0942(.A(new_n704), .B1(new_n1133), .B2(new_n1142), .ZN(new_n1143));
  AOI211_X1 g0943(.A(new_n885), .B(new_n954), .C1(new_n886), .C2(new_n887), .ZN(new_n1144));
  NAND4_X1  g0944(.A1(new_n1144), .A2(new_n1127), .A3(new_n1132), .A4(new_n1141), .ZN(new_n1145));
  NAND2_X1  g0945(.A1(new_n1143), .A2(new_n1145), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n941), .A2(new_n768), .ZN(new_n1147));
  OAI21_X1  g0947(.A(new_n757), .B1(new_n258), .B2(new_n850), .ZN(new_n1148));
  NOR2_X1   g0948(.A1(new_n794), .A2(new_n205), .ZN(new_n1149));
  OAI22_X1  g0949(.A1(new_n784), .A2(new_n206), .B1(new_n778), .B2(new_n852), .ZN(new_n1150));
  AOI211_X1 g0950(.A(new_n1149), .B(new_n1150), .C1(G283), .C2(new_n800), .ZN(new_n1151));
  INV_X1    g0951(.A(new_n860), .ZN(new_n1152));
  AOI211_X1 g0952(.A(new_n352), .B(new_n1094), .C1(new_n792), .C2(G294), .ZN(new_n1153));
  NAND4_X1  g0953(.A1(new_n1151), .A2(new_n820), .A3(new_n1152), .A4(new_n1153), .ZN(new_n1154));
  NOR2_X1   g0954(.A1(new_n797), .A2(new_n1087), .ZN(new_n1155));
  OAI21_X1  g0955(.A(new_n352), .B1(new_n778), .B2(new_n862), .ZN(new_n1156));
  AOI211_X1 g0956(.A(new_n1155), .B(new_n1156), .C1(G128), .C2(new_n800), .ZN(new_n1157));
  OR3_X1    g0957(.A1(new_n984), .A2(KEYINPUT53), .A3(new_n1068), .ZN(new_n1158));
  OAI21_X1  g0958(.A(KEYINPUT53), .B1(new_n984), .B2(new_n1068), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n792), .A2(G125), .ZN(new_n1160));
  NAND4_X1  g0960(.A1(new_n1157), .A2(new_n1158), .A3(new_n1159), .A4(new_n1160), .ZN(new_n1161));
  XNOR2_X1  g0961(.A(KEYINPUT54), .B(G143), .ZN(new_n1162));
  INV_X1    g0962(.A(new_n1162), .ZN(new_n1163));
  AOI22_X1  g0963(.A1(new_n783), .A2(G137), .B1(new_n814), .B2(new_n1163), .ZN(new_n1164));
  INV_X1    g0964(.A(KEYINPUT116), .ZN(new_n1165));
  AOI22_X1  g0965(.A1(new_n1164), .A2(new_n1165), .B1(G50), .B2(new_n807), .ZN(new_n1166));
  OAI21_X1  g0966(.A(new_n1166), .B1(new_n1165), .B2(new_n1164), .ZN(new_n1167));
  OAI21_X1  g0967(.A(new_n1154), .B1(new_n1161), .B2(new_n1167), .ZN(new_n1168));
  AOI21_X1  g0968(.A(new_n1148), .B1(new_n1168), .B2(new_n771), .ZN(new_n1169));
  NAND2_X1  g0969(.A1(new_n1147), .A2(new_n1169), .ZN(new_n1170));
  INV_X1    g0970(.A(new_n756), .ZN(new_n1171));
  OAI21_X1  g0971(.A(new_n1170), .B1(new_n1133), .B2(new_n1171), .ZN(new_n1172));
  INV_X1    g0972(.A(new_n1172), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n1146), .A2(new_n1173), .ZN(G378));
  AOI21_X1  g0974(.A(new_n727), .B1(new_n830), .B2(new_n717), .ZN(new_n1175));
  INV_X1    g0975(.A(new_n728), .ZN(new_n1176));
  OAI21_X1  g0976(.A(new_n887), .B1(new_n1175), .B2(new_n1176), .ZN(new_n1177));
  NAND3_X1  g0977(.A1(new_n1177), .A2(new_n641), .A3(new_n955), .ZN(new_n1178));
  AOI21_X1  g0978(.A(new_n1126), .B1(new_n1120), .B2(new_n1125), .ZN(new_n1179));
  NOR3_X1   g0979(.A1(new_n1131), .A2(new_n1128), .A3(new_n1124), .ZN(new_n1180));
  NOR2_X1   g0980(.A1(new_n1179), .A2(new_n1180), .ZN(new_n1181));
  AOI21_X1  g0981(.A(new_n1178), .B1(new_n1181), .B2(new_n1141), .ZN(new_n1182));
  XOR2_X1   g0982(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1183));
  INV_X1    g0983(.A(new_n1183), .ZN(new_n1184));
  NOR2_X1   g0984(.A1(new_n271), .A2(new_n678), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n307), .A2(new_n1185), .ZN(new_n1186));
  INV_X1    g0986(.A(KEYINPUT119), .ZN(new_n1187));
  OAI211_X1 g0987(.A(new_n299), .B(new_n306), .C1(new_n271), .C2(new_n678), .ZN(new_n1188));
  NAND3_X1  g0988(.A1(new_n1186), .A2(new_n1187), .A3(new_n1188), .ZN(new_n1189));
  INV_X1    g0989(.A(new_n1189), .ZN(new_n1190));
  AOI21_X1  g0990(.A(new_n1187), .B1(new_n1186), .B2(new_n1188), .ZN(new_n1191));
  OAI21_X1  g0991(.A(new_n1184), .B1(new_n1190), .B2(new_n1191), .ZN(new_n1192));
  NAND2_X1  g0992(.A1(new_n1186), .A2(new_n1188), .ZN(new_n1193));
  NAND2_X1  g0993(.A1(new_n1193), .A2(KEYINPUT119), .ZN(new_n1194));
  NAND3_X1  g0994(.A1(new_n1194), .A2(new_n1189), .A3(new_n1183), .ZN(new_n1195));
  AND2_X1   g0995(.A1(new_n1192), .A2(new_n1195), .ZN(new_n1196));
  NOR2_X1   g0996(.A1(new_n953), .A2(new_n1196), .ZN(new_n1197));
  NAND2_X1  g0997(.A1(new_n1192), .A2(new_n1195), .ZN(new_n1198));
  AOI21_X1  g0998(.A(new_n1198), .B1(new_n958), .B2(G330), .ZN(new_n1199));
  OAI21_X1  g0999(.A(new_n944), .B1(new_n1197), .B2(new_n1199), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(new_n953), .A2(new_n1196), .ZN(new_n1201));
  AOI22_X1  g1001(.A1(new_n1129), .A2(new_n942), .B1(new_n922), .B2(new_n678), .ZN(new_n1202));
  NAND3_X1  g1002(.A1(new_n958), .A2(G330), .A3(new_n1198), .ZN(new_n1203));
  NAND4_X1  g1003(.A1(new_n1201), .A2(new_n1202), .A3(new_n1203), .A4(new_n921), .ZN(new_n1204));
  NAND3_X1  g1004(.A1(new_n1200), .A2(KEYINPUT57), .A3(new_n1204), .ZN(new_n1205));
  OAI21_X1  g1005(.A(new_n703), .B1(new_n1182), .B2(new_n1205), .ZN(new_n1206));
  INV_X1    g1006(.A(new_n1141), .ZN(new_n1207));
  OAI21_X1  g1007(.A(new_n1144), .B1(new_n1133), .B2(new_n1207), .ZN(new_n1208));
  AND2_X1   g1008(.A1(new_n1200), .A2(new_n1204), .ZN(new_n1209));
  AOI21_X1  g1009(.A(KEYINPUT57), .B1(new_n1208), .B2(new_n1209), .ZN(new_n1210));
  OR2_X1    g1010(.A1(new_n1206), .A2(new_n1210), .ZN(new_n1211));
  NAND2_X1  g1011(.A1(new_n1209), .A2(new_n756), .ZN(new_n1212));
  NAND2_X1  g1012(.A1(new_n807), .A2(G58), .ZN(new_n1213));
  AOI21_X1  g1013(.A(new_n979), .B1(new_n779), .B2(G107), .ZN(new_n1214));
  OAI21_X1  g1014(.A(new_n1214), .B1(new_n852), .B2(new_n854), .ZN(new_n1215));
  AOI21_X1  g1015(.A(new_n1215), .B1(G283), .B2(new_n792), .ZN(new_n1216));
  AOI22_X1  g1016(.A1(new_n783), .A2(G97), .B1(new_n814), .B2(new_n343), .ZN(new_n1217));
  XNOR2_X1  g1017(.A(new_n1217), .B(KEYINPUT117), .ZN(new_n1218));
  NAND2_X1  g1018(.A1(new_n1092), .A2(new_n288), .ZN(new_n1219));
  AOI21_X1  g1019(.A(new_n1219), .B1(G77), .B2(new_n808), .ZN(new_n1220));
  AND4_X1   g1020(.A1(new_n1213), .A2(new_n1216), .A3(new_n1218), .A4(new_n1220), .ZN(new_n1221));
  NAND2_X1  g1021(.A1(new_n1221), .A2(KEYINPUT58), .ZN(new_n1222));
  OAI211_X1 g1022(.A(new_n1219), .B(new_n202), .C1(G33), .C2(G41), .ZN(new_n1223));
  AND2_X1   g1023(.A1(new_n1222), .A2(new_n1223), .ZN(new_n1224));
  AOI22_X1  g1024(.A1(new_n800), .A2(G125), .B1(new_n816), .B2(G150), .ZN(new_n1225));
  INV_X1    g1025(.A(G128), .ZN(new_n1226));
  OAI21_X1  g1026(.A(new_n1225), .B1(new_n1226), .B2(new_n778), .ZN(new_n1227));
  AOI22_X1  g1027(.A1(new_n783), .A2(G132), .B1(new_n814), .B2(G137), .ZN(new_n1228));
  XOR2_X1   g1028(.A(new_n1228), .B(KEYINPUT118), .Z(new_n1229));
  AOI211_X1 g1029(.A(new_n1227), .B(new_n1229), .C1(new_n808), .C2(new_n1163), .ZN(new_n1230));
  INV_X1    g1030(.A(new_n1230), .ZN(new_n1231));
  NAND2_X1  g1031(.A1(new_n1231), .A2(KEYINPUT59), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(new_n807), .A2(new_n811), .ZN(new_n1233));
  AOI211_X1 g1033(.A(G33), .B(G41), .C1(new_n792), .C2(G124), .ZN(new_n1234));
  NAND3_X1  g1034(.A1(new_n1232), .A2(new_n1233), .A3(new_n1234), .ZN(new_n1235));
  NOR2_X1   g1035(.A1(new_n1231), .A2(KEYINPUT59), .ZN(new_n1236));
  OAI221_X1 g1036(.A(new_n1224), .B1(KEYINPUT58), .B2(new_n1221), .C1(new_n1235), .C2(new_n1236), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(new_n1237), .A2(new_n771), .ZN(new_n1238));
  OAI211_X1 g1038(.A(new_n1238), .B(new_n757), .C1(G50), .C2(new_n850), .ZN(new_n1239));
  AOI21_X1  g1039(.A(new_n1239), .B1(new_n1198), .B2(new_n768), .ZN(new_n1240));
  XNOR2_X1  g1040(.A(new_n1240), .B(KEYINPUT120), .ZN(new_n1241));
  AND2_X1   g1041(.A1(new_n1212), .A2(new_n1241), .ZN(new_n1242));
  NAND2_X1  g1042(.A1(new_n1211), .A2(new_n1242), .ZN(G375));
  INV_X1    g1043(.A(KEYINPUT124), .ZN(new_n1244));
  NAND2_X1  g1044(.A1(new_n1141), .A2(new_n756), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n1115), .A2(new_n768), .ZN(new_n1246));
  OAI21_X1  g1046(.A(new_n757), .B1(G68), .B2(new_n850), .ZN(new_n1247));
  AOI22_X1  g1047(.A1(new_n779), .A2(G137), .B1(new_n783), .B2(new_n1163), .ZN(new_n1248));
  OAI21_X1  g1048(.A(new_n1248), .B1(new_n862), .B2(new_n854), .ZN(new_n1249));
  XNOR2_X1  g1049(.A(new_n1249), .B(KEYINPUT123), .ZN(new_n1250));
  OAI22_X1  g1050(.A1(new_n794), .A2(new_n1068), .B1(new_n797), .B2(new_n202), .ZN(new_n1251));
  AOI211_X1 g1051(.A(new_n1092), .B(new_n1251), .C1(new_n792), .C2(G128), .ZN(new_n1252));
  OAI211_X1 g1052(.A(new_n1252), .B(new_n1213), .C1(new_n1087), .C2(new_n984), .ZN(new_n1253));
  AOI21_X1  g1053(.A(new_n352), .B1(new_n807), .B2(G77), .ZN(new_n1254));
  XNOR2_X1  g1054(.A(new_n1254), .B(KEYINPUT122), .ZN(new_n1255));
  OAI22_X1  g1055(.A1(new_n854), .A2(new_n798), .B1(new_n206), .B2(new_n794), .ZN(new_n1256));
  AOI21_X1  g1056(.A(new_n1256), .B1(G116), .B2(new_n783), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(new_n808), .A2(G97), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(new_n792), .A2(G303), .ZN(new_n1259));
  AOI22_X1  g1059(.A1(new_n779), .A2(G283), .B1(new_n343), .B2(new_n816), .ZN(new_n1260));
  NAND4_X1  g1060(.A1(new_n1257), .A2(new_n1258), .A3(new_n1259), .A4(new_n1260), .ZN(new_n1261));
  OAI22_X1  g1061(.A1(new_n1250), .A2(new_n1253), .B1(new_n1255), .B2(new_n1261), .ZN(new_n1262));
  AOI21_X1  g1062(.A(new_n1247), .B1(new_n1262), .B2(new_n771), .ZN(new_n1263));
  AND2_X1   g1063(.A1(new_n1246), .A2(new_n1263), .ZN(new_n1264));
  INV_X1    g1064(.A(new_n1264), .ZN(new_n1265));
  AOI21_X1  g1065(.A(new_n1244), .B1(new_n1245), .B2(new_n1265), .ZN(new_n1266));
  AOI211_X1 g1066(.A(KEYINPUT124), .B(new_n1264), .C1(new_n1141), .C2(new_n756), .ZN(new_n1267));
  OR2_X1    g1067(.A1(new_n1266), .A2(new_n1267), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1178), .A2(new_n1207), .ZN(new_n1269));
  XNOR2_X1  g1069(.A(new_n1023), .B(KEYINPUT121), .ZN(new_n1270));
  NAND3_X1  g1070(.A1(new_n1269), .A2(new_n1142), .A3(new_n1270), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(new_n1268), .A2(new_n1271), .ZN(G381));
  NAND3_X1  g1072(.A1(new_n1044), .A2(new_n826), .A3(new_n1076), .ZN(new_n1273));
  INV_X1    g1073(.A(new_n1273), .ZN(new_n1274));
  NAND3_X1  g1074(.A1(new_n1274), .A2(new_n1268), .A3(new_n1271), .ZN(new_n1275));
  AOI21_X1  g1075(.A(new_n1112), .B1(new_n1080), .B2(new_n1081), .ZN(new_n1276));
  INV_X1    g1076(.A(G384), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(new_n1276), .A2(new_n1277), .ZN(new_n1278));
  NOR4_X1   g1078(.A1(new_n1275), .A2(new_n1278), .A3(G378), .A4(G387), .ZN(new_n1279));
  NAND4_X1  g1079(.A1(new_n1279), .A2(new_n1241), .A3(new_n1212), .A4(new_n1211), .ZN(G407));
  AOI21_X1  g1080(.A(new_n1172), .B1(new_n1145), .B2(new_n1143), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(new_n1281), .A2(new_n679), .ZN(new_n1282));
  OAI211_X1 g1082(.A(G407), .B(G213), .C1(G375), .C2(new_n1282), .ZN(G409));
  INV_X1    g1083(.A(G213), .ZN(new_n1284));
  NOR2_X1   g1084(.A1(new_n1284), .A2(G343), .ZN(new_n1285));
  NAND2_X1  g1085(.A1(new_n1285), .A2(G2897), .ZN(new_n1286));
  INV_X1    g1086(.A(new_n1286), .ZN(new_n1287));
  INV_X1    g1087(.A(KEYINPUT60), .ZN(new_n1288));
  AOI21_X1  g1088(.A(new_n1288), .B1(new_n1269), .B2(new_n1142), .ZN(new_n1289));
  AOI21_X1  g1089(.A(new_n1141), .B1(new_n888), .B2(new_n955), .ZN(new_n1290));
  OAI21_X1  g1090(.A(new_n703), .B1(new_n1290), .B2(KEYINPUT60), .ZN(new_n1291));
  OAI21_X1  g1091(.A(new_n1268), .B1(new_n1289), .B2(new_n1291), .ZN(new_n1292));
  NAND2_X1  g1092(.A1(new_n1292), .A2(new_n1277), .ZN(new_n1293));
  INV_X1    g1093(.A(KEYINPUT125), .ZN(new_n1294));
  OAI211_X1 g1094(.A(G384), .B(new_n1268), .C1(new_n1289), .C2(new_n1291), .ZN(new_n1295));
  AND3_X1   g1095(.A1(new_n1293), .A2(new_n1294), .A3(new_n1295), .ZN(new_n1296));
  AOI21_X1  g1096(.A(new_n1294), .B1(new_n1293), .B2(new_n1295), .ZN(new_n1297));
  OAI21_X1  g1097(.A(new_n1287), .B1(new_n1296), .B2(new_n1297), .ZN(new_n1298));
  OAI211_X1 g1098(.A(G378), .B(new_n1242), .C1(new_n1206), .C2(new_n1210), .ZN(new_n1299));
  AND3_X1   g1099(.A1(new_n1208), .A2(new_n1209), .A3(new_n1270), .ZN(new_n1300));
  NAND2_X1  g1100(.A1(new_n1212), .A2(new_n1241), .ZN(new_n1301));
  OAI21_X1  g1101(.A(new_n1281), .B1(new_n1300), .B2(new_n1301), .ZN(new_n1302));
  AOI21_X1  g1102(.A(new_n1285), .B1(new_n1299), .B2(new_n1302), .ZN(new_n1303));
  INV_X1    g1103(.A(new_n1303), .ZN(new_n1304));
  NOR2_X1   g1104(.A1(new_n1178), .A2(new_n1207), .ZN(new_n1305));
  OAI21_X1  g1105(.A(KEYINPUT60), .B1(new_n1305), .B2(new_n1290), .ZN(new_n1306));
  AOI21_X1  g1106(.A(new_n704), .B1(new_n1269), .B2(new_n1288), .ZN(new_n1307));
  NAND2_X1  g1107(.A1(new_n1306), .A2(new_n1307), .ZN(new_n1308));
  AOI21_X1  g1108(.A(G384), .B1(new_n1308), .B2(new_n1268), .ZN(new_n1309));
  INV_X1    g1109(.A(new_n1295), .ZN(new_n1310));
  OAI21_X1  g1110(.A(KEYINPUT125), .B1(new_n1309), .B2(new_n1310), .ZN(new_n1311));
  NAND2_X1  g1111(.A1(new_n1311), .A2(new_n1286), .ZN(new_n1312));
  NAND3_X1  g1112(.A1(new_n1298), .A2(new_n1304), .A3(new_n1312), .ZN(new_n1313));
  INV_X1    g1113(.A(KEYINPUT61), .ZN(new_n1314));
  NAND2_X1  g1114(.A1(new_n1299), .A2(new_n1302), .ZN(new_n1315));
  INV_X1    g1115(.A(new_n1285), .ZN(new_n1316));
  NOR2_X1   g1116(.A1(new_n1309), .A2(new_n1310), .ZN(new_n1317));
  NAND3_X1  g1117(.A1(new_n1315), .A2(new_n1316), .A3(new_n1317), .ZN(new_n1318));
  NAND2_X1  g1118(.A1(new_n1318), .A2(KEYINPUT62), .ZN(new_n1319));
  INV_X1    g1119(.A(KEYINPUT62), .ZN(new_n1320));
  NAND3_X1  g1120(.A1(new_n1303), .A2(new_n1320), .A3(new_n1317), .ZN(new_n1321));
  NAND4_X1  g1121(.A1(new_n1313), .A2(new_n1314), .A3(new_n1319), .A4(new_n1321), .ZN(new_n1322));
  AOI21_X1  g1122(.A(new_n826), .B1(new_n1044), .B2(new_n1076), .ZN(new_n1323));
  NOR2_X1   g1123(.A1(new_n1274), .A2(new_n1323), .ZN(new_n1324));
  AND2_X1   g1124(.A1(G387), .A2(G390), .ZN(new_n1325));
  NOR2_X1   g1125(.A1(G387), .A2(G390), .ZN(new_n1326));
  OAI211_X1 g1126(.A(KEYINPUT127), .B(new_n1324), .C1(new_n1325), .C2(new_n1326), .ZN(new_n1327));
  INV_X1    g1127(.A(KEYINPUT127), .ZN(new_n1328));
  OAI21_X1  g1128(.A(new_n1328), .B1(new_n1274), .B2(new_n1323), .ZN(new_n1329));
  INV_X1    g1129(.A(new_n1323), .ZN(new_n1330));
  NAND3_X1  g1130(.A1(new_n1330), .A2(KEYINPUT127), .A3(new_n1273), .ZN(new_n1331));
  NAND2_X1  g1131(.A1(G387), .A2(G390), .ZN(new_n1332));
  OAI211_X1 g1132(.A(new_n1276), .B(new_n991), .C1(new_n1025), .C2(new_n1039), .ZN(new_n1333));
  NAND4_X1  g1133(.A1(new_n1329), .A2(new_n1331), .A3(new_n1332), .A4(new_n1333), .ZN(new_n1334));
  NAND2_X1  g1134(.A1(new_n1327), .A2(new_n1334), .ZN(new_n1335));
  NAND2_X1  g1135(.A1(new_n1322), .A2(new_n1335), .ZN(new_n1336));
  INV_X1    g1136(.A(KEYINPUT126), .ZN(new_n1337));
  NAND3_X1  g1137(.A1(new_n1293), .A2(new_n1294), .A3(new_n1295), .ZN(new_n1338));
  AOI21_X1  g1138(.A(new_n1286), .B1(new_n1311), .B2(new_n1338), .ZN(new_n1339));
  NOR2_X1   g1139(.A1(new_n1297), .A2(new_n1287), .ZN(new_n1340));
  OAI21_X1  g1140(.A(new_n1337), .B1(new_n1339), .B2(new_n1340), .ZN(new_n1341));
  NAND3_X1  g1141(.A1(new_n1298), .A2(KEYINPUT126), .A3(new_n1312), .ZN(new_n1342));
  NAND3_X1  g1142(.A1(new_n1341), .A2(new_n1342), .A3(new_n1304), .ZN(new_n1343));
  AND3_X1   g1143(.A1(new_n1303), .A2(KEYINPUT63), .A3(new_n1317), .ZN(new_n1344));
  AOI21_X1  g1144(.A(KEYINPUT63), .B1(new_n1303), .B2(new_n1317), .ZN(new_n1345));
  NAND3_X1  g1145(.A1(new_n1327), .A2(new_n1314), .A3(new_n1334), .ZN(new_n1346));
  NOR3_X1   g1146(.A1(new_n1344), .A2(new_n1345), .A3(new_n1346), .ZN(new_n1347));
  NAND2_X1  g1147(.A1(new_n1343), .A2(new_n1347), .ZN(new_n1348));
  NAND2_X1  g1148(.A1(new_n1336), .A2(new_n1348), .ZN(G405));
  AOI21_X1  g1149(.A(G378), .B1(new_n1211), .B2(new_n1242), .ZN(new_n1350));
  INV_X1    g1150(.A(new_n1350), .ZN(new_n1351));
  INV_X1    g1151(.A(new_n1317), .ZN(new_n1352));
  NAND3_X1  g1152(.A1(new_n1351), .A2(new_n1352), .A3(new_n1299), .ZN(new_n1353));
  INV_X1    g1153(.A(new_n1299), .ZN(new_n1354));
  OAI21_X1  g1154(.A(new_n1317), .B1(new_n1350), .B2(new_n1354), .ZN(new_n1355));
  NAND2_X1  g1155(.A1(new_n1353), .A2(new_n1355), .ZN(new_n1356));
  XNOR2_X1  g1156(.A(new_n1356), .B(new_n1335), .ZN(G402));
endmodule


