//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 0 0 1 0 1 0 0 1 0 1 0 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 0 1 0 1 1 1 0 1 1 0 1 0 1 1 1 1 0 1 0 1 1 1 1 0 1 1 0 1 1 0 1 1 1 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:20:44 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n718, new_n719, new_n720, new_n721,
    new_n723, new_n724, new_n725, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n758, new_n759,
    new_n760, new_n761, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n788, new_n789, new_n790, new_n791, new_n792,
    new_n793, new_n794, new_n796, new_n798, new_n799, new_n800, new_n801,
    new_n802, new_n803, new_n804, new_n805, new_n806, new_n807, new_n808,
    new_n809, new_n810, new_n811, new_n812, new_n813, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n825, new_n826, new_n827, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n895, new_n896, new_n898,
    new_n899, new_n900, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n912, new_n913,
    new_n914, new_n915, new_n916, new_n917, new_n918, new_n919, new_n920,
    new_n921, new_n922, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n952, new_n953, new_n954, new_n956, new_n957, new_n959,
    new_n960, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n973, new_n974, new_n976,
    new_n977, new_n978, new_n979, new_n980, new_n981, new_n982, new_n984,
    new_n985, new_n986, new_n987, new_n988, new_n990, new_n991, new_n992,
    new_n993, new_n994, new_n995, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1003, new_n1004, new_n1005, new_n1006, new_n1008,
    new_n1009, new_n1010;
  INV_X1    g000(.A(G155gat), .ZN(new_n202));
  INV_X1    g001(.A(G162gat), .ZN(new_n203));
  NAND2_X1  g002(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  NAND2_X1  g003(.A1(G155gat), .A2(G162gat), .ZN(new_n205));
  NAND2_X1  g004(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  INV_X1    g005(.A(KEYINPUT76), .ZN(new_n207));
  NAND2_X1  g006(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  NAND3_X1  g007(.A1(new_n204), .A2(KEYINPUT76), .A3(new_n205), .ZN(new_n209));
  INV_X1    g008(.A(G141gat), .ZN(new_n210));
  NAND2_X1  g009(.A1(new_n210), .A2(G148gat), .ZN(new_n211));
  INV_X1    g010(.A(G148gat), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n212), .A2(G141gat), .ZN(new_n213));
  AOI22_X1  g012(.A1(new_n211), .A2(new_n213), .B1(KEYINPUT2), .B2(new_n205), .ZN(new_n214));
  NAND3_X1  g013(.A1(new_n208), .A2(new_n209), .A3(new_n214), .ZN(new_n215));
  XNOR2_X1  g014(.A(G141gat), .B(G148gat), .ZN(new_n216));
  AND2_X1   g015(.A1(new_n205), .A2(KEYINPUT2), .ZN(new_n217));
  OAI211_X1 g016(.A(new_n207), .B(new_n206), .C1(new_n216), .C2(new_n217), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n215), .A2(new_n218), .ZN(new_n219));
  XNOR2_X1  g018(.A(G113gat), .B(G120gat), .ZN(new_n220));
  OAI211_X1 g019(.A(KEYINPUT68), .B(G134gat), .C1(new_n220), .C2(KEYINPUT1), .ZN(new_n221));
  INV_X1    g020(.A(G120gat), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n222), .A2(G113gat), .ZN(new_n223));
  INV_X1    g022(.A(G113gat), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n224), .A2(G120gat), .ZN(new_n225));
  AOI21_X1  g024(.A(KEYINPUT1), .B1(new_n223), .B2(new_n225), .ZN(new_n226));
  INV_X1    g025(.A(G134gat), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  INV_X1    g027(.A(G127gat), .ZN(new_n229));
  AND3_X1   g028(.A1(new_n221), .A2(new_n228), .A3(new_n229), .ZN(new_n230));
  AOI21_X1  g029(.A(new_n229), .B1(new_n221), .B2(new_n228), .ZN(new_n231));
  OAI21_X1  g030(.A(new_n219), .B1(new_n230), .B2(new_n231), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n232), .A2(KEYINPUT78), .ZN(new_n233));
  NAND2_X1  g032(.A1(KEYINPUT68), .A2(G134gat), .ZN(new_n234));
  NOR2_X1   g033(.A1(new_n226), .A2(new_n234), .ZN(new_n235));
  NOR3_X1   g034(.A1(new_n220), .A2(KEYINPUT1), .A3(G134gat), .ZN(new_n236));
  OAI21_X1  g035(.A(G127gat), .B1(new_n235), .B2(new_n236), .ZN(new_n237));
  NAND3_X1  g036(.A1(new_n221), .A2(new_n228), .A3(new_n229), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n237), .A2(new_n238), .ZN(new_n239));
  INV_X1    g038(.A(KEYINPUT78), .ZN(new_n240));
  NAND3_X1  g039(.A1(new_n239), .A2(new_n240), .A3(new_n219), .ZN(new_n241));
  NAND3_X1  g040(.A1(new_n233), .A2(KEYINPUT4), .A3(new_n241), .ZN(new_n242));
  XNOR2_X1  g041(.A(KEYINPUT77), .B(KEYINPUT4), .ZN(new_n243));
  NAND3_X1  g042(.A1(new_n239), .A2(new_n219), .A3(new_n243), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n242), .A2(new_n244), .ZN(new_n245));
  INV_X1    g044(.A(KEYINPUT5), .ZN(new_n246));
  INV_X1    g045(.A(new_n219), .ZN(new_n247));
  AOI21_X1  g046(.A(new_n239), .B1(KEYINPUT3), .B2(new_n247), .ZN(new_n248));
  INV_X1    g047(.A(KEYINPUT3), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n219), .A2(new_n249), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n248), .A2(new_n250), .ZN(new_n251));
  NAND2_X1  g050(.A1(G225gat), .A2(G233gat), .ZN(new_n252));
  NAND4_X1  g051(.A1(new_n245), .A2(new_n246), .A3(new_n251), .A4(new_n252), .ZN(new_n253));
  INV_X1    g052(.A(new_n252), .ZN(new_n254));
  AOI21_X1  g053(.A(new_n254), .B1(new_n248), .B2(new_n250), .ZN(new_n255));
  AOI21_X1  g054(.A(KEYINPUT4), .B1(new_n233), .B2(new_n241), .ZN(new_n256));
  AOI21_X1  g055(.A(new_n243), .B1(new_n239), .B2(new_n219), .ZN(new_n257));
  OAI21_X1  g056(.A(new_n255), .B1(new_n256), .B2(new_n257), .ZN(new_n258));
  NAND3_X1  g057(.A1(new_n247), .A2(new_n237), .A3(new_n238), .ZN(new_n259));
  NAND3_X1  g058(.A1(new_n233), .A2(new_n259), .A3(new_n241), .ZN(new_n260));
  AOI21_X1  g059(.A(new_n246), .B1(new_n260), .B2(new_n254), .ZN(new_n261));
  OAI21_X1  g060(.A(new_n258), .B1(new_n261), .B2(KEYINPUT79), .ZN(new_n262));
  INV_X1    g061(.A(KEYINPUT79), .ZN(new_n263));
  AOI211_X1 g062(.A(new_n263), .B(new_n246), .C1(new_n260), .C2(new_n254), .ZN(new_n264));
  OAI21_X1  g063(.A(new_n253), .B1(new_n262), .B2(new_n264), .ZN(new_n265));
  XNOR2_X1  g064(.A(G1gat), .B(G29gat), .ZN(new_n266));
  XNOR2_X1  g065(.A(new_n266), .B(KEYINPUT0), .ZN(new_n267));
  XNOR2_X1  g066(.A(G57gat), .B(G85gat), .ZN(new_n268));
  XOR2_X1   g067(.A(new_n267), .B(new_n268), .Z(new_n269));
  INV_X1    g068(.A(new_n269), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n265), .A2(new_n270), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n271), .A2(KEYINPUT81), .ZN(new_n272));
  OAI211_X1 g071(.A(new_n269), .B(new_n253), .C1(new_n262), .C2(new_n264), .ZN(new_n273));
  INV_X1    g072(.A(KEYINPUT6), .ZN(new_n274));
  AND2_X1   g073(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  INV_X1    g074(.A(KEYINPUT81), .ZN(new_n276));
  NAND3_X1  g075(.A1(new_n265), .A2(new_n276), .A3(new_n270), .ZN(new_n277));
  NAND3_X1  g076(.A1(new_n272), .A2(new_n275), .A3(new_n277), .ZN(new_n278));
  NAND3_X1  g077(.A1(new_n265), .A2(KEYINPUT6), .A3(new_n270), .ZN(new_n279));
  XNOR2_X1  g078(.A(G197gat), .B(G204gat), .ZN(new_n280));
  INV_X1    g079(.A(G218gat), .ZN(new_n281));
  OR2_X1    g080(.A1(KEYINPUT70), .A2(G211gat), .ZN(new_n282));
  NAND2_X1  g081(.A1(KEYINPUT70), .A2(G211gat), .ZN(new_n283));
  AOI21_X1  g082(.A(new_n281), .B1(new_n282), .B2(new_n283), .ZN(new_n284));
  OAI21_X1  g083(.A(new_n280), .B1(new_n284), .B2(KEYINPUT22), .ZN(new_n285));
  XNOR2_X1  g084(.A(G211gat), .B(G218gat), .ZN(new_n286));
  INV_X1    g085(.A(new_n286), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n285), .A2(new_n287), .ZN(new_n288));
  OAI211_X1 g087(.A(new_n280), .B(new_n286), .C1(new_n284), .C2(KEYINPUT22), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  INV_X1    g089(.A(G226gat), .ZN(new_n291));
  INV_X1    g090(.A(G233gat), .ZN(new_n292));
  NOR2_X1   g091(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  INV_X1    g092(.A(new_n293), .ZN(new_n294));
  INV_X1    g093(.A(G169gat), .ZN(new_n295));
  INV_X1    g094(.A(G176gat), .ZN(new_n296));
  NOR2_X1   g095(.A1(new_n295), .A2(new_n296), .ZN(new_n297));
  INV_X1    g096(.A(KEYINPUT26), .ZN(new_n298));
  NOR2_X1   g097(.A1(G169gat), .A2(G176gat), .ZN(new_n299));
  AOI21_X1  g098(.A(new_n297), .B1(new_n298), .B2(new_n299), .ZN(new_n300));
  INV_X1    g099(.A(KEYINPUT67), .ZN(new_n301));
  OAI21_X1  g100(.A(new_n301), .B1(new_n299), .B2(new_n298), .ZN(new_n302));
  OAI211_X1 g101(.A(KEYINPUT67), .B(KEYINPUT26), .C1(G169gat), .C2(G176gat), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n300), .A2(new_n304), .ZN(new_n305));
  INV_X1    g104(.A(G183gat), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n306), .A2(KEYINPUT27), .ZN(new_n307));
  INV_X1    g106(.A(KEYINPUT27), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n308), .A2(G183gat), .ZN(new_n309));
  INV_X1    g108(.A(G190gat), .ZN(new_n310));
  NAND3_X1  g109(.A1(new_n307), .A2(new_n309), .A3(new_n310), .ZN(new_n311));
  OR2_X1    g110(.A1(new_n311), .A2(KEYINPUT28), .ZN(new_n312));
  AOI22_X1  g111(.A1(new_n311), .A2(KEYINPUT28), .B1(G183gat), .B2(G190gat), .ZN(new_n313));
  NAND3_X1  g112(.A1(new_n305), .A2(new_n312), .A3(new_n313), .ZN(new_n314));
  OAI21_X1  g113(.A(KEYINPUT23), .B1(new_n295), .B2(new_n296), .ZN(new_n315));
  INV_X1    g114(.A(new_n299), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n315), .A2(new_n316), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n299), .A2(KEYINPUT23), .ZN(new_n318));
  NOR2_X1   g117(.A1(G183gat), .A2(G190gat), .ZN(new_n319));
  INV_X1    g118(.A(KEYINPUT66), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  NAND2_X1  g120(.A1(G183gat), .A2(G190gat), .ZN(new_n322));
  INV_X1    g121(.A(KEYINPUT24), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n321), .A2(new_n324), .ZN(new_n325));
  NAND3_X1  g124(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n326));
  OAI21_X1  g125(.A(new_n326), .B1(new_n319), .B2(new_n320), .ZN(new_n327));
  OAI211_X1 g126(.A(new_n317), .B(new_n318), .C1(new_n325), .C2(new_n327), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n328), .A2(KEYINPUT25), .ZN(new_n329));
  INV_X1    g128(.A(KEYINPUT23), .ZN(new_n330));
  NOR3_X1   g129(.A1(new_n330), .A2(G169gat), .A3(G176gat), .ZN(new_n331));
  AOI21_X1  g130(.A(new_n331), .B1(new_n316), .B2(new_n315), .ZN(new_n332));
  INV_X1    g131(.A(KEYINPUT25), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n324), .A2(KEYINPUT64), .ZN(new_n334));
  INV_X1    g133(.A(KEYINPUT64), .ZN(new_n335));
  NAND3_X1  g134(.A1(new_n322), .A2(new_n335), .A3(new_n323), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n334), .A2(new_n336), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n319), .A2(KEYINPUT65), .ZN(new_n338));
  INV_X1    g137(.A(KEYINPUT65), .ZN(new_n339));
  OAI21_X1  g138(.A(new_n339), .B1(G183gat), .B2(G190gat), .ZN(new_n340));
  NAND3_X1  g139(.A1(new_n338), .A2(new_n340), .A3(new_n326), .ZN(new_n341));
  OAI211_X1 g140(.A(new_n332), .B(new_n333), .C1(new_n337), .C2(new_n341), .ZN(new_n342));
  NAND3_X1  g141(.A1(new_n314), .A2(new_n329), .A3(new_n342), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n343), .A2(KEYINPUT71), .ZN(new_n344));
  AND2_X1   g143(.A1(new_n340), .A2(new_n326), .ZN(new_n345));
  NAND4_X1  g144(.A1(new_n345), .A2(new_n338), .A3(new_n336), .A4(new_n334), .ZN(new_n346));
  AND3_X1   g145(.A1(new_n317), .A2(new_n333), .A3(new_n318), .ZN(new_n347));
  AOI22_X1  g146(.A1(new_n346), .A2(new_n347), .B1(new_n328), .B2(KEYINPUT25), .ZN(new_n348));
  INV_X1    g147(.A(KEYINPUT71), .ZN(new_n349));
  NAND3_X1  g148(.A1(new_n348), .A2(new_n349), .A3(new_n314), .ZN(new_n350));
  AOI21_X1  g149(.A(new_n294), .B1(new_n344), .B2(new_n350), .ZN(new_n351));
  NOR2_X1   g150(.A1(new_n293), .A2(KEYINPUT29), .ZN(new_n352));
  INV_X1    g151(.A(new_n352), .ZN(new_n353));
  INV_X1    g152(.A(KEYINPUT72), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n343), .A2(new_n354), .ZN(new_n355));
  NAND3_X1  g154(.A1(new_n348), .A2(KEYINPUT72), .A3(new_n314), .ZN(new_n356));
  AOI21_X1  g155(.A(new_n353), .B1(new_n355), .B2(new_n356), .ZN(new_n357));
  OAI21_X1  g156(.A(new_n290), .B1(new_n351), .B2(new_n357), .ZN(new_n358));
  XNOR2_X1  g157(.A(G8gat), .B(G36gat), .ZN(new_n359));
  XNOR2_X1  g158(.A(new_n359), .B(KEYINPUT74), .ZN(new_n360));
  XNOR2_X1  g159(.A(G64gat), .B(G92gat), .ZN(new_n361));
  XNOR2_X1  g160(.A(new_n360), .B(new_n361), .ZN(new_n362));
  NAND3_X1  g161(.A1(new_n344), .A2(new_n350), .A3(new_n352), .ZN(new_n363));
  NAND3_X1  g162(.A1(new_n355), .A2(new_n356), .A3(new_n293), .ZN(new_n364));
  INV_X1    g163(.A(new_n290), .ZN(new_n365));
  NAND3_X1  g164(.A1(new_n363), .A2(new_n364), .A3(new_n365), .ZN(new_n366));
  NAND3_X1  g165(.A1(new_n358), .A2(new_n362), .A3(new_n366), .ZN(new_n367));
  INV_X1    g166(.A(KEYINPUT37), .ZN(new_n368));
  NAND3_X1  g167(.A1(new_n358), .A2(new_n368), .A3(new_n366), .ZN(new_n369));
  INV_X1    g168(.A(new_n362), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n369), .A2(new_n370), .ZN(new_n371));
  XOR2_X1   g170(.A(KEYINPUT82), .B(KEYINPUT38), .Z(new_n372));
  INV_X1    g171(.A(new_n351), .ZN(new_n373));
  INV_X1    g172(.A(new_n357), .ZN(new_n374));
  AOI21_X1  g173(.A(new_n290), .B1(new_n373), .B2(new_n374), .ZN(new_n375));
  NAND3_X1  g174(.A1(new_n363), .A2(new_n364), .A3(new_n290), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n376), .A2(KEYINPUT37), .ZN(new_n377));
  OAI21_X1  g176(.A(new_n372), .B1(new_n375), .B2(new_n377), .ZN(new_n378));
  OAI21_X1  g177(.A(new_n367), .B1(new_n371), .B2(new_n378), .ZN(new_n379));
  INV_X1    g178(.A(KEYINPUT73), .ZN(new_n380));
  AND3_X1   g179(.A1(new_n358), .A2(new_n380), .A3(new_n366), .ZN(new_n381));
  AOI21_X1  g180(.A(new_n380), .B1(new_n358), .B2(new_n366), .ZN(new_n382));
  OAI21_X1  g181(.A(KEYINPUT37), .B1(new_n381), .B2(new_n382), .ZN(new_n383));
  INV_X1    g182(.A(new_n371), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  INV_X1    g184(.A(new_n372), .ZN(new_n386));
  AOI21_X1  g185(.A(new_n379), .B1(new_n385), .B2(new_n386), .ZN(new_n387));
  NAND3_X1  g186(.A1(new_n278), .A2(new_n279), .A3(new_n387), .ZN(new_n388));
  AND2_X1   g187(.A1(G228gat), .A2(G233gat), .ZN(new_n389));
  INV_X1    g188(.A(new_n389), .ZN(new_n390));
  NOR2_X1   g189(.A1(new_n390), .A2(KEYINPUT80), .ZN(new_n391));
  XNOR2_X1  g190(.A(G78gat), .B(G106gat), .ZN(new_n392));
  XNOR2_X1  g191(.A(new_n391), .B(new_n392), .ZN(new_n393));
  INV_X1    g192(.A(new_n393), .ZN(new_n394));
  INV_X1    g193(.A(KEYINPUT29), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n250), .A2(new_n395), .ZN(new_n396));
  AOI22_X1  g195(.A1(new_n396), .A2(new_n365), .B1(KEYINPUT80), .B2(new_n390), .ZN(new_n397));
  INV_X1    g196(.A(G22gat), .ZN(new_n398));
  AOI21_X1  g197(.A(KEYINPUT29), .B1(new_n288), .B2(new_n289), .ZN(new_n399));
  OAI21_X1  g198(.A(new_n247), .B1(new_n399), .B2(KEYINPUT3), .ZN(new_n400));
  NAND3_X1  g199(.A1(new_n397), .A2(new_n398), .A3(new_n400), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n290), .A2(new_n395), .ZN(new_n402));
  AOI21_X1  g201(.A(new_n219), .B1(new_n402), .B2(new_n249), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n390), .A2(KEYINPUT80), .ZN(new_n404));
  AOI21_X1  g203(.A(KEYINPUT29), .B1(new_n219), .B2(new_n249), .ZN(new_n405));
  OAI21_X1  g204(.A(new_n404), .B1(new_n405), .B2(new_n290), .ZN(new_n406));
  OAI21_X1  g205(.A(G22gat), .B1(new_n403), .B2(new_n406), .ZN(new_n407));
  XNOR2_X1  g206(.A(KEYINPUT31), .B(G50gat), .ZN(new_n408));
  INV_X1    g207(.A(new_n408), .ZN(new_n409));
  AND3_X1   g208(.A1(new_n401), .A2(new_n407), .A3(new_n409), .ZN(new_n410));
  AOI21_X1  g209(.A(new_n409), .B1(new_n401), .B2(new_n407), .ZN(new_n411));
  OAI21_X1  g210(.A(new_n394), .B1(new_n410), .B2(new_n411), .ZN(new_n412));
  NAND2_X1  g211(.A1(new_n401), .A2(new_n407), .ZN(new_n413));
  NAND2_X1  g212(.A1(new_n413), .A2(new_n408), .ZN(new_n414));
  NAND3_X1  g213(.A1(new_n401), .A2(new_n407), .A3(new_n409), .ZN(new_n415));
  NAND3_X1  g214(.A1(new_n414), .A2(new_n393), .A3(new_n415), .ZN(new_n416));
  AND2_X1   g215(.A1(new_n412), .A2(new_n416), .ZN(new_n417));
  INV_X1    g216(.A(KEYINPUT40), .ZN(new_n418));
  AOI21_X1  g217(.A(new_n252), .B1(new_n245), .B2(new_n251), .ZN(new_n419));
  INV_X1    g218(.A(KEYINPUT39), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  INV_X1    g220(.A(new_n421), .ZN(new_n422));
  OAI21_X1  g221(.A(KEYINPUT39), .B1(new_n260), .B2(new_n254), .ZN(new_n423));
  OAI21_X1  g222(.A(new_n269), .B1(new_n419), .B2(new_n423), .ZN(new_n424));
  OAI21_X1  g223(.A(new_n418), .B1(new_n422), .B2(new_n424), .ZN(new_n425));
  OR2_X1    g224(.A1(new_n419), .A2(new_n423), .ZN(new_n426));
  NAND4_X1  g225(.A1(new_n426), .A2(KEYINPUT40), .A3(new_n269), .A4(new_n421), .ZN(new_n427));
  AND2_X1   g226(.A1(new_n425), .A2(new_n427), .ZN(new_n428));
  OAI21_X1  g227(.A(new_n370), .B1(new_n381), .B2(new_n382), .ZN(new_n429));
  NAND4_X1  g228(.A1(new_n358), .A2(KEYINPUT30), .A3(new_n362), .A4(new_n366), .ZN(new_n430));
  INV_X1    g229(.A(KEYINPUT75), .ZN(new_n431));
  OR2_X1    g230(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  INV_X1    g231(.A(KEYINPUT30), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n367), .A2(new_n433), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n430), .A2(new_n431), .ZN(new_n435));
  NAND4_X1  g234(.A1(new_n429), .A2(new_n432), .A3(new_n434), .A4(new_n435), .ZN(new_n436));
  NAND4_X1  g235(.A1(new_n428), .A2(new_n272), .A3(new_n277), .A4(new_n436), .ZN(new_n437));
  NAND3_X1  g236(.A1(new_n388), .A2(new_n417), .A3(new_n437), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n273), .A2(new_n274), .ZN(new_n439));
  AND2_X1   g238(.A1(new_n260), .A2(new_n254), .ZN(new_n440));
  OAI21_X1  g239(.A(new_n263), .B1(new_n440), .B2(new_n246), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n261), .A2(KEYINPUT79), .ZN(new_n442));
  NAND3_X1  g241(.A1(new_n441), .A2(new_n442), .A3(new_n258), .ZN(new_n443));
  AOI21_X1  g242(.A(new_n269), .B1(new_n443), .B2(new_n253), .ZN(new_n444));
  OAI21_X1  g243(.A(new_n279), .B1(new_n439), .B2(new_n444), .ZN(new_n445));
  INV_X1    g244(.A(new_n436), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  INV_X1    g246(.A(new_n417), .ZN(new_n448));
  INV_X1    g247(.A(KEYINPUT34), .ZN(new_n449));
  INV_X1    g248(.A(G227gat), .ZN(new_n450));
  NOR2_X1   g249(.A1(new_n450), .A2(new_n292), .ZN(new_n451));
  INV_X1    g250(.A(new_n451), .ZN(new_n452));
  AOI21_X1  g251(.A(new_n449), .B1(new_n452), .B2(KEYINPUT69), .ZN(new_n453));
  INV_X1    g252(.A(new_n453), .ZN(new_n454));
  NAND4_X1  g253(.A1(new_n348), .A2(new_n237), .A3(new_n238), .A4(new_n314), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n343), .A2(new_n239), .ZN(new_n456));
  NAND3_X1  g255(.A1(new_n455), .A2(new_n456), .A3(new_n451), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n457), .A2(KEYINPUT32), .ZN(new_n458));
  INV_X1    g257(.A(KEYINPUT33), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n457), .A2(new_n459), .ZN(new_n460));
  XOR2_X1   g259(.A(G15gat), .B(G43gat), .Z(new_n461));
  XNOR2_X1  g260(.A(G71gat), .B(G99gat), .ZN(new_n462));
  XNOR2_X1  g261(.A(new_n461), .B(new_n462), .ZN(new_n463));
  NAND3_X1  g262(.A1(new_n458), .A2(new_n460), .A3(new_n463), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n455), .A2(new_n456), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n465), .A2(new_n452), .ZN(new_n466));
  INV_X1    g265(.A(new_n463), .ZN(new_n467));
  OAI211_X1 g266(.A(new_n457), .B(KEYINPUT32), .C1(new_n459), .C2(new_n467), .ZN(new_n468));
  AND3_X1   g267(.A1(new_n464), .A2(new_n466), .A3(new_n468), .ZN(new_n469));
  AOI21_X1  g268(.A(new_n466), .B1(new_n464), .B2(new_n468), .ZN(new_n470));
  OAI21_X1  g269(.A(new_n454), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n464), .A2(new_n468), .ZN(new_n472));
  INV_X1    g271(.A(new_n466), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  NAND3_X1  g273(.A1(new_n464), .A2(new_n466), .A3(new_n468), .ZN(new_n475));
  NAND3_X1  g274(.A1(new_n474), .A2(new_n453), .A3(new_n475), .ZN(new_n476));
  NAND3_X1  g275(.A1(new_n471), .A2(new_n476), .A3(KEYINPUT36), .ZN(new_n477));
  INV_X1    g276(.A(KEYINPUT36), .ZN(new_n478));
  NOR3_X1   g277(.A1(new_n469), .A2(new_n470), .A3(new_n454), .ZN(new_n479));
  AOI21_X1  g278(.A(new_n453), .B1(new_n474), .B2(new_n475), .ZN(new_n480));
  OAI21_X1  g279(.A(new_n478), .B1(new_n479), .B2(new_n480), .ZN(new_n481));
  AOI22_X1  g280(.A1(new_n447), .A2(new_n448), .B1(new_n477), .B2(new_n481), .ZN(new_n482));
  NAND3_X1  g281(.A1(new_n417), .A2(new_n471), .A3(new_n476), .ZN(new_n483));
  INV_X1    g282(.A(new_n483), .ZN(new_n484));
  NAND3_X1  g283(.A1(new_n484), .A2(new_n445), .A3(new_n446), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n485), .A2(KEYINPUT35), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n278), .A2(new_n279), .ZN(new_n487));
  XOR2_X1   g286(.A(KEYINPUT83), .B(KEYINPUT35), .Z(new_n488));
  NOR3_X1   g287(.A1(new_n483), .A2(new_n436), .A3(new_n488), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n487), .A2(new_n489), .ZN(new_n490));
  AOI22_X1  g289(.A1(new_n438), .A2(new_n482), .B1(new_n486), .B2(new_n490), .ZN(new_n491));
  XNOR2_X1  g290(.A(G113gat), .B(G141gat), .ZN(new_n492));
  XNOR2_X1  g291(.A(new_n492), .B(G197gat), .ZN(new_n493));
  XOR2_X1   g292(.A(KEYINPUT11), .B(G169gat), .Z(new_n494));
  XNOR2_X1  g293(.A(new_n493), .B(new_n494), .ZN(new_n495));
  XOR2_X1   g294(.A(new_n495), .B(KEYINPUT12), .Z(new_n496));
  NOR2_X1   g295(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n497));
  INV_X1    g296(.A(G36gat), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  OAI21_X1  g298(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  NAND2_X1  g300(.A1(G43gat), .A2(G50gat), .ZN(new_n502));
  INV_X1    g301(.A(new_n502), .ZN(new_n503));
  NOR2_X1   g302(.A1(G43gat), .A2(G50gat), .ZN(new_n504));
  OAI21_X1  g303(.A(KEYINPUT15), .B1(new_n503), .B2(new_n504), .ZN(new_n505));
  AND2_X1   g304(.A1(KEYINPUT85), .A2(G29gat), .ZN(new_n506));
  NOR2_X1   g305(.A1(KEYINPUT85), .A2(G29gat), .ZN(new_n507));
  OAI21_X1  g306(.A(G36gat), .B1(new_n506), .B2(new_n507), .ZN(new_n508));
  INV_X1    g307(.A(G43gat), .ZN(new_n509));
  INV_X1    g308(.A(G50gat), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  INV_X1    g310(.A(KEYINPUT15), .ZN(new_n512));
  NAND3_X1  g311(.A1(new_n511), .A2(new_n512), .A3(new_n502), .ZN(new_n513));
  NAND4_X1  g312(.A1(new_n501), .A2(new_n505), .A3(new_n508), .A4(new_n513), .ZN(new_n514));
  INV_X1    g313(.A(KEYINPUT84), .ZN(new_n515));
  AOI22_X1  g314(.A1(new_n500), .A2(new_n515), .B1(new_n497), .B2(new_n498), .ZN(new_n516));
  OAI211_X1 g315(.A(KEYINPUT84), .B(KEYINPUT14), .C1(G29gat), .C2(G36gat), .ZN(new_n517));
  XNOR2_X1  g316(.A(KEYINPUT85), .B(G29gat), .ZN(new_n518));
  AOI22_X1  g317(.A1(new_n516), .A2(new_n517), .B1(G36gat), .B2(new_n518), .ZN(new_n519));
  OAI21_X1  g318(.A(new_n514), .B1(new_n519), .B2(new_n505), .ZN(new_n520));
  INV_X1    g319(.A(G1gat), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n521), .A2(KEYINPUT16), .ZN(new_n522));
  INV_X1    g321(.A(G15gat), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n523), .A2(G22gat), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n398), .A2(G15gat), .ZN(new_n525));
  NAND3_X1  g324(.A1(new_n522), .A2(new_n524), .A3(new_n525), .ZN(new_n526));
  INV_X1    g325(.A(new_n526), .ZN(new_n527));
  AOI21_X1  g326(.A(G1gat), .B1(new_n524), .B2(new_n525), .ZN(new_n528));
  OAI21_X1  g327(.A(G8gat), .B1(new_n527), .B2(new_n528), .ZN(new_n529));
  INV_X1    g328(.A(G8gat), .ZN(new_n530));
  XNOR2_X1  g329(.A(G15gat), .B(G22gat), .ZN(new_n531));
  OAI211_X1 g330(.A(new_n526), .B(new_n530), .C1(G1gat), .C2(new_n531), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n529), .A2(new_n532), .ZN(new_n533));
  AOI22_X1  g332(.A1(new_n520), .A2(new_n533), .B1(G229gat), .B2(G233gat), .ZN(new_n534));
  AND2_X1   g333(.A1(new_n534), .A2(KEYINPUT18), .ZN(new_n535));
  INV_X1    g334(.A(KEYINPUT17), .ZN(new_n536));
  OAI21_X1  g335(.A(KEYINPUT87), .B1(new_n520), .B2(new_n536), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n500), .A2(new_n515), .ZN(new_n538));
  NAND3_X1  g337(.A1(new_n538), .A2(new_n517), .A3(new_n499), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n539), .A2(new_n508), .ZN(new_n540));
  INV_X1    g339(.A(new_n505), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  INV_X1    g341(.A(KEYINPUT87), .ZN(new_n543));
  NAND4_X1  g342(.A1(new_n542), .A2(new_n543), .A3(KEYINPUT17), .A4(new_n514), .ZN(new_n544));
  INV_X1    g343(.A(KEYINPUT86), .ZN(new_n545));
  INV_X1    g344(.A(new_n514), .ZN(new_n546));
  AOI21_X1  g345(.A(new_n505), .B1(new_n539), .B2(new_n508), .ZN(new_n547));
  OAI211_X1 g346(.A(new_n545), .B(new_n536), .C1(new_n546), .C2(new_n547), .ZN(new_n548));
  INV_X1    g347(.A(new_n548), .ZN(new_n549));
  AOI21_X1  g348(.A(new_n545), .B1(new_n520), .B2(new_n536), .ZN(new_n550));
  OAI211_X1 g349(.A(new_n537), .B(new_n544), .C1(new_n549), .C2(new_n550), .ZN(new_n551));
  OAI21_X1  g350(.A(new_n535), .B1(new_n551), .B2(new_n533), .ZN(new_n552));
  NAND2_X1  g351(.A1(G229gat), .A2(G233gat), .ZN(new_n553));
  XOR2_X1   g352(.A(new_n553), .B(KEYINPUT13), .Z(new_n554));
  NOR2_X1   g353(.A1(new_n520), .A2(new_n533), .ZN(new_n555));
  AOI22_X1  g354(.A1(new_n542), .A2(new_n514), .B1(new_n529), .B2(new_n532), .ZN(new_n556));
  OAI21_X1  g355(.A(new_n554), .B1(new_n555), .B2(new_n556), .ZN(new_n557));
  INV_X1    g356(.A(KEYINPUT88), .ZN(new_n558));
  NAND2_X1  g357(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  OAI211_X1 g358(.A(KEYINPUT88), .B(new_n554), .C1(new_n555), .C2(new_n556), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n552), .A2(new_n561), .ZN(new_n562));
  OAI21_X1  g361(.A(new_n536), .B1(new_n546), .B2(new_n547), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n563), .A2(KEYINPUT86), .ZN(new_n564));
  NAND2_X1  g363(.A1(new_n564), .A2(new_n548), .ZN(new_n565));
  INV_X1    g364(.A(new_n533), .ZN(new_n566));
  NAND4_X1  g365(.A1(new_n565), .A2(new_n566), .A3(new_n537), .A4(new_n544), .ZN(new_n567));
  AOI21_X1  g366(.A(KEYINPUT18), .B1(new_n567), .B2(new_n534), .ZN(new_n568));
  OAI21_X1  g367(.A(new_n496), .B1(new_n562), .B2(new_n568), .ZN(new_n569));
  OAI21_X1  g368(.A(new_n534), .B1(new_n551), .B2(new_n533), .ZN(new_n570));
  INV_X1    g369(.A(KEYINPUT18), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  AOI22_X1  g371(.A1(new_n567), .A2(new_n535), .B1(new_n559), .B2(new_n560), .ZN(new_n573));
  INV_X1    g372(.A(new_n496), .ZN(new_n574));
  NAND3_X1  g373(.A1(new_n572), .A2(new_n573), .A3(new_n574), .ZN(new_n575));
  NAND3_X1  g374(.A1(new_n569), .A2(KEYINPUT89), .A3(new_n575), .ZN(new_n576));
  INV_X1    g375(.A(KEYINPUT89), .ZN(new_n577));
  OAI211_X1 g376(.A(new_n577), .B(new_n496), .C1(new_n562), .C2(new_n568), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n576), .A2(new_n578), .ZN(new_n579));
  NOR2_X1   g378(.A1(new_n491), .A2(new_n579), .ZN(new_n580));
  INV_X1    g379(.A(KEYINPUT98), .ZN(new_n581));
  XOR2_X1   g380(.A(G99gat), .B(G106gat), .Z(new_n582));
  INV_X1    g381(.A(new_n582), .ZN(new_n583));
  INV_X1    g382(.A(KEYINPUT8), .ZN(new_n584));
  AOI21_X1  g383(.A(new_n584), .B1(G99gat), .B2(G106gat), .ZN(new_n585));
  NOR2_X1   g384(.A1(G85gat), .A2(G92gat), .ZN(new_n586));
  OAI21_X1  g385(.A(KEYINPUT94), .B1(new_n585), .B2(new_n586), .ZN(new_n587));
  NAND2_X1  g386(.A1(G99gat), .A2(G106gat), .ZN(new_n588));
  NAND2_X1  g387(.A1(new_n588), .A2(KEYINPUT8), .ZN(new_n589));
  INV_X1    g388(.A(KEYINPUT94), .ZN(new_n590));
  INV_X1    g389(.A(G85gat), .ZN(new_n591));
  INV_X1    g390(.A(G92gat), .ZN(new_n592));
  NAND2_X1  g391(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  NAND3_X1  g392(.A1(new_n589), .A2(new_n590), .A3(new_n593), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n587), .A2(new_n594), .ZN(new_n595));
  NAND2_X1  g394(.A1(G85gat), .A2(G92gat), .ZN(new_n596));
  INV_X1    g395(.A(KEYINPUT7), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  NAND3_X1  g397(.A1(KEYINPUT7), .A2(G85gat), .A3(G92gat), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  INV_X1    g399(.A(new_n600), .ZN(new_n601));
  AOI21_X1  g400(.A(new_n583), .B1(new_n595), .B2(new_n601), .ZN(new_n602));
  AOI211_X1 g401(.A(new_n582), .B(new_n600), .C1(new_n587), .C2(new_n594), .ZN(new_n603));
  NOR2_X1   g402(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  AND2_X1   g403(.A1(G232gat), .A2(G233gat), .ZN(new_n605));
  AOI22_X1  g404(.A1(new_n604), .A2(new_n520), .B1(KEYINPUT41), .B2(new_n605), .ZN(new_n606));
  OAI21_X1  g405(.A(new_n606), .B1(new_n551), .B2(new_n604), .ZN(new_n607));
  XNOR2_X1  g406(.A(G190gat), .B(G218gat), .ZN(new_n608));
  XNOR2_X1  g407(.A(new_n608), .B(KEYINPUT95), .ZN(new_n609));
  INV_X1    g408(.A(new_n609), .ZN(new_n610));
  NAND2_X1  g409(.A1(new_n607), .A2(new_n610), .ZN(new_n611));
  OAI211_X1 g410(.A(new_n606), .B(new_n609), .C1(new_n551), .C2(new_n604), .ZN(new_n612));
  NAND3_X1  g411(.A1(new_n611), .A2(KEYINPUT96), .A3(new_n612), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n613), .A2(KEYINPUT97), .ZN(new_n614));
  INV_X1    g413(.A(KEYINPUT97), .ZN(new_n615));
  NAND4_X1  g414(.A1(new_n611), .A2(KEYINPUT96), .A3(new_n615), .A4(new_n612), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n614), .A2(new_n616), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n611), .A2(new_n612), .ZN(new_n618));
  INV_X1    g417(.A(KEYINPUT96), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  NOR2_X1   g419(.A1(new_n605), .A2(KEYINPUT41), .ZN(new_n621));
  XNOR2_X1  g420(.A(new_n621), .B(G134gat), .ZN(new_n622));
  XNOR2_X1  g421(.A(new_n622), .B(new_n203), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n620), .A2(new_n623), .ZN(new_n624));
  NAND2_X1  g423(.A1(new_n617), .A2(new_n624), .ZN(new_n625));
  INV_X1    g424(.A(new_n623), .ZN(new_n626));
  AOI21_X1  g425(.A(new_n626), .B1(new_n618), .B2(new_n619), .ZN(new_n627));
  NAND3_X1  g426(.A1(new_n627), .A2(new_n614), .A3(new_n616), .ZN(new_n628));
  NAND2_X1  g427(.A1(new_n625), .A2(new_n628), .ZN(new_n629));
  INV_X1    g428(.A(KEYINPUT90), .ZN(new_n630));
  INV_X1    g429(.A(G64gat), .ZN(new_n631));
  NOR2_X1   g430(.A1(new_n631), .A2(G57gat), .ZN(new_n632));
  INV_X1    g431(.A(G57gat), .ZN(new_n633));
  NOR2_X1   g432(.A1(new_n633), .A2(G64gat), .ZN(new_n634));
  OAI21_X1  g433(.A(new_n630), .B1(new_n632), .B2(new_n634), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n633), .A2(G64gat), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n631), .A2(G57gat), .ZN(new_n637));
  NAND3_X1  g436(.A1(new_n636), .A2(new_n637), .A3(KEYINPUT90), .ZN(new_n638));
  NAND2_X1  g437(.A1(G71gat), .A2(G78gat), .ZN(new_n639));
  INV_X1    g438(.A(KEYINPUT9), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  NAND3_X1  g440(.A1(new_n635), .A2(new_n638), .A3(new_n641), .ZN(new_n642));
  OR2_X1    g441(.A1(G71gat), .A2(G78gat), .ZN(new_n643));
  AND2_X1   g442(.A1(new_n643), .A2(new_n639), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n634), .A2(KEYINPUT91), .ZN(new_n645));
  INV_X1    g444(.A(KEYINPUT91), .ZN(new_n646));
  NAND2_X1  g445(.A1(new_n637), .A2(new_n646), .ZN(new_n647));
  NAND3_X1  g446(.A1(new_n645), .A2(new_n636), .A3(new_n647), .ZN(new_n648));
  OAI21_X1  g447(.A(new_n639), .B1(new_n643), .B2(new_n640), .ZN(new_n649));
  AOI22_X1  g448(.A1(new_n642), .A2(new_n644), .B1(new_n648), .B2(new_n649), .ZN(new_n650));
  AOI21_X1  g449(.A(new_n533), .B1(new_n650), .B2(KEYINPUT21), .ZN(new_n651));
  XNOR2_X1  g450(.A(new_n651), .B(KEYINPUT93), .ZN(new_n652));
  NOR2_X1   g451(.A1(new_n650), .A2(KEYINPUT21), .ZN(new_n653));
  XOR2_X1   g452(.A(G127gat), .B(G155gat), .Z(new_n654));
  XNOR2_X1  g453(.A(new_n653), .B(new_n654), .ZN(new_n655));
  XNOR2_X1  g454(.A(new_n652), .B(new_n655), .ZN(new_n656));
  NAND2_X1  g455(.A1(G231gat), .A2(G233gat), .ZN(new_n657));
  XNOR2_X1  g456(.A(new_n657), .B(KEYINPUT92), .ZN(new_n658));
  XOR2_X1   g457(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n659));
  XNOR2_X1  g458(.A(new_n658), .B(new_n659), .ZN(new_n660));
  XNOR2_X1  g459(.A(G183gat), .B(G211gat), .ZN(new_n661));
  XNOR2_X1  g460(.A(new_n660), .B(new_n661), .ZN(new_n662));
  XOR2_X1   g461(.A(new_n656), .B(new_n662), .Z(new_n663));
  OAI21_X1  g462(.A(new_n581), .B1(new_n629), .B2(new_n663), .ZN(new_n664));
  INV_X1    g463(.A(new_n663), .ZN(new_n665));
  NAND4_X1  g464(.A1(new_n665), .A2(KEYINPUT98), .A3(new_n628), .A4(new_n625), .ZN(new_n666));
  XNOR2_X1  g465(.A(G57gat), .B(G64gat), .ZN(new_n667));
  OAI21_X1  g466(.A(new_n641), .B1(new_n667), .B2(KEYINPUT90), .ZN(new_n668));
  INV_X1    g467(.A(new_n638), .ZN(new_n669));
  OAI21_X1  g468(.A(new_n644), .B1(new_n668), .B2(new_n669), .ZN(new_n670));
  NAND2_X1  g469(.A1(new_n648), .A2(new_n649), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  OAI21_X1  g471(.A(new_n672), .B1(new_n602), .B2(new_n603), .ZN(new_n673));
  AND3_X1   g472(.A1(new_n589), .A2(new_n590), .A3(new_n593), .ZN(new_n674));
  AOI21_X1  g473(.A(new_n590), .B1(new_n589), .B2(new_n593), .ZN(new_n675));
  OAI21_X1  g474(.A(new_n601), .B1(new_n674), .B2(new_n675), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n676), .A2(new_n582), .ZN(new_n677));
  NAND3_X1  g476(.A1(new_n595), .A2(new_n583), .A3(new_n601), .ZN(new_n678));
  NAND3_X1  g477(.A1(new_n650), .A2(new_n677), .A3(new_n678), .ZN(new_n679));
  NAND2_X1  g478(.A1(new_n673), .A2(new_n679), .ZN(new_n680));
  NAND2_X1  g479(.A1(G230gat), .A2(G233gat), .ZN(new_n681));
  INV_X1    g480(.A(new_n681), .ZN(new_n682));
  NAND2_X1  g481(.A1(new_n680), .A2(new_n682), .ZN(new_n683));
  XNOR2_X1  g482(.A(new_n683), .B(KEYINPUT99), .ZN(new_n684));
  INV_X1    g483(.A(KEYINPUT10), .ZN(new_n685));
  NAND3_X1  g484(.A1(new_n673), .A2(new_n685), .A3(new_n679), .ZN(new_n686));
  NAND3_X1  g485(.A1(new_n604), .A2(KEYINPUT10), .A3(new_n650), .ZN(new_n687));
  AOI21_X1  g486(.A(new_n682), .B1(new_n686), .B2(new_n687), .ZN(new_n688));
  XNOR2_X1  g487(.A(G120gat), .B(G148gat), .ZN(new_n689));
  XNOR2_X1  g488(.A(G176gat), .B(G204gat), .ZN(new_n690));
  XOR2_X1   g489(.A(new_n689), .B(new_n690), .Z(new_n691));
  INV_X1    g490(.A(new_n691), .ZN(new_n692));
  NOR2_X1   g491(.A1(new_n688), .A2(new_n692), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n684), .A2(new_n693), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n686), .A2(new_n687), .ZN(new_n695));
  NAND2_X1  g494(.A1(new_n695), .A2(new_n681), .ZN(new_n696));
  NAND2_X1  g495(.A1(new_n696), .A2(new_n683), .ZN(new_n697));
  NAND2_X1  g496(.A1(new_n697), .A2(new_n692), .ZN(new_n698));
  NAND2_X1  g497(.A1(new_n694), .A2(new_n698), .ZN(new_n699));
  INV_X1    g498(.A(new_n699), .ZN(new_n700));
  NAND3_X1  g499(.A1(new_n664), .A2(new_n666), .A3(new_n700), .ZN(new_n701));
  NAND2_X1  g500(.A1(new_n701), .A2(KEYINPUT100), .ZN(new_n702));
  INV_X1    g501(.A(KEYINPUT100), .ZN(new_n703));
  NAND4_X1  g502(.A1(new_n664), .A2(new_n703), .A3(new_n666), .A4(new_n700), .ZN(new_n704));
  AND2_X1   g503(.A1(new_n702), .A2(new_n704), .ZN(new_n705));
  NAND2_X1  g504(.A1(new_n580), .A2(new_n705), .ZN(new_n706));
  NOR2_X1   g505(.A1(new_n706), .A2(new_n445), .ZN(new_n707));
  XNOR2_X1  g506(.A(new_n707), .B(new_n521), .ZN(G1324gat));
  OR3_X1    g507(.A1(new_n706), .A2(KEYINPUT101), .A3(new_n446), .ZN(new_n709));
  OAI21_X1  g508(.A(KEYINPUT101), .B1(new_n706), .B2(new_n446), .ZN(new_n710));
  NAND3_X1  g509(.A1(new_n709), .A2(G8gat), .A3(new_n710), .ZN(new_n711));
  INV_X1    g510(.A(new_n706), .ZN(new_n712));
  XOR2_X1   g511(.A(KEYINPUT16), .B(G8gat), .Z(new_n713));
  NAND4_X1  g512(.A1(new_n712), .A2(KEYINPUT42), .A3(new_n436), .A4(new_n713), .ZN(new_n714));
  INV_X1    g513(.A(new_n713), .ZN(new_n715));
  AOI21_X1  g514(.A(new_n715), .B1(new_n709), .B2(new_n710), .ZN(new_n716));
  OAI211_X1 g515(.A(new_n711), .B(new_n714), .C1(new_n716), .C2(KEYINPUT42), .ZN(G1325gat));
  NAND2_X1  g516(.A1(new_n481), .A2(new_n477), .ZN(new_n718));
  OAI21_X1  g517(.A(G15gat), .B1(new_n706), .B2(new_n718), .ZN(new_n719));
  NOR2_X1   g518(.A1(new_n479), .A2(new_n480), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n720), .A2(new_n523), .ZN(new_n721));
  OAI21_X1  g520(.A(new_n719), .B1(new_n706), .B2(new_n721), .ZN(G1326gat));
  NAND2_X1  g521(.A1(new_n712), .A2(new_n448), .ZN(new_n723));
  XNOR2_X1  g522(.A(new_n723), .B(KEYINPUT102), .ZN(new_n724));
  XNOR2_X1  g523(.A(KEYINPUT43), .B(G22gat), .ZN(new_n725));
  XNOR2_X1  g524(.A(new_n724), .B(new_n725), .ZN(G1327gat));
  AND3_X1   g525(.A1(new_n627), .A2(new_n614), .A3(new_n616), .ZN(new_n727));
  AOI22_X1  g526(.A1(new_n614), .A2(new_n616), .B1(new_n620), .B2(new_n623), .ZN(new_n728));
  NOR2_X1   g527(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  NOR2_X1   g528(.A1(new_n491), .A2(new_n729), .ZN(new_n730));
  NOR3_X1   g529(.A1(new_n665), .A2(new_n579), .A3(new_n699), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  NOR3_X1   g531(.A1(new_n732), .A2(new_n445), .A3(new_n518), .ZN(new_n733));
  INV_X1    g532(.A(KEYINPUT45), .ZN(new_n734));
  XNOR2_X1  g533(.A(new_n733), .B(new_n734), .ZN(new_n735));
  INV_X1    g534(.A(KEYINPUT44), .ZN(new_n736));
  OAI21_X1  g535(.A(new_n736), .B1(new_n491), .B2(new_n729), .ZN(new_n737));
  NAND3_X1  g536(.A1(new_n271), .A2(new_n274), .A3(new_n273), .ZN(new_n738));
  AOI21_X1  g537(.A(new_n436), .B1(new_n738), .B2(new_n279), .ZN(new_n739));
  OAI21_X1  g538(.A(new_n718), .B1(new_n739), .B2(new_n417), .ZN(new_n740));
  AND3_X1   g539(.A1(new_n436), .A2(new_n425), .A3(new_n427), .ZN(new_n741));
  AND2_X1   g540(.A1(new_n272), .A2(new_n277), .ZN(new_n742));
  AOI21_X1  g541(.A(new_n448), .B1(new_n741), .B2(new_n742), .ZN(new_n743));
  AOI21_X1  g542(.A(new_n740), .B1(new_n388), .B2(new_n743), .ZN(new_n744));
  AOI22_X1  g543(.A1(KEYINPUT35), .A2(new_n485), .B1(new_n487), .B2(new_n489), .ZN(new_n745));
  OAI211_X1 g544(.A(KEYINPUT44), .B(new_n629), .C1(new_n744), .C2(new_n745), .ZN(new_n746));
  AND2_X1   g545(.A1(new_n737), .A2(new_n746), .ZN(new_n747));
  INV_X1    g546(.A(new_n445), .ZN(new_n748));
  NAND3_X1  g547(.A1(new_n747), .A2(new_n748), .A3(new_n731), .ZN(new_n749));
  NAND2_X1  g548(.A1(new_n749), .A2(KEYINPUT103), .ZN(new_n750));
  NAND2_X1  g549(.A1(new_n750), .A2(new_n518), .ZN(new_n751));
  NOR2_X1   g550(.A1(new_n749), .A2(KEYINPUT103), .ZN(new_n752));
  OAI21_X1  g551(.A(new_n735), .B1(new_n751), .B2(new_n752), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n753), .A2(KEYINPUT104), .ZN(new_n754));
  INV_X1    g553(.A(KEYINPUT104), .ZN(new_n755));
  OAI211_X1 g554(.A(new_n735), .B(new_n755), .C1(new_n751), .C2(new_n752), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n754), .A2(new_n756), .ZN(G1328gat));
  NOR3_X1   g556(.A1(new_n732), .A2(G36gat), .A3(new_n446), .ZN(new_n758));
  XNOR2_X1  g557(.A(new_n758), .B(KEYINPUT46), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n747), .A2(new_n731), .ZN(new_n760));
  OAI21_X1  g559(.A(G36gat), .B1(new_n760), .B2(new_n446), .ZN(new_n761));
  NAND2_X1  g560(.A1(new_n759), .A2(new_n761), .ZN(G1329gat));
  INV_X1    g561(.A(new_n720), .ZN(new_n763));
  OAI21_X1  g562(.A(new_n509), .B1(new_n732), .B2(new_n763), .ZN(new_n764));
  INV_X1    g563(.A(new_n718), .ZN(new_n765));
  NAND2_X1  g564(.A1(new_n765), .A2(G43gat), .ZN(new_n766));
  OAI21_X1  g565(.A(new_n764), .B1(new_n760), .B2(new_n766), .ZN(new_n767));
  XNOR2_X1  g566(.A(new_n767), .B(KEYINPUT47), .ZN(G1330gat));
  OAI21_X1  g567(.A(G50gat), .B1(new_n760), .B2(new_n417), .ZN(new_n769));
  INV_X1    g568(.A(KEYINPUT105), .ZN(new_n770));
  AOI21_X1  g569(.A(KEYINPUT48), .B1(new_n769), .B2(new_n770), .ZN(new_n771));
  NAND2_X1  g570(.A1(new_n448), .A2(new_n510), .ZN(new_n772));
  OAI21_X1  g571(.A(new_n769), .B1(new_n732), .B2(new_n772), .ZN(new_n773));
  XNOR2_X1  g572(.A(new_n771), .B(new_n773), .ZN(G1331gat));
  INV_X1    g573(.A(new_n491), .ZN(new_n775));
  AND2_X1   g574(.A1(new_n664), .A2(new_n666), .ZN(new_n776));
  AND3_X1   g575(.A1(new_n776), .A2(new_n699), .A3(new_n579), .ZN(new_n777));
  AND2_X1   g576(.A1(new_n775), .A2(new_n777), .ZN(new_n778));
  NAND2_X1  g577(.A1(new_n778), .A2(new_n748), .ZN(new_n779));
  XNOR2_X1  g578(.A(KEYINPUT106), .B(G57gat), .ZN(new_n780));
  XNOR2_X1  g579(.A(new_n779), .B(new_n780), .ZN(G1332gat));
  INV_X1    g580(.A(new_n778), .ZN(new_n782));
  NOR2_X1   g581(.A1(new_n782), .A2(new_n446), .ZN(new_n783));
  NOR2_X1   g582(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n784));
  AND2_X1   g583(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n785));
  OAI21_X1  g584(.A(new_n783), .B1(new_n784), .B2(new_n785), .ZN(new_n786));
  OAI21_X1  g585(.A(new_n786), .B1(new_n783), .B2(new_n784), .ZN(G1333gat));
  INV_X1    g586(.A(KEYINPUT107), .ZN(new_n788));
  OAI21_X1  g587(.A(new_n788), .B1(new_n782), .B2(new_n763), .ZN(new_n789));
  INV_X1    g588(.A(G71gat), .ZN(new_n790));
  NAND3_X1  g589(.A1(new_n778), .A2(KEYINPUT107), .A3(new_n720), .ZN(new_n791));
  NAND3_X1  g590(.A1(new_n789), .A2(new_n790), .A3(new_n791), .ZN(new_n792));
  NAND3_X1  g591(.A1(new_n778), .A2(G71gat), .A3(new_n765), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n792), .A2(new_n793), .ZN(new_n794));
  XNOR2_X1  g593(.A(new_n794), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g594(.A1(new_n778), .A2(new_n448), .ZN(new_n796));
  XNOR2_X1  g595(.A(new_n796), .B(G78gat), .ZN(G1335gat));
  AND2_X1   g596(.A1(new_n576), .A2(new_n578), .ZN(new_n798));
  NOR2_X1   g597(.A1(new_n665), .A2(new_n798), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n799), .A2(new_n699), .ZN(new_n800));
  XNOR2_X1  g599(.A(new_n800), .B(KEYINPUT108), .ZN(new_n801));
  NAND3_X1  g600(.A1(new_n737), .A2(new_n746), .A3(new_n801), .ZN(new_n802));
  NAND2_X1  g601(.A1(new_n802), .A2(KEYINPUT109), .ZN(new_n803));
  INV_X1    g602(.A(KEYINPUT109), .ZN(new_n804));
  NAND4_X1  g603(.A1(new_n737), .A2(new_n746), .A3(new_n804), .A4(new_n801), .ZN(new_n805));
  NAND3_X1  g604(.A1(new_n803), .A2(new_n748), .A3(new_n805), .ZN(new_n806));
  AOI21_X1  g605(.A(new_n591), .B1(new_n806), .B2(KEYINPUT110), .ZN(new_n807));
  OAI21_X1  g606(.A(new_n807), .B1(KEYINPUT110), .B2(new_n806), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n730), .A2(new_n799), .ZN(new_n809));
  OR2_X1    g608(.A1(new_n809), .A2(KEYINPUT51), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n809), .A2(KEYINPUT51), .ZN(new_n811));
  NAND3_X1  g610(.A1(new_n810), .A2(new_n699), .A3(new_n811), .ZN(new_n812));
  NAND2_X1  g611(.A1(new_n748), .A2(new_n591), .ZN(new_n813));
  OAI21_X1  g612(.A(new_n808), .B1(new_n812), .B2(new_n813), .ZN(G1336gat));
  INV_X1    g613(.A(new_n812), .ZN(new_n815));
  NOR2_X1   g614(.A1(new_n446), .A2(G92gat), .ZN(new_n816));
  NAND3_X1  g615(.A1(new_n803), .A2(new_n436), .A3(new_n805), .ZN(new_n817));
  AOI22_X1  g616(.A1(new_n815), .A2(new_n816), .B1(G92gat), .B2(new_n817), .ZN(new_n818));
  INV_X1    g617(.A(KEYINPUT52), .ZN(new_n819));
  INV_X1    g618(.A(new_n816), .ZN(new_n820));
  OAI21_X1  g619(.A(new_n819), .B1(new_n812), .B2(new_n820), .ZN(new_n821));
  INV_X1    g620(.A(new_n802), .ZN(new_n822));
  AOI21_X1  g621(.A(new_n592), .B1(new_n822), .B2(new_n436), .ZN(new_n823));
  OAI22_X1  g622(.A1(new_n818), .A2(new_n819), .B1(new_n821), .B2(new_n823), .ZN(G1337gat));
  XNOR2_X1  g623(.A(KEYINPUT111), .B(G99gat), .ZN(new_n825));
  NOR2_X1   g624(.A1(new_n763), .A2(new_n825), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n815), .A2(new_n826), .ZN(new_n827));
  NAND3_X1  g626(.A1(new_n803), .A2(new_n765), .A3(new_n805), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n828), .A2(new_n825), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n827), .A2(new_n829), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n830), .A2(KEYINPUT112), .ZN(new_n831));
  INV_X1    g630(.A(KEYINPUT112), .ZN(new_n832));
  NAND3_X1  g631(.A1(new_n827), .A2(new_n832), .A3(new_n829), .ZN(new_n833));
  NAND2_X1  g632(.A1(new_n831), .A2(new_n833), .ZN(G1338gat));
  NOR2_X1   g633(.A1(new_n417), .A2(G106gat), .ZN(new_n835));
  AND4_X1   g634(.A1(new_n699), .A2(new_n810), .A3(new_n811), .A4(new_n835), .ZN(new_n836));
  NOR2_X1   g635(.A1(new_n836), .A2(KEYINPUT53), .ZN(new_n837));
  OAI21_X1  g636(.A(G106gat), .B1(new_n802), .B2(new_n417), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n837), .A2(new_n838), .ZN(new_n839));
  NAND3_X1  g638(.A1(new_n803), .A2(new_n448), .A3(new_n805), .ZN(new_n840));
  AND3_X1   g639(.A1(new_n840), .A2(KEYINPUT113), .A3(G106gat), .ZN(new_n841));
  AOI21_X1  g640(.A(KEYINPUT113), .B1(new_n840), .B2(G106gat), .ZN(new_n842));
  NOR3_X1   g641(.A1(new_n841), .A2(new_n842), .A3(new_n836), .ZN(new_n843));
  INV_X1    g642(.A(KEYINPUT53), .ZN(new_n844));
  OAI21_X1  g643(.A(new_n839), .B1(new_n843), .B2(new_n844), .ZN(G1339gat));
  NAND3_X1  g644(.A1(new_n686), .A2(new_n687), .A3(new_n682), .ZN(new_n846));
  NAND3_X1  g645(.A1(new_n696), .A2(KEYINPUT54), .A3(new_n846), .ZN(new_n847));
  XOR2_X1   g646(.A(KEYINPUT114), .B(KEYINPUT54), .Z(new_n848));
  AOI21_X1  g647(.A(new_n691), .B1(new_n688), .B2(new_n848), .ZN(new_n849));
  NAND2_X1  g648(.A1(new_n847), .A2(new_n849), .ZN(new_n850));
  INV_X1    g649(.A(KEYINPUT55), .ZN(new_n851));
  AOI22_X1  g650(.A1(new_n850), .A2(new_n851), .B1(new_n684), .B2(new_n693), .ZN(new_n852));
  INV_X1    g651(.A(KEYINPUT115), .ZN(new_n853));
  NAND4_X1  g652(.A1(new_n847), .A2(new_n849), .A3(new_n853), .A4(KEYINPUT55), .ZN(new_n854));
  NAND3_X1  g653(.A1(new_n847), .A2(KEYINPUT55), .A3(new_n849), .ZN(new_n855));
  NAND2_X1  g654(.A1(new_n855), .A2(KEYINPUT115), .ZN(new_n856));
  NAND3_X1  g655(.A1(new_n852), .A2(new_n854), .A3(new_n856), .ZN(new_n857));
  INV_X1    g656(.A(new_n556), .ZN(new_n858));
  AOI21_X1  g657(.A(new_n553), .B1(new_n567), .B2(new_n858), .ZN(new_n859));
  NOR3_X1   g658(.A1(new_n555), .A2(new_n556), .A3(new_n554), .ZN(new_n860));
  OAI21_X1  g659(.A(new_n495), .B1(new_n859), .B2(new_n860), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n575), .A2(new_n861), .ZN(new_n862));
  NOR2_X1   g661(.A1(new_n857), .A2(new_n862), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n629), .A2(new_n863), .ZN(new_n864));
  AND3_X1   g663(.A1(new_n852), .A2(new_n854), .A3(new_n856), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n865), .A2(new_n798), .ZN(new_n866));
  NAND3_X1  g665(.A1(new_n699), .A2(new_n575), .A3(new_n861), .ZN(new_n867));
  AOI21_X1  g666(.A(KEYINPUT116), .B1(new_n866), .B2(new_n867), .ZN(new_n868));
  OAI211_X1 g667(.A(KEYINPUT116), .B(new_n867), .C1(new_n857), .C2(new_n579), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n869), .A2(new_n729), .ZN(new_n870));
  OAI21_X1  g669(.A(new_n864), .B1(new_n868), .B2(new_n870), .ZN(new_n871));
  INV_X1    g670(.A(KEYINPUT117), .ZN(new_n872));
  NAND2_X1  g671(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  OAI211_X1 g672(.A(KEYINPUT117), .B(new_n864), .C1(new_n868), .C2(new_n870), .ZN(new_n874));
  NAND3_X1  g673(.A1(new_n873), .A2(new_n663), .A3(new_n874), .ZN(new_n875));
  NAND3_X1  g674(.A1(new_n776), .A2(new_n700), .A3(new_n579), .ZN(new_n876));
  NAND2_X1  g675(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  NAND3_X1  g676(.A1(new_n877), .A2(new_n748), .A3(new_n484), .ZN(new_n878));
  INV_X1    g677(.A(KEYINPUT119), .ZN(new_n879));
  NAND2_X1  g678(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  AOI21_X1  g679(.A(new_n445), .B1(new_n875), .B2(new_n876), .ZN(new_n881));
  NAND3_X1  g680(.A1(new_n881), .A2(KEYINPUT119), .A3(new_n484), .ZN(new_n882));
  AOI21_X1  g681(.A(new_n436), .B1(new_n880), .B2(new_n882), .ZN(new_n883));
  AOI21_X1  g682(.A(G113gat), .B1(new_n883), .B2(new_n798), .ZN(new_n884));
  INV_X1    g683(.A(KEYINPUT118), .ZN(new_n885));
  AOI21_X1  g684(.A(new_n885), .B1(new_n877), .B2(new_n417), .ZN(new_n886));
  AOI211_X1 g685(.A(KEYINPUT118), .B(new_n448), .C1(new_n875), .C2(new_n876), .ZN(new_n887));
  NOR2_X1   g686(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  NAND2_X1  g687(.A1(new_n748), .A2(new_n446), .ZN(new_n889));
  NOR2_X1   g688(.A1(new_n889), .A2(new_n763), .ZN(new_n890));
  INV_X1    g689(.A(new_n890), .ZN(new_n891));
  NOR2_X1   g690(.A1(new_n888), .A2(new_n891), .ZN(new_n892));
  NOR2_X1   g691(.A1(new_n579), .A2(new_n224), .ZN(new_n893));
  AOI21_X1  g692(.A(new_n884), .B1(new_n892), .B2(new_n893), .ZN(G1340gat));
  AOI21_X1  g693(.A(G120gat), .B1(new_n883), .B2(new_n699), .ZN(new_n895));
  NOR2_X1   g694(.A1(new_n700), .A2(new_n222), .ZN(new_n896));
  AOI21_X1  g695(.A(new_n895), .B1(new_n892), .B2(new_n896), .ZN(G1341gat));
  XOR2_X1   g696(.A(KEYINPUT68), .B(G127gat), .Z(new_n898));
  INV_X1    g697(.A(new_n882), .ZN(new_n899));
  AOI21_X1  g698(.A(KEYINPUT119), .B1(new_n881), .B2(new_n484), .ZN(new_n900));
  OAI21_X1  g699(.A(new_n446), .B1(new_n899), .B2(new_n900), .ZN(new_n901));
  OAI21_X1  g700(.A(new_n898), .B1(new_n901), .B2(new_n663), .ZN(new_n902));
  NOR2_X1   g701(.A1(new_n663), .A2(new_n898), .ZN(new_n903));
  NAND2_X1  g702(.A1(new_n892), .A2(new_n903), .ZN(new_n904));
  NAND3_X1  g703(.A1(new_n902), .A2(new_n904), .A3(KEYINPUT120), .ZN(new_n905));
  INV_X1    g704(.A(KEYINPUT120), .ZN(new_n906));
  INV_X1    g705(.A(new_n898), .ZN(new_n907));
  AOI21_X1  g706(.A(new_n907), .B1(new_n883), .B2(new_n665), .ZN(new_n908));
  NOR4_X1   g707(.A1(new_n888), .A2(new_n663), .A3(new_n891), .A4(new_n898), .ZN(new_n909));
  OAI21_X1  g708(.A(new_n906), .B1(new_n908), .B2(new_n909), .ZN(new_n910));
  NAND2_X1  g709(.A1(new_n905), .A2(new_n910), .ZN(G1342gat));
  NOR2_X1   g710(.A1(new_n729), .A2(new_n436), .ZN(new_n912));
  XNOR2_X1  g711(.A(new_n912), .B(KEYINPUT121), .ZN(new_n913));
  INV_X1    g712(.A(new_n913), .ZN(new_n914));
  OAI211_X1 g713(.A(new_n227), .B(new_n914), .C1(new_n899), .C2(new_n900), .ZN(new_n915));
  XNOR2_X1  g714(.A(KEYINPUT122), .B(KEYINPUT56), .ZN(new_n916));
  OR2_X1    g715(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  NAND2_X1  g716(.A1(new_n915), .A2(new_n916), .ZN(new_n918));
  OAI211_X1 g717(.A(new_n629), .B(new_n890), .C1(new_n886), .C2(new_n887), .ZN(new_n919));
  INV_X1    g718(.A(KEYINPUT123), .ZN(new_n920));
  AND3_X1   g719(.A1(new_n919), .A2(new_n920), .A3(G134gat), .ZN(new_n921));
  AOI21_X1  g720(.A(new_n920), .B1(new_n919), .B2(G134gat), .ZN(new_n922));
  OAI211_X1 g721(.A(new_n917), .B(new_n918), .C1(new_n921), .C2(new_n922), .ZN(G1343gat));
  NOR2_X1   g722(.A1(new_n889), .A2(new_n765), .ZN(new_n924));
  INV_X1    g723(.A(new_n864), .ZN(new_n925));
  AOI21_X1  g724(.A(new_n629), .B1(new_n866), .B2(new_n867), .ZN(new_n926));
  OAI21_X1  g725(.A(new_n663), .B1(new_n925), .B2(new_n926), .ZN(new_n927));
  AOI21_X1  g726(.A(new_n417), .B1(new_n876), .B2(new_n927), .ZN(new_n928));
  INV_X1    g727(.A(KEYINPUT57), .ZN(new_n929));
  OAI21_X1  g728(.A(new_n924), .B1(new_n928), .B2(new_n929), .ZN(new_n930));
  AOI21_X1  g729(.A(new_n417), .B1(new_n875), .B2(new_n876), .ZN(new_n931));
  AOI21_X1  g730(.A(new_n930), .B1(new_n929), .B2(new_n931), .ZN(new_n932));
  AOI21_X1  g731(.A(new_n210), .B1(new_n932), .B2(new_n798), .ZN(new_n933));
  NOR2_X1   g732(.A1(new_n765), .A2(new_n417), .ZN(new_n934));
  AND2_X1   g733(.A1(new_n881), .A2(new_n934), .ZN(new_n935));
  NOR2_X1   g734(.A1(new_n579), .A2(G141gat), .ZN(new_n936));
  XNOR2_X1  g735(.A(new_n936), .B(KEYINPUT124), .ZN(new_n937));
  AND3_X1   g736(.A1(new_n935), .A2(new_n446), .A3(new_n937), .ZN(new_n938));
  NOR2_X1   g737(.A1(new_n933), .A2(new_n938), .ZN(new_n939));
  INV_X1    g738(.A(KEYINPUT58), .ZN(new_n940));
  XNOR2_X1  g739(.A(new_n939), .B(new_n940), .ZN(G1344gat));
  NAND4_X1  g740(.A1(new_n935), .A2(new_n212), .A3(new_n699), .A4(new_n446), .ZN(new_n942));
  XNOR2_X1  g741(.A(new_n942), .B(KEYINPUT125), .ZN(new_n943));
  INV_X1    g742(.A(KEYINPUT59), .ZN(new_n944));
  NAND3_X1  g743(.A1(new_n702), .A2(new_n704), .A3(new_n579), .ZN(new_n945));
  NAND2_X1  g744(.A1(new_n945), .A2(new_n927), .ZN(new_n946));
  NAND2_X1  g745(.A1(new_n946), .A2(new_n448), .ZN(new_n947));
  NAND2_X1  g746(.A1(new_n947), .A2(new_n929), .ZN(new_n948));
  AOI211_X1 g747(.A(new_n929), .B(new_n417), .C1(new_n875), .C2(new_n876), .ZN(new_n949));
  OAI21_X1  g748(.A(new_n948), .B1(new_n949), .B2(KEYINPUT126), .ZN(new_n950));
  AND3_X1   g749(.A1(new_n931), .A2(KEYINPUT126), .A3(KEYINPUT57), .ZN(new_n951));
  OAI211_X1 g750(.A(new_n699), .B(new_n924), .C1(new_n950), .C2(new_n951), .ZN(new_n952));
  AOI21_X1  g751(.A(new_n944), .B1(new_n952), .B2(G148gat), .ZN(new_n953));
  AOI211_X1 g752(.A(KEYINPUT59), .B(new_n212), .C1(new_n932), .C2(new_n699), .ZN(new_n954));
  OAI21_X1  g753(.A(new_n943), .B1(new_n953), .B2(new_n954), .ZN(G1345gat));
  NAND4_X1  g754(.A1(new_n935), .A2(new_n202), .A3(new_n665), .A4(new_n446), .ZN(new_n956));
  AND2_X1   g755(.A1(new_n932), .A2(new_n665), .ZN(new_n957));
  OAI21_X1  g756(.A(new_n956), .B1(new_n957), .B2(new_n202), .ZN(G1346gat));
  NAND3_X1  g757(.A1(new_n935), .A2(new_n203), .A3(new_n914), .ZN(new_n959));
  AND2_X1   g758(.A1(new_n932), .A2(new_n629), .ZN(new_n960));
  OAI21_X1  g759(.A(new_n959), .B1(new_n960), .B2(new_n203), .ZN(G1347gat));
  AOI21_X1  g760(.A(new_n748), .B1(new_n875), .B2(new_n876), .ZN(new_n962));
  NOR2_X1   g761(.A1(new_n446), .A2(new_n483), .ZN(new_n963));
  AND2_X1   g762(.A1(new_n962), .A2(new_n963), .ZN(new_n964));
  AOI21_X1  g763(.A(G169gat), .B1(new_n964), .B2(new_n798), .ZN(new_n965));
  NOR2_X1   g764(.A1(new_n748), .A2(new_n446), .ZN(new_n966));
  INV_X1    g765(.A(new_n966), .ZN(new_n967));
  NOR2_X1   g766(.A1(new_n967), .A2(new_n763), .ZN(new_n968));
  INV_X1    g767(.A(new_n968), .ZN(new_n969));
  NOR2_X1   g768(.A1(new_n888), .A2(new_n969), .ZN(new_n970));
  NOR2_X1   g769(.A1(new_n579), .A2(new_n295), .ZN(new_n971));
  AOI21_X1  g770(.A(new_n965), .B1(new_n970), .B2(new_n971), .ZN(G1348gat));
  NAND3_X1  g771(.A1(new_n964), .A2(new_n296), .A3(new_n699), .ZN(new_n973));
  NOR3_X1   g772(.A1(new_n888), .A2(new_n700), .A3(new_n969), .ZN(new_n974));
  OAI21_X1  g773(.A(new_n973), .B1(new_n974), .B2(new_n296), .ZN(G1349gat));
  AND3_X1   g774(.A1(new_n665), .A2(new_n307), .A3(new_n309), .ZN(new_n976));
  NAND3_X1  g775(.A1(new_n962), .A2(new_n963), .A3(new_n976), .ZN(new_n977));
  NAND2_X1  g776(.A1(KEYINPUT127), .A2(KEYINPUT60), .ZN(new_n978));
  NAND2_X1  g777(.A1(new_n977), .A2(new_n978), .ZN(new_n979));
  OAI211_X1 g778(.A(new_n665), .B(new_n968), .C1(new_n886), .C2(new_n887), .ZN(new_n980));
  AOI21_X1  g779(.A(new_n979), .B1(new_n980), .B2(G183gat), .ZN(new_n981));
  NOR2_X1   g780(.A1(KEYINPUT127), .A2(KEYINPUT60), .ZN(new_n982));
  XNOR2_X1  g781(.A(new_n981), .B(new_n982), .ZN(G1350gat));
  NAND3_X1  g782(.A1(new_n964), .A2(new_n310), .A3(new_n629), .ZN(new_n984));
  OAI211_X1 g783(.A(new_n629), .B(new_n968), .C1(new_n886), .C2(new_n887), .ZN(new_n985));
  INV_X1    g784(.A(KEYINPUT61), .ZN(new_n986));
  AND3_X1   g785(.A1(new_n985), .A2(new_n986), .A3(G190gat), .ZN(new_n987));
  AOI21_X1  g786(.A(new_n986), .B1(new_n985), .B2(G190gat), .ZN(new_n988));
  OAI21_X1  g787(.A(new_n984), .B1(new_n987), .B2(new_n988), .ZN(G1351gat));
  AND3_X1   g788(.A1(new_n962), .A2(new_n436), .A3(new_n934), .ZN(new_n990));
  AOI21_X1  g789(.A(G197gat), .B1(new_n990), .B2(new_n798), .ZN(new_n991));
  OR2_X1    g790(.A1(new_n950), .A2(new_n951), .ZN(new_n992));
  NOR2_X1   g791(.A1(new_n967), .A2(new_n765), .ZN(new_n993));
  AND2_X1   g792(.A1(new_n992), .A2(new_n993), .ZN(new_n994));
  AND2_X1   g793(.A1(new_n798), .A2(G197gat), .ZN(new_n995));
  AOI21_X1  g794(.A(new_n991), .B1(new_n994), .B2(new_n995), .ZN(G1352gat));
  NAND3_X1  g795(.A1(new_n992), .A2(new_n699), .A3(new_n993), .ZN(new_n997));
  NAND2_X1  g796(.A1(new_n997), .A2(G204gat), .ZN(new_n998));
  INV_X1    g797(.A(G204gat), .ZN(new_n999));
  NAND3_X1  g798(.A1(new_n990), .A2(new_n999), .A3(new_n699), .ZN(new_n1000));
  XOR2_X1   g799(.A(new_n1000), .B(KEYINPUT62), .Z(new_n1001));
  NAND2_X1  g800(.A1(new_n998), .A2(new_n1001), .ZN(G1353gat));
  NAND4_X1  g801(.A1(new_n990), .A2(new_n665), .A3(new_n282), .A4(new_n283), .ZN(new_n1003));
  OAI211_X1 g802(.A(new_n665), .B(new_n993), .C1(new_n950), .C2(new_n951), .ZN(new_n1004));
  AND3_X1   g803(.A1(new_n1004), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n1005));
  AOI21_X1  g804(.A(KEYINPUT63), .B1(new_n1004), .B2(G211gat), .ZN(new_n1006));
  OAI21_X1  g805(.A(new_n1003), .B1(new_n1005), .B2(new_n1006), .ZN(G1354gat));
  NAND3_X1  g806(.A1(new_n992), .A2(new_n629), .A3(new_n993), .ZN(new_n1008));
  NAND2_X1  g807(.A1(new_n1008), .A2(G218gat), .ZN(new_n1009));
  NAND3_X1  g808(.A1(new_n990), .A2(new_n281), .A3(new_n629), .ZN(new_n1010));
  NAND2_X1  g809(.A1(new_n1009), .A2(new_n1010), .ZN(G1355gat));
endmodule


