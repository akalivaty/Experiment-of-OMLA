

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
         n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706,
         n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717,
         n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
         n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739,
         n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750,
         n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761,
         n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772,
         n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783,
         n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n794,
         n795, n796, n797, n798, n799, n800, n801, n802, n803, n804, n805,
         n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n816,
         n817, n818, n819, n820, n821, n822, n823, n824, n825, n826, n827,
         n828, n829, n830, n831, n832, n833, n834, n835, n836, n837, n838,
         n839, n840, n841, n842, n843, n844, n845, n846, n847, n848, n849,
         n850, n851, n852, n853, n854, n855, n856, n857, n858, n859, n860,
         n861, n862, n863, n864, n865, n866, n867, n868, n869, n870, n871,
         n872, n873, n874, n875, n876, n877, n878, n879, n880, n881, n882,
         n883, n884, n885, n886, n887, n888, n889, n890, n891, n892, n893,
         n894, n895, n896, n897, n898, n899, n900, n901, n902, n903, n904,
         n905, n906, n907, n908, n909, n910, n911, n912, n913, n914, n915,
         n916, n917, n918, n919, n920, n921, n922, n923, n924, n925, n926,
         n927, n928, n929, n930, n931, n932, n933, n934, n935, n936, n937,
         n938, n939, n940, n941, n942, n943, n944, n945, n946, n947, n948,
         n949, n950, n951, n952, n953, n954, n955, n956, n957, n958, n959,
         n960, n961, n962, n963, n964, n965, n966, n967, n968, n969, n970,
         n971, n972, n973, n974, n975, n976, n977, n978, n979, n980, n981,
         n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, n992,
         n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003,
         n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013,
         n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023,
         n1024, n1025;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  AND2_X1 U551 ( .A1(n1009), .A2(n824), .ZN(n516) );
  XNOR2_X1 U552 ( .A(KEYINPUT102), .B(KEYINPUT30), .ZN(n719) );
  XNOR2_X1 U553 ( .A(n720), .B(n719), .ZN(n721) );
  NOR2_X1 U554 ( .A1(n716), .A2(n715), .ZN(n717) );
  AND2_X1 U555 ( .A1(n738), .A2(n737), .ZN(n739) );
  NOR2_X1 U556 ( .A1(G164), .A2(G1384), .ZN(n796) );
  INV_X1 U557 ( .A(G2104), .ZN(n521) );
  NOR2_X2 U558 ( .A1(G2105), .A2(n521), .ZN(n878) );
  NOR2_X1 U559 ( .A1(n810), .A2(n516), .ZN(n811) );
  XNOR2_X1 U560 ( .A(n522), .B(KEYINPUT65), .ZN(n884) );
  NOR2_X1 U561 ( .A1(G651), .A2(n627), .ZN(n642) );
  AND2_X1 U562 ( .A1(G2104), .A2(G2105), .ZN(n882) );
  NAND2_X1 U563 ( .A1(n882), .A2(G113), .ZN(n519) );
  NAND2_X1 U564 ( .A1(G101), .A2(n878), .ZN(n517) );
  XOR2_X1 U565 ( .A(KEYINPUT23), .B(n517), .Z(n518) );
  NAND2_X1 U566 ( .A1(n519), .A2(n518), .ZN(n526) );
  OR2_X1 U567 ( .A1(G2105), .A2(G2104), .ZN(n520) );
  XNOR2_X2 U568 ( .A(n520), .B(KEYINPUT17), .ZN(n879) );
  NAND2_X1 U569 ( .A1(G137), .A2(n879), .ZN(n524) );
  NAND2_X1 U570 ( .A1(n521), .A2(G2105), .ZN(n522) );
  NAND2_X1 U571 ( .A1(G125), .A2(n884), .ZN(n523) );
  NAND2_X1 U572 ( .A1(n524), .A2(n523), .ZN(n525) );
  NOR2_X1 U573 ( .A1(n526), .A2(n525), .ZN(G160) );
  NAND2_X1 U574 ( .A1(G114), .A2(n882), .ZN(n528) );
  NAND2_X1 U575 ( .A1(G126), .A2(n884), .ZN(n527) );
  NAND2_X1 U576 ( .A1(n528), .A2(n527), .ZN(n534) );
  NAND2_X1 U577 ( .A1(G138), .A2(n879), .ZN(n530) );
  NAND2_X1 U578 ( .A1(G102), .A2(n878), .ZN(n529) );
  NAND2_X1 U579 ( .A1(n530), .A2(n529), .ZN(n532) );
  INV_X1 U580 ( .A(KEYINPUT87), .ZN(n531) );
  XNOR2_X1 U581 ( .A(n532), .B(n531), .ZN(n533) );
  NOR2_X1 U582 ( .A1(n534), .A2(n533), .ZN(G164) );
  NOR2_X1 U583 ( .A1(G651), .A2(G543), .ZN(n633) );
  NAND2_X1 U584 ( .A1(G90), .A2(n633), .ZN(n536) );
  XOR2_X1 U585 ( .A(KEYINPUT0), .B(G543), .Z(n627) );
  XOR2_X1 U586 ( .A(G651), .B(KEYINPUT66), .Z(n538) );
  NOR2_X1 U587 ( .A1(n627), .A2(n538), .ZN(n638) );
  NAND2_X1 U588 ( .A1(G77), .A2(n638), .ZN(n535) );
  NAND2_X1 U589 ( .A1(n536), .A2(n535), .ZN(n537) );
  XNOR2_X1 U590 ( .A(KEYINPUT9), .B(n537), .ZN(n544) );
  NAND2_X1 U591 ( .A1(n642), .A2(G52), .ZN(n541) );
  NOR2_X1 U592 ( .A1(G543), .A2(n538), .ZN(n539) );
  XOR2_X1 U593 ( .A(KEYINPUT1), .B(n539), .Z(n634) );
  NAND2_X1 U594 ( .A1(G64), .A2(n634), .ZN(n540) );
  NAND2_X1 U595 ( .A1(n541), .A2(n540), .ZN(n542) );
  XOR2_X1 U596 ( .A(KEYINPUT68), .B(n542), .Z(n543) );
  NAND2_X1 U597 ( .A1(n544), .A2(n543), .ZN(G301) );
  INV_X1 U598 ( .A(G301), .ZN(G171) );
  AND2_X1 U599 ( .A1(G452), .A2(G94), .ZN(G173) );
  NAND2_X1 U600 ( .A1(G99), .A2(n878), .ZN(n546) );
  NAND2_X1 U601 ( .A1(G111), .A2(n882), .ZN(n545) );
  NAND2_X1 U602 ( .A1(n546), .A2(n545), .ZN(n549) );
  NAND2_X1 U603 ( .A1(n884), .A2(G123), .ZN(n547) );
  XOR2_X1 U604 ( .A(KEYINPUT18), .B(n547), .Z(n548) );
  NOR2_X1 U605 ( .A1(n549), .A2(n548), .ZN(n551) );
  NAND2_X1 U606 ( .A1(n879), .A2(G135), .ZN(n550) );
  NAND2_X1 U607 ( .A1(n551), .A2(n550), .ZN(n926) );
  XNOR2_X1 U608 ( .A(G2096), .B(n926), .ZN(n552) );
  OR2_X1 U609 ( .A1(G2100), .A2(n552), .ZN(G156) );
  INV_X1 U610 ( .A(G120), .ZN(G236) );
  INV_X1 U611 ( .A(G69), .ZN(G235) );
  INV_X1 U612 ( .A(G108), .ZN(G238) );
  NAND2_X1 U613 ( .A1(n642), .A2(G51), .ZN(n554) );
  NAND2_X1 U614 ( .A1(G63), .A2(n634), .ZN(n553) );
  NAND2_X1 U615 ( .A1(n554), .A2(n553), .ZN(n555) );
  XNOR2_X1 U616 ( .A(KEYINPUT6), .B(n555), .ZN(n562) );
  NAND2_X1 U617 ( .A1(n633), .A2(G89), .ZN(n556) );
  XNOR2_X1 U618 ( .A(n556), .B(KEYINPUT4), .ZN(n558) );
  NAND2_X1 U619 ( .A1(G76), .A2(n638), .ZN(n557) );
  NAND2_X1 U620 ( .A1(n558), .A2(n557), .ZN(n559) );
  XNOR2_X1 U621 ( .A(KEYINPUT5), .B(n559), .ZN(n560) );
  XNOR2_X1 U622 ( .A(KEYINPUT73), .B(n560), .ZN(n561) );
  NOR2_X1 U623 ( .A1(n562), .A2(n561), .ZN(n563) );
  XOR2_X1 U624 ( .A(KEYINPUT7), .B(n563), .Z(G168) );
  XOR2_X1 U625 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U626 ( .A1(G7), .A2(G661), .ZN(n564) );
  XNOR2_X1 U627 ( .A(n564), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U628 ( .A(G223), .ZN(n829) );
  NAND2_X1 U629 ( .A1(n829), .A2(G567), .ZN(n565) );
  XOR2_X1 U630 ( .A(KEYINPUT11), .B(n565), .Z(G234) );
  NAND2_X1 U631 ( .A1(n633), .A2(G81), .ZN(n566) );
  XNOR2_X1 U632 ( .A(n566), .B(KEYINPUT12), .ZN(n568) );
  NAND2_X1 U633 ( .A1(G68), .A2(n638), .ZN(n567) );
  NAND2_X1 U634 ( .A1(n568), .A2(n567), .ZN(n569) );
  XNOR2_X1 U635 ( .A(KEYINPUT13), .B(n569), .ZN(n575) );
  NAND2_X1 U636 ( .A1(n634), .A2(G56), .ZN(n570) );
  XOR2_X1 U637 ( .A(KEYINPUT14), .B(n570), .Z(n573) );
  NAND2_X1 U638 ( .A1(n642), .A2(G43), .ZN(n571) );
  XOR2_X1 U639 ( .A(KEYINPUT70), .B(n571), .Z(n572) );
  NOR2_X1 U640 ( .A1(n573), .A2(n572), .ZN(n574) );
  NAND2_X1 U641 ( .A1(n575), .A2(n574), .ZN(n999) );
  XNOR2_X1 U642 ( .A(G860), .B(KEYINPUT71), .ZN(n595) );
  OR2_X1 U643 ( .A1(n999), .A2(n595), .ZN(G153) );
  NAND2_X1 U644 ( .A1(G92), .A2(n633), .ZN(n577) );
  NAND2_X1 U645 ( .A1(G79), .A2(n638), .ZN(n576) );
  NAND2_X1 U646 ( .A1(n577), .A2(n576), .ZN(n581) );
  NAND2_X1 U647 ( .A1(n642), .A2(G54), .ZN(n579) );
  NAND2_X1 U648 ( .A1(G66), .A2(n634), .ZN(n578) );
  NAND2_X1 U649 ( .A1(n579), .A2(n578), .ZN(n580) );
  NOR2_X1 U650 ( .A1(n581), .A2(n580), .ZN(n582) );
  XOR2_X1 U651 ( .A(KEYINPUT15), .B(n582), .Z(n583) );
  XNOR2_X1 U652 ( .A(KEYINPUT72), .B(n583), .ZN(n700) );
  INV_X1 U653 ( .A(n700), .ZN(n1000) );
  NOR2_X1 U654 ( .A1(n1000), .A2(G868), .ZN(n585) );
  INV_X1 U655 ( .A(G868), .ZN(n645) );
  NOR2_X1 U656 ( .A1(n645), .A2(G301), .ZN(n584) );
  NOR2_X1 U657 ( .A1(n585), .A2(n584), .ZN(G284) );
  NAND2_X1 U658 ( .A1(G91), .A2(n633), .ZN(n587) );
  NAND2_X1 U659 ( .A1(G78), .A2(n638), .ZN(n586) );
  NAND2_X1 U660 ( .A1(n587), .A2(n586), .ZN(n590) );
  NAND2_X1 U661 ( .A1(G65), .A2(n634), .ZN(n588) );
  XNOR2_X1 U662 ( .A(KEYINPUT69), .B(n588), .ZN(n589) );
  NOR2_X1 U663 ( .A1(n590), .A2(n589), .ZN(n592) );
  NAND2_X1 U664 ( .A1(n642), .A2(G53), .ZN(n591) );
  NAND2_X1 U665 ( .A1(n592), .A2(n591), .ZN(G299) );
  NOR2_X1 U666 ( .A1(G286), .A2(n645), .ZN(n594) );
  NOR2_X1 U667 ( .A1(G868), .A2(G299), .ZN(n593) );
  NOR2_X1 U668 ( .A1(n594), .A2(n593), .ZN(G297) );
  NAND2_X1 U669 ( .A1(G559), .A2(n595), .ZN(n596) );
  XNOR2_X1 U670 ( .A(n596), .B(KEYINPUT74), .ZN(n597) );
  NAND2_X1 U671 ( .A1(n597), .A2(n700), .ZN(n598) );
  XNOR2_X1 U672 ( .A(KEYINPUT16), .B(n598), .ZN(G148) );
  NOR2_X1 U673 ( .A1(G868), .A2(n999), .ZN(n599) );
  XOR2_X1 U674 ( .A(KEYINPUT75), .B(n599), .Z(n602) );
  NAND2_X1 U675 ( .A1(G868), .A2(n700), .ZN(n600) );
  NOR2_X1 U676 ( .A1(G559), .A2(n600), .ZN(n601) );
  NOR2_X1 U677 ( .A1(n602), .A2(n601), .ZN(G282) );
  NAND2_X1 U678 ( .A1(G93), .A2(n633), .ZN(n603) );
  XNOR2_X1 U679 ( .A(n603), .B(KEYINPUT76), .ZN(n610) );
  NAND2_X1 U680 ( .A1(G67), .A2(n634), .ZN(n605) );
  NAND2_X1 U681 ( .A1(G80), .A2(n638), .ZN(n604) );
  NAND2_X1 U682 ( .A1(n605), .A2(n604), .ZN(n608) );
  NAND2_X1 U683 ( .A1(G55), .A2(n642), .ZN(n606) );
  XNOR2_X1 U684 ( .A(KEYINPUT77), .B(n606), .ZN(n607) );
  NOR2_X1 U685 ( .A1(n608), .A2(n607), .ZN(n609) );
  NAND2_X1 U686 ( .A1(n610), .A2(n609), .ZN(n647) );
  NAND2_X1 U687 ( .A1(G559), .A2(n700), .ZN(n656) );
  XNOR2_X1 U688 ( .A(n999), .B(n656), .ZN(n611) );
  NOR2_X1 U689 ( .A1(G860), .A2(n611), .ZN(n612) );
  XOR2_X1 U690 ( .A(n647), .B(n612), .Z(G145) );
  NAND2_X1 U691 ( .A1(G85), .A2(n633), .ZN(n614) );
  NAND2_X1 U692 ( .A1(G72), .A2(n638), .ZN(n613) );
  NAND2_X1 U693 ( .A1(n614), .A2(n613), .ZN(n617) );
  NAND2_X1 U694 ( .A1(G60), .A2(n634), .ZN(n615) );
  XNOR2_X1 U695 ( .A(KEYINPUT67), .B(n615), .ZN(n616) );
  NOR2_X1 U696 ( .A1(n617), .A2(n616), .ZN(n619) );
  NAND2_X1 U697 ( .A1(n642), .A2(G47), .ZN(n618) );
  NAND2_X1 U698 ( .A1(n619), .A2(n618), .ZN(G290) );
  NAND2_X1 U699 ( .A1(G62), .A2(n634), .ZN(n621) );
  NAND2_X1 U700 ( .A1(G75), .A2(n638), .ZN(n620) );
  NAND2_X1 U701 ( .A1(n621), .A2(n620), .ZN(n624) );
  NAND2_X1 U702 ( .A1(G88), .A2(n633), .ZN(n622) );
  XNOR2_X1 U703 ( .A(KEYINPUT79), .B(n622), .ZN(n623) );
  NOR2_X1 U704 ( .A1(n624), .A2(n623), .ZN(n626) );
  NAND2_X1 U705 ( .A1(n642), .A2(G50), .ZN(n625) );
  NAND2_X1 U706 ( .A1(n626), .A2(n625), .ZN(G303) );
  INV_X1 U707 ( .A(G303), .ZN(G166) );
  NAND2_X1 U708 ( .A1(G87), .A2(n627), .ZN(n629) );
  NAND2_X1 U709 ( .A1(G74), .A2(G651), .ZN(n628) );
  NAND2_X1 U710 ( .A1(n629), .A2(n628), .ZN(n630) );
  NOR2_X1 U711 ( .A1(n634), .A2(n630), .ZN(n632) );
  NAND2_X1 U712 ( .A1(n642), .A2(G49), .ZN(n631) );
  NAND2_X1 U713 ( .A1(n632), .A2(n631), .ZN(G288) );
  NAND2_X1 U714 ( .A1(n633), .A2(G86), .ZN(n636) );
  NAND2_X1 U715 ( .A1(G61), .A2(n634), .ZN(n635) );
  NAND2_X1 U716 ( .A1(n636), .A2(n635), .ZN(n637) );
  XNOR2_X1 U717 ( .A(KEYINPUT78), .B(n637), .ZN(n641) );
  NAND2_X1 U718 ( .A1(G73), .A2(n638), .ZN(n639) );
  XOR2_X1 U719 ( .A(KEYINPUT2), .B(n639), .Z(n640) );
  NOR2_X1 U720 ( .A1(n641), .A2(n640), .ZN(n644) );
  NAND2_X1 U721 ( .A1(n642), .A2(G48), .ZN(n643) );
  NAND2_X1 U722 ( .A1(n644), .A2(n643), .ZN(G305) );
  NAND2_X1 U723 ( .A1(n645), .A2(n647), .ZN(n646) );
  XNOR2_X1 U724 ( .A(n646), .B(KEYINPUT82), .ZN(n659) );
  INV_X1 U725 ( .A(G299), .ZN(n1005) );
  XNOR2_X1 U726 ( .A(n1005), .B(n647), .ZN(n653) );
  XOR2_X1 U727 ( .A(KEYINPUT19), .B(KEYINPUT81), .Z(n649) );
  XNOR2_X1 U728 ( .A(G166), .B(KEYINPUT80), .ZN(n648) );
  XNOR2_X1 U729 ( .A(n649), .B(n648), .ZN(n650) );
  XOR2_X1 U730 ( .A(n650), .B(G288), .Z(n651) );
  XNOR2_X1 U731 ( .A(G290), .B(n651), .ZN(n652) );
  XNOR2_X1 U732 ( .A(n653), .B(n652), .ZN(n654) );
  XNOR2_X1 U733 ( .A(n654), .B(n999), .ZN(n655) );
  XNOR2_X1 U734 ( .A(n655), .B(G305), .ZN(n894) );
  XNOR2_X1 U735 ( .A(n894), .B(n656), .ZN(n657) );
  NAND2_X1 U736 ( .A1(G868), .A2(n657), .ZN(n658) );
  NAND2_X1 U737 ( .A1(n659), .A2(n658), .ZN(n660) );
  XOR2_X1 U738 ( .A(KEYINPUT83), .B(n660), .Z(G295) );
  NAND2_X1 U739 ( .A1(G2084), .A2(G2078), .ZN(n661) );
  XOR2_X1 U740 ( .A(KEYINPUT20), .B(n661), .Z(n662) );
  NAND2_X1 U741 ( .A1(G2090), .A2(n662), .ZN(n663) );
  XNOR2_X1 U742 ( .A(KEYINPUT21), .B(n663), .ZN(n664) );
  NAND2_X1 U743 ( .A1(n664), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U744 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U745 ( .A1(G235), .A2(G236), .ZN(n665) );
  XNOR2_X1 U746 ( .A(n665), .B(KEYINPUT85), .ZN(n666) );
  NOR2_X1 U747 ( .A1(G238), .A2(n666), .ZN(n667) );
  NAND2_X1 U748 ( .A1(G57), .A2(n667), .ZN(n915) );
  NAND2_X1 U749 ( .A1(G567), .A2(n915), .ZN(n673) );
  NAND2_X1 U750 ( .A1(G132), .A2(G82), .ZN(n668) );
  XNOR2_X1 U751 ( .A(n668), .B(KEYINPUT84), .ZN(n669) );
  XNOR2_X1 U752 ( .A(n669), .B(KEYINPUT22), .ZN(n670) );
  NOR2_X1 U753 ( .A1(G218), .A2(n670), .ZN(n671) );
  NAND2_X1 U754 ( .A1(G96), .A2(n671), .ZN(n914) );
  NAND2_X1 U755 ( .A1(G2106), .A2(n914), .ZN(n672) );
  NAND2_X1 U756 ( .A1(n673), .A2(n672), .ZN(n674) );
  XOR2_X1 U757 ( .A(KEYINPUT86), .B(n674), .Z(G319) );
  INV_X1 U758 ( .A(G319), .ZN(n676) );
  NAND2_X1 U759 ( .A1(G661), .A2(G483), .ZN(n675) );
  NOR2_X1 U760 ( .A1(n676), .A2(n675), .ZN(n833) );
  NAND2_X1 U761 ( .A1(n833), .A2(G36), .ZN(G176) );
  NAND2_X1 U762 ( .A1(G160), .A2(G40), .ZN(n795) );
  XNOR2_X1 U763 ( .A(KEYINPUT95), .B(n795), .ZN(n677) );
  NAND2_X1 U764 ( .A1(n677), .A2(n796), .ZN(n678) );
  XNOR2_X1 U765 ( .A(n678), .B(KEYINPUT64), .ZN(n712) );
  NAND2_X1 U766 ( .A1(n712), .A2(G8), .ZN(n771) );
  NOR2_X1 U767 ( .A1(G1981), .A2(G305), .ZN(n679) );
  XOR2_X1 U768 ( .A(n679), .B(KEYINPUT24), .Z(n680) );
  XNOR2_X1 U769 ( .A(KEYINPUT96), .B(n680), .ZN(n681) );
  OR2_X1 U770 ( .A1(n771), .A2(n681), .ZN(n764) );
  INV_X1 U771 ( .A(n712), .ZN(n710) );
  NAND2_X1 U772 ( .A1(G2072), .A2(n710), .ZN(n682) );
  XNOR2_X1 U773 ( .A(n682), .B(KEYINPUT27), .ZN(n684) );
  AND2_X1 U774 ( .A1(n712), .A2(G1956), .ZN(n683) );
  NOR2_X1 U775 ( .A1(n684), .A2(n683), .ZN(n703) );
  NOR2_X1 U776 ( .A1(n1005), .A2(n703), .ZN(n685) );
  XOR2_X1 U777 ( .A(n685), .B(KEYINPUT28), .Z(n707) );
  NAND2_X1 U778 ( .A1(n710), .A2(G1996), .ZN(n686) );
  NAND2_X1 U779 ( .A1(n686), .A2(KEYINPUT26), .ZN(n690) );
  INV_X1 U780 ( .A(n686), .ZN(n688) );
  INV_X1 U781 ( .A(KEYINPUT26), .ZN(n687) );
  NAND2_X1 U782 ( .A1(n688), .A2(n687), .ZN(n689) );
  NAND2_X1 U783 ( .A1(n690), .A2(n689), .ZN(n692) );
  INV_X1 U784 ( .A(n710), .ZN(n731) );
  NAND2_X1 U785 ( .A1(n731), .A2(G1341), .ZN(n691) );
  NAND2_X1 U786 ( .A1(n692), .A2(n691), .ZN(n693) );
  NOR2_X1 U787 ( .A1(n999), .A2(n693), .ZN(n699) );
  NAND2_X1 U788 ( .A1(n700), .A2(n699), .ZN(n698) );
  AND2_X1 U789 ( .A1(n710), .A2(G2067), .ZN(n694) );
  XNOR2_X1 U790 ( .A(n694), .B(KEYINPUT99), .ZN(n696) );
  NAND2_X1 U791 ( .A1(n731), .A2(G1348), .ZN(n695) );
  NAND2_X1 U792 ( .A1(n696), .A2(n695), .ZN(n697) );
  NAND2_X1 U793 ( .A1(n698), .A2(n697), .ZN(n702) );
  OR2_X1 U794 ( .A1(n700), .A2(n699), .ZN(n701) );
  NAND2_X1 U795 ( .A1(n702), .A2(n701), .ZN(n705) );
  NAND2_X1 U796 ( .A1(n1005), .A2(n703), .ZN(n704) );
  NAND2_X1 U797 ( .A1(n705), .A2(n704), .ZN(n706) );
  NAND2_X1 U798 ( .A1(n707), .A2(n706), .ZN(n709) );
  XNOR2_X1 U799 ( .A(KEYINPUT29), .B(KEYINPUT100), .ZN(n708) );
  XNOR2_X1 U800 ( .A(n709), .B(n708), .ZN(n716) );
  XNOR2_X1 U801 ( .A(KEYINPUT25), .B(G2078), .ZN(n950) );
  NAND2_X1 U802 ( .A1(n710), .A2(n950), .ZN(n711) );
  XNOR2_X1 U803 ( .A(n711), .B(KEYINPUT98), .ZN(n714) );
  INV_X1 U804 ( .A(G1961), .ZN(n967) );
  NAND2_X1 U805 ( .A1(n712), .A2(n967), .ZN(n713) );
  NAND2_X1 U806 ( .A1(n714), .A2(n713), .ZN(n722) );
  AND2_X1 U807 ( .A1(n722), .A2(G171), .ZN(n715) );
  XNOR2_X1 U808 ( .A(n717), .B(KEYINPUT101), .ZN(n728) );
  NOR2_X1 U809 ( .A1(G1966), .A2(n771), .ZN(n743) );
  NOR2_X1 U810 ( .A1(n731), .A2(G2084), .ZN(n740) );
  NOR2_X1 U811 ( .A1(n743), .A2(n740), .ZN(n718) );
  NAND2_X1 U812 ( .A1(G8), .A2(n718), .ZN(n720) );
  NOR2_X1 U813 ( .A1(G168), .A2(n721), .ZN(n724) );
  NOR2_X1 U814 ( .A1(G171), .A2(n722), .ZN(n723) );
  NOR2_X1 U815 ( .A1(n724), .A2(n723), .ZN(n725) );
  XNOR2_X1 U816 ( .A(n725), .B(KEYINPUT103), .ZN(n726) );
  XNOR2_X1 U817 ( .A(n726), .B(KEYINPUT31), .ZN(n727) );
  NAND2_X1 U818 ( .A1(n728), .A2(n727), .ZN(n742) );
  AND2_X1 U819 ( .A1(G286), .A2(G8), .ZN(n729) );
  NAND2_X1 U820 ( .A1(n742), .A2(n729), .ZN(n738) );
  INV_X1 U821 ( .A(G8), .ZN(n736) );
  NOR2_X1 U822 ( .A1(G1971), .A2(n771), .ZN(n730) );
  XNOR2_X1 U823 ( .A(n730), .B(KEYINPUT104), .ZN(n733) );
  NOR2_X1 U824 ( .A1(n731), .A2(G2090), .ZN(n732) );
  NOR2_X1 U825 ( .A1(n733), .A2(n732), .ZN(n734) );
  NAND2_X1 U826 ( .A1(n734), .A2(G303), .ZN(n735) );
  OR2_X1 U827 ( .A1(n736), .A2(n735), .ZN(n737) );
  XNOR2_X1 U828 ( .A(n739), .B(KEYINPUT32), .ZN(n766) );
  NAND2_X1 U829 ( .A1(G8), .A2(n740), .ZN(n741) );
  XOR2_X1 U830 ( .A(KEYINPUT97), .B(n741), .Z(n746) );
  INV_X1 U831 ( .A(n742), .ZN(n744) );
  NOR2_X1 U832 ( .A1(n744), .A2(n743), .ZN(n745) );
  NAND2_X1 U833 ( .A1(n746), .A2(n745), .ZN(n765) );
  NAND2_X1 U834 ( .A1(G1976), .A2(G288), .ZN(n1011) );
  AND2_X1 U835 ( .A1(n765), .A2(n1011), .ZN(n747) );
  NAND2_X1 U836 ( .A1(n766), .A2(n747), .ZN(n753) );
  INV_X1 U837 ( .A(n1011), .ZN(n751) );
  NOR2_X1 U838 ( .A1(G1976), .A2(G288), .ZN(n748) );
  XOR2_X1 U839 ( .A(KEYINPUT105), .B(n748), .Z(n754) );
  NOR2_X1 U840 ( .A1(G1971), .A2(G303), .ZN(n749) );
  NOR2_X1 U841 ( .A1(n754), .A2(n749), .ZN(n750) );
  OR2_X1 U842 ( .A1(n751), .A2(n750), .ZN(n752) );
  AND2_X1 U843 ( .A1(n753), .A2(n752), .ZN(n758) );
  INV_X1 U844 ( .A(n754), .ZN(n1012) );
  NOR2_X1 U845 ( .A1(n771), .A2(n1012), .ZN(n755) );
  AND2_X1 U846 ( .A1(KEYINPUT33), .A2(n755), .ZN(n756) );
  XNOR2_X1 U847 ( .A(G1981), .B(G305), .ZN(n996) );
  OR2_X1 U848 ( .A1(n756), .A2(n996), .ZN(n759) );
  OR2_X1 U849 ( .A1(n771), .A2(n759), .ZN(n757) );
  NOR2_X1 U850 ( .A1(n758), .A2(n757), .ZN(n762) );
  INV_X1 U851 ( .A(n759), .ZN(n760) );
  AND2_X1 U852 ( .A1(n760), .A2(KEYINPUT33), .ZN(n761) );
  NOR2_X1 U853 ( .A1(n762), .A2(n761), .ZN(n763) );
  NAND2_X1 U854 ( .A1(n764), .A2(n763), .ZN(n774) );
  NAND2_X1 U855 ( .A1(n766), .A2(n765), .ZN(n769) );
  NOR2_X1 U856 ( .A1(G2090), .A2(G303), .ZN(n767) );
  NAND2_X1 U857 ( .A1(G8), .A2(n767), .ZN(n768) );
  NAND2_X1 U858 ( .A1(n769), .A2(n768), .ZN(n770) );
  XNOR2_X1 U859 ( .A(n770), .B(KEYINPUT106), .ZN(n772) );
  AND2_X1 U860 ( .A1(n772), .A2(n771), .ZN(n773) );
  NOR2_X1 U861 ( .A1(n774), .A2(n773), .ZN(n775) );
  INV_X1 U862 ( .A(n775), .ZN(n812) );
  XNOR2_X1 U863 ( .A(KEYINPUT92), .B(G1991), .ZN(n956) );
  NAND2_X1 U864 ( .A1(G95), .A2(n878), .ZN(n777) );
  NAND2_X1 U865 ( .A1(G131), .A2(n879), .ZN(n776) );
  NAND2_X1 U866 ( .A1(n777), .A2(n776), .ZN(n783) );
  NAND2_X1 U867 ( .A1(G119), .A2(n884), .ZN(n778) );
  XNOR2_X1 U868 ( .A(n778), .B(KEYINPUT90), .ZN(n781) );
  NAND2_X1 U869 ( .A1(G107), .A2(n882), .ZN(n779) );
  XOR2_X1 U870 ( .A(KEYINPUT91), .B(n779), .Z(n780) );
  NAND2_X1 U871 ( .A1(n781), .A2(n780), .ZN(n782) );
  OR2_X1 U872 ( .A1(n783), .A2(n782), .ZN(n873) );
  AND2_X1 U873 ( .A1(n956), .A2(n873), .ZN(n794) );
  NAND2_X1 U874 ( .A1(G105), .A2(n878), .ZN(n784) );
  XNOR2_X1 U875 ( .A(n784), .B(KEYINPUT38), .ZN(n791) );
  NAND2_X1 U876 ( .A1(G141), .A2(n879), .ZN(n786) );
  NAND2_X1 U877 ( .A1(G117), .A2(n882), .ZN(n785) );
  NAND2_X1 U878 ( .A1(n786), .A2(n785), .ZN(n789) );
  NAND2_X1 U879 ( .A1(G129), .A2(n884), .ZN(n787) );
  XNOR2_X1 U880 ( .A(KEYINPUT93), .B(n787), .ZN(n788) );
  NOR2_X1 U881 ( .A1(n789), .A2(n788), .ZN(n790) );
  NAND2_X1 U882 ( .A1(n791), .A2(n790), .ZN(n867) );
  NAND2_X1 U883 ( .A1(G1996), .A2(n867), .ZN(n792) );
  XOR2_X1 U884 ( .A(KEYINPUT94), .B(n792), .Z(n793) );
  NOR2_X1 U885 ( .A1(n794), .A2(n793), .ZN(n934) );
  NOR2_X1 U886 ( .A1(n796), .A2(n795), .ZN(n824) );
  INV_X1 U887 ( .A(n824), .ZN(n797) );
  NOR2_X1 U888 ( .A1(n934), .A2(n797), .ZN(n815) );
  INV_X1 U889 ( .A(n815), .ZN(n809) );
  NAND2_X1 U890 ( .A1(G104), .A2(n878), .ZN(n799) );
  NAND2_X1 U891 ( .A1(G140), .A2(n879), .ZN(n798) );
  NAND2_X1 U892 ( .A1(n799), .A2(n798), .ZN(n800) );
  XNOR2_X1 U893 ( .A(KEYINPUT34), .B(n800), .ZN(n806) );
  NAND2_X1 U894 ( .A1(n884), .A2(G128), .ZN(n801) );
  XNOR2_X1 U895 ( .A(n801), .B(KEYINPUT88), .ZN(n803) );
  NAND2_X1 U896 ( .A1(G116), .A2(n882), .ZN(n802) );
  NAND2_X1 U897 ( .A1(n803), .A2(n802), .ZN(n804) );
  XOR2_X1 U898 ( .A(n804), .B(KEYINPUT35), .Z(n805) );
  NOR2_X1 U899 ( .A1(n806), .A2(n805), .ZN(n807) );
  XOR2_X1 U900 ( .A(KEYINPUT36), .B(n807), .Z(n808) );
  XNOR2_X1 U901 ( .A(KEYINPUT89), .B(n808), .ZN(n890) );
  XNOR2_X1 U902 ( .A(G2067), .B(KEYINPUT37), .ZN(n821) );
  NOR2_X1 U903 ( .A1(n890), .A2(n821), .ZN(n925) );
  NAND2_X1 U904 ( .A1(n824), .A2(n925), .ZN(n819) );
  NAND2_X1 U905 ( .A1(n809), .A2(n819), .ZN(n810) );
  XNOR2_X1 U906 ( .A(G1986), .B(G290), .ZN(n1009) );
  NAND2_X1 U907 ( .A1(n812), .A2(n811), .ZN(n827) );
  NOR2_X1 U908 ( .A1(G1996), .A2(n867), .ZN(n929) );
  NOR2_X1 U909 ( .A1(G1986), .A2(G290), .ZN(n813) );
  NOR2_X1 U910 ( .A1(n956), .A2(n873), .ZN(n935) );
  NOR2_X1 U911 ( .A1(n813), .A2(n935), .ZN(n814) );
  NOR2_X1 U912 ( .A1(n815), .A2(n814), .ZN(n816) );
  XOR2_X1 U913 ( .A(KEYINPUT107), .B(n816), .Z(n817) );
  NOR2_X1 U914 ( .A1(n929), .A2(n817), .ZN(n818) );
  XNOR2_X1 U915 ( .A(n818), .B(KEYINPUT39), .ZN(n820) );
  NAND2_X1 U916 ( .A1(n820), .A2(n819), .ZN(n822) );
  NAND2_X1 U917 ( .A1(n890), .A2(n821), .ZN(n922) );
  NAND2_X1 U918 ( .A1(n822), .A2(n922), .ZN(n823) );
  NAND2_X1 U919 ( .A1(n824), .A2(n823), .ZN(n825) );
  XNOR2_X1 U920 ( .A(KEYINPUT108), .B(n825), .ZN(n826) );
  NAND2_X1 U921 ( .A1(n827), .A2(n826), .ZN(n828) );
  XNOR2_X1 U922 ( .A(n828), .B(KEYINPUT40), .ZN(G329) );
  NAND2_X1 U923 ( .A1(n829), .A2(G2106), .ZN(n830) );
  XNOR2_X1 U924 ( .A(n830), .B(KEYINPUT110), .ZN(G217) );
  AND2_X1 U925 ( .A1(G15), .A2(G2), .ZN(n831) );
  NAND2_X1 U926 ( .A1(G661), .A2(n831), .ZN(G259) );
  NAND2_X1 U927 ( .A1(G3), .A2(G1), .ZN(n832) );
  NAND2_X1 U928 ( .A1(n833), .A2(n832), .ZN(G188) );
  XOR2_X1 U929 ( .A(G2096), .B(KEYINPUT112), .Z(n835) );
  XNOR2_X1 U930 ( .A(G2072), .B(KEYINPUT43), .ZN(n834) );
  XNOR2_X1 U931 ( .A(n835), .B(n834), .ZN(n836) );
  XOR2_X1 U932 ( .A(n836), .B(KEYINPUT42), .Z(n838) );
  XNOR2_X1 U933 ( .A(G2067), .B(G2090), .ZN(n837) );
  XNOR2_X1 U934 ( .A(n838), .B(n837), .ZN(n842) );
  XOR2_X1 U935 ( .A(G2678), .B(G2100), .Z(n840) );
  XNOR2_X1 U936 ( .A(G2084), .B(G2078), .ZN(n839) );
  XNOR2_X1 U937 ( .A(n840), .B(n839), .ZN(n841) );
  XNOR2_X1 U938 ( .A(n842), .B(n841), .ZN(G227) );
  XOR2_X1 U939 ( .A(G1976), .B(G1971), .Z(n844) );
  XNOR2_X1 U940 ( .A(G1961), .B(G1956), .ZN(n843) );
  XNOR2_X1 U941 ( .A(n844), .B(n843), .ZN(n845) );
  XOR2_X1 U942 ( .A(n845), .B(KEYINPUT41), .Z(n847) );
  XNOR2_X1 U943 ( .A(G1966), .B(G1981), .ZN(n846) );
  XNOR2_X1 U944 ( .A(n847), .B(n846), .ZN(n851) );
  XOR2_X1 U945 ( .A(G2474), .B(G1986), .Z(n849) );
  XNOR2_X1 U946 ( .A(G1996), .B(G1991), .ZN(n848) );
  XNOR2_X1 U947 ( .A(n849), .B(n848), .ZN(n850) );
  XNOR2_X1 U948 ( .A(n851), .B(n850), .ZN(G229) );
  NAND2_X1 U949 ( .A1(n884), .A2(G124), .ZN(n852) );
  XNOR2_X1 U950 ( .A(n852), .B(KEYINPUT44), .ZN(n854) );
  NAND2_X1 U951 ( .A1(G136), .A2(n879), .ZN(n853) );
  NAND2_X1 U952 ( .A1(n854), .A2(n853), .ZN(n859) );
  NAND2_X1 U953 ( .A1(G100), .A2(n878), .ZN(n856) );
  NAND2_X1 U954 ( .A1(G112), .A2(n882), .ZN(n855) );
  NAND2_X1 U955 ( .A1(n856), .A2(n855), .ZN(n857) );
  XOR2_X1 U956 ( .A(KEYINPUT113), .B(n857), .Z(n858) );
  NOR2_X1 U957 ( .A1(n859), .A2(n858), .ZN(G162) );
  NAND2_X1 U958 ( .A1(G118), .A2(n882), .ZN(n861) );
  NAND2_X1 U959 ( .A1(G130), .A2(n884), .ZN(n860) );
  NAND2_X1 U960 ( .A1(n861), .A2(n860), .ZN(n866) );
  NAND2_X1 U961 ( .A1(G106), .A2(n878), .ZN(n863) );
  NAND2_X1 U962 ( .A1(G142), .A2(n879), .ZN(n862) );
  NAND2_X1 U963 ( .A1(n863), .A2(n862), .ZN(n864) );
  XOR2_X1 U964 ( .A(KEYINPUT45), .B(n864), .Z(n865) );
  NOR2_X1 U965 ( .A1(n866), .A2(n865), .ZN(n877) );
  XNOR2_X1 U966 ( .A(G162), .B(n867), .ZN(n868) );
  XNOR2_X1 U967 ( .A(n868), .B(n926), .ZN(n872) );
  XOR2_X1 U968 ( .A(KEYINPUT114), .B(KEYINPUT46), .Z(n870) );
  XNOR2_X1 U969 ( .A(G160), .B(KEYINPUT48), .ZN(n869) );
  XNOR2_X1 U970 ( .A(n870), .B(n869), .ZN(n871) );
  XOR2_X1 U971 ( .A(n872), .B(n871), .Z(n875) );
  XOR2_X1 U972 ( .A(G164), .B(n873), .Z(n874) );
  XNOR2_X1 U973 ( .A(n875), .B(n874), .ZN(n876) );
  XNOR2_X1 U974 ( .A(n877), .B(n876), .ZN(n892) );
  NAND2_X1 U975 ( .A1(G103), .A2(n878), .ZN(n881) );
  NAND2_X1 U976 ( .A1(G139), .A2(n879), .ZN(n880) );
  NAND2_X1 U977 ( .A1(n881), .A2(n880), .ZN(n889) );
  NAND2_X1 U978 ( .A1(n882), .A2(G115), .ZN(n883) );
  XOR2_X1 U979 ( .A(KEYINPUT115), .B(n883), .Z(n886) );
  NAND2_X1 U980 ( .A1(n884), .A2(G127), .ZN(n885) );
  NAND2_X1 U981 ( .A1(n886), .A2(n885), .ZN(n887) );
  XOR2_X1 U982 ( .A(KEYINPUT47), .B(n887), .Z(n888) );
  NOR2_X1 U983 ( .A1(n889), .A2(n888), .ZN(n918) );
  XNOR2_X1 U984 ( .A(n890), .B(n918), .ZN(n891) );
  XNOR2_X1 U985 ( .A(n892), .B(n891), .ZN(n893) );
  NOR2_X1 U986 ( .A1(G37), .A2(n893), .ZN(G395) );
  XNOR2_X1 U987 ( .A(n1000), .B(G286), .ZN(n895) );
  XNOR2_X1 U988 ( .A(n895), .B(n894), .ZN(n896) );
  XNOR2_X1 U989 ( .A(n896), .B(G171), .ZN(n897) );
  NOR2_X1 U990 ( .A1(G37), .A2(n897), .ZN(G397) );
  NOR2_X1 U991 ( .A1(G227), .A2(G229), .ZN(n899) );
  XNOR2_X1 U992 ( .A(KEYINPUT116), .B(KEYINPUT49), .ZN(n898) );
  XNOR2_X1 U993 ( .A(n899), .B(n898), .ZN(n911) );
  XOR2_X1 U994 ( .A(G2430), .B(G2451), .Z(n901) );
  XNOR2_X1 U995 ( .A(G2446), .B(G2427), .ZN(n900) );
  XNOR2_X1 U996 ( .A(n901), .B(n900), .ZN(n908) );
  XOR2_X1 U997 ( .A(G2438), .B(G2435), .Z(n903) );
  XNOR2_X1 U998 ( .A(G2443), .B(KEYINPUT109), .ZN(n902) );
  XNOR2_X1 U999 ( .A(n903), .B(n902), .ZN(n904) );
  XOR2_X1 U1000 ( .A(n904), .B(G2454), .Z(n906) );
  XNOR2_X1 U1001 ( .A(G1341), .B(G1348), .ZN(n905) );
  XNOR2_X1 U1002 ( .A(n906), .B(n905), .ZN(n907) );
  XNOR2_X1 U1003 ( .A(n908), .B(n907), .ZN(n909) );
  NAND2_X1 U1004 ( .A1(n909), .A2(G14), .ZN(n917) );
  NAND2_X1 U1005 ( .A1(n917), .A2(G319), .ZN(n910) );
  NOR2_X1 U1006 ( .A1(n911), .A2(n910), .ZN(n913) );
  NOR2_X1 U1007 ( .A1(G395), .A2(G397), .ZN(n912) );
  NAND2_X1 U1008 ( .A1(n913), .A2(n912), .ZN(G225) );
  XNOR2_X1 U1009 ( .A(KEYINPUT117), .B(G225), .ZN(G308) );
  INV_X1 U1011 ( .A(G132), .ZN(G219) );
  INV_X1 U1012 ( .A(G82), .ZN(G220) );
  NOR2_X1 U1013 ( .A1(n915), .A2(n914), .ZN(n916) );
  XNOR2_X1 U1014 ( .A(n916), .B(KEYINPUT111), .ZN(G261) );
  INV_X1 U1015 ( .A(G261), .ZN(G325) );
  INV_X1 U1016 ( .A(G96), .ZN(G221) );
  INV_X1 U1017 ( .A(G57), .ZN(G237) );
  INV_X1 U1018 ( .A(n917), .ZN(G401) );
  XOR2_X1 U1019 ( .A(G2072), .B(n918), .Z(n920) );
  XOR2_X1 U1020 ( .A(G164), .B(G2078), .Z(n919) );
  NOR2_X1 U1021 ( .A1(n920), .A2(n919), .ZN(n921) );
  XNOR2_X1 U1022 ( .A(n921), .B(KEYINPUT50), .ZN(n923) );
  NAND2_X1 U1023 ( .A1(n923), .A2(n922), .ZN(n924) );
  NOR2_X1 U1024 ( .A1(n925), .A2(n924), .ZN(n938) );
  XNOR2_X1 U1025 ( .A(G160), .B(G2084), .ZN(n927) );
  NAND2_X1 U1026 ( .A1(n927), .A2(n926), .ZN(n932) );
  XOR2_X1 U1027 ( .A(G2090), .B(G162), .Z(n928) );
  NOR2_X1 U1028 ( .A1(n929), .A2(n928), .ZN(n930) );
  XNOR2_X1 U1029 ( .A(n930), .B(KEYINPUT51), .ZN(n931) );
  NOR2_X1 U1030 ( .A1(n932), .A2(n931), .ZN(n933) );
  NAND2_X1 U1031 ( .A1(n934), .A2(n933), .ZN(n936) );
  NOR2_X1 U1032 ( .A1(n936), .A2(n935), .ZN(n937) );
  NAND2_X1 U1033 ( .A1(n938), .A2(n937), .ZN(n939) );
  XNOR2_X1 U1034 ( .A(KEYINPUT52), .B(n939), .ZN(n940) );
  XNOR2_X1 U1035 ( .A(n940), .B(KEYINPUT118), .ZN(n941) );
  NOR2_X1 U1036 ( .A1(KEYINPUT55), .A2(n941), .ZN(n942) );
  XNOR2_X1 U1037 ( .A(KEYINPUT119), .B(n942), .ZN(n943) );
  NAND2_X1 U1038 ( .A1(n943), .A2(G29), .ZN(n944) );
  XNOR2_X1 U1039 ( .A(n944), .B(KEYINPUT120), .ZN(n994) );
  XNOR2_X1 U1040 ( .A(G2084), .B(G34), .ZN(n945) );
  XNOR2_X1 U1041 ( .A(n945), .B(KEYINPUT54), .ZN(n964) );
  XNOR2_X1 U1042 ( .A(G2090), .B(G35), .ZN(n961) );
  XNOR2_X1 U1043 ( .A(KEYINPUT121), .B(G2067), .ZN(n946) );
  XNOR2_X1 U1044 ( .A(n946), .B(G26), .ZN(n955) );
  XNOR2_X1 U1045 ( .A(G1996), .B(G32), .ZN(n948) );
  XNOR2_X1 U1046 ( .A(G33), .B(G2072), .ZN(n947) );
  NOR2_X1 U1047 ( .A1(n948), .A2(n947), .ZN(n949) );
  NAND2_X1 U1048 ( .A1(G28), .A2(n949), .ZN(n953) );
  XOR2_X1 U1049 ( .A(G27), .B(n950), .Z(n951) );
  XNOR2_X1 U1050 ( .A(KEYINPUT122), .B(n951), .ZN(n952) );
  NOR2_X1 U1051 ( .A1(n953), .A2(n952), .ZN(n954) );
  NAND2_X1 U1052 ( .A1(n955), .A2(n954), .ZN(n958) );
  XNOR2_X1 U1053 ( .A(G25), .B(n956), .ZN(n957) );
  NOR2_X1 U1054 ( .A1(n958), .A2(n957), .ZN(n959) );
  XNOR2_X1 U1055 ( .A(KEYINPUT53), .B(n959), .ZN(n960) );
  NOR2_X1 U1056 ( .A1(n961), .A2(n960), .ZN(n962) );
  XNOR2_X1 U1057 ( .A(n962), .B(KEYINPUT123), .ZN(n963) );
  NOR2_X1 U1058 ( .A1(n964), .A2(n963), .ZN(n965) );
  XOR2_X1 U1059 ( .A(KEYINPUT55), .B(n965), .Z(n966) );
  NOR2_X1 U1060 ( .A1(G29), .A2(n966), .ZN(n992) );
  XNOR2_X1 U1061 ( .A(G5), .B(n967), .ZN(n979) );
  XOR2_X1 U1062 ( .A(G20), .B(G1956), .Z(n971) );
  XNOR2_X1 U1063 ( .A(G1341), .B(G19), .ZN(n969) );
  XNOR2_X1 U1064 ( .A(G6), .B(G1981), .ZN(n968) );
  NOR2_X1 U1065 ( .A1(n969), .A2(n968), .ZN(n970) );
  NAND2_X1 U1066 ( .A1(n971), .A2(n970), .ZN(n974) );
  XOR2_X1 U1067 ( .A(KEYINPUT59), .B(G1348), .Z(n972) );
  XNOR2_X1 U1068 ( .A(G4), .B(n972), .ZN(n973) );
  NOR2_X1 U1069 ( .A1(n974), .A2(n973), .ZN(n975) );
  XOR2_X1 U1070 ( .A(KEYINPUT60), .B(n975), .Z(n977) );
  XNOR2_X1 U1071 ( .A(G1966), .B(G21), .ZN(n976) );
  NOR2_X1 U1072 ( .A1(n977), .A2(n976), .ZN(n978) );
  NAND2_X1 U1073 ( .A1(n979), .A2(n978), .ZN(n986) );
  XNOR2_X1 U1074 ( .A(G1971), .B(G22), .ZN(n981) );
  XNOR2_X1 U1075 ( .A(G24), .B(G1986), .ZN(n980) );
  NOR2_X1 U1076 ( .A1(n981), .A2(n980), .ZN(n983) );
  XOR2_X1 U1077 ( .A(G1976), .B(G23), .Z(n982) );
  NAND2_X1 U1078 ( .A1(n983), .A2(n982), .ZN(n984) );
  XNOR2_X1 U1079 ( .A(KEYINPUT58), .B(n984), .ZN(n985) );
  NOR2_X1 U1080 ( .A1(n986), .A2(n985), .ZN(n987) );
  XNOR2_X1 U1081 ( .A(KEYINPUT61), .B(n987), .ZN(n989) );
  INV_X1 U1082 ( .A(G16), .ZN(n988) );
  NAND2_X1 U1083 ( .A1(n989), .A2(n988), .ZN(n990) );
  NAND2_X1 U1084 ( .A1(n990), .A2(G11), .ZN(n991) );
  NOR2_X1 U1085 ( .A1(n992), .A2(n991), .ZN(n993) );
  NAND2_X1 U1086 ( .A1(n994), .A2(n993), .ZN(n1024) );
  XOR2_X1 U1087 ( .A(KEYINPUT56), .B(G16), .Z(n1022) );
  XOR2_X1 U1088 ( .A(G168), .B(G1966), .Z(n995) );
  NOR2_X1 U1089 ( .A1(n996), .A2(n995), .ZN(n997) );
  XOR2_X1 U1090 ( .A(KEYINPUT57), .B(n997), .Z(n998) );
  XNOR2_X1 U1091 ( .A(KEYINPUT124), .B(n998), .ZN(n1004) );
  XNOR2_X1 U1092 ( .A(n999), .B(G1341), .ZN(n1002) );
  XNOR2_X1 U1093 ( .A(n1000), .B(G1348), .ZN(n1001) );
  NOR2_X1 U1094 ( .A1(n1002), .A2(n1001), .ZN(n1003) );
  NAND2_X1 U1095 ( .A1(n1004), .A2(n1003), .ZN(n1020) );
  XNOR2_X1 U1096 ( .A(n1005), .B(G1956), .ZN(n1007) );
  XNOR2_X1 U1097 ( .A(G171), .B(G1961), .ZN(n1006) );
  NAND2_X1 U1098 ( .A1(n1007), .A2(n1006), .ZN(n1008) );
  NOR2_X1 U1099 ( .A1(n1009), .A2(n1008), .ZN(n1018) );
  XNOR2_X1 U1100 ( .A(G166), .B(G1971), .ZN(n1010) );
  XNOR2_X1 U1101 ( .A(n1010), .B(KEYINPUT126), .ZN(n1015) );
  NAND2_X1 U1102 ( .A1(n1012), .A2(n1011), .ZN(n1013) );
  XNOR2_X1 U1103 ( .A(KEYINPUT125), .B(n1013), .ZN(n1014) );
  NAND2_X1 U1104 ( .A1(n1015), .A2(n1014), .ZN(n1016) );
  XNOR2_X1 U1105 ( .A(n1016), .B(KEYINPUT127), .ZN(n1017) );
  NAND2_X1 U1106 ( .A1(n1018), .A2(n1017), .ZN(n1019) );
  NOR2_X1 U1107 ( .A1(n1020), .A2(n1019), .ZN(n1021) );
  NOR2_X1 U1108 ( .A1(n1022), .A2(n1021), .ZN(n1023) );
  NOR2_X1 U1109 ( .A1(n1024), .A2(n1023), .ZN(n1025) );
  XNOR2_X1 U1110 ( .A(n1025), .B(KEYINPUT62), .ZN(G311) );
  INV_X1 U1111 ( .A(G311), .ZN(G150) );
endmodule

