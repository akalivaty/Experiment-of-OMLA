//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 0 1 1 0 0 0 1 0 0 0 0 0 0 0 1 1 0 1 0 0 1 0 1 1 0 0 1 1 0 0 1 1 1 1 0 0 1 0 1 1 0 1 0 0 0 1 1 1 1 1 1 1 0 0 1 0 1 0 1 0 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:38:03 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n204, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n223, new_n224,
    new_n225, new_n226, new_n227, new_n228, new_n229, new_n230, new_n232,
    new_n233, new_n234, new_n235, new_n236, new_n237, new_n239, new_n240,
    new_n241, new_n242, new_n243, new_n244, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1248,
    new_n1249, new_n1250, new_n1251, new_n1252, new_n1253, new_n1254,
    new_n1255, new_n1256, new_n1257, new_n1259, new_n1260, new_n1261,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1329,
    new_n1330, new_n1331, new_n1332, new_n1333, new_n1334, new_n1335,
    new_n1336, new_n1337, new_n1338;
  OR2_X1    g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  NOR3_X1   g0001(.A1(new_n201), .A2(G50), .A3(G77), .ZN(G353));
  OAI21_X1  g0002(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0003(.A1(G1), .A2(G20), .ZN(new_n204));
  NOR2_X1   g0004(.A1(new_n204), .A2(G13), .ZN(new_n205));
  OAI211_X1 g0005(.A(new_n205), .B(G250), .C1(G257), .C2(G264), .ZN(new_n206));
  XNOR2_X1  g0006(.A(new_n206), .B(KEYINPUT0), .ZN(new_n207));
  AND2_X1   g0007(.A1(G1), .A2(G13), .ZN(new_n208));
  NAND2_X1  g0008(.A1(new_n208), .A2(G20), .ZN(new_n209));
  NAND2_X1  g0009(.A1(new_n201), .A2(G50), .ZN(new_n210));
  AOI22_X1  g0010(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n211));
  INV_X1    g0011(.A(G68), .ZN(new_n212));
  INV_X1    g0012(.A(G238), .ZN(new_n213));
  INV_X1    g0013(.A(G87), .ZN(new_n214));
  INV_X1    g0014(.A(G250), .ZN(new_n215));
  OAI221_X1 g0015(.A(new_n211), .B1(new_n212), .B2(new_n213), .C1(new_n214), .C2(new_n215), .ZN(new_n216));
  AOI22_X1  g0016(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n217));
  AOI22_X1  g0017(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n218));
  NAND2_X1  g0018(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  OAI21_X1  g0019(.A(new_n204), .B1(new_n216), .B2(new_n219), .ZN(new_n220));
  OAI221_X1 g0020(.A(new_n207), .B1(new_n209), .B2(new_n210), .C1(KEYINPUT1), .C2(new_n220), .ZN(new_n221));
  AOI21_X1  g0021(.A(new_n221), .B1(KEYINPUT1), .B2(new_n220), .ZN(G361));
  XNOR2_X1  g0022(.A(G238), .B(G244), .ZN(new_n223));
  INV_X1    g0023(.A(G232), .ZN(new_n224));
  XNOR2_X1  g0024(.A(new_n223), .B(new_n224), .ZN(new_n225));
  XOR2_X1   g0025(.A(KEYINPUT2), .B(G226), .Z(new_n226));
  XNOR2_X1  g0026(.A(new_n225), .B(new_n226), .ZN(new_n227));
  XOR2_X1   g0027(.A(G264), .B(G270), .Z(new_n228));
  XNOR2_X1  g0028(.A(G250), .B(G257), .ZN(new_n229));
  XNOR2_X1  g0029(.A(new_n228), .B(new_n229), .ZN(new_n230));
  XNOR2_X1  g0030(.A(new_n227), .B(new_n230), .ZN(G358));
  XNOR2_X1  g0031(.A(G50), .B(G68), .ZN(new_n232));
  XNOR2_X1  g0032(.A(G58), .B(G77), .ZN(new_n233));
  XOR2_X1   g0033(.A(new_n232), .B(new_n233), .Z(new_n234));
  XOR2_X1   g0034(.A(G87), .B(G97), .Z(new_n235));
  XNOR2_X1  g0035(.A(G107), .B(G116), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n234), .B(new_n237), .ZN(G351));
  INV_X1    g0038(.A(KEYINPUT13), .ZN(new_n239));
  INV_X1    g0039(.A(KEYINPUT3), .ZN(new_n240));
  INV_X1    g0040(.A(G33), .ZN(new_n241));
  NAND2_X1  g0041(.A1(new_n240), .A2(new_n241), .ZN(new_n242));
  NAND2_X1  g0042(.A1(KEYINPUT3), .A2(G33), .ZN(new_n243));
  NAND2_X1  g0043(.A1(new_n242), .A2(new_n243), .ZN(new_n244));
  NAND3_X1  g0044(.A1(new_n244), .A2(G232), .A3(G1698), .ZN(new_n245));
  INV_X1    g0045(.A(G1698), .ZN(new_n246));
  NAND3_X1  g0046(.A1(new_n244), .A2(G226), .A3(new_n246), .ZN(new_n247));
  NAND2_X1  g0047(.A1(G33), .A2(G97), .ZN(new_n248));
  NAND3_X1  g0048(.A1(new_n245), .A2(new_n247), .A3(new_n248), .ZN(new_n249));
  NAND2_X1  g0049(.A1(G33), .A2(G41), .ZN(new_n250));
  NAND3_X1  g0050(.A1(new_n250), .A2(G1), .A3(G13), .ZN(new_n251));
  INV_X1    g0051(.A(new_n251), .ZN(new_n252));
  NAND2_X1  g0052(.A1(new_n249), .A2(new_n252), .ZN(new_n253));
  INV_X1    g0053(.A(G274), .ZN(new_n254));
  AOI21_X1  g0054(.A(new_n254), .B1(new_n208), .B2(new_n250), .ZN(new_n255));
  INV_X1    g0055(.A(G1), .ZN(new_n256));
  OAI21_X1  g0056(.A(new_n256), .B1(G41), .B2(G45), .ZN(new_n257));
  INV_X1    g0057(.A(new_n257), .ZN(new_n258));
  AND2_X1   g0058(.A1(new_n255), .A2(new_n258), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n251), .A2(new_n257), .ZN(new_n260));
  INV_X1    g0060(.A(new_n260), .ZN(new_n261));
  AOI21_X1  g0061(.A(new_n259), .B1(G238), .B2(new_n261), .ZN(new_n262));
  AOI21_X1  g0062(.A(new_n239), .B1(new_n253), .B2(new_n262), .ZN(new_n263));
  INV_X1    g0063(.A(new_n263), .ZN(new_n264));
  NAND3_X1  g0064(.A1(new_n253), .A2(new_n262), .A3(new_n239), .ZN(new_n265));
  NAND3_X1  g0065(.A1(new_n264), .A2(G190), .A3(new_n265), .ZN(new_n266));
  INV_X1    g0066(.A(new_n265), .ZN(new_n267));
  OAI21_X1  g0067(.A(G200), .B1(new_n267), .B2(new_n263), .ZN(new_n268));
  INV_X1    g0068(.A(G20), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n269), .A2(new_n241), .ZN(new_n270));
  INV_X1    g0070(.A(new_n270), .ZN(new_n271));
  AOI22_X1  g0071(.A1(new_n271), .A2(G50), .B1(G20), .B2(new_n212), .ZN(new_n272));
  INV_X1    g0072(.A(G77), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n269), .A2(G33), .ZN(new_n274));
  OAI21_X1  g0074(.A(new_n272), .B1(new_n273), .B2(new_n274), .ZN(new_n275));
  OAI21_X1  g0075(.A(KEYINPUT64), .B1(new_n204), .B2(new_n241), .ZN(new_n276));
  NAND2_X1  g0076(.A1(G1), .A2(G13), .ZN(new_n277));
  INV_X1    g0077(.A(KEYINPUT64), .ZN(new_n278));
  NAND4_X1  g0078(.A1(new_n278), .A2(G1), .A3(G20), .A4(G33), .ZN(new_n279));
  NAND3_X1  g0079(.A1(new_n276), .A2(new_n277), .A3(new_n279), .ZN(new_n280));
  NAND3_X1  g0080(.A1(new_n275), .A2(KEYINPUT11), .A3(new_n280), .ZN(new_n281));
  INV_X1    g0081(.A(G13), .ZN(new_n282));
  NOR3_X1   g0082(.A1(new_n282), .A2(new_n269), .A3(G1), .ZN(new_n283));
  NOR2_X1   g0083(.A1(new_n280), .A2(new_n283), .ZN(new_n284));
  NOR2_X1   g0084(.A1(new_n269), .A2(G1), .ZN(new_n285));
  INV_X1    g0085(.A(new_n285), .ZN(new_n286));
  NAND3_X1  g0086(.A1(new_n284), .A2(G68), .A3(new_n286), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n281), .A2(new_n287), .ZN(new_n288));
  AOI21_X1  g0088(.A(KEYINPUT11), .B1(new_n275), .B2(new_n280), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n283), .A2(new_n212), .ZN(new_n290));
  NOR2_X1   g0090(.A1(KEYINPUT70), .A2(KEYINPUT12), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  XNOR2_X1  g0092(.A(KEYINPUT70), .B(KEYINPUT12), .ZN(new_n293));
  OAI21_X1  g0093(.A(new_n292), .B1(new_n290), .B2(new_n293), .ZN(new_n294));
  NOR3_X1   g0094(.A1(new_n288), .A2(new_n289), .A3(new_n294), .ZN(new_n295));
  NAND3_X1  g0095(.A1(new_n266), .A2(new_n268), .A3(new_n295), .ZN(new_n296));
  INV_X1    g0096(.A(KEYINPUT71), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n296), .A2(new_n297), .ZN(new_n298));
  NAND4_X1  g0098(.A1(new_n266), .A2(new_n268), .A3(KEYINPUT71), .A4(new_n295), .ZN(new_n299));
  NAND2_X1  g0099(.A1(KEYINPUT72), .A2(G169), .ZN(new_n300));
  INV_X1    g0100(.A(new_n300), .ZN(new_n301));
  OAI21_X1  g0101(.A(new_n301), .B1(new_n267), .B2(new_n263), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n302), .A2(KEYINPUT14), .ZN(new_n303));
  INV_X1    g0103(.A(KEYINPUT14), .ZN(new_n304));
  OAI211_X1 g0104(.A(new_n304), .B(new_n301), .C1(new_n267), .C2(new_n263), .ZN(new_n305));
  NAND3_X1  g0105(.A1(new_n264), .A2(G179), .A3(new_n265), .ZN(new_n306));
  NAND3_X1  g0106(.A1(new_n303), .A2(new_n305), .A3(new_n306), .ZN(new_n307));
  INV_X1    g0107(.A(new_n295), .ZN(new_n308));
  AOI22_X1  g0108(.A1(new_n298), .A2(new_n299), .B1(new_n307), .B2(new_n308), .ZN(new_n309));
  INV_X1    g0109(.A(KEYINPUT75), .ZN(new_n310));
  INV_X1    g0110(.A(G159), .ZN(new_n311));
  NOR2_X1   g0111(.A1(new_n270), .A2(new_n311), .ZN(new_n312));
  NAND2_X1  g0112(.A1(G58), .A2(G68), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n313), .A2(KEYINPUT74), .ZN(new_n314));
  INV_X1    g0114(.A(KEYINPUT74), .ZN(new_n315));
  NAND3_X1  g0115(.A1(new_n315), .A2(G58), .A3(G68), .ZN(new_n316));
  NAND3_X1  g0116(.A1(new_n314), .A2(new_n316), .A3(new_n201), .ZN(new_n317));
  AOI21_X1  g0117(.A(new_n312), .B1(new_n317), .B2(G20), .ZN(new_n318));
  AND2_X1   g0118(.A1(KEYINPUT3), .A2(G33), .ZN(new_n319));
  NOR2_X1   g0119(.A1(KEYINPUT3), .A2(G33), .ZN(new_n320));
  NOR3_X1   g0120(.A1(new_n319), .A2(new_n320), .A3(G20), .ZN(new_n321));
  INV_X1    g0121(.A(KEYINPUT7), .ZN(new_n322));
  OAI21_X1  g0122(.A(G68), .B1(new_n321), .B2(new_n322), .ZN(new_n323));
  NAND3_X1  g0123(.A1(new_n242), .A2(new_n269), .A3(new_n243), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n322), .A2(KEYINPUT73), .ZN(new_n325));
  INV_X1    g0125(.A(KEYINPUT73), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n326), .A2(KEYINPUT7), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n325), .A2(new_n327), .ZN(new_n328));
  NOR2_X1   g0128(.A1(new_n324), .A2(new_n328), .ZN(new_n329));
  OAI211_X1 g0129(.A(KEYINPUT16), .B(new_n318), .C1(new_n323), .C2(new_n329), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n330), .A2(new_n280), .ZN(new_n331));
  NAND4_X1  g0131(.A1(new_n242), .A2(KEYINPUT7), .A3(new_n269), .A4(new_n243), .ZN(new_n332));
  OAI21_X1  g0132(.A(new_n332), .B1(new_n321), .B2(new_n328), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n333), .A2(G68), .ZN(new_n334));
  AOI21_X1  g0134(.A(KEYINPUT16), .B1(new_n334), .B2(new_n318), .ZN(new_n335));
  OAI21_X1  g0135(.A(new_n310), .B1(new_n331), .B2(new_n335), .ZN(new_n336));
  INV_X1    g0136(.A(KEYINPUT16), .ZN(new_n337));
  INV_X1    g0137(.A(new_n318), .ZN(new_n338));
  XNOR2_X1  g0138(.A(KEYINPUT73), .B(KEYINPUT7), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n324), .A2(new_n339), .ZN(new_n340));
  AOI21_X1  g0140(.A(new_n212), .B1(new_n340), .B2(new_n332), .ZN(new_n341));
  OAI21_X1  g0141(.A(new_n337), .B1(new_n338), .B2(new_n341), .ZN(new_n342));
  NAND4_X1  g0142(.A1(new_n342), .A2(KEYINPUT75), .A3(new_n280), .A4(new_n330), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n336), .A2(new_n343), .ZN(new_n344));
  XNOR2_X1  g0144(.A(KEYINPUT8), .B(G58), .ZN(new_n345));
  NOR2_X1   g0145(.A1(new_n345), .A2(new_n285), .ZN(new_n346));
  AOI22_X1  g0146(.A1(new_n284), .A2(new_n346), .B1(new_n283), .B2(new_n345), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n344), .A2(new_n347), .ZN(new_n348));
  INV_X1    g0148(.A(KEYINPUT76), .ZN(new_n349));
  OAI21_X1  g0149(.A(new_n349), .B1(new_n260), .B2(new_n224), .ZN(new_n350));
  NAND4_X1  g0150(.A1(new_n251), .A2(new_n257), .A3(KEYINPUT76), .A4(G232), .ZN(new_n351));
  AOI21_X1  g0151(.A(new_n259), .B1(new_n350), .B2(new_n351), .ZN(new_n352));
  OAI211_X1 g0152(.A(G223), .B(new_n246), .C1(new_n319), .C2(new_n320), .ZN(new_n353));
  OAI211_X1 g0153(.A(G226), .B(G1698), .C1(new_n319), .C2(new_n320), .ZN(new_n354));
  OAI211_X1 g0154(.A(new_n353), .B(new_n354), .C1(new_n241), .C2(new_n214), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n355), .A2(new_n252), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n352), .A2(new_n356), .ZN(new_n357));
  INV_X1    g0157(.A(G179), .ZN(new_n358));
  NOR2_X1   g0158(.A1(new_n357), .A2(new_n358), .ZN(new_n359));
  INV_X1    g0159(.A(G169), .ZN(new_n360));
  AOI21_X1  g0160(.A(new_n360), .B1(new_n352), .B2(new_n356), .ZN(new_n361));
  NOR2_X1   g0161(.A1(new_n359), .A2(new_n361), .ZN(new_n362));
  INV_X1    g0162(.A(new_n362), .ZN(new_n363));
  NAND3_X1  g0163(.A1(new_n348), .A2(KEYINPUT18), .A3(new_n363), .ZN(new_n364));
  INV_X1    g0164(.A(KEYINPUT18), .ZN(new_n365));
  INV_X1    g0165(.A(new_n347), .ZN(new_n366));
  AOI21_X1  g0166(.A(new_n366), .B1(new_n336), .B2(new_n343), .ZN(new_n367));
  OAI21_X1  g0167(.A(new_n365), .B1(new_n367), .B2(new_n362), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n364), .A2(new_n368), .ZN(new_n369));
  INV_X1    g0169(.A(G190), .ZN(new_n370));
  NAND3_X1  g0170(.A1(new_n352), .A2(new_n370), .A3(new_n356), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n371), .A2(KEYINPUT77), .ZN(new_n372));
  INV_X1    g0172(.A(G200), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n357), .A2(new_n373), .ZN(new_n374));
  INV_X1    g0174(.A(KEYINPUT77), .ZN(new_n375));
  NAND4_X1  g0175(.A1(new_n352), .A2(new_n356), .A3(new_n375), .A4(new_n370), .ZN(new_n376));
  NAND3_X1  g0176(.A1(new_n372), .A2(new_n374), .A3(new_n376), .ZN(new_n377));
  AND4_X1   g0177(.A1(KEYINPUT17), .A2(new_n344), .A3(new_n347), .A4(new_n377), .ZN(new_n378));
  AOI21_X1  g0178(.A(KEYINPUT17), .B1(new_n367), .B2(new_n377), .ZN(new_n379));
  NOR2_X1   g0179(.A1(new_n378), .A2(new_n379), .ZN(new_n380));
  NAND3_X1  g0180(.A1(new_n309), .A2(new_n369), .A3(new_n380), .ZN(new_n381));
  NAND3_X1  g0181(.A1(new_n284), .A2(G50), .A3(new_n286), .ZN(new_n382));
  INV_X1    g0182(.A(G150), .ZN(new_n383));
  OAI22_X1  g0183(.A1(new_n345), .A2(new_n274), .B1(new_n383), .B2(new_n270), .ZN(new_n384));
  NOR2_X1   g0184(.A1(new_n201), .A2(G50), .ZN(new_n385));
  NOR2_X1   g0185(.A1(new_n385), .A2(new_n269), .ZN(new_n386));
  OAI21_X1  g0186(.A(new_n280), .B1(new_n384), .B2(new_n386), .ZN(new_n387));
  INV_X1    g0187(.A(G50), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n283), .A2(new_n388), .ZN(new_n389));
  NAND3_X1  g0189(.A1(new_n382), .A2(new_n387), .A3(new_n389), .ZN(new_n390));
  XNOR2_X1  g0190(.A(new_n390), .B(KEYINPUT9), .ZN(new_n391));
  NAND3_X1  g0191(.A1(new_n244), .A2(G222), .A3(new_n246), .ZN(new_n392));
  NAND3_X1  g0192(.A1(new_n244), .A2(G223), .A3(G1698), .ZN(new_n393));
  OAI211_X1 g0193(.A(new_n392), .B(new_n393), .C1(new_n273), .C2(new_n244), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n394), .A2(new_n252), .ZN(new_n395));
  AOI21_X1  g0195(.A(new_n259), .B1(G226), .B2(new_n261), .ZN(new_n396));
  AOI21_X1  g0196(.A(new_n373), .B1(new_n395), .B2(new_n396), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n395), .A2(new_n396), .ZN(new_n398));
  INV_X1    g0198(.A(new_n398), .ZN(new_n399));
  AOI21_X1  g0199(.A(new_n397), .B1(new_n399), .B2(G190), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n391), .A2(new_n400), .ZN(new_n401));
  OAI21_X1  g0201(.A(KEYINPUT10), .B1(new_n397), .B2(KEYINPUT68), .ZN(new_n402));
  INV_X1    g0202(.A(new_n402), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n401), .A2(new_n403), .ZN(new_n404));
  NAND3_X1  g0204(.A1(new_n391), .A2(new_n400), .A3(new_n402), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n404), .A2(new_n405), .ZN(new_n406));
  OAI21_X1  g0206(.A(new_n390), .B1(new_n399), .B2(G169), .ZN(new_n407));
  NOR2_X1   g0207(.A1(new_n398), .A2(G179), .ZN(new_n408));
  NOR2_X1   g0208(.A1(new_n407), .A2(new_n408), .ZN(new_n409));
  INV_X1    g0209(.A(new_n409), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n406), .A2(new_n410), .ZN(new_n411));
  INV_X1    g0211(.A(new_n411), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n255), .A2(new_n258), .ZN(new_n413));
  INV_X1    g0213(.A(G244), .ZN(new_n414));
  OAI21_X1  g0214(.A(new_n413), .B1(new_n414), .B2(new_n260), .ZN(new_n415));
  NAND3_X1  g0215(.A1(new_n244), .A2(G232), .A3(new_n246), .ZN(new_n416));
  NAND3_X1  g0216(.A1(new_n244), .A2(G238), .A3(G1698), .ZN(new_n417));
  INV_X1    g0217(.A(G107), .ZN(new_n418));
  OAI211_X1 g0218(.A(new_n416), .B(new_n417), .C1(new_n418), .C2(new_n244), .ZN(new_n419));
  AOI21_X1  g0219(.A(new_n415), .B1(new_n419), .B2(new_n252), .ZN(new_n420));
  INV_X1    g0220(.A(new_n420), .ZN(new_n421));
  NOR2_X1   g0221(.A1(new_n421), .A2(new_n370), .ZN(new_n422));
  INV_X1    g0222(.A(KEYINPUT15), .ZN(new_n423));
  NOR2_X1   g0223(.A1(new_n423), .A2(G87), .ZN(new_n424));
  NOR2_X1   g0224(.A1(new_n214), .A2(KEYINPUT15), .ZN(new_n425));
  OAI21_X1  g0225(.A(KEYINPUT65), .B1(new_n424), .B2(new_n425), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n214), .A2(KEYINPUT15), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n423), .A2(G87), .ZN(new_n428));
  INV_X1    g0228(.A(KEYINPUT65), .ZN(new_n429));
  NAND3_X1  g0229(.A1(new_n427), .A2(new_n428), .A3(new_n429), .ZN(new_n430));
  NAND4_X1  g0230(.A1(new_n426), .A2(new_n269), .A3(G33), .A4(new_n430), .ZN(new_n431));
  XOR2_X1   g0231(.A(KEYINPUT8), .B(G58), .Z(new_n432));
  AOI22_X1  g0232(.A1(new_n432), .A2(new_n271), .B1(G20), .B2(G77), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n431), .A2(new_n433), .ZN(new_n434));
  AOI22_X1  g0234(.A1(new_n434), .A2(new_n280), .B1(new_n273), .B2(new_n283), .ZN(new_n435));
  NAND3_X1  g0235(.A1(new_n284), .A2(G77), .A3(new_n286), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n435), .A2(new_n436), .ZN(new_n437));
  INV_X1    g0237(.A(KEYINPUT66), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n437), .A2(new_n438), .ZN(new_n439));
  NAND3_X1  g0239(.A1(new_n435), .A2(KEYINPUT66), .A3(new_n436), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n421), .A2(G200), .ZN(new_n441));
  NAND3_X1  g0241(.A1(new_n439), .A2(new_n440), .A3(new_n441), .ZN(new_n442));
  AOI21_X1  g0242(.A(new_n422), .B1(new_n442), .B2(KEYINPUT67), .ZN(new_n443));
  INV_X1    g0243(.A(KEYINPUT67), .ZN(new_n444));
  NAND4_X1  g0244(.A1(new_n439), .A2(new_n441), .A3(new_n444), .A4(new_n440), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n443), .A2(new_n445), .ZN(new_n446));
  INV_X1    g0246(.A(KEYINPUT69), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n420), .A2(new_n358), .ZN(new_n448));
  OAI21_X1  g0248(.A(new_n448), .B1(G169), .B2(new_n420), .ZN(new_n449));
  AOI21_X1  g0249(.A(new_n449), .B1(new_n439), .B2(new_n440), .ZN(new_n450));
  INV_X1    g0250(.A(new_n450), .ZN(new_n451));
  NAND4_X1  g0251(.A1(new_n412), .A2(new_n446), .A3(new_n447), .A4(new_n451), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n446), .A2(new_n451), .ZN(new_n453));
  OAI21_X1  g0253(.A(KEYINPUT69), .B1(new_n453), .B2(new_n411), .ZN(new_n454));
  AOI21_X1  g0254(.A(new_n381), .B1(new_n452), .B2(new_n454), .ZN(new_n455));
  INV_X1    g0255(.A(G45), .ZN(new_n456));
  NOR2_X1   g0256(.A1(new_n456), .A2(G1), .ZN(new_n457));
  XNOR2_X1  g0257(.A(KEYINPUT5), .B(G41), .ZN(new_n458));
  AOI21_X1  g0258(.A(new_n252), .B1(new_n457), .B2(new_n458), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n459), .A2(G264), .ZN(new_n460));
  NAND3_X1  g0260(.A1(new_n255), .A2(new_n457), .A3(new_n458), .ZN(new_n461));
  AND2_X1   g0261(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n244), .A2(G257), .ZN(new_n463));
  INV_X1    g0263(.A(G294), .ZN(new_n464));
  OAI22_X1  g0264(.A1(new_n463), .A2(new_n246), .B1(new_n241), .B2(new_n464), .ZN(new_n465));
  NAND3_X1  g0265(.A1(new_n244), .A2(G250), .A3(new_n246), .ZN(new_n466));
  INV_X1    g0266(.A(KEYINPUT84), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  NAND4_X1  g0268(.A1(new_n244), .A2(KEYINPUT84), .A3(G250), .A4(new_n246), .ZN(new_n469));
  AOI21_X1  g0269(.A(new_n465), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  OAI211_X1 g0270(.A(new_n462), .B(new_n358), .C1(new_n470), .C2(new_n251), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n468), .A2(new_n469), .ZN(new_n472));
  AND2_X1   g0272(.A1(new_n244), .A2(G257), .ZN(new_n473));
  AOI22_X1  g0273(.A1(new_n473), .A2(G1698), .B1(G33), .B2(G294), .ZN(new_n474));
  AOI21_X1  g0274(.A(new_n251), .B1(new_n472), .B2(new_n474), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n460), .A2(new_n461), .ZN(new_n476));
  OAI21_X1  g0276(.A(new_n360), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  NOR2_X1   g0277(.A1(new_n241), .A2(G1), .ZN(new_n478));
  NOR3_X1   g0278(.A1(new_n280), .A2(new_n283), .A3(new_n478), .ZN(new_n479));
  AND2_X1   g0279(.A1(new_n479), .A2(G107), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n283), .A2(new_n418), .ZN(new_n481));
  XNOR2_X1  g0281(.A(new_n481), .B(KEYINPUT25), .ZN(new_n482));
  NOR2_X1   g0282(.A1(new_n480), .A2(new_n482), .ZN(new_n483));
  INV_X1    g0283(.A(new_n483), .ZN(new_n484));
  INV_X1    g0284(.A(new_n280), .ZN(new_n485));
  NAND2_X1  g0285(.A1(G33), .A2(G116), .ZN(new_n486));
  NOR2_X1   g0286(.A1(new_n486), .A2(G20), .ZN(new_n487));
  INV_X1    g0287(.A(KEYINPUT23), .ZN(new_n488));
  OAI21_X1  g0288(.A(new_n488), .B1(new_n269), .B2(G107), .ZN(new_n489));
  NAND3_X1  g0289(.A1(new_n418), .A2(KEYINPUT23), .A3(G20), .ZN(new_n490));
  AOI21_X1  g0290(.A(new_n487), .B1(new_n489), .B2(new_n490), .ZN(new_n491));
  OAI211_X1 g0291(.A(new_n269), .B(G87), .C1(new_n319), .C2(new_n320), .ZN(new_n492));
  AND2_X1   g0292(.A1(KEYINPUT83), .A2(KEYINPUT22), .ZN(new_n493));
  AND2_X1   g0293(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  NOR2_X1   g0294(.A1(new_n492), .A2(new_n493), .ZN(new_n495));
  OAI21_X1  g0295(.A(new_n491), .B1(new_n494), .B2(new_n495), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n496), .A2(KEYINPUT24), .ZN(new_n497));
  XNOR2_X1  g0297(.A(new_n492), .B(new_n493), .ZN(new_n498));
  INV_X1    g0298(.A(KEYINPUT24), .ZN(new_n499));
  NAND3_X1  g0299(.A1(new_n498), .A2(new_n499), .A3(new_n491), .ZN(new_n500));
  AOI21_X1  g0300(.A(new_n485), .B1(new_n497), .B2(new_n500), .ZN(new_n501));
  OAI211_X1 g0301(.A(new_n471), .B(new_n477), .C1(new_n484), .C2(new_n501), .ZN(new_n502));
  NAND3_X1  g0302(.A1(new_n244), .A2(G264), .A3(G1698), .ZN(new_n503));
  NAND3_X1  g0303(.A1(new_n244), .A2(G257), .A3(new_n246), .ZN(new_n504));
  NOR2_X1   g0304(.A1(new_n319), .A2(new_n320), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n505), .A2(G303), .ZN(new_n506));
  NAND3_X1  g0306(.A1(new_n503), .A2(new_n504), .A3(new_n506), .ZN(new_n507));
  AOI22_X1  g0307(.A1(new_n507), .A2(new_n252), .B1(G270), .B2(new_n459), .ZN(new_n508));
  AOI21_X1  g0308(.A(new_n360), .B1(new_n508), .B2(new_n461), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n479), .A2(G116), .ZN(new_n510));
  INV_X1    g0310(.A(new_n283), .ZN(new_n511));
  NOR2_X1   g0311(.A1(new_n511), .A2(G116), .ZN(new_n512));
  INV_X1    g0312(.A(new_n512), .ZN(new_n513));
  AOI21_X1  g0313(.A(G20), .B1(new_n241), .B2(G97), .ZN(new_n514));
  NAND2_X1  g0314(.A1(G33), .A2(G283), .ZN(new_n515));
  INV_X1    g0315(.A(KEYINPUT79), .ZN(new_n516));
  NOR2_X1   g0316(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  AOI21_X1  g0317(.A(KEYINPUT79), .B1(G33), .B2(G283), .ZN(new_n518));
  OAI21_X1  g0318(.A(new_n514), .B1(new_n517), .B2(new_n518), .ZN(new_n519));
  INV_X1    g0319(.A(G116), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n520), .A2(G20), .ZN(new_n521));
  AND2_X1   g0321(.A1(new_n519), .A2(new_n521), .ZN(new_n522));
  AOI21_X1  g0322(.A(KEYINPUT20), .B1(new_n522), .B2(new_n280), .ZN(new_n523));
  AND4_X1   g0323(.A1(KEYINPUT20), .A2(new_n280), .A3(new_n519), .A4(new_n521), .ZN(new_n524));
  OAI211_X1 g0324(.A(new_n510), .B(new_n513), .C1(new_n523), .C2(new_n524), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n509), .A2(new_n525), .ZN(new_n526));
  INV_X1    g0326(.A(KEYINPUT21), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  NAND4_X1  g0328(.A1(new_n525), .A2(G179), .A3(new_n461), .A4(new_n508), .ZN(new_n529));
  NAND3_X1  g0329(.A1(new_n509), .A2(new_n525), .A3(KEYINPUT21), .ZN(new_n530));
  NAND4_X1  g0330(.A1(new_n502), .A2(new_n528), .A3(new_n529), .A4(new_n530), .ZN(new_n531));
  INV_X1    g0331(.A(new_n531), .ZN(new_n532));
  OAI211_X1 g0332(.A(G244), .B(new_n246), .C1(new_n319), .C2(new_n320), .ZN(new_n533));
  INV_X1    g0333(.A(KEYINPUT4), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  NAND4_X1  g0335(.A1(new_n244), .A2(KEYINPUT4), .A3(G244), .A4(new_n246), .ZN(new_n536));
  XNOR2_X1  g0336(.A(new_n515), .B(new_n516), .ZN(new_n537));
  NAND3_X1  g0337(.A1(new_n244), .A2(G250), .A3(G1698), .ZN(new_n538));
  NAND4_X1  g0338(.A1(new_n535), .A2(new_n536), .A3(new_n537), .A4(new_n538), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n539), .A2(new_n252), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n458), .A2(new_n457), .ZN(new_n541));
  NAND3_X1  g0341(.A1(new_n541), .A2(G257), .A3(new_n251), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n542), .A2(new_n461), .ZN(new_n543));
  INV_X1    g0343(.A(new_n543), .ZN(new_n544));
  NAND3_X1  g0344(.A1(new_n540), .A2(G179), .A3(new_n544), .ZN(new_n545));
  AOI21_X1  g0345(.A(new_n543), .B1(new_n539), .B2(new_n252), .ZN(new_n546));
  OAI21_X1  g0346(.A(new_n545), .B1(new_n360), .B2(new_n546), .ZN(new_n547));
  INV_X1    g0347(.A(KEYINPUT78), .ZN(new_n548));
  INV_X1    g0348(.A(KEYINPUT6), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  AND2_X1   g0350(.A1(G97), .A2(G107), .ZN(new_n551));
  NOR2_X1   g0351(.A1(G97), .A2(G107), .ZN(new_n552));
  OAI21_X1  g0352(.A(new_n550), .B1(new_n551), .B2(new_n552), .ZN(new_n553));
  NOR2_X1   g0353(.A1(KEYINPUT78), .A2(KEYINPUT6), .ZN(new_n554));
  INV_X1    g0354(.A(G97), .ZN(new_n555));
  AOI21_X1  g0355(.A(new_n554), .B1(KEYINPUT6), .B2(new_n555), .ZN(new_n556));
  XNOR2_X1  g0356(.A(G97), .B(G107), .ZN(new_n557));
  OAI211_X1 g0357(.A(G20), .B(new_n553), .C1(new_n556), .C2(new_n557), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n271), .A2(G77), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  AOI21_X1  g0360(.A(new_n418), .B1(new_n340), .B2(new_n332), .ZN(new_n561));
  OAI21_X1  g0361(.A(new_n280), .B1(new_n560), .B2(new_n561), .ZN(new_n562));
  NOR2_X1   g0362(.A1(new_n511), .A2(G97), .ZN(new_n563));
  AOI21_X1  g0363(.A(new_n563), .B1(new_n479), .B2(G97), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n562), .A2(new_n564), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n565), .A2(KEYINPUT81), .ZN(new_n566));
  INV_X1    g0366(.A(KEYINPUT81), .ZN(new_n567));
  NAND3_X1  g0367(.A1(new_n562), .A2(new_n567), .A3(new_n564), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n566), .A2(new_n568), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n540), .A2(new_n544), .ZN(new_n570));
  INV_X1    g0370(.A(KEYINPUT80), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n546), .A2(KEYINPUT80), .ZN(new_n573));
  NAND3_X1  g0373(.A1(new_n572), .A2(G200), .A3(new_n573), .ZN(new_n574));
  AOI21_X1  g0374(.A(new_n565), .B1(G190), .B2(new_n546), .ZN(new_n575));
  AOI22_X1  g0375(.A1(new_n547), .A2(new_n569), .B1(new_n574), .B2(new_n575), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n497), .A2(new_n500), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n577), .A2(new_n280), .ZN(new_n578));
  OAI21_X1  g0378(.A(G200), .B1(new_n475), .B2(new_n476), .ZN(new_n579));
  OAI211_X1 g0379(.A(new_n462), .B(G190), .C1(new_n470), .C2(new_n251), .ZN(new_n580));
  NAND4_X1  g0380(.A1(new_n578), .A2(new_n579), .A3(new_n580), .A4(new_n483), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n213), .A2(new_n246), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n414), .A2(G1698), .ZN(new_n583));
  OAI211_X1 g0383(.A(new_n582), .B(new_n583), .C1(new_n319), .C2(new_n320), .ZN(new_n584));
  AOI21_X1  g0384(.A(new_n251), .B1(new_n584), .B2(new_n486), .ZN(new_n585));
  NAND3_X1  g0385(.A1(new_n251), .A2(G274), .A3(new_n457), .ZN(new_n586));
  AOI21_X1  g0386(.A(new_n215), .B1(new_n256), .B2(G45), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n587), .A2(new_n251), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n586), .A2(new_n588), .ZN(new_n589));
  OAI21_X1  g0389(.A(G200), .B1(new_n585), .B2(new_n589), .ZN(new_n590));
  INV_X1    g0390(.A(KEYINPUT19), .ZN(new_n591));
  OAI21_X1  g0391(.A(new_n269), .B1(new_n248), .B2(new_n591), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n552), .A2(new_n214), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  OAI211_X1 g0394(.A(new_n269), .B(G68), .C1(new_n319), .C2(new_n320), .ZN(new_n595));
  OAI21_X1  g0395(.A(new_n591), .B1(new_n274), .B2(new_n555), .ZN(new_n596));
  NAND3_X1  g0396(.A1(new_n594), .A2(new_n595), .A3(new_n596), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n426), .A2(new_n430), .ZN(new_n598));
  AOI22_X1  g0398(.A1(new_n280), .A2(new_n597), .B1(new_n598), .B2(new_n283), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n479), .A2(G87), .ZN(new_n600));
  AOI22_X1  g0400(.A1(new_n255), .A2(new_n457), .B1(new_n251), .B2(new_n587), .ZN(new_n601));
  NOR2_X1   g0401(.A1(G238), .A2(G1698), .ZN(new_n602));
  AOI21_X1  g0402(.A(new_n602), .B1(new_n414), .B2(G1698), .ZN(new_n603));
  AOI22_X1  g0403(.A1(new_n603), .A2(new_n244), .B1(G33), .B2(G116), .ZN(new_n604));
  OAI211_X1 g0404(.A(G190), .B(new_n601), .C1(new_n604), .C2(new_n251), .ZN(new_n605));
  AND4_X1   g0405(.A1(new_n590), .A2(new_n599), .A3(new_n600), .A4(new_n605), .ZN(new_n606));
  OAI211_X1 g0406(.A(new_n358), .B(new_n601), .C1(new_n604), .C2(new_n251), .ZN(new_n607));
  OAI21_X1  g0407(.A(new_n360), .B1(new_n585), .B2(new_n589), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  INV_X1    g0409(.A(KEYINPUT82), .ZN(new_n610));
  AND2_X1   g0410(.A1(new_n426), .A2(new_n430), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n479), .A2(new_n611), .ZN(new_n612));
  AOI22_X1  g0412(.A1(new_n609), .A2(new_n610), .B1(new_n599), .B2(new_n612), .ZN(new_n613));
  NAND3_X1  g0413(.A1(new_n607), .A2(new_n608), .A3(KEYINPUT82), .ZN(new_n614));
  AOI21_X1  g0414(.A(new_n606), .B1(new_n613), .B2(new_n614), .ZN(new_n615));
  INV_X1    g0415(.A(new_n525), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n508), .A2(new_n461), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n617), .A2(G200), .ZN(new_n618));
  NAND3_X1  g0418(.A1(new_n508), .A2(G190), .A3(new_n461), .ZN(new_n619));
  NAND3_X1  g0419(.A1(new_n616), .A2(new_n618), .A3(new_n619), .ZN(new_n620));
  AND3_X1   g0420(.A1(new_n581), .A2(new_n615), .A3(new_n620), .ZN(new_n621));
  AND4_X1   g0421(.A1(new_n455), .A2(new_n532), .A3(new_n576), .A4(new_n621), .ZN(G372));
  AOI21_X1  g0422(.A(KEYINPUT18), .B1(new_n348), .B2(new_n363), .ZN(new_n623));
  NOR3_X1   g0423(.A1(new_n367), .A2(new_n362), .A3(new_n365), .ZN(new_n624));
  NOR2_X1   g0424(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n298), .A2(new_n299), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n626), .A2(new_n450), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n307), .A2(new_n308), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  AOI21_X1  g0429(.A(new_n625), .B1(new_n629), .B2(new_n380), .ZN(new_n630));
  INV_X1    g0430(.A(new_n406), .ZN(new_n631));
  OAI21_X1  g0431(.A(new_n410), .B1(new_n630), .B2(new_n631), .ZN(new_n632));
  INV_X1    g0432(.A(new_n632), .ZN(new_n633));
  INV_X1    g0433(.A(new_n455), .ZN(new_n634));
  INV_X1    g0434(.A(KEYINPUT87), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n584), .A2(new_n486), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n636), .A2(new_n252), .ZN(new_n637));
  INV_X1    g0437(.A(KEYINPUT85), .ZN(new_n638));
  AND3_X1   g0438(.A1(new_n586), .A2(new_n588), .A3(new_n638), .ZN(new_n639));
  AOI21_X1  g0439(.A(new_n638), .B1(new_n586), .B2(new_n588), .ZN(new_n640));
  OAI21_X1  g0440(.A(new_n637), .B1(new_n639), .B2(new_n640), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n641), .A2(new_n360), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n599), .A2(new_n612), .ZN(new_n643));
  AND4_X1   g0443(.A1(KEYINPUT86), .A2(new_n642), .A3(new_n607), .A4(new_n643), .ZN(new_n644));
  NOR3_X1   g0444(.A1(new_n585), .A2(new_n589), .A3(G179), .ZN(new_n645));
  AOI21_X1  g0445(.A(new_n645), .B1(new_n599), .B2(new_n612), .ZN(new_n646));
  AOI21_X1  g0446(.A(KEYINPUT86), .B1(new_n646), .B2(new_n642), .ZN(new_n647));
  NOR2_X1   g0447(.A1(new_n644), .A2(new_n647), .ZN(new_n648));
  AND3_X1   g0448(.A1(new_n599), .A2(new_n600), .A3(new_n605), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n641), .A2(G200), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  NAND3_X1  g0451(.A1(new_n642), .A2(new_n643), .A3(new_n607), .ZN(new_n652));
  NAND4_X1  g0452(.A1(new_n547), .A2(new_n651), .A3(new_n565), .A4(new_n652), .ZN(new_n653));
  OAI21_X1  g0453(.A(new_n648), .B1(new_n653), .B2(KEYINPUT26), .ZN(new_n654));
  INV_X1    g0454(.A(KEYINPUT26), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n570), .A2(G169), .ZN(new_n656));
  AOI22_X1  g0456(.A1(new_n566), .A2(new_n568), .B1(new_n656), .B2(new_n545), .ZN(new_n657));
  AOI21_X1  g0457(.A(new_n655), .B1(new_n657), .B2(new_n615), .ZN(new_n658));
  OAI21_X1  g0458(.A(new_n635), .B1(new_n654), .B2(new_n658), .ZN(new_n659));
  INV_X1    g0459(.A(new_n568), .ZN(new_n660));
  AOI21_X1  g0460(.A(new_n567), .B1(new_n562), .B2(new_n564), .ZN(new_n661));
  OAI21_X1  g0461(.A(new_n547), .B1(new_n660), .B2(new_n661), .ZN(new_n662));
  AOI21_X1  g0462(.A(G169), .B1(new_n637), .B2(new_n601), .ZN(new_n663));
  OAI21_X1  g0463(.A(new_n610), .B1(new_n663), .B2(new_n645), .ZN(new_n664));
  NAND3_X1  g0464(.A1(new_n664), .A2(new_n614), .A3(new_n643), .ZN(new_n665));
  INV_X1    g0465(.A(new_n606), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  OAI21_X1  g0467(.A(KEYINPUT26), .B1(new_n662), .B2(new_n667), .ZN(new_n668));
  AOI22_X1  g0468(.A1(new_n649), .A2(new_n650), .B1(new_n646), .B2(new_n642), .ZN(new_n669));
  NAND4_X1  g0469(.A1(new_n669), .A2(new_n655), .A3(new_n547), .A4(new_n565), .ZN(new_n670));
  NAND4_X1  g0470(.A1(new_n668), .A2(KEYINPUT87), .A3(new_n670), .A4(new_n648), .ZN(new_n671));
  AND2_X1   g0471(.A1(new_n581), .A2(new_n669), .ZN(new_n672));
  NAND3_X1  g0472(.A1(new_n672), .A2(new_n531), .A3(new_n576), .ZN(new_n673));
  NAND3_X1  g0473(.A1(new_n659), .A2(new_n671), .A3(new_n673), .ZN(new_n674));
  INV_X1    g0474(.A(new_n674), .ZN(new_n675));
  OAI21_X1  g0475(.A(new_n633), .B1(new_n634), .B2(new_n675), .ZN(G369));
  NAND3_X1  g0476(.A1(new_n256), .A2(new_n269), .A3(G13), .ZN(new_n677));
  OR2_X1    g0477(.A1(new_n677), .A2(KEYINPUT27), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n677), .A2(KEYINPUT27), .ZN(new_n679));
  NAND3_X1  g0479(.A1(new_n678), .A2(G213), .A3(new_n679), .ZN(new_n680));
  INV_X1    g0480(.A(G343), .ZN(new_n681));
  NOR2_X1   g0481(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n525), .A2(new_n682), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n620), .A2(new_n683), .ZN(new_n684));
  NAND4_X1  g0484(.A1(new_n684), .A2(new_n528), .A3(new_n529), .A4(new_n530), .ZN(new_n685));
  NAND3_X1  g0485(.A1(new_n528), .A2(new_n529), .A3(new_n530), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n686), .A2(new_n683), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n685), .A2(new_n687), .ZN(new_n688));
  INV_X1    g0488(.A(KEYINPUT88), .ZN(new_n689));
  XNOR2_X1  g0489(.A(new_n688), .B(new_n689), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n690), .A2(G330), .ZN(new_n691));
  NOR2_X1   g0491(.A1(new_n502), .A2(new_n682), .ZN(new_n692));
  INV_X1    g0492(.A(new_n502), .ZN(new_n693));
  OAI21_X1  g0493(.A(new_n682), .B1(new_n484), .B2(new_n501), .ZN(new_n694));
  AOI21_X1  g0494(.A(new_n693), .B1(new_n694), .B2(new_n581), .ZN(new_n695));
  NOR3_X1   g0495(.A1(new_n691), .A2(new_n692), .A3(new_n695), .ZN(new_n696));
  INV_X1    g0496(.A(new_n696), .ZN(new_n697));
  INV_X1    g0497(.A(new_n682), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n686), .A2(new_n698), .ZN(new_n699));
  OAI22_X1  g0499(.A1(new_n695), .A2(new_n699), .B1(new_n502), .B2(new_n682), .ZN(new_n700));
  INV_X1    g0500(.A(new_n700), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n697), .A2(new_n701), .ZN(G399));
  INV_X1    g0502(.A(new_n205), .ZN(new_n703));
  NOR2_X1   g0503(.A1(new_n703), .A2(G41), .ZN(new_n704));
  INV_X1    g0504(.A(new_n704), .ZN(new_n705));
  NOR2_X1   g0505(.A1(new_n593), .A2(G116), .ZN(new_n706));
  NAND3_X1  g0506(.A1(new_n705), .A2(G1), .A3(new_n706), .ZN(new_n707));
  INV_X1    g0507(.A(KEYINPUT89), .ZN(new_n708));
  OAI22_X1  g0508(.A1(new_n707), .A2(new_n708), .B1(new_n210), .B2(new_n705), .ZN(new_n709));
  AOI21_X1  g0509(.A(new_n709), .B1(new_n708), .B2(new_n707), .ZN(new_n710));
  XOR2_X1   g0510(.A(new_n710), .B(KEYINPUT28), .Z(new_n711));
  INV_X1    g0511(.A(KEYINPUT29), .ZN(new_n712));
  INV_X1    g0512(.A(new_n648), .ZN(new_n713));
  NOR3_X1   g0513(.A1(new_n662), .A2(new_n667), .A3(KEYINPUT26), .ZN(new_n714));
  AOI211_X1 g0514(.A(new_n713), .B(new_n714), .C1(KEYINPUT26), .C2(new_n653), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n576), .A2(KEYINPUT90), .ZN(new_n716));
  INV_X1    g0516(.A(KEYINPUT90), .ZN(new_n717));
  AND2_X1   g0517(.A1(new_n574), .A2(new_n575), .ZN(new_n718));
  OAI21_X1  g0518(.A(new_n717), .B1(new_n718), .B2(new_n657), .ZN(new_n719));
  NAND4_X1  g0519(.A1(new_n716), .A2(new_n719), .A3(new_n531), .A4(new_n672), .ZN(new_n720));
  AOI211_X1 g0520(.A(new_n712), .B(new_n682), .C1(new_n715), .C2(new_n720), .ZN(new_n721));
  AOI21_X1  g0521(.A(KEYINPUT29), .B1(new_n674), .B2(new_n698), .ZN(new_n722));
  NOR2_X1   g0522(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  NAND4_X1  g0523(.A1(new_n532), .A2(new_n576), .A3(new_n621), .A4(new_n698), .ZN(new_n724));
  INV_X1    g0524(.A(new_n545), .ZN(new_n725));
  NAND2_X1  g0525(.A1(new_n472), .A2(new_n474), .ZN(new_n726));
  AOI21_X1  g0526(.A(new_n476), .B1(new_n726), .B2(new_n252), .ZN(new_n727));
  NOR2_X1   g0527(.A1(new_n585), .A2(new_n589), .ZN(new_n728));
  AND2_X1   g0528(.A1(new_n508), .A2(new_n728), .ZN(new_n729));
  NAND3_X1  g0529(.A1(new_n725), .A2(new_n727), .A3(new_n729), .ZN(new_n730));
  INV_X1    g0530(.A(KEYINPUT30), .ZN(new_n731));
  NAND2_X1  g0531(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  NAND4_X1  g0532(.A1(new_n725), .A2(new_n729), .A3(new_n727), .A4(KEYINPUT30), .ZN(new_n733));
  INV_X1    g0533(.A(new_n727), .ZN(new_n734));
  AND2_X1   g0534(.A1(new_n641), .A2(new_n358), .ZN(new_n735));
  NAND4_X1  g0535(.A1(new_n734), .A2(new_n617), .A3(new_n570), .A4(new_n735), .ZN(new_n736));
  NAND3_X1  g0536(.A1(new_n732), .A2(new_n733), .A3(new_n736), .ZN(new_n737));
  NAND2_X1  g0537(.A1(new_n737), .A2(new_n682), .ZN(new_n738));
  INV_X1    g0538(.A(KEYINPUT31), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  NAND3_X1  g0540(.A1(new_n737), .A2(KEYINPUT31), .A3(new_n682), .ZN(new_n741));
  NAND3_X1  g0541(.A1(new_n724), .A2(new_n740), .A3(new_n741), .ZN(new_n742));
  NAND2_X1  g0542(.A1(new_n742), .A2(G330), .ZN(new_n743));
  INV_X1    g0543(.A(new_n743), .ZN(new_n744));
  NOR2_X1   g0544(.A1(new_n723), .A2(new_n744), .ZN(new_n745));
  OAI21_X1  g0545(.A(new_n711), .B1(new_n745), .B2(G1), .ZN(G364));
  NOR2_X1   g0546(.A1(new_n690), .A2(G330), .ZN(new_n747));
  AND2_X1   g0547(.A1(new_n690), .A2(G330), .ZN(new_n748));
  NOR2_X1   g0548(.A1(new_n282), .A2(G20), .ZN(new_n749));
  AOI21_X1  g0549(.A(new_n256), .B1(new_n749), .B2(G45), .ZN(new_n750));
  AOI211_X1 g0550(.A(new_n747), .B(new_n748), .C1(new_n705), .C2(new_n750), .ZN(new_n751));
  INV_X1    g0551(.A(new_n750), .ZN(new_n752));
  NOR2_X1   g0552(.A1(new_n704), .A2(new_n752), .ZN(new_n753));
  XOR2_X1   g0553(.A(new_n753), .B(KEYINPUT91), .Z(new_n754));
  NAND2_X1  g0554(.A1(new_n244), .A2(new_n205), .ZN(new_n755));
  INV_X1    g0555(.A(G355), .ZN(new_n756));
  OAI22_X1  g0556(.A1(new_n755), .A2(new_n756), .B1(G116), .B2(new_n205), .ZN(new_n757));
  OR2_X1    g0557(.A1(new_n234), .A2(new_n456), .ZN(new_n758));
  NOR2_X1   g0558(.A1(new_n703), .A2(new_n244), .ZN(new_n759));
  INV_X1    g0559(.A(new_n759), .ZN(new_n760));
  INV_X1    g0560(.A(new_n210), .ZN(new_n761));
  AOI21_X1  g0561(.A(new_n760), .B1(new_n456), .B2(new_n761), .ZN(new_n762));
  AOI21_X1  g0562(.A(new_n757), .B1(new_n758), .B2(new_n762), .ZN(new_n763));
  OAI21_X1  g0563(.A(new_n208), .B1(new_n269), .B2(G169), .ZN(new_n764));
  XNOR2_X1  g0564(.A(new_n764), .B(KEYINPUT92), .ZN(new_n765));
  INV_X1    g0565(.A(new_n765), .ZN(new_n766));
  NOR2_X1   g0566(.A1(G13), .A2(G33), .ZN(new_n767));
  INV_X1    g0567(.A(new_n767), .ZN(new_n768));
  NOR2_X1   g0568(.A1(new_n768), .A2(G20), .ZN(new_n769));
  NOR2_X1   g0569(.A1(new_n766), .A2(new_n769), .ZN(new_n770));
  INV_X1    g0570(.A(new_n770), .ZN(new_n771));
  OAI21_X1  g0571(.A(new_n754), .B1(new_n763), .B2(new_n771), .ZN(new_n772));
  NOR2_X1   g0572(.A1(new_n269), .A2(new_n358), .ZN(new_n773));
  INV_X1    g0573(.A(new_n773), .ZN(new_n774));
  NOR3_X1   g0574(.A1(new_n774), .A2(new_n370), .A3(new_n373), .ZN(new_n775));
  INV_X1    g0575(.A(new_n775), .ZN(new_n776));
  NOR2_X1   g0576(.A1(G190), .A2(G200), .ZN(new_n777));
  NAND2_X1  g0577(.A1(new_n773), .A2(new_n777), .ZN(new_n778));
  OAI22_X1  g0578(.A1(new_n776), .A2(new_n388), .B1(new_n778), .B2(new_n273), .ZN(new_n779));
  NAND3_X1  g0579(.A1(new_n773), .A2(new_n370), .A3(G200), .ZN(new_n780));
  INV_X1    g0580(.A(new_n780), .ZN(new_n781));
  AOI211_X1 g0581(.A(new_n505), .B(new_n779), .C1(G68), .C2(new_n781), .ZN(new_n782));
  NOR2_X1   g0582(.A1(new_n269), .A2(G179), .ZN(new_n783));
  NAND3_X1  g0583(.A1(new_n783), .A2(G190), .A3(G200), .ZN(new_n784));
  NOR2_X1   g0584(.A1(new_n784), .A2(new_n214), .ZN(new_n785));
  NAND2_X1  g0585(.A1(new_n783), .A2(new_n777), .ZN(new_n786));
  NOR2_X1   g0586(.A1(new_n786), .A2(new_n311), .ZN(new_n787));
  INV_X1    g0587(.A(new_n787), .ZN(new_n788));
  NOR2_X1   g0588(.A1(new_n788), .A2(KEYINPUT32), .ZN(new_n789));
  NAND3_X1  g0589(.A1(new_n783), .A2(new_n370), .A3(G200), .ZN(new_n790));
  INV_X1    g0590(.A(new_n790), .ZN(new_n791));
  AOI211_X1 g0591(.A(new_n785), .B(new_n789), .C1(G107), .C2(new_n791), .ZN(new_n792));
  NOR3_X1   g0592(.A1(new_n774), .A2(new_n370), .A3(G200), .ZN(new_n793));
  XOR2_X1   g0593(.A(new_n793), .B(KEYINPUT93), .Z(new_n794));
  INV_X1    g0594(.A(new_n794), .ZN(new_n795));
  NAND2_X1  g0595(.A1(new_n795), .A2(G58), .ZN(new_n796));
  NOR3_X1   g0596(.A1(new_n370), .A2(G179), .A3(G200), .ZN(new_n797));
  NOR2_X1   g0597(.A1(new_n797), .A2(new_n269), .ZN(new_n798));
  INV_X1    g0598(.A(new_n798), .ZN(new_n799));
  AOI22_X1  g0599(.A1(new_n788), .A2(KEYINPUT32), .B1(new_n799), .B2(G97), .ZN(new_n800));
  NAND4_X1  g0600(.A1(new_n782), .A2(new_n792), .A3(new_n796), .A4(new_n800), .ZN(new_n801));
  OR2_X1    g0601(.A1(new_n801), .A2(KEYINPUT94), .ZN(new_n802));
  INV_X1    g0602(.A(G303), .ZN(new_n803));
  NOR2_X1   g0603(.A1(new_n784), .A2(new_n803), .ZN(new_n804));
  AOI211_X1 g0604(.A(new_n244), .B(new_n804), .C1(G326), .C2(new_n775), .ZN(new_n805));
  INV_X1    g0605(.A(new_n786), .ZN(new_n806));
  AOI22_X1  g0606(.A1(new_n793), .A2(G322), .B1(G329), .B2(new_n806), .ZN(new_n807));
  XNOR2_X1  g0607(.A(KEYINPUT33), .B(G317), .ZN(new_n808));
  INV_X1    g0608(.A(new_n778), .ZN(new_n809));
  AOI22_X1  g0609(.A1(new_n781), .A2(new_n808), .B1(new_n809), .B2(G311), .ZN(new_n810));
  AOI22_X1  g0610(.A1(new_n799), .A2(G294), .B1(new_n791), .B2(G283), .ZN(new_n811));
  NAND4_X1  g0611(.A1(new_n805), .A2(new_n807), .A3(new_n810), .A4(new_n811), .ZN(new_n812));
  NAND2_X1  g0612(.A1(new_n801), .A2(KEYINPUT94), .ZN(new_n813));
  NAND3_X1  g0613(.A1(new_n802), .A2(new_n812), .A3(new_n813), .ZN(new_n814));
  AOI21_X1  g0614(.A(new_n772), .B1(new_n814), .B2(new_n766), .ZN(new_n815));
  INV_X1    g0615(.A(new_n769), .ZN(new_n816));
  OAI21_X1  g0616(.A(new_n815), .B1(new_n690), .B2(new_n816), .ZN(new_n817));
  XNOR2_X1  g0617(.A(new_n817), .B(KEYINPUT95), .ZN(new_n818));
  NOR2_X1   g0618(.A1(new_n751), .A2(new_n818), .ZN(new_n819));
  INV_X1    g0619(.A(new_n819), .ZN(G396));
  NAND2_X1  g0620(.A1(new_n450), .A2(new_n698), .ZN(new_n821));
  INV_X1    g0621(.A(new_n821), .ZN(new_n822));
  AOI21_X1  g0622(.A(new_n698), .B1(new_n439), .B2(new_n440), .ZN(new_n823));
  INV_X1    g0623(.A(new_n823), .ZN(new_n824));
  NAND2_X1  g0624(.A1(new_n446), .A2(new_n824), .ZN(new_n825));
  AOI21_X1  g0625(.A(new_n822), .B1(new_n825), .B2(new_n451), .ZN(new_n826));
  AOI21_X1  g0626(.A(new_n826), .B1(new_n674), .B2(new_n698), .ZN(new_n827));
  INV_X1    g0627(.A(KEYINPUT97), .ZN(new_n828));
  AOI211_X1 g0628(.A(new_n682), .B(new_n450), .C1(new_n443), .C2(new_n445), .ZN(new_n829));
  NAND3_X1  g0629(.A1(new_n674), .A2(new_n828), .A3(new_n829), .ZN(new_n830));
  NAND2_X1  g0630(.A1(new_n674), .A2(new_n829), .ZN(new_n831));
  NAND2_X1  g0631(.A1(new_n831), .A2(KEYINPUT97), .ZN(new_n832));
  AOI21_X1  g0632(.A(new_n827), .B1(new_n830), .B2(new_n832), .ZN(new_n833));
  NAND2_X1  g0633(.A1(new_n833), .A2(new_n744), .ZN(new_n834));
  INV_X1    g0634(.A(new_n834), .ZN(new_n835));
  OAI22_X1  g0635(.A1(new_n833), .A2(new_n744), .B1(new_n704), .B2(new_n752), .ZN(new_n836));
  NOR2_X1   g0636(.A1(new_n826), .A2(new_n768), .ZN(new_n837));
  NAND2_X1  g0637(.A1(new_n765), .A2(new_n768), .ZN(new_n838));
  XNOR2_X1  g0638(.A(new_n838), .B(KEYINPUT96), .ZN(new_n839));
  AOI22_X1  g0639(.A1(G116), .A2(new_n809), .B1(new_n806), .B2(G311), .ZN(new_n840));
  INV_X1    g0640(.A(G283), .ZN(new_n841));
  INV_X1    g0641(.A(new_n793), .ZN(new_n842));
  OAI221_X1 g0642(.A(new_n840), .B1(new_n841), .B2(new_n780), .C1(new_n464), .C2(new_n842), .ZN(new_n843));
  OAI221_X1 g0643(.A(new_n505), .B1(new_n555), .B2(new_n798), .C1(new_n776), .C2(new_n803), .ZN(new_n844));
  NOR2_X1   g0644(.A1(new_n784), .A2(new_n418), .ZN(new_n845));
  NOR2_X1   g0645(.A1(new_n790), .A2(new_n214), .ZN(new_n846));
  NOR4_X1   g0646(.A1(new_n843), .A2(new_n844), .A3(new_n845), .A4(new_n846), .ZN(new_n847));
  AOI22_X1  g0647(.A1(new_n775), .A2(G137), .B1(G159), .B2(new_n809), .ZN(new_n848));
  INV_X1    g0648(.A(G143), .ZN(new_n849));
  OAI221_X1 g0649(.A(new_n848), .B1(new_n383), .B2(new_n780), .C1(new_n794), .C2(new_n849), .ZN(new_n850));
  XNOR2_X1  g0650(.A(new_n850), .B(KEYINPUT34), .ZN(new_n851));
  INV_X1    g0651(.A(G132), .ZN(new_n852));
  OAI21_X1  g0652(.A(new_n244), .B1(new_n786), .B2(new_n852), .ZN(new_n853));
  OAI22_X1  g0653(.A1(new_n388), .A2(new_n784), .B1(new_n790), .B2(new_n212), .ZN(new_n854));
  AOI211_X1 g0654(.A(new_n853), .B(new_n854), .C1(G58), .C2(new_n799), .ZN(new_n855));
  AOI21_X1  g0655(.A(new_n847), .B1(new_n851), .B2(new_n855), .ZN(new_n856));
  OAI221_X1 g0656(.A(new_n754), .B1(G77), .B2(new_n839), .C1(new_n856), .C2(new_n765), .ZN(new_n857));
  OAI22_X1  g0657(.A1(new_n835), .A2(new_n836), .B1(new_n837), .B2(new_n857), .ZN(G384));
  NOR2_X1   g0658(.A1(new_n749), .A2(new_n256), .ZN(new_n859));
  AOI21_X1  g0659(.A(new_n823), .B1(new_n443), .B2(new_n445), .ZN(new_n860));
  OAI21_X1  g0660(.A(new_n821), .B1(new_n860), .B2(new_n450), .ZN(new_n861));
  OAI211_X1 g0661(.A(new_n626), .B(new_n628), .C1(new_n295), .C2(new_n698), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n626), .A2(new_n628), .ZN(new_n863));
  NOR2_X1   g0663(.A1(new_n295), .A2(new_n698), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  AOI21_X1  g0665(.A(new_n861), .B1(new_n862), .B2(new_n865), .ZN(new_n866));
  INV_X1    g0666(.A(KEYINPUT102), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n742), .A2(new_n867), .ZN(new_n868));
  NAND4_X1  g0668(.A1(new_n724), .A2(new_n740), .A3(KEYINPUT102), .A4(new_n741), .ZN(new_n869));
  NAND4_X1  g0669(.A1(new_n866), .A2(new_n868), .A3(KEYINPUT40), .A4(new_n869), .ZN(new_n870));
  INV_X1    g0670(.A(new_n680), .ZN(new_n871));
  OAI21_X1  g0671(.A(new_n318), .B1(new_n323), .B2(new_n329), .ZN(new_n872));
  AND2_X1   g0672(.A1(new_n872), .A2(new_n337), .ZN(new_n873));
  OAI21_X1  g0673(.A(new_n347), .B1(new_n873), .B2(new_n331), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n367), .A2(new_n377), .ZN(new_n875));
  INV_X1    g0675(.A(KEYINPUT17), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  NAND3_X1  g0677(.A1(new_n367), .A2(KEYINPUT17), .A3(new_n377), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n877), .A2(new_n878), .ZN(new_n879));
  OAI211_X1 g0679(.A(new_n871), .B(new_n874), .C1(new_n625), .C2(new_n879), .ZN(new_n880));
  NOR3_X1   g0680(.A1(new_n359), .A2(new_n361), .A3(new_n871), .ZN(new_n881));
  INV_X1    g0681(.A(new_n881), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n348), .A2(new_n882), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n883), .A2(new_n875), .ZN(new_n884));
  INV_X1    g0684(.A(KEYINPUT37), .ZN(new_n885));
  AOI21_X1  g0685(.A(new_n885), .B1(new_n882), .B2(new_n874), .ZN(new_n886));
  AOI22_X1  g0686(.A1(new_n884), .A2(new_n885), .B1(new_n886), .B2(new_n875), .ZN(new_n887));
  AND3_X1   g0687(.A1(new_n880), .A2(KEYINPUT38), .A3(new_n887), .ZN(new_n888));
  OAI21_X1  g0688(.A(KEYINPUT100), .B1(new_n367), .B2(new_n881), .ZN(new_n889));
  AND4_X1   g0689(.A1(KEYINPUT37), .A2(new_n883), .A3(new_n889), .A4(new_n875), .ZN(new_n890));
  AOI22_X1  g0690(.A1(new_n875), .A2(new_n883), .B1(new_n889), .B2(KEYINPUT37), .ZN(new_n891));
  NOR2_X1   g0691(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  OAI211_X1 g0692(.A(new_n348), .B(new_n871), .C1(new_n625), .C2(new_n879), .ZN(new_n893));
  AOI21_X1  g0693(.A(KEYINPUT38), .B1(new_n892), .B2(new_n893), .ZN(new_n894));
  NOR2_X1   g0694(.A1(new_n888), .A2(new_n894), .ZN(new_n895));
  NOR2_X1   g0695(.A1(new_n870), .A2(new_n895), .ZN(new_n896));
  AND3_X1   g0696(.A1(new_n866), .A2(new_n868), .A3(new_n869), .ZN(new_n897));
  AOI21_X1  g0697(.A(KEYINPUT38), .B1(new_n880), .B2(new_n887), .ZN(new_n898));
  NOR3_X1   g0698(.A1(new_n888), .A2(new_n898), .A3(KEYINPUT99), .ZN(new_n899));
  INV_X1    g0699(.A(KEYINPUT99), .ZN(new_n900));
  INV_X1    g0700(.A(KEYINPUT38), .ZN(new_n901));
  INV_X1    g0701(.A(new_n874), .ZN(new_n902));
  AOI211_X1 g0702(.A(new_n680), .B(new_n902), .C1(new_n380), .C2(new_n369), .ZN(new_n903));
  INV_X1    g0703(.A(new_n887), .ZN(new_n904));
  OAI21_X1  g0704(.A(new_n901), .B1(new_n903), .B2(new_n904), .ZN(new_n905));
  NAND3_X1  g0705(.A1(new_n880), .A2(KEYINPUT38), .A3(new_n887), .ZN(new_n906));
  AOI21_X1  g0706(.A(new_n900), .B1(new_n905), .B2(new_n906), .ZN(new_n907));
  OAI21_X1  g0707(.A(new_n897), .B1(new_n899), .B2(new_n907), .ZN(new_n908));
  INV_X1    g0708(.A(KEYINPUT40), .ZN(new_n909));
  AOI21_X1  g0709(.A(new_n896), .B1(new_n908), .B2(new_n909), .ZN(new_n910));
  INV_X1    g0710(.A(new_n910), .ZN(new_n911));
  AND2_X1   g0711(.A1(new_n868), .A2(new_n869), .ZN(new_n912));
  INV_X1    g0712(.A(new_n912), .ZN(new_n913));
  OAI21_X1  g0713(.A(new_n911), .B1(new_n634), .B2(new_n913), .ZN(new_n914));
  NAND3_X1  g0714(.A1(new_n910), .A2(new_n455), .A3(new_n912), .ZN(new_n915));
  NAND3_X1  g0715(.A1(new_n914), .A2(G330), .A3(new_n915), .ZN(new_n916));
  XNOR2_X1  g0716(.A(new_n916), .B(KEYINPUT103), .ZN(new_n917));
  INV_X1    g0717(.A(new_n917), .ZN(new_n918));
  INV_X1    g0718(.A(KEYINPUT39), .ZN(new_n919));
  OAI21_X1  g0719(.A(new_n919), .B1(new_n888), .B2(new_n894), .ZN(new_n920));
  NOR2_X1   g0720(.A1(new_n628), .A2(new_n682), .ZN(new_n921));
  NAND3_X1  g0721(.A1(new_n905), .A2(KEYINPUT39), .A3(new_n906), .ZN(new_n922));
  NAND3_X1  g0722(.A1(new_n920), .A2(new_n921), .A3(new_n922), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n625), .A2(new_n680), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  INV_X1    g0725(.A(new_n925), .ZN(new_n926));
  INV_X1    g0726(.A(KEYINPUT101), .ZN(new_n927));
  AND2_X1   g0727(.A1(new_n865), .A2(new_n862), .ZN(new_n928));
  INV_X1    g0728(.A(new_n928), .ZN(new_n929));
  OAI21_X1  g0729(.A(KEYINPUT99), .B1(new_n888), .B2(new_n898), .ZN(new_n930));
  NAND3_X1  g0730(.A1(new_n905), .A2(new_n900), .A3(new_n906), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  INV_X1    g0732(.A(KEYINPUT98), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n832), .A2(new_n830), .ZN(new_n934));
  AOI21_X1  g0734(.A(new_n933), .B1(new_n934), .B2(new_n821), .ZN(new_n935));
  AND3_X1   g0735(.A1(new_n674), .A2(new_n828), .A3(new_n829), .ZN(new_n936));
  AOI21_X1  g0736(.A(new_n828), .B1(new_n674), .B2(new_n829), .ZN(new_n937));
  OAI211_X1 g0737(.A(new_n933), .B(new_n821), .C1(new_n936), .C2(new_n937), .ZN(new_n938));
  INV_X1    g0738(.A(new_n938), .ZN(new_n939));
  OAI211_X1 g0739(.A(new_n929), .B(new_n932), .C1(new_n935), .C2(new_n939), .ZN(new_n940));
  AND3_X1   g0740(.A1(new_n926), .A2(new_n927), .A3(new_n940), .ZN(new_n941));
  AOI21_X1  g0741(.A(new_n927), .B1(new_n926), .B2(new_n940), .ZN(new_n942));
  NOR2_X1   g0742(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  AOI21_X1  g0743(.A(new_n632), .B1(new_n723), .B2(new_n455), .ZN(new_n944));
  XOR2_X1   g0744(.A(new_n943), .B(new_n944), .Z(new_n945));
  AOI21_X1  g0745(.A(new_n859), .B1(new_n918), .B2(new_n945), .ZN(new_n946));
  OAI21_X1  g0746(.A(new_n946), .B1(new_n918), .B2(new_n945), .ZN(new_n947));
  NOR2_X1   g0747(.A1(new_n209), .A2(new_n520), .ZN(new_n948));
  OAI21_X1  g0748(.A(new_n553), .B1(new_n556), .B2(new_n557), .ZN(new_n949));
  INV_X1    g0749(.A(KEYINPUT35), .ZN(new_n950));
  OAI21_X1  g0750(.A(new_n948), .B1(new_n949), .B2(new_n950), .ZN(new_n951));
  AOI21_X1  g0751(.A(new_n951), .B1(new_n950), .B2(new_n949), .ZN(new_n952));
  XOR2_X1   g0752(.A(new_n952), .B(KEYINPUT36), .Z(new_n953));
  NAND4_X1  g0753(.A1(new_n761), .A2(G77), .A3(new_n316), .A4(new_n314), .ZN(new_n954));
  OAI21_X1  g0754(.A(new_n954), .B1(G50), .B2(new_n212), .ZN(new_n955));
  NAND3_X1  g0755(.A1(new_n955), .A2(G1), .A3(new_n282), .ZN(new_n956));
  NAND3_X1  g0756(.A1(new_n947), .A2(new_n953), .A3(new_n956), .ZN(new_n957));
  XNOR2_X1  g0757(.A(new_n957), .B(KEYINPUT104), .ZN(G367));
  OAI221_X1 g0758(.A(new_n770), .B1(new_n205), .B2(new_n598), .C1(new_n230), .C2(new_n760), .ZN(new_n959));
  AND2_X1   g0759(.A1(new_n959), .A2(new_n754), .ZN(new_n960));
  OAI21_X1  g0760(.A(new_n244), .B1(new_n780), .B2(new_n311), .ZN(new_n961));
  INV_X1    g0761(.A(new_n784), .ZN(new_n962));
  AOI21_X1  g0762(.A(new_n961), .B1(G58), .B2(new_n962), .ZN(new_n963));
  AOI22_X1  g0763(.A1(new_n793), .A2(G150), .B1(new_n775), .B2(G143), .ZN(new_n964));
  AOI22_X1  g0764(.A1(G50), .A2(new_n809), .B1(new_n806), .B2(G137), .ZN(new_n965));
  NOR2_X1   g0765(.A1(new_n790), .A2(new_n273), .ZN(new_n966));
  AOI21_X1  g0766(.A(new_n966), .B1(G68), .B2(new_n799), .ZN(new_n967));
  NAND4_X1  g0767(.A1(new_n963), .A2(new_n964), .A3(new_n965), .A4(new_n967), .ZN(new_n968));
  AOI22_X1  g0768(.A1(new_n775), .A2(G311), .B1(new_n781), .B2(G294), .ZN(new_n969));
  INV_X1    g0769(.A(G317), .ZN(new_n970));
  OAI21_X1  g0770(.A(new_n969), .B1(new_n970), .B2(new_n786), .ZN(new_n971));
  NOR2_X1   g0771(.A1(new_n784), .A2(new_n520), .ZN(new_n972));
  AOI21_X1  g0772(.A(new_n971), .B1(KEYINPUT46), .B2(new_n972), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n791), .A2(G97), .ZN(new_n974));
  OAI211_X1 g0774(.A(new_n974), .B(new_n505), .C1(new_n841), .C2(new_n778), .ZN(new_n975));
  AOI21_X1  g0775(.A(new_n975), .B1(G107), .B2(new_n799), .ZN(new_n976));
  OAI211_X1 g0776(.A(new_n973), .B(new_n976), .C1(new_n803), .C2(new_n794), .ZN(new_n977));
  NOR2_X1   g0777(.A1(new_n972), .A2(KEYINPUT46), .ZN(new_n978));
  XNOR2_X1  g0778(.A(new_n978), .B(KEYINPUT107), .ZN(new_n979));
  OAI21_X1  g0779(.A(new_n968), .B1(new_n977), .B2(new_n979), .ZN(new_n980));
  INV_X1    g0780(.A(KEYINPUT47), .ZN(new_n981));
  AND2_X1   g0781(.A1(new_n980), .A2(new_n981), .ZN(new_n982));
  OAI21_X1  g0782(.A(new_n766), .B1(new_n980), .B2(new_n981), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n599), .A2(new_n600), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n984), .A2(new_n682), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n669), .A2(new_n985), .ZN(new_n986));
  OR2_X1    g0786(.A1(new_n986), .A2(KEYINPUT105), .ZN(new_n987));
  OAI211_X1 g0787(.A(new_n986), .B(KEYINPUT105), .C1(new_n648), .C2(new_n985), .ZN(new_n988));
  NAND2_X1  g0788(.A1(new_n987), .A2(new_n988), .ZN(new_n989));
  INV_X1    g0789(.A(new_n989), .ZN(new_n990));
  OAI221_X1 g0790(.A(new_n960), .B1(new_n982), .B2(new_n983), .C1(new_n990), .C2(new_n816), .ZN(new_n991));
  NAND2_X1  g0791(.A1(new_n565), .A2(new_n682), .ZN(new_n992));
  NAND3_X1  g0792(.A1(new_n716), .A2(new_n719), .A3(new_n992), .ZN(new_n993));
  NAND3_X1  g0793(.A1(new_n547), .A2(new_n565), .A3(new_n682), .ZN(new_n994));
  AND2_X1   g0794(.A1(new_n993), .A2(new_n994), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n995), .A2(new_n700), .ZN(new_n996));
  XOR2_X1   g0796(.A(new_n996), .B(KEYINPUT44), .Z(new_n997));
  NAND2_X1  g0797(.A1(new_n993), .A2(new_n994), .ZN(new_n998));
  NAND3_X1  g0798(.A1(new_n701), .A2(new_n998), .A3(KEYINPUT45), .ZN(new_n999));
  INV_X1    g0799(.A(new_n999), .ZN(new_n1000));
  AOI21_X1  g0800(.A(KEYINPUT45), .B1(new_n701), .B2(new_n998), .ZN(new_n1001));
  NOR2_X1   g0801(.A1(new_n1000), .A2(new_n1001), .ZN(new_n1002));
  INV_X1    g0802(.A(new_n1002), .ZN(new_n1003));
  AOI21_X1  g0803(.A(new_n697), .B1(new_n997), .B2(new_n1003), .ZN(new_n1004));
  XNOR2_X1  g0804(.A(new_n996), .B(KEYINPUT44), .ZN(new_n1005));
  NOR3_X1   g0805(.A1(new_n1005), .A2(new_n696), .A3(new_n1002), .ZN(new_n1006));
  NOR2_X1   g0806(.A1(new_n1004), .A2(new_n1006), .ZN(new_n1007));
  NOR2_X1   g0807(.A1(new_n695), .A2(new_n692), .ZN(new_n1008));
  XNOR2_X1  g0808(.A(new_n1008), .B(new_n699), .ZN(new_n1009));
  XNOR2_X1  g0809(.A(new_n691), .B(new_n1009), .ZN(new_n1010));
  NAND2_X1  g0810(.A1(new_n745), .A2(new_n1010), .ZN(new_n1011));
  INV_X1    g0811(.A(new_n1011), .ZN(new_n1012));
  NAND2_X1  g0812(.A1(new_n1007), .A2(new_n1012), .ZN(new_n1013));
  NAND2_X1  g0813(.A1(new_n1013), .A2(new_n745), .ZN(new_n1014));
  XNOR2_X1  g0814(.A(new_n704), .B(KEYINPUT41), .ZN(new_n1015));
  AOI21_X1  g0815(.A(new_n752), .B1(new_n1014), .B2(new_n1015), .ZN(new_n1016));
  NAND4_X1  g0816(.A1(new_n998), .A2(new_n686), .A3(new_n698), .A4(new_n1008), .ZN(new_n1017));
  INV_X1    g0817(.A(KEYINPUT42), .ZN(new_n1018));
  AND2_X1   g0818(.A1(new_n1017), .A2(new_n1018), .ZN(new_n1019));
  NOR2_X1   g0819(.A1(new_n1017), .A2(new_n1018), .ZN(new_n1020));
  AOI21_X1  g0820(.A(new_n657), .B1(new_n998), .B2(new_n693), .ZN(new_n1021));
  OAI22_X1  g0821(.A1(new_n1019), .A2(new_n1020), .B1(new_n1021), .B2(new_n682), .ZN(new_n1022));
  OR3_X1    g0822(.A1(new_n1022), .A2(KEYINPUT43), .A3(new_n990), .ZN(new_n1023));
  XNOR2_X1  g0823(.A(new_n989), .B(KEYINPUT43), .ZN(new_n1024));
  NAND2_X1  g0824(.A1(new_n1022), .A2(new_n1024), .ZN(new_n1025));
  NAND2_X1  g0825(.A1(new_n1025), .A2(KEYINPUT106), .ZN(new_n1026));
  INV_X1    g0826(.A(KEYINPUT106), .ZN(new_n1027));
  NAND3_X1  g0827(.A1(new_n1022), .A2(new_n1027), .A3(new_n1024), .ZN(new_n1028));
  NAND3_X1  g0828(.A1(new_n1023), .A2(new_n1026), .A3(new_n1028), .ZN(new_n1029));
  OAI21_X1  g0829(.A(new_n1029), .B1(new_n697), .B2(new_n995), .ZN(new_n1030));
  NOR2_X1   g0830(.A1(new_n697), .A2(new_n995), .ZN(new_n1031));
  NAND4_X1  g0831(.A1(new_n1023), .A2(new_n1026), .A3(new_n1031), .A4(new_n1028), .ZN(new_n1032));
  NAND2_X1  g0832(.A1(new_n1030), .A2(new_n1032), .ZN(new_n1033));
  OAI21_X1  g0833(.A(new_n991), .B1(new_n1016), .B2(new_n1033), .ZN(G387));
  OAI21_X1  g0834(.A(KEYINPUT108), .B1(new_n745), .B2(new_n1010), .ZN(new_n1035));
  OR2_X1    g0835(.A1(new_n721), .A2(new_n722), .ZN(new_n1036));
  NAND2_X1  g0836(.A1(new_n1036), .A2(new_n743), .ZN(new_n1037));
  XNOR2_X1  g0837(.A(new_n748), .B(new_n1009), .ZN(new_n1038));
  INV_X1    g0838(.A(KEYINPUT108), .ZN(new_n1039));
  NAND3_X1  g0839(.A1(new_n1037), .A2(new_n1038), .A3(new_n1039), .ZN(new_n1040));
  NAND4_X1  g0840(.A1(new_n1035), .A2(new_n704), .A3(new_n1011), .A4(new_n1040), .ZN(new_n1041));
  INV_X1    g0841(.A(new_n754), .ZN(new_n1042));
  INV_X1    g0842(.A(new_n706), .ZN(new_n1043));
  AOI211_X1 g0843(.A(G45), .B(new_n1043), .C1(G68), .C2(G77), .ZN(new_n1044));
  NOR2_X1   g0844(.A1(new_n345), .A2(G50), .ZN(new_n1045));
  XNOR2_X1  g0845(.A(new_n1045), .B(KEYINPUT50), .ZN(new_n1046));
  AOI21_X1  g0846(.A(new_n760), .B1(new_n1044), .B2(new_n1046), .ZN(new_n1047));
  OAI21_X1  g0847(.A(new_n1047), .B1(new_n227), .B2(new_n456), .ZN(new_n1048));
  OAI221_X1 g0848(.A(new_n1048), .B1(G107), .B2(new_n205), .C1(new_n706), .C2(new_n755), .ZN(new_n1049));
  AOI21_X1  g0849(.A(new_n1042), .B1(new_n1049), .B2(new_n770), .ZN(new_n1050));
  AOI21_X1  g0850(.A(new_n505), .B1(new_n775), .B2(G159), .ZN(new_n1051));
  NAND2_X1  g0851(.A1(new_n962), .A2(G77), .ZN(new_n1052));
  NAND3_X1  g0852(.A1(new_n1051), .A2(new_n974), .A3(new_n1052), .ZN(new_n1053));
  OAI22_X1  g0853(.A1(new_n842), .A2(new_n388), .B1(new_n345), .B2(new_n780), .ZN(new_n1054));
  NOR2_X1   g0854(.A1(new_n598), .A2(new_n798), .ZN(new_n1055));
  OAI22_X1  g0855(.A1(new_n778), .A2(new_n212), .B1(new_n786), .B2(new_n383), .ZN(new_n1056));
  NOR4_X1   g0856(.A1(new_n1053), .A2(new_n1054), .A3(new_n1055), .A4(new_n1056), .ZN(new_n1057));
  AOI22_X1  g0857(.A1(new_n781), .A2(G311), .B1(new_n809), .B2(G303), .ZN(new_n1058));
  INV_X1    g0858(.A(G322), .ZN(new_n1059));
  OAI221_X1 g0859(.A(new_n1058), .B1(new_n1059), .B2(new_n776), .C1(new_n794), .C2(new_n970), .ZN(new_n1060));
  INV_X1    g0860(.A(KEYINPUT48), .ZN(new_n1061));
  OR2_X1    g0861(.A1(new_n1060), .A2(new_n1061), .ZN(new_n1062));
  NAND2_X1  g0862(.A1(new_n1060), .A2(new_n1061), .ZN(new_n1063));
  AOI22_X1  g0863(.A1(new_n799), .A2(G283), .B1(new_n962), .B2(G294), .ZN(new_n1064));
  NAND3_X1  g0864(.A1(new_n1062), .A2(new_n1063), .A3(new_n1064), .ZN(new_n1065));
  INV_X1    g0865(.A(KEYINPUT49), .ZN(new_n1066));
  NOR2_X1   g0866(.A1(new_n1065), .A2(new_n1066), .ZN(new_n1067));
  AOI21_X1  g0867(.A(new_n244), .B1(new_n806), .B2(G326), .ZN(new_n1068));
  OAI21_X1  g0868(.A(new_n1068), .B1(new_n520), .B2(new_n790), .ZN(new_n1069));
  NOR2_X1   g0869(.A1(new_n1067), .A2(new_n1069), .ZN(new_n1070));
  NAND2_X1  g0870(.A1(new_n1065), .A2(new_n1066), .ZN(new_n1071));
  AOI21_X1  g0871(.A(new_n1057), .B1(new_n1070), .B2(new_n1071), .ZN(new_n1072));
  OAI221_X1 g0872(.A(new_n1050), .B1(new_n1008), .B2(new_n816), .C1(new_n1072), .C2(new_n765), .ZN(new_n1073));
  OAI21_X1  g0873(.A(new_n1073), .B1(new_n1038), .B2(new_n750), .ZN(new_n1074));
  INV_X1    g0874(.A(new_n1074), .ZN(new_n1075));
  NAND2_X1  g0875(.A1(new_n1041), .A2(new_n1075), .ZN(G393));
  OAI21_X1  g0876(.A(new_n1011), .B1(new_n1004), .B2(new_n1006), .ZN(new_n1077));
  NAND3_X1  g0877(.A1(new_n1013), .A2(new_n704), .A3(new_n1077), .ZN(new_n1078));
  NAND2_X1  g0878(.A1(new_n995), .A2(new_n769), .ZN(new_n1079));
  OAI221_X1 g0879(.A(new_n770), .B1(new_n555), .B2(new_n205), .C1(new_n237), .C2(new_n760), .ZN(new_n1080));
  OAI21_X1  g0880(.A(new_n754), .B1(new_n1080), .B2(KEYINPUT109), .ZN(new_n1081));
  AOI22_X1  g0881(.A1(new_n793), .A2(G159), .B1(new_n775), .B2(G150), .ZN(new_n1082));
  XOR2_X1   g0882(.A(new_n1082), .B(KEYINPUT51), .Z(new_n1083));
  OAI22_X1  g0883(.A1(new_n778), .A2(new_n345), .B1(new_n786), .B2(new_n849), .ZN(new_n1084));
  AOI211_X1 g0884(.A(new_n505), .B(new_n1084), .C1(G50), .C2(new_n781), .ZN(new_n1085));
  NOR2_X1   g0885(.A1(new_n784), .A2(new_n212), .ZN(new_n1086));
  AOI211_X1 g0886(.A(new_n846), .B(new_n1086), .C1(G77), .C2(new_n799), .ZN(new_n1087));
  NAND3_X1  g0887(.A1(new_n1083), .A2(new_n1085), .A3(new_n1087), .ZN(new_n1088));
  AOI22_X1  g0888(.A1(new_n793), .A2(G311), .B1(new_n775), .B2(G317), .ZN(new_n1089));
  XOR2_X1   g0889(.A(new_n1089), .B(KEYINPUT52), .Z(new_n1090));
  OAI22_X1  g0890(.A1(new_n778), .A2(new_n464), .B1(new_n786), .B2(new_n1059), .ZN(new_n1091));
  AOI211_X1 g0891(.A(new_n244), .B(new_n1091), .C1(G303), .C2(new_n781), .ZN(new_n1092));
  OAI22_X1  g0892(.A1(new_n418), .A2(new_n790), .B1(new_n784), .B2(new_n841), .ZN(new_n1093));
  AOI21_X1  g0893(.A(new_n1093), .B1(G116), .B2(new_n799), .ZN(new_n1094));
  NAND3_X1  g0894(.A1(new_n1090), .A2(new_n1092), .A3(new_n1094), .ZN(new_n1095));
  AOI21_X1  g0895(.A(new_n765), .B1(new_n1088), .B2(new_n1095), .ZN(new_n1096));
  AOI211_X1 g0896(.A(new_n1081), .B(new_n1096), .C1(KEYINPUT109), .C2(new_n1080), .ZN(new_n1097));
  AOI22_X1  g0897(.A1(new_n1007), .A2(new_n752), .B1(new_n1079), .B2(new_n1097), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n1078), .A2(new_n1098), .ZN(G390));
  NAND2_X1  g0899(.A1(new_n826), .A2(G330), .ZN(new_n1100));
  OAI21_X1  g0900(.A(new_n928), .B1(new_n913), .B2(new_n1100), .ZN(new_n1101));
  AOI21_X1  g0901(.A(new_n682), .B1(new_n715), .B2(new_n720), .ZN(new_n1102));
  NAND2_X1  g0902(.A1(new_n825), .A2(new_n451), .ZN(new_n1103));
  AOI21_X1  g0903(.A(new_n822), .B1(new_n1102), .B2(new_n1103), .ZN(new_n1104));
  NAND3_X1  g0904(.A1(new_n826), .A2(new_n742), .A3(G330), .ZN(new_n1105));
  NOR2_X1   g0905(.A1(new_n1105), .A2(new_n928), .ZN(new_n1106));
  NOR2_X1   g0906(.A1(new_n1106), .A2(KEYINPUT110), .ZN(new_n1107));
  AND2_X1   g0907(.A1(new_n1106), .A2(KEYINPUT110), .ZN(new_n1108));
  OAI211_X1 g0908(.A(new_n1101), .B(new_n1104), .C1(new_n1107), .C2(new_n1108), .ZN(new_n1109));
  NAND4_X1  g0909(.A1(new_n912), .A2(G330), .A3(new_n826), .A4(new_n929), .ZN(new_n1110));
  INV_X1    g0910(.A(new_n1105), .ZN(new_n1111));
  OAI21_X1  g0911(.A(new_n1110), .B1(new_n929), .B2(new_n1111), .ZN(new_n1112));
  OAI21_X1  g0912(.A(new_n821), .B1(new_n936), .B2(new_n937), .ZN(new_n1113));
  NAND2_X1  g0913(.A1(new_n1113), .A2(KEYINPUT98), .ZN(new_n1114));
  NAND2_X1  g0914(.A1(new_n1114), .A2(new_n938), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n1112), .A2(new_n1115), .ZN(new_n1116));
  NAND2_X1  g0916(.A1(new_n1109), .A2(new_n1116), .ZN(new_n1117));
  NAND4_X1  g0917(.A1(new_n455), .A2(G330), .A3(new_n868), .A4(new_n869), .ZN(new_n1118));
  NAND2_X1  g0918(.A1(new_n1118), .A2(KEYINPUT111), .ZN(new_n1119));
  INV_X1    g0919(.A(KEYINPUT111), .ZN(new_n1120));
  NAND4_X1  g0920(.A1(new_n912), .A2(new_n1120), .A3(G330), .A4(new_n455), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n1119), .A2(new_n1121), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n1122), .A2(new_n944), .ZN(new_n1123));
  INV_X1    g0923(.A(new_n1123), .ZN(new_n1124));
  NAND2_X1  g0924(.A1(new_n1117), .A2(new_n1124), .ZN(new_n1125));
  OR2_X1    g0925(.A1(new_n888), .A2(new_n894), .ZN(new_n1126));
  INV_X1    g0926(.A(new_n921), .ZN(new_n1127));
  OAI211_X1 g0927(.A(new_n1126), .B(new_n1127), .C1(new_n1104), .C2(new_n928), .ZN(new_n1128));
  INV_X1    g0928(.A(new_n1128), .ZN(new_n1129));
  OAI21_X1  g0929(.A(new_n929), .B1(new_n935), .B2(new_n939), .ZN(new_n1130));
  NAND2_X1  g0930(.A1(new_n1130), .A2(new_n1127), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n920), .A2(new_n922), .ZN(new_n1132));
  AOI21_X1  g0932(.A(new_n1129), .B1(new_n1131), .B2(new_n1132), .ZN(new_n1133));
  NOR2_X1   g0933(.A1(new_n1133), .A2(new_n1110), .ZN(new_n1134));
  OR2_X1    g0934(.A1(new_n1108), .A2(new_n1107), .ZN(new_n1135));
  AOI21_X1  g0935(.A(new_n921), .B1(new_n1115), .B2(new_n929), .ZN(new_n1136));
  INV_X1    g0936(.A(new_n1132), .ZN(new_n1137));
  OAI211_X1 g0937(.A(new_n1135), .B(new_n1128), .C1(new_n1136), .C2(new_n1137), .ZN(new_n1138));
  INV_X1    g0938(.A(new_n1138), .ZN(new_n1139));
  OAI21_X1  g0939(.A(new_n1125), .B1(new_n1134), .B2(new_n1139), .ZN(new_n1140));
  AOI21_X1  g0940(.A(new_n1123), .B1(new_n1109), .B2(new_n1116), .ZN(new_n1141));
  OAI211_X1 g0941(.A(new_n1141), .B(new_n1138), .C1(new_n1133), .C2(new_n1110), .ZN(new_n1142));
  NAND3_X1  g0942(.A1(new_n1140), .A2(new_n704), .A3(new_n1142), .ZN(new_n1143));
  AOI22_X1  g0943(.A1(new_n781), .A2(G107), .B1(new_n809), .B2(G97), .ZN(new_n1144));
  OAI221_X1 g0944(.A(new_n1144), .B1(new_n464), .B2(new_n786), .C1(new_n520), .C2(new_n842), .ZN(new_n1145));
  OAI21_X1  g0945(.A(new_n505), .B1(new_n776), .B2(new_n841), .ZN(new_n1146));
  OAI22_X1  g0946(.A1(new_n798), .A2(new_n273), .B1(new_n790), .B2(new_n212), .ZN(new_n1147));
  NOR4_X1   g0947(.A1(new_n1145), .A2(new_n785), .A3(new_n1146), .A4(new_n1147), .ZN(new_n1148));
  XOR2_X1   g0948(.A(new_n1148), .B(KEYINPUT112), .Z(new_n1149));
  AOI22_X1  g0949(.A1(new_n793), .A2(G132), .B1(new_n781), .B2(G137), .ZN(new_n1150));
  AOI22_X1  g0950(.A1(new_n775), .A2(G128), .B1(G125), .B2(new_n806), .ZN(new_n1151));
  NAND2_X1  g0951(.A1(new_n1150), .A2(new_n1151), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n962), .A2(G150), .ZN(new_n1153));
  AOI21_X1  g0953(.A(new_n1152), .B1(KEYINPUT53), .B2(new_n1153), .ZN(new_n1154));
  NOR2_X1   g0954(.A1(new_n790), .A2(new_n388), .ZN(new_n1155));
  XNOR2_X1  g0955(.A(KEYINPUT54), .B(G143), .ZN(new_n1156));
  OAI21_X1  g0956(.A(new_n244), .B1(new_n778), .B2(new_n1156), .ZN(new_n1157));
  AOI211_X1 g0957(.A(new_n1155), .B(new_n1157), .C1(G159), .C2(new_n799), .ZN(new_n1158));
  OAI211_X1 g0958(.A(new_n1154), .B(new_n1158), .C1(KEYINPUT53), .C2(new_n1153), .ZN(new_n1159));
  AOI21_X1  g0959(.A(new_n765), .B1(new_n1149), .B2(new_n1159), .ZN(new_n1160));
  OAI21_X1  g0960(.A(new_n754), .B1(new_n839), .B2(new_n432), .ZN(new_n1161));
  AOI211_X1 g0961(.A(new_n1160), .B(new_n1161), .C1(new_n1132), .C2(new_n767), .ZN(new_n1162));
  NOR2_X1   g0962(.A1(new_n1134), .A2(new_n1139), .ZN(new_n1163));
  AOI21_X1  g0963(.A(new_n1162), .B1(new_n1163), .B2(new_n752), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n1143), .A2(new_n1164), .ZN(G378));
  NAND2_X1  g0965(.A1(new_n390), .A2(new_n871), .ZN(new_n1166));
  XNOR2_X1  g0966(.A(new_n411), .B(new_n1166), .ZN(new_n1167));
  XNOR2_X1  g0967(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1168));
  XOR2_X1   g0968(.A(new_n1167), .B(new_n1168), .Z(new_n1169));
  INV_X1    g0969(.A(new_n1169), .ZN(new_n1170));
  AOI21_X1  g0970(.A(new_n1170), .B1(new_n910), .B2(G330), .ZN(new_n1171));
  NAND3_X1  g0971(.A1(new_n1126), .A2(new_n897), .A3(KEYINPUT40), .ZN(new_n1172));
  NAND3_X1  g0972(.A1(new_n866), .A2(new_n868), .A3(new_n869), .ZN(new_n1173));
  AOI21_X1  g0973(.A(new_n1173), .B1(new_n930), .B2(new_n931), .ZN(new_n1174));
  OAI211_X1 g0974(.A(new_n1172), .B(G330), .C1(new_n1174), .C2(KEYINPUT40), .ZN(new_n1175));
  NOR2_X1   g0975(.A1(new_n1175), .A2(new_n1169), .ZN(new_n1176));
  OAI22_X1  g0976(.A1(new_n941), .A2(new_n942), .B1(new_n1171), .B2(new_n1176), .ZN(new_n1177));
  AOI221_X4 g0977(.A(new_n928), .B1(new_n930), .B2(new_n931), .C1(new_n1114), .C2(new_n938), .ZN(new_n1178));
  OAI21_X1  g0978(.A(KEYINPUT101), .B1(new_n1178), .B2(new_n925), .ZN(new_n1179));
  NAND3_X1  g0979(.A1(new_n926), .A2(new_n940), .A3(new_n927), .ZN(new_n1180));
  NAND3_X1  g0980(.A1(new_n910), .A2(G330), .A3(new_n1170), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n1175), .A2(new_n1169), .ZN(new_n1182));
  NAND4_X1  g0982(.A1(new_n1179), .A2(new_n1180), .A3(new_n1181), .A4(new_n1182), .ZN(new_n1183));
  NAND3_X1  g0983(.A1(new_n1177), .A2(new_n752), .A3(new_n1183), .ZN(new_n1184));
  OAI21_X1  g0984(.A(new_n753), .B1(new_n839), .B2(G50), .ZN(new_n1185));
  INV_X1    g0985(.A(G41), .ZN(new_n1186));
  NAND2_X1  g0986(.A1(new_n505), .A2(new_n1186), .ZN(new_n1187));
  OAI211_X1 g0987(.A(new_n1187), .B(new_n388), .C1(G33), .C2(G41), .ZN(new_n1188));
  OAI22_X1  g0988(.A1(new_n776), .A2(new_n520), .B1(new_n786), .B2(new_n841), .ZN(new_n1189));
  AOI211_X1 g0989(.A(new_n1187), .B(new_n1189), .C1(G107), .C2(new_n793), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n799), .A2(G68), .ZN(new_n1191));
  NAND2_X1  g0991(.A1(new_n791), .A2(G58), .ZN(new_n1192));
  XNOR2_X1  g0992(.A(new_n1192), .B(KEYINPUT113), .ZN(new_n1193));
  NAND4_X1  g0993(.A1(new_n1190), .A2(new_n1191), .A3(new_n1052), .A4(new_n1193), .ZN(new_n1194));
  OAI22_X1  g0994(.A1(new_n598), .A2(new_n778), .B1(new_n555), .B2(new_n780), .ZN(new_n1195));
  XNOR2_X1  g0995(.A(new_n1195), .B(KEYINPUT114), .ZN(new_n1196));
  NOR2_X1   g0996(.A1(new_n1194), .A2(new_n1196), .ZN(new_n1197));
  OAI21_X1  g0997(.A(new_n1188), .B1(new_n1197), .B2(KEYINPUT58), .ZN(new_n1198));
  XOR2_X1   g0998(.A(new_n1198), .B(KEYINPUT115), .Z(new_n1199));
  NAND2_X1  g0999(.A1(new_n1197), .A2(KEYINPUT58), .ZN(new_n1200));
  AOI22_X1  g1000(.A1(new_n775), .A2(G125), .B1(new_n781), .B2(G132), .ZN(new_n1201));
  AOI22_X1  g1001(.A1(new_n793), .A2(G128), .B1(G137), .B2(new_n809), .ZN(new_n1202));
  NAND2_X1  g1002(.A1(new_n1201), .A2(new_n1202), .ZN(new_n1203));
  OAI22_X1  g1003(.A1(new_n798), .A2(new_n383), .B1(new_n784), .B2(new_n1156), .ZN(new_n1204));
  NOR2_X1   g1004(.A1(new_n1203), .A2(new_n1204), .ZN(new_n1205));
  INV_X1    g1005(.A(new_n1205), .ZN(new_n1206));
  NOR2_X1   g1006(.A1(new_n1206), .A2(KEYINPUT59), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n1206), .A2(KEYINPUT59), .ZN(new_n1208));
  NAND2_X1  g1008(.A1(new_n791), .A2(G159), .ZN(new_n1209));
  AOI211_X1 g1009(.A(G33), .B(G41), .C1(new_n806), .C2(G124), .ZN(new_n1210));
  NAND3_X1  g1010(.A1(new_n1208), .A2(new_n1209), .A3(new_n1210), .ZN(new_n1211));
  OAI211_X1 g1011(.A(new_n1199), .B(new_n1200), .C1(new_n1207), .C2(new_n1211), .ZN(new_n1212));
  AOI21_X1  g1012(.A(new_n1185), .B1(new_n1212), .B2(new_n766), .ZN(new_n1213));
  OAI21_X1  g1013(.A(new_n1213), .B1(new_n1170), .B2(new_n768), .ZN(new_n1214));
  NAND2_X1  g1014(.A1(new_n1184), .A2(new_n1214), .ZN(new_n1215));
  INV_X1    g1015(.A(new_n1215), .ZN(new_n1216));
  NAND2_X1  g1016(.A1(new_n1142), .A2(new_n1124), .ZN(new_n1217));
  NAND4_X1  g1017(.A1(new_n1217), .A2(KEYINPUT57), .A3(new_n1183), .A4(new_n1177), .ZN(new_n1218));
  NAND2_X1  g1018(.A1(new_n1218), .A2(new_n704), .ZN(new_n1219));
  AND2_X1   g1019(.A1(new_n1177), .A2(new_n1183), .ZN(new_n1220));
  AOI21_X1  g1020(.A(KEYINPUT57), .B1(new_n1220), .B2(new_n1217), .ZN(new_n1221));
  OAI21_X1  g1021(.A(new_n1216), .B1(new_n1219), .B2(new_n1221), .ZN(G375));
  NOR2_X1   g1022(.A1(new_n1117), .A2(new_n1124), .ZN(new_n1223));
  INV_X1    g1023(.A(new_n1223), .ZN(new_n1224));
  NAND3_X1  g1024(.A1(new_n1224), .A2(new_n1015), .A3(new_n1125), .ZN(new_n1225));
  XNOR2_X1  g1025(.A(new_n1225), .B(KEYINPUT116), .ZN(new_n1226));
  OAI21_X1  g1026(.A(new_n754), .B1(new_n839), .B2(G68), .ZN(new_n1227));
  AOI22_X1  g1027(.A1(new_n793), .A2(G283), .B1(new_n781), .B2(G116), .ZN(new_n1228));
  OAI221_X1 g1028(.A(new_n1228), .B1(new_n464), .B2(new_n776), .C1(new_n803), .C2(new_n786), .ZN(new_n1229));
  NOR2_X1   g1029(.A1(new_n1229), .A2(new_n1055), .ZN(new_n1230));
  AOI211_X1 g1030(.A(new_n244), .B(new_n966), .C1(G107), .C2(new_n809), .ZN(new_n1231));
  OAI211_X1 g1031(.A(new_n1230), .B(new_n1231), .C1(new_n555), .C2(new_n784), .ZN(new_n1232));
  OAI21_X1  g1032(.A(new_n244), .B1(new_n780), .B2(new_n1156), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(new_n806), .A2(G128), .ZN(new_n1234));
  OAI21_X1  g1034(.A(new_n1234), .B1(new_n776), .B2(new_n852), .ZN(new_n1235));
  AOI211_X1 g1035(.A(new_n1233), .B(new_n1235), .C1(G159), .C2(new_n962), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n795), .A2(G137), .ZN(new_n1237));
  OAI22_X1  g1037(.A1(new_n798), .A2(new_n388), .B1(new_n778), .B2(new_n383), .ZN(new_n1238));
  XOR2_X1   g1038(.A(new_n1238), .B(KEYINPUT117), .Z(new_n1239));
  NAND4_X1  g1039(.A1(new_n1236), .A2(new_n1237), .A3(new_n1193), .A4(new_n1239), .ZN(new_n1240));
  NAND2_X1  g1040(.A1(new_n1232), .A2(new_n1240), .ZN(new_n1241));
  AOI21_X1  g1041(.A(new_n1227), .B1(new_n1241), .B2(new_n766), .ZN(new_n1242));
  XOR2_X1   g1042(.A(new_n1242), .B(KEYINPUT118), .Z(new_n1243));
  OAI21_X1  g1043(.A(new_n1243), .B1(new_n929), .B2(new_n768), .ZN(new_n1244));
  INV_X1    g1044(.A(new_n1244), .ZN(new_n1245));
  AOI21_X1  g1045(.A(new_n1245), .B1(new_n1117), .B2(new_n752), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(new_n1226), .A2(new_n1246), .ZN(G381));
  INV_X1    g1047(.A(G387), .ZN(new_n1248));
  INV_X1    g1048(.A(G390), .ZN(new_n1249));
  NAND3_X1  g1049(.A1(new_n1041), .A2(new_n819), .A3(new_n1075), .ZN(new_n1250));
  OR2_X1    g1050(.A1(new_n1250), .A2(G384), .ZN(new_n1251));
  INV_X1    g1051(.A(KEYINPUT119), .ZN(new_n1252));
  OAI211_X1 g1052(.A(new_n1248), .B(new_n1249), .C1(new_n1251), .C2(new_n1252), .ZN(new_n1253));
  AOI21_X1  g1053(.A(new_n1253), .B1(new_n1252), .B2(new_n1251), .ZN(new_n1254));
  INV_X1    g1054(.A(G378), .ZN(new_n1255));
  INV_X1    g1055(.A(G375), .ZN(new_n1256));
  INV_X1    g1056(.A(G381), .ZN(new_n1257));
  NAND4_X1  g1057(.A1(new_n1254), .A2(new_n1255), .A3(new_n1256), .A4(new_n1257), .ZN(G407));
  NAND2_X1  g1058(.A1(new_n681), .A2(G213), .ZN(new_n1259));
  INV_X1    g1059(.A(new_n1259), .ZN(new_n1260));
  NAND3_X1  g1060(.A1(new_n1256), .A2(new_n1255), .A3(new_n1260), .ZN(new_n1261));
  NAND3_X1  g1061(.A1(G407), .A2(G213), .A3(new_n1261), .ZN(G409));
  NAND2_X1  g1062(.A1(new_n1215), .A2(KEYINPUT120), .ZN(new_n1263));
  INV_X1    g1063(.A(KEYINPUT120), .ZN(new_n1264));
  NAND3_X1  g1064(.A1(new_n1184), .A2(new_n1264), .A3(new_n1214), .ZN(new_n1265));
  NAND3_X1  g1065(.A1(new_n1220), .A2(new_n1015), .A3(new_n1217), .ZN(new_n1266));
  NAND3_X1  g1066(.A1(new_n1263), .A2(new_n1265), .A3(new_n1266), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(new_n1267), .A2(new_n1255), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1268), .A2(KEYINPUT121), .ZN(new_n1269));
  OAI211_X1 g1069(.A(G378), .B(new_n1216), .C1(new_n1219), .C2(new_n1221), .ZN(new_n1270));
  INV_X1    g1070(.A(KEYINPUT121), .ZN(new_n1271));
  NAND3_X1  g1071(.A1(new_n1267), .A2(new_n1271), .A3(new_n1255), .ZN(new_n1272));
  NAND3_X1  g1072(.A1(new_n1269), .A2(new_n1270), .A3(new_n1272), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(new_n1273), .A2(new_n1259), .ZN(new_n1274));
  INV_X1    g1074(.A(G384), .ZN(new_n1275));
  NAND3_X1  g1075(.A1(new_n1223), .A2(KEYINPUT60), .A3(new_n1125), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(new_n1276), .A2(new_n704), .ZN(new_n1277));
  AOI21_X1  g1077(.A(new_n1223), .B1(KEYINPUT60), .B2(new_n1125), .ZN(new_n1278));
  NOR2_X1   g1078(.A1(new_n1277), .A2(new_n1278), .ZN(new_n1279));
  INV_X1    g1079(.A(new_n1246), .ZN(new_n1280));
  OAI21_X1  g1080(.A(new_n1275), .B1(new_n1279), .B2(new_n1280), .ZN(new_n1281));
  OAI211_X1 g1081(.A(G384), .B(new_n1246), .C1(new_n1277), .C2(new_n1278), .ZN(new_n1282));
  NAND2_X1  g1082(.A1(new_n1281), .A2(new_n1282), .ZN(new_n1283));
  NAND2_X1  g1083(.A1(new_n1260), .A2(G2897), .ZN(new_n1284));
  XNOR2_X1  g1084(.A(new_n1283), .B(new_n1284), .ZN(new_n1285));
  AOI21_X1  g1085(.A(KEYINPUT61), .B1(new_n1274), .B2(new_n1285), .ZN(new_n1286));
  AND2_X1   g1086(.A1(new_n1281), .A2(new_n1282), .ZN(new_n1287));
  NAND3_X1  g1087(.A1(new_n1273), .A2(new_n1259), .A3(new_n1287), .ZN(new_n1288));
  INV_X1    g1088(.A(KEYINPUT63), .ZN(new_n1289));
  NAND2_X1  g1089(.A1(G387), .A2(new_n1249), .ZN(new_n1290));
  NAND2_X1  g1090(.A1(new_n1290), .A2(KEYINPUT123), .ZN(new_n1291));
  OAI211_X1 g1091(.A(new_n991), .B(G390), .C1(new_n1016), .C2(new_n1033), .ZN(new_n1292));
  NAND2_X1  g1092(.A1(G393), .A2(G396), .ZN(new_n1293));
  NAND2_X1  g1093(.A1(new_n1293), .A2(new_n1250), .ZN(new_n1294));
  AND2_X1   g1094(.A1(new_n1292), .A2(new_n1294), .ZN(new_n1295));
  INV_X1    g1095(.A(KEYINPUT123), .ZN(new_n1296));
  NAND3_X1  g1096(.A1(G387), .A2(new_n1296), .A3(new_n1249), .ZN(new_n1297));
  NAND3_X1  g1097(.A1(new_n1291), .A2(new_n1295), .A3(new_n1297), .ZN(new_n1298));
  NAND3_X1  g1098(.A1(new_n1290), .A2(KEYINPUT122), .A3(new_n1292), .ZN(new_n1299));
  INV_X1    g1099(.A(new_n1294), .ZN(new_n1300));
  INV_X1    g1100(.A(KEYINPUT122), .ZN(new_n1301));
  NAND3_X1  g1101(.A1(new_n1248), .A2(new_n1301), .A3(G390), .ZN(new_n1302));
  NAND3_X1  g1102(.A1(new_n1299), .A2(new_n1300), .A3(new_n1302), .ZN(new_n1303));
  AOI22_X1  g1103(.A1(new_n1288), .A2(new_n1289), .B1(new_n1298), .B2(new_n1303), .ZN(new_n1304));
  NAND4_X1  g1104(.A1(new_n1273), .A2(KEYINPUT63), .A3(new_n1259), .A4(new_n1287), .ZN(new_n1305));
  AND2_X1   g1105(.A1(new_n1305), .A2(KEYINPUT124), .ZN(new_n1306));
  NOR2_X1   g1106(.A1(new_n1305), .A2(KEYINPUT124), .ZN(new_n1307));
  OAI211_X1 g1107(.A(new_n1286), .B(new_n1304), .C1(new_n1306), .C2(new_n1307), .ZN(new_n1308));
  NAND2_X1  g1108(.A1(new_n1288), .A2(KEYINPUT62), .ZN(new_n1309));
  INV_X1    g1109(.A(KEYINPUT61), .ZN(new_n1310));
  INV_X1    g1110(.A(new_n1272), .ZN(new_n1311));
  INV_X1    g1111(.A(new_n1270), .ZN(new_n1312));
  AOI21_X1  g1112(.A(new_n1271), .B1(new_n1267), .B2(new_n1255), .ZN(new_n1313));
  NOR3_X1   g1113(.A1(new_n1311), .A2(new_n1312), .A3(new_n1313), .ZN(new_n1314));
  OAI21_X1  g1114(.A(new_n1285), .B1(new_n1314), .B2(new_n1260), .ZN(new_n1315));
  INV_X1    g1115(.A(KEYINPUT62), .ZN(new_n1316));
  NAND4_X1  g1116(.A1(new_n1273), .A2(new_n1316), .A3(new_n1259), .A4(new_n1287), .ZN(new_n1317));
  NAND4_X1  g1117(.A1(new_n1309), .A2(new_n1310), .A3(new_n1315), .A4(new_n1317), .ZN(new_n1318));
  AOI21_X1  g1118(.A(KEYINPUT125), .B1(new_n1303), .B2(new_n1298), .ZN(new_n1319));
  INV_X1    g1119(.A(new_n1319), .ZN(new_n1320));
  INV_X1    g1120(.A(KEYINPUT126), .ZN(new_n1321));
  NAND3_X1  g1121(.A1(new_n1303), .A2(KEYINPUT125), .A3(new_n1298), .ZN(new_n1322));
  NAND3_X1  g1122(.A1(new_n1320), .A2(new_n1321), .A3(new_n1322), .ZN(new_n1323));
  AND3_X1   g1123(.A1(new_n1303), .A2(KEYINPUT125), .A3(new_n1298), .ZN(new_n1324));
  OAI21_X1  g1124(.A(KEYINPUT126), .B1(new_n1324), .B2(new_n1319), .ZN(new_n1325));
  AND2_X1   g1125(.A1(new_n1323), .A2(new_n1325), .ZN(new_n1326));
  NAND2_X1  g1126(.A1(new_n1318), .A2(new_n1326), .ZN(new_n1327));
  NAND2_X1  g1127(.A1(new_n1308), .A2(new_n1327), .ZN(G405));
  NOR2_X1   g1128(.A1(new_n1324), .A2(new_n1319), .ZN(new_n1329));
  NAND2_X1  g1129(.A1(G375), .A2(new_n1255), .ZN(new_n1330));
  NAND3_X1  g1130(.A1(new_n1330), .A2(new_n1283), .A3(new_n1270), .ZN(new_n1331));
  NAND2_X1  g1131(.A1(new_n1330), .A2(new_n1270), .ZN(new_n1332));
  NAND2_X1  g1132(.A1(new_n1332), .A2(new_n1287), .ZN(new_n1333));
  NAND3_X1  g1133(.A1(new_n1329), .A2(new_n1331), .A3(new_n1333), .ZN(new_n1334));
  AOI21_X1  g1134(.A(new_n1329), .B1(new_n1333), .B2(new_n1331), .ZN(new_n1335));
  INV_X1    g1135(.A(KEYINPUT127), .ZN(new_n1336));
  OAI21_X1  g1136(.A(new_n1334), .B1(new_n1335), .B2(new_n1336), .ZN(new_n1337));
  AOI211_X1 g1137(.A(KEYINPUT127), .B(new_n1329), .C1(new_n1333), .C2(new_n1331), .ZN(new_n1338));
  NOR2_X1   g1138(.A1(new_n1337), .A2(new_n1338), .ZN(G402));
endmodule


