//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 0 1 1 1 1 1 1 0 1 1 0 0 0 0 0 0 0 1 1 1 0 0 1 0 1 1 0 1 1 0 0 0 1 0 1 0 1 0 1 1 0 0 0 1 0 0 1 0 1 0 1 0 1 1 0 1 0 0 0 0 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:25:43 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n603, new_n604, new_n605, new_n606, new_n607, new_n608,
    new_n609, new_n610, new_n611, new_n612, new_n614, new_n615, new_n616,
    new_n617, new_n618, new_n619, new_n620, new_n621, new_n622, new_n624,
    new_n625, new_n626, new_n627, new_n628, new_n629, new_n630, new_n631,
    new_n632, new_n633, new_n634, new_n635, new_n636, new_n637, new_n638,
    new_n639, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n687, new_n688, new_n690, new_n691, new_n692,
    new_n693, new_n695, new_n696, new_n697, new_n698, new_n699, new_n700,
    new_n701, new_n702, new_n703, new_n704, new_n705, new_n706, new_n707,
    new_n708, new_n709, new_n710, new_n711, new_n712, new_n713, new_n714,
    new_n715, new_n716, new_n718, new_n719, new_n720, new_n721, new_n722,
    new_n723, new_n724, new_n725, new_n726, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n756, new_n757, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n785, new_n786, new_n787, new_n788, new_n789,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n911, new_n912, new_n913, new_n914, new_n915, new_n916, new_n917,
    new_n918, new_n919, new_n920, new_n921, new_n922, new_n923, new_n924,
    new_n925, new_n926, new_n927, new_n928, new_n929, new_n930, new_n931,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n947, new_n948,
    new_n949, new_n950, new_n951, new_n952, new_n954, new_n955, new_n956,
    new_n957, new_n958, new_n959, new_n960, new_n961, new_n962, new_n963,
    new_n964, new_n965, new_n966, new_n967, new_n968, new_n969, new_n970,
    new_n971, new_n973, new_n974, new_n975, new_n976, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013;
  INV_X1    g000(.A(G221), .ZN(new_n187));
  XNOR2_X1  g001(.A(KEYINPUT9), .B(G234), .ZN(new_n188));
  XOR2_X1   g002(.A(new_n188), .B(KEYINPUT73), .Z(new_n189));
  INV_X1    g003(.A(new_n189), .ZN(new_n190));
  INV_X1    g004(.A(G902), .ZN(new_n191));
  AOI21_X1  g005(.A(new_n187), .B1(new_n190), .B2(new_n191), .ZN(new_n192));
  XNOR2_X1  g006(.A(G110), .B(G140), .ZN(new_n193));
  INV_X1    g007(.A(G227), .ZN(new_n194));
  NOR2_X1   g008(.A1(new_n194), .A2(G953), .ZN(new_n195));
  XNOR2_X1  g009(.A(new_n193), .B(new_n195), .ZN(new_n196));
  INV_X1    g010(.A(new_n196), .ZN(new_n197));
  INV_X1    g011(.A(G128), .ZN(new_n198));
  NOR2_X1   g012(.A1(new_n198), .A2(KEYINPUT1), .ZN(new_n199));
  INV_X1    g013(.A(G146), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n200), .A2(G143), .ZN(new_n201));
  INV_X1    g015(.A(G143), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n202), .A2(G146), .ZN(new_n203));
  NAND3_X1  g017(.A1(new_n199), .A2(new_n201), .A3(new_n203), .ZN(new_n204));
  INV_X1    g018(.A(KEYINPUT65), .ZN(new_n205));
  NOR2_X1   g019(.A1(new_n202), .A2(G146), .ZN(new_n206));
  NOR2_X1   g020(.A1(new_n200), .A2(G143), .ZN(new_n207));
  OAI21_X1  g021(.A(new_n198), .B1(new_n206), .B2(new_n207), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n207), .A2(KEYINPUT1), .ZN(new_n209));
  AOI21_X1  g023(.A(new_n205), .B1(new_n208), .B2(new_n209), .ZN(new_n210));
  AOI21_X1  g024(.A(G128), .B1(new_n201), .B2(new_n203), .ZN(new_n211));
  AND3_X1   g025(.A1(new_n202), .A2(KEYINPUT1), .A3(G146), .ZN(new_n212));
  NOR3_X1   g026(.A1(new_n211), .A2(KEYINPUT65), .A3(new_n212), .ZN(new_n213));
  OAI21_X1  g027(.A(new_n204), .B1(new_n210), .B2(new_n213), .ZN(new_n214));
  INV_X1    g028(.A(KEYINPUT10), .ZN(new_n215));
  INV_X1    g029(.A(G101), .ZN(new_n216));
  INV_X1    g030(.A(G107), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n217), .A2(G104), .ZN(new_n218));
  INV_X1    g032(.A(G104), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n219), .A2(G107), .ZN(new_n220));
  AOI21_X1  g034(.A(new_n216), .B1(new_n218), .B2(new_n220), .ZN(new_n221));
  NAND3_X1  g035(.A1(new_n217), .A2(KEYINPUT74), .A3(G104), .ZN(new_n222));
  INV_X1    g036(.A(KEYINPUT3), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  NAND4_X1  g038(.A1(new_n217), .A2(KEYINPUT74), .A3(KEYINPUT3), .A4(G104), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  NOR2_X1   g040(.A1(new_n217), .A2(G104), .ZN(new_n227));
  AND2_X1   g041(.A1(KEYINPUT75), .A2(G101), .ZN(new_n228));
  NOR2_X1   g042(.A1(KEYINPUT75), .A2(G101), .ZN(new_n229));
  NOR3_X1   g043(.A1(new_n227), .A2(new_n228), .A3(new_n229), .ZN(new_n230));
  AOI211_X1 g044(.A(new_n215), .B(new_n221), .C1(new_n226), .C2(new_n230), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n226), .A2(new_n230), .ZN(new_n232));
  NAND3_X1  g046(.A1(new_n208), .A2(new_n204), .A3(new_n209), .ZN(new_n233));
  INV_X1    g047(.A(new_n221), .ZN(new_n234));
  NAND3_X1  g048(.A1(new_n232), .A2(new_n233), .A3(new_n234), .ZN(new_n235));
  AOI22_X1  g049(.A1(new_n214), .A2(new_n231), .B1(new_n235), .B2(new_n215), .ZN(new_n236));
  AOI21_X1  g050(.A(new_n227), .B1(new_n224), .B2(new_n225), .ZN(new_n237));
  OAI211_X1 g051(.A(new_n232), .B(KEYINPUT4), .C1(new_n216), .C2(new_n237), .ZN(new_n238));
  XNOR2_X1  g052(.A(G143), .B(G146), .ZN(new_n239));
  INV_X1    g053(.A(KEYINPUT0), .ZN(new_n240));
  OAI21_X1  g054(.A(new_n239), .B1(new_n240), .B2(new_n198), .ZN(new_n241));
  XOR2_X1   g055(.A(KEYINPUT0), .B(G128), .Z(new_n242));
  OAI21_X1  g056(.A(new_n241), .B1(new_n239), .B2(new_n242), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n226), .A2(new_n220), .ZN(new_n244));
  INV_X1    g058(.A(KEYINPUT4), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n245), .A2(G101), .ZN(new_n246));
  INV_X1    g060(.A(new_n246), .ZN(new_n247));
  AOI21_X1  g061(.A(KEYINPUT76), .B1(new_n244), .B2(new_n247), .ZN(new_n248));
  INV_X1    g062(.A(KEYINPUT76), .ZN(new_n249));
  NOR3_X1   g063(.A1(new_n237), .A2(new_n249), .A3(new_n246), .ZN(new_n250));
  OAI211_X1 g064(.A(new_n238), .B(new_n243), .C1(new_n248), .C2(new_n250), .ZN(new_n251));
  INV_X1    g065(.A(KEYINPUT11), .ZN(new_n252));
  INV_X1    g066(.A(G134), .ZN(new_n253));
  OAI21_X1  g067(.A(new_n252), .B1(new_n253), .B2(G137), .ZN(new_n254));
  INV_X1    g068(.A(G137), .ZN(new_n255));
  NAND3_X1  g069(.A1(new_n255), .A2(KEYINPUT11), .A3(G134), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n253), .A2(G137), .ZN(new_n257));
  NAND3_X1  g071(.A1(new_n254), .A2(new_n256), .A3(new_n257), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n258), .A2(G131), .ZN(new_n259));
  INV_X1    g073(.A(G131), .ZN(new_n260));
  NAND4_X1  g074(.A1(new_n254), .A2(new_n256), .A3(new_n260), .A4(new_n257), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n259), .A2(new_n261), .ZN(new_n262));
  INV_X1    g076(.A(new_n262), .ZN(new_n263));
  NAND3_X1  g077(.A1(new_n236), .A2(new_n251), .A3(new_n263), .ZN(new_n264));
  INV_X1    g078(.A(KEYINPUT77), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  NAND4_X1  g080(.A1(new_n236), .A2(new_n251), .A3(KEYINPUT77), .A4(new_n263), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n236), .A2(new_n251), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n269), .A2(new_n262), .ZN(new_n270));
  AOI21_X1  g084(.A(new_n197), .B1(new_n268), .B2(new_n270), .ZN(new_n271));
  INV_X1    g085(.A(new_n271), .ZN(new_n272));
  NAND3_X1  g086(.A1(new_n268), .A2(KEYINPUT78), .A3(new_n197), .ZN(new_n273));
  AOI21_X1  g087(.A(new_n221), .B1(new_n226), .B2(new_n230), .ZN(new_n274));
  OAI21_X1  g088(.A(new_n235), .B1(new_n214), .B2(new_n274), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n275), .A2(new_n262), .ZN(new_n276));
  INV_X1    g090(.A(KEYINPUT12), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  NAND3_X1  g092(.A1(new_n275), .A2(KEYINPUT12), .A3(new_n262), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n273), .A2(new_n280), .ZN(new_n281));
  AOI21_X1  g095(.A(new_n196), .B1(new_n266), .B2(new_n267), .ZN(new_n282));
  NOR2_X1   g096(.A1(new_n282), .A2(KEYINPUT78), .ZN(new_n283));
  OAI21_X1  g097(.A(new_n272), .B1(new_n281), .B2(new_n283), .ZN(new_n284));
  INV_X1    g098(.A(G469), .ZN(new_n285));
  NAND3_X1  g099(.A1(new_n284), .A2(new_n285), .A3(new_n191), .ZN(new_n286));
  INV_X1    g100(.A(KEYINPUT79), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n268), .A2(new_n197), .ZN(new_n289));
  INV_X1    g103(.A(KEYINPUT78), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  AND2_X1   g105(.A1(new_n278), .A2(new_n279), .ZN(new_n292));
  AOI21_X1  g106(.A(new_n292), .B1(new_n282), .B2(KEYINPUT78), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n291), .A2(new_n293), .ZN(new_n294));
  AOI21_X1  g108(.A(G902), .B1(new_n294), .B2(new_n272), .ZN(new_n295));
  NAND3_X1  g109(.A1(new_n295), .A2(KEYINPUT79), .A3(new_n285), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n288), .A2(new_n296), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n268), .A2(new_n280), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n298), .A2(new_n196), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n282), .A2(new_n270), .ZN(new_n300));
  AND2_X1   g114(.A1(new_n299), .A2(new_n300), .ZN(new_n301));
  OAI21_X1  g115(.A(G469), .B1(new_n301), .B2(G902), .ZN(new_n302));
  AOI21_X1  g116(.A(new_n192), .B1(new_n297), .B2(new_n302), .ZN(new_n303));
  INV_X1    g117(.A(KEYINPUT28), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n262), .A2(new_n243), .ZN(new_n305));
  OAI21_X1  g119(.A(KEYINPUT65), .B1(new_n211), .B2(new_n212), .ZN(new_n306));
  OAI211_X1 g120(.A(new_n209), .B(new_n205), .C1(new_n239), .C2(G128), .ZN(new_n307));
  AOI22_X1  g121(.A1(new_n306), .A2(new_n307), .B1(new_n239), .B2(new_n199), .ZN(new_n308));
  INV_X1    g122(.A(new_n257), .ZN(new_n309));
  NOR2_X1   g123(.A1(new_n253), .A2(G137), .ZN(new_n310));
  OAI21_X1  g124(.A(G131), .B1(new_n309), .B2(new_n310), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n311), .A2(new_n261), .ZN(new_n312));
  OAI21_X1  g126(.A(new_n305), .B1(new_n308), .B2(new_n312), .ZN(new_n313));
  XOR2_X1   g127(.A(KEYINPUT2), .B(G113), .Z(new_n314));
  XNOR2_X1  g128(.A(G116), .B(G119), .ZN(new_n315));
  XNOR2_X1  g129(.A(new_n314), .B(new_n315), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n313), .A2(new_n316), .ZN(new_n317));
  INV_X1    g131(.A(new_n316), .ZN(new_n318));
  OAI211_X1 g132(.A(new_n318), .B(new_n305), .C1(new_n308), .C2(new_n312), .ZN(new_n319));
  AOI21_X1  g133(.A(new_n304), .B1(new_n317), .B2(new_n319), .ZN(new_n320));
  OR2_X1    g134(.A1(new_n320), .A2(KEYINPUT67), .ZN(new_n321));
  INV_X1    g135(.A(new_n319), .ZN(new_n322));
  NOR2_X1   g136(.A1(new_n322), .A2(KEYINPUT28), .ZN(new_n323));
  OAI21_X1  g137(.A(KEYINPUT67), .B1(new_n320), .B2(new_n323), .ZN(new_n324));
  NOR2_X1   g138(.A1(G237), .A2(G953), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n325), .A2(G210), .ZN(new_n326));
  XNOR2_X1  g140(.A(new_n326), .B(KEYINPUT27), .ZN(new_n327));
  XNOR2_X1  g141(.A(KEYINPUT26), .B(G101), .ZN(new_n328));
  XNOR2_X1  g142(.A(new_n327), .B(new_n328), .ZN(new_n329));
  NAND4_X1  g143(.A1(new_n321), .A2(new_n324), .A3(KEYINPUT29), .A4(new_n329), .ZN(new_n330));
  INV_X1    g144(.A(new_n329), .ZN(new_n331));
  NOR3_X1   g145(.A1(new_n320), .A2(new_n323), .A3(new_n331), .ZN(new_n332));
  OR2_X1    g146(.A1(new_n332), .A2(KEYINPUT29), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n313), .A2(KEYINPUT64), .ZN(new_n334));
  INV_X1    g148(.A(KEYINPUT30), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  NAND3_X1  g150(.A1(new_n313), .A2(KEYINPUT64), .A3(KEYINPUT30), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n336), .A2(new_n337), .ZN(new_n338));
  AOI21_X1  g152(.A(new_n322), .B1(new_n338), .B2(new_n316), .ZN(new_n339));
  NOR2_X1   g153(.A1(new_n339), .A2(new_n329), .ZN(new_n340));
  OAI211_X1 g154(.A(new_n330), .B(new_n191), .C1(new_n333), .C2(new_n340), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n341), .A2(G472), .ZN(new_n342));
  AND3_X1   g156(.A1(new_n313), .A2(KEYINPUT64), .A3(KEYINPUT30), .ZN(new_n343));
  AOI21_X1  g157(.A(KEYINPUT30), .B1(new_n313), .B2(KEYINPUT64), .ZN(new_n344));
  OAI21_X1  g158(.A(new_n316), .B1(new_n343), .B2(new_n344), .ZN(new_n345));
  NAND3_X1  g159(.A1(new_n345), .A2(new_n319), .A3(new_n329), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n346), .A2(KEYINPUT31), .ZN(new_n347));
  OAI21_X1  g161(.A(new_n331), .B1(new_n320), .B2(new_n323), .ZN(new_n348));
  INV_X1    g162(.A(KEYINPUT31), .ZN(new_n349));
  NAND4_X1  g163(.A1(new_n345), .A2(new_n349), .A3(new_n319), .A4(new_n329), .ZN(new_n350));
  NAND3_X1  g164(.A1(new_n347), .A2(new_n348), .A3(new_n350), .ZN(new_n351));
  INV_X1    g165(.A(KEYINPUT32), .ZN(new_n352));
  INV_X1    g166(.A(G472), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n353), .A2(new_n191), .ZN(new_n354));
  XNOR2_X1  g168(.A(new_n354), .B(KEYINPUT66), .ZN(new_n355));
  AND3_X1   g169(.A1(new_n351), .A2(new_n352), .A3(new_n355), .ZN(new_n356));
  AOI21_X1  g170(.A(new_n352), .B1(new_n351), .B2(new_n355), .ZN(new_n357));
  OAI21_X1  g171(.A(new_n342), .B1(new_n356), .B2(new_n357), .ZN(new_n358));
  INV_X1    g172(.A(G217), .ZN(new_n359));
  AOI21_X1  g173(.A(new_n359), .B1(G234), .B2(new_n191), .ZN(new_n360));
  INV_X1    g174(.A(new_n360), .ZN(new_n361));
  INV_X1    g175(.A(G140), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n362), .A2(G125), .ZN(new_n363));
  OAI21_X1  g177(.A(KEYINPUT71), .B1(new_n363), .B2(KEYINPUT16), .ZN(new_n364));
  INV_X1    g178(.A(KEYINPUT71), .ZN(new_n365));
  INV_X1    g179(.A(KEYINPUT16), .ZN(new_n366));
  NAND4_X1  g180(.A1(new_n365), .A2(new_n366), .A3(new_n362), .A4(G125), .ZN(new_n367));
  AND2_X1   g181(.A1(new_n364), .A2(new_n367), .ZN(new_n368));
  INV_X1    g182(.A(G125), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n369), .A2(G140), .ZN(new_n370));
  NAND3_X1  g184(.A1(new_n370), .A2(new_n363), .A3(KEYINPUT70), .ZN(new_n371));
  OR3_X1    g185(.A1(new_n362), .A2(KEYINPUT70), .A3(G125), .ZN(new_n372));
  AOI21_X1  g186(.A(new_n366), .B1(new_n371), .B2(new_n372), .ZN(new_n373));
  OAI21_X1  g187(.A(new_n200), .B1(new_n368), .B2(new_n373), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n364), .A2(new_n367), .ZN(new_n375));
  NOR3_X1   g189(.A1(new_n362), .A2(KEYINPUT70), .A3(G125), .ZN(new_n376));
  XNOR2_X1  g190(.A(G125), .B(G140), .ZN(new_n377));
  AOI21_X1  g191(.A(new_n376), .B1(new_n377), .B2(KEYINPUT70), .ZN(new_n378));
  OAI211_X1 g192(.A(G146), .B(new_n375), .C1(new_n378), .C2(new_n366), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n374), .A2(new_n379), .ZN(new_n380));
  INV_X1    g194(.A(G110), .ZN(new_n381));
  OAI211_X1 g195(.A(KEYINPUT69), .B(KEYINPUT23), .C1(new_n198), .C2(G119), .ZN(new_n382));
  INV_X1    g196(.A(G119), .ZN(new_n383));
  NOR2_X1   g197(.A1(new_n383), .A2(G128), .ZN(new_n384));
  OAI211_X1 g198(.A(new_n382), .B(new_n384), .C1(KEYINPUT69), .C2(KEYINPUT23), .ZN(new_n385));
  OAI21_X1  g199(.A(new_n385), .B1(new_n384), .B2(new_n382), .ZN(new_n386));
  INV_X1    g200(.A(KEYINPUT68), .ZN(new_n387));
  AOI21_X1  g201(.A(new_n387), .B1(new_n383), .B2(G128), .ZN(new_n388));
  NOR3_X1   g202(.A1(new_n198), .A2(KEYINPUT68), .A3(G119), .ZN(new_n389));
  OAI22_X1  g203(.A1(new_n388), .A2(new_n389), .B1(new_n383), .B2(G128), .ZN(new_n390));
  XNOR2_X1  g204(.A(KEYINPUT24), .B(G110), .ZN(new_n391));
  OAI221_X1 g205(.A(new_n380), .B1(new_n381), .B2(new_n386), .C1(new_n390), .C2(new_n391), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n386), .A2(new_n381), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n390), .A2(new_n391), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n393), .A2(new_n394), .ZN(new_n395));
  INV_X1    g209(.A(KEYINPUT72), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n379), .A2(new_n396), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n371), .A2(new_n372), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n398), .A2(KEYINPUT16), .ZN(new_n399));
  NAND4_X1  g213(.A1(new_n399), .A2(KEYINPUT72), .A3(G146), .A4(new_n375), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n377), .A2(new_n200), .ZN(new_n401));
  NAND4_X1  g215(.A1(new_n395), .A2(new_n397), .A3(new_n400), .A4(new_n401), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n392), .A2(new_n402), .ZN(new_n403));
  XNOR2_X1  g217(.A(KEYINPUT22), .B(G137), .ZN(new_n404));
  INV_X1    g218(.A(G234), .ZN(new_n405));
  NOR3_X1   g219(.A1(new_n187), .A2(new_n405), .A3(G953), .ZN(new_n406));
  XOR2_X1   g220(.A(new_n404), .B(new_n406), .Z(new_n407));
  INV_X1    g221(.A(new_n407), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n403), .A2(new_n408), .ZN(new_n409));
  NAND3_X1  g223(.A1(new_n392), .A2(new_n402), .A3(new_n407), .ZN(new_n410));
  NAND3_X1  g224(.A1(new_n409), .A2(new_n191), .A3(new_n410), .ZN(new_n411));
  INV_X1    g225(.A(KEYINPUT25), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n411), .A2(new_n412), .ZN(new_n413));
  NAND4_X1  g227(.A1(new_n409), .A2(KEYINPUT25), .A3(new_n191), .A4(new_n410), .ZN(new_n414));
  AOI21_X1  g228(.A(new_n361), .B1(new_n413), .B2(new_n414), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n409), .A2(new_n410), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n361), .A2(new_n191), .ZN(new_n417));
  NOR2_X1   g231(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  NOR2_X1   g232(.A1(new_n415), .A2(new_n418), .ZN(new_n419));
  XNOR2_X1  g233(.A(G110), .B(G122), .ZN(new_n420));
  OAI211_X1 g234(.A(new_n238), .B(new_n316), .C1(new_n248), .C2(new_n250), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n314), .A2(new_n315), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n315), .A2(KEYINPUT5), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n383), .A2(G116), .ZN(new_n424));
  OR2_X1    g238(.A1(new_n424), .A2(KEYINPUT5), .ZN(new_n425));
  NAND3_X1  g239(.A1(new_n423), .A2(G113), .A3(new_n425), .ZN(new_n426));
  AND3_X1   g240(.A1(new_n274), .A2(new_n422), .A3(new_n426), .ZN(new_n427));
  INV_X1    g241(.A(new_n427), .ZN(new_n428));
  AOI21_X1  g242(.A(new_n420), .B1(new_n421), .B2(new_n428), .ZN(new_n429));
  INV_X1    g243(.A(new_n429), .ZN(new_n430));
  NAND3_X1  g244(.A1(new_n421), .A2(new_n420), .A3(new_n428), .ZN(new_n431));
  NAND3_X1  g245(.A1(new_n430), .A2(KEYINPUT6), .A3(new_n431), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n243), .A2(G125), .ZN(new_n433));
  OAI21_X1  g247(.A(new_n433), .B1(new_n308), .B2(G125), .ZN(new_n434));
  XNOR2_X1  g248(.A(KEYINPUT81), .B(G224), .ZN(new_n435));
  NOR2_X1   g249(.A1(new_n435), .A2(G953), .ZN(new_n436));
  OR2_X1    g250(.A1(new_n434), .A2(new_n436), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n434), .A2(new_n436), .ZN(new_n438));
  AND2_X1   g252(.A1(new_n437), .A2(new_n438), .ZN(new_n439));
  INV_X1    g253(.A(KEYINPUT6), .ZN(new_n440));
  AND3_X1   g254(.A1(new_n429), .A2(KEYINPUT80), .A3(new_n440), .ZN(new_n441));
  AOI21_X1  g255(.A(KEYINPUT80), .B1(new_n429), .B2(new_n440), .ZN(new_n442));
  OAI211_X1 g256(.A(new_n432), .B(new_n439), .C1(new_n441), .C2(new_n442), .ZN(new_n443));
  XNOR2_X1  g257(.A(new_n420), .B(KEYINPUT8), .ZN(new_n444));
  AOI21_X1  g258(.A(new_n274), .B1(new_n422), .B2(new_n426), .ZN(new_n445));
  OAI21_X1  g259(.A(new_n444), .B1(new_n427), .B2(new_n445), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n431), .A2(new_n446), .ZN(new_n447));
  NOR3_X1   g261(.A1(new_n434), .A2(KEYINPUT7), .A3(new_n436), .ZN(new_n448));
  NOR2_X1   g262(.A1(new_n447), .A2(new_n448), .ZN(new_n449));
  OAI211_X1 g263(.A(new_n437), .B(new_n438), .C1(KEYINPUT7), .C2(new_n436), .ZN(new_n450));
  AOI21_X1  g264(.A(G902), .B1(new_n449), .B2(new_n450), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n443), .A2(new_n451), .ZN(new_n452));
  OAI21_X1  g266(.A(G210), .B1(G237), .B2(G902), .ZN(new_n453));
  NOR2_X1   g267(.A1(new_n453), .A2(KEYINPUT82), .ZN(new_n454));
  OR2_X1    g268(.A1(new_n452), .A2(new_n454), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n452), .A2(new_n454), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n455), .A2(new_n456), .ZN(new_n457));
  INV_X1    g271(.A(G953), .ZN(new_n458));
  AND2_X1   g272(.A1(new_n458), .A2(G952), .ZN(new_n459));
  INV_X1    g273(.A(G237), .ZN(new_n460));
  OAI21_X1  g274(.A(new_n459), .B1(new_n405), .B2(new_n460), .ZN(new_n461));
  INV_X1    g275(.A(new_n461), .ZN(new_n462));
  INV_X1    g276(.A(G898), .ZN(new_n463));
  AOI21_X1  g277(.A(new_n458), .B1(KEYINPUT21), .B2(new_n463), .ZN(new_n464));
  OAI21_X1  g278(.A(new_n464), .B1(KEYINPUT21), .B2(new_n463), .ZN(new_n465));
  INV_X1    g279(.A(new_n465), .ZN(new_n466));
  AOI21_X1  g280(.A(new_n191), .B1(G234), .B2(G237), .ZN(new_n467));
  AOI21_X1  g281(.A(new_n462), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  INV_X1    g282(.A(new_n468), .ZN(new_n469));
  OAI21_X1  g283(.A(G214), .B1(G237), .B2(G902), .ZN(new_n470));
  NAND3_X1  g284(.A1(new_n457), .A2(new_n469), .A3(new_n470), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n202), .A2(G128), .ZN(new_n472));
  INV_X1    g286(.A(KEYINPUT13), .ZN(new_n473));
  OAI21_X1  g287(.A(KEYINPUT89), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  INV_X1    g288(.A(KEYINPUT89), .ZN(new_n475));
  NAND4_X1  g289(.A1(new_n475), .A2(new_n202), .A3(KEYINPUT13), .A4(G128), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n198), .A2(G143), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n472), .A2(new_n473), .ZN(new_n478));
  NAND4_X1  g292(.A1(new_n474), .A2(new_n476), .A3(new_n477), .A4(new_n478), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n479), .A2(G134), .ZN(new_n480));
  AND2_X1   g294(.A1(new_n472), .A2(new_n477), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n481), .A2(new_n253), .ZN(new_n482));
  XNOR2_X1  g296(.A(G116), .B(G122), .ZN(new_n483));
  INV_X1    g297(.A(new_n483), .ZN(new_n484));
  NOR2_X1   g298(.A1(new_n484), .A2(G107), .ZN(new_n485));
  NOR2_X1   g299(.A1(new_n483), .A2(new_n217), .ZN(new_n486));
  OAI211_X1 g300(.A(new_n480), .B(new_n482), .C1(new_n485), .C2(new_n486), .ZN(new_n487));
  XNOR2_X1  g301(.A(new_n481), .B(new_n253), .ZN(new_n488));
  INV_X1    g302(.A(new_n485), .ZN(new_n489));
  INV_X1    g303(.A(G116), .ZN(new_n490));
  NAND3_X1  g304(.A1(new_n490), .A2(KEYINPUT14), .A3(G122), .ZN(new_n491));
  OAI211_X1 g305(.A(G107), .B(new_n491), .C1(new_n484), .C2(KEYINPUT14), .ZN(new_n492));
  NAND3_X1  g306(.A1(new_n488), .A2(new_n489), .A3(new_n492), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n487), .A2(new_n493), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n494), .A2(KEYINPUT90), .ZN(new_n495));
  INV_X1    g309(.A(KEYINPUT90), .ZN(new_n496));
  NAND3_X1  g310(.A1(new_n487), .A2(new_n493), .A3(new_n496), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n495), .A2(new_n497), .ZN(new_n498));
  NOR3_X1   g312(.A1(new_n189), .A2(new_n359), .A3(G953), .ZN(new_n499));
  INV_X1    g313(.A(new_n499), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n498), .A2(new_n500), .ZN(new_n501));
  NAND3_X1  g315(.A1(new_n495), .A2(new_n499), .A3(new_n497), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n503), .A2(new_n191), .ZN(new_n504));
  INV_X1    g318(.A(G478), .ZN(new_n505));
  NOR2_X1   g319(.A1(new_n505), .A2(KEYINPUT15), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n504), .A2(new_n506), .ZN(new_n507));
  OAI211_X1 g321(.A(new_n503), .B(new_n191), .C1(KEYINPUT15), .C2(new_n505), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  NAND3_X1  g323(.A1(new_n325), .A2(G143), .A3(G214), .ZN(new_n510));
  INV_X1    g324(.A(new_n510), .ZN(new_n511));
  AOI21_X1  g325(.A(G143), .B1(new_n325), .B2(G214), .ZN(new_n512));
  OAI21_X1  g326(.A(G131), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  INV_X1    g327(.A(new_n512), .ZN(new_n514));
  NAND3_X1  g328(.A1(new_n514), .A2(new_n260), .A3(new_n510), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n513), .A2(new_n515), .ZN(new_n516));
  INV_X1    g330(.A(KEYINPUT84), .ZN(new_n517));
  NOR2_X1   g331(.A1(new_n517), .A2(KEYINPUT19), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n377), .A2(new_n518), .ZN(new_n519));
  AOI22_X1  g333(.A1(new_n371), .A2(new_n372), .B1(new_n377), .B2(new_n517), .ZN(new_n520));
  INV_X1    g334(.A(KEYINPUT19), .ZN(new_n521));
  OAI211_X1 g335(.A(new_n200), .B(new_n519), .C1(new_n520), .C2(new_n521), .ZN(new_n522));
  NAND4_X1  g336(.A1(new_n397), .A2(new_n400), .A3(new_n516), .A4(new_n522), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n514), .A2(new_n510), .ZN(new_n524));
  NAND3_X1  g338(.A1(new_n524), .A2(KEYINPUT18), .A3(G131), .ZN(new_n525));
  OAI21_X1  g339(.A(new_n401), .B1(new_n398), .B2(new_n200), .ZN(new_n526));
  NAND2_X1  g340(.A1(KEYINPUT18), .A2(G131), .ZN(new_n527));
  NAND3_X1  g341(.A1(new_n514), .A2(new_n510), .A3(new_n527), .ZN(new_n528));
  NAND3_X1  g342(.A1(new_n525), .A2(new_n526), .A3(new_n528), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n523), .A2(new_n529), .ZN(new_n530));
  XOR2_X1   g344(.A(G113), .B(G122), .Z(new_n531));
  XOR2_X1   g345(.A(KEYINPUT85), .B(G104), .Z(new_n532));
  XOR2_X1   g346(.A(new_n531), .B(new_n532), .Z(new_n533));
  INV_X1    g347(.A(new_n533), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n530), .A2(new_n534), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n535), .A2(KEYINPUT86), .ZN(new_n536));
  INV_X1    g350(.A(KEYINPUT87), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n380), .A2(new_n537), .ZN(new_n538));
  NAND3_X1  g352(.A1(new_n374), .A2(KEYINPUT87), .A3(new_n379), .ZN(new_n539));
  INV_X1    g353(.A(KEYINPUT17), .ZN(new_n540));
  NOR2_X1   g354(.A1(new_n513), .A2(new_n540), .ZN(new_n541));
  AND2_X1   g355(.A1(new_n513), .A2(new_n515), .ZN(new_n542));
  AOI21_X1  g356(.A(new_n541), .B1(new_n542), .B2(new_n540), .ZN(new_n543));
  NAND3_X1  g357(.A1(new_n538), .A2(new_n539), .A3(new_n543), .ZN(new_n544));
  NAND3_X1  g358(.A1(new_n544), .A2(new_n533), .A3(new_n529), .ZN(new_n545));
  INV_X1    g359(.A(KEYINPUT86), .ZN(new_n546));
  NAND3_X1  g360(.A1(new_n530), .A2(new_n546), .A3(new_n534), .ZN(new_n547));
  NAND3_X1  g361(.A1(new_n536), .A2(new_n545), .A3(new_n547), .ZN(new_n548));
  INV_X1    g362(.A(KEYINPUT88), .ZN(new_n549));
  INV_X1    g363(.A(KEYINPUT20), .ZN(new_n550));
  NOR2_X1   g364(.A1(G475), .A2(G902), .ZN(new_n551));
  NAND4_X1  g365(.A1(new_n548), .A2(new_n549), .A3(new_n550), .A4(new_n551), .ZN(new_n552));
  INV_X1    g366(.A(new_n545), .ZN(new_n553));
  AOI21_X1  g367(.A(new_n533), .B1(new_n544), .B2(new_n529), .ZN(new_n554));
  OAI21_X1  g368(.A(new_n191), .B1(new_n553), .B2(new_n554), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n555), .A2(G475), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n545), .A2(new_n547), .ZN(new_n557));
  AOI21_X1  g371(.A(new_n546), .B1(new_n530), .B2(new_n534), .ZN(new_n558));
  OAI211_X1 g372(.A(new_n550), .B(new_n551), .C1(new_n557), .C2(new_n558), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n559), .A2(KEYINPUT88), .ZN(new_n560));
  XOR2_X1   g374(.A(KEYINPUT83), .B(KEYINPUT20), .Z(new_n561));
  AOI21_X1  g375(.A(new_n561), .B1(new_n548), .B2(new_n551), .ZN(new_n562));
  OAI211_X1 g376(.A(new_n552), .B(new_n556), .C1(new_n560), .C2(new_n562), .ZN(new_n563));
  NOR3_X1   g377(.A1(new_n471), .A2(new_n509), .A3(new_n563), .ZN(new_n564));
  NAND4_X1  g378(.A1(new_n303), .A2(new_n358), .A3(new_n419), .A4(new_n564), .ZN(new_n565));
  XNOR2_X1  g379(.A(new_n565), .B(KEYINPUT91), .ZN(new_n566));
  NOR2_X1   g380(.A1(new_n228), .A2(new_n229), .ZN(new_n567));
  XOR2_X1   g381(.A(new_n566), .B(new_n567), .Z(G3));
  AOI21_X1  g382(.A(KEYINPUT79), .B1(new_n295), .B2(new_n285), .ZN(new_n569));
  AOI21_X1  g383(.A(new_n271), .B1(new_n291), .B2(new_n293), .ZN(new_n570));
  NOR4_X1   g384(.A1(new_n570), .A2(new_n287), .A3(G469), .A4(G902), .ZN(new_n571));
  OAI21_X1  g385(.A(new_n302), .B1(new_n569), .B2(new_n571), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n351), .A2(new_n355), .ZN(new_n573));
  AND2_X1   g387(.A1(new_n351), .A2(new_n191), .ZN(new_n574));
  OAI21_X1  g388(.A(new_n573), .B1(new_n574), .B2(new_n353), .ZN(new_n575));
  INV_X1    g389(.A(new_n419), .ZN(new_n576));
  NOR2_X1   g390(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  INV_X1    g391(.A(new_n192), .ZN(new_n578));
  NAND3_X1  g392(.A1(new_n572), .A2(new_n577), .A3(new_n578), .ZN(new_n579));
  INV_X1    g393(.A(KEYINPUT92), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  NAND3_X1  g395(.A1(new_n303), .A2(KEYINPUT92), .A3(new_n577), .ZN(new_n582));
  AND2_X1   g396(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  INV_X1    g397(.A(new_n563), .ZN(new_n584));
  INV_X1    g398(.A(KEYINPUT33), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n503), .A2(new_n585), .ZN(new_n586));
  NAND3_X1  g400(.A1(new_n501), .A2(KEYINPUT33), .A3(new_n502), .ZN(new_n587));
  NAND4_X1  g401(.A1(new_n586), .A2(G478), .A3(new_n191), .A4(new_n587), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n504), .A2(new_n505), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  INV_X1    g404(.A(new_n590), .ZN(new_n591));
  NOR2_X1   g405(.A1(new_n584), .A2(new_n591), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n452), .A2(new_n453), .ZN(new_n593));
  INV_X1    g407(.A(new_n453), .ZN(new_n594));
  NAND3_X1  g408(.A1(new_n443), .A2(new_n451), .A3(new_n594), .ZN(new_n595));
  NAND3_X1  g409(.A1(new_n593), .A2(new_n470), .A3(new_n595), .ZN(new_n596));
  NOR2_X1   g410(.A1(new_n596), .A2(new_n468), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n592), .A2(new_n597), .ZN(new_n598));
  INV_X1    g412(.A(new_n598), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n583), .A2(new_n599), .ZN(new_n600));
  XOR2_X1   g414(.A(KEYINPUT34), .B(G104), .Z(new_n601));
  XNOR2_X1  g415(.A(new_n600), .B(new_n601), .ZN(G6));
  OAI21_X1  g416(.A(new_n551), .B1(new_n557), .B2(new_n558), .ZN(new_n603));
  INV_X1    g417(.A(new_n561), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  NAND3_X1  g419(.A1(new_n548), .A2(new_n551), .A3(new_n561), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n607), .A2(new_n556), .ZN(new_n608));
  AND2_X1   g422(.A1(new_n507), .A2(new_n508), .ZN(new_n609));
  NOR4_X1   g423(.A1(new_n596), .A2(new_n608), .A3(new_n609), .A4(new_n468), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n583), .A2(new_n610), .ZN(new_n611));
  XOR2_X1   g425(.A(KEYINPUT35), .B(G107), .Z(new_n612));
  XNOR2_X1  g426(.A(new_n611), .B(new_n612), .ZN(G9));
  NOR3_X1   g427(.A1(new_n403), .A2(KEYINPUT36), .A3(new_n408), .ZN(new_n614));
  NOR2_X1   g428(.A1(new_n408), .A2(KEYINPUT36), .ZN(new_n615));
  AOI21_X1  g429(.A(new_n615), .B1(new_n392), .B2(new_n402), .ZN(new_n616));
  OR2_X1    g430(.A1(new_n614), .A2(new_n616), .ZN(new_n617));
  NOR2_X1   g431(.A1(new_n617), .A2(new_n417), .ZN(new_n618));
  NOR2_X1   g432(.A1(new_n415), .A2(new_n618), .ZN(new_n619));
  NOR2_X1   g433(.A1(new_n575), .A2(new_n619), .ZN(new_n620));
  NAND3_X1  g434(.A1(new_n303), .A2(new_n564), .A3(new_n620), .ZN(new_n621));
  XOR2_X1   g435(.A(KEYINPUT37), .B(G110), .Z(new_n622));
  XNOR2_X1  g436(.A(new_n621), .B(new_n622), .ZN(G12));
  NOR2_X1   g437(.A1(new_n458), .A2(G900), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n467), .A2(new_n624), .ZN(new_n625));
  INV_X1    g439(.A(KEYINPUT93), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  NAND3_X1  g441(.A1(new_n467), .A2(KEYINPUT93), .A3(new_n624), .ZN(new_n628));
  AND3_X1   g442(.A1(new_n627), .A2(new_n461), .A3(new_n628), .ZN(new_n629));
  INV_X1    g443(.A(new_n629), .ZN(new_n630));
  NAND4_X1  g444(.A1(new_n607), .A2(new_n509), .A3(new_n556), .A4(new_n630), .ZN(new_n631));
  NOR2_X1   g445(.A1(new_n631), .A2(new_n596), .ZN(new_n632));
  INV_X1    g446(.A(new_n619), .ZN(new_n633));
  AND3_X1   g447(.A1(new_n632), .A2(new_n358), .A3(new_n633), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n303), .A2(new_n634), .ZN(new_n635));
  NAND2_X1  g449(.A1(new_n635), .A2(KEYINPUT94), .ZN(new_n636));
  INV_X1    g450(.A(KEYINPUT94), .ZN(new_n637));
  NAND3_X1  g451(.A1(new_n303), .A2(new_n634), .A3(new_n637), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n636), .A2(new_n638), .ZN(new_n639));
  XNOR2_X1  g453(.A(new_n639), .B(G128), .ZN(G30));
  XOR2_X1   g454(.A(new_n629), .B(KEYINPUT39), .Z(new_n641));
  NAND2_X1  g455(.A1(new_n303), .A2(new_n641), .ZN(new_n642));
  OR2_X1    g456(.A1(new_n642), .A2(KEYINPUT40), .ZN(new_n643));
  XNOR2_X1  g457(.A(KEYINPUT96), .B(KEYINPUT38), .ZN(new_n644));
  XNOR2_X1  g458(.A(new_n644), .B(KEYINPUT95), .ZN(new_n645));
  XNOR2_X1  g459(.A(new_n457), .B(new_n645), .ZN(new_n646));
  AND3_X1   g460(.A1(new_n563), .A2(new_n470), .A3(new_n509), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n647), .A2(new_n619), .ZN(new_n648));
  INV_X1    g462(.A(KEYINPUT99), .ZN(new_n649));
  OAI21_X1  g463(.A(new_n646), .B1(new_n648), .B2(new_n649), .ZN(new_n650));
  AOI21_X1  g464(.A(new_n650), .B1(new_n649), .B2(new_n648), .ZN(new_n651));
  NAND2_X1  g465(.A1(new_n642), .A2(KEYINPUT40), .ZN(new_n652));
  OR2_X1    g466(.A1(new_n356), .A2(new_n357), .ZN(new_n653));
  AND2_X1   g467(.A1(new_n317), .A2(new_n319), .ZN(new_n654));
  OAI21_X1  g468(.A(new_n346), .B1(new_n654), .B2(new_n329), .ZN(new_n655));
  AOI21_X1  g469(.A(G902), .B1(new_n655), .B2(KEYINPUT97), .ZN(new_n656));
  OAI21_X1  g470(.A(new_n656), .B1(KEYINPUT97), .B2(new_n655), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n657), .A2(G472), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n653), .A2(new_n658), .ZN(new_n659));
  NAND2_X1  g473(.A1(new_n659), .A2(KEYINPUT98), .ZN(new_n660));
  INV_X1    g474(.A(KEYINPUT98), .ZN(new_n661));
  NAND3_X1  g475(.A1(new_n653), .A2(new_n661), .A3(new_n658), .ZN(new_n662));
  NAND2_X1  g476(.A1(new_n660), .A2(new_n662), .ZN(new_n663));
  NAND4_X1  g477(.A1(new_n643), .A2(new_n651), .A3(new_n652), .A4(new_n663), .ZN(new_n664));
  XNOR2_X1  g478(.A(new_n664), .B(G143), .ZN(G45));
  NAND3_X1  g479(.A1(new_n563), .A2(new_n590), .A3(new_n630), .ZN(new_n666));
  NAND2_X1  g480(.A1(new_n666), .A2(KEYINPUT100), .ZN(new_n667));
  INV_X1    g481(.A(new_n596), .ZN(new_n668));
  INV_X1    g482(.A(KEYINPUT100), .ZN(new_n669));
  NAND4_X1  g483(.A1(new_n563), .A2(new_n669), .A3(new_n590), .A4(new_n630), .ZN(new_n670));
  NAND3_X1  g484(.A1(new_n667), .A2(new_n668), .A3(new_n670), .ZN(new_n671));
  INV_X1    g485(.A(KEYINPUT101), .ZN(new_n672));
  NAND2_X1  g486(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  INV_X1    g487(.A(new_n358), .ZN(new_n674));
  NOR2_X1   g488(.A1(new_n674), .A2(new_n619), .ZN(new_n675));
  NAND4_X1  g489(.A1(new_n667), .A2(KEYINPUT101), .A3(new_n668), .A4(new_n670), .ZN(new_n676));
  NAND4_X1  g490(.A1(new_n673), .A2(new_n303), .A3(new_n675), .A4(new_n676), .ZN(new_n677));
  XNOR2_X1  g491(.A(new_n677), .B(G146), .ZN(G48));
  OAI21_X1  g492(.A(G469), .B1(new_n570), .B2(G902), .ZN(new_n679));
  OAI211_X1 g493(.A(new_n578), .B(new_n679), .C1(new_n569), .C2(new_n571), .ZN(new_n680));
  NAND2_X1  g494(.A1(new_n358), .A2(new_n419), .ZN(new_n681));
  NOR3_X1   g495(.A1(new_n680), .A2(new_n598), .A3(new_n681), .ZN(new_n682));
  INV_X1    g496(.A(KEYINPUT102), .ZN(new_n683));
  XNOR2_X1  g497(.A(new_n682), .B(new_n683), .ZN(new_n684));
  XNOR2_X1  g498(.A(KEYINPUT41), .B(G113), .ZN(new_n685));
  XNOR2_X1  g499(.A(new_n684), .B(new_n685), .ZN(G15));
  NOR2_X1   g500(.A1(new_n680), .A2(new_n681), .ZN(new_n687));
  NAND2_X1  g501(.A1(new_n687), .A2(new_n610), .ZN(new_n688));
  XNOR2_X1  g502(.A(new_n688), .B(G116), .ZN(G18));
  INV_X1    g503(.A(new_n680), .ZN(new_n690));
  NOR2_X1   g504(.A1(new_n563), .A2(new_n509), .ZN(new_n691));
  AND4_X1   g505(.A1(new_n358), .A2(new_n597), .A3(new_n691), .A4(new_n633), .ZN(new_n692));
  NAND2_X1  g506(.A1(new_n690), .A2(new_n692), .ZN(new_n693));
  XNOR2_X1  g507(.A(new_n693), .B(G119), .ZN(G21));
  NAND2_X1  g508(.A1(new_n413), .A2(new_n414), .ZN(new_n695));
  NAND2_X1  g509(.A1(new_n695), .A2(new_n360), .ZN(new_n696));
  INV_X1    g510(.A(new_n418), .ZN(new_n697));
  NAND3_X1  g511(.A1(new_n696), .A2(KEYINPUT104), .A3(new_n697), .ZN(new_n698));
  INV_X1    g512(.A(KEYINPUT104), .ZN(new_n699));
  OAI21_X1  g513(.A(new_n699), .B1(new_n415), .B2(new_n418), .ZN(new_n700));
  NAND2_X1  g514(.A1(new_n698), .A2(new_n700), .ZN(new_n701));
  XOR2_X1   g515(.A(new_n355), .B(KEYINPUT103), .Z(new_n702));
  INV_X1    g516(.A(new_n702), .ZN(new_n703));
  AND2_X1   g517(.A1(new_n347), .A2(new_n350), .ZN(new_n704));
  NAND2_X1  g518(.A1(new_n321), .A2(new_n324), .ZN(new_n705));
  NAND2_X1  g519(.A1(new_n705), .A2(new_n331), .ZN(new_n706));
  AOI21_X1  g520(.A(new_n703), .B1(new_n704), .B2(new_n706), .ZN(new_n707));
  AOI21_X1  g521(.A(new_n353), .B1(new_n351), .B2(new_n191), .ZN(new_n708));
  NOR2_X1   g522(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  NAND2_X1  g523(.A1(new_n701), .A2(new_n709), .ZN(new_n710));
  INV_X1    g524(.A(KEYINPUT105), .ZN(new_n711));
  XNOR2_X1  g525(.A(new_n710), .B(new_n711), .ZN(new_n712));
  NAND3_X1  g526(.A1(new_n647), .A2(new_n593), .A3(new_n595), .ZN(new_n713));
  NOR3_X1   g527(.A1(new_n680), .A2(new_n713), .A3(new_n468), .ZN(new_n714));
  NAND2_X1  g528(.A1(new_n712), .A2(new_n714), .ZN(new_n715));
  XOR2_X1   g529(.A(KEYINPUT106), .B(G122), .Z(new_n716));
  XNOR2_X1  g530(.A(new_n715), .B(new_n716), .ZN(G24));
  NOR2_X1   g531(.A1(new_n680), .A2(new_n596), .ZN(new_n718));
  NOR3_X1   g532(.A1(new_n619), .A2(new_n707), .A3(new_n708), .ZN(new_n719));
  AND3_X1   g533(.A1(new_n719), .A2(new_n667), .A3(new_n670), .ZN(new_n720));
  AOI21_X1  g534(.A(KEYINPUT107), .B1(new_n718), .B2(new_n720), .ZN(new_n721));
  NAND4_X1  g535(.A1(new_n297), .A2(new_n578), .A3(new_n668), .A4(new_n679), .ZN(new_n722));
  NAND3_X1  g536(.A1(new_n719), .A2(new_n667), .A3(new_n670), .ZN(new_n723));
  INV_X1    g537(.A(KEYINPUT107), .ZN(new_n724));
  NOR3_X1   g538(.A1(new_n722), .A2(new_n723), .A3(new_n724), .ZN(new_n725));
  NOR2_X1   g539(.A1(new_n721), .A2(new_n725), .ZN(new_n726));
  XNOR2_X1  g540(.A(new_n726), .B(new_n369), .ZN(G27));
  INV_X1    g541(.A(KEYINPUT108), .ZN(new_n728));
  NAND3_X1  g542(.A1(new_n298), .A2(new_n728), .A3(new_n196), .ZN(new_n729));
  AOI22_X1  g543(.A1(new_n266), .A2(new_n267), .B1(new_n278), .B2(new_n279), .ZN(new_n730));
  OAI21_X1  g544(.A(KEYINPUT108), .B1(new_n730), .B2(new_n197), .ZN(new_n731));
  NAND3_X1  g545(.A1(new_n729), .A2(new_n731), .A3(new_n300), .ZN(new_n732));
  AOI21_X1  g546(.A(new_n285), .B1(new_n732), .B2(new_n191), .ZN(new_n733));
  AOI21_X1  g547(.A(new_n733), .B1(new_n288), .B2(new_n296), .ZN(new_n734));
  OAI21_X1  g548(.A(KEYINPUT109), .B1(new_n734), .B2(new_n192), .ZN(new_n735));
  INV_X1    g549(.A(new_n733), .ZN(new_n736));
  OAI21_X1  g550(.A(new_n736), .B1(new_n569), .B2(new_n571), .ZN(new_n737));
  INV_X1    g551(.A(KEYINPUT109), .ZN(new_n738));
  NAND3_X1  g552(.A1(new_n737), .A2(new_n738), .A3(new_n578), .ZN(new_n739));
  NAND2_X1  g553(.A1(new_n667), .A2(new_n670), .ZN(new_n740));
  INV_X1    g554(.A(new_n740), .ZN(new_n741));
  NAND3_X1  g555(.A1(new_n455), .A2(new_n456), .A3(new_n470), .ZN(new_n742));
  NOR2_X1   g556(.A1(new_n681), .A2(new_n742), .ZN(new_n743));
  NAND4_X1  g557(.A1(new_n735), .A2(new_n739), .A3(new_n741), .A4(new_n743), .ZN(new_n744));
  INV_X1    g558(.A(KEYINPUT42), .ZN(new_n745));
  NAND2_X1  g559(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  NAND3_X1  g560(.A1(new_n358), .A2(new_n701), .A3(KEYINPUT42), .ZN(new_n747));
  NOR2_X1   g561(.A1(new_n740), .A2(new_n747), .ZN(new_n748));
  INV_X1    g562(.A(new_n742), .ZN(new_n749));
  NAND4_X1  g563(.A1(new_n748), .A2(new_n735), .A3(new_n739), .A4(new_n749), .ZN(new_n750));
  INV_X1    g564(.A(KEYINPUT110), .ZN(new_n751));
  AND2_X1   g565(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  NOR2_X1   g566(.A1(new_n750), .A2(new_n751), .ZN(new_n753));
  OAI21_X1  g567(.A(new_n746), .B1(new_n752), .B2(new_n753), .ZN(new_n754));
  XNOR2_X1  g568(.A(new_n754), .B(G131), .ZN(G33));
  INV_X1    g569(.A(new_n631), .ZN(new_n756));
  NAND4_X1  g570(.A1(new_n735), .A2(new_n739), .A3(new_n756), .A4(new_n743), .ZN(new_n757));
  XNOR2_X1  g571(.A(new_n757), .B(G134), .ZN(G36));
  NAND2_X1  g572(.A1(new_n584), .A2(new_n590), .ZN(new_n759));
  INV_X1    g573(.A(KEYINPUT43), .ZN(new_n760));
  OR3_X1    g574(.A1(new_n759), .A2(KEYINPUT112), .A3(new_n760), .ZN(new_n761));
  OAI21_X1  g575(.A(KEYINPUT112), .B1(new_n759), .B2(new_n760), .ZN(new_n762));
  NAND2_X1  g576(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  AOI21_X1  g577(.A(KEYINPUT43), .B1(new_n584), .B2(new_n590), .ZN(new_n764));
  NOR2_X1   g578(.A1(new_n764), .A2(KEYINPUT111), .ZN(new_n765));
  AND2_X1   g579(.A1(new_n764), .A2(KEYINPUT111), .ZN(new_n766));
  OAI21_X1  g580(.A(new_n763), .B1(new_n765), .B2(new_n766), .ZN(new_n767));
  AND3_X1   g581(.A1(new_n767), .A2(new_n575), .A3(new_n633), .ZN(new_n768));
  OR3_X1    g582(.A1(new_n768), .A2(KEYINPUT113), .A3(KEYINPUT44), .ZN(new_n769));
  OAI21_X1  g583(.A(KEYINPUT113), .B1(new_n768), .B2(KEYINPUT44), .ZN(new_n770));
  NAND2_X1  g584(.A1(new_n768), .A2(KEYINPUT44), .ZN(new_n771));
  OAI21_X1  g585(.A(G469), .B1(new_n301), .B2(KEYINPUT45), .ZN(new_n772));
  INV_X1    g586(.A(new_n732), .ZN(new_n773));
  AOI21_X1  g587(.A(new_n772), .B1(KEYINPUT45), .B2(new_n773), .ZN(new_n774));
  NOR2_X1   g588(.A1(new_n285), .A2(new_n191), .ZN(new_n775));
  NOR2_X1   g589(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  OR2_X1    g590(.A1(new_n776), .A2(KEYINPUT46), .ZN(new_n777));
  NAND2_X1  g591(.A1(new_n776), .A2(KEYINPUT46), .ZN(new_n778));
  NAND3_X1  g592(.A1(new_n777), .A2(new_n297), .A3(new_n778), .ZN(new_n779));
  NAND2_X1  g593(.A1(new_n779), .A2(new_n578), .ZN(new_n780));
  INV_X1    g594(.A(new_n641), .ZN(new_n781));
  NOR3_X1   g595(.A1(new_n780), .A2(new_n781), .A3(new_n742), .ZN(new_n782));
  NAND4_X1  g596(.A1(new_n769), .A2(new_n770), .A3(new_n771), .A4(new_n782), .ZN(new_n783));
  XNOR2_X1  g597(.A(new_n783), .B(G137), .ZN(G39));
  NAND4_X1  g598(.A1(new_n741), .A2(new_n674), .A3(new_n576), .A4(new_n749), .ZN(new_n785));
  INV_X1    g599(.A(KEYINPUT47), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n780), .A2(new_n786), .ZN(new_n787));
  NAND3_X1  g601(.A1(new_n779), .A2(KEYINPUT47), .A3(new_n578), .ZN(new_n788));
  AOI21_X1  g602(.A(new_n785), .B1(new_n787), .B2(new_n788), .ZN(new_n789));
  XNOR2_X1  g603(.A(new_n789), .B(new_n362), .ZN(G42));
  NAND2_X1  g604(.A1(new_n767), .A2(new_n462), .ZN(new_n791));
  INV_X1    g605(.A(KEYINPUT118), .ZN(new_n792));
  NAND2_X1  g606(.A1(new_n791), .A2(new_n792), .ZN(new_n793));
  NAND3_X1  g607(.A1(new_n767), .A2(KEYINPUT118), .A3(new_n462), .ZN(new_n794));
  AOI211_X1 g608(.A(new_n680), .B(new_n742), .C1(new_n793), .C2(new_n794), .ZN(new_n795));
  NOR3_X1   g609(.A1(new_n663), .A2(new_n576), .A3(new_n461), .ZN(new_n796));
  NOR2_X1   g610(.A1(new_n680), .A2(new_n742), .ZN(new_n797));
  AND2_X1   g611(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  NOR2_X1   g612(.A1(new_n563), .A2(new_n590), .ZN(new_n799));
  AOI22_X1  g613(.A1(new_n795), .A2(new_n719), .B1(new_n798), .B2(new_n799), .ZN(new_n800));
  INV_X1    g614(.A(new_n712), .ZN(new_n801));
  AOI21_X1  g615(.A(new_n801), .B1(new_n793), .B2(new_n794), .ZN(new_n802));
  INV_X1    g616(.A(new_n679), .ZN(new_n803));
  AOI21_X1  g617(.A(new_n803), .B1(new_n288), .B2(new_n296), .ZN(new_n804));
  NAND2_X1  g618(.A1(new_n804), .A2(new_n192), .ZN(new_n805));
  NAND3_X1  g619(.A1(new_n787), .A2(new_n788), .A3(new_n805), .ZN(new_n806));
  NAND3_X1  g620(.A1(new_n802), .A2(new_n806), .A3(new_n749), .ZN(new_n807));
  NOR3_X1   g621(.A1(new_n646), .A2(new_n680), .A3(new_n470), .ZN(new_n808));
  XNOR2_X1  g622(.A(new_n808), .B(KEYINPUT119), .ZN(new_n809));
  NAND2_X1  g623(.A1(new_n802), .A2(new_n809), .ZN(new_n810));
  XOR2_X1   g624(.A(KEYINPUT120), .B(KEYINPUT50), .Z(new_n811));
  NAND2_X1  g625(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  NOR2_X1   g626(.A1(KEYINPUT120), .A2(KEYINPUT50), .ZN(new_n813));
  NAND3_X1  g627(.A1(new_n802), .A2(new_n809), .A3(new_n813), .ZN(new_n814));
  NAND4_X1  g628(.A1(new_n800), .A2(new_n807), .A3(new_n812), .A4(new_n814), .ZN(new_n815));
  INV_X1    g629(.A(KEYINPUT51), .ZN(new_n816));
  NAND2_X1  g630(.A1(new_n815), .A2(new_n816), .ZN(new_n817));
  NAND2_X1  g631(.A1(new_n802), .A2(new_n718), .ZN(new_n818));
  INV_X1    g632(.A(new_n592), .ZN(new_n819));
  INV_X1    g633(.A(new_n798), .ZN(new_n820));
  OAI21_X1  g634(.A(new_n818), .B1(new_n819), .B2(new_n820), .ZN(new_n821));
  NAND3_X1  g635(.A1(new_n795), .A2(new_n358), .A3(new_n701), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n822), .A2(KEYINPUT48), .ZN(new_n823));
  INV_X1    g637(.A(KEYINPUT48), .ZN(new_n824));
  NAND4_X1  g638(.A1(new_n795), .A2(new_n824), .A3(new_n358), .A4(new_n701), .ZN(new_n825));
  AOI21_X1  g639(.A(new_n821), .B1(new_n823), .B2(new_n825), .ZN(new_n826));
  NAND2_X1  g640(.A1(new_n817), .A2(new_n826), .ZN(new_n827));
  NOR2_X1   g641(.A1(new_n815), .A2(new_n816), .ZN(new_n828));
  NOR2_X1   g642(.A1(new_n827), .A2(new_n828), .ZN(new_n829));
  AND2_X1   g643(.A1(new_n735), .A2(new_n739), .ZN(new_n830));
  NAND4_X1  g644(.A1(new_n830), .A2(KEYINPUT115), .A3(new_n720), .A4(new_n749), .ZN(new_n831));
  NAND4_X1  g645(.A1(new_n735), .A2(new_n720), .A3(new_n739), .A4(new_n749), .ZN(new_n832));
  INV_X1    g646(.A(KEYINPUT115), .ZN(new_n833));
  NAND2_X1  g647(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  NAND2_X1  g648(.A1(new_n831), .A2(new_n834), .ZN(new_n835));
  NOR3_X1   g649(.A1(new_n608), .A2(new_n509), .A3(new_n629), .ZN(new_n836));
  NAND4_X1  g650(.A1(new_n303), .A2(new_n675), .A3(new_n749), .A4(new_n836), .ZN(new_n837));
  NAND2_X1  g651(.A1(new_n757), .A2(new_n837), .ZN(new_n838));
  INV_X1    g652(.A(new_n838), .ZN(new_n839));
  AOI21_X1  g653(.A(KEYINPUT116), .B1(new_n835), .B2(new_n839), .ZN(new_n840));
  INV_X1    g654(.A(KEYINPUT116), .ZN(new_n841));
  AOI211_X1 g655(.A(new_n841), .B(new_n838), .C1(new_n831), .C2(new_n834), .ZN(new_n842));
  NOR2_X1   g656(.A1(new_n840), .A2(new_n842), .ZN(new_n843));
  INV_X1    g657(.A(KEYINPUT114), .ZN(new_n844));
  NAND2_X1  g658(.A1(new_n584), .A2(new_n509), .ZN(new_n845));
  NOR2_X1   g659(.A1(new_n471), .A2(new_n845), .ZN(new_n846));
  NAND3_X1  g660(.A1(new_n581), .A2(new_n582), .A3(new_n846), .ZN(new_n847));
  AOI21_X1  g661(.A(new_n844), .B1(new_n847), .B2(new_n621), .ZN(new_n848));
  NOR2_X1   g662(.A1(new_n819), .A2(new_n471), .ZN(new_n849));
  NAND3_X1  g663(.A1(new_n581), .A2(new_n582), .A3(new_n849), .ZN(new_n850));
  NAND2_X1  g664(.A1(new_n850), .A2(new_n565), .ZN(new_n851));
  NOR2_X1   g665(.A1(new_n848), .A2(new_n851), .ZN(new_n852));
  AND3_X1   g666(.A1(new_n847), .A2(new_n844), .A3(new_n621), .ZN(new_n853));
  INV_X1    g667(.A(new_n853), .ZN(new_n854));
  AOI22_X1  g668(.A1(new_n687), .A2(new_n610), .B1(new_n690), .B2(new_n692), .ZN(new_n855));
  NOR2_X1   g669(.A1(new_n682), .A2(new_n683), .ZN(new_n856));
  NOR4_X1   g670(.A1(new_n680), .A2(new_n598), .A3(new_n681), .A4(KEYINPUT102), .ZN(new_n857));
  OAI211_X1 g671(.A(new_n715), .B(new_n855), .C1(new_n856), .C2(new_n857), .ZN(new_n858));
  INV_X1    g672(.A(new_n858), .ZN(new_n859));
  NAND4_X1  g673(.A1(new_n852), .A2(new_n754), .A3(new_n854), .A4(new_n859), .ZN(new_n860));
  NOR2_X1   g674(.A1(new_n843), .A2(new_n860), .ZN(new_n861));
  INV_X1    g675(.A(KEYINPUT117), .ZN(new_n862));
  NAND3_X1  g676(.A1(new_n619), .A2(new_n578), .A3(new_n630), .ZN(new_n863));
  NOR3_X1   g677(.A1(new_n713), .A2(new_n734), .A3(new_n863), .ZN(new_n864));
  NAND2_X1  g678(.A1(new_n663), .A2(new_n864), .ZN(new_n865));
  OAI21_X1  g679(.A(new_n865), .B1(new_n721), .B2(new_n725), .ZN(new_n866));
  AND3_X1   g680(.A1(new_n303), .A2(new_n634), .A3(new_n637), .ZN(new_n867));
  AOI21_X1  g681(.A(new_n637), .B1(new_n303), .B2(new_n634), .ZN(new_n868));
  NAND3_X1  g682(.A1(new_n303), .A2(new_n675), .A3(new_n676), .ZN(new_n869));
  AND2_X1   g683(.A1(new_n671), .A2(new_n672), .ZN(new_n870));
  OAI22_X1  g684(.A1(new_n867), .A2(new_n868), .B1(new_n869), .B2(new_n870), .ZN(new_n871));
  OAI21_X1  g685(.A(KEYINPUT52), .B1(new_n866), .B2(new_n871), .ZN(new_n872));
  NAND3_X1  g686(.A1(new_n718), .A2(KEYINPUT107), .A3(new_n720), .ZN(new_n873));
  OAI21_X1  g687(.A(new_n724), .B1(new_n722), .B2(new_n723), .ZN(new_n874));
  AOI22_X1  g688(.A1(new_n873), .A2(new_n874), .B1(new_n864), .B2(new_n663), .ZN(new_n875));
  INV_X1    g689(.A(KEYINPUT52), .ZN(new_n876));
  NAND4_X1  g690(.A1(new_n875), .A2(new_n876), .A3(new_n639), .A4(new_n677), .ZN(new_n877));
  AOI21_X1  g691(.A(new_n862), .B1(new_n872), .B2(new_n877), .ZN(new_n878));
  INV_X1    g692(.A(new_n878), .ZN(new_n879));
  NAND3_X1  g693(.A1(new_n872), .A2(new_n877), .A3(new_n862), .ZN(new_n880));
  NAND2_X1  g694(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  NAND3_X1  g695(.A1(new_n861), .A2(KEYINPUT53), .A3(new_n881), .ZN(new_n882));
  INV_X1    g696(.A(KEYINPUT53), .ZN(new_n883));
  NOR3_X1   g697(.A1(new_n853), .A2(new_n848), .A3(new_n851), .ZN(new_n884));
  XNOR2_X1  g698(.A(new_n750), .B(new_n751), .ZN(new_n885));
  AOI21_X1  g699(.A(new_n858), .B1(new_n885), .B2(new_n746), .ZN(new_n886));
  OAI211_X1 g700(.A(new_n884), .B(new_n886), .C1(new_n840), .C2(new_n842), .ZN(new_n887));
  NAND2_X1  g701(.A1(new_n872), .A2(new_n877), .ZN(new_n888));
  OAI21_X1  g702(.A(new_n883), .B1(new_n887), .B2(new_n888), .ZN(new_n889));
  NAND2_X1  g703(.A1(new_n882), .A2(new_n889), .ZN(new_n890));
  NAND2_X1  g704(.A1(new_n890), .A2(KEYINPUT54), .ZN(new_n891));
  AND3_X1   g705(.A1(new_n872), .A2(new_n862), .A3(new_n877), .ZN(new_n892));
  NOR2_X1   g706(.A1(new_n892), .A2(new_n878), .ZN(new_n893));
  OAI21_X1  g707(.A(new_n883), .B1(new_n893), .B2(new_n887), .ZN(new_n894));
  INV_X1    g708(.A(new_n860), .ZN(new_n895));
  AOI21_X1  g709(.A(new_n838), .B1(new_n831), .B2(new_n834), .ZN(new_n896));
  XNOR2_X1  g710(.A(new_n896), .B(KEYINPUT116), .ZN(new_n897));
  INV_X1    g711(.A(new_n888), .ZN(new_n898));
  NAND4_X1  g712(.A1(new_n895), .A2(new_n897), .A3(KEYINPUT53), .A4(new_n898), .ZN(new_n899));
  NAND2_X1  g713(.A1(new_n894), .A2(new_n899), .ZN(new_n900));
  OR2_X1    g714(.A1(new_n900), .A2(KEYINPUT54), .ZN(new_n901));
  NAND3_X1  g715(.A1(new_n829), .A2(new_n891), .A3(new_n901), .ZN(new_n902));
  OAI21_X1  g716(.A(G953), .B1(new_n902), .B2(KEYINPUT121), .ZN(new_n903));
  NAND4_X1  g717(.A1(new_n829), .A2(KEYINPUT121), .A3(new_n891), .A4(new_n901), .ZN(new_n904));
  NAND2_X1  g718(.A1(new_n904), .A2(new_n459), .ZN(new_n905));
  XOR2_X1   g719(.A(new_n804), .B(KEYINPUT49), .Z(new_n906));
  NAND3_X1  g720(.A1(new_n701), .A2(new_n578), .A3(new_n470), .ZN(new_n907));
  OR2_X1    g721(.A1(new_n646), .A2(new_n907), .ZN(new_n908));
  OR4_X1    g722(.A1(new_n663), .A2(new_n906), .A3(new_n759), .A4(new_n908), .ZN(new_n909));
  NAND3_X1  g723(.A1(new_n903), .A2(new_n905), .A3(new_n909), .ZN(G75));
  OAI21_X1  g724(.A(new_n432), .B1(new_n441), .B2(new_n442), .ZN(new_n911));
  XNOR2_X1  g725(.A(new_n911), .B(new_n439), .ZN(new_n912));
  XOR2_X1   g726(.A(new_n912), .B(KEYINPUT55), .Z(new_n913));
  AOI21_X1  g727(.A(new_n191), .B1(new_n894), .B2(new_n899), .ZN(new_n914));
  AND2_X1   g728(.A1(new_n914), .A2(G210), .ZN(new_n915));
  OAI211_X1 g729(.A(KEYINPUT122), .B(new_n913), .C1(new_n915), .C2(KEYINPUT56), .ZN(new_n916));
  INV_X1    g730(.A(KEYINPUT122), .ZN(new_n917));
  AOI21_X1  g731(.A(KEYINPUT56), .B1(new_n914), .B2(G210), .ZN(new_n918));
  INV_X1    g732(.A(new_n913), .ZN(new_n919));
  OAI21_X1  g733(.A(new_n917), .B1(new_n918), .B2(new_n919), .ZN(new_n920));
  NAND2_X1  g734(.A1(new_n916), .A2(new_n920), .ZN(new_n921));
  NOR2_X1   g735(.A1(new_n458), .A2(G952), .ZN(new_n922));
  XNOR2_X1  g736(.A(new_n922), .B(KEYINPUT124), .ZN(new_n923));
  INV_X1    g737(.A(new_n923), .ZN(new_n924));
  NAND2_X1  g738(.A1(new_n900), .A2(G902), .ZN(new_n925));
  INV_X1    g739(.A(KEYINPUT123), .ZN(new_n926));
  NAND2_X1  g740(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  NAND2_X1  g741(.A1(new_n914), .A2(KEYINPUT123), .ZN(new_n928));
  NAND3_X1  g742(.A1(new_n927), .A2(new_n594), .A3(new_n928), .ZN(new_n929));
  NOR2_X1   g743(.A1(new_n913), .A2(KEYINPUT56), .ZN(new_n930));
  AOI21_X1  g744(.A(new_n924), .B1(new_n929), .B2(new_n930), .ZN(new_n931));
  AND2_X1   g745(.A1(new_n921), .A2(new_n931), .ZN(G51));
  XNOR2_X1  g746(.A(new_n900), .B(KEYINPUT54), .ZN(new_n933));
  XNOR2_X1  g747(.A(new_n775), .B(KEYINPUT57), .ZN(new_n934));
  NAND2_X1  g748(.A1(new_n933), .A2(new_n934), .ZN(new_n935));
  NAND2_X1  g749(.A1(new_n935), .A2(new_n284), .ZN(new_n936));
  NAND3_X1  g750(.A1(new_n927), .A2(new_n774), .A3(new_n928), .ZN(new_n937));
  AOI21_X1  g751(.A(new_n922), .B1(new_n936), .B2(new_n937), .ZN(G54));
  AND2_X1   g752(.A1(KEYINPUT58), .A2(G475), .ZN(new_n939));
  NAND3_X1  g753(.A1(new_n927), .A2(new_n928), .A3(new_n939), .ZN(new_n940));
  INV_X1    g754(.A(new_n548), .ZN(new_n941));
  NAND2_X1  g755(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  INV_X1    g756(.A(new_n922), .ZN(new_n943));
  NAND2_X1  g757(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  NOR2_X1   g758(.A1(new_n940), .A2(new_n941), .ZN(new_n945));
  NOR2_X1   g759(.A1(new_n944), .A2(new_n945), .ZN(G60));
  AND2_X1   g760(.A1(new_n586), .A2(new_n587), .ZN(new_n947));
  NAND2_X1  g761(.A1(G478), .A2(G902), .ZN(new_n948));
  XNOR2_X1  g762(.A(new_n948), .B(KEYINPUT59), .ZN(new_n949));
  AND3_X1   g763(.A1(new_n933), .A2(new_n947), .A3(new_n949), .ZN(new_n950));
  NAND2_X1  g764(.A1(new_n901), .A2(new_n891), .ZN(new_n951));
  AOI21_X1  g765(.A(new_n947), .B1(new_n951), .B2(new_n949), .ZN(new_n952));
  NOR3_X1   g766(.A1(new_n950), .A2(new_n952), .A3(new_n924), .ZN(G63));
  NAND2_X1  g767(.A1(G217), .A2(G902), .ZN(new_n954));
  XNOR2_X1  g768(.A(new_n954), .B(KEYINPUT60), .ZN(new_n955));
  INV_X1    g769(.A(new_n955), .ZN(new_n956));
  AOI21_X1  g770(.A(KEYINPUT53), .B1(new_n861), .B2(new_n881), .ZN(new_n957));
  NOR3_X1   g771(.A1(new_n887), .A2(new_n883), .A3(new_n888), .ZN(new_n958));
  OAI21_X1  g772(.A(new_n956), .B1(new_n957), .B2(new_n958), .ZN(new_n959));
  NAND2_X1  g773(.A1(new_n959), .A2(KEYINPUT125), .ZN(new_n960));
  INV_X1    g774(.A(KEYINPUT125), .ZN(new_n961));
  NAND3_X1  g775(.A1(new_n900), .A2(new_n961), .A3(new_n956), .ZN(new_n962));
  NAND3_X1  g776(.A1(new_n960), .A2(new_n416), .A3(new_n962), .ZN(new_n963));
  INV_X1    g777(.A(new_n617), .ZN(new_n964));
  AOI21_X1  g778(.A(new_n961), .B1(new_n900), .B2(new_n956), .ZN(new_n965));
  AOI211_X1 g779(.A(KEYINPUT125), .B(new_n955), .C1(new_n894), .C2(new_n899), .ZN(new_n966));
  OAI21_X1  g780(.A(new_n964), .B1(new_n965), .B2(new_n966), .ZN(new_n967));
  NAND3_X1  g781(.A1(new_n963), .A2(new_n967), .A3(new_n923), .ZN(new_n968));
  INV_X1    g782(.A(KEYINPUT61), .ZN(new_n969));
  NAND2_X1  g783(.A1(new_n968), .A2(new_n969), .ZN(new_n970));
  NAND4_X1  g784(.A1(new_n963), .A2(new_n967), .A3(KEYINPUT61), .A4(new_n923), .ZN(new_n971));
  NAND2_X1  g785(.A1(new_n970), .A2(new_n971), .ZN(G66));
  AND2_X1   g786(.A1(new_n435), .A2(G953), .ZN(new_n973));
  NAND2_X1  g787(.A1(new_n884), .A2(new_n859), .ZN(new_n974));
  AOI211_X1 g788(.A(new_n466), .B(new_n973), .C1(new_n974), .C2(new_n458), .ZN(new_n975));
  OAI21_X1  g789(.A(new_n911), .B1(G898), .B2(new_n458), .ZN(new_n976));
  XOR2_X1   g790(.A(new_n975), .B(new_n976), .Z(G69));
  OAI21_X1  g791(.A(new_n519), .B1(new_n520), .B2(new_n521), .ZN(new_n978));
  XNOR2_X1  g792(.A(new_n338), .B(new_n978), .ZN(new_n979));
  AOI211_X1 g793(.A(new_n674), .B(new_n713), .C1(new_n700), .C2(new_n698), .ZN(new_n980));
  NAND4_X1  g794(.A1(new_n779), .A2(new_n578), .A3(new_n641), .A4(new_n980), .ZN(new_n981));
  NAND2_X1  g795(.A1(new_n981), .A2(new_n757), .ZN(new_n982));
  NOR2_X1   g796(.A1(new_n789), .A2(new_n982), .ZN(new_n983));
  NOR2_X1   g797(.A1(new_n871), .A2(new_n726), .ZN(new_n984));
  NAND3_X1  g798(.A1(new_n783), .A2(new_n983), .A3(new_n984), .ZN(new_n985));
  INV_X1    g799(.A(new_n754), .ZN(new_n986));
  OAI21_X1  g800(.A(new_n458), .B1(new_n985), .B2(new_n986), .ZN(new_n987));
  XNOR2_X1  g801(.A(new_n624), .B(KEYINPUT127), .ZN(new_n988));
  AOI21_X1  g802(.A(new_n979), .B1(new_n987), .B2(new_n988), .ZN(new_n989));
  INV_X1    g803(.A(new_n743), .ZN(new_n990));
  AOI211_X1 g804(.A(new_n990), .B(new_n642), .C1(new_n819), .C2(new_n845), .ZN(new_n991));
  NOR2_X1   g805(.A1(new_n789), .A2(new_n991), .ZN(new_n992));
  NAND2_X1  g806(.A1(new_n984), .A2(new_n664), .ZN(new_n993));
  OR2_X1    g807(.A1(new_n993), .A2(KEYINPUT62), .ZN(new_n994));
  NAND2_X1  g808(.A1(new_n993), .A2(KEYINPUT62), .ZN(new_n995));
  NAND4_X1  g809(.A1(new_n783), .A2(new_n992), .A3(new_n994), .A4(new_n995), .ZN(new_n996));
  NAND2_X1  g810(.A1(new_n996), .A2(new_n458), .ZN(new_n997));
  AOI21_X1  g811(.A(new_n989), .B1(new_n997), .B2(new_n979), .ZN(new_n998));
  INV_X1    g812(.A(G900), .ZN(new_n999));
  OAI21_X1  g813(.A(G953), .B1(new_n194), .B2(new_n999), .ZN(new_n1000));
  OAI21_X1  g814(.A(new_n1000), .B1(new_n989), .B2(KEYINPUT126), .ZN(new_n1001));
  XOR2_X1   g815(.A(new_n998), .B(new_n1001), .Z(G72));
  NAND2_X1  g816(.A1(G472), .A2(G902), .ZN(new_n1003));
  XOR2_X1   g817(.A(new_n1003), .B(KEYINPUT63), .Z(new_n1004));
  OR2_X1    g818(.A1(new_n985), .A2(new_n986), .ZN(new_n1005));
  OAI21_X1  g819(.A(new_n1004), .B1(new_n1005), .B2(new_n974), .ZN(new_n1006));
  NAND3_X1  g820(.A1(new_n1006), .A2(new_n331), .A3(new_n339), .ZN(new_n1007));
  NOR2_X1   g821(.A1(new_n339), .A2(new_n331), .ZN(new_n1008));
  INV_X1    g822(.A(new_n1008), .ZN(new_n1009));
  NAND2_X1  g823(.A1(new_n339), .A2(new_n331), .ZN(new_n1010));
  NAND4_X1  g824(.A1(new_n890), .A2(new_n1009), .A3(new_n1004), .A4(new_n1010), .ZN(new_n1011));
  OAI21_X1  g825(.A(new_n1004), .B1(new_n996), .B2(new_n974), .ZN(new_n1012));
  NAND2_X1  g826(.A1(new_n1012), .A2(new_n1008), .ZN(new_n1013));
  AND4_X1   g827(.A1(new_n943), .A2(new_n1007), .A3(new_n1011), .A4(new_n1013), .ZN(G57));
endmodule


