

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372,
         n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383,
         n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394,
         n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405,
         n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416,
         n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427,
         n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438,
         n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449,
         n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460,
         n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471,
         n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482,
         n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493,
         n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504,
         n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515,
         n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526,
         n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537,
         n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
         n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559,
         n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570,
         n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581,
         n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592,
         n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603,
         n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614,
         n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625,
         n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636,
         n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647,
         n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658,
         n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669,
         n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680,
         n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691,
         n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702,
         n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713,
         n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724,
         n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735,
         n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746,
         n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757,
         n758, n759, n760, n761, n762, n763, n764, n765;

  XNOR2_X1 U383 ( .A(n398), .B(KEYINPUT65), .ZN(n446) );
  INV_X4 U384 ( .A(G953), .ZN(n756) );
  NOR2_X1 U385 ( .A1(n667), .A2(n761), .ZN(n619) );
  XNOR2_X1 U386 ( .A(KEYINPUT64), .B(KEYINPUT4), .ZN(n438) );
  XNOR2_X1 U387 ( .A(G113), .B(G116), .ZN(n428) );
  AND2_X4 U388 ( .A1(n391), .A2(n390), .ZN(n648) );
  XNOR2_X2 U389 ( .A(n577), .B(n370), .ZN(n717) );
  XNOR2_X2 U390 ( .A(n380), .B(KEYINPUT22), .ZN(n615) );
  NOR2_X1 U391 ( .A1(n763), .A2(n764), .ZN(n532) );
  AND2_X1 U392 ( .A1(n411), .A2(n409), .ZN(n408) );
  NAND2_X1 U393 ( .A1(n404), .A2(n405), .ZN(n407) );
  NOR2_X1 U394 ( .A1(n557), .A2(n401), .ZN(n400) );
  NOR2_X1 U395 ( .A1(n547), .A2(n680), .ZN(n402) );
  XNOR2_X1 U396 ( .A(n532), .B(KEYINPUT46), .ZN(n399) );
  XNOR2_X1 U397 ( .A(n522), .B(n521), .ZN(n706) );
  AND2_X1 U398 ( .A1(n425), .A2(n695), .ZN(n575) );
  XNOR2_X1 U399 ( .A(n540), .B(n422), .ZN(n425) );
  XNOR2_X1 U400 ( .A(n426), .B(n475), .ZN(n540) );
  XNOR2_X1 U401 ( .A(n379), .B(n374), .ZN(n652) );
  XNOR2_X1 U402 ( .A(n378), .B(n375), .ZN(n374) );
  XNOR2_X1 U403 ( .A(n472), .B(n741), .ZN(n379) );
  XNOR2_X1 U404 ( .A(n397), .B(n368), .ZN(n378) );
  XNOR2_X1 U405 ( .A(n377), .B(n376), .ZN(n375) );
  XNOR2_X1 U406 ( .A(n446), .B(n432), .ZN(n377) );
  XNOR2_X1 U407 ( .A(n436), .B(n438), .ZN(n376) );
  XNOR2_X1 U408 ( .A(G902), .B(KEYINPUT15), .ZN(n624) );
  XNOR2_X1 U409 ( .A(G104), .B(G107), .ZN(n430) );
  INV_X1 U410 ( .A(n569), .ZN(n362) );
  AND2_X1 U411 ( .A1(n387), .A2(n372), .ZN(n386) );
  XOR2_X2 U412 ( .A(G110), .B(KEYINPUT90), .Z(n364) );
  XOR2_X1 U413 ( .A(KEYINPUT99), .B(KEYINPUT5), .Z(n440) );
  XNOR2_X1 U414 ( .A(n445), .B(G125), .ZN(n453) );
  XNOR2_X1 U415 ( .A(n508), .B(n439), .ZN(n473) );
  INV_X1 U416 ( .A(G101), .ZN(n398) );
  XNOR2_X1 U417 ( .A(G137), .B(G140), .ZN(n459) );
  XNOR2_X1 U418 ( .A(n458), .B(n454), .ZN(n396) );
  XNOR2_X1 U419 ( .A(KEYINPUT96), .B(KEYINPUT72), .ZN(n454) );
  AND2_X1 U420 ( .A1(n506), .A2(G221), .ZN(n393) );
  XNOR2_X1 U421 ( .A(n436), .B(G134), .ZN(n508) );
  XNOR2_X1 U422 ( .A(KEYINPUT9), .B(KEYINPUT104), .ZN(n501) );
  XOR2_X1 U423 ( .A(G107), .B(KEYINPUT7), .Z(n502) );
  XNOR2_X1 U424 ( .A(G143), .B(G113), .ZN(n489) );
  XNOR2_X1 U425 ( .A(n453), .B(n395), .ZN(n485) );
  INV_X1 U426 ( .A(KEYINPUT10), .ZN(n395) );
  XNOR2_X1 U427 ( .A(n487), .B(G122), .ZN(n488) );
  NAND2_X1 U428 ( .A1(n624), .A2(n623), .ZN(n415) );
  XNOR2_X1 U429 ( .A(n534), .B(KEYINPUT86), .ZN(n552) );
  NOR2_X1 U430 ( .A1(n593), .A2(n482), .ZN(n542) );
  AND2_X1 U431 ( .A1(n603), .A2(n363), .ZN(n404) );
  OR2_X1 U432 ( .A1(G237), .A2(G902), .ZN(n449) );
  NAND2_X1 U433 ( .A1(n623), .A2(n421), .ZN(n419) );
  INV_X1 U434 ( .A(n624), .ZN(n420) );
  INV_X1 U435 ( .A(n453), .ZN(n397) );
  NOR2_X1 U436 ( .A1(n708), .A2(n709), .ZN(n518) );
  XNOR2_X1 U437 ( .A(n533), .B(KEYINPUT38), .ZN(n708) );
  INV_X1 U438 ( .A(G902), .ZN(n498) );
  INV_X1 U439 ( .A(KEYINPUT1), .ZN(n422) );
  XNOR2_X1 U440 ( .A(n444), .B(n373), .ZN(n630) );
  XNOR2_X1 U441 ( .A(n443), .B(n470), .ZN(n373) );
  XNOR2_X1 U442 ( .A(KEYINPUT69), .B(KEYINPUT70), .ZN(n431) );
  INV_X1 U443 ( .A(KEYINPUT19), .ZN(n551) );
  BUF_X1 U444 ( .A(n523), .Z(n699) );
  XNOR2_X1 U445 ( .A(G122), .B(KEYINPUT16), .ZN(n429) );
  XNOR2_X1 U446 ( .A(n393), .B(n460), .ZN(n392) );
  XNOR2_X1 U447 ( .A(n396), .B(n485), .ZN(n394) );
  XNOR2_X1 U448 ( .A(G116), .B(G122), .ZN(n504) );
  XNOR2_X1 U449 ( .A(n485), .B(n488), .ZN(n497) );
  NAND2_X1 U450 ( .A1(n386), .A2(n385), .ZN(n391) );
  XNOR2_X1 U451 ( .A(n516), .B(KEYINPUT40), .ZN(n763) );
  NAND2_X1 U452 ( .A1(n588), .A2(n587), .ZN(n589) );
  XNOR2_X1 U453 ( .A(n586), .B(n585), .ZN(n588) );
  INV_X1 U454 ( .A(KEYINPUT34), .ZN(n585) );
  XNOR2_X1 U455 ( .A(n515), .B(KEYINPUT107), .ZN(n671) );
  NAND2_X1 U456 ( .A1(n543), .A2(n388), .ZN(n544) );
  AND2_X1 U457 ( .A1(n389), .A2(n542), .ZN(n388) );
  AND2_X1 U458 ( .A1(n587), .A2(n362), .ZN(n389) );
  AND2_X1 U459 ( .A1(n602), .A2(KEYINPUT84), .ZN(n363) );
  XOR2_X1 U460 ( .A(n434), .B(n433), .Z(n365) );
  AND2_X1 U461 ( .A1(n491), .A2(G210), .ZN(n366) );
  XOR2_X1 U462 ( .A(KEYINPUT23), .B(G110), .Z(n367) );
  XNOR2_X1 U463 ( .A(n622), .B(n621), .ZN(n735) );
  INV_X1 U464 ( .A(n735), .ZN(n383) );
  XNOR2_X1 U465 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n368) );
  INV_X1 U466 ( .A(n425), .ZN(n694) );
  INV_X1 U467 ( .A(G146), .ZN(n445) );
  XOR2_X1 U468 ( .A(KEYINPUT88), .B(KEYINPUT0), .Z(n369) );
  XOR2_X1 U469 ( .A(n576), .B(KEYINPUT33), .Z(n370) );
  XNOR2_X1 U470 ( .A(n394), .B(n392), .ZN(n731) );
  XNOR2_X1 U471 ( .A(KEYINPUT48), .B(KEYINPUT83), .ZN(n371) );
  AND2_X1 U472 ( .A1(n416), .A2(n415), .ZN(n372) );
  INV_X1 U473 ( .A(n418), .ZN(n417) );
  NAND2_X1 U474 ( .A1(n420), .A2(n419), .ZN(n418) );
  NAND2_X1 U475 ( .A1(n648), .A2(G210), .ZN(n654) );
  XNOR2_X2 U476 ( .A(n442), .B(n429), .ZN(n741) );
  XNOR2_X2 U477 ( .A(n427), .B(n428), .ZN(n442) );
  XNOR2_X2 U478 ( .A(n740), .B(n431), .ZN(n472) );
  XNOR2_X2 U479 ( .A(n364), .B(n430), .ZN(n740) );
  NAND2_X1 U480 ( .A1(n599), .A2(n598), .ZN(n380) );
  XNOR2_X2 U481 ( .A(n381), .B(n369), .ZN(n599) );
  OR2_X2 U482 ( .A1(n584), .A2(n583), .ZN(n381) );
  NAND2_X1 U483 ( .A1(n383), .A2(n384), .ZN(n687) );
  NAND2_X1 U484 ( .A1(n382), .A2(n383), .ZN(n387) );
  NOR2_X1 U485 ( .A1(n753), .A2(n418), .ZN(n382) );
  INV_X1 U486 ( .A(n753), .ZN(n384) );
  NAND2_X1 U487 ( .A1(n687), .A2(n623), .ZN(n385) );
  XNOR2_X1 U488 ( .A(n451), .B(KEYINPUT30), .ZN(n543) );
  INV_X1 U489 ( .A(n689), .ZN(n390) );
  NAND2_X1 U490 ( .A1(n414), .A2(n413), .ZN(n622) );
  NOR2_X2 U491 ( .A1(n641), .A2(n734), .ZN(n642) );
  NOR2_X2 U492 ( .A1(n634), .A2(n734), .ZN(n636) );
  NOR2_X2 U493 ( .A1(n655), .A2(n734), .ZN(n657) );
  NAND2_X1 U494 ( .A1(n400), .A2(n399), .ZN(n563) );
  NAND2_X1 U495 ( .A1(n562), .A2(n402), .ZN(n401) );
  NAND2_X1 U496 ( .A1(n603), .A2(n602), .ZN(n412) );
  NAND2_X1 U497 ( .A1(n403), .A2(n618), .ZN(n406) );
  NAND2_X1 U498 ( .A1(n619), .A2(n617), .ZN(n403) );
  NAND2_X1 U499 ( .A1(n637), .A2(KEYINPUT44), .ZN(n405) );
  NAND2_X1 U500 ( .A1(n406), .A2(n620), .ZN(n414) );
  NAND2_X1 U501 ( .A1(n408), .A2(n407), .ZN(n413) );
  NAND2_X1 U502 ( .A1(n637), .A2(n410), .ZN(n409) );
  AND2_X1 U503 ( .A1(n604), .A2(KEYINPUT44), .ZN(n410) );
  NAND2_X1 U504 ( .A1(n412), .A2(n604), .ZN(n411) );
  NAND2_X1 U505 ( .A1(n417), .A2(KEYINPUT2), .ZN(n416) );
  INV_X1 U506 ( .A(KEYINPUT2), .ZN(n421) );
  XNOR2_X2 U507 ( .A(n424), .B(n423), .ZN(n695) );
  INV_X1 U508 ( .A(KEYINPUT66), .ZN(n423) );
  NAND2_X1 U509 ( .A1(n524), .A2(n691), .ZN(n424) );
  NAND2_X1 U510 ( .A1(n644), .A2(n498), .ZN(n426) );
  XNOR2_X2 U511 ( .A(KEYINPUT110), .B(n544), .ZN(n762) );
  XOR2_X2 U512 ( .A(G119), .B(KEYINPUT3), .Z(n427) );
  XNOR2_X1 U513 ( .A(n442), .B(n366), .ZN(n443) );
  NOR2_X1 U514 ( .A1(n590), .A2(n610), .ZN(n577) );
  INV_X1 U515 ( .A(KEYINPUT112), .ZN(n519) );
  BUF_X1 U516 ( .A(n524), .Z(n605) );
  BUF_X1 U517 ( .A(n753), .Z(n754) );
  XNOR2_X1 U518 ( .A(n520), .B(n519), .ZN(n521) );
  XNOR2_X1 U519 ( .A(n448), .B(n447), .ZN(n523) );
  INV_X1 U520 ( .A(n671), .ZN(n675) );
  INV_X1 U521 ( .A(KEYINPUT63), .ZN(n635) );
  NAND2_X1 U522 ( .A1(G224), .A2(n756), .ZN(n432) );
  XNOR2_X2 U523 ( .A(G143), .B(G128), .ZN(n436) );
  NAND2_X1 U524 ( .A1(n652), .A2(n624), .ZN(n435) );
  XOR2_X1 U525 ( .A(KEYINPUT91), .B(KEYINPUT92), .Z(n434) );
  NAND2_X1 U526 ( .A1(G210), .A2(n449), .ZN(n433) );
  XNOR2_X2 U527 ( .A(n435), .B(n365), .ZN(n533) );
  INV_X1 U528 ( .A(n708), .ZN(n452) );
  XNOR2_X1 U529 ( .A(KEYINPUT67), .B(G137), .ZN(n437) );
  XNOR2_X1 U530 ( .A(n438), .B(n437), .ZN(n439) );
  XNOR2_X1 U531 ( .A(n440), .B(G131), .ZN(n441) );
  XNOR2_X1 U532 ( .A(n473), .B(n441), .ZN(n444) );
  NOR2_X1 U533 ( .A1(G953), .A2(G237), .ZN(n491) );
  XNOR2_X1 U534 ( .A(n446), .B(G146), .ZN(n470) );
  NAND2_X1 U535 ( .A1(n630), .A2(n498), .ZN(n448) );
  XOR2_X1 U536 ( .A(G472), .B(KEYINPUT100), .Z(n447) );
  NAND2_X1 U537 ( .A1(n449), .A2(G214), .ZN(n450) );
  XNOR2_X1 U538 ( .A(KEYINPUT93), .B(n450), .ZN(n709) );
  NOR2_X1 U539 ( .A1(n523), .A2(n709), .ZN(n451) );
  AND2_X1 U540 ( .A1(n452), .A2(n543), .ZN(n483) );
  NAND2_X1 U541 ( .A1(n756), .A2(G234), .ZN(n456) );
  XNOR2_X1 U542 ( .A(KEYINPUT79), .B(KEYINPUT8), .ZN(n455) );
  XNOR2_X1 U543 ( .A(n456), .B(n455), .ZN(n506) );
  XNOR2_X1 U544 ( .A(G128), .B(G119), .ZN(n457) );
  XNOR2_X1 U545 ( .A(n367), .B(n457), .ZN(n458) );
  XNOR2_X1 U546 ( .A(n459), .B(KEYINPUT24), .ZN(n460) );
  NOR2_X1 U547 ( .A1(n731), .A2(G902), .ZN(n465) );
  XOR2_X1 U548 ( .A(KEYINPUT25), .B(KEYINPUT97), .Z(n463) );
  NAND2_X1 U549 ( .A1(n624), .A2(G234), .ZN(n461) );
  XNOR2_X1 U550 ( .A(n461), .B(KEYINPUT20), .ZN(n466) );
  NAND2_X1 U551 ( .A1(n466), .A2(G217), .ZN(n462) );
  XNOR2_X1 U552 ( .A(n463), .B(n462), .ZN(n464) );
  XNOR2_X1 U553 ( .A(n465), .B(n464), .ZN(n524) );
  NAND2_X1 U554 ( .A1(G221), .A2(n466), .ZN(n467) );
  XOR2_X1 U555 ( .A(KEYINPUT21), .B(n467), .Z(n691) );
  NAND2_X1 U556 ( .A1(n756), .A2(G227), .ZN(n468) );
  XNOR2_X1 U557 ( .A(n468), .B(KEYINPUT73), .ZN(n469) );
  XNOR2_X1 U558 ( .A(n470), .B(n469), .ZN(n471) );
  XNOR2_X1 U559 ( .A(n472), .B(n471), .ZN(n474) );
  XNOR2_X1 U560 ( .A(G140), .B(G131), .ZN(n486) );
  XNOR2_X1 U561 ( .A(n473), .B(n486), .ZN(n747) );
  XNOR2_X1 U562 ( .A(n474), .B(n747), .ZN(n644) );
  INV_X1 U563 ( .A(G469), .ZN(n475) );
  INV_X1 U564 ( .A(n540), .ZN(n529) );
  NAND2_X1 U565 ( .A1(n695), .A2(n529), .ZN(n593) );
  NAND2_X1 U566 ( .A1(G234), .A2(G237), .ZN(n476) );
  XNOR2_X1 U567 ( .A(n476), .B(KEYINPUT14), .ZN(n478) );
  NAND2_X1 U568 ( .A1(G952), .A2(n478), .ZN(n722) );
  NOR2_X1 U569 ( .A1(G953), .A2(n722), .ZN(n477) );
  XNOR2_X1 U570 ( .A(KEYINPUT94), .B(n477), .ZN(n582) );
  INV_X1 U571 ( .A(n582), .ZN(n481) );
  NAND2_X1 U572 ( .A1(G902), .A2(n478), .ZN(n578) );
  NOR2_X1 U573 ( .A1(G900), .A2(n578), .ZN(n479) );
  NAND2_X1 U574 ( .A1(G953), .A2(n479), .ZN(n480) );
  NAND2_X1 U575 ( .A1(n481), .A2(n480), .ZN(n525) );
  INV_X1 U576 ( .A(n525), .ZN(n482) );
  AND2_X1 U577 ( .A1(n483), .A2(n542), .ZN(n484) );
  XNOR2_X1 U578 ( .A(n484), .B(KEYINPUT39), .ZN(n564) );
  XNOR2_X1 U579 ( .A(KEYINPUT12), .B(n486), .ZN(n487) );
  XOR2_X1 U580 ( .A(KEYINPUT102), .B(KEYINPUT11), .Z(n490) );
  XNOR2_X1 U581 ( .A(n490), .B(n489), .ZN(n495) );
  XOR2_X1 U582 ( .A(G104), .B(KEYINPUT103), .Z(n493) );
  NAND2_X1 U583 ( .A1(G214), .A2(n491), .ZN(n492) );
  XNOR2_X1 U584 ( .A(n493), .B(n492), .ZN(n494) );
  XOR2_X1 U585 ( .A(n495), .B(n494), .Z(n496) );
  XNOR2_X1 U586 ( .A(n497), .B(n496), .ZN(n638) );
  NAND2_X1 U587 ( .A1(n638), .A2(n498), .ZN(n500) );
  XOR2_X1 U588 ( .A(KEYINPUT13), .B(G475), .Z(n499) );
  XNOR2_X1 U589 ( .A(n500), .B(n499), .ZN(n548) );
  XNOR2_X1 U590 ( .A(n502), .B(n501), .ZN(n503) );
  XOR2_X1 U591 ( .A(n503), .B(KEYINPUT105), .Z(n505) );
  XNOR2_X1 U592 ( .A(n505), .B(n504), .ZN(n510) );
  NAND2_X1 U593 ( .A1(G217), .A2(n506), .ZN(n507) );
  XOR2_X1 U594 ( .A(n508), .B(n507), .Z(n509) );
  XNOR2_X1 U595 ( .A(n510), .B(n509), .ZN(n728) );
  NOR2_X1 U596 ( .A1(G902), .A2(n728), .ZN(n511) );
  XNOR2_X1 U597 ( .A(n511), .B(KEYINPUT106), .ZN(n513) );
  INV_X1 U598 ( .A(G478), .ZN(n512) );
  XNOR2_X1 U599 ( .A(n513), .B(n512), .ZN(n550) );
  INV_X1 U600 ( .A(n550), .ZN(n514) );
  NAND2_X1 U601 ( .A1(n548), .A2(n514), .ZN(n515) );
  NOR2_X1 U602 ( .A1(n564), .A2(n675), .ZN(n516) );
  INV_X1 U603 ( .A(KEYINPUT111), .ZN(n517) );
  XNOR2_X1 U604 ( .A(n518), .B(n517), .ZN(n713) );
  NOR2_X1 U605 ( .A1(n548), .A2(n550), .ZN(n711) );
  NAND2_X1 U606 ( .A1(n713), .A2(n711), .ZN(n522) );
  XOR2_X1 U607 ( .A(KEYINPUT113), .B(KEYINPUT41), .Z(n520) );
  NAND2_X1 U608 ( .A1(n525), .A2(n691), .ZN(n526) );
  NOR2_X1 U609 ( .A1(n524), .A2(n526), .ZN(n527) );
  XOR2_X1 U610 ( .A(KEYINPUT68), .B(n527), .Z(n536) );
  NOR2_X1 U611 ( .A1(n699), .A2(n536), .ZN(n528) );
  XNOR2_X1 U612 ( .A(n528), .B(KEYINPUT28), .ZN(n530) );
  NAND2_X1 U613 ( .A1(n530), .A2(n529), .ZN(n553) );
  NOR2_X1 U614 ( .A1(n706), .A2(n553), .ZN(n531) );
  XNOR2_X1 U615 ( .A(n531), .B(KEYINPUT42), .ZN(n764) );
  INV_X1 U616 ( .A(n709), .ZN(n565) );
  NAND2_X1 U617 ( .A1(n533), .A2(n565), .ZN(n534) );
  INV_X1 U618 ( .A(KEYINPUT6), .ZN(n535) );
  XNOR2_X1 U619 ( .A(n699), .B(n535), .ZN(n610) );
  NOR2_X1 U620 ( .A1(n536), .A2(n610), .ZN(n537) );
  NAND2_X1 U621 ( .A1(n671), .A2(n537), .ZN(n567) );
  NOR2_X1 U622 ( .A1(n552), .A2(n567), .ZN(n539) );
  XNOR2_X1 U623 ( .A(KEYINPUT85), .B(KEYINPUT36), .ZN(n538) );
  XNOR2_X1 U624 ( .A(n539), .B(n538), .ZN(n541) );
  XOR2_X1 U625 ( .A(KEYINPUT89), .B(n694), .Z(n611) );
  NOR2_X1 U626 ( .A1(n541), .A2(n611), .ZN(n680) );
  AND2_X1 U627 ( .A1(n550), .A2(n548), .ZN(n587) );
  INV_X1 U628 ( .A(n533), .ZN(n569) );
  XNOR2_X1 U629 ( .A(KEYINPUT78), .B(n762), .ZN(n546) );
  INV_X1 U630 ( .A(KEYINPUT77), .ZN(n559) );
  OR2_X1 U631 ( .A1(n559), .A2(KEYINPUT47), .ZN(n545) );
  NAND2_X1 U632 ( .A1(n546), .A2(n545), .ZN(n547) );
  INV_X1 U633 ( .A(n548), .ZN(n549) );
  NAND2_X1 U634 ( .A1(n550), .A2(n549), .ZN(n678) );
  NAND2_X1 U635 ( .A1(n675), .A2(n678), .ZN(n712) );
  INV_X1 U636 ( .A(n712), .ZN(n558) );
  XNOR2_X1 U637 ( .A(n552), .B(n551), .ZN(n584) );
  NOR2_X1 U638 ( .A1(n553), .A2(n584), .ZN(n554) );
  XNOR2_X1 U639 ( .A(n554), .B(KEYINPUT75), .ZN(n668) );
  NOR2_X1 U640 ( .A1(KEYINPUT47), .A2(n668), .ZN(n555) );
  NOR2_X1 U641 ( .A1(n555), .A2(KEYINPUT77), .ZN(n556) );
  NOR2_X1 U642 ( .A1(n558), .A2(n556), .ZN(n557) );
  NAND2_X1 U643 ( .A1(n559), .A2(n558), .ZN(n560) );
  INV_X1 U644 ( .A(n668), .ZN(n672) );
  NAND2_X1 U645 ( .A1(n560), .A2(n672), .ZN(n561) );
  NAND2_X1 U646 ( .A1(n561), .A2(KEYINPUT47), .ZN(n562) );
  XNOR2_X1 U647 ( .A(n563), .B(n371), .ZN(n573) );
  NOR2_X1 U648 ( .A1(n678), .A2(n564), .ZN(n682) );
  NAND2_X1 U649 ( .A1(n694), .A2(n565), .ZN(n566) );
  OR2_X1 U650 ( .A1(n567), .A2(n566), .ZN(n568) );
  XNOR2_X1 U651 ( .A(n568), .B(KEYINPUT43), .ZN(n570) );
  NAND2_X1 U652 ( .A1(n570), .A2(n569), .ZN(n684) );
  INV_X1 U653 ( .A(n684), .ZN(n571) );
  NOR2_X1 U654 ( .A1(n682), .A2(n571), .ZN(n572) );
  NAND2_X1 U655 ( .A1(n573), .A2(n572), .ZN(n625) );
  INV_X1 U656 ( .A(KEYINPUT81), .ZN(n574) );
  XNOR2_X1 U657 ( .A(n625), .B(n574), .ZN(n753) );
  XNOR2_X1 U658 ( .A(n575), .B(KEYINPUT71), .ZN(n590) );
  INV_X1 U659 ( .A(KEYINPUT109), .ZN(n576) );
  INV_X1 U660 ( .A(n578), .ZN(n579) );
  NOR2_X1 U661 ( .A1(G898), .A2(n756), .ZN(n744) );
  NAND2_X1 U662 ( .A1(n579), .A2(n744), .ZN(n580) );
  XNOR2_X1 U663 ( .A(KEYINPUT95), .B(n580), .ZN(n581) );
  NOR2_X1 U664 ( .A1(n582), .A2(n581), .ZN(n583) );
  NAND2_X1 U665 ( .A1(n599), .A2(n717), .ZN(n586) );
  XNOR2_X2 U666 ( .A(n589), .B(KEYINPUT35), .ZN(n637) );
  NOR2_X1 U667 ( .A1(n590), .A2(n699), .ZN(n591) );
  XNOR2_X1 U668 ( .A(n591), .B(KEYINPUT101), .ZN(n701) );
  INV_X1 U669 ( .A(n599), .ZN(n594) );
  NOR2_X1 U670 ( .A1(n701), .A2(n594), .ZN(n592) );
  XNOR2_X1 U671 ( .A(n592), .B(KEYINPUT31), .ZN(n677) );
  NOR2_X2 U672 ( .A1(n594), .A2(n593), .ZN(n595) );
  XNOR2_X1 U673 ( .A(KEYINPUT98), .B(n595), .ZN(n596) );
  NAND2_X1 U674 ( .A1(n596), .A2(n699), .ZN(n664) );
  NAND2_X1 U675 ( .A1(n677), .A2(n664), .ZN(n597) );
  NAND2_X1 U676 ( .A1(n597), .A2(n712), .ZN(n603) );
  AND2_X1 U677 ( .A1(n711), .A2(n691), .ZN(n598) );
  XNOR2_X1 U678 ( .A(n605), .B(KEYINPUT108), .ZN(n692) );
  AND2_X1 U679 ( .A1(n692), .A2(n694), .ZN(n600) );
  NAND2_X1 U680 ( .A1(n610), .A2(n600), .ZN(n601) );
  NOR2_X1 U681 ( .A1(n615), .A2(n601), .ZN(n658) );
  INV_X1 U682 ( .A(n658), .ZN(n602) );
  INV_X1 U683 ( .A(KEYINPUT84), .ZN(n604) );
  INV_X1 U684 ( .A(n637), .ZN(n617) );
  INV_X1 U685 ( .A(n605), .ZN(n606) );
  AND2_X1 U686 ( .A1(n606), .A2(n699), .ZN(n607) );
  NAND2_X1 U687 ( .A1(n607), .A2(n694), .ZN(n608) );
  NOR2_X1 U688 ( .A1(n615), .A2(n608), .ZN(n667) );
  INV_X1 U689 ( .A(n692), .ZN(n609) );
  NAND2_X1 U690 ( .A1(n610), .A2(n609), .ZN(n612) );
  NOR2_X1 U691 ( .A1(n612), .A2(n611), .ZN(n613) );
  XOR2_X1 U692 ( .A(KEYINPUT74), .B(n613), .Z(n614) );
  NOR2_X1 U693 ( .A1(n615), .A2(n614), .ZN(n616) );
  XNOR2_X1 U694 ( .A(n616), .B(KEYINPUT32), .ZN(n761) );
  INV_X1 U695 ( .A(KEYINPUT44), .ZN(n618) );
  NAND2_X1 U696 ( .A1(n619), .A2(KEYINPUT44), .ZN(n620) );
  INV_X1 U697 ( .A(KEYINPUT45), .ZN(n621) );
  INV_X1 U698 ( .A(KEYINPUT80), .ZN(n623) );
  INV_X1 U699 ( .A(n625), .ZN(n626) );
  NAND2_X1 U700 ( .A1(n626), .A2(KEYINPUT2), .ZN(n627) );
  NOR2_X1 U701 ( .A1(n735), .A2(n627), .ZN(n689) );
  NAND2_X1 U702 ( .A1(n648), .A2(G472), .ZN(n632) );
  XNOR2_X1 U703 ( .A(KEYINPUT114), .B(KEYINPUT115), .ZN(n628) );
  XNOR2_X1 U704 ( .A(n628), .B(KEYINPUT62), .ZN(n629) );
  XNOR2_X1 U705 ( .A(n630), .B(n629), .ZN(n631) );
  XNOR2_X1 U706 ( .A(n632), .B(n631), .ZN(n634) );
  INV_X1 U707 ( .A(G952), .ZN(n633) );
  AND2_X1 U708 ( .A1(n633), .A2(G953), .ZN(n734) );
  XNOR2_X1 U709 ( .A(n636), .B(n635), .ZN(G57) );
  XOR2_X1 U710 ( .A(n637), .B(G122), .Z(G24) );
  NAND2_X1 U711 ( .A1(n648), .A2(G475), .ZN(n640) );
  XNOR2_X1 U712 ( .A(n638), .B(KEYINPUT59), .ZN(n639) );
  XNOR2_X1 U713 ( .A(n640), .B(n639), .ZN(n641) );
  XNOR2_X1 U714 ( .A(n642), .B(KEYINPUT60), .ZN(G60) );
  NAND2_X1 U715 ( .A1(n648), .A2(G469), .ZN(n646) );
  XNOR2_X1 U716 ( .A(KEYINPUT57), .B(KEYINPUT58), .ZN(n643) );
  XNOR2_X1 U717 ( .A(n644), .B(n643), .ZN(n645) );
  XNOR2_X1 U718 ( .A(n646), .B(n645), .ZN(n647) );
  NOR2_X1 U719 ( .A1(n647), .A2(n734), .ZN(G54) );
  XOR2_X1 U720 ( .A(KEYINPUT87), .B(KEYINPUT54), .Z(n650) );
  XNOR2_X1 U721 ( .A(KEYINPUT55), .B(KEYINPUT76), .ZN(n649) );
  XNOR2_X1 U722 ( .A(n650), .B(n649), .ZN(n651) );
  XNOR2_X1 U723 ( .A(n652), .B(n651), .ZN(n653) );
  XNOR2_X1 U724 ( .A(n654), .B(n653), .ZN(n655) );
  XNOR2_X1 U725 ( .A(KEYINPUT82), .B(KEYINPUT56), .ZN(n656) );
  XNOR2_X1 U726 ( .A(n657), .B(n656), .ZN(G51) );
  XOR2_X1 U727 ( .A(G101), .B(n658), .Z(n659) );
  XNOR2_X1 U728 ( .A(KEYINPUT116), .B(n659), .ZN(G3) );
  NOR2_X1 U729 ( .A1(n675), .A2(n664), .ZN(n661) );
  XNOR2_X1 U730 ( .A(G104), .B(KEYINPUT117), .ZN(n660) );
  XNOR2_X1 U731 ( .A(n661), .B(n660), .ZN(G6) );
  XOR2_X1 U732 ( .A(KEYINPUT118), .B(KEYINPUT26), .Z(n663) );
  XNOR2_X1 U733 ( .A(G107), .B(KEYINPUT27), .ZN(n662) );
  XNOR2_X1 U734 ( .A(n663), .B(n662), .ZN(n666) );
  NOR2_X1 U735 ( .A1(n678), .A2(n664), .ZN(n665) );
  XOR2_X1 U736 ( .A(n666), .B(n665), .Z(G9) );
  XOR2_X1 U737 ( .A(G110), .B(n667), .Z(G12) );
  XOR2_X1 U738 ( .A(G128), .B(KEYINPUT29), .Z(n670) );
  OR2_X1 U739 ( .A1(n668), .A2(n678), .ZN(n669) );
  XNOR2_X1 U740 ( .A(n670), .B(n669), .ZN(G30) );
  XOR2_X1 U741 ( .A(G146), .B(KEYINPUT119), .Z(n674) );
  NAND2_X1 U742 ( .A1(n672), .A2(n671), .ZN(n673) );
  XNOR2_X1 U743 ( .A(n674), .B(n673), .ZN(G48) );
  NOR2_X1 U744 ( .A1(n675), .A2(n677), .ZN(n676) );
  XOR2_X1 U745 ( .A(G113), .B(n676), .Z(G15) );
  NOR2_X1 U746 ( .A1(n678), .A2(n677), .ZN(n679) );
  XOR2_X1 U747 ( .A(G116), .B(n679), .Z(G18) );
  XNOR2_X1 U748 ( .A(G125), .B(n680), .ZN(n681) );
  XNOR2_X1 U749 ( .A(n681), .B(KEYINPUT37), .ZN(G27) );
  XOR2_X1 U750 ( .A(G134), .B(n682), .Z(n683) );
  XNOR2_X1 U751 ( .A(KEYINPUT120), .B(n683), .ZN(G36) );
  XNOR2_X1 U752 ( .A(G140), .B(n684), .ZN(G42) );
  INV_X1 U753 ( .A(n706), .ZN(n685) );
  NAND2_X1 U754 ( .A1(n685), .A2(n717), .ZN(n686) );
  AND2_X1 U755 ( .A1(n686), .A2(n756), .ZN(n726) );
  INV_X1 U756 ( .A(n687), .ZN(n688) );
  NOR2_X1 U757 ( .A1(n688), .A2(KEYINPUT2), .ZN(n690) );
  NOR2_X1 U758 ( .A1(n690), .A2(n689), .ZN(n724) );
  OR2_X1 U759 ( .A1(n692), .A2(n691), .ZN(n693) );
  XNOR2_X1 U760 ( .A(n693), .B(KEYINPUT49), .ZN(n698) );
  NOR2_X1 U761 ( .A1(n695), .A2(n425), .ZN(n696) );
  XNOR2_X1 U762 ( .A(n696), .B(KEYINPUT50), .ZN(n697) );
  NOR2_X1 U763 ( .A1(n698), .A2(n697), .ZN(n700) );
  NAND2_X1 U764 ( .A1(n700), .A2(n699), .ZN(n702) );
  NAND2_X1 U765 ( .A1(n702), .A2(n701), .ZN(n703) );
  XNOR2_X1 U766 ( .A(n703), .B(KEYINPUT51), .ZN(n704) );
  XOR2_X1 U767 ( .A(KEYINPUT121), .B(n704), .Z(n705) );
  NOR2_X1 U768 ( .A1(n706), .A2(n705), .ZN(n707) );
  XOR2_X1 U769 ( .A(KEYINPUT122), .B(n707), .Z(n719) );
  NAND2_X1 U770 ( .A1(n709), .A2(n708), .ZN(n710) );
  NAND2_X1 U771 ( .A1(n711), .A2(n710), .ZN(n715) );
  NAND2_X1 U772 ( .A1(n713), .A2(n712), .ZN(n714) );
  NAND2_X1 U773 ( .A1(n715), .A2(n714), .ZN(n716) );
  NAND2_X1 U774 ( .A1(n717), .A2(n716), .ZN(n718) );
  NAND2_X1 U775 ( .A1(n719), .A2(n718), .ZN(n720) );
  XOR2_X1 U776 ( .A(KEYINPUT52), .B(n720), .Z(n721) );
  NOR2_X1 U777 ( .A1(n722), .A2(n721), .ZN(n723) );
  NOR2_X1 U778 ( .A1(n724), .A2(n723), .ZN(n725) );
  NAND2_X1 U779 ( .A1(n726), .A2(n725), .ZN(n727) );
  XOR2_X1 U780 ( .A(KEYINPUT53), .B(n727), .Z(G75) );
  NAND2_X1 U781 ( .A1(n648), .A2(G478), .ZN(n729) );
  XNOR2_X1 U782 ( .A(n729), .B(n728), .ZN(n730) );
  NOR2_X1 U783 ( .A1(n734), .A2(n730), .ZN(G63) );
  NAND2_X1 U784 ( .A1(n648), .A2(G217), .ZN(n732) );
  XNOR2_X1 U785 ( .A(n732), .B(n731), .ZN(n733) );
  NOR2_X1 U786 ( .A1(n734), .A2(n733), .ZN(G66) );
  NAND2_X1 U787 ( .A1(n383), .A2(n756), .ZN(n739) );
  NAND2_X1 U788 ( .A1(G953), .A2(G224), .ZN(n736) );
  XNOR2_X1 U789 ( .A(KEYINPUT61), .B(n736), .ZN(n737) );
  NAND2_X1 U790 ( .A1(n737), .A2(G898), .ZN(n738) );
  NAND2_X1 U791 ( .A1(n739), .A2(n738), .ZN(n746) );
  XNOR2_X1 U792 ( .A(G101), .B(n740), .ZN(n742) );
  XNOR2_X1 U793 ( .A(n742), .B(n741), .ZN(n743) );
  NOR2_X1 U794 ( .A1(n744), .A2(n743), .ZN(n745) );
  XNOR2_X1 U795 ( .A(n746), .B(n745), .ZN(G69) );
  XOR2_X1 U796 ( .A(n485), .B(KEYINPUT123), .Z(n748) );
  XNOR2_X1 U797 ( .A(n748), .B(n747), .ZN(n755) );
  XNOR2_X1 U798 ( .A(G227), .B(n755), .ZN(n749) );
  NAND2_X1 U799 ( .A1(n749), .A2(G900), .ZN(n750) );
  XOR2_X1 U800 ( .A(KEYINPUT124), .B(n750), .Z(n751) );
  NOR2_X1 U801 ( .A1(n756), .A2(n751), .ZN(n752) );
  XNOR2_X1 U802 ( .A(KEYINPUT125), .B(n752), .ZN(n759) );
  XNOR2_X1 U803 ( .A(n755), .B(n754), .ZN(n757) );
  NAND2_X1 U804 ( .A1(n757), .A2(n756), .ZN(n758) );
  NAND2_X1 U805 ( .A1(n759), .A2(n758), .ZN(n760) );
  XNOR2_X1 U806 ( .A(n760), .B(KEYINPUT126), .ZN(G72) );
  XOR2_X1 U807 ( .A(G119), .B(n761), .Z(G21) );
  XNOR2_X1 U808 ( .A(G143), .B(n762), .ZN(G45) );
  XOR2_X1 U809 ( .A(G131), .B(n763), .Z(G33) );
  XNOR2_X1 U810 ( .A(G137), .B(KEYINPUT127), .ZN(n765) );
  XNOR2_X1 U811 ( .A(n765), .B(n764), .ZN(G39) );
endmodule

