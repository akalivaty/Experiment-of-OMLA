//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 1 1 0 0 0 0 1 0 1 1 1 1 1 0 0 1 0 0 1 1 1 1 0 0 0 0 1 0 1 0 0 0 1 0 0 1 1 0 0 1 1 0 0 1 0 0 0 1 0 1 1 0 1 0 0 1 0 0 1 0 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:37:53 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1247, new_n1248,
    new_n1249, new_n1250, new_n1251, new_n1253, new_n1254, new_n1255,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1312, new_n1313;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(new_n201), .ZN(new_n202));
  NOR2_X1   g0002(.A1(new_n202), .A2(G50), .ZN(new_n203));
  INV_X1    g0003(.A(new_n203), .ZN(new_n204));
  NOR2_X1   g0004(.A1(new_n204), .A2(G77), .ZN(G353));
  OAI21_X1  g0005(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0006(.A(G1), .ZN(new_n207));
  INV_X1    g0007(.A(G20), .ZN(new_n208));
  NOR2_X1   g0008(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  INV_X1    g0009(.A(new_n209), .ZN(new_n210));
  NOR2_X1   g0010(.A1(new_n210), .A2(G13), .ZN(new_n211));
  OAI211_X1 g0011(.A(new_n211), .B(G250), .C1(G257), .C2(G264), .ZN(new_n212));
  INV_X1    g0012(.A(KEYINPUT0), .ZN(new_n213));
  NAND2_X1  g0013(.A1(G1), .A2(G13), .ZN(new_n214));
  NOR2_X1   g0014(.A1(new_n214), .A2(new_n208), .ZN(new_n215));
  NAND2_X1  g0015(.A1(new_n202), .A2(G50), .ZN(new_n216));
  INV_X1    g0016(.A(new_n216), .ZN(new_n217));
  AOI22_X1  g0017(.A1(new_n212), .A2(new_n213), .B1(new_n215), .B2(new_n217), .ZN(new_n218));
  XNOR2_X1  g0018(.A(KEYINPUT64), .B(G238), .ZN(new_n219));
  INV_X1    g0019(.A(G68), .ZN(new_n220));
  NOR2_X1   g0020(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  AOI22_X1  g0021(.A1(G58), .A2(G232), .B1(G87), .B2(G250), .ZN(new_n222));
  AOI22_X1  g0022(.A1(G77), .A2(G244), .B1(G116), .B2(G270), .ZN(new_n223));
  AOI22_X1  g0023(.A1(G50), .A2(G226), .B1(G97), .B2(G257), .ZN(new_n224));
  NAND2_X1  g0024(.A1(G107), .A2(G264), .ZN(new_n225));
  NAND4_X1  g0025(.A1(new_n222), .A2(new_n223), .A3(new_n224), .A4(new_n225), .ZN(new_n226));
  OAI21_X1  g0026(.A(new_n210), .B1(new_n221), .B2(new_n226), .ZN(new_n227));
  OAI221_X1 g0027(.A(new_n218), .B1(new_n213), .B2(new_n212), .C1(new_n227), .C2(KEYINPUT1), .ZN(new_n228));
  AOI21_X1  g0028(.A(new_n228), .B1(KEYINPUT1), .B2(new_n227), .ZN(G361));
  XNOR2_X1  g0029(.A(G238), .B(G244), .ZN(new_n230));
  XNOR2_X1  g0030(.A(new_n230), .B(KEYINPUT2), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n231), .B(G226), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n232), .B(G232), .ZN(new_n233));
  XOR2_X1   g0033(.A(G250), .B(G257), .Z(new_n234));
  XNOR2_X1  g0034(.A(G264), .B(G270), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n233), .B(new_n236), .ZN(G358));
  XOR2_X1   g0037(.A(G68), .B(G77), .Z(new_n238));
  XNOR2_X1  g0038(.A(G50), .B(G58), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XOR2_X1   g0040(.A(G87), .B(G97), .Z(new_n241));
  XNOR2_X1  g0041(.A(G107), .B(G116), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n240), .B(new_n243), .ZN(G351));
  INV_X1    g0044(.A(G33), .ZN(new_n245));
  NOR2_X1   g0045(.A1(new_n245), .A2(KEYINPUT3), .ZN(new_n246));
  INV_X1    g0046(.A(KEYINPUT3), .ZN(new_n247));
  NOR2_X1   g0047(.A1(new_n247), .A2(G33), .ZN(new_n248));
  NOR2_X1   g0048(.A1(new_n246), .A2(new_n248), .ZN(new_n249));
  NAND3_X1  g0049(.A1(new_n249), .A2(G223), .A3(G1698), .ZN(new_n250));
  INV_X1    g0050(.A(G1698), .ZN(new_n251));
  NAND3_X1  g0051(.A1(new_n249), .A2(G222), .A3(new_n251), .ZN(new_n252));
  INV_X1    g0052(.A(G77), .ZN(new_n253));
  OAI211_X1 g0053(.A(new_n250), .B(new_n252), .C1(new_n253), .C2(new_n249), .ZN(new_n254));
  NAND2_X1  g0054(.A1(G33), .A2(G41), .ZN(new_n255));
  NAND3_X1  g0055(.A1(new_n255), .A2(G1), .A3(G13), .ZN(new_n256));
  INV_X1    g0056(.A(new_n256), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n254), .A2(new_n257), .ZN(new_n258));
  OAI21_X1  g0058(.A(new_n207), .B1(G41), .B2(G45), .ZN(new_n259));
  INV_X1    g0059(.A(G274), .ZN(new_n260));
  NOR2_X1   g0060(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n256), .A2(new_n259), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n262), .A2(KEYINPUT65), .ZN(new_n263));
  INV_X1    g0063(.A(KEYINPUT65), .ZN(new_n264));
  NAND3_X1  g0064(.A1(new_n256), .A2(new_n264), .A3(new_n259), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n263), .A2(new_n265), .ZN(new_n266));
  AOI21_X1  g0066(.A(new_n261), .B1(new_n266), .B2(G226), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n258), .A2(new_n267), .ZN(new_n268));
  INV_X1    g0068(.A(KEYINPUT66), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  NAND3_X1  g0070(.A1(new_n258), .A2(KEYINPUT66), .A3(new_n267), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  INV_X1    g0072(.A(G179), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  XOR2_X1   g0074(.A(new_n274), .B(KEYINPUT69), .Z(new_n275));
  NAND3_X1  g0075(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n276), .A2(new_n214), .ZN(new_n277));
  NAND3_X1  g0077(.A1(new_n204), .A2(KEYINPUT67), .A3(G20), .ZN(new_n278));
  INV_X1    g0078(.A(G150), .ZN(new_n279));
  NOR2_X1   g0079(.A1(G20), .A2(G33), .ZN(new_n280));
  INV_X1    g0080(.A(new_n280), .ZN(new_n281));
  XNOR2_X1  g0081(.A(KEYINPUT8), .B(G58), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n208), .A2(G33), .ZN(new_n283));
  OAI221_X1 g0083(.A(new_n278), .B1(new_n279), .B2(new_n281), .C1(new_n282), .C2(new_n283), .ZN(new_n284));
  AOI21_X1  g0084(.A(KEYINPUT67), .B1(new_n204), .B2(G20), .ZN(new_n285));
  OAI21_X1  g0085(.A(new_n277), .B1(new_n284), .B2(new_n285), .ZN(new_n286));
  NOR2_X1   g0086(.A1(new_n208), .A2(G1), .ZN(new_n287));
  XNOR2_X1  g0087(.A(new_n287), .B(KEYINPUT68), .ZN(new_n288));
  AND2_X1   g0088(.A1(new_n276), .A2(new_n214), .ZN(new_n289));
  INV_X1    g0089(.A(G13), .ZN(new_n290));
  NOR2_X1   g0090(.A1(new_n290), .A2(G1), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n291), .A2(G20), .ZN(new_n292));
  NAND3_X1  g0092(.A1(new_n288), .A2(new_n289), .A3(new_n292), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n293), .A2(G50), .ZN(new_n294));
  INV_X1    g0094(.A(new_n292), .ZN(new_n295));
  OAI21_X1  g0095(.A(new_n294), .B1(G50), .B2(new_n295), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n286), .A2(new_n296), .ZN(new_n297));
  OAI211_X1 g0097(.A(new_n275), .B(new_n297), .C1(G169), .C2(new_n272), .ZN(new_n298));
  NOR2_X1   g0098(.A1(KEYINPUT72), .A2(KEYINPUT10), .ZN(new_n299));
  XNOR2_X1  g0099(.A(new_n297), .B(KEYINPUT9), .ZN(new_n300));
  INV_X1    g0100(.A(G190), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n272), .A2(new_n301), .ZN(new_n302));
  OAI21_X1  g0102(.A(new_n302), .B1(G200), .B2(new_n272), .ZN(new_n303));
  AOI21_X1  g0103(.A(new_n299), .B1(new_n300), .B2(new_n303), .ZN(new_n304));
  NAND2_X1  g0104(.A1(KEYINPUT72), .A2(KEYINPUT10), .ZN(new_n305));
  OR2_X1    g0105(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n304), .A2(new_n305), .ZN(new_n307));
  NAND3_X1  g0107(.A1(new_n298), .A2(new_n306), .A3(new_n307), .ZN(new_n308));
  INV_X1    g0108(.A(new_n282), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n293), .A2(new_n309), .ZN(new_n310));
  OAI21_X1  g0110(.A(new_n310), .B1(new_n295), .B2(new_n309), .ZN(new_n311));
  NAND3_X1  g0111(.A1(new_n256), .A2(G232), .A3(new_n259), .ZN(new_n312));
  OR2_X1    g0112(.A1(new_n312), .A2(KEYINPUT79), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n312), .A2(KEYINPUT79), .ZN(new_n314));
  INV_X1    g0114(.A(new_n261), .ZN(new_n315));
  NAND3_X1  g0115(.A1(new_n313), .A2(new_n314), .A3(new_n315), .ZN(new_n316));
  INV_X1    g0116(.A(KEYINPUT76), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n317), .A2(new_n245), .ZN(new_n318));
  NAND2_X1  g0118(.A1(KEYINPUT76), .A2(G33), .ZN(new_n319));
  NAND3_X1  g0119(.A1(new_n318), .A2(KEYINPUT3), .A3(new_n319), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n247), .A2(G33), .ZN(new_n321));
  AND2_X1   g0121(.A1(G226), .A2(G1698), .ZN(new_n322));
  NAND3_X1  g0122(.A1(new_n320), .A2(new_n321), .A3(new_n322), .ZN(new_n323));
  NAND2_X1  g0123(.A1(G33), .A2(G87), .ZN(new_n324));
  AND2_X1   g0124(.A1(new_n323), .A2(new_n324), .ZN(new_n325));
  AND2_X1   g0125(.A1(KEYINPUT76), .A2(G33), .ZN(new_n326));
  NOR2_X1   g0126(.A1(KEYINPUT76), .A2(G33), .ZN(new_n327));
  NOR2_X1   g0127(.A1(new_n326), .A2(new_n327), .ZN(new_n328));
  AOI21_X1  g0128(.A(new_n246), .B1(new_n328), .B2(KEYINPUT3), .ZN(new_n329));
  NAND4_X1  g0129(.A1(new_n329), .A2(KEYINPUT78), .A3(G223), .A4(new_n251), .ZN(new_n330));
  NAND4_X1  g0130(.A1(new_n320), .A2(G223), .A3(new_n251), .A4(new_n321), .ZN(new_n331));
  INV_X1    g0131(.A(KEYINPUT78), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n331), .A2(new_n332), .ZN(new_n333));
  NAND3_X1  g0133(.A1(new_n325), .A2(new_n330), .A3(new_n333), .ZN(new_n334));
  AOI211_X1 g0134(.A(G190), .B(new_n316), .C1(new_n334), .C2(new_n257), .ZN(new_n335));
  OAI211_X1 g0135(.A(new_n324), .B(new_n323), .C1(new_n331), .C2(new_n332), .ZN(new_n336));
  AND2_X1   g0136(.A1(new_n331), .A2(new_n332), .ZN(new_n337));
  OAI21_X1  g0137(.A(new_n257), .B1(new_n336), .B2(new_n337), .ZN(new_n338));
  INV_X1    g0138(.A(new_n316), .ZN(new_n339));
  AOI21_X1  g0139(.A(G200), .B1(new_n338), .B2(new_n339), .ZN(new_n340));
  OAI21_X1  g0140(.A(new_n311), .B1(new_n335), .B2(new_n340), .ZN(new_n341));
  INV_X1    g0141(.A(KEYINPUT77), .ZN(new_n342));
  INV_X1    g0142(.A(KEYINPUT7), .ZN(new_n343));
  NOR3_X1   g0143(.A1(new_n326), .A2(new_n327), .A3(new_n247), .ZN(new_n344));
  OAI211_X1 g0144(.A(new_n343), .B(new_n208), .C1(new_n344), .C2(new_n246), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n345), .A2(G68), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n320), .A2(new_n321), .ZN(new_n347));
  AOI21_X1  g0147(.A(new_n343), .B1(new_n347), .B2(new_n208), .ZN(new_n348));
  OAI21_X1  g0148(.A(new_n342), .B1(new_n346), .B2(new_n348), .ZN(new_n349));
  NAND2_X1  g0149(.A1(G58), .A2(G68), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n202), .A2(new_n350), .ZN(new_n351));
  AOI22_X1  g0151(.A1(new_n351), .A2(G20), .B1(G159), .B2(new_n280), .ZN(new_n352));
  OAI21_X1  g0152(.A(KEYINPUT7), .B1(new_n329), .B2(G20), .ZN(new_n353));
  NAND4_X1  g0153(.A1(new_n353), .A2(KEYINPUT77), .A3(G68), .A4(new_n345), .ZN(new_n354));
  NAND4_X1  g0154(.A1(new_n349), .A2(KEYINPUT16), .A3(new_n352), .A4(new_n354), .ZN(new_n355));
  INV_X1    g0155(.A(KEYINPUT16), .ZN(new_n356));
  AOI21_X1  g0156(.A(KEYINPUT3), .B1(new_n318), .B2(new_n319), .ZN(new_n357));
  OAI211_X1 g0157(.A(KEYINPUT7), .B(new_n208), .C1(new_n357), .C2(new_n248), .ZN(new_n358));
  OAI21_X1  g0158(.A(new_n343), .B1(new_n249), .B2(G20), .ZN(new_n359));
  AOI21_X1  g0159(.A(new_n220), .B1(new_n358), .B2(new_n359), .ZN(new_n360));
  INV_X1    g0160(.A(new_n352), .ZN(new_n361));
  OAI21_X1  g0161(.A(new_n356), .B1(new_n360), .B2(new_n361), .ZN(new_n362));
  AND3_X1   g0162(.A1(new_n355), .A2(new_n362), .A3(new_n277), .ZN(new_n363));
  OAI21_X1  g0163(.A(KEYINPUT80), .B1(new_n341), .B2(new_n363), .ZN(new_n364));
  NAND3_X1  g0164(.A1(new_n338), .A2(new_n301), .A3(new_n339), .ZN(new_n365));
  AOI21_X1  g0165(.A(new_n316), .B1(new_n334), .B2(new_n257), .ZN(new_n366));
  OAI21_X1  g0166(.A(new_n365), .B1(G200), .B2(new_n366), .ZN(new_n367));
  NAND3_X1  g0167(.A1(new_n355), .A2(new_n362), .A3(new_n277), .ZN(new_n368));
  INV_X1    g0168(.A(KEYINPUT80), .ZN(new_n369));
  NAND4_X1  g0169(.A1(new_n367), .A2(new_n368), .A3(new_n369), .A4(new_n311), .ZN(new_n370));
  NAND3_X1  g0170(.A1(new_n364), .A2(KEYINPUT17), .A3(new_n370), .ZN(new_n371));
  NAND3_X1  g0171(.A1(new_n367), .A2(new_n368), .A3(new_n311), .ZN(new_n372));
  OR2_X1    g0172(.A1(new_n372), .A2(KEYINPUT17), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n371), .A2(new_n373), .ZN(new_n374));
  NAND3_X1  g0174(.A1(new_n338), .A2(new_n273), .A3(new_n339), .ZN(new_n375));
  OAI21_X1  g0175(.A(new_n375), .B1(G169), .B2(new_n366), .ZN(new_n376));
  AOI21_X1  g0176(.A(new_n376), .B1(new_n368), .B2(new_n311), .ZN(new_n377));
  XNOR2_X1  g0177(.A(new_n377), .B(KEYINPUT18), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n374), .A2(new_n378), .ZN(new_n379));
  NAND3_X1  g0179(.A1(new_n291), .A2(G20), .A3(new_n220), .ZN(new_n380));
  XNOR2_X1  g0180(.A(new_n380), .B(KEYINPUT12), .ZN(new_n381));
  AOI22_X1  g0181(.A1(new_n280), .A2(G50), .B1(G20), .B2(new_n220), .ZN(new_n382));
  OAI21_X1  g0182(.A(new_n382), .B1(new_n253), .B2(new_n283), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n383), .A2(new_n277), .ZN(new_n384));
  INV_X1    g0184(.A(new_n384), .ZN(new_n385));
  OAI21_X1  g0185(.A(new_n381), .B1(new_n385), .B2(KEYINPUT11), .ZN(new_n386));
  INV_X1    g0186(.A(KEYINPUT11), .ZN(new_n387));
  OAI22_X1  g0187(.A1(new_n293), .A2(new_n220), .B1(new_n384), .B2(new_n387), .ZN(new_n388));
  NOR2_X1   g0188(.A1(new_n386), .A2(new_n388), .ZN(new_n389));
  AND3_X1   g0189(.A1(new_n256), .A2(new_n264), .A3(new_n259), .ZN(new_n390));
  AOI21_X1  g0190(.A(new_n264), .B1(new_n256), .B2(new_n259), .ZN(new_n391));
  NOR3_X1   g0191(.A1(new_n390), .A2(new_n391), .A3(KEYINPUT74), .ZN(new_n392));
  INV_X1    g0192(.A(KEYINPUT74), .ZN(new_n393));
  AOI21_X1  g0193(.A(new_n393), .B1(new_n263), .B2(new_n265), .ZN(new_n394));
  OAI21_X1  g0194(.A(G238), .B1(new_n392), .B2(new_n394), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n245), .A2(KEYINPUT3), .ZN(new_n396));
  NAND4_X1  g0196(.A1(new_n321), .A2(new_n396), .A3(G232), .A4(G1698), .ZN(new_n397));
  NAND4_X1  g0197(.A1(new_n321), .A2(new_n396), .A3(G226), .A4(new_n251), .ZN(new_n398));
  NAND2_X1  g0198(.A1(G33), .A2(G97), .ZN(new_n399));
  NAND3_X1  g0199(.A1(new_n397), .A2(new_n398), .A3(new_n399), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n400), .A2(KEYINPUT73), .ZN(new_n401));
  INV_X1    g0201(.A(KEYINPUT73), .ZN(new_n402));
  NAND4_X1  g0202(.A1(new_n397), .A2(new_n398), .A3(new_n402), .A4(new_n399), .ZN(new_n403));
  NAND3_X1  g0203(.A1(new_n401), .A2(new_n257), .A3(new_n403), .ZN(new_n404));
  NAND3_X1  g0204(.A1(new_n395), .A2(new_n315), .A3(new_n404), .ZN(new_n405));
  NOR2_X1   g0205(.A1(new_n405), .A2(KEYINPUT13), .ZN(new_n406));
  INV_X1    g0206(.A(KEYINPUT13), .ZN(new_n407));
  OAI21_X1  g0207(.A(KEYINPUT74), .B1(new_n390), .B2(new_n391), .ZN(new_n408));
  NAND3_X1  g0208(.A1(new_n263), .A2(new_n393), .A3(new_n265), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n408), .A2(new_n409), .ZN(new_n410));
  AOI21_X1  g0210(.A(new_n261), .B1(new_n410), .B2(G238), .ZN(new_n411));
  AOI21_X1  g0211(.A(new_n407), .B1(new_n411), .B2(new_n404), .ZN(new_n412));
  NOR3_X1   g0212(.A1(new_n406), .A2(new_n412), .A3(G190), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n405), .A2(KEYINPUT13), .ZN(new_n414));
  NAND3_X1  g0214(.A1(new_n411), .A2(new_n407), .A3(new_n404), .ZN(new_n415));
  AOI21_X1  g0215(.A(G200), .B1(new_n414), .B2(new_n415), .ZN(new_n416));
  OAI21_X1  g0216(.A(new_n389), .B1(new_n413), .B2(new_n416), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n417), .A2(KEYINPUT75), .ZN(new_n418));
  INV_X1    g0218(.A(G200), .ZN(new_n419));
  OAI21_X1  g0219(.A(new_n419), .B1(new_n406), .B2(new_n412), .ZN(new_n420));
  NAND3_X1  g0220(.A1(new_n414), .A2(new_n301), .A3(new_n415), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n420), .A2(new_n421), .ZN(new_n422));
  INV_X1    g0222(.A(KEYINPUT75), .ZN(new_n423));
  NAND3_X1  g0223(.A1(new_n422), .A2(new_n423), .A3(new_n389), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n418), .A2(new_n424), .ZN(new_n425));
  INV_X1    g0225(.A(new_n389), .ZN(new_n426));
  NAND3_X1  g0226(.A1(new_n414), .A2(G179), .A3(new_n415), .ZN(new_n427));
  INV_X1    g0227(.A(G169), .ZN(new_n428));
  AOI21_X1  g0228(.A(new_n428), .B1(new_n414), .B2(new_n415), .ZN(new_n429));
  INV_X1    g0229(.A(KEYINPUT14), .ZN(new_n430));
  OAI21_X1  g0230(.A(new_n427), .B1(new_n429), .B2(new_n430), .ZN(new_n431));
  AOI211_X1 g0231(.A(KEYINPUT14), .B(new_n428), .C1(new_n414), .C2(new_n415), .ZN(new_n432));
  OAI21_X1  g0232(.A(new_n426), .B1(new_n431), .B2(new_n432), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n425), .A2(new_n433), .ZN(new_n434));
  XNOR2_X1  g0234(.A(KEYINPUT15), .B(G87), .ZN(new_n435));
  OAI22_X1  g0235(.A1(new_n435), .A2(new_n283), .B1(new_n208), .B2(new_n253), .ZN(new_n436));
  NOR2_X1   g0236(.A1(new_n282), .A2(new_n281), .ZN(new_n437));
  OAI21_X1  g0237(.A(new_n277), .B1(new_n436), .B2(new_n437), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n295), .A2(new_n253), .ZN(new_n439));
  OAI211_X1 g0239(.A(new_n438), .B(new_n439), .C1(new_n293), .C2(new_n253), .ZN(new_n440));
  XNOR2_X1  g0240(.A(new_n440), .B(KEYINPUT71), .ZN(new_n441));
  INV_X1    g0241(.A(new_n441), .ZN(new_n442));
  NAND3_X1  g0242(.A1(new_n249), .A2(G232), .A3(new_n251), .ZN(new_n443));
  INV_X1    g0243(.A(G107), .ZN(new_n444));
  OAI21_X1  g0244(.A(new_n443), .B1(new_n444), .B2(new_n249), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n321), .A2(new_n396), .ZN(new_n446));
  NOR3_X1   g0246(.A1(new_n446), .A2(new_n219), .A3(new_n251), .ZN(new_n447));
  OAI21_X1  g0247(.A(new_n257), .B1(new_n445), .B2(new_n447), .ZN(new_n448));
  INV_X1    g0248(.A(KEYINPUT70), .ZN(new_n449));
  AOI21_X1  g0249(.A(new_n261), .B1(new_n266), .B2(G244), .ZN(new_n450));
  NAND3_X1  g0250(.A1(new_n448), .A2(new_n449), .A3(new_n450), .ZN(new_n451));
  INV_X1    g0251(.A(new_n451), .ZN(new_n452));
  AOI21_X1  g0252(.A(new_n449), .B1(new_n448), .B2(new_n450), .ZN(new_n453));
  OAI21_X1  g0253(.A(new_n301), .B1(new_n452), .B2(new_n453), .ZN(new_n454));
  INV_X1    g0254(.A(new_n453), .ZN(new_n455));
  NAND3_X1  g0255(.A1(new_n455), .A2(new_n419), .A3(new_n451), .ZN(new_n456));
  AOI21_X1  g0256(.A(new_n442), .B1(new_n454), .B2(new_n456), .ZN(new_n457));
  OAI21_X1  g0257(.A(G179), .B1(new_n452), .B2(new_n453), .ZN(new_n458));
  NAND3_X1  g0258(.A1(new_n455), .A2(G169), .A3(new_n451), .ZN(new_n459));
  AOI21_X1  g0259(.A(new_n441), .B1(new_n458), .B2(new_n459), .ZN(new_n460));
  NOR2_X1   g0260(.A1(new_n457), .A2(new_n460), .ZN(new_n461));
  INV_X1    g0261(.A(new_n461), .ZN(new_n462));
  NOR4_X1   g0262(.A1(new_n308), .A2(new_n379), .A3(new_n434), .A4(new_n462), .ZN(new_n463));
  INV_X1    g0263(.A(KEYINPUT6), .ZN(new_n464));
  INV_X1    g0264(.A(G97), .ZN(new_n465));
  NOR2_X1   g0265(.A1(new_n465), .A2(new_n444), .ZN(new_n466));
  NOR2_X1   g0266(.A1(G97), .A2(G107), .ZN(new_n467));
  OAI21_X1  g0267(.A(new_n464), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  NAND3_X1  g0268(.A1(new_n444), .A2(KEYINPUT6), .A3(G97), .ZN(new_n469));
  AND2_X1   g0269(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  OAI22_X1  g0270(.A1(new_n470), .A2(new_n208), .B1(new_n253), .B2(new_n281), .ZN(new_n471));
  AOI21_X1  g0271(.A(new_n444), .B1(new_n358), .B2(new_n359), .ZN(new_n472));
  OAI21_X1  g0272(.A(new_n277), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  OAI211_X1 g0273(.A(new_n289), .B(new_n292), .C1(G1), .C2(new_n245), .ZN(new_n474));
  MUX2_X1   g0274(.A(new_n292), .B(new_n474), .S(G97), .Z(new_n475));
  NAND2_X1  g0275(.A1(new_n473), .A2(new_n475), .ZN(new_n476));
  NAND4_X1  g0276(.A1(new_n320), .A2(G244), .A3(new_n251), .A4(new_n321), .ZN(new_n477));
  INV_X1    g0277(.A(KEYINPUT4), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  NAND4_X1  g0279(.A1(new_n321), .A2(new_n396), .A3(G250), .A4(G1698), .ZN(new_n480));
  AND2_X1   g0280(.A1(KEYINPUT4), .A2(G244), .ZN(new_n481));
  NAND4_X1  g0281(.A1(new_n321), .A2(new_n396), .A3(new_n481), .A4(new_n251), .ZN(new_n482));
  NAND2_X1  g0282(.A1(G33), .A2(G283), .ZN(new_n483));
  AND3_X1   g0283(.A1(new_n480), .A2(new_n482), .A3(new_n483), .ZN(new_n484));
  AOI21_X1  g0284(.A(new_n256), .B1(new_n479), .B2(new_n484), .ZN(new_n485));
  INV_X1    g0285(.A(G45), .ZN(new_n486));
  NOR2_X1   g0286(.A1(new_n486), .A2(G1), .ZN(new_n487));
  AND2_X1   g0287(.A1(KEYINPUT5), .A2(G41), .ZN(new_n488));
  NOR2_X1   g0288(.A1(KEYINPUT5), .A2(G41), .ZN(new_n489));
  OAI21_X1  g0289(.A(new_n487), .B1(new_n488), .B2(new_n489), .ZN(new_n490));
  OR2_X1    g0290(.A1(new_n490), .A2(new_n260), .ZN(new_n491));
  INV_X1    g0291(.A(G257), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n490), .A2(new_n256), .ZN(new_n493));
  OAI21_X1  g0293(.A(new_n491), .B1(new_n492), .B2(new_n493), .ZN(new_n494));
  OAI21_X1  g0294(.A(new_n419), .B1(new_n485), .B2(new_n494), .ZN(new_n495));
  INV_X1    g0295(.A(new_n494), .ZN(new_n496));
  AND2_X1   g0296(.A1(new_n479), .A2(new_n484), .ZN(new_n497));
  OAI211_X1 g0297(.A(new_n496), .B(new_n301), .C1(new_n497), .C2(new_n256), .ZN(new_n498));
  AOI21_X1  g0298(.A(new_n476), .B1(new_n495), .B2(new_n498), .ZN(new_n499));
  OAI211_X1 g0299(.A(new_n496), .B(G179), .C1(new_n497), .C2(new_n256), .ZN(new_n500));
  OAI21_X1  g0300(.A(G169), .B1(new_n485), .B2(new_n494), .ZN(new_n501));
  AOI22_X1  g0301(.A1(new_n500), .A2(new_n501), .B1(new_n473), .B2(new_n475), .ZN(new_n502));
  OAI21_X1  g0302(.A(KEYINPUT81), .B1(new_n499), .B2(new_n502), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n500), .A2(new_n501), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n504), .A2(new_n476), .ZN(new_n505));
  INV_X1    g0305(.A(KEYINPUT81), .ZN(new_n506));
  AND2_X1   g0306(.A1(new_n498), .A2(new_n495), .ZN(new_n507));
  OAI211_X1 g0307(.A(new_n505), .B(new_n506), .C1(new_n476), .C2(new_n507), .ZN(new_n508));
  AND2_X1   g0308(.A1(new_n503), .A2(new_n508), .ZN(new_n509));
  NAND3_X1  g0309(.A1(new_n291), .A2(G20), .A3(new_n444), .ZN(new_n510));
  OR2_X1    g0310(.A1(new_n510), .A2(KEYINPUT25), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n510), .A2(KEYINPUT25), .ZN(new_n512));
  OAI211_X1 g0312(.A(new_n511), .B(new_n512), .C1(new_n474), .C2(new_n444), .ZN(new_n513));
  INV_X1    g0313(.A(new_n513), .ZN(new_n514));
  INV_X1    g0314(.A(G87), .ZN(new_n515));
  OR4_X1    g0315(.A1(KEYINPUT22), .A2(new_n446), .A3(G20), .A4(new_n515), .ZN(new_n516));
  NAND3_X1  g0316(.A1(new_n329), .A2(new_n208), .A3(G87), .ZN(new_n517));
  INV_X1    g0317(.A(KEYINPUT92), .ZN(new_n518));
  OAI21_X1  g0318(.A(KEYINPUT22), .B1(new_n517), .B2(new_n518), .ZN(new_n519));
  NOR2_X1   g0319(.A1(new_n347), .A2(G20), .ZN(new_n520));
  AOI21_X1  g0320(.A(KEYINPUT92), .B1(new_n520), .B2(G87), .ZN(new_n521));
  OAI21_X1  g0321(.A(new_n516), .B1(new_n519), .B2(new_n521), .ZN(new_n522));
  OAI21_X1  g0322(.A(G116), .B1(new_n326), .B2(new_n327), .ZN(new_n523));
  INV_X1    g0323(.A(new_n523), .ZN(new_n524));
  INV_X1    g0324(.A(KEYINPUT23), .ZN(new_n525));
  OAI21_X1  g0325(.A(new_n525), .B1(new_n208), .B2(G107), .ZN(new_n526));
  NAND3_X1  g0326(.A1(new_n444), .A2(KEYINPUT23), .A3(G20), .ZN(new_n527));
  AOI22_X1  g0327(.A1(new_n524), .A2(new_n208), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  NAND3_X1  g0328(.A1(new_n522), .A2(KEYINPUT24), .A3(new_n528), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n529), .A2(new_n277), .ZN(new_n530));
  AOI21_X1  g0330(.A(KEYINPUT24), .B1(new_n522), .B2(new_n528), .ZN(new_n531));
  OAI21_X1  g0331(.A(new_n514), .B1(new_n530), .B2(new_n531), .ZN(new_n532));
  INV_X1    g0332(.A(G250), .ZN(new_n533));
  MUX2_X1   g0333(.A(new_n533), .B(new_n492), .S(G1698), .Z(new_n534));
  INV_X1    g0334(.A(G294), .ZN(new_n535));
  OAI22_X1  g0335(.A1(new_n347), .A2(new_n534), .B1(new_n535), .B2(new_n328), .ZN(new_n536));
  INV_X1    g0336(.A(new_n493), .ZN(new_n537));
  AOI22_X1  g0337(.A1(new_n536), .A2(new_n257), .B1(G264), .B2(new_n537), .ZN(new_n538));
  AND2_X1   g0338(.A1(new_n538), .A2(new_n491), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n539), .A2(G179), .ZN(new_n540));
  OAI21_X1  g0340(.A(new_n540), .B1(new_n428), .B2(new_n539), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n532), .A2(new_n541), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n539), .A2(new_n301), .ZN(new_n543));
  OAI21_X1  g0343(.A(new_n543), .B1(new_n539), .B2(G200), .ZN(new_n544));
  OAI211_X1 g0344(.A(new_n544), .B(new_n514), .C1(new_n530), .C2(new_n531), .ZN(new_n545));
  NAND4_X1  g0345(.A1(new_n320), .A2(new_n208), .A3(G68), .A4(new_n321), .ZN(new_n546));
  INV_X1    g0346(.A(KEYINPUT19), .ZN(new_n547));
  OAI21_X1  g0347(.A(new_n208), .B1(new_n399), .B2(new_n547), .ZN(new_n548));
  NOR2_X1   g0348(.A1(G87), .A2(G97), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n549), .A2(new_n444), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n548), .A2(new_n550), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n551), .A2(KEYINPUT83), .ZN(new_n552));
  INV_X1    g0352(.A(KEYINPUT83), .ZN(new_n553));
  NAND3_X1  g0353(.A1(new_n548), .A2(new_n550), .A3(new_n553), .ZN(new_n554));
  OAI21_X1  g0354(.A(new_n547), .B1(new_n399), .B2(G20), .ZN(new_n555));
  NAND4_X1  g0355(.A1(new_n546), .A2(new_n552), .A3(new_n554), .A4(new_n555), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n556), .A2(new_n277), .ZN(new_n557));
  INV_X1    g0357(.A(new_n435), .ZN(new_n558));
  NOR2_X1   g0358(.A1(new_n558), .A2(new_n292), .ZN(new_n559));
  INV_X1    g0359(.A(new_n559), .ZN(new_n560));
  OAI211_X1 g0360(.A(new_n557), .B(new_n560), .C1(new_n435), .C2(new_n474), .ZN(new_n561));
  NAND4_X1  g0361(.A1(new_n320), .A2(G238), .A3(new_n251), .A4(new_n321), .ZN(new_n562));
  NAND4_X1  g0362(.A1(new_n320), .A2(G244), .A3(G1698), .A4(new_n321), .ZN(new_n563));
  NAND3_X1  g0363(.A1(new_n562), .A2(new_n563), .A3(new_n523), .ZN(new_n564));
  NOR2_X1   g0364(.A1(new_n487), .A2(new_n533), .ZN(new_n565));
  NOR3_X1   g0365(.A1(new_n486), .A2(new_n260), .A3(G1), .ZN(new_n566));
  OAI21_X1  g0366(.A(new_n256), .B1(new_n565), .B2(new_n566), .ZN(new_n567));
  INV_X1    g0367(.A(KEYINPUT82), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  OAI211_X1 g0369(.A(KEYINPUT82), .B(new_n256), .C1(new_n565), .C2(new_n566), .ZN(new_n570));
  AOI22_X1  g0370(.A1(new_n564), .A2(new_n257), .B1(new_n569), .B2(new_n570), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n571), .A2(new_n273), .ZN(new_n572));
  OAI211_X1 g0372(.A(new_n561), .B(new_n572), .C1(G169), .C2(new_n571), .ZN(new_n573));
  NOR2_X1   g0373(.A1(new_n474), .A2(new_n515), .ZN(new_n574));
  AOI211_X1 g0374(.A(new_n559), .B(new_n574), .C1(new_n556), .C2(new_n277), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n571), .A2(G190), .ZN(new_n576));
  OAI211_X1 g0376(.A(new_n575), .B(new_n576), .C1(new_n419), .C2(new_n571), .ZN(new_n577));
  INV_X1    g0377(.A(KEYINPUT84), .ZN(new_n578));
  AND3_X1   g0378(.A1(new_n573), .A2(new_n577), .A3(new_n578), .ZN(new_n579));
  AOI21_X1  g0379(.A(new_n578), .B1(new_n573), .B2(new_n577), .ZN(new_n580));
  NOR2_X1   g0380(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  NAND4_X1  g0381(.A1(new_n509), .A2(new_n542), .A3(new_n545), .A4(new_n581), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n446), .A2(G303), .ZN(new_n583));
  NAND4_X1  g0383(.A1(new_n320), .A2(G264), .A3(G1698), .A4(new_n321), .ZN(new_n584));
  NAND4_X1  g0384(.A1(new_n320), .A2(G257), .A3(new_n251), .A4(new_n321), .ZN(new_n585));
  INV_X1    g0385(.A(KEYINPUT85), .ZN(new_n586));
  OAI211_X1 g0386(.A(new_n583), .B(new_n584), .C1(new_n585), .C2(new_n586), .ZN(new_n587));
  AND2_X1   g0387(.A1(new_n585), .A2(new_n586), .ZN(new_n588));
  OAI21_X1  g0388(.A(new_n257), .B1(new_n587), .B2(new_n588), .ZN(new_n589));
  INV_X1    g0389(.A(G270), .ZN(new_n590));
  OAI21_X1  g0390(.A(new_n491), .B1(new_n590), .B2(new_n493), .ZN(new_n591));
  INV_X1    g0391(.A(new_n591), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n589), .A2(new_n592), .ZN(new_n593));
  NOR2_X1   g0393(.A1(new_n593), .A2(new_n273), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n474), .A2(G116), .ZN(new_n595));
  OAI21_X1  g0395(.A(new_n595), .B1(G116), .B2(new_n295), .ZN(new_n596));
  OAI21_X1  g0396(.A(new_n208), .B1(new_n465), .B2(G33), .ZN(new_n597));
  INV_X1    g0397(.A(new_n483), .ZN(new_n598));
  OAI21_X1  g0398(.A(KEYINPUT87), .B1(new_n597), .B2(new_n598), .ZN(new_n599));
  AOI21_X1  g0399(.A(G20), .B1(new_n245), .B2(G97), .ZN(new_n600));
  INV_X1    g0400(.A(KEYINPUT87), .ZN(new_n601));
  NAND3_X1  g0401(.A1(new_n600), .A2(new_n601), .A3(new_n483), .ZN(new_n602));
  INV_X1    g0402(.A(G116), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n603), .A2(G20), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n277), .A2(new_n604), .ZN(new_n605));
  AOI22_X1  g0405(.A1(new_n599), .A2(new_n602), .B1(new_n605), .B2(KEYINPUT86), .ZN(new_n606));
  INV_X1    g0406(.A(KEYINPUT86), .ZN(new_n607));
  NAND3_X1  g0407(.A1(new_n277), .A2(new_n607), .A3(new_n604), .ZN(new_n608));
  AOI21_X1  g0408(.A(KEYINPUT20), .B1(new_n606), .B2(new_n608), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n599), .A2(new_n602), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n605), .A2(KEYINPUT86), .ZN(new_n611));
  AND4_X1   g0411(.A1(KEYINPUT20), .A2(new_n610), .A3(new_n608), .A4(new_n611), .ZN(new_n612));
  OAI21_X1  g0412(.A(new_n596), .B1(new_n609), .B2(new_n612), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n594), .A2(new_n613), .ZN(new_n614));
  NAND3_X1  g0414(.A1(new_n610), .A2(new_n608), .A3(new_n611), .ZN(new_n615));
  INV_X1    g0415(.A(KEYINPUT20), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n615), .A2(new_n616), .ZN(new_n617));
  NAND3_X1  g0417(.A1(new_n606), .A2(KEYINPUT20), .A3(new_n608), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  AOI21_X1  g0419(.A(new_n428), .B1(new_n619), .B2(new_n596), .ZN(new_n620));
  NAND3_X1  g0420(.A1(new_n620), .A2(KEYINPUT21), .A3(new_n593), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n614), .A2(new_n621), .ZN(new_n622));
  INV_X1    g0422(.A(new_n622), .ZN(new_n623));
  NAND3_X1  g0423(.A1(new_n589), .A2(new_n301), .A3(new_n592), .ZN(new_n624));
  NAND4_X1  g0424(.A1(new_n329), .A2(KEYINPUT85), .A3(G257), .A4(new_n251), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n585), .A2(new_n586), .ZN(new_n626));
  NAND4_X1  g0426(.A1(new_n625), .A2(new_n626), .A3(new_n583), .A4(new_n584), .ZN(new_n627));
  AOI21_X1  g0427(.A(new_n591), .B1(new_n627), .B2(new_n257), .ZN(new_n628));
  OAI21_X1  g0428(.A(new_n624), .B1(new_n628), .B2(G200), .ZN(new_n629));
  INV_X1    g0429(.A(KEYINPUT90), .ZN(new_n630));
  INV_X1    g0430(.A(new_n613), .ZN(new_n631));
  NAND3_X1  g0431(.A1(new_n629), .A2(new_n630), .A3(new_n631), .ZN(new_n632));
  INV_X1    g0432(.A(new_n632), .ZN(new_n633));
  AOI21_X1  g0433(.A(new_n630), .B1(new_n629), .B2(new_n631), .ZN(new_n634));
  NOR2_X1   g0434(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  NAND3_X1  g0435(.A1(new_n593), .A2(G169), .A3(new_n613), .ZN(new_n636));
  INV_X1    g0436(.A(KEYINPUT88), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  NAND3_X1  g0438(.A1(new_n620), .A2(KEYINPUT88), .A3(new_n593), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  INV_X1    g0440(.A(KEYINPUT21), .ZN(new_n641));
  AOI21_X1  g0441(.A(KEYINPUT89), .B1(new_n640), .B2(new_n641), .ZN(new_n642));
  INV_X1    g0442(.A(KEYINPUT89), .ZN(new_n643));
  AOI211_X1 g0443(.A(new_n643), .B(KEYINPUT21), .C1(new_n638), .C2(new_n639), .ZN(new_n644));
  OAI211_X1 g0444(.A(new_n623), .B(new_n635), .C1(new_n642), .C2(new_n644), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n645), .A2(KEYINPUT91), .ZN(new_n646));
  AND4_X1   g0446(.A1(KEYINPUT88), .A2(new_n593), .A3(G169), .A4(new_n613), .ZN(new_n647));
  AOI21_X1  g0447(.A(KEYINPUT88), .B1(new_n620), .B2(new_n593), .ZN(new_n648));
  OAI21_X1  g0448(.A(new_n641), .B1(new_n647), .B2(new_n648), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n649), .A2(new_n643), .ZN(new_n650));
  NAND3_X1  g0450(.A1(new_n640), .A2(KEYINPUT89), .A3(new_n641), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  INV_X1    g0452(.A(KEYINPUT91), .ZN(new_n653));
  NAND4_X1  g0453(.A1(new_n652), .A2(new_n653), .A3(new_n623), .A4(new_n635), .ZN(new_n654));
  AOI21_X1  g0454(.A(new_n582), .B1(new_n646), .B2(new_n654), .ZN(new_n655));
  AND2_X1   g0455(.A1(new_n463), .A2(new_n655), .ZN(G372));
  INV_X1    g0456(.A(new_n433), .ZN(new_n657));
  AOI21_X1  g0457(.A(new_n657), .B1(new_n425), .B2(new_n460), .ZN(new_n658));
  INV_X1    g0458(.A(new_n374), .ZN(new_n659));
  OAI21_X1  g0459(.A(new_n378), .B1(new_n658), .B2(new_n659), .ZN(new_n660));
  NAND3_X1  g0460(.A1(new_n660), .A2(new_n306), .A3(new_n307), .ZN(new_n661));
  AND2_X1   g0461(.A1(new_n661), .A2(new_n298), .ZN(new_n662));
  NOR2_X1   g0462(.A1(new_n571), .A2(new_n419), .ZN(new_n663));
  OAI211_X1 g0463(.A(new_n557), .B(new_n560), .C1(new_n515), .C2(new_n474), .ZN(new_n664));
  OAI21_X1  g0464(.A(KEYINPUT94), .B1(new_n663), .B2(new_n664), .ZN(new_n665));
  INV_X1    g0465(.A(KEYINPUT94), .ZN(new_n666));
  OAI211_X1 g0466(.A(new_n575), .B(new_n666), .C1(new_n419), .C2(new_n571), .ZN(new_n667));
  NAND3_X1  g0467(.A1(new_n665), .A2(new_n667), .A3(new_n576), .ZN(new_n668));
  INV_X1    g0468(.A(KEYINPUT26), .ZN(new_n669));
  OR3_X1    g0469(.A1(new_n571), .A2(KEYINPUT93), .A3(G169), .ZN(new_n670));
  OAI21_X1  g0470(.A(KEYINPUT93), .B1(new_n571), .B2(G169), .ZN(new_n671));
  NAND4_X1  g0471(.A1(new_n670), .A2(new_n671), .A3(new_n561), .A4(new_n572), .ZN(new_n672));
  NAND4_X1  g0472(.A1(new_n668), .A2(new_n669), .A3(new_n502), .A4(new_n672), .ZN(new_n673));
  INV_X1    g0473(.A(KEYINPUT95), .ZN(new_n674));
  XNOR2_X1  g0474(.A(new_n672), .B(new_n674), .ZN(new_n675));
  NOR3_X1   g0475(.A1(new_n579), .A2(new_n580), .A3(new_n505), .ZN(new_n676));
  OAI211_X1 g0476(.A(new_n673), .B(new_n675), .C1(new_n676), .C2(new_n669), .ZN(new_n677));
  INV_X1    g0477(.A(new_n677), .ZN(new_n678));
  OAI211_X1 g0478(.A(new_n623), .B(new_n542), .C1(new_n642), .C2(new_n644), .ZN(new_n679));
  NOR2_X1   g0479(.A1(new_n499), .A2(new_n502), .ZN(new_n680));
  AND4_X1   g0480(.A1(new_n680), .A2(new_n545), .A3(new_n672), .A4(new_n668), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n679), .A2(new_n681), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n678), .A2(new_n682), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n463), .A2(new_n683), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n662), .A2(new_n684), .ZN(G369));
  INV_X1    g0485(.A(new_n291), .ZN(new_n686));
  OR3_X1    g0486(.A1(new_n686), .A2(KEYINPUT27), .A3(G20), .ZN(new_n687));
  OAI21_X1  g0487(.A(KEYINPUT27), .B1(new_n686), .B2(G20), .ZN(new_n688));
  NAND3_X1  g0488(.A1(new_n687), .A2(G213), .A3(new_n688), .ZN(new_n689));
  INV_X1    g0489(.A(G343), .ZN(new_n690));
  NOR2_X1   g0490(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n613), .A2(new_n691), .ZN(new_n692));
  NAND3_X1  g0492(.A1(new_n646), .A2(new_n654), .A3(new_n692), .ZN(new_n693));
  AOI21_X1  g0493(.A(new_n622), .B1(new_n650), .B2(new_n651), .ZN(new_n694));
  NAND3_X1  g0494(.A1(new_n694), .A2(new_n613), .A3(new_n691), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n693), .A2(new_n695), .ZN(new_n696));
  INV_X1    g0496(.A(G330), .ZN(new_n697));
  NOR2_X1   g0497(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  NOR2_X1   g0498(.A1(new_n542), .A2(new_n691), .ZN(new_n699));
  INV_X1    g0499(.A(new_n532), .ZN(new_n700));
  INV_X1    g0500(.A(new_n691), .ZN(new_n701));
  OAI21_X1  g0501(.A(new_n545), .B1(new_n700), .B2(new_n701), .ZN(new_n702));
  AOI21_X1  g0502(.A(new_n699), .B1(new_n702), .B2(new_n542), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n698), .A2(new_n703), .ZN(new_n704));
  NOR2_X1   g0504(.A1(new_n694), .A2(new_n691), .ZN(new_n705));
  AOI21_X1  g0505(.A(new_n699), .B1(new_n705), .B2(new_n703), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n704), .A2(new_n706), .ZN(G399));
  INV_X1    g0507(.A(G41), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n211), .A2(new_n708), .ZN(new_n709));
  INV_X1    g0509(.A(new_n709), .ZN(new_n710));
  NAND3_X1  g0510(.A1(new_n549), .A2(new_n444), .A3(new_n603), .ZN(new_n711));
  NOR3_X1   g0511(.A1(new_n710), .A2(new_n207), .A3(new_n711), .ZN(new_n712));
  AOI21_X1  g0512(.A(new_n712), .B1(new_n217), .B2(new_n710), .ZN(new_n713));
  XOR2_X1   g0513(.A(new_n713), .B(KEYINPUT28), .Z(new_n714));
  NAND3_X1  g0514(.A1(new_n581), .A2(new_n669), .A3(new_n502), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n668), .A2(new_n672), .ZN(new_n716));
  OAI21_X1  g0516(.A(KEYINPUT26), .B1(new_n716), .B2(new_n505), .ZN(new_n717));
  NAND3_X1  g0517(.A1(new_n715), .A2(new_n717), .A3(new_n675), .ZN(new_n718));
  AOI21_X1  g0518(.A(new_n718), .B1(new_n682), .B2(KEYINPUT96), .ZN(new_n719));
  INV_X1    g0519(.A(KEYINPUT96), .ZN(new_n720));
  NAND3_X1  g0520(.A1(new_n679), .A2(new_n720), .A3(new_n681), .ZN(new_n721));
  AOI21_X1  g0521(.A(new_n691), .B1(new_n719), .B2(new_n721), .ZN(new_n722));
  NAND2_X1  g0522(.A1(new_n722), .A2(KEYINPUT29), .ZN(new_n723));
  AOI21_X1  g0523(.A(new_n691), .B1(new_n678), .B2(new_n682), .ZN(new_n724));
  OR2_X1    g0524(.A1(new_n724), .A2(KEYINPUT29), .ZN(new_n725));
  NAND2_X1  g0525(.A1(new_n723), .A2(new_n725), .ZN(new_n726));
  INV_X1    g0526(.A(new_n582), .ZN(new_n727));
  INV_X1    g0527(.A(new_n654), .ZN(new_n728));
  AOI21_X1  g0528(.A(new_n653), .B1(new_n694), .B2(new_n635), .ZN(new_n729));
  OAI211_X1 g0529(.A(new_n727), .B(new_n701), .C1(new_n728), .C2(new_n729), .ZN(new_n730));
  NOR2_X1   g0530(.A1(new_n485), .A2(new_n494), .ZN(new_n731));
  NAND4_X1  g0531(.A1(new_n594), .A2(new_n538), .A3(new_n731), .A4(new_n571), .ZN(new_n732));
  INV_X1    g0532(.A(KEYINPUT30), .ZN(new_n733));
  OR2_X1    g0533(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n732), .A2(new_n733), .ZN(new_n735));
  NOR4_X1   g0535(.A1(new_n539), .A2(new_n731), .A3(G179), .A4(new_n571), .ZN(new_n736));
  NAND2_X1  g0536(.A1(new_n736), .A2(new_n593), .ZN(new_n737));
  NAND3_X1  g0537(.A1(new_n734), .A2(new_n735), .A3(new_n737), .ZN(new_n738));
  NAND2_X1  g0538(.A1(new_n738), .A2(new_n691), .ZN(new_n739));
  INV_X1    g0539(.A(KEYINPUT31), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  NAND3_X1  g0541(.A1(new_n738), .A2(KEYINPUT31), .A3(new_n691), .ZN(new_n742));
  NAND2_X1  g0542(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  INV_X1    g0543(.A(new_n743), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n730), .A2(new_n744), .ZN(new_n745));
  NAND2_X1  g0545(.A1(new_n745), .A2(G330), .ZN(new_n746));
  NAND2_X1  g0546(.A1(new_n726), .A2(new_n746), .ZN(new_n747));
  INV_X1    g0547(.A(new_n747), .ZN(new_n748));
  OAI21_X1  g0548(.A(new_n714), .B1(new_n748), .B2(G1), .ZN(G364));
  NOR2_X1   g0549(.A1(new_n290), .A2(G20), .ZN(new_n750));
  NAND2_X1  g0550(.A1(new_n750), .A2(G45), .ZN(new_n751));
  NAND3_X1  g0551(.A1(new_n709), .A2(G1), .A3(new_n751), .ZN(new_n752));
  INV_X1    g0552(.A(new_n696), .ZN(new_n753));
  NOR2_X1   g0553(.A1(new_n753), .A2(G330), .ZN(new_n754));
  OAI21_X1  g0554(.A(new_n752), .B1(new_n754), .B2(new_n698), .ZN(new_n755));
  INV_X1    g0555(.A(new_n752), .ZN(new_n756));
  NOR2_X1   g0556(.A1(G13), .A2(G33), .ZN(new_n757));
  INV_X1    g0557(.A(new_n757), .ZN(new_n758));
  NOR2_X1   g0558(.A1(new_n758), .A2(G20), .ZN(new_n759));
  AND2_X1   g0559(.A1(new_n696), .A2(new_n759), .ZN(new_n760));
  NOR2_X1   g0560(.A1(new_n208), .A2(G190), .ZN(new_n761));
  NOR2_X1   g0561(.A1(G179), .A2(G200), .ZN(new_n762));
  NAND2_X1  g0562(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  INV_X1    g0563(.A(G159), .ZN(new_n764));
  NOR2_X1   g0564(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  XNOR2_X1  g0565(.A(new_n765), .B(KEYINPUT32), .ZN(new_n766));
  NOR2_X1   g0566(.A1(new_n273), .A2(G200), .ZN(new_n767));
  NAND2_X1  g0567(.A1(new_n761), .A2(new_n767), .ZN(new_n768));
  INV_X1    g0568(.A(new_n768), .ZN(new_n769));
  NOR2_X1   g0569(.A1(new_n419), .A2(G179), .ZN(new_n770));
  NAND2_X1  g0570(.A1(new_n761), .A2(new_n770), .ZN(new_n771));
  INV_X1    g0571(.A(new_n771), .ZN(new_n772));
  AOI22_X1  g0572(.A1(G77), .A2(new_n769), .B1(new_n772), .B2(G107), .ZN(new_n773));
  INV_X1    g0573(.A(G50), .ZN(new_n774));
  NOR2_X1   g0574(.A1(new_n273), .A2(new_n419), .ZN(new_n775));
  NOR2_X1   g0575(.A1(new_n208), .A2(new_n301), .ZN(new_n776));
  NAND2_X1  g0576(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  OAI211_X1 g0577(.A(new_n766), .B(new_n773), .C1(new_n774), .C2(new_n777), .ZN(new_n778));
  NAND2_X1  g0578(.A1(new_n762), .A2(G190), .ZN(new_n779));
  NAND2_X1  g0579(.A1(new_n779), .A2(G20), .ZN(new_n780));
  INV_X1    g0580(.A(new_n780), .ZN(new_n781));
  NOR2_X1   g0581(.A1(new_n781), .A2(new_n465), .ZN(new_n782));
  INV_X1    g0582(.A(G58), .ZN(new_n783));
  NAND2_X1  g0583(.A1(new_n776), .A2(new_n767), .ZN(new_n784));
  NAND2_X1  g0584(.A1(new_n776), .A2(new_n770), .ZN(new_n785));
  OAI22_X1  g0585(.A1(new_n783), .A2(new_n784), .B1(new_n785), .B2(new_n515), .ZN(new_n786));
  NAND2_X1  g0586(.A1(new_n775), .A2(new_n761), .ZN(new_n787));
  OAI21_X1  g0587(.A(new_n249), .B1(new_n787), .B2(new_n220), .ZN(new_n788));
  OR3_X1    g0588(.A1(new_n782), .A2(new_n786), .A3(new_n788), .ZN(new_n789));
  INV_X1    g0589(.A(new_n777), .ZN(new_n790));
  INV_X1    g0590(.A(new_n785), .ZN(new_n791));
  AOI22_X1  g0591(.A1(G326), .A2(new_n790), .B1(new_n791), .B2(G303), .ZN(new_n792));
  INV_X1    g0592(.A(G311), .ZN(new_n793));
  XOR2_X1   g0593(.A(KEYINPUT33), .B(G317), .Z(new_n794));
  OAI221_X1 g0594(.A(new_n792), .B1(new_n793), .B2(new_n768), .C1(new_n787), .C2(new_n794), .ZN(new_n795));
  INV_X1    g0595(.A(new_n763), .ZN(new_n796));
  AOI22_X1  g0596(.A1(G283), .A2(new_n772), .B1(new_n796), .B2(G329), .ZN(new_n797));
  INV_X1    g0597(.A(new_n784), .ZN(new_n798));
  AOI21_X1  g0598(.A(new_n249), .B1(new_n798), .B2(G322), .ZN(new_n799));
  OAI211_X1 g0599(.A(new_n797), .B(new_n799), .C1(new_n535), .C2(new_n781), .ZN(new_n800));
  OAI22_X1  g0600(.A1(new_n778), .A2(new_n789), .B1(new_n795), .B2(new_n800), .ZN(new_n801));
  AOI21_X1  g0601(.A(new_n214), .B1(G20), .B2(new_n428), .ZN(new_n802));
  NAND2_X1  g0602(.A1(new_n801), .A2(new_n802), .ZN(new_n803));
  NAND3_X1  g0603(.A1(new_n211), .A2(G355), .A3(new_n249), .ZN(new_n804));
  NOR2_X1   g0604(.A1(new_n217), .A2(G45), .ZN(new_n805));
  AOI21_X1  g0605(.A(new_n805), .B1(new_n240), .B2(G45), .ZN(new_n806));
  NAND2_X1  g0606(.A1(new_n211), .A2(new_n347), .ZN(new_n807));
  OAI221_X1 g0607(.A(new_n804), .B1(G116), .B2(new_n211), .C1(new_n806), .C2(new_n807), .ZN(new_n808));
  NOR2_X1   g0608(.A1(new_n759), .A2(new_n802), .ZN(new_n809));
  XOR2_X1   g0609(.A(new_n809), .B(KEYINPUT97), .Z(new_n810));
  NAND2_X1  g0610(.A1(new_n808), .A2(new_n810), .ZN(new_n811));
  NAND2_X1  g0611(.A1(new_n803), .A2(new_n811), .ZN(new_n812));
  OAI21_X1  g0612(.A(new_n756), .B1(new_n760), .B2(new_n812), .ZN(new_n813));
  NAND2_X1  g0613(.A1(new_n755), .A2(new_n813), .ZN(new_n814));
  INV_X1    g0614(.A(new_n814), .ZN(G396));
  INV_X1    g0615(.A(new_n802), .ZN(new_n816));
  NAND2_X1  g0616(.A1(new_n816), .A2(new_n758), .ZN(new_n817));
  AOI21_X1  g0617(.A(new_n249), .B1(new_n796), .B2(G311), .ZN(new_n818));
  OAI221_X1 g0618(.A(new_n818), .B1(new_n444), .B2(new_n785), .C1(new_n603), .C2(new_n768), .ZN(new_n819));
  NAND2_X1  g0619(.A1(new_n772), .A2(G87), .ZN(new_n820));
  OAI21_X1  g0620(.A(new_n820), .B1(new_n535), .B2(new_n784), .ZN(new_n821));
  INV_X1    g0621(.A(G303), .ZN(new_n822));
  INV_X1    g0622(.A(G283), .ZN(new_n823));
  OAI22_X1  g0623(.A1(new_n777), .A2(new_n822), .B1(new_n787), .B2(new_n823), .ZN(new_n824));
  NOR4_X1   g0624(.A1(new_n819), .A2(new_n782), .A3(new_n821), .A4(new_n824), .ZN(new_n825));
  INV_X1    g0625(.A(G132), .ZN(new_n826));
  OAI21_X1  g0626(.A(new_n329), .B1(new_n826), .B2(new_n763), .ZN(new_n827));
  INV_X1    g0627(.A(G137), .ZN(new_n828));
  NOR2_X1   g0628(.A1(new_n777), .A2(new_n828), .ZN(new_n829));
  INV_X1    g0629(.A(G143), .ZN(new_n830));
  OAI22_X1  g0630(.A1(new_n830), .A2(new_n784), .B1(new_n787), .B2(new_n279), .ZN(new_n831));
  AOI211_X1 g0631(.A(new_n829), .B(new_n831), .C1(G159), .C2(new_n769), .ZN(new_n832));
  NOR2_X1   g0632(.A1(new_n832), .A2(KEYINPUT34), .ZN(new_n833));
  AOI211_X1 g0633(.A(new_n827), .B(new_n833), .C1(G58), .C2(new_n780), .ZN(new_n834));
  OAI22_X1  g0634(.A1(new_n785), .A2(new_n774), .B1(new_n771), .B2(new_n220), .ZN(new_n835));
  XNOR2_X1  g0635(.A(new_n835), .B(KEYINPUT98), .ZN(new_n836));
  AOI21_X1  g0636(.A(new_n836), .B1(new_n832), .B2(KEYINPUT34), .ZN(new_n837));
  AOI21_X1  g0637(.A(new_n825), .B1(new_n834), .B2(new_n837), .ZN(new_n838));
  OAI221_X1 g0638(.A(new_n756), .B1(G77), .B2(new_n817), .C1(new_n838), .C2(new_n816), .ZN(new_n839));
  INV_X1    g0639(.A(new_n460), .ZN(new_n840));
  NOR2_X1   g0640(.A1(new_n840), .A2(new_n701), .ZN(new_n841));
  INV_X1    g0641(.A(new_n841), .ZN(new_n842));
  NOR2_X1   g0642(.A1(new_n441), .A2(new_n701), .ZN(new_n843));
  INV_X1    g0643(.A(new_n843), .ZN(new_n844));
  AOI21_X1  g0644(.A(KEYINPUT99), .B1(new_n461), .B2(new_n844), .ZN(new_n845));
  INV_X1    g0645(.A(KEYINPUT99), .ZN(new_n846));
  NOR4_X1   g0646(.A1(new_n457), .A2(new_n460), .A3(new_n846), .A4(new_n843), .ZN(new_n847));
  OAI21_X1  g0647(.A(new_n842), .B1(new_n845), .B2(new_n847), .ZN(new_n848));
  INV_X1    g0648(.A(new_n848), .ZN(new_n849));
  AOI21_X1  g0649(.A(new_n839), .B1(new_n849), .B2(new_n757), .ZN(new_n850));
  XOR2_X1   g0650(.A(new_n850), .B(KEYINPUT100), .Z(new_n851));
  XNOR2_X1  g0651(.A(new_n724), .B(new_n848), .ZN(new_n852));
  OAI21_X1  g0652(.A(new_n752), .B1(new_n852), .B2(new_n746), .ZN(new_n853));
  INV_X1    g0653(.A(new_n853), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n852), .A2(new_n746), .ZN(new_n855));
  AOI21_X1  g0655(.A(new_n851), .B1(new_n854), .B2(new_n855), .ZN(new_n856));
  INV_X1    g0656(.A(new_n856), .ZN(G384));
  INV_X1    g0657(.A(new_n470), .ZN(new_n858));
  OAI211_X1 g0658(.A(G116), .B(new_n215), .C1(new_n858), .C2(KEYINPUT35), .ZN(new_n859));
  AOI21_X1  g0659(.A(new_n859), .B1(KEYINPUT35), .B2(new_n858), .ZN(new_n860));
  XNOR2_X1  g0660(.A(KEYINPUT101), .B(KEYINPUT36), .ZN(new_n861));
  XNOR2_X1  g0661(.A(new_n860), .B(new_n861), .ZN(new_n862));
  NAND3_X1  g0662(.A1(new_n217), .A2(G77), .A3(new_n350), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n774), .A2(G68), .ZN(new_n864));
  XNOR2_X1  g0664(.A(new_n864), .B(KEYINPUT102), .ZN(new_n865));
  AOI211_X1 g0665(.A(new_n207), .B(G13), .C1(new_n863), .C2(new_n865), .ZN(new_n866));
  NOR2_X1   g0666(.A1(new_n862), .A2(new_n866), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n657), .A2(new_n701), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n368), .A2(new_n311), .ZN(new_n869));
  INV_X1    g0669(.A(new_n376), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n871), .A2(KEYINPUT18), .ZN(new_n872));
  INV_X1    g0672(.A(KEYINPUT18), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n377), .A2(new_n873), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n872), .A2(new_n874), .ZN(new_n875));
  AOI21_X1  g0675(.A(new_n875), .B1(new_n373), .B2(new_n371), .ZN(new_n876));
  AND2_X1   g0676(.A1(new_n354), .A2(new_n352), .ZN(new_n877));
  AOI21_X1  g0677(.A(KEYINPUT16), .B1(new_n877), .B2(new_n349), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n355), .A2(new_n277), .ZN(new_n879));
  OAI21_X1  g0679(.A(new_n311), .B1(new_n878), .B2(new_n879), .ZN(new_n880));
  INV_X1    g0680(.A(new_n689), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  OAI21_X1  g0682(.A(KEYINPUT103), .B1(new_n876), .B2(new_n882), .ZN(new_n883));
  INV_X1    g0683(.A(KEYINPUT103), .ZN(new_n884));
  INV_X1    g0684(.A(new_n882), .ZN(new_n885));
  NAND3_X1  g0685(.A1(new_n379), .A2(new_n884), .A3(new_n885), .ZN(new_n886));
  AND2_X1   g0686(.A1(new_n364), .A2(new_n370), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n869), .A2(new_n881), .ZN(new_n888));
  INV_X1    g0688(.A(KEYINPUT37), .ZN(new_n889));
  AND3_X1   g0689(.A1(new_n871), .A2(new_n888), .A3(new_n889), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n376), .A2(new_n689), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n880), .A2(new_n891), .ZN(new_n892));
  NAND3_X1  g0692(.A1(new_n892), .A2(new_n364), .A3(new_n370), .ZN(new_n893));
  AOI22_X1  g0693(.A1(new_n887), .A2(new_n890), .B1(new_n893), .B2(KEYINPUT37), .ZN(new_n894));
  INV_X1    g0694(.A(new_n894), .ZN(new_n895));
  NAND4_X1  g0695(.A1(new_n883), .A2(KEYINPUT38), .A3(new_n886), .A4(new_n895), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n896), .A2(KEYINPUT104), .ZN(new_n897));
  INV_X1    g0697(.A(KEYINPUT39), .ZN(new_n898));
  AOI21_X1  g0698(.A(new_n882), .B1(new_n374), .B2(new_n378), .ZN(new_n899));
  AOI21_X1  g0699(.A(new_n894), .B1(new_n899), .B2(new_n884), .ZN(new_n900));
  INV_X1    g0700(.A(KEYINPUT104), .ZN(new_n901));
  NAND4_X1  g0701(.A1(new_n900), .A2(new_n901), .A3(new_n883), .A4(KEYINPUT38), .ZN(new_n902));
  INV_X1    g0702(.A(KEYINPUT38), .ZN(new_n903));
  NOR2_X1   g0703(.A1(new_n876), .A2(new_n888), .ZN(new_n904));
  NAND3_X1  g0704(.A1(new_n871), .A2(new_n888), .A3(new_n372), .ZN(new_n905));
  AOI22_X1  g0705(.A1(new_n890), .A2(new_n887), .B1(KEYINPUT37), .B2(new_n905), .ZN(new_n906));
  OAI21_X1  g0706(.A(new_n903), .B1(new_n904), .B2(new_n906), .ZN(new_n907));
  NAND4_X1  g0707(.A1(new_n897), .A2(new_n898), .A3(new_n902), .A4(new_n907), .ZN(new_n908));
  AND3_X1   g0708(.A1(new_n900), .A2(KEYINPUT38), .A3(new_n883), .ZN(new_n909));
  AOI21_X1  g0709(.A(KEYINPUT38), .B1(new_n900), .B2(new_n883), .ZN(new_n910));
  OAI21_X1  g0710(.A(KEYINPUT39), .B1(new_n909), .B2(new_n910), .ZN(new_n911));
  AOI21_X1  g0711(.A(new_n868), .B1(new_n908), .B2(new_n911), .ZN(new_n912));
  NOR2_X1   g0712(.A1(new_n840), .A2(new_n691), .ZN(new_n913));
  AOI21_X1  g0713(.A(new_n913), .B1(new_n724), .B2(new_n848), .ZN(new_n914));
  INV_X1    g0714(.A(new_n914), .ZN(new_n915));
  NOR2_X1   g0715(.A1(new_n389), .A2(new_n701), .ZN(new_n916));
  INV_X1    g0716(.A(new_n916), .ZN(new_n917));
  NOR2_X1   g0717(.A1(new_n417), .A2(KEYINPUT75), .ZN(new_n918));
  AOI21_X1  g0718(.A(new_n423), .B1(new_n422), .B2(new_n389), .ZN(new_n919));
  OAI211_X1 g0719(.A(new_n433), .B(new_n917), .C1(new_n918), .C2(new_n919), .ZN(new_n920));
  INV_X1    g0720(.A(new_n920), .ZN(new_n921));
  AOI21_X1  g0721(.A(new_n917), .B1(new_n425), .B2(new_n433), .ZN(new_n922));
  NOR2_X1   g0722(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  INV_X1    g0723(.A(new_n923), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n915), .A2(new_n924), .ZN(new_n925));
  NOR2_X1   g0725(.A1(new_n909), .A2(new_n910), .ZN(new_n926));
  OAI22_X1  g0726(.A1(new_n925), .A2(new_n926), .B1(new_n378), .B2(new_n881), .ZN(new_n927));
  OR2_X1    g0727(.A1(new_n912), .A2(new_n927), .ZN(new_n928));
  NAND3_X1  g0728(.A1(new_n723), .A2(new_n463), .A3(new_n725), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n929), .A2(new_n662), .ZN(new_n930));
  XNOR2_X1  g0730(.A(new_n928), .B(new_n930), .ZN(new_n931));
  AND2_X1   g0731(.A1(new_n745), .A2(new_n463), .ZN(new_n932));
  XOR2_X1   g0732(.A(new_n932), .B(KEYINPUT105), .Z(new_n933));
  INV_X1    g0733(.A(KEYINPUT40), .ZN(new_n934));
  OAI21_X1  g0734(.A(new_n848), .B1(new_n921), .B2(new_n922), .ZN(new_n935));
  INV_X1    g0735(.A(new_n935), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n745), .A2(new_n936), .ZN(new_n937));
  OAI21_X1  g0737(.A(new_n934), .B1(new_n926), .B2(new_n937), .ZN(new_n938));
  NAND3_X1  g0738(.A1(new_n897), .A2(new_n902), .A3(new_n907), .ZN(new_n939));
  AOI21_X1  g0739(.A(new_n743), .B1(new_n655), .B2(new_n701), .ZN(new_n940));
  NOR3_X1   g0740(.A1(new_n940), .A2(new_n934), .A3(new_n935), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n939), .A2(new_n941), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n938), .A2(new_n942), .ZN(new_n943));
  OR2_X1    g0743(.A1(new_n933), .A2(new_n943), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n933), .A2(new_n943), .ZN(new_n945));
  NAND3_X1  g0745(.A1(new_n944), .A2(G330), .A3(new_n945), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n931), .A2(new_n946), .ZN(new_n947));
  OAI21_X1  g0747(.A(new_n947), .B1(new_n207), .B2(new_n750), .ZN(new_n948));
  NOR2_X1   g0748(.A1(new_n931), .A2(new_n946), .ZN(new_n949));
  OAI21_X1  g0749(.A(new_n867), .B1(new_n948), .B2(new_n949), .ZN(G367));
  NOR2_X1   g0750(.A1(new_n575), .A2(new_n701), .ZN(new_n951));
  XNOR2_X1  g0751(.A(new_n951), .B(KEYINPUT106), .ZN(new_n952));
  MUX2_X1   g0752(.A(new_n716), .B(new_n675), .S(new_n952), .Z(new_n953));
  INV_X1    g0753(.A(KEYINPUT43), .ZN(new_n954));
  NOR2_X1   g0754(.A1(new_n953), .A2(new_n954), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n476), .A2(new_n691), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n680), .A2(new_n956), .ZN(new_n957));
  XOR2_X1   g0757(.A(new_n957), .B(KEYINPUT107), .Z(new_n958));
  OAI21_X1  g0758(.A(new_n958), .B1(new_n505), .B2(new_n701), .ZN(new_n959));
  NAND3_X1  g0759(.A1(new_n959), .A2(new_n703), .A3(new_n705), .ZN(new_n960));
  NOR2_X1   g0760(.A1(new_n960), .A2(KEYINPUT42), .ZN(new_n961));
  OR2_X1    g0761(.A1(new_n958), .A2(new_n542), .ZN(new_n962));
  AOI21_X1  g0762(.A(new_n691), .B1(new_n962), .B2(new_n505), .ZN(new_n963));
  NOR2_X1   g0763(.A1(new_n961), .A2(new_n963), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n960), .A2(KEYINPUT42), .ZN(new_n965));
  AOI21_X1  g0765(.A(new_n955), .B1(new_n964), .B2(new_n965), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n953), .A2(new_n954), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n966), .A2(new_n967), .ZN(new_n968));
  NAND4_X1  g0768(.A1(new_n964), .A2(new_n954), .A3(new_n953), .A4(new_n965), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n968), .A2(new_n969), .ZN(new_n970));
  INV_X1    g0770(.A(new_n959), .ZN(new_n971));
  NOR2_X1   g0771(.A1(new_n704), .A2(new_n971), .ZN(new_n972));
  INV_X1    g0772(.A(new_n972), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n970), .A2(new_n973), .ZN(new_n974));
  INV_X1    g0774(.A(KEYINPUT108), .ZN(new_n975));
  NAND4_X1  g0775(.A1(new_n968), .A2(new_n975), .A3(new_n972), .A4(new_n969), .ZN(new_n976));
  AND2_X1   g0776(.A1(new_n974), .A2(new_n976), .ZN(new_n977));
  OAI21_X1  g0777(.A(KEYINPUT108), .B1(new_n970), .B2(new_n973), .ZN(new_n978));
  XNOR2_X1  g0778(.A(new_n709), .B(KEYINPUT41), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n706), .A2(new_n959), .ZN(new_n980));
  XNOR2_X1  g0780(.A(new_n980), .B(KEYINPUT45), .ZN(new_n981));
  INV_X1    g0781(.A(new_n981), .ZN(new_n982));
  OR3_X1    g0782(.A1(new_n706), .A2(new_n959), .A3(KEYINPUT44), .ZN(new_n983));
  OAI21_X1  g0783(.A(KEYINPUT44), .B1(new_n706), .B2(new_n959), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n983), .A2(new_n984), .ZN(new_n985));
  INV_X1    g0785(.A(new_n985), .ZN(new_n986));
  AOI21_X1  g0786(.A(new_n704), .B1(new_n982), .B2(new_n986), .ZN(new_n987));
  INV_X1    g0787(.A(new_n704), .ZN(new_n988));
  NOR3_X1   g0788(.A1(new_n988), .A2(new_n981), .A3(new_n985), .ZN(new_n989));
  NOR2_X1   g0789(.A1(new_n987), .A2(new_n989), .ZN(new_n990));
  XNOR2_X1  g0790(.A(new_n705), .B(new_n703), .ZN(new_n991));
  XNOR2_X1  g0791(.A(new_n698), .B(new_n991), .ZN(new_n992));
  INV_X1    g0792(.A(new_n992), .ZN(new_n993));
  NOR2_X1   g0793(.A1(new_n993), .A2(new_n747), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n990), .A2(new_n994), .ZN(new_n995));
  AOI21_X1  g0795(.A(new_n979), .B1(new_n995), .B2(new_n748), .ZN(new_n996));
  NAND2_X1  g0796(.A1(new_n751), .A2(G1), .ZN(new_n997));
  OAI211_X1 g0797(.A(new_n977), .B(new_n978), .C1(new_n996), .C2(new_n997), .ZN(new_n998));
  OAI221_X1 g0798(.A(new_n809), .B1(new_n211), .B2(new_n435), .C1(new_n236), .C2(new_n807), .ZN(new_n999));
  INV_X1    g0799(.A(KEYINPUT109), .ZN(new_n1000));
  OAI21_X1  g0800(.A(new_n756), .B1(new_n999), .B2(new_n1000), .ZN(new_n1001));
  AOI21_X1  g0801(.A(new_n1001), .B1(new_n1000), .B2(new_n999), .ZN(new_n1002));
  NOR2_X1   g0802(.A1(new_n771), .A2(new_n465), .ZN(new_n1003));
  OAI22_X1  g0803(.A1(new_n784), .A2(new_n822), .B1(new_n768), .B2(new_n823), .ZN(new_n1004));
  AOI211_X1 g0804(.A(new_n1003), .B(new_n1004), .C1(G317), .C2(new_n796), .ZN(new_n1005));
  NAND2_X1  g0805(.A1(new_n780), .A2(G107), .ZN(new_n1006));
  OAI22_X1  g0806(.A1(new_n777), .A2(new_n793), .B1(new_n787), .B2(new_n535), .ZN(new_n1007));
  NOR2_X1   g0807(.A1(new_n1007), .A2(new_n329), .ZN(new_n1008));
  NAND2_X1  g0808(.A1(new_n791), .A2(G116), .ZN(new_n1009));
  XNOR2_X1  g0809(.A(new_n1009), .B(KEYINPUT46), .ZN(new_n1010));
  NAND4_X1  g0810(.A1(new_n1005), .A2(new_n1006), .A3(new_n1008), .A4(new_n1010), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n772), .A2(G77), .ZN(new_n1012));
  OAI21_X1  g0812(.A(new_n1012), .B1(new_n830), .B2(new_n777), .ZN(new_n1013));
  NOR2_X1   g0813(.A1(new_n781), .A2(new_n220), .ZN(new_n1014));
  OAI21_X1  g0814(.A(new_n249), .B1(new_n784), .B2(new_n279), .ZN(new_n1015));
  OR3_X1    g0815(.A1(new_n1013), .A2(new_n1014), .A3(new_n1015), .ZN(new_n1016));
  INV_X1    g0816(.A(new_n787), .ZN(new_n1017));
  AOI22_X1  g0817(.A1(G159), .A2(new_n1017), .B1(new_n769), .B2(G50), .ZN(new_n1018));
  OR2_X1    g0818(.A1(new_n1018), .A2(KEYINPUT110), .ZN(new_n1019));
  OAI22_X1  g0819(.A1(new_n785), .A2(new_n783), .B1(new_n763), .B2(new_n828), .ZN(new_n1020));
  XNOR2_X1  g0820(.A(new_n1020), .B(KEYINPUT111), .ZN(new_n1021));
  NAND2_X1  g0821(.A1(new_n1018), .A2(KEYINPUT110), .ZN(new_n1022));
  NAND3_X1  g0822(.A1(new_n1019), .A2(new_n1021), .A3(new_n1022), .ZN(new_n1023));
  OAI21_X1  g0823(.A(new_n1011), .B1(new_n1016), .B2(new_n1023), .ZN(new_n1024));
  INV_X1    g0824(.A(KEYINPUT47), .ZN(new_n1025));
  AND2_X1   g0825(.A1(new_n1024), .A2(new_n1025), .ZN(new_n1026));
  OAI21_X1  g0826(.A(new_n802), .B1(new_n1024), .B2(new_n1025), .ZN(new_n1027));
  OAI21_X1  g0827(.A(new_n1002), .B1(new_n1026), .B2(new_n1027), .ZN(new_n1028));
  XOR2_X1   g0828(.A(new_n1028), .B(KEYINPUT112), .Z(new_n1029));
  AOI21_X1  g0829(.A(new_n1029), .B1(new_n759), .B2(new_n953), .ZN(new_n1030));
  XOR2_X1   g0830(.A(new_n1030), .B(KEYINPUT113), .Z(new_n1031));
  NAND2_X1  g0831(.A1(new_n998), .A2(new_n1031), .ZN(G387));
  INV_X1    g0832(.A(new_n994), .ZN(new_n1033));
  NAND2_X1  g0833(.A1(new_n993), .A2(new_n747), .ZN(new_n1034));
  NAND3_X1  g0834(.A1(new_n1033), .A2(new_n1034), .A3(new_n710), .ZN(new_n1035));
  NOR2_X1   g0835(.A1(new_n282), .A2(G50), .ZN(new_n1036));
  XNOR2_X1  g0836(.A(new_n1036), .B(KEYINPUT50), .ZN(new_n1037));
  AOI211_X1 g0837(.A(G45), .B(new_n711), .C1(G68), .C2(G77), .ZN(new_n1038));
  AOI21_X1  g0838(.A(new_n807), .B1(new_n1037), .B2(new_n1038), .ZN(new_n1039));
  OAI21_X1  g0839(.A(new_n1039), .B1(new_n233), .B2(new_n486), .ZN(new_n1040));
  NAND3_X1  g0840(.A1(new_n211), .A2(new_n249), .A3(new_n711), .ZN(new_n1041));
  OAI211_X1 g0841(.A(new_n1040), .B(new_n1041), .C1(G107), .C2(new_n211), .ZN(new_n1042));
  NAND2_X1  g0842(.A1(new_n1042), .A2(new_n810), .ZN(new_n1043));
  NAND2_X1  g0843(.A1(new_n1043), .A2(new_n756), .ZN(new_n1044));
  NOR3_X1   g0844(.A1(new_n703), .A2(G20), .A3(new_n758), .ZN(new_n1045));
  NAND2_X1  g0845(.A1(new_n558), .A2(new_n780), .ZN(new_n1046));
  OAI21_X1  g0846(.A(new_n1046), .B1(new_n774), .B2(new_n784), .ZN(new_n1047));
  XNOR2_X1  g0847(.A(new_n1047), .B(KEYINPUT114), .ZN(new_n1048));
  AOI22_X1  g0848(.A1(G77), .A2(new_n791), .B1(new_n1017), .B2(new_n309), .ZN(new_n1049));
  AOI22_X1  g0849(.A1(G68), .A2(new_n769), .B1(new_n796), .B2(G150), .ZN(new_n1050));
  AOI211_X1 g0850(.A(new_n347), .B(new_n1003), .C1(G159), .C2(new_n790), .ZN(new_n1051));
  NAND4_X1  g0851(.A1(new_n1048), .A2(new_n1049), .A3(new_n1050), .A4(new_n1051), .ZN(new_n1052));
  AOI22_X1  g0852(.A1(G116), .A2(new_n772), .B1(new_n796), .B2(G326), .ZN(new_n1053));
  OAI22_X1  g0853(.A1(new_n781), .A2(new_n823), .B1(new_n785), .B2(new_n535), .ZN(new_n1054));
  NOR2_X1   g0854(.A1(new_n768), .A2(new_n822), .ZN(new_n1055));
  INV_X1    g0855(.A(G317), .ZN(new_n1056));
  OAI22_X1  g0856(.A1(new_n793), .A2(new_n787), .B1(new_n784), .B2(new_n1056), .ZN(new_n1057));
  AOI211_X1 g0857(.A(new_n1055), .B(new_n1057), .C1(G322), .C2(new_n790), .ZN(new_n1058));
  AOI21_X1  g0858(.A(new_n1054), .B1(new_n1058), .B2(KEYINPUT48), .ZN(new_n1059));
  OAI21_X1  g0859(.A(new_n1059), .B1(KEYINPUT48), .B2(new_n1058), .ZN(new_n1060));
  INV_X1    g0860(.A(KEYINPUT49), .ZN(new_n1061));
  OAI211_X1 g0861(.A(new_n347), .B(new_n1053), .C1(new_n1060), .C2(new_n1061), .ZN(new_n1062));
  AND2_X1   g0862(.A1(new_n1060), .A2(new_n1061), .ZN(new_n1063));
  OAI21_X1  g0863(.A(new_n1052), .B1(new_n1062), .B2(new_n1063), .ZN(new_n1064));
  AOI211_X1 g0864(.A(new_n1044), .B(new_n1045), .C1(new_n802), .C2(new_n1064), .ZN(new_n1065));
  AOI21_X1  g0865(.A(new_n1065), .B1(new_n992), .B2(new_n997), .ZN(new_n1066));
  NAND2_X1  g0866(.A1(new_n1035), .A2(new_n1066), .ZN(G393));
  NAND2_X1  g0867(.A1(new_n990), .A2(new_n997), .ZN(new_n1068));
  NAND2_X1  g0868(.A1(new_n971), .A2(new_n759), .ZN(new_n1069));
  NAND2_X1  g0869(.A1(new_n1017), .A2(G50), .ZN(new_n1070));
  NAND2_X1  g0870(.A1(new_n780), .A2(G77), .ZN(new_n1071));
  NAND4_X1  g0871(.A1(new_n1070), .A2(new_n820), .A3(new_n1071), .A4(new_n329), .ZN(new_n1072));
  OAI22_X1  g0872(.A1(new_n777), .A2(new_n279), .B1(new_n784), .B2(new_n764), .ZN(new_n1073));
  XOR2_X1   g0873(.A(KEYINPUT115), .B(KEYINPUT51), .Z(new_n1074));
  OR2_X1    g0874(.A1(new_n1073), .A2(new_n1074), .ZN(new_n1075));
  NAND2_X1  g0875(.A1(new_n1073), .A2(new_n1074), .ZN(new_n1076));
  NAND2_X1  g0876(.A1(new_n769), .A2(new_n309), .ZN(new_n1077));
  AOI22_X1  g0877(.A1(G68), .A2(new_n791), .B1(new_n796), .B2(G143), .ZN(new_n1078));
  NAND4_X1  g0878(.A1(new_n1075), .A2(new_n1076), .A3(new_n1077), .A4(new_n1078), .ZN(new_n1079));
  OAI22_X1  g0879(.A1(new_n777), .A2(new_n1056), .B1(new_n784), .B2(new_n793), .ZN(new_n1080));
  XOR2_X1   g0880(.A(new_n1080), .B(KEYINPUT52), .Z(new_n1081));
  AOI22_X1  g0881(.A1(G283), .A2(new_n791), .B1(new_n769), .B2(G294), .ZN(new_n1082));
  AOI22_X1  g0882(.A1(G303), .A2(new_n1017), .B1(new_n796), .B2(G322), .ZN(new_n1083));
  NAND2_X1  g0883(.A1(new_n780), .A2(G116), .ZN(new_n1084));
  AOI21_X1  g0884(.A(new_n249), .B1(new_n772), .B2(G107), .ZN(new_n1085));
  NAND4_X1  g0885(.A1(new_n1082), .A2(new_n1083), .A3(new_n1084), .A4(new_n1085), .ZN(new_n1086));
  OAI22_X1  g0886(.A1(new_n1072), .A2(new_n1079), .B1(new_n1081), .B2(new_n1086), .ZN(new_n1087));
  NAND2_X1  g0887(.A1(new_n1087), .A2(new_n802), .ZN(new_n1088));
  OAI221_X1 g0888(.A(new_n809), .B1(new_n465), .B2(new_n211), .C1(new_n243), .C2(new_n807), .ZN(new_n1089));
  NAND4_X1  g0889(.A1(new_n1069), .A2(new_n756), .A3(new_n1088), .A4(new_n1089), .ZN(new_n1090));
  NAND2_X1  g0890(.A1(new_n1068), .A2(new_n1090), .ZN(new_n1091));
  AOI21_X1  g0891(.A(new_n709), .B1(new_n990), .B2(new_n994), .ZN(new_n1092));
  OAI21_X1  g0892(.A(new_n1033), .B1(new_n989), .B2(new_n987), .ZN(new_n1093));
  AOI21_X1  g0893(.A(new_n1091), .B1(new_n1092), .B2(new_n1093), .ZN(new_n1094));
  INV_X1    g0894(.A(new_n1094), .ZN(G390));
  AOI211_X1 g0895(.A(new_n582), .B(new_n691), .C1(new_n646), .C2(new_n654), .ZN(new_n1096));
  OAI211_X1 g0896(.A(G330), .B(new_n848), .C1(new_n1096), .C2(new_n743), .ZN(new_n1097));
  NAND2_X1  g0897(.A1(new_n1097), .A2(new_n923), .ZN(new_n1098));
  NOR2_X1   g0898(.A1(new_n845), .A2(new_n847), .ZN(new_n1099));
  AOI21_X1  g0899(.A(new_n913), .B1(new_n722), .B2(new_n1099), .ZN(new_n1100));
  AND2_X1   g0900(.A1(new_n1098), .A2(new_n1100), .ZN(new_n1101));
  AOI21_X1  g0901(.A(new_n697), .B1(new_n730), .B2(new_n744), .ZN(new_n1102));
  AOI21_X1  g0902(.A(KEYINPUT116), .B1(new_n1102), .B2(new_n936), .ZN(new_n1103));
  INV_X1    g0903(.A(KEYINPUT116), .ZN(new_n1104));
  NOR4_X1   g0904(.A1(new_n940), .A2(new_n1104), .A3(new_n697), .A4(new_n935), .ZN(new_n1105));
  NOR2_X1   g0905(.A1(new_n1103), .A2(new_n1105), .ZN(new_n1106));
  NAND2_X1  g0906(.A1(new_n1101), .A2(new_n1106), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n1102), .A2(new_n936), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n1098), .A2(new_n1108), .ZN(new_n1109));
  AOI21_X1  g0909(.A(KEYINPUT117), .B1(new_n1109), .B2(new_n915), .ZN(new_n1110));
  AOI22_X1  g0910(.A1(new_n1097), .A2(new_n923), .B1(new_n1102), .B2(new_n936), .ZN(new_n1111));
  INV_X1    g0911(.A(KEYINPUT117), .ZN(new_n1112));
  NOR3_X1   g0912(.A1(new_n1111), .A2(new_n1112), .A3(new_n914), .ZN(new_n1113));
  OAI21_X1  g0913(.A(new_n1107), .B1(new_n1110), .B2(new_n1113), .ZN(new_n1114));
  OAI211_X1 g0914(.A(new_n939), .B(new_n868), .C1(new_n923), .C2(new_n1100), .ZN(new_n1115));
  OAI21_X1  g0915(.A(new_n868), .B1(new_n914), .B2(new_n923), .ZN(new_n1116));
  NAND3_X1  g0916(.A1(new_n908), .A2(new_n911), .A3(new_n1116), .ZN(new_n1117));
  NAND2_X1  g0917(.A1(new_n1115), .A2(new_n1117), .ZN(new_n1118));
  INV_X1    g0918(.A(new_n1108), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n1118), .A2(new_n1119), .ZN(new_n1120));
  NAND3_X1  g0920(.A1(new_n1115), .A2(new_n1106), .A3(new_n1117), .ZN(new_n1121));
  AOI21_X1  g0921(.A(new_n930), .B1(G330), .B2(new_n932), .ZN(new_n1122));
  NAND4_X1  g0922(.A1(new_n1114), .A2(new_n1120), .A3(new_n1121), .A4(new_n1122), .ZN(new_n1123));
  OAI21_X1  g0923(.A(new_n1112), .B1(new_n1111), .B2(new_n914), .ZN(new_n1124));
  AOI21_X1  g0924(.A(new_n924), .B1(new_n1102), .B2(new_n848), .ZN(new_n1125));
  OAI211_X1 g0925(.A(KEYINPUT117), .B(new_n915), .C1(new_n1119), .C2(new_n1125), .ZN(new_n1126));
  AOI22_X1  g0926(.A1(new_n1124), .A2(new_n1126), .B1(new_n1106), .B2(new_n1101), .ZN(new_n1127));
  INV_X1    g0927(.A(new_n1122), .ZN(new_n1128));
  AND3_X1   g0928(.A1(new_n1115), .A2(new_n1106), .A3(new_n1117), .ZN(new_n1129));
  AOI21_X1  g0929(.A(new_n1108), .B1(new_n1115), .B2(new_n1117), .ZN(new_n1130));
  OAI22_X1  g0930(.A1(new_n1127), .A2(new_n1128), .B1(new_n1129), .B2(new_n1130), .ZN(new_n1131));
  NAND3_X1  g0931(.A1(new_n1123), .A2(new_n1131), .A3(new_n710), .ZN(new_n1132));
  INV_X1    g0932(.A(KEYINPUT118), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n1132), .A2(new_n1133), .ZN(new_n1134));
  NAND4_X1  g0934(.A1(new_n1123), .A2(new_n1131), .A3(KEYINPUT118), .A4(new_n710), .ZN(new_n1135));
  NOR2_X1   g0935(.A1(new_n1129), .A2(new_n1130), .ZN(new_n1136));
  NAND3_X1  g0936(.A1(new_n908), .A2(new_n757), .A3(new_n911), .ZN(new_n1137));
  OAI21_X1  g0937(.A(new_n756), .B1(new_n309), .B2(new_n817), .ZN(new_n1138));
  OAI22_X1  g0938(.A1(new_n777), .A2(new_n823), .B1(new_n771), .B2(new_n220), .ZN(new_n1139));
  AOI211_X1 g0939(.A(new_n249), .B(new_n1139), .C1(G87), .C2(new_n791), .ZN(new_n1140));
  AOI22_X1  g0940(.A1(G107), .A2(new_n1017), .B1(new_n798), .B2(G116), .ZN(new_n1141));
  AOI22_X1  g0941(.A1(G97), .A2(new_n769), .B1(new_n796), .B2(G294), .ZN(new_n1142));
  NAND4_X1  g0942(.A1(new_n1140), .A2(new_n1071), .A3(new_n1141), .A4(new_n1142), .ZN(new_n1143));
  OAI21_X1  g0943(.A(new_n249), .B1(new_n771), .B2(new_n774), .ZN(new_n1144));
  AOI21_X1  g0944(.A(new_n1144), .B1(G125), .B2(new_n796), .ZN(new_n1145));
  XNOR2_X1  g0945(.A(new_n1145), .B(KEYINPUT120), .ZN(new_n1146));
  XOR2_X1   g0946(.A(KEYINPUT121), .B(KEYINPUT53), .Z(new_n1147));
  AOI21_X1  g0947(.A(new_n1147), .B1(new_n791), .B2(G150), .ZN(new_n1148));
  AOI21_X1  g0948(.A(new_n1148), .B1(G159), .B2(new_n780), .ZN(new_n1149));
  NAND3_X1  g0949(.A1(new_n791), .A2(G150), .A3(new_n1147), .ZN(new_n1150));
  INV_X1    g0950(.A(G128), .ZN(new_n1151));
  OAI22_X1  g0951(.A1(new_n777), .A2(new_n1151), .B1(new_n784), .B2(new_n826), .ZN(new_n1152));
  AOI21_X1  g0952(.A(new_n1152), .B1(G137), .B2(new_n1017), .ZN(new_n1153));
  XNOR2_X1  g0953(.A(KEYINPUT54), .B(G143), .ZN(new_n1154));
  XNOR2_X1  g0954(.A(new_n1154), .B(KEYINPUT119), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n1155), .A2(new_n769), .ZN(new_n1156));
  NAND4_X1  g0956(.A1(new_n1149), .A2(new_n1150), .A3(new_n1153), .A4(new_n1156), .ZN(new_n1157));
  OAI21_X1  g0957(.A(new_n1143), .B1(new_n1146), .B2(new_n1157), .ZN(new_n1158));
  AOI21_X1  g0958(.A(new_n1138), .B1(new_n1158), .B2(new_n802), .ZN(new_n1159));
  AOI22_X1  g0959(.A1(new_n1136), .A2(new_n997), .B1(new_n1137), .B2(new_n1159), .ZN(new_n1160));
  NAND3_X1  g0960(.A1(new_n1134), .A2(new_n1135), .A3(new_n1160), .ZN(G378));
  AOI21_X1  g0961(.A(new_n1128), .B1(new_n1136), .B2(new_n1114), .ZN(new_n1162));
  XOR2_X1   g0962(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1163));
  INV_X1    g0963(.A(new_n1163), .ZN(new_n1164));
  OR2_X1    g0964(.A1(new_n308), .A2(new_n1164), .ZN(new_n1165));
  NAND2_X1  g0965(.A1(new_n308), .A2(new_n1164), .ZN(new_n1166));
  NAND2_X1  g0966(.A1(new_n1165), .A2(new_n1166), .ZN(new_n1167));
  NAND2_X1  g0967(.A1(new_n297), .A2(new_n881), .ZN(new_n1168));
  XOR2_X1   g0968(.A(new_n1168), .B(KEYINPUT125), .Z(new_n1169));
  INV_X1    g0969(.A(new_n1169), .ZN(new_n1170));
  NAND2_X1  g0970(.A1(new_n1167), .A2(new_n1170), .ZN(new_n1171));
  NAND3_X1  g0971(.A1(new_n1165), .A2(new_n1169), .A3(new_n1166), .ZN(new_n1172));
  NAND2_X1  g0972(.A1(new_n1171), .A2(new_n1172), .ZN(new_n1173));
  OAI211_X1 g0973(.A(new_n745), .B(new_n936), .C1(new_n909), .C2(new_n910), .ZN(new_n1174));
  AOI22_X1  g0974(.A1(new_n934), .A2(new_n1174), .B1(new_n939), .B2(new_n941), .ZN(new_n1175));
  AOI21_X1  g0975(.A(new_n1173), .B1(new_n1175), .B2(G330), .ZN(new_n1176));
  AND4_X1   g0976(.A1(G330), .A2(new_n938), .A3(new_n942), .A4(new_n1173), .ZN(new_n1177));
  OAI21_X1  g0977(.A(new_n928), .B1(new_n1176), .B2(new_n1177), .ZN(new_n1178));
  INV_X1    g0978(.A(new_n1173), .ZN(new_n1179));
  OAI21_X1  g0979(.A(new_n1179), .B1(new_n943), .B2(new_n697), .ZN(new_n1180));
  NOR2_X1   g0980(.A1(new_n912), .A2(new_n927), .ZN(new_n1181));
  NAND3_X1  g0981(.A1(new_n1175), .A2(G330), .A3(new_n1173), .ZN(new_n1182));
  NAND3_X1  g0982(.A1(new_n1180), .A2(new_n1181), .A3(new_n1182), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n1178), .A2(new_n1183), .ZN(new_n1184));
  OAI21_X1  g0984(.A(KEYINPUT57), .B1(new_n1162), .B2(new_n1184), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n1120), .A2(new_n1121), .ZN(new_n1186));
  OAI21_X1  g0986(.A(new_n1122), .B1(new_n1186), .B2(new_n1127), .ZN(new_n1187));
  INV_X1    g0987(.A(KEYINPUT57), .ZN(new_n1188));
  NAND4_X1  g0988(.A1(new_n1187), .A2(new_n1188), .A3(new_n1183), .A4(new_n1178), .ZN(new_n1189));
  AOI21_X1  g0989(.A(new_n709), .B1(new_n1185), .B2(new_n1189), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n1173), .A2(new_n757), .ZN(new_n1191));
  OAI21_X1  g0991(.A(new_n756), .B1(G50), .B2(new_n817), .ZN(new_n1192));
  NOR2_X1   g0992(.A1(new_n329), .A2(G41), .ZN(new_n1193));
  AOI211_X1 g0993(.A(G50), .B(new_n1193), .C1(new_n245), .C2(new_n708), .ZN(new_n1194));
  OAI22_X1  g0994(.A1(new_n768), .A2(new_n435), .B1(new_n763), .B2(new_n823), .ZN(new_n1195));
  INV_X1    g0995(.A(new_n1195), .ZN(new_n1196));
  OAI211_X1 g0996(.A(new_n1196), .B(new_n1193), .C1(new_n465), .C2(new_n787), .ZN(new_n1197));
  OAI22_X1  g0997(.A1(new_n785), .A2(new_n253), .B1(new_n771), .B2(new_n783), .ZN(new_n1198));
  OAI22_X1  g0998(.A1(new_n777), .A2(new_n603), .B1(new_n784), .B2(new_n444), .ZN(new_n1199));
  NOR4_X1   g0999(.A1(new_n1197), .A2(new_n1014), .A3(new_n1198), .A4(new_n1199), .ZN(new_n1200));
  XNOR2_X1  g1000(.A(new_n1200), .B(KEYINPUT122), .ZN(new_n1201));
  XNOR2_X1  g1001(.A(KEYINPUT123), .B(KEYINPUT58), .ZN(new_n1202));
  AOI21_X1  g1002(.A(new_n1194), .B1(new_n1201), .B2(new_n1202), .ZN(new_n1203));
  AOI22_X1  g1003(.A1(G125), .A2(new_n790), .B1(new_n1017), .B2(G132), .ZN(new_n1204));
  OAI221_X1 g1004(.A(new_n1204), .B1(new_n828), .B2(new_n768), .C1(new_n279), .C2(new_n781), .ZN(new_n1205));
  AOI22_X1  g1005(.A1(new_n1155), .A2(new_n791), .B1(G128), .B2(new_n798), .ZN(new_n1206));
  OR2_X1    g1006(.A1(new_n1206), .A2(KEYINPUT124), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n1206), .A2(KEYINPUT124), .ZN(new_n1208));
  AOI21_X1  g1008(.A(new_n1205), .B1(new_n1207), .B2(new_n1208), .ZN(new_n1209));
  INV_X1    g1009(.A(KEYINPUT59), .ZN(new_n1210));
  AND2_X1   g1010(.A1(new_n1209), .A2(new_n1210), .ZN(new_n1211));
  OAI211_X1 g1011(.A(new_n245), .B(new_n708), .C1(new_n771), .C2(new_n764), .ZN(new_n1212));
  AOI21_X1  g1012(.A(new_n1212), .B1(G124), .B2(new_n796), .ZN(new_n1213));
  OAI21_X1  g1013(.A(new_n1213), .B1(new_n1209), .B2(new_n1210), .ZN(new_n1214));
  OAI221_X1 g1014(.A(new_n1203), .B1(new_n1211), .B2(new_n1214), .C1(new_n1201), .C2(new_n1202), .ZN(new_n1215));
  AOI21_X1  g1015(.A(new_n1192), .B1(new_n1215), .B2(new_n802), .ZN(new_n1216));
  NAND2_X1  g1016(.A1(new_n1191), .A2(new_n1216), .ZN(new_n1217));
  INV_X1    g1017(.A(new_n997), .ZN(new_n1218));
  OAI21_X1  g1018(.A(new_n1217), .B1(new_n1184), .B2(new_n1218), .ZN(new_n1219));
  NOR2_X1   g1019(.A1(new_n1190), .A2(new_n1219), .ZN(new_n1220));
  INV_X1    g1020(.A(new_n1220), .ZN(G375));
  INV_X1    g1021(.A(KEYINPUT126), .ZN(new_n1222));
  OAI21_X1  g1022(.A(new_n1222), .B1(new_n1114), .B2(new_n1122), .ZN(new_n1223));
  INV_X1    g1023(.A(new_n979), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(new_n1114), .A2(new_n1122), .ZN(new_n1225));
  NAND3_X1  g1025(.A1(new_n1127), .A2(new_n1128), .A3(KEYINPUT126), .ZN(new_n1226));
  NAND4_X1  g1026(.A1(new_n1223), .A2(new_n1224), .A3(new_n1225), .A4(new_n1226), .ZN(new_n1227));
  INV_X1    g1027(.A(KEYINPUT127), .ZN(new_n1228));
  OR2_X1    g1028(.A1(new_n1227), .A2(new_n1228), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n1227), .A2(new_n1228), .ZN(new_n1230));
  NAND2_X1  g1030(.A1(new_n923), .A2(new_n757), .ZN(new_n1231));
  OAI21_X1  g1031(.A(new_n756), .B1(G68), .B2(new_n817), .ZN(new_n1232));
  AOI22_X1  g1032(.A1(G97), .A2(new_n791), .B1(new_n796), .B2(G303), .ZN(new_n1233));
  OAI221_X1 g1033(.A(new_n1233), .B1(new_n444), .B2(new_n768), .C1(new_n535), .C2(new_n777), .ZN(new_n1234));
  AOI22_X1  g1034(.A1(G116), .A2(new_n1017), .B1(new_n798), .B2(G283), .ZN(new_n1235));
  NAND4_X1  g1035(.A1(new_n1235), .A2(new_n446), .A3(new_n1012), .A4(new_n1046), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n1155), .A2(new_n1017), .ZN(new_n1237));
  AOI22_X1  g1037(.A1(G137), .A2(new_n798), .B1(new_n769), .B2(G150), .ZN(new_n1238));
  AOI22_X1  g1038(.A1(G132), .A2(new_n790), .B1(new_n791), .B2(G159), .ZN(new_n1239));
  NAND3_X1  g1039(.A1(new_n1237), .A2(new_n1238), .A3(new_n1239), .ZN(new_n1240));
  AOI22_X1  g1040(.A1(G58), .A2(new_n772), .B1(new_n796), .B2(G128), .ZN(new_n1241));
  OAI211_X1 g1041(.A(new_n1241), .B(new_n329), .C1(new_n774), .C2(new_n781), .ZN(new_n1242));
  OAI22_X1  g1042(.A1(new_n1234), .A2(new_n1236), .B1(new_n1240), .B2(new_n1242), .ZN(new_n1243));
  AOI21_X1  g1043(.A(new_n1232), .B1(new_n1243), .B2(new_n802), .ZN(new_n1244));
  AOI22_X1  g1044(.A1(new_n1114), .A2(new_n997), .B1(new_n1231), .B2(new_n1244), .ZN(new_n1245));
  NAND3_X1  g1045(.A1(new_n1229), .A2(new_n1230), .A3(new_n1245), .ZN(G381));
  NAND2_X1  g1046(.A1(new_n1132), .A2(new_n1160), .ZN(new_n1247));
  NOR2_X1   g1047(.A1(G375), .A2(new_n1247), .ZN(new_n1248));
  NAND3_X1  g1048(.A1(new_n998), .A2(new_n1031), .A3(new_n1094), .ZN(new_n1249));
  NAND3_X1  g1049(.A1(new_n1035), .A2(new_n814), .A3(new_n1066), .ZN(new_n1250));
  NOR4_X1   g1050(.A1(G381), .A2(G384), .A3(new_n1249), .A4(new_n1250), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n1248), .A2(new_n1251), .ZN(G407));
  INV_X1    g1052(.A(G213), .ZN(new_n1253));
  NOR2_X1   g1053(.A1(new_n1253), .A2(G343), .ZN(new_n1254));
  NAND2_X1  g1054(.A1(new_n1248), .A2(new_n1254), .ZN(new_n1255));
  NAND3_X1  g1055(.A1(G407), .A2(new_n1255), .A3(G213), .ZN(G409));
  INV_X1    g1056(.A(new_n1254), .ZN(new_n1257));
  OAI21_X1  g1057(.A(KEYINPUT60), .B1(new_n1127), .B2(new_n1128), .ZN(new_n1258));
  NAND3_X1  g1058(.A1(new_n1223), .A2(new_n1258), .A3(new_n1226), .ZN(new_n1259));
  NOR2_X1   g1059(.A1(new_n1114), .A2(new_n1122), .ZN(new_n1260));
  AOI21_X1  g1060(.A(new_n709), .B1(new_n1260), .B2(KEYINPUT60), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(new_n1259), .A2(new_n1261), .ZN(new_n1262));
  AOI21_X1  g1062(.A(G384), .B1(new_n1262), .B2(new_n1245), .ZN(new_n1263));
  INV_X1    g1063(.A(new_n1245), .ZN(new_n1264));
  AOI211_X1 g1064(.A(new_n856), .B(new_n1264), .C1(new_n1259), .C2(new_n1261), .ZN(new_n1265));
  NOR2_X1   g1065(.A1(new_n1263), .A2(new_n1265), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(new_n1135), .A2(new_n1160), .ZN(new_n1267));
  AOI21_X1  g1067(.A(new_n709), .B1(new_n1225), .B2(new_n1186), .ZN(new_n1268));
  AOI21_X1  g1068(.A(KEYINPUT118), .B1(new_n1268), .B2(new_n1123), .ZN(new_n1269));
  NOR2_X1   g1069(.A1(new_n1267), .A2(new_n1269), .ZN(new_n1270));
  NOR3_X1   g1070(.A1(new_n1270), .A2(new_n1190), .A3(new_n1219), .ZN(new_n1271));
  INV_X1    g1071(.A(new_n1219), .ZN(new_n1272));
  NAND4_X1  g1072(.A1(new_n1187), .A2(new_n1224), .A3(new_n1183), .A4(new_n1178), .ZN(new_n1273));
  AOI21_X1  g1073(.A(new_n1247), .B1(new_n1272), .B2(new_n1273), .ZN(new_n1274));
  OAI211_X1 g1074(.A(new_n1257), .B(new_n1266), .C1(new_n1271), .C2(new_n1274), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(new_n1275), .A2(KEYINPUT62), .ZN(new_n1276));
  INV_X1    g1076(.A(KEYINPUT61), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(new_n1262), .A2(new_n1245), .ZN(new_n1278));
  NAND2_X1  g1078(.A1(new_n1278), .A2(new_n856), .ZN(new_n1279));
  NAND3_X1  g1079(.A1(new_n1262), .A2(G384), .A3(new_n1245), .ZN(new_n1280));
  NAND2_X1  g1080(.A1(new_n1254), .A2(G2897), .ZN(new_n1281));
  NAND3_X1  g1081(.A1(new_n1279), .A2(new_n1280), .A3(new_n1281), .ZN(new_n1282));
  INV_X1    g1082(.A(new_n1281), .ZN(new_n1283));
  OAI21_X1  g1083(.A(new_n1283), .B1(new_n1263), .B2(new_n1265), .ZN(new_n1284));
  AOI21_X1  g1084(.A(new_n1274), .B1(new_n1220), .B2(G378), .ZN(new_n1285));
  OAI211_X1 g1085(.A(new_n1282), .B(new_n1284), .C1(new_n1285), .C2(new_n1254), .ZN(new_n1286));
  AND2_X1   g1086(.A1(new_n1185), .A2(new_n1189), .ZN(new_n1287));
  OAI211_X1 g1087(.A(G378), .B(new_n1272), .C1(new_n1287), .C2(new_n709), .ZN(new_n1288));
  INV_X1    g1088(.A(new_n1274), .ZN(new_n1289));
  NAND2_X1  g1089(.A1(new_n1288), .A2(new_n1289), .ZN(new_n1290));
  INV_X1    g1090(.A(KEYINPUT62), .ZN(new_n1291));
  NAND4_X1  g1091(.A1(new_n1290), .A2(new_n1291), .A3(new_n1257), .A4(new_n1266), .ZN(new_n1292));
  NAND4_X1  g1092(.A1(new_n1276), .A2(new_n1277), .A3(new_n1286), .A4(new_n1292), .ZN(new_n1293));
  NAND2_X1  g1093(.A1(G393), .A2(G396), .ZN(new_n1294));
  NAND2_X1  g1094(.A1(new_n1294), .A2(new_n1250), .ZN(new_n1295));
  INV_X1    g1095(.A(new_n1295), .ZN(new_n1296));
  INV_X1    g1096(.A(new_n1249), .ZN(new_n1297));
  AOI21_X1  g1097(.A(new_n1094), .B1(new_n998), .B2(new_n1031), .ZN(new_n1298));
  OAI21_X1  g1098(.A(new_n1296), .B1(new_n1297), .B2(new_n1298), .ZN(new_n1299));
  NAND2_X1  g1099(.A1(G387), .A2(G390), .ZN(new_n1300));
  NAND3_X1  g1100(.A1(new_n1300), .A2(new_n1249), .A3(new_n1295), .ZN(new_n1301));
  NAND2_X1  g1101(.A1(new_n1299), .A2(new_n1301), .ZN(new_n1302));
  NAND2_X1  g1102(.A1(new_n1293), .A2(new_n1302), .ZN(new_n1303));
  AOI21_X1  g1103(.A(new_n1254), .B1(new_n1288), .B2(new_n1289), .ZN(new_n1304));
  NAND2_X1  g1104(.A1(new_n1282), .A2(new_n1284), .ZN(new_n1305));
  OAI21_X1  g1105(.A(KEYINPUT63), .B1(new_n1304), .B2(new_n1305), .ZN(new_n1306));
  NAND2_X1  g1106(.A1(new_n1306), .A2(new_n1275), .ZN(new_n1307));
  NAND3_X1  g1107(.A1(new_n1304), .A2(KEYINPUT63), .A3(new_n1266), .ZN(new_n1308));
  NOR2_X1   g1108(.A1(new_n1302), .A2(KEYINPUT61), .ZN(new_n1309));
  NAND3_X1  g1109(.A1(new_n1307), .A2(new_n1308), .A3(new_n1309), .ZN(new_n1310));
  NAND2_X1  g1110(.A1(new_n1303), .A2(new_n1310), .ZN(G405));
  XNOR2_X1  g1111(.A(new_n1302), .B(new_n1266), .ZN(new_n1312));
  OAI21_X1  g1112(.A(new_n1288), .B1(new_n1220), .B2(new_n1247), .ZN(new_n1313));
  XNOR2_X1  g1113(.A(new_n1312), .B(new_n1313), .ZN(G402));
endmodule


