//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 0 0 0 1 1 0 0 1 0 1 1 0 1 1 0 1 1 1 1 1 1 0 0 0 1 0 0 1 1 0 0 1 0 1 1 1 0 1 1 0 0 1 0 0 1 1 1 1 0 1 1 0 1 0 1 0 1 0 0 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:20:51 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n670, new_n671, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n692, new_n693, new_n694, new_n695, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n704, new_n705,
    new_n706, new_n708, new_n709, new_n710, new_n711, new_n712, new_n714,
    new_n715, new_n716, new_n717, new_n718, new_n719, new_n721, new_n722,
    new_n723, new_n725, new_n727, new_n728, new_n729, new_n730, new_n731,
    new_n732, new_n733, new_n734, new_n735, new_n736, new_n737, new_n738,
    new_n739, new_n740, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n844, new_n845, new_n846, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n854, new_n856, new_n857,
    new_n858, new_n859, new_n860, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n919, new_n920, new_n922, new_n923, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n937, new_n938, new_n940, new_n941,
    new_n942, new_n944, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n951, new_n952, new_n954, new_n955, new_n956, new_n957,
    new_n958, new_n959, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n974, new_n975, new_n976, new_n977, new_n978, new_n980, new_n981;
  XOR2_X1   g000(.A(G197gat), .B(G204gat), .Z(new_n202));
  INV_X1    g001(.A(new_n202), .ZN(new_n203));
  XNOR2_X1  g002(.A(G211gat), .B(G218gat), .ZN(new_n204));
  XNOR2_X1  g003(.A(KEYINPUT73), .B(G218gat), .ZN(new_n205));
  AND2_X1   g004(.A1(new_n205), .A2(G211gat), .ZN(new_n206));
  OAI211_X1 g005(.A(new_n203), .B(new_n204), .C1(new_n206), .C2(KEYINPUT22), .ZN(new_n207));
  INV_X1    g006(.A(new_n204), .ZN(new_n208));
  AOI21_X1  g007(.A(KEYINPUT22), .B1(new_n205), .B2(G211gat), .ZN(new_n209));
  OAI21_X1  g008(.A(new_n208), .B1(new_n209), .B2(new_n202), .ZN(new_n210));
  NAND2_X1  g009(.A1(new_n207), .A2(new_n210), .ZN(new_n211));
  INV_X1    g010(.A(new_n211), .ZN(new_n212));
  INV_X1    g011(.A(G226gat), .ZN(new_n213));
  INV_X1    g012(.A(G233gat), .ZN(new_n214));
  NOR2_X1   g013(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  INV_X1    g014(.A(G183gat), .ZN(new_n216));
  OAI21_X1  g015(.A(KEYINPUT27), .B1(new_n216), .B2(KEYINPUT66), .ZN(new_n217));
  INV_X1    g016(.A(G190gat), .ZN(new_n218));
  INV_X1    g017(.A(KEYINPUT27), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n219), .A2(G183gat), .ZN(new_n220));
  OAI211_X1 g019(.A(new_n217), .B(new_n218), .C1(KEYINPUT66), .C2(new_n220), .ZN(new_n221));
  XNOR2_X1  g020(.A(KEYINPUT67), .B(KEYINPUT28), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  XNOR2_X1  g022(.A(KEYINPUT27), .B(G183gat), .ZN(new_n224));
  NAND3_X1  g023(.A1(new_n224), .A2(KEYINPUT28), .A3(new_n218), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n223), .A2(new_n225), .ZN(new_n226));
  INV_X1    g025(.A(G169gat), .ZN(new_n227));
  INV_X1    g026(.A(G176gat), .ZN(new_n228));
  NOR2_X1   g027(.A1(new_n227), .A2(new_n228), .ZN(new_n229));
  NOR2_X1   g028(.A1(G169gat), .A2(G176gat), .ZN(new_n230));
  NOR3_X1   g029(.A1(new_n229), .A2(KEYINPUT26), .A3(new_n230), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n230), .A2(KEYINPUT26), .ZN(new_n232));
  NAND2_X1  g031(.A1(G183gat), .A2(G190gat), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n232), .A2(new_n233), .ZN(new_n234));
  NOR2_X1   g033(.A1(new_n231), .A2(new_n234), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n226), .A2(new_n235), .ZN(new_n236));
  INV_X1    g035(.A(KEYINPUT25), .ZN(new_n237));
  AOI22_X1  g036(.A1(new_n237), .A2(KEYINPUT65), .B1(G169gat), .B2(G176gat), .ZN(new_n238));
  NAND3_X1  g037(.A1(new_n227), .A2(new_n228), .A3(KEYINPUT23), .ZN(new_n239));
  INV_X1    g038(.A(KEYINPUT23), .ZN(new_n240));
  OAI21_X1  g039(.A(new_n240), .B1(G169gat), .B2(G176gat), .ZN(new_n241));
  INV_X1    g040(.A(KEYINPUT24), .ZN(new_n242));
  NAND3_X1  g041(.A1(new_n242), .A2(G183gat), .A3(G190gat), .ZN(new_n243));
  NAND4_X1  g042(.A1(new_n238), .A2(new_n239), .A3(new_n241), .A4(new_n243), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n216), .A2(new_n218), .ZN(new_n245));
  AND3_X1   g044(.A1(new_n245), .A2(KEYINPUT24), .A3(new_n233), .ZN(new_n246));
  OAI22_X1  g045(.A1(new_n244), .A2(new_n246), .B1(KEYINPUT65), .B2(new_n237), .ZN(new_n247));
  AND2_X1   g046(.A1(new_n238), .A2(new_n243), .ZN(new_n248));
  AND2_X1   g047(.A1(new_n239), .A2(new_n241), .ZN(new_n249));
  NOR2_X1   g048(.A1(new_n237), .A2(KEYINPUT65), .ZN(new_n250));
  NAND3_X1  g049(.A1(new_n245), .A2(KEYINPUT24), .A3(new_n233), .ZN(new_n251));
  NAND4_X1  g050(.A1(new_n248), .A2(new_n249), .A3(new_n250), .A4(new_n251), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n247), .A2(new_n252), .ZN(new_n253));
  NAND2_X1  g052(.A1(new_n236), .A2(new_n253), .ZN(new_n254));
  INV_X1    g053(.A(KEYINPUT29), .ZN(new_n255));
  AOI21_X1  g054(.A(new_n215), .B1(new_n254), .B2(new_n255), .ZN(new_n256));
  AOI22_X1  g055(.A1(new_n226), .A2(new_n235), .B1(new_n247), .B2(new_n252), .ZN(new_n257));
  NOR3_X1   g056(.A1(new_n257), .A2(new_n213), .A3(new_n214), .ZN(new_n258));
  OAI21_X1  g057(.A(new_n212), .B1(new_n256), .B2(new_n258), .ZN(new_n259));
  XNOR2_X1  g058(.A(G8gat), .B(G36gat), .ZN(new_n260));
  XNOR2_X1  g059(.A(G64gat), .B(G92gat), .ZN(new_n261));
  XOR2_X1   g060(.A(new_n260), .B(new_n261), .Z(new_n262));
  OAI22_X1  g061(.A1(new_n257), .A2(KEYINPUT29), .B1(new_n213), .B2(new_n214), .ZN(new_n263));
  NAND2_X1  g062(.A1(new_n254), .A2(new_n215), .ZN(new_n264));
  NAND3_X1  g063(.A1(new_n263), .A2(new_n211), .A3(new_n264), .ZN(new_n265));
  NAND3_X1  g064(.A1(new_n259), .A2(new_n262), .A3(new_n265), .ZN(new_n266));
  INV_X1    g065(.A(KEYINPUT30), .ZN(new_n267));
  NAND2_X1  g066(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  INV_X1    g067(.A(new_n262), .ZN(new_n269));
  INV_X1    g068(.A(new_n265), .ZN(new_n270));
  AOI21_X1  g069(.A(new_n211), .B1(new_n263), .B2(new_n264), .ZN(new_n271));
  OAI21_X1  g070(.A(new_n269), .B1(new_n270), .B2(new_n271), .ZN(new_n272));
  NAND4_X1  g071(.A1(new_n259), .A2(KEYINPUT30), .A3(new_n265), .A4(new_n262), .ZN(new_n273));
  NAND3_X1  g072(.A1(new_n268), .A2(new_n272), .A3(new_n273), .ZN(new_n274));
  OR2_X1    g073(.A1(new_n274), .A2(KEYINPUT35), .ZN(new_n275));
  AND2_X1   g074(.A1(new_n226), .A2(new_n235), .ZN(new_n276));
  AND2_X1   g075(.A1(new_n247), .A2(new_n252), .ZN(new_n277));
  INV_X1    g076(.A(G127gat), .ZN(new_n278));
  OAI21_X1  g077(.A(KEYINPUT68), .B1(new_n278), .B2(G134gat), .ZN(new_n279));
  XNOR2_X1  g078(.A(G113gat), .B(G120gat), .ZN(new_n280));
  OAI21_X1  g079(.A(new_n279), .B1(new_n280), .B2(KEYINPUT1), .ZN(new_n281));
  XNOR2_X1  g080(.A(G127gat), .B(G134gat), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  INV_X1    g082(.A(new_n282), .ZN(new_n284));
  OAI211_X1 g083(.A(new_n284), .B(new_n279), .C1(KEYINPUT1), .C2(new_n280), .ZN(new_n285));
  AND3_X1   g084(.A1(new_n283), .A2(new_n285), .A3(KEYINPUT69), .ZN(new_n286));
  AOI21_X1  g085(.A(KEYINPUT69), .B1(new_n283), .B2(new_n285), .ZN(new_n287));
  OAI22_X1  g086(.A1(new_n276), .A2(new_n277), .B1(new_n286), .B2(new_n287), .ZN(new_n288));
  NAND3_X1  g087(.A1(new_n283), .A2(new_n285), .A3(KEYINPUT69), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n283), .A2(new_n285), .ZN(new_n290));
  INV_X1    g089(.A(KEYINPUT69), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  NAND3_X1  g091(.A1(new_n257), .A2(new_n289), .A3(new_n292), .ZN(new_n293));
  NAND2_X1  g092(.A1(G227gat), .A2(G233gat), .ZN(new_n294));
  XNOR2_X1  g093(.A(new_n294), .B(KEYINPUT64), .ZN(new_n295));
  NAND3_X1  g094(.A1(new_n288), .A2(new_n293), .A3(new_n295), .ZN(new_n296));
  AND2_X1   g095(.A1(new_n296), .A2(KEYINPUT32), .ZN(new_n297));
  INV_X1    g096(.A(new_n294), .ZN(new_n298));
  AOI21_X1  g097(.A(new_n298), .B1(new_n288), .B2(new_n293), .ZN(new_n299));
  XOR2_X1   g098(.A(KEYINPUT70), .B(KEYINPUT34), .Z(new_n300));
  NOR2_X1   g099(.A1(new_n299), .A2(new_n300), .ZN(new_n301));
  AOI211_X1 g100(.A(KEYINPUT34), .B(new_n295), .C1(new_n288), .C2(new_n293), .ZN(new_n302));
  OAI21_X1  g101(.A(new_n297), .B1(new_n301), .B2(new_n302), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n296), .A2(KEYINPUT32), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n288), .A2(new_n293), .ZN(new_n305));
  INV_X1    g104(.A(KEYINPUT34), .ZN(new_n306));
  INV_X1    g105(.A(new_n295), .ZN(new_n307));
  NAND3_X1  g106(.A1(new_n305), .A2(new_n306), .A3(new_n307), .ZN(new_n308));
  OAI211_X1 g107(.A(new_n304), .B(new_n308), .C1(new_n299), .C2(new_n300), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n303), .A2(new_n309), .ZN(new_n310));
  INV_X1    g109(.A(KEYINPUT71), .ZN(new_n311));
  INV_X1    g110(.A(KEYINPUT33), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n296), .A2(new_n312), .ZN(new_n313));
  XOR2_X1   g112(.A(G15gat), .B(G43gat), .Z(new_n314));
  XNOR2_X1  g113(.A(G71gat), .B(G99gat), .ZN(new_n315));
  XNOR2_X1  g114(.A(new_n314), .B(new_n315), .ZN(new_n316));
  AOI21_X1  g115(.A(new_n311), .B1(new_n313), .B2(new_n316), .ZN(new_n317));
  INV_X1    g116(.A(new_n316), .ZN(new_n318));
  AOI211_X1 g117(.A(KEYINPUT71), .B(new_n318), .C1(new_n296), .C2(new_n312), .ZN(new_n319));
  NOR2_X1   g118(.A1(new_n317), .A2(new_n319), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n310), .A2(new_n320), .ZN(new_n321));
  OAI211_X1 g120(.A(new_n303), .B(new_n309), .C1(new_n317), .C2(new_n319), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  INV_X1    g122(.A(G155gat), .ZN(new_n324));
  INV_X1    g123(.A(G162gat), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n324), .A2(new_n325), .ZN(new_n326));
  NAND2_X1  g125(.A1(G155gat), .A2(G162gat), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n326), .A2(new_n327), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n328), .A2(KEYINPUT75), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n327), .A2(KEYINPUT2), .ZN(new_n330));
  INV_X1    g129(.A(G141gat), .ZN(new_n331));
  INV_X1    g130(.A(G148gat), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n331), .A2(new_n332), .ZN(new_n333));
  NAND2_X1  g132(.A1(G141gat), .A2(G148gat), .ZN(new_n334));
  NAND3_X1  g133(.A1(new_n330), .A2(new_n333), .A3(new_n334), .ZN(new_n335));
  INV_X1    g134(.A(KEYINPUT75), .ZN(new_n336));
  NAND3_X1  g135(.A1(new_n326), .A2(new_n336), .A3(new_n327), .ZN(new_n337));
  NAND3_X1  g136(.A1(new_n329), .A2(new_n335), .A3(new_n337), .ZN(new_n338));
  AND2_X1   g137(.A1(new_n333), .A2(new_n334), .ZN(new_n339));
  INV_X1    g138(.A(KEYINPUT76), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n330), .A2(new_n340), .ZN(new_n341));
  NAND3_X1  g140(.A1(new_n327), .A2(KEYINPUT76), .A3(KEYINPUT2), .ZN(new_n342));
  NAND4_X1  g141(.A1(new_n339), .A2(new_n328), .A3(new_n341), .A4(new_n342), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n338), .A2(new_n343), .ZN(new_n344));
  AOI21_X1  g143(.A(KEYINPUT29), .B1(new_n207), .B2(new_n210), .ZN(new_n345));
  OAI21_X1  g144(.A(new_n344), .B1(new_n345), .B2(KEYINPUT3), .ZN(new_n346));
  INV_X1    g145(.A(G228gat), .ZN(new_n347));
  NOR2_X1   g146(.A1(new_n347), .A2(new_n214), .ZN(new_n348));
  INV_X1    g147(.A(KEYINPUT3), .ZN(new_n349));
  NAND3_X1  g148(.A1(new_n338), .A2(new_n343), .A3(new_n349), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n350), .A2(new_n255), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n212), .A2(new_n351), .ZN(new_n352));
  NAND3_X1  g151(.A1(new_n346), .A2(new_n348), .A3(new_n352), .ZN(new_n353));
  INV_X1    g152(.A(new_n353), .ZN(new_n354));
  AOI21_X1  g153(.A(new_n348), .B1(new_n346), .B2(new_n352), .ZN(new_n355));
  OAI21_X1  g154(.A(KEYINPUT78), .B1(new_n354), .B2(new_n355), .ZN(new_n356));
  INV_X1    g155(.A(new_n348), .ZN(new_n357));
  INV_X1    g156(.A(new_n344), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n211), .A2(new_n255), .ZN(new_n359));
  AOI21_X1  g158(.A(new_n358), .B1(new_n359), .B2(new_n349), .ZN(new_n360));
  AOI21_X1  g159(.A(new_n211), .B1(new_n255), .B2(new_n350), .ZN(new_n361));
  OAI21_X1  g160(.A(new_n357), .B1(new_n360), .B2(new_n361), .ZN(new_n362));
  INV_X1    g161(.A(KEYINPUT78), .ZN(new_n363));
  NAND3_X1  g162(.A1(new_n362), .A2(new_n353), .A3(new_n363), .ZN(new_n364));
  NAND3_X1  g163(.A1(new_n356), .A2(G22gat), .A3(new_n364), .ZN(new_n365));
  XNOR2_X1  g164(.A(G78gat), .B(G106gat), .ZN(new_n366));
  XNOR2_X1  g165(.A(KEYINPUT31), .B(G50gat), .ZN(new_n367));
  XOR2_X1   g166(.A(new_n366), .B(new_n367), .Z(new_n368));
  INV_X1    g167(.A(new_n368), .ZN(new_n369));
  AOI21_X1  g168(.A(new_n363), .B1(new_n362), .B2(new_n353), .ZN(new_n370));
  INV_X1    g169(.A(G22gat), .ZN(new_n371));
  AOI21_X1  g170(.A(new_n369), .B1(new_n370), .B2(new_n371), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n362), .A2(new_n353), .ZN(new_n373));
  AND2_X1   g172(.A1(KEYINPUT79), .A2(G22gat), .ZN(new_n374));
  OR2_X1    g173(.A1(new_n373), .A2(new_n374), .ZN(new_n375));
  AOI21_X1  g174(.A(new_n368), .B1(new_n373), .B2(new_n374), .ZN(new_n376));
  AOI22_X1  g175(.A1(new_n365), .A2(new_n372), .B1(new_n375), .B2(new_n376), .ZN(new_n377));
  INV_X1    g176(.A(KEYINPUT6), .ZN(new_n378));
  XOR2_X1   g177(.A(G1gat), .B(G29gat), .Z(new_n379));
  XNOR2_X1  g178(.A(new_n379), .B(KEYINPUT0), .ZN(new_n380));
  XNOR2_X1  g179(.A(G57gat), .B(G85gat), .ZN(new_n381));
  XNOR2_X1  g180(.A(new_n380), .B(new_n381), .ZN(new_n382));
  OAI211_X1 g181(.A(KEYINPUT4), .B(new_n358), .C1(new_n286), .C2(new_n287), .ZN(new_n383));
  AOI21_X1  g182(.A(new_n349), .B1(new_n338), .B2(new_n343), .ZN(new_n384));
  INV_X1    g183(.A(new_n384), .ZN(new_n385));
  NAND3_X1  g184(.A1(new_n385), .A2(new_n290), .A3(new_n350), .ZN(new_n386));
  NAND2_X1  g185(.A1(G225gat), .A2(G233gat), .ZN(new_n387));
  NAND4_X1  g186(.A1(new_n283), .A2(new_n285), .A3(new_n338), .A4(new_n343), .ZN(new_n388));
  INV_X1    g187(.A(KEYINPUT4), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n388), .A2(new_n389), .ZN(new_n390));
  NAND4_X1  g189(.A1(new_n383), .A2(new_n386), .A3(new_n387), .A4(new_n390), .ZN(new_n391));
  INV_X1    g190(.A(KEYINPUT5), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n290), .A2(new_n344), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n393), .A2(new_n388), .ZN(new_n394));
  INV_X1    g193(.A(new_n387), .ZN(new_n395));
  AOI21_X1  g194(.A(new_n392), .B1(new_n394), .B2(new_n395), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n391), .A2(new_n396), .ZN(new_n397));
  NOR2_X1   g196(.A1(new_n388), .A2(new_n389), .ZN(new_n398));
  OAI21_X1  g197(.A(new_n358), .B1(new_n286), .B2(new_n287), .ZN(new_n399));
  AOI21_X1  g198(.A(new_n398), .B1(new_n399), .B2(new_n389), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n350), .A2(new_n290), .ZN(new_n401));
  OAI211_X1 g200(.A(new_n392), .B(new_n387), .C1(new_n401), .C2(new_n384), .ZN(new_n402));
  INV_X1    g201(.A(new_n402), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n400), .A2(new_n403), .ZN(new_n404));
  AOI211_X1 g203(.A(new_n378), .B(new_n382), .C1(new_n397), .C2(new_n404), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n397), .A2(new_n404), .ZN(new_n406));
  INV_X1    g205(.A(new_n382), .ZN(new_n407));
  AOI21_X1  g206(.A(KEYINPUT6), .B1(new_n406), .B2(new_n407), .ZN(new_n408));
  AOI22_X1  g207(.A1(new_n391), .A2(new_n396), .B1(new_n400), .B2(new_n403), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n409), .A2(new_n382), .ZN(new_n410));
  AOI21_X1  g209(.A(new_n405), .B1(new_n408), .B2(new_n410), .ZN(new_n411));
  NOR4_X1   g210(.A1(new_n275), .A2(new_n323), .A3(new_n377), .A4(new_n411), .ZN(new_n412));
  OAI21_X1  g211(.A(KEYINPUT81), .B1(new_n323), .B2(new_n377), .ZN(new_n413));
  NAND2_X1  g212(.A1(new_n372), .A2(new_n365), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n375), .A2(new_n376), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n414), .A2(new_n415), .ZN(new_n416));
  INV_X1    g215(.A(KEYINPUT81), .ZN(new_n417));
  NAND4_X1  g216(.A1(new_n416), .A2(new_n417), .A3(new_n321), .A4(new_n322), .ZN(new_n418));
  OAI21_X1  g217(.A(new_n378), .B1(new_n409), .B2(new_n382), .ZN(new_n419));
  NOR2_X1   g218(.A1(new_n406), .A2(new_n407), .ZN(new_n420));
  OAI21_X1  g219(.A(KEYINPUT77), .B1(new_n419), .B2(new_n420), .ZN(new_n421));
  INV_X1    g220(.A(KEYINPUT77), .ZN(new_n422));
  NAND3_X1  g221(.A1(new_n408), .A2(new_n422), .A3(new_n410), .ZN(new_n423));
  INV_X1    g222(.A(new_n405), .ZN(new_n424));
  NAND3_X1  g223(.A1(new_n421), .A2(new_n423), .A3(new_n424), .ZN(new_n425));
  AND3_X1   g224(.A1(new_n272), .A2(KEYINPUT74), .A3(new_n273), .ZN(new_n426));
  AOI21_X1  g225(.A(KEYINPUT74), .B1(new_n272), .B2(new_n273), .ZN(new_n427));
  INV_X1    g226(.A(new_n268), .ZN(new_n428));
  NOR3_X1   g227(.A1(new_n426), .A2(new_n427), .A3(new_n428), .ZN(new_n429));
  NAND4_X1  g228(.A1(new_n413), .A2(new_n418), .A3(new_n425), .A4(new_n429), .ZN(new_n430));
  AOI21_X1  g229(.A(new_n412), .B1(new_n430), .B2(KEYINPUT35), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n425), .A2(new_n429), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n432), .A2(new_n377), .ZN(new_n433));
  INV_X1    g232(.A(KEYINPUT40), .ZN(new_n434));
  AOI21_X1  g233(.A(new_n387), .B1(new_n400), .B2(new_n386), .ZN(new_n435));
  INV_X1    g234(.A(KEYINPUT39), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n435), .A2(new_n436), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n437), .A2(new_n382), .ZN(new_n438));
  OAI21_X1  g237(.A(KEYINPUT39), .B1(new_n394), .B2(new_n395), .ZN(new_n439));
  NOR2_X1   g238(.A1(new_n435), .A2(new_n439), .ZN(new_n440));
  OAI21_X1  g239(.A(new_n434), .B1(new_n438), .B2(new_n440), .ZN(new_n441));
  AOI21_X1  g240(.A(new_n407), .B1(new_n435), .B2(new_n436), .ZN(new_n442));
  OAI211_X1 g241(.A(new_n442), .B(KEYINPUT40), .C1(new_n435), .C2(new_n439), .ZN(new_n443));
  NOR2_X1   g242(.A1(new_n409), .A2(new_n382), .ZN(new_n444));
  INV_X1    g243(.A(new_n444), .ZN(new_n445));
  NAND4_X1  g244(.A1(new_n441), .A2(new_n443), .A3(new_n274), .A4(new_n445), .ZN(new_n446));
  INV_X1    g245(.A(KEYINPUT80), .ZN(new_n447));
  NAND3_X1  g246(.A1(new_n259), .A2(new_n447), .A3(new_n265), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n448), .A2(KEYINPUT37), .ZN(new_n449));
  INV_X1    g248(.A(KEYINPUT37), .ZN(new_n450));
  NAND4_X1  g249(.A1(new_n259), .A2(new_n447), .A3(new_n265), .A4(new_n450), .ZN(new_n451));
  NAND3_X1  g250(.A1(new_n449), .A2(new_n269), .A3(new_n451), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n452), .A2(KEYINPUT38), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n453), .A2(new_n411), .ZN(new_n454));
  OAI21_X1  g253(.A(new_n266), .B1(new_n452), .B2(KEYINPUT38), .ZN(new_n455));
  OAI211_X1 g254(.A(new_n416), .B(new_n446), .C1(new_n454), .C2(new_n455), .ZN(new_n456));
  INV_X1    g255(.A(KEYINPUT72), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n323), .A2(new_n457), .ZN(new_n458));
  INV_X1    g257(.A(KEYINPUT36), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  NAND3_X1  g259(.A1(new_n323), .A2(new_n457), .A3(KEYINPUT36), .ZN(new_n461));
  AND4_X1   g260(.A1(new_n433), .A2(new_n456), .A3(new_n460), .A4(new_n461), .ZN(new_n462));
  OR2_X1    g261(.A1(new_n431), .A2(new_n462), .ZN(new_n463));
  INV_X1    g262(.A(G8gat), .ZN(new_n464));
  XNOR2_X1  g263(.A(G15gat), .B(G22gat), .ZN(new_n465));
  INV_X1    g264(.A(G1gat), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n466), .A2(KEYINPUT16), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n465), .A2(new_n467), .ZN(new_n468));
  AOI21_X1  g267(.A(new_n464), .B1(new_n468), .B2(KEYINPUT88), .ZN(new_n469));
  OAI21_X1  g268(.A(new_n468), .B1(G1gat), .B2(new_n465), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  OAI221_X1 g270(.A(new_n468), .B1(KEYINPUT88), .B2(new_n464), .C1(G1gat), .C2(new_n465), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  INV_X1    g272(.A(new_n473), .ZN(new_n474));
  INV_X1    g273(.A(G29gat), .ZN(new_n475));
  INV_X1    g274(.A(G36gat), .ZN(new_n476));
  NAND3_X1  g275(.A1(new_n475), .A2(new_n476), .A3(KEYINPUT14), .ZN(new_n477));
  INV_X1    g276(.A(KEYINPUT14), .ZN(new_n478));
  OAI21_X1  g277(.A(new_n478), .B1(G29gat), .B2(G36gat), .ZN(new_n479));
  NAND2_X1  g278(.A1(G29gat), .A2(G36gat), .ZN(new_n480));
  NAND4_X1  g279(.A1(new_n477), .A2(new_n479), .A3(KEYINPUT85), .A4(new_n480), .ZN(new_n481));
  INV_X1    g280(.A(G50gat), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n482), .A2(G43gat), .ZN(new_n483));
  INV_X1    g282(.A(G43gat), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n484), .A2(G50gat), .ZN(new_n485));
  NAND3_X1  g284(.A1(new_n483), .A2(new_n485), .A3(KEYINPUT15), .ZN(new_n486));
  XNOR2_X1  g285(.A(new_n481), .B(new_n486), .ZN(new_n487));
  AND3_X1   g286(.A1(new_n477), .A2(new_n479), .A3(new_n480), .ZN(new_n488));
  INV_X1    g287(.A(KEYINPUT87), .ZN(new_n489));
  NAND3_X1  g288(.A1(new_n483), .A2(new_n485), .A3(new_n489), .ZN(new_n490));
  NAND3_X1  g289(.A1(new_n484), .A2(KEYINPUT87), .A3(G50gat), .ZN(new_n491));
  OR2_X1    g290(.A1(KEYINPUT86), .A2(KEYINPUT15), .ZN(new_n492));
  NAND2_X1  g291(.A1(KEYINPUT86), .A2(KEYINPUT15), .ZN(new_n493));
  AND3_X1   g292(.A1(new_n491), .A2(new_n492), .A3(new_n493), .ZN(new_n494));
  AND3_X1   g293(.A1(new_n488), .A2(new_n490), .A3(new_n494), .ZN(new_n495));
  INV_X1    g294(.A(KEYINPUT17), .ZN(new_n496));
  NOR3_X1   g295(.A1(new_n487), .A2(new_n495), .A3(new_n496), .ZN(new_n497));
  NAND3_X1  g296(.A1(new_n488), .A2(KEYINPUT85), .A3(new_n486), .ZN(new_n498));
  INV_X1    g297(.A(new_n486), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n499), .A2(new_n481), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n498), .A2(new_n500), .ZN(new_n501));
  NAND3_X1  g300(.A1(new_n488), .A2(new_n494), .A3(new_n490), .ZN(new_n502));
  AOI21_X1  g301(.A(KEYINPUT17), .B1(new_n501), .B2(new_n502), .ZN(new_n503));
  OAI21_X1  g302(.A(new_n474), .B1(new_n497), .B2(new_n503), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n504), .A2(KEYINPUT89), .ZN(new_n505));
  NAND2_X1  g304(.A1(G229gat), .A2(G233gat), .ZN(new_n506));
  NAND3_X1  g305(.A1(new_n473), .A2(new_n501), .A3(new_n502), .ZN(new_n507));
  INV_X1    g306(.A(KEYINPUT89), .ZN(new_n508));
  OAI211_X1 g307(.A(new_n508), .B(new_n474), .C1(new_n497), .C2(new_n503), .ZN(new_n509));
  NAND4_X1  g308(.A1(new_n505), .A2(new_n506), .A3(new_n507), .A4(new_n509), .ZN(new_n510));
  INV_X1    g309(.A(KEYINPUT18), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  AND2_X1   g311(.A1(new_n509), .A2(new_n507), .ZN(new_n513));
  NAND4_X1  g312(.A1(new_n513), .A2(KEYINPUT18), .A3(new_n506), .A4(new_n505), .ZN(new_n514));
  AND2_X1   g313(.A1(new_n499), .A2(new_n481), .ZN(new_n515));
  NOR2_X1   g314(.A1(new_n499), .A2(new_n481), .ZN(new_n516));
  OAI21_X1  g315(.A(new_n502), .B1(new_n515), .B2(new_n516), .ZN(new_n517));
  XNOR2_X1  g316(.A(new_n473), .B(new_n517), .ZN(new_n518));
  XOR2_X1   g317(.A(new_n506), .B(KEYINPUT13), .Z(new_n519));
  INV_X1    g318(.A(new_n519), .ZN(new_n520));
  OAI21_X1  g319(.A(KEYINPUT90), .B1(new_n518), .B2(new_n520), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n474), .A2(new_n517), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n522), .A2(new_n507), .ZN(new_n523));
  INV_X1    g322(.A(KEYINPUT90), .ZN(new_n524));
  NAND3_X1  g323(.A1(new_n523), .A2(new_n524), .A3(new_n519), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n521), .A2(new_n525), .ZN(new_n526));
  NAND3_X1  g325(.A1(new_n512), .A2(new_n514), .A3(new_n526), .ZN(new_n527));
  XNOR2_X1  g326(.A(G169gat), .B(G197gat), .ZN(new_n528));
  XNOR2_X1  g327(.A(KEYINPUT82), .B(KEYINPUT11), .ZN(new_n529));
  XNOR2_X1  g328(.A(new_n528), .B(new_n529), .ZN(new_n530));
  XOR2_X1   g329(.A(G113gat), .B(G141gat), .Z(new_n531));
  XNOR2_X1  g330(.A(new_n530), .B(new_n531), .ZN(new_n532));
  XNOR2_X1  g331(.A(KEYINPUT83), .B(KEYINPUT84), .ZN(new_n533));
  XNOR2_X1  g332(.A(new_n532), .B(new_n533), .ZN(new_n534));
  XNOR2_X1  g333(.A(new_n534), .B(KEYINPUT12), .ZN(new_n535));
  INV_X1    g334(.A(new_n535), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n527), .A2(new_n536), .ZN(new_n537));
  NAND4_X1  g336(.A1(new_n535), .A2(new_n514), .A3(new_n512), .A4(new_n526), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  INV_X1    g338(.A(KEYINPUT96), .ZN(new_n540));
  AND2_X1   g339(.A1(G232gat), .A2(G233gat), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n541), .A2(KEYINPUT41), .ZN(new_n542));
  NAND2_X1  g341(.A1(G99gat), .A2(G106gat), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n543), .A2(KEYINPUT8), .ZN(new_n544));
  NAND2_X1  g343(.A1(G85gat), .A2(G92gat), .ZN(new_n545));
  INV_X1    g344(.A(KEYINPUT7), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  INV_X1    g346(.A(G85gat), .ZN(new_n548));
  INV_X1    g347(.A(G92gat), .ZN(new_n549));
  NAND2_X1  g348(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  NAND3_X1  g349(.A1(KEYINPUT7), .A2(G85gat), .A3(G92gat), .ZN(new_n551));
  NAND4_X1  g350(.A1(new_n544), .A2(new_n547), .A3(new_n550), .A4(new_n551), .ZN(new_n552));
  XNOR2_X1  g351(.A(G99gat), .B(G106gat), .ZN(new_n553));
  INV_X1    g352(.A(new_n553), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n552), .A2(new_n554), .ZN(new_n555));
  AOI22_X1  g354(.A1(KEYINPUT8), .A2(new_n543), .B1(new_n548), .B2(new_n549), .ZN(new_n556));
  NAND4_X1  g355(.A1(new_n556), .A2(new_n553), .A3(new_n547), .A4(new_n551), .ZN(new_n557));
  NAND3_X1  g356(.A1(new_n555), .A2(KEYINPUT93), .A3(new_n557), .ZN(new_n558));
  AND2_X1   g357(.A1(new_n547), .A2(new_n551), .ZN(new_n559));
  INV_X1    g358(.A(KEYINPUT93), .ZN(new_n560));
  NAND4_X1  g359(.A1(new_n559), .A2(new_n560), .A3(new_n553), .A4(new_n556), .ZN(new_n561));
  AND2_X1   g360(.A1(new_n558), .A2(new_n561), .ZN(new_n562));
  OAI21_X1  g361(.A(new_n542), .B1(new_n562), .B2(new_n517), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n558), .A2(new_n561), .ZN(new_n564));
  NAND2_X1  g363(.A1(new_n564), .A2(KEYINPUT94), .ZN(new_n565));
  INV_X1    g364(.A(KEYINPUT94), .ZN(new_n566));
  NAND3_X1  g365(.A1(new_n558), .A2(new_n566), .A3(new_n561), .ZN(new_n567));
  OAI211_X1 g366(.A(new_n565), .B(new_n567), .C1(new_n497), .C2(new_n503), .ZN(new_n568));
  INV_X1    g367(.A(KEYINPUT95), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  NAND2_X1  g369(.A1(new_n517), .A2(new_n496), .ZN(new_n571));
  NAND3_X1  g370(.A1(new_n501), .A2(KEYINPUT17), .A3(new_n502), .ZN(new_n572));
  NAND2_X1  g371(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  NAND4_X1  g372(.A1(new_n573), .A2(KEYINPUT95), .A3(new_n565), .A4(new_n567), .ZN(new_n574));
  AOI21_X1  g373(.A(new_n563), .B1(new_n570), .B2(new_n574), .ZN(new_n575));
  XNOR2_X1  g374(.A(G190gat), .B(G218gat), .ZN(new_n576));
  INV_X1    g375(.A(new_n576), .ZN(new_n577));
  AOI21_X1  g376(.A(new_n540), .B1(new_n575), .B2(new_n577), .ZN(new_n578));
  NOR2_X1   g377(.A1(new_n541), .A2(KEYINPUT41), .ZN(new_n579));
  XNOR2_X1  g378(.A(G134gat), .B(G162gat), .ZN(new_n580));
  XNOR2_X1  g379(.A(new_n579), .B(new_n580), .ZN(new_n581));
  INV_X1    g380(.A(new_n581), .ZN(new_n582));
  NOR2_X1   g381(.A1(new_n575), .A2(new_n577), .ZN(new_n583));
  AOI211_X1 g382(.A(new_n576), .B(new_n563), .C1(new_n570), .C2(new_n574), .ZN(new_n584));
  OAI22_X1  g383(.A1(new_n578), .A2(new_n582), .B1(new_n583), .B2(new_n584), .ZN(new_n585));
  INV_X1    g384(.A(G57gat), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n586), .A2(KEYINPUT91), .ZN(new_n587));
  INV_X1    g386(.A(KEYINPUT91), .ZN(new_n588));
  NAND2_X1  g387(.A1(new_n588), .A2(G57gat), .ZN(new_n589));
  NAND3_X1  g388(.A1(new_n587), .A2(new_n589), .A3(G64gat), .ZN(new_n590));
  NOR2_X1   g389(.A1(new_n586), .A2(G64gat), .ZN(new_n591));
  INV_X1    g390(.A(new_n591), .ZN(new_n592));
  NAND2_X1  g391(.A1(new_n590), .A2(new_n592), .ZN(new_n593));
  NAND2_X1  g392(.A1(G71gat), .A2(G78gat), .ZN(new_n594));
  OR2_X1    g393(.A1(G71gat), .A2(G78gat), .ZN(new_n595));
  INV_X1    g394(.A(KEYINPUT9), .ZN(new_n596));
  OAI21_X1  g395(.A(new_n594), .B1(new_n595), .B2(new_n596), .ZN(new_n597));
  INV_X1    g396(.A(G64gat), .ZN(new_n598));
  NOR2_X1   g397(.A1(new_n598), .A2(G57gat), .ZN(new_n599));
  OAI21_X1  g398(.A(KEYINPUT9), .B1(new_n591), .B2(new_n599), .ZN(new_n600));
  AND2_X1   g399(.A1(new_n595), .A2(new_n594), .ZN(new_n601));
  AOI22_X1  g400(.A1(new_n593), .A2(new_n597), .B1(new_n600), .B2(new_n601), .ZN(new_n602));
  NOR2_X1   g401(.A1(new_n602), .A2(KEYINPUT21), .ZN(new_n603));
  XNOR2_X1  g402(.A(G127gat), .B(G155gat), .ZN(new_n604));
  XNOR2_X1  g403(.A(new_n603), .B(new_n604), .ZN(new_n605));
  AOI21_X1  g404(.A(new_n473), .B1(KEYINPUT21), .B2(new_n602), .ZN(new_n606));
  XOR2_X1   g405(.A(new_n605), .B(new_n606), .Z(new_n607));
  NAND2_X1  g406(.A1(G231gat), .A2(G233gat), .ZN(new_n608));
  XNOR2_X1  g407(.A(new_n608), .B(KEYINPUT92), .ZN(new_n609));
  XOR2_X1   g408(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n610));
  XNOR2_X1  g409(.A(new_n609), .B(new_n610), .ZN(new_n611));
  XNOR2_X1  g410(.A(G183gat), .B(G211gat), .ZN(new_n612));
  XNOR2_X1  g411(.A(new_n611), .B(new_n612), .ZN(new_n613));
  XNOR2_X1  g412(.A(new_n607), .B(new_n613), .ZN(new_n614));
  AND2_X1   g413(.A1(new_n570), .A2(new_n574), .ZN(new_n615));
  OAI21_X1  g414(.A(new_n576), .B1(new_n615), .B2(new_n563), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n575), .A2(new_n577), .ZN(new_n617));
  NAND4_X1  g416(.A1(new_n616), .A2(new_n540), .A3(new_n617), .A4(new_n581), .ZN(new_n618));
  NAND2_X1  g417(.A1(G230gat), .A2(G233gat), .ZN(new_n619));
  INV_X1    g418(.A(new_n602), .ZN(new_n620));
  NAND2_X1  g419(.A1(new_n564), .A2(new_n620), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n555), .A2(new_n557), .ZN(new_n622));
  NAND2_X1  g421(.A1(new_n622), .A2(new_n602), .ZN(new_n623));
  AOI21_X1  g422(.A(KEYINPUT10), .B1(new_n621), .B2(new_n623), .ZN(new_n624));
  NAND3_X1  g423(.A1(new_n564), .A2(KEYINPUT10), .A3(new_n602), .ZN(new_n625));
  INV_X1    g424(.A(new_n625), .ZN(new_n626));
  OAI21_X1  g425(.A(new_n619), .B1(new_n624), .B2(new_n626), .ZN(new_n627));
  INV_X1    g426(.A(new_n619), .ZN(new_n628));
  NAND3_X1  g427(.A1(new_n621), .A2(new_n628), .A3(new_n623), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n627), .A2(new_n629), .ZN(new_n630));
  XNOR2_X1  g429(.A(G120gat), .B(G148gat), .ZN(new_n631));
  XNOR2_X1  g430(.A(G176gat), .B(G204gat), .ZN(new_n632));
  XOR2_X1   g431(.A(new_n631), .B(new_n632), .Z(new_n633));
  INV_X1    g432(.A(new_n633), .ZN(new_n634));
  NAND2_X1  g433(.A1(new_n630), .A2(new_n634), .ZN(new_n635));
  NAND3_X1  g434(.A1(new_n627), .A2(new_n629), .A3(new_n633), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  INV_X1    g436(.A(new_n637), .ZN(new_n638));
  NAND4_X1  g437(.A1(new_n585), .A2(new_n614), .A3(new_n618), .A4(new_n638), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n639), .A2(KEYINPUT97), .ZN(new_n640));
  AND2_X1   g439(.A1(new_n585), .A2(new_n618), .ZN(new_n641));
  INV_X1    g440(.A(KEYINPUT97), .ZN(new_n642));
  NAND4_X1  g441(.A1(new_n641), .A2(new_n642), .A3(new_n614), .A4(new_n638), .ZN(new_n643));
  NAND4_X1  g442(.A1(new_n463), .A2(new_n539), .A3(new_n640), .A4(new_n643), .ZN(new_n644));
  INV_X1    g443(.A(new_n644), .ZN(new_n645));
  INV_X1    g444(.A(new_n425), .ZN(new_n646));
  NAND2_X1  g445(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  XNOR2_X1  g446(.A(new_n647), .B(G1gat), .ZN(G1324gat));
  NAND2_X1  g447(.A1(new_n645), .A2(new_n274), .ZN(new_n649));
  INV_X1    g448(.A(new_n649), .ZN(new_n650));
  NOR2_X1   g449(.A1(KEYINPUT98), .A2(KEYINPUT42), .ZN(new_n651));
  XNOR2_X1  g450(.A(KEYINPUT16), .B(G8gat), .ZN(new_n652));
  MUX2_X1   g451(.A(new_n651), .B(KEYINPUT98), .S(new_n652), .Z(new_n653));
  NAND2_X1  g452(.A1(new_n650), .A2(new_n653), .ZN(new_n654));
  NOR2_X1   g453(.A1(new_n650), .A2(new_n464), .ZN(new_n655));
  OAI21_X1  g454(.A(KEYINPUT42), .B1(new_n649), .B2(new_n652), .ZN(new_n656));
  OAI21_X1  g455(.A(new_n654), .B1(new_n655), .B2(new_n656), .ZN(new_n657));
  INV_X1    g456(.A(KEYINPUT99), .ZN(new_n658));
  XNOR2_X1  g457(.A(new_n657), .B(new_n658), .ZN(G1325gat));
  INV_X1    g458(.A(G15gat), .ZN(new_n660));
  INV_X1    g459(.A(new_n323), .ZN(new_n661));
  NAND3_X1  g460(.A1(new_n645), .A2(new_n660), .A3(new_n661), .ZN(new_n662));
  INV_X1    g461(.A(new_n460), .ZN(new_n663));
  INV_X1    g462(.A(new_n461), .ZN(new_n664));
  NOR2_X1   g463(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  INV_X1    g464(.A(new_n665), .ZN(new_n666));
  NAND2_X1  g465(.A1(new_n645), .A2(new_n666), .ZN(new_n667));
  INV_X1    g466(.A(new_n667), .ZN(new_n668));
  OAI21_X1  g467(.A(new_n662), .B1(new_n668), .B2(new_n660), .ZN(G1326gat));
  NAND2_X1  g468(.A1(new_n645), .A2(new_n377), .ZN(new_n670));
  XNOR2_X1  g469(.A(KEYINPUT43), .B(G22gat), .ZN(new_n671));
  XNOR2_X1  g470(.A(new_n670), .B(new_n671), .ZN(G1327gat));
  NAND2_X1  g471(.A1(new_n585), .A2(new_n618), .ZN(new_n673));
  OAI21_X1  g472(.A(new_n673), .B1(new_n431), .B2(new_n462), .ZN(new_n674));
  INV_X1    g473(.A(KEYINPUT44), .ZN(new_n675));
  NAND2_X1  g474(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  OAI211_X1 g475(.A(KEYINPUT44), .B(new_n673), .C1(new_n431), .C2(new_n462), .ZN(new_n677));
  AND2_X1   g476(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  INV_X1    g477(.A(new_n539), .ZN(new_n679));
  NOR3_X1   g478(.A1(new_n679), .A2(new_n614), .A3(new_n637), .ZN(new_n680));
  NAND2_X1  g479(.A1(new_n678), .A2(new_n680), .ZN(new_n681));
  OAI21_X1  g480(.A(G29gat), .B1(new_n681), .B2(new_n425), .ZN(new_n682));
  INV_X1    g481(.A(new_n674), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n683), .A2(new_n680), .ZN(new_n684));
  NAND2_X1  g483(.A1(new_n646), .A2(new_n475), .ZN(new_n685));
  OR3_X1    g484(.A1(new_n684), .A2(KEYINPUT100), .A3(new_n685), .ZN(new_n686));
  INV_X1    g485(.A(KEYINPUT45), .ZN(new_n687));
  OAI21_X1  g486(.A(KEYINPUT100), .B1(new_n684), .B2(new_n685), .ZN(new_n688));
  AND3_X1   g487(.A1(new_n686), .A2(new_n687), .A3(new_n688), .ZN(new_n689));
  AOI21_X1  g488(.A(new_n687), .B1(new_n686), .B2(new_n688), .ZN(new_n690));
  OAI21_X1  g489(.A(new_n682), .B1(new_n689), .B2(new_n690), .ZN(G1328gat));
  INV_X1    g490(.A(new_n274), .ZN(new_n692));
  NOR3_X1   g491(.A1(new_n684), .A2(G36gat), .A3(new_n692), .ZN(new_n693));
  XNOR2_X1  g492(.A(new_n693), .B(KEYINPUT46), .ZN(new_n694));
  OAI21_X1  g493(.A(G36gat), .B1(new_n681), .B2(new_n692), .ZN(new_n695));
  NAND2_X1  g494(.A1(new_n694), .A2(new_n695), .ZN(G1329gat));
  INV_X1    g495(.A(KEYINPUT101), .ZN(new_n697));
  NAND2_X1  g496(.A1(new_n697), .A2(KEYINPUT47), .ZN(new_n698));
  NOR2_X1   g497(.A1(new_n684), .A2(new_n323), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n666), .A2(G43gat), .ZN(new_n700));
  OAI221_X1 g499(.A(new_n698), .B1(new_n699), .B2(G43gat), .C1(new_n681), .C2(new_n700), .ZN(new_n701));
  NOR2_X1   g500(.A1(new_n697), .A2(KEYINPUT47), .ZN(new_n702));
  XOR2_X1   g501(.A(new_n701), .B(new_n702), .Z(G1330gat));
  OAI21_X1  g502(.A(new_n482), .B1(new_n684), .B2(new_n416), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n377), .A2(G50gat), .ZN(new_n705));
  OAI21_X1  g504(.A(new_n704), .B1(new_n681), .B2(new_n705), .ZN(new_n706));
  XNOR2_X1  g505(.A(new_n706), .B(KEYINPUT48), .ZN(G1331gat));
  INV_X1    g506(.A(new_n614), .ZN(new_n708));
  NOR4_X1   g507(.A1(new_n673), .A2(new_n539), .A3(new_n708), .A4(new_n638), .ZN(new_n709));
  AND2_X1   g508(.A1(new_n463), .A2(new_n709), .ZN(new_n710));
  NAND2_X1  g509(.A1(new_n710), .A2(new_n646), .ZN(new_n711));
  AND2_X1   g510(.A1(new_n587), .A2(new_n589), .ZN(new_n712));
  XOR2_X1   g511(.A(new_n711), .B(new_n712), .Z(G1332gat));
  INV_X1    g512(.A(KEYINPUT102), .ZN(new_n714));
  XNOR2_X1  g513(.A(new_n710), .B(new_n714), .ZN(new_n715));
  AND2_X1   g514(.A1(new_n715), .A2(new_n274), .ZN(new_n716));
  NOR2_X1   g515(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n717));
  AND2_X1   g516(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n718));
  OAI21_X1  g517(.A(new_n716), .B1(new_n717), .B2(new_n718), .ZN(new_n719));
  OAI21_X1  g518(.A(new_n719), .B1(new_n716), .B2(new_n717), .ZN(G1333gat));
  NAND2_X1  g519(.A1(new_n715), .A2(new_n666), .ZN(new_n721));
  NOR2_X1   g520(.A1(new_n323), .A2(G71gat), .ZN(new_n722));
  AOI22_X1  g521(.A1(new_n721), .A2(G71gat), .B1(new_n710), .B2(new_n722), .ZN(new_n723));
  XNOR2_X1  g522(.A(new_n723), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g523(.A1(new_n715), .A2(new_n377), .ZN(new_n725));
  XNOR2_X1  g524(.A(new_n725), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g525(.A1(new_n539), .A2(new_n614), .ZN(new_n727));
  NAND3_X1  g526(.A1(new_n463), .A2(new_n673), .A3(new_n727), .ZN(new_n728));
  INV_X1    g527(.A(KEYINPUT51), .ZN(new_n729));
  XNOR2_X1  g528(.A(new_n728), .B(new_n729), .ZN(new_n730));
  NAND2_X1  g529(.A1(new_n730), .A2(new_n637), .ZN(new_n731));
  INV_X1    g530(.A(new_n731), .ZN(new_n732));
  NAND3_X1  g531(.A1(new_n732), .A2(new_n548), .A3(new_n646), .ZN(new_n733));
  NAND2_X1  g532(.A1(new_n727), .A2(new_n637), .ZN(new_n734));
  XOR2_X1   g533(.A(new_n734), .B(KEYINPUT103), .Z(new_n735));
  NAND3_X1  g534(.A1(new_n676), .A2(new_n677), .A3(new_n735), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n736), .A2(KEYINPUT104), .ZN(new_n737));
  INV_X1    g536(.A(KEYINPUT104), .ZN(new_n738));
  NAND4_X1  g537(.A1(new_n676), .A2(new_n738), .A3(new_n677), .A4(new_n735), .ZN(new_n739));
  AND3_X1   g538(.A1(new_n737), .A2(new_n646), .A3(new_n739), .ZN(new_n740));
  OAI21_X1  g539(.A(new_n733), .B1(new_n548), .B2(new_n740), .ZN(G1336gat));
  NOR2_X1   g540(.A1(new_n692), .A2(G92gat), .ZN(new_n742));
  NOR2_X1   g541(.A1(new_n728), .A2(new_n729), .ZN(new_n743));
  AOI21_X1  g542(.A(KEYINPUT51), .B1(new_n683), .B2(new_n727), .ZN(new_n744));
  OAI211_X1 g543(.A(new_n637), .B(new_n742), .C1(new_n743), .C2(new_n744), .ZN(new_n745));
  AOI21_X1  g544(.A(KEYINPUT52), .B1(new_n745), .B2(KEYINPUT106), .ZN(new_n746));
  NAND3_X1  g545(.A1(new_n678), .A2(new_n274), .A3(new_n735), .ZN(new_n747));
  INV_X1    g546(.A(KEYINPUT107), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  NAND2_X1  g548(.A1(new_n749), .A2(G92gat), .ZN(new_n750));
  NOR2_X1   g549(.A1(new_n747), .A2(new_n748), .ZN(new_n751));
  OAI221_X1 g550(.A(new_n746), .B1(KEYINPUT106), .B2(new_n745), .C1(new_n750), .C2(new_n751), .ZN(new_n752));
  NAND3_X1  g551(.A1(new_n737), .A2(new_n274), .A3(new_n739), .ZN(new_n753));
  INV_X1    g552(.A(KEYINPUT105), .ZN(new_n754));
  AND3_X1   g553(.A1(new_n753), .A2(new_n754), .A3(G92gat), .ZN(new_n755));
  AOI21_X1  g554(.A(new_n754), .B1(new_n753), .B2(G92gat), .ZN(new_n756));
  INV_X1    g555(.A(new_n745), .ZN(new_n757));
  NOR3_X1   g556(.A1(new_n755), .A2(new_n756), .A3(new_n757), .ZN(new_n758));
  INV_X1    g557(.A(KEYINPUT52), .ZN(new_n759));
  OAI21_X1  g558(.A(new_n752), .B1(new_n758), .B2(new_n759), .ZN(G1337gat));
  INV_X1    g559(.A(G99gat), .ZN(new_n761));
  NAND3_X1  g560(.A1(new_n737), .A2(new_n666), .A3(new_n739), .ZN(new_n762));
  AOI21_X1  g561(.A(new_n761), .B1(new_n762), .B2(KEYINPUT108), .ZN(new_n763));
  OAI21_X1  g562(.A(new_n763), .B1(KEYINPUT108), .B2(new_n762), .ZN(new_n764));
  NAND3_X1  g563(.A1(new_n732), .A2(new_n761), .A3(new_n661), .ZN(new_n765));
  NAND2_X1  g564(.A1(new_n764), .A2(new_n765), .ZN(G1338gat));
  INV_X1    g565(.A(KEYINPUT53), .ZN(new_n767));
  OAI21_X1  g566(.A(G106gat), .B1(new_n736), .B2(new_n416), .ZN(new_n768));
  OR2_X1    g567(.A1(new_n416), .A2(G106gat), .ZN(new_n769));
  OAI211_X1 g568(.A(new_n767), .B(new_n768), .C1(new_n731), .C2(new_n769), .ZN(new_n770));
  NOR2_X1   g569(.A1(new_n731), .A2(new_n769), .ZN(new_n771));
  NAND3_X1  g570(.A1(new_n737), .A2(new_n377), .A3(new_n739), .ZN(new_n772));
  AOI21_X1  g571(.A(new_n771), .B1(G106gat), .B2(new_n772), .ZN(new_n773));
  OAI21_X1  g572(.A(new_n770), .B1(new_n773), .B2(new_n767), .ZN(G1339gat));
  INV_X1    g573(.A(KEYINPUT111), .ZN(new_n775));
  INV_X1    g574(.A(new_n506), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n509), .A2(new_n507), .ZN(new_n777));
  AOI21_X1  g576(.A(new_n508), .B1(new_n573), .B2(new_n474), .ZN(new_n778));
  OAI21_X1  g577(.A(new_n776), .B1(new_n777), .B2(new_n778), .ZN(new_n779));
  NAND2_X1  g578(.A1(new_n518), .A2(new_n520), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  AOI21_X1  g580(.A(new_n775), .B1(new_n781), .B2(new_n534), .ZN(new_n782));
  INV_X1    g581(.A(new_n534), .ZN(new_n783));
  AOI211_X1 g582(.A(KEYINPUT111), .B(new_n783), .C1(new_n779), .C2(new_n780), .ZN(new_n784));
  OAI211_X1 g583(.A(new_n538), .B(new_n637), .C1(new_n782), .C2(new_n784), .ZN(new_n785));
  XNOR2_X1  g584(.A(new_n785), .B(KEYINPUT112), .ZN(new_n786));
  INV_X1    g585(.A(KEYINPUT55), .ZN(new_n787));
  INV_X1    g586(.A(KEYINPUT10), .ZN(new_n788));
  AOI21_X1  g587(.A(new_n602), .B1(new_n558), .B2(new_n561), .ZN(new_n789));
  AND2_X1   g588(.A1(new_n622), .A2(new_n602), .ZN(new_n790));
  OAI21_X1  g589(.A(new_n788), .B1(new_n789), .B2(new_n790), .ZN(new_n791));
  AOI21_X1  g590(.A(new_n628), .B1(new_n791), .B2(new_n625), .ZN(new_n792));
  INV_X1    g591(.A(KEYINPUT54), .ZN(new_n793));
  AOI211_X1 g592(.A(new_n787), .B(new_n633), .C1(new_n792), .C2(new_n793), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n791), .A2(new_n625), .ZN(new_n795));
  AOI21_X1  g594(.A(new_n793), .B1(new_n795), .B2(new_n619), .ZN(new_n796));
  NAND3_X1  g595(.A1(new_n791), .A2(new_n628), .A3(new_n625), .ZN(new_n797));
  AND3_X1   g596(.A1(new_n796), .A2(KEYINPUT109), .A3(new_n797), .ZN(new_n798));
  AOI21_X1  g597(.A(KEYINPUT109), .B1(new_n796), .B2(new_n797), .ZN(new_n799));
  OAI21_X1  g598(.A(new_n794), .B1(new_n798), .B2(new_n799), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n800), .A2(new_n636), .ZN(new_n801));
  NAND3_X1  g600(.A1(new_n627), .A2(KEYINPUT54), .A3(new_n797), .ZN(new_n802));
  INV_X1    g601(.A(KEYINPUT109), .ZN(new_n803));
  NAND2_X1  g602(.A1(new_n802), .A2(new_n803), .ZN(new_n804));
  NAND3_X1  g603(.A1(new_n796), .A2(KEYINPUT109), .A3(new_n797), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  AOI21_X1  g605(.A(new_n633), .B1(new_n792), .B2(new_n793), .ZN(new_n807));
  AOI21_X1  g606(.A(KEYINPUT55), .B1(new_n806), .B2(new_n807), .ZN(new_n808));
  OAI21_X1  g607(.A(KEYINPUT110), .B1(new_n801), .B2(new_n808), .ZN(new_n809));
  OAI21_X1  g608(.A(new_n807), .B1(new_n798), .B2(new_n799), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n810), .A2(new_n787), .ZN(new_n811));
  INV_X1    g610(.A(new_n636), .ZN(new_n812));
  AOI21_X1  g611(.A(new_n812), .B1(new_n806), .B2(new_n794), .ZN(new_n813));
  INV_X1    g612(.A(KEYINPUT110), .ZN(new_n814));
  NAND3_X1  g613(.A1(new_n811), .A2(new_n813), .A3(new_n814), .ZN(new_n815));
  NAND3_X1  g614(.A1(new_n809), .A2(new_n539), .A3(new_n815), .ZN(new_n816));
  AOI21_X1  g615(.A(new_n673), .B1(new_n786), .B2(new_n816), .ZN(new_n817));
  OR2_X1    g616(.A1(new_n782), .A2(new_n784), .ZN(new_n818));
  AND2_X1   g617(.A1(new_n818), .A2(new_n538), .ZN(new_n819));
  NAND4_X1  g618(.A1(new_n819), .A2(new_n809), .A3(new_n673), .A4(new_n815), .ZN(new_n820));
  INV_X1    g619(.A(new_n820), .ZN(new_n821));
  OAI21_X1  g620(.A(new_n708), .B1(new_n817), .B2(new_n821), .ZN(new_n822));
  NOR2_X1   g621(.A1(new_n639), .A2(new_n539), .ZN(new_n823));
  INV_X1    g622(.A(new_n823), .ZN(new_n824));
  AOI21_X1  g623(.A(new_n425), .B1(new_n822), .B2(new_n824), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n413), .A2(new_n418), .ZN(new_n826));
  INV_X1    g625(.A(new_n826), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n825), .A2(new_n827), .ZN(new_n828));
  INV_X1    g627(.A(KEYINPUT114), .ZN(new_n829));
  NOR2_X1   g628(.A1(new_n828), .A2(new_n829), .ZN(new_n830));
  AOI21_X1  g629(.A(KEYINPUT114), .B1(new_n825), .B2(new_n827), .ZN(new_n831));
  NOR3_X1   g630(.A1(new_n830), .A2(new_n274), .A3(new_n831), .ZN(new_n832));
  NOR2_X1   g631(.A1(new_n679), .A2(G113gat), .ZN(new_n833));
  XNOR2_X1  g632(.A(new_n833), .B(KEYINPUT115), .ZN(new_n834));
  NAND2_X1  g633(.A1(new_n832), .A2(new_n834), .ZN(new_n835));
  NOR2_X1   g634(.A1(new_n425), .A2(new_n274), .ZN(new_n836));
  NAND2_X1  g635(.A1(new_n822), .A2(new_n824), .ZN(new_n837));
  AOI21_X1  g636(.A(KEYINPUT113), .B1(new_n837), .B2(new_n416), .ZN(new_n838));
  INV_X1    g637(.A(KEYINPUT113), .ZN(new_n839));
  AOI211_X1 g638(.A(new_n839), .B(new_n377), .C1(new_n822), .C2(new_n824), .ZN(new_n840));
  OAI211_X1 g639(.A(new_n661), .B(new_n836), .C1(new_n838), .C2(new_n840), .ZN(new_n841));
  OAI21_X1  g640(.A(G113gat), .B1(new_n841), .B2(new_n679), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n835), .A2(new_n842), .ZN(G1340gat));
  AOI21_X1  g642(.A(G120gat), .B1(new_n832), .B2(new_n637), .ZN(new_n844));
  INV_X1    g643(.A(new_n841), .ZN(new_n845));
  AND2_X1   g644(.A1(new_n637), .A2(G120gat), .ZN(new_n846));
  AOI21_X1  g645(.A(new_n844), .B1(new_n845), .B2(new_n846), .ZN(G1341gat));
  NOR2_X1   g646(.A1(new_n708), .A2(G127gat), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n832), .A2(new_n848), .ZN(new_n849));
  OAI21_X1  g648(.A(G127gat), .B1(new_n841), .B2(new_n708), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n849), .A2(new_n850), .ZN(new_n851));
  NAND2_X1  g650(.A1(new_n851), .A2(KEYINPUT116), .ZN(new_n852));
  INV_X1    g651(.A(KEYINPUT116), .ZN(new_n853));
  NAND3_X1  g652(.A1(new_n849), .A2(new_n853), .A3(new_n850), .ZN(new_n854));
  NAND2_X1  g653(.A1(new_n852), .A2(new_n854), .ZN(G1342gat));
  INV_X1    g654(.A(G134gat), .ZN(new_n856));
  NAND3_X1  g655(.A1(new_n832), .A2(new_n856), .A3(new_n673), .ZN(new_n857));
  OR2_X1    g656(.A1(new_n857), .A2(KEYINPUT56), .ZN(new_n858));
  OAI21_X1  g657(.A(G134gat), .B1(new_n841), .B2(new_n641), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n857), .A2(KEYINPUT56), .ZN(new_n860));
  NAND3_X1  g659(.A1(new_n858), .A2(new_n859), .A3(new_n860), .ZN(G1343gat));
  AND2_X1   g660(.A1(new_n665), .A2(new_n836), .ZN(new_n862));
  AOI21_X1  g661(.A(new_n416), .B1(new_n822), .B2(new_n824), .ZN(new_n863));
  NOR2_X1   g662(.A1(new_n863), .A2(KEYINPUT57), .ZN(new_n864));
  INV_X1    g663(.A(KEYINPUT57), .ZN(new_n865));
  INV_X1    g664(.A(new_n807), .ZN(new_n866));
  AOI21_X1  g665(.A(new_n866), .B1(new_n804), .B2(new_n805), .ZN(new_n867));
  OAI21_X1  g666(.A(KEYINPUT117), .B1(new_n867), .B2(KEYINPUT55), .ZN(new_n868));
  INV_X1    g667(.A(KEYINPUT117), .ZN(new_n869));
  NAND3_X1  g668(.A1(new_n810), .A2(new_n869), .A3(new_n787), .ZN(new_n870));
  NAND2_X1  g669(.A1(new_n868), .A2(new_n870), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n539), .A2(new_n813), .ZN(new_n872));
  OAI21_X1  g671(.A(new_n785), .B1(new_n871), .B2(new_n872), .ZN(new_n873));
  NAND2_X1  g672(.A1(new_n873), .A2(new_n641), .ZN(new_n874));
  INV_X1    g673(.A(new_n874), .ZN(new_n875));
  OAI21_X1  g674(.A(new_n708), .B1(new_n875), .B2(new_n821), .ZN(new_n876));
  AOI211_X1 g675(.A(new_n865), .B(new_n416), .C1(new_n876), .C2(new_n824), .ZN(new_n877));
  OAI21_X1  g676(.A(new_n862), .B1(new_n864), .B2(new_n877), .ZN(new_n878));
  OAI21_X1  g677(.A(G141gat), .B1(new_n878), .B2(new_n679), .ZN(new_n879));
  NAND4_X1  g678(.A1(new_n825), .A2(new_n377), .A3(new_n692), .A4(new_n665), .ZN(new_n880));
  INV_X1    g679(.A(new_n880), .ZN(new_n881));
  NAND3_X1  g680(.A1(new_n881), .A2(new_n331), .A3(new_n539), .ZN(new_n882));
  NAND2_X1  g681(.A1(new_n879), .A2(new_n882), .ZN(new_n883));
  XNOR2_X1  g682(.A(new_n883), .B(KEYINPUT58), .ZN(G1344gat));
  NAND3_X1  g683(.A1(new_n881), .A2(new_n332), .A3(new_n637), .ZN(new_n885));
  INV_X1    g684(.A(KEYINPUT59), .ZN(new_n886));
  NOR2_X1   g685(.A1(new_n416), .A2(new_n865), .ZN(new_n887));
  AND3_X1   g686(.A1(new_n809), .A2(new_n539), .A3(new_n815), .ZN(new_n888));
  NAND4_X1  g687(.A1(new_n818), .A2(KEYINPUT112), .A3(new_n538), .A4(new_n637), .ZN(new_n889));
  INV_X1    g688(.A(KEYINPUT112), .ZN(new_n890));
  NAND2_X1  g689(.A1(new_n785), .A2(new_n890), .ZN(new_n891));
  NAND2_X1  g690(.A1(new_n889), .A2(new_n891), .ZN(new_n892));
  OAI21_X1  g691(.A(new_n641), .B1(new_n888), .B2(new_n892), .ZN(new_n893));
  AOI21_X1  g692(.A(new_n614), .B1(new_n893), .B2(new_n820), .ZN(new_n894));
  OAI21_X1  g693(.A(new_n887), .B1(new_n894), .B2(new_n823), .ZN(new_n895));
  NAND3_X1  g694(.A1(new_n643), .A2(new_n679), .A3(new_n640), .ZN(new_n896));
  INV_X1    g695(.A(KEYINPUT120), .ZN(new_n897));
  NAND2_X1  g696(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  NAND4_X1  g697(.A1(new_n643), .A2(KEYINPUT120), .A3(new_n679), .A4(new_n640), .ZN(new_n899));
  NAND2_X1  g698(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  INV_X1    g699(.A(KEYINPUT121), .ZN(new_n901));
  OAI211_X1 g700(.A(new_n800), .B(new_n636), .C1(new_n867), .C2(KEYINPUT55), .ZN(new_n902));
  OAI21_X1  g701(.A(new_n901), .B1(new_n641), .B2(new_n902), .ZN(new_n903));
  NAND4_X1  g702(.A1(new_n673), .A2(KEYINPUT121), .A3(new_n813), .A4(new_n811), .ZN(new_n904));
  NAND3_X1  g703(.A1(new_n903), .A2(new_n819), .A3(new_n904), .ZN(new_n905));
  AOI21_X1  g704(.A(new_n614), .B1(new_n874), .B2(new_n905), .ZN(new_n906));
  OAI21_X1  g705(.A(new_n377), .B1(new_n900), .B2(new_n906), .ZN(new_n907));
  AOI22_X1  g706(.A1(new_n895), .A2(KEYINPUT119), .B1(new_n865), .B2(new_n907), .ZN(new_n908));
  INV_X1    g707(.A(KEYINPUT119), .ZN(new_n909));
  NAND3_X1  g708(.A1(new_n837), .A2(new_n909), .A3(new_n887), .ZN(new_n910));
  NAND2_X1  g709(.A1(new_n908), .A2(new_n910), .ZN(new_n911));
  INV_X1    g710(.A(new_n862), .ZN(new_n912));
  AOI21_X1  g711(.A(new_n638), .B1(new_n912), .B2(KEYINPUT118), .ZN(new_n913));
  OAI211_X1 g712(.A(new_n911), .B(new_n913), .C1(KEYINPUT118), .C2(new_n912), .ZN(new_n914));
  AOI21_X1  g713(.A(new_n886), .B1(new_n914), .B2(G148gat), .ZN(new_n915));
  NOR2_X1   g714(.A1(new_n878), .A2(new_n638), .ZN(new_n916));
  NOR3_X1   g715(.A1(new_n916), .A2(KEYINPUT59), .A3(new_n332), .ZN(new_n917));
  OAI21_X1  g716(.A(new_n885), .B1(new_n915), .B2(new_n917), .ZN(G1345gat));
  OAI21_X1  g717(.A(G155gat), .B1(new_n878), .B2(new_n708), .ZN(new_n919));
  NAND3_X1  g718(.A1(new_n881), .A2(new_n324), .A3(new_n614), .ZN(new_n920));
  NAND2_X1  g719(.A1(new_n919), .A2(new_n920), .ZN(G1346gat));
  NOR3_X1   g720(.A1(new_n878), .A2(new_n325), .A3(new_n641), .ZN(new_n922));
  AOI21_X1  g721(.A(G162gat), .B1(new_n881), .B2(new_n673), .ZN(new_n923));
  NOR2_X1   g722(.A1(new_n922), .A2(new_n923), .ZN(G1347gat));
  NOR2_X1   g723(.A1(new_n646), .A2(new_n692), .ZN(new_n925));
  NAND2_X1  g724(.A1(new_n925), .A2(new_n661), .ZN(new_n926));
  XNOR2_X1  g725(.A(new_n926), .B(KEYINPUT123), .ZN(new_n927));
  OAI21_X1  g726(.A(new_n927), .B1(new_n838), .B2(new_n840), .ZN(new_n928));
  OAI21_X1  g727(.A(G169gat), .B1(new_n928), .B2(new_n679), .ZN(new_n929));
  OR2_X1    g728(.A1(new_n929), .A2(KEYINPUT124), .ZN(new_n930));
  NAND2_X1  g729(.A1(new_n929), .A2(KEYINPUT124), .ZN(new_n931));
  NAND3_X1  g730(.A1(new_n837), .A2(new_n827), .A3(new_n925), .ZN(new_n932));
  INV_X1    g731(.A(new_n932), .ZN(new_n933));
  NAND3_X1  g732(.A1(new_n933), .A2(new_n227), .A3(new_n539), .ZN(new_n934));
  XNOR2_X1  g733(.A(new_n934), .B(KEYINPUT122), .ZN(new_n935));
  NAND3_X1  g734(.A1(new_n930), .A2(new_n931), .A3(new_n935), .ZN(G1348gat));
  OAI21_X1  g735(.A(G176gat), .B1(new_n928), .B2(new_n638), .ZN(new_n937));
  NAND3_X1  g736(.A1(new_n933), .A2(new_n228), .A3(new_n637), .ZN(new_n938));
  NAND2_X1  g737(.A1(new_n937), .A2(new_n938), .ZN(G1349gat));
  OAI21_X1  g738(.A(G183gat), .B1(new_n928), .B2(new_n708), .ZN(new_n940));
  NAND3_X1  g739(.A1(new_n933), .A2(new_n224), .A3(new_n614), .ZN(new_n941));
  NAND2_X1  g740(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  XNOR2_X1  g741(.A(new_n942), .B(KEYINPUT60), .ZN(G1350gat));
  NAND3_X1  g742(.A1(new_n933), .A2(new_n218), .A3(new_n673), .ZN(new_n944));
  OAI211_X1 g743(.A(new_n673), .B(new_n927), .C1(new_n838), .C2(new_n840), .ZN(new_n945));
  INV_X1    g744(.A(KEYINPUT61), .ZN(new_n946));
  AND3_X1   g745(.A1(new_n945), .A2(new_n946), .A3(G190gat), .ZN(new_n947));
  AOI21_X1  g746(.A(new_n946), .B1(new_n945), .B2(G190gat), .ZN(new_n948));
  OAI21_X1  g747(.A(new_n944), .B1(new_n947), .B2(new_n948), .ZN(new_n949));
  NAND2_X1  g748(.A1(new_n949), .A2(KEYINPUT125), .ZN(new_n950));
  INV_X1    g749(.A(KEYINPUT125), .ZN(new_n951));
  OAI211_X1 g750(.A(new_n944), .B(new_n951), .C1(new_n947), .C2(new_n948), .ZN(new_n952));
  NAND2_X1  g751(.A1(new_n950), .A2(new_n952), .ZN(G1351gat));
  NAND2_X1  g752(.A1(new_n665), .A2(new_n925), .ZN(new_n954));
  INV_X1    g753(.A(new_n954), .ZN(new_n955));
  AND2_X1   g754(.A1(new_n863), .A2(new_n955), .ZN(new_n956));
  AOI21_X1  g755(.A(G197gat), .B1(new_n956), .B2(new_n539), .ZN(new_n957));
  AOI21_X1  g756(.A(new_n954), .B1(new_n908), .B2(new_n910), .ZN(new_n958));
  AND2_X1   g757(.A1(new_n539), .A2(G197gat), .ZN(new_n959));
  AOI21_X1  g758(.A(new_n957), .B1(new_n958), .B2(new_n959), .ZN(G1352gat));
  NAND2_X1  g759(.A1(new_n955), .A2(new_n637), .ZN(new_n961));
  NOR2_X1   g760(.A1(new_n961), .A2(G204gat), .ZN(new_n962));
  NAND2_X1  g761(.A1(new_n962), .A2(new_n863), .ZN(new_n963));
  XOR2_X1   g762(.A(new_n963), .B(KEYINPUT62), .Z(new_n964));
  AOI21_X1  g763(.A(new_n961), .B1(new_n908), .B2(new_n910), .ZN(new_n965));
  INV_X1    g764(.A(KEYINPUT126), .ZN(new_n966));
  OAI21_X1  g765(.A(G204gat), .B1(new_n965), .B2(new_n966), .ZN(new_n967));
  AOI211_X1 g766(.A(KEYINPUT126), .B(new_n961), .C1(new_n908), .C2(new_n910), .ZN(new_n968));
  OAI21_X1  g767(.A(new_n964), .B1(new_n967), .B2(new_n968), .ZN(new_n969));
  NAND2_X1  g768(.A1(new_n969), .A2(KEYINPUT127), .ZN(new_n970));
  INV_X1    g769(.A(KEYINPUT127), .ZN(new_n971));
  OAI211_X1 g770(.A(new_n971), .B(new_n964), .C1(new_n967), .C2(new_n968), .ZN(new_n972));
  NAND2_X1  g771(.A1(new_n970), .A2(new_n972), .ZN(G1353gat));
  INV_X1    g772(.A(G211gat), .ZN(new_n974));
  NAND3_X1  g773(.A1(new_n956), .A2(new_n974), .A3(new_n614), .ZN(new_n975));
  NAND2_X1  g774(.A1(new_n958), .A2(new_n614), .ZN(new_n976));
  AND3_X1   g775(.A1(new_n976), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n977));
  AOI21_X1  g776(.A(KEYINPUT63), .B1(new_n976), .B2(G211gat), .ZN(new_n978));
  OAI21_X1  g777(.A(new_n975), .B1(new_n977), .B2(new_n978), .ZN(G1354gat));
  AOI21_X1  g778(.A(G218gat), .B1(new_n956), .B2(new_n673), .ZN(new_n980));
  AND2_X1   g779(.A1(new_n673), .A2(new_n205), .ZN(new_n981));
  AOI21_X1  g780(.A(new_n980), .B1(new_n958), .B2(new_n981), .ZN(G1355gat));
endmodule


