//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 1 1 0 1 1 0 1 0 0 1 1 1 0 1 1 0 0 0 0 1 0 0 0 1 1 0 1 1 0 0 0 0 1 0 1 0 1 1 0 0 0 0 0 1 0 1 0 1 1 1 1 1 1 1 1 0 0 1 0 0 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:24:22 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n564, new_n565, new_n566,
    new_n567, new_n568, new_n569, new_n570, new_n572, new_n573, new_n574,
    new_n575, new_n576, new_n577, new_n578, new_n579, new_n581, new_n582,
    new_n583, new_n584, new_n585, new_n586, new_n587, new_n588, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n623, new_n624, new_n625, new_n626,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n636, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n657, new_n658, new_n659,
    new_n660, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n691, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n831, new_n832, new_n833, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n846, new_n847, new_n848, new_n849, new_n850,
    new_n851, new_n852, new_n853, new_n854, new_n855, new_n856, new_n857,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n868, new_n869, new_n870, new_n871, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n912, new_n913, new_n914, new_n915, new_n916, new_n917,
    new_n918, new_n919, new_n920;
  XOR2_X1   g000(.A(KEYINPUT9), .B(G234), .Z(new_n187));
  XNOR2_X1  g001(.A(new_n187), .B(KEYINPUT77), .ZN(new_n188));
  INV_X1    g002(.A(G902), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n188), .A2(new_n189), .ZN(new_n190));
  AND2_X1   g004(.A1(new_n190), .A2(G221), .ZN(new_n191));
  INV_X1    g005(.A(G104), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n192), .A2(G107), .ZN(new_n193));
  INV_X1    g007(.A(G107), .ZN(new_n194));
  INV_X1    g008(.A(KEYINPUT3), .ZN(new_n195));
  OAI211_X1 g009(.A(G104), .B(new_n194), .C1(new_n195), .C2(KEYINPUT78), .ZN(new_n196));
  XNOR2_X1  g010(.A(KEYINPUT78), .B(KEYINPUT3), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n194), .A2(G104), .ZN(new_n198));
  INV_X1    g012(.A(new_n198), .ZN(new_n199));
  OAI211_X1 g013(.A(new_n193), .B(new_n196), .C1(new_n197), .C2(new_n199), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n200), .A2(G101), .ZN(new_n201));
  NOR2_X1   g015(.A1(new_n195), .A2(KEYINPUT78), .ZN(new_n202));
  INV_X1    g016(.A(KEYINPUT78), .ZN(new_n203));
  NOR2_X1   g017(.A1(new_n203), .A2(KEYINPUT3), .ZN(new_n204));
  OAI21_X1  g018(.A(new_n198), .B1(new_n202), .B2(new_n204), .ZN(new_n205));
  INV_X1    g019(.A(G101), .ZN(new_n206));
  NAND4_X1  g020(.A1(new_n205), .A2(new_n206), .A3(new_n193), .A4(new_n196), .ZN(new_n207));
  NAND3_X1  g021(.A1(new_n201), .A2(KEYINPUT4), .A3(new_n207), .ZN(new_n208));
  INV_X1    g022(.A(G119), .ZN(new_n209));
  OAI21_X1  g023(.A(KEYINPUT70), .B1(new_n209), .B2(G116), .ZN(new_n210));
  INV_X1    g024(.A(KEYINPUT70), .ZN(new_n211));
  INV_X1    g025(.A(G116), .ZN(new_n212));
  NAND3_X1  g026(.A1(new_n211), .A2(new_n212), .A3(G119), .ZN(new_n213));
  AOI22_X1  g027(.A1(new_n210), .A2(new_n213), .B1(G116), .B2(new_n209), .ZN(new_n214));
  XOR2_X1   g028(.A(KEYINPUT2), .B(G113), .Z(new_n215));
  XNOR2_X1  g029(.A(new_n214), .B(new_n215), .ZN(new_n216));
  INV_X1    g030(.A(KEYINPUT4), .ZN(new_n217));
  NAND3_X1  g031(.A1(new_n200), .A2(new_n217), .A3(G101), .ZN(new_n218));
  NAND3_X1  g032(.A1(new_n208), .A2(new_n216), .A3(new_n218), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n219), .A2(KEYINPUT84), .ZN(new_n220));
  NAND3_X1  g034(.A1(new_n198), .A2(new_n193), .A3(KEYINPUT79), .ZN(new_n221));
  OR3_X1    g035(.A1(new_n192), .A2(KEYINPUT79), .A3(G107), .ZN(new_n222));
  NAND3_X1  g036(.A1(new_n221), .A2(new_n222), .A3(G101), .ZN(new_n223));
  INV_X1    g037(.A(KEYINPUT80), .ZN(new_n224));
  NOR2_X1   g038(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  OAI21_X1  g039(.A(KEYINPUT80), .B1(new_n200), .B2(G101), .ZN(new_n226));
  AOI21_X1  g040(.A(new_n225), .B1(new_n226), .B2(new_n223), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n214), .A2(new_n215), .ZN(new_n228));
  NOR3_X1   g042(.A1(new_n212), .A2(KEYINPUT5), .A3(G119), .ZN(new_n229));
  AOI21_X1  g043(.A(new_n229), .B1(new_n214), .B2(KEYINPUT5), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n230), .A2(G113), .ZN(new_n231));
  NAND3_X1  g045(.A1(new_n227), .A2(new_n228), .A3(new_n231), .ZN(new_n232));
  INV_X1    g046(.A(KEYINPUT84), .ZN(new_n233));
  NAND4_X1  g047(.A1(new_n208), .A2(new_n216), .A3(new_n233), .A4(new_n218), .ZN(new_n234));
  NAND3_X1  g048(.A1(new_n220), .A2(new_n232), .A3(new_n234), .ZN(new_n235));
  XOR2_X1   g049(.A(G110), .B(G122), .Z(new_n236));
  NAND2_X1  g050(.A1(new_n235), .A2(new_n236), .ZN(new_n237));
  INV_X1    g051(.A(new_n236), .ZN(new_n238));
  NAND4_X1  g052(.A1(new_n220), .A2(new_n232), .A3(new_n238), .A4(new_n234), .ZN(new_n239));
  NAND3_X1  g053(.A1(new_n237), .A2(KEYINPUT6), .A3(new_n239), .ZN(new_n240));
  INV_X1    g054(.A(KEYINPUT0), .ZN(new_n241));
  INV_X1    g055(.A(G128), .ZN(new_n242));
  NOR2_X1   g056(.A1(new_n241), .A2(new_n242), .ZN(new_n243));
  NOR2_X1   g057(.A1(KEYINPUT0), .A2(G128), .ZN(new_n244));
  NOR2_X1   g058(.A1(new_n243), .A2(new_n244), .ZN(new_n245));
  XNOR2_X1  g059(.A(G143), .B(G146), .ZN(new_n246));
  OR2_X1    g060(.A1(new_n245), .A2(new_n246), .ZN(new_n247));
  OAI21_X1  g061(.A(new_n246), .B1(new_n241), .B2(new_n242), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n247), .A2(new_n248), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n249), .A2(G125), .ZN(new_n250));
  INV_X1    g064(.A(G146), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n251), .A2(G143), .ZN(new_n252));
  NOR2_X1   g066(.A1(new_n252), .A2(G128), .ZN(new_n253));
  NOR2_X1   g067(.A1(new_n242), .A2(KEYINPUT1), .ZN(new_n254));
  INV_X1    g068(.A(G143), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n255), .A2(G146), .ZN(new_n256));
  NOR2_X1   g070(.A1(new_n254), .A2(new_n256), .ZN(new_n257));
  NAND3_X1  g071(.A1(new_n254), .A2(new_n252), .A3(new_n256), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n258), .A2(KEYINPUT69), .ZN(new_n259));
  INV_X1    g073(.A(KEYINPUT69), .ZN(new_n260));
  NAND3_X1  g074(.A1(new_n246), .A2(new_n260), .A3(new_n254), .ZN(new_n261));
  AOI211_X1 g075(.A(new_n253), .B(new_n257), .C1(new_n259), .C2(new_n261), .ZN(new_n262));
  OAI21_X1  g076(.A(new_n250), .B1(new_n262), .B2(G125), .ZN(new_n263));
  INV_X1    g077(.A(G224), .ZN(new_n264));
  NOR2_X1   g078(.A1(new_n264), .A2(G953), .ZN(new_n265));
  INV_X1    g079(.A(new_n265), .ZN(new_n266));
  XNOR2_X1  g080(.A(new_n263), .B(new_n266), .ZN(new_n267));
  INV_X1    g081(.A(KEYINPUT6), .ZN(new_n268));
  NAND3_X1  g082(.A1(new_n235), .A2(new_n268), .A3(new_n236), .ZN(new_n269));
  NAND3_X1  g083(.A1(new_n240), .A2(new_n267), .A3(new_n269), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n231), .A2(new_n228), .ZN(new_n271));
  XOR2_X1   g085(.A(new_n227), .B(new_n271), .Z(new_n272));
  XOR2_X1   g086(.A(KEYINPUT85), .B(KEYINPUT8), .Z(new_n273));
  XNOR2_X1  g087(.A(new_n236), .B(new_n273), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n272), .A2(new_n274), .ZN(new_n275));
  AOI21_X1  g089(.A(new_n263), .B1(KEYINPUT86), .B2(new_n266), .ZN(new_n276));
  INV_X1    g090(.A(KEYINPUT7), .ZN(new_n277));
  OAI21_X1  g091(.A(new_n276), .B1(new_n277), .B2(new_n265), .ZN(new_n278));
  OAI211_X1 g092(.A(KEYINPUT7), .B(new_n266), .C1(new_n263), .C2(KEYINPUT86), .ZN(new_n279));
  NAND4_X1  g093(.A1(new_n275), .A2(new_n278), .A3(new_n239), .A4(new_n279), .ZN(new_n280));
  NAND3_X1  g094(.A1(new_n270), .A2(new_n280), .A3(new_n189), .ZN(new_n281));
  OAI21_X1  g095(.A(G210), .B1(G237), .B2(G902), .ZN(new_n282));
  INV_X1    g096(.A(new_n282), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n281), .A2(new_n283), .ZN(new_n284));
  NAND4_X1  g098(.A1(new_n270), .A2(new_n280), .A3(new_n189), .A4(new_n282), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  OAI21_X1  g100(.A(G214), .B1(G237), .B2(G902), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  INV_X1    g102(.A(KEYINPUT66), .ZN(new_n289));
  AND2_X1   g103(.A1(KEYINPUT65), .A2(G134), .ZN(new_n290));
  NOR2_X1   g104(.A1(KEYINPUT65), .A2(G134), .ZN(new_n291));
  NOR3_X1   g105(.A1(new_n290), .A2(new_n291), .A3(G137), .ZN(new_n292));
  OAI21_X1  g106(.A(new_n289), .B1(new_n292), .B2(KEYINPUT11), .ZN(new_n293));
  INV_X1    g107(.A(G137), .ZN(new_n294));
  AND3_X1   g108(.A1(new_n294), .A2(KEYINPUT11), .A3(G134), .ZN(new_n295));
  XNOR2_X1  g109(.A(KEYINPUT65), .B(G134), .ZN(new_n296));
  AOI21_X1  g110(.A(new_n295), .B1(new_n296), .B2(G137), .ZN(new_n297));
  INV_X1    g111(.A(KEYINPUT11), .ZN(new_n298));
  OAI211_X1 g112(.A(KEYINPUT66), .B(new_n298), .C1(new_n296), .C2(G137), .ZN(new_n299));
  NAND3_X1  g113(.A1(new_n293), .A2(new_n297), .A3(new_n299), .ZN(new_n300));
  INV_X1    g114(.A(KEYINPUT67), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  NAND4_X1  g116(.A1(new_n293), .A2(KEYINPUT67), .A3(new_n297), .A4(new_n299), .ZN(new_n303));
  NAND3_X1  g117(.A1(new_n302), .A2(G131), .A3(new_n303), .ZN(new_n304));
  AND3_X1   g118(.A1(new_n293), .A2(new_n297), .A3(new_n299), .ZN(new_n305));
  INV_X1    g119(.A(G131), .ZN(new_n306));
  AOI21_X1  g120(.A(KEYINPUT68), .B1(new_n305), .B2(new_n306), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n304), .A2(new_n307), .ZN(new_n308));
  NAND4_X1  g122(.A1(new_n302), .A2(KEYINPUT68), .A3(G131), .A4(new_n303), .ZN(new_n309));
  AND2_X1   g123(.A1(new_n308), .A2(new_n309), .ZN(new_n310));
  AOI21_X1  g124(.A(new_n257), .B1(new_n259), .B2(new_n261), .ZN(new_n311));
  OAI21_X1  g125(.A(new_n311), .B1(G128), .B2(new_n252), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n226), .A2(new_n223), .ZN(new_n313));
  INV_X1    g127(.A(new_n225), .ZN(new_n314));
  NAND3_X1  g128(.A1(new_n312), .A2(new_n313), .A3(new_n314), .ZN(new_n315));
  INV_X1    g129(.A(KEYINPUT10), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n315), .A2(new_n316), .ZN(new_n317));
  AND2_X1   g131(.A1(new_n208), .A2(new_n218), .ZN(new_n318));
  INV_X1    g132(.A(KEYINPUT71), .ZN(new_n319));
  AOI21_X1  g133(.A(new_n319), .B1(new_n247), .B2(new_n248), .ZN(new_n320));
  OAI211_X1 g134(.A(new_n248), .B(new_n319), .C1(new_n245), .C2(new_n246), .ZN(new_n321));
  INV_X1    g135(.A(new_n321), .ZN(new_n322));
  NOR2_X1   g136(.A1(new_n320), .A2(new_n322), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n318), .A2(new_n323), .ZN(new_n324));
  NAND3_X1  g138(.A1(new_n227), .A2(KEYINPUT10), .A3(new_n312), .ZN(new_n325));
  NAND3_X1  g139(.A1(new_n317), .A2(new_n324), .A3(new_n325), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n310), .A2(new_n326), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n308), .A2(new_n309), .ZN(new_n328));
  AOI22_X1  g142(.A1(new_n316), .A2(new_n315), .B1(new_n318), .B2(new_n323), .ZN(new_n329));
  NAND3_X1  g143(.A1(new_n328), .A2(new_n329), .A3(new_n325), .ZN(new_n330));
  INV_X1    g144(.A(KEYINPUT82), .ZN(new_n331));
  NAND3_X1  g145(.A1(new_n327), .A2(new_n330), .A3(new_n331), .ZN(new_n332));
  XNOR2_X1  g146(.A(G110), .B(G140), .ZN(new_n333));
  INV_X1    g147(.A(G953), .ZN(new_n334));
  AND2_X1   g148(.A1(new_n334), .A2(G227), .ZN(new_n335));
  XOR2_X1   g149(.A(new_n333), .B(new_n335), .Z(new_n336));
  INV_X1    g150(.A(new_n336), .ZN(new_n337));
  NAND3_X1  g151(.A1(new_n310), .A2(KEYINPUT82), .A3(new_n326), .ZN(new_n338));
  NAND3_X1  g152(.A1(new_n332), .A2(new_n337), .A3(new_n338), .ZN(new_n339));
  AND3_X1   g153(.A1(new_n221), .A2(G101), .A3(new_n222), .ZN(new_n340));
  AOI21_X1  g154(.A(new_n340), .B1(new_n207), .B2(KEYINPUT80), .ZN(new_n341));
  OAI21_X1  g155(.A(new_n262), .B1(new_n341), .B2(new_n225), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n315), .A2(new_n342), .ZN(new_n343));
  NAND3_X1  g157(.A1(new_n308), .A2(new_n343), .A3(new_n309), .ZN(new_n344));
  NOR2_X1   g158(.A1(KEYINPUT81), .A2(KEYINPUT12), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n344), .A2(new_n345), .ZN(new_n346));
  NAND2_X1  g160(.A1(KEYINPUT81), .A2(KEYINPUT12), .ZN(new_n347));
  INV_X1    g161(.A(new_n345), .ZN(new_n348));
  NAND4_X1  g162(.A1(new_n308), .A2(new_n343), .A3(new_n309), .A4(new_n348), .ZN(new_n349));
  NAND3_X1  g163(.A1(new_n346), .A2(new_n347), .A3(new_n349), .ZN(new_n350));
  NAND3_X1  g164(.A1(new_n350), .A2(new_n330), .A3(new_n336), .ZN(new_n351));
  AOI211_X1 g165(.A(G469), .B(G902), .C1(new_n339), .C2(new_n351), .ZN(new_n352));
  AOI21_X1  g166(.A(new_n337), .B1(new_n332), .B2(new_n338), .ZN(new_n353));
  AOI21_X1  g167(.A(new_n336), .B1(new_n350), .B2(new_n330), .ZN(new_n354));
  OAI21_X1  g168(.A(new_n189), .B1(new_n353), .B2(new_n354), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n355), .A2(G469), .ZN(new_n356));
  AOI21_X1  g170(.A(new_n352), .B1(new_n356), .B2(KEYINPUT83), .ZN(new_n357));
  INV_X1    g171(.A(KEYINPUT83), .ZN(new_n358));
  NAND3_X1  g172(.A1(new_n355), .A2(new_n358), .A3(G469), .ZN(new_n359));
  AOI211_X1 g173(.A(new_n191), .B(new_n288), .C1(new_n357), .C2(new_n359), .ZN(new_n360));
  NAND3_X1  g174(.A1(new_n308), .A2(new_n309), .A3(new_n323), .ZN(new_n361));
  INV_X1    g175(.A(new_n216), .ZN(new_n362));
  NOR2_X1   g176(.A1(new_n294), .A2(G134), .ZN(new_n363));
  OAI21_X1  g177(.A(G131), .B1(new_n292), .B2(new_n363), .ZN(new_n364));
  OAI211_X1 g178(.A(new_n312), .B(new_n364), .C1(G131), .C2(new_n300), .ZN(new_n365));
  NAND3_X1  g179(.A1(new_n361), .A2(new_n362), .A3(new_n365), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n366), .A2(KEYINPUT28), .ZN(new_n367));
  INV_X1    g181(.A(KEYINPUT28), .ZN(new_n368));
  NAND4_X1  g182(.A1(new_n361), .A2(new_n368), .A3(new_n362), .A4(new_n365), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n361), .A2(new_n365), .ZN(new_n370));
  AOI22_X1  g184(.A1(new_n367), .A2(new_n369), .B1(new_n216), .B2(new_n370), .ZN(new_n371));
  INV_X1    g185(.A(G237), .ZN(new_n372));
  NAND3_X1  g186(.A1(new_n372), .A2(new_n334), .A3(G210), .ZN(new_n373));
  XOR2_X1   g187(.A(new_n373), .B(KEYINPUT73), .Z(new_n374));
  XNOR2_X1  g188(.A(KEYINPUT26), .B(G101), .ZN(new_n375));
  XNOR2_X1  g189(.A(new_n374), .B(new_n375), .ZN(new_n376));
  XNOR2_X1  g190(.A(KEYINPUT72), .B(KEYINPUT27), .ZN(new_n377));
  XNOR2_X1  g191(.A(new_n376), .B(new_n377), .ZN(new_n378));
  INV_X1    g192(.A(new_n378), .ZN(new_n379));
  INV_X1    g193(.A(KEYINPUT29), .ZN(new_n380));
  NOR2_X1   g194(.A1(new_n379), .A2(new_n380), .ZN(new_n381));
  AOI21_X1  g195(.A(G902), .B1(new_n371), .B2(new_n381), .ZN(new_n382));
  NAND3_X1  g196(.A1(new_n308), .A2(new_n309), .A3(new_n249), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n383), .A2(new_n365), .ZN(new_n384));
  XOR2_X1   g198(.A(KEYINPUT64), .B(KEYINPUT30), .Z(new_n385));
  NAND2_X1  g199(.A1(new_n384), .A2(new_n385), .ZN(new_n386));
  NAND3_X1  g200(.A1(new_n361), .A2(KEYINPUT30), .A3(new_n365), .ZN(new_n387));
  NAND3_X1  g201(.A1(new_n386), .A2(new_n216), .A3(new_n387), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n388), .A2(new_n366), .ZN(new_n389));
  INV_X1    g203(.A(new_n389), .ZN(new_n390));
  NOR2_X1   g204(.A1(new_n390), .A2(new_n378), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n367), .A2(new_n369), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n384), .A2(new_n216), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n392), .A2(new_n393), .ZN(new_n394));
  OAI21_X1  g208(.A(new_n380), .B1(new_n394), .B2(new_n379), .ZN(new_n395));
  OAI21_X1  g209(.A(new_n382), .B1(new_n391), .B2(new_n395), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n396), .A2(G472), .ZN(new_n397));
  NAND3_X1  g211(.A1(new_n388), .A2(new_n366), .A3(new_n378), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n398), .A2(KEYINPUT31), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n394), .A2(new_n379), .ZN(new_n400));
  INV_X1    g214(.A(KEYINPUT31), .ZN(new_n401));
  NAND4_X1  g215(.A1(new_n388), .A2(new_n401), .A3(new_n366), .A4(new_n378), .ZN(new_n402));
  NAND3_X1  g216(.A1(new_n399), .A2(new_n400), .A3(new_n402), .ZN(new_n403));
  INV_X1    g217(.A(KEYINPUT32), .ZN(new_n404));
  NOR2_X1   g218(.A1(G472), .A2(G902), .ZN(new_n405));
  AND3_X1   g219(.A1(new_n403), .A2(new_n404), .A3(new_n405), .ZN(new_n406));
  AOI21_X1  g220(.A(new_n404), .B1(new_n403), .B2(new_n405), .ZN(new_n407));
  OAI21_X1  g221(.A(new_n397), .B1(new_n406), .B2(new_n407), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n209), .A2(G128), .ZN(new_n409));
  XNOR2_X1  g223(.A(new_n409), .B(KEYINPUT76), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n242), .A2(G119), .ZN(new_n411));
  XNOR2_X1  g225(.A(new_n411), .B(KEYINPUT75), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n410), .A2(new_n412), .ZN(new_n413));
  XNOR2_X1  g227(.A(KEYINPUT24), .B(G110), .ZN(new_n414));
  INV_X1    g228(.A(G110), .ZN(new_n415));
  NAND3_X1  g229(.A1(new_n411), .A2(new_n409), .A3(KEYINPUT23), .ZN(new_n416));
  OAI21_X1  g230(.A(new_n416), .B1(KEYINPUT23), .B2(new_n411), .ZN(new_n417));
  AOI22_X1  g231(.A1(new_n413), .A2(new_n414), .B1(new_n415), .B2(new_n417), .ZN(new_n418));
  INV_X1    g232(.A(G125), .ZN(new_n419));
  NOR3_X1   g233(.A1(new_n419), .A2(KEYINPUT16), .A3(G140), .ZN(new_n420));
  XNOR2_X1  g234(.A(G125), .B(G140), .ZN(new_n421));
  AOI21_X1  g235(.A(new_n420), .B1(new_n421), .B2(KEYINPUT16), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n422), .A2(G146), .ZN(new_n423));
  INV_X1    g237(.A(new_n421), .ZN(new_n424));
  OAI21_X1  g238(.A(new_n423), .B1(G146), .B2(new_n424), .ZN(new_n425));
  OR2_X1    g239(.A1(new_n418), .A2(new_n425), .ZN(new_n426));
  OAI22_X1  g240(.A1(new_n413), .A2(new_n414), .B1(new_n415), .B2(new_n417), .ZN(new_n427));
  XNOR2_X1  g241(.A(new_n422), .B(new_n251), .ZN(new_n428));
  OR2_X1    g242(.A1(new_n427), .A2(new_n428), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n426), .A2(new_n429), .ZN(new_n430));
  NAND3_X1  g244(.A1(new_n334), .A2(G221), .A3(G234), .ZN(new_n431));
  XNOR2_X1  g245(.A(new_n431), .B(KEYINPUT22), .ZN(new_n432));
  XNOR2_X1  g246(.A(new_n432), .B(G137), .ZN(new_n433));
  INV_X1    g247(.A(new_n433), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n430), .A2(new_n434), .ZN(new_n435));
  NAND3_X1  g249(.A1(new_n426), .A2(new_n429), .A3(new_n433), .ZN(new_n436));
  AND2_X1   g250(.A1(new_n435), .A2(new_n436), .ZN(new_n437));
  INV_X1    g251(.A(new_n437), .ZN(new_n438));
  OR3_X1    g252(.A1(new_n438), .A2(KEYINPUT25), .A3(G902), .ZN(new_n439));
  OAI21_X1  g253(.A(KEYINPUT25), .B1(new_n438), .B2(G902), .ZN(new_n440));
  INV_X1    g254(.A(G234), .ZN(new_n441));
  OAI21_X1  g255(.A(G217), .B1(new_n441), .B2(G902), .ZN(new_n442));
  XNOR2_X1  g256(.A(new_n442), .B(KEYINPUT74), .ZN(new_n443));
  NAND3_X1  g257(.A1(new_n439), .A2(new_n440), .A3(new_n443), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n442), .A2(new_n189), .ZN(new_n445));
  INV_X1    g259(.A(new_n445), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n437), .A2(new_n446), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n444), .A2(new_n447), .ZN(new_n448));
  INV_X1    g262(.A(new_n448), .ZN(new_n449));
  XNOR2_X1  g263(.A(new_n421), .B(G146), .ZN(new_n450));
  OR2_X1    g264(.A1(new_n450), .A2(KEYINPUT87), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n450), .A2(KEYINPUT87), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n451), .A2(new_n452), .ZN(new_n453));
  NAND3_X1  g267(.A1(new_n372), .A2(new_n334), .A3(G214), .ZN(new_n454));
  XNOR2_X1  g268(.A(new_n454), .B(new_n255), .ZN(new_n455));
  AND2_X1   g269(.A1(KEYINPUT18), .A2(G131), .ZN(new_n456));
  XNOR2_X1  g270(.A(new_n455), .B(new_n456), .ZN(new_n457));
  INV_X1    g271(.A(new_n457), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n453), .A2(new_n458), .ZN(new_n459));
  NAND3_X1  g273(.A1(new_n455), .A2(KEYINPUT17), .A3(G131), .ZN(new_n460));
  XNOR2_X1  g274(.A(new_n455), .B(G131), .ZN(new_n461));
  OAI211_X1 g275(.A(new_n428), .B(new_n460), .C1(new_n461), .C2(KEYINPUT17), .ZN(new_n462));
  XNOR2_X1  g276(.A(G113), .B(G122), .ZN(new_n463));
  XNOR2_X1  g277(.A(new_n463), .B(new_n192), .ZN(new_n464));
  XNOR2_X1  g278(.A(new_n464), .B(KEYINPUT89), .ZN(new_n465));
  NAND3_X1  g279(.A1(new_n459), .A2(new_n462), .A3(new_n465), .ZN(new_n466));
  INV_X1    g280(.A(new_n466), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n459), .A2(new_n462), .ZN(new_n468));
  INV_X1    g282(.A(KEYINPUT90), .ZN(new_n469));
  AOI21_X1  g283(.A(new_n464), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  NAND3_X1  g284(.A1(new_n459), .A2(new_n462), .A3(KEYINPUT90), .ZN(new_n471));
  AOI21_X1  g285(.A(new_n467), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  OAI21_X1  g286(.A(G475), .B1(new_n472), .B2(G902), .ZN(new_n473));
  INV_X1    g287(.A(new_n464), .ZN(new_n474));
  NAND2_X1  g288(.A1(KEYINPUT88), .A2(KEYINPUT19), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n421), .A2(new_n475), .ZN(new_n476));
  NOR2_X1   g290(.A1(KEYINPUT88), .A2(KEYINPUT19), .ZN(new_n477));
  XNOR2_X1  g291(.A(new_n476), .B(new_n477), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n478), .A2(new_n251), .ZN(new_n479));
  AND3_X1   g293(.A1(new_n479), .A2(new_n461), .A3(new_n423), .ZN(new_n480));
  AOI21_X1  g294(.A(new_n457), .B1(new_n451), .B2(new_n452), .ZN(new_n481));
  OAI21_X1  g295(.A(new_n474), .B1(new_n480), .B2(new_n481), .ZN(new_n482));
  AOI21_X1  g296(.A(G475), .B1(new_n482), .B2(new_n466), .ZN(new_n483));
  AOI21_X1  g297(.A(KEYINPUT20), .B1(new_n483), .B2(new_n189), .ZN(new_n484));
  INV_X1    g298(.A(new_n484), .ZN(new_n485));
  NAND3_X1  g299(.A1(new_n483), .A2(KEYINPUT20), .A3(new_n189), .ZN(new_n486));
  NAND3_X1  g300(.A1(new_n473), .A2(new_n485), .A3(new_n486), .ZN(new_n487));
  AND2_X1   g301(.A1(new_n334), .A2(G952), .ZN(new_n488));
  NAND2_X1  g302(.A1(G234), .A2(G237), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  INV_X1    g304(.A(new_n490), .ZN(new_n491));
  XOR2_X1   g305(.A(KEYINPUT21), .B(G898), .Z(new_n492));
  INV_X1    g306(.A(new_n492), .ZN(new_n493));
  NAND3_X1  g307(.A1(new_n489), .A2(G902), .A3(G953), .ZN(new_n494));
  INV_X1    g308(.A(new_n494), .ZN(new_n495));
  AOI21_X1  g309(.A(new_n491), .B1(new_n493), .B2(new_n495), .ZN(new_n496));
  AOI21_X1  g310(.A(KEYINPUT13), .B1(new_n255), .B2(G128), .ZN(new_n497));
  OR2_X1    g311(.A1(new_n497), .A2(KEYINPUT92), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n242), .A2(G143), .ZN(new_n499));
  NAND3_X1  g313(.A1(new_n255), .A2(KEYINPUT13), .A3(G128), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n497), .A2(KEYINPUT92), .ZN(new_n501));
  NAND4_X1  g315(.A1(new_n498), .A2(new_n499), .A3(new_n500), .A4(new_n501), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n502), .A2(G134), .ZN(new_n503));
  XNOR2_X1  g317(.A(G128), .B(G143), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n296), .A2(new_n504), .ZN(new_n505));
  AND2_X1   g319(.A1(KEYINPUT91), .A2(G122), .ZN(new_n506));
  NOR2_X1   g320(.A1(KEYINPUT91), .A2(G122), .ZN(new_n507));
  OAI21_X1  g321(.A(G116), .B1(new_n506), .B2(new_n507), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n212), .A2(G122), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  NOR2_X1   g324(.A1(new_n510), .A2(G107), .ZN(new_n511));
  AOI21_X1  g325(.A(new_n194), .B1(new_n508), .B2(new_n509), .ZN(new_n512));
  OAI211_X1 g326(.A(new_n503), .B(new_n505), .C1(new_n511), .C2(new_n512), .ZN(new_n513));
  AOI21_X1  g327(.A(new_n194), .B1(new_n508), .B2(KEYINPUT14), .ZN(new_n514));
  OR2_X1    g328(.A1(new_n514), .A2(new_n510), .ZN(new_n515));
  XNOR2_X1  g329(.A(new_n296), .B(new_n504), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n514), .A2(new_n510), .ZN(new_n517));
  NAND3_X1  g331(.A1(new_n515), .A2(new_n516), .A3(new_n517), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n513), .A2(new_n518), .ZN(new_n519));
  NAND3_X1  g333(.A1(new_n188), .A2(G217), .A3(new_n334), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  INV_X1    g335(.A(new_n520), .ZN(new_n522));
  NAND3_X1  g336(.A1(new_n513), .A2(new_n518), .A3(new_n522), .ZN(new_n523));
  NAND3_X1  g337(.A1(new_n521), .A2(KEYINPUT93), .A3(new_n523), .ZN(new_n524));
  INV_X1    g338(.A(KEYINPUT93), .ZN(new_n525));
  NAND3_X1  g339(.A1(new_n519), .A2(new_n525), .A3(new_n520), .ZN(new_n526));
  NAND3_X1  g340(.A1(new_n524), .A2(new_n189), .A3(new_n526), .ZN(new_n527));
  INV_X1    g341(.A(G478), .ZN(new_n528));
  NOR2_X1   g342(.A1(new_n528), .A2(KEYINPUT15), .ZN(new_n529));
  XNOR2_X1  g343(.A(new_n527), .B(new_n529), .ZN(new_n530));
  NOR3_X1   g344(.A1(new_n487), .A2(new_n496), .A3(new_n530), .ZN(new_n531));
  NAND4_X1  g345(.A1(new_n360), .A2(new_n408), .A3(new_n449), .A4(new_n531), .ZN(new_n532));
  XOR2_X1   g346(.A(KEYINPUT94), .B(G101), .Z(new_n533));
  XNOR2_X1  g347(.A(new_n532), .B(new_n533), .ZN(G3));
  AOI211_X1 g348(.A(new_n448), .B(new_n191), .C1(new_n357), .C2(new_n359), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n403), .A2(new_n405), .ZN(new_n536));
  INV_X1    g350(.A(new_n536), .ZN(new_n537));
  INV_X1    g351(.A(G472), .ZN(new_n538));
  AOI21_X1  g352(.A(new_n538), .B1(new_n403), .B2(new_n189), .ZN(new_n539));
  NOR2_X1   g353(.A1(new_n537), .A2(new_n539), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n535), .A2(new_n540), .ZN(new_n541));
  XNOR2_X1  g355(.A(new_n541), .B(KEYINPUT95), .ZN(new_n542));
  INV_X1    g356(.A(KEYINPUT33), .ZN(new_n543));
  NAND3_X1  g357(.A1(new_n524), .A2(new_n543), .A3(new_n526), .ZN(new_n544));
  NAND3_X1  g358(.A1(new_n521), .A2(KEYINPUT33), .A3(new_n523), .ZN(new_n545));
  NAND3_X1  g359(.A1(new_n544), .A2(new_n189), .A3(new_n545), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n546), .A2(G478), .ZN(new_n547));
  OR2_X1    g361(.A1(new_n527), .A2(G478), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n549), .A2(KEYINPUT97), .ZN(new_n550));
  INV_X1    g364(.A(KEYINPUT97), .ZN(new_n551));
  NAND3_X1  g365(.A1(new_n547), .A2(new_n551), .A3(new_n548), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n550), .A2(new_n552), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n553), .A2(new_n487), .ZN(new_n554));
  INV_X1    g368(.A(KEYINPUT96), .ZN(new_n555));
  NAND3_X1  g369(.A1(new_n284), .A2(new_n555), .A3(new_n285), .ZN(new_n556));
  INV_X1    g370(.A(new_n496), .ZN(new_n557));
  NAND3_X1  g371(.A1(new_n281), .A2(KEYINPUT96), .A3(new_n283), .ZN(new_n558));
  NAND4_X1  g372(.A1(new_n556), .A2(new_n557), .A3(new_n287), .A4(new_n558), .ZN(new_n559));
  NOR2_X1   g373(.A1(new_n554), .A2(new_n559), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n542), .A2(new_n560), .ZN(new_n561));
  XOR2_X1   g375(.A(KEYINPUT34), .B(G104), .Z(new_n562));
  XNOR2_X1  g376(.A(new_n561), .B(new_n562), .ZN(G6));
  INV_X1    g377(.A(new_n487), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n564), .A2(new_n530), .ZN(new_n565));
  NOR2_X1   g379(.A1(new_n559), .A2(new_n565), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n542), .A2(new_n566), .ZN(new_n567));
  XNOR2_X1  g381(.A(KEYINPUT35), .B(G107), .ZN(new_n568));
  XNOR2_X1  g382(.A(new_n567), .B(new_n568), .ZN(new_n569));
  XNOR2_X1  g383(.A(KEYINPUT98), .B(KEYINPUT99), .ZN(new_n570));
  XNOR2_X1  g384(.A(new_n569), .B(new_n570), .ZN(G9));
  XOR2_X1   g385(.A(new_n430), .B(KEYINPUT100), .Z(new_n572));
  NOR2_X1   g386(.A1(new_n434), .A2(KEYINPUT36), .ZN(new_n573));
  OR2_X1    g387(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n572), .A2(new_n573), .ZN(new_n575));
  NAND3_X1  g389(.A1(new_n574), .A2(new_n446), .A3(new_n575), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n444), .A2(new_n576), .ZN(new_n577));
  NAND4_X1  g391(.A1(new_n360), .A2(new_n531), .A3(new_n540), .A4(new_n577), .ZN(new_n578));
  XNOR2_X1  g392(.A(new_n578), .B(KEYINPUT37), .ZN(new_n579));
  XNOR2_X1  g393(.A(new_n579), .B(new_n415), .ZN(G12));
  AOI21_X1  g394(.A(new_n191), .B1(new_n357), .B2(new_n359), .ZN(new_n581));
  XNOR2_X1  g395(.A(KEYINPUT101), .B(G900), .ZN(new_n582));
  AOI21_X1  g396(.A(new_n491), .B1(new_n495), .B2(new_n582), .ZN(new_n583));
  NOR2_X1   g397(.A1(new_n565), .A2(new_n583), .ZN(new_n584));
  NAND3_X1  g398(.A1(new_n556), .A2(new_n287), .A3(new_n558), .ZN(new_n585));
  INV_X1    g399(.A(new_n577), .ZN(new_n586));
  NOR2_X1   g400(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  NAND4_X1  g401(.A1(new_n408), .A2(new_n581), .A3(new_n584), .A4(new_n587), .ZN(new_n588));
  XNOR2_X1  g402(.A(new_n588), .B(G128), .ZN(G30));
  NAND2_X1  g403(.A1(new_n356), .A2(KEYINPUT83), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n339), .A2(new_n351), .ZN(new_n591));
  INV_X1    g405(.A(G469), .ZN(new_n592));
  NAND3_X1  g406(.A1(new_n591), .A2(new_n592), .A3(new_n189), .ZN(new_n593));
  NAND3_X1  g407(.A1(new_n590), .A2(new_n359), .A3(new_n593), .ZN(new_n594));
  INV_X1    g408(.A(new_n191), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  XNOR2_X1  g410(.A(new_n583), .B(KEYINPUT39), .ZN(new_n597));
  NOR2_X1   g411(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n598), .A2(KEYINPUT40), .ZN(new_n599));
  INV_X1    g413(.A(KEYINPUT40), .ZN(new_n600));
  OAI21_X1  g414(.A(new_n600), .B1(new_n596), .B2(new_n597), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n599), .A2(new_n601), .ZN(new_n602));
  INV_X1    g416(.A(KEYINPUT102), .ZN(new_n603));
  XNOR2_X1  g417(.A(new_n286), .B(new_n603), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n604), .A2(KEYINPUT38), .ZN(new_n605));
  XNOR2_X1  g419(.A(new_n286), .B(KEYINPUT102), .ZN(new_n606));
  INV_X1    g420(.A(KEYINPUT38), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n605), .A2(new_n608), .ZN(new_n609));
  NAND3_X1  g423(.A1(new_n487), .A2(new_n530), .A3(new_n287), .ZN(new_n610));
  OAI21_X1  g424(.A(KEYINPUT104), .B1(new_n577), .B2(new_n610), .ZN(new_n611));
  OR3_X1    g425(.A1(new_n577), .A2(KEYINPUT104), .A3(new_n610), .ZN(new_n612));
  AOI21_X1  g426(.A(new_n609), .B1(new_n611), .B2(new_n612), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n370), .A2(new_n216), .ZN(new_n614));
  AOI21_X1  g428(.A(new_n378), .B1(new_n614), .B2(new_n366), .ZN(new_n615));
  OR2_X1    g429(.A1(new_n615), .A2(KEYINPUT103), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n615), .A2(KEYINPUT103), .ZN(new_n617));
  AND3_X1   g431(.A1(new_n616), .A2(new_n398), .A3(new_n617), .ZN(new_n618));
  OAI21_X1  g432(.A(G472), .B1(new_n618), .B2(G902), .ZN(new_n619));
  OAI21_X1  g433(.A(new_n619), .B1(new_n406), .B2(new_n407), .ZN(new_n620));
  NAND3_X1  g434(.A1(new_n602), .A2(new_n613), .A3(new_n620), .ZN(new_n621));
  XNOR2_X1  g435(.A(new_n621), .B(G143), .ZN(G45));
  INV_X1    g436(.A(new_n583), .ZN(new_n623));
  NAND3_X1  g437(.A1(new_n553), .A2(new_n487), .A3(new_n623), .ZN(new_n624));
  INV_X1    g438(.A(new_n624), .ZN(new_n625));
  NAND4_X1  g439(.A1(new_n408), .A2(new_n581), .A3(new_n587), .A4(new_n625), .ZN(new_n626));
  XNOR2_X1  g440(.A(new_n626), .B(G146), .ZN(G48));
  NOR2_X1   g441(.A1(new_n592), .A2(KEYINPUT105), .ZN(new_n628));
  INV_X1    g442(.A(new_n628), .ZN(new_n629));
  AOI21_X1  g443(.A(new_n629), .B1(new_n591), .B2(new_n189), .ZN(new_n630));
  AOI211_X1 g444(.A(G902), .B(new_n628), .C1(new_n339), .C2(new_n351), .ZN(new_n631));
  NOR3_X1   g445(.A1(new_n630), .A2(new_n631), .A3(new_n191), .ZN(new_n632));
  NAND4_X1  g446(.A1(new_n408), .A2(new_n449), .A3(new_n560), .A4(new_n632), .ZN(new_n633));
  XNOR2_X1  g447(.A(KEYINPUT41), .B(G113), .ZN(new_n634));
  XNOR2_X1  g448(.A(new_n633), .B(new_n634), .ZN(G15));
  NAND4_X1  g449(.A1(new_n408), .A2(new_n449), .A3(new_n566), .A4(new_n632), .ZN(new_n636));
  XNOR2_X1  g450(.A(new_n636), .B(G116), .ZN(G18));
  INV_X1    g451(.A(new_n630), .ZN(new_n638));
  NAND3_X1  g452(.A1(new_n591), .A2(new_n189), .A3(new_n629), .ZN(new_n639));
  NAND3_X1  g453(.A1(new_n638), .A2(new_n595), .A3(new_n639), .ZN(new_n640));
  OAI21_X1  g454(.A(KEYINPUT106), .B1(new_n640), .B2(new_n585), .ZN(new_n641));
  AND3_X1   g455(.A1(new_n556), .A2(new_n287), .A3(new_n558), .ZN(new_n642));
  INV_X1    g456(.A(KEYINPUT106), .ZN(new_n643));
  NAND3_X1  g457(.A1(new_n642), .A2(new_n632), .A3(new_n643), .ZN(new_n644));
  NAND2_X1  g458(.A1(new_n641), .A2(new_n644), .ZN(new_n645));
  NAND4_X1  g459(.A1(new_n645), .A2(new_n408), .A3(new_n531), .A4(new_n577), .ZN(new_n646));
  XNOR2_X1  g460(.A(new_n646), .B(G119), .ZN(G21));
  OR2_X1    g461(.A1(new_n371), .A2(new_n378), .ZN(new_n648));
  NAND3_X1  g462(.A1(new_n648), .A2(new_n399), .A3(new_n402), .ZN(new_n649));
  AND2_X1   g463(.A1(new_n649), .A2(new_n405), .ZN(new_n650));
  NOR3_X1   g464(.A1(new_n650), .A2(new_n539), .A3(new_n448), .ZN(new_n651));
  NAND2_X1  g465(.A1(new_n487), .A2(new_n530), .ZN(new_n652));
  NOR2_X1   g466(.A1(new_n640), .A2(new_n652), .ZN(new_n653));
  NAND4_X1  g467(.A1(new_n651), .A2(new_n557), .A3(new_n642), .A4(new_n653), .ZN(new_n654));
  XNOR2_X1  g468(.A(new_n654), .B(KEYINPUT107), .ZN(new_n655));
  XOR2_X1   g469(.A(new_n655), .B(G122), .Z(G24));
  NOR3_X1   g470(.A1(new_n650), .A2(new_n539), .A3(new_n586), .ZN(new_n657));
  NOR3_X1   g471(.A1(new_n640), .A2(new_n585), .A3(KEYINPUT106), .ZN(new_n658));
  AOI21_X1  g472(.A(new_n643), .B1(new_n642), .B2(new_n632), .ZN(new_n659));
  OAI211_X1 g473(.A(new_n657), .B(new_n625), .C1(new_n658), .C2(new_n659), .ZN(new_n660));
  XNOR2_X1  g474(.A(new_n660), .B(G125), .ZN(G27));
  INV_X1    g475(.A(KEYINPUT109), .ZN(new_n662));
  NOR2_X1   g476(.A1(new_n662), .A2(KEYINPUT42), .ZN(new_n663));
  INV_X1    g477(.A(new_n663), .ZN(new_n664));
  NAND2_X1  g478(.A1(new_n332), .A2(new_n338), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n665), .A2(new_n336), .ZN(new_n666));
  NAND2_X1  g480(.A1(new_n666), .A2(KEYINPUT108), .ZN(new_n667));
  INV_X1    g481(.A(new_n354), .ZN(new_n668));
  INV_X1    g482(.A(KEYINPUT108), .ZN(new_n669));
  NAND2_X1  g483(.A1(new_n353), .A2(new_n669), .ZN(new_n670));
  NAND4_X1  g484(.A1(new_n667), .A2(G469), .A3(new_n668), .A4(new_n670), .ZN(new_n671));
  NOR2_X1   g485(.A1(new_n592), .A2(new_n189), .ZN(new_n672));
  INV_X1    g486(.A(new_n672), .ZN(new_n673));
  NAND3_X1  g487(.A1(new_n671), .A2(new_n593), .A3(new_n673), .ZN(new_n674));
  AND2_X1   g488(.A1(new_n674), .A2(new_n595), .ZN(new_n675));
  INV_X1    g489(.A(new_n287), .ZN(new_n676));
  NOR2_X1   g490(.A1(new_n286), .A2(new_n676), .ZN(new_n677));
  NAND4_X1  g491(.A1(new_n408), .A2(new_n675), .A3(new_n449), .A4(new_n677), .ZN(new_n678));
  NOR2_X1   g492(.A1(new_n678), .A2(new_n624), .ZN(new_n679));
  NAND2_X1  g493(.A1(new_n662), .A2(KEYINPUT42), .ZN(new_n680));
  INV_X1    g494(.A(new_n680), .ZN(new_n681));
  OAI21_X1  g495(.A(new_n664), .B1(new_n679), .B2(new_n681), .ZN(new_n682));
  INV_X1    g496(.A(new_n407), .ZN(new_n683));
  NAND3_X1  g497(.A1(new_n403), .A2(new_n404), .A3(new_n405), .ZN(new_n684));
  NAND2_X1  g498(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  AOI21_X1  g499(.A(new_n448), .B1(new_n685), .B2(new_n397), .ZN(new_n686));
  NAND4_X1  g500(.A1(new_n686), .A2(new_n625), .A3(new_n677), .A4(new_n675), .ZN(new_n687));
  NAND2_X1  g501(.A1(new_n687), .A2(new_n663), .ZN(new_n688));
  NAND2_X1  g502(.A1(new_n682), .A2(new_n688), .ZN(new_n689));
  XNOR2_X1  g503(.A(new_n689), .B(G131), .ZN(G33));
  NAND4_X1  g504(.A1(new_n686), .A2(new_n584), .A3(new_n677), .A4(new_n675), .ZN(new_n691));
  XNOR2_X1  g505(.A(new_n691), .B(G134), .ZN(G36));
  INV_X1    g506(.A(new_n540), .ZN(new_n693));
  INV_X1    g507(.A(KEYINPUT110), .ZN(new_n694));
  NAND2_X1  g508(.A1(new_n487), .A2(new_n694), .ZN(new_n695));
  NAND4_X1  g509(.A1(new_n473), .A2(KEYINPUT110), .A3(new_n485), .A4(new_n486), .ZN(new_n696));
  INV_X1    g510(.A(new_n552), .ZN(new_n697));
  AOI21_X1  g511(.A(new_n551), .B1(new_n547), .B2(new_n548), .ZN(new_n698));
  OAI211_X1 g512(.A(new_n695), .B(new_n696), .C1(new_n697), .C2(new_n698), .ZN(new_n699));
  NAND2_X1  g513(.A1(new_n699), .A2(KEYINPUT43), .ZN(new_n700));
  INV_X1    g514(.A(KEYINPUT43), .ZN(new_n701));
  NAND3_X1  g515(.A1(new_n553), .A2(new_n701), .A3(new_n564), .ZN(new_n702));
  AND3_X1   g516(.A1(new_n700), .A2(KEYINPUT111), .A3(new_n702), .ZN(new_n703));
  AOI21_X1  g517(.A(KEYINPUT111), .B1(new_n700), .B2(new_n702), .ZN(new_n704));
  OAI211_X1 g518(.A(new_n693), .B(new_n577), .C1(new_n703), .C2(new_n704), .ZN(new_n705));
  INV_X1    g519(.A(KEYINPUT44), .ZN(new_n706));
  NAND2_X1  g520(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  INV_X1    g521(.A(KEYINPUT111), .ZN(new_n708));
  AOI22_X1  g522(.A1(new_n550), .A2(new_n552), .B1(new_n694), .B2(new_n487), .ZN(new_n709));
  AOI21_X1  g523(.A(new_n701), .B1(new_n709), .B2(new_n696), .ZN(new_n710));
  INV_X1    g524(.A(new_n702), .ZN(new_n711));
  OAI21_X1  g525(.A(new_n708), .B1(new_n710), .B2(new_n711), .ZN(new_n712));
  NAND3_X1  g526(.A1(new_n700), .A2(KEYINPUT111), .A3(new_n702), .ZN(new_n713));
  NAND2_X1  g527(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  NAND4_X1  g528(.A1(new_n714), .A2(KEYINPUT44), .A3(new_n693), .A4(new_n577), .ZN(new_n715));
  INV_X1    g529(.A(new_n597), .ZN(new_n716));
  NAND2_X1  g530(.A1(new_n668), .A2(new_n666), .ZN(new_n717));
  INV_X1    g531(.A(KEYINPUT45), .ZN(new_n718));
  AOI21_X1  g532(.A(new_n592), .B1(new_n717), .B2(new_n718), .ZN(new_n719));
  NAND4_X1  g533(.A1(new_n667), .A2(KEYINPUT45), .A3(new_n668), .A4(new_n670), .ZN(new_n720));
  AOI21_X1  g534(.A(new_n672), .B1(new_n719), .B2(new_n720), .ZN(new_n721));
  NAND2_X1  g535(.A1(new_n721), .A2(KEYINPUT46), .ZN(new_n722));
  INV_X1    g536(.A(new_n722), .ZN(new_n723));
  OAI21_X1  g537(.A(new_n593), .B1(new_n721), .B2(KEYINPUT46), .ZN(new_n724));
  OAI211_X1 g538(.A(new_n595), .B(new_n716), .C1(new_n723), .C2(new_n724), .ZN(new_n725));
  INV_X1    g539(.A(new_n725), .ZN(new_n726));
  NAND4_X1  g540(.A1(new_n707), .A2(new_n715), .A3(new_n677), .A4(new_n726), .ZN(new_n727));
  XNOR2_X1  g541(.A(new_n727), .B(G137), .ZN(G39));
  OAI21_X1  g542(.A(new_n595), .B1(new_n723), .B2(new_n724), .ZN(new_n729));
  XNOR2_X1  g543(.A(KEYINPUT112), .B(KEYINPUT47), .ZN(new_n730));
  INV_X1    g544(.A(new_n730), .ZN(new_n731));
  NAND2_X1  g545(.A1(new_n729), .A2(new_n731), .ZN(new_n732));
  OAI211_X1 g546(.A(new_n595), .B(new_n730), .C1(new_n723), .C2(new_n724), .ZN(new_n733));
  NOR4_X1   g547(.A1(new_n408), .A2(new_n449), .A3(new_n676), .A4(new_n286), .ZN(new_n734));
  NAND4_X1  g548(.A1(new_n732), .A2(new_n625), .A3(new_n733), .A4(new_n734), .ZN(new_n735));
  XNOR2_X1  g549(.A(new_n735), .B(G140), .ZN(G42));
  NOR2_X1   g550(.A1(new_n630), .A2(new_n631), .ZN(new_n737));
  XNOR2_X1  g551(.A(new_n737), .B(KEYINPUT49), .ZN(new_n738));
  NAND4_X1  g552(.A1(new_n609), .A2(new_n449), .A3(new_n287), .A4(new_n738), .ZN(new_n739));
  OR4_X1    g553(.A1(new_n191), .A2(new_n739), .A3(new_n620), .A4(new_n699), .ZN(new_n740));
  INV_X1    g554(.A(KEYINPUT53), .ZN(new_n741));
  NAND4_X1  g555(.A1(new_n646), .A2(new_n633), .A3(new_n636), .A4(new_n654), .ZN(new_n742));
  NAND2_X1  g556(.A1(new_n554), .A2(new_n565), .ZN(new_n743));
  NAND4_X1  g557(.A1(new_n535), .A2(new_n557), .A3(new_n540), .A4(new_n743), .ZN(new_n744));
  OAI211_X1 g558(.A(new_n532), .B(new_n578), .C1(new_n744), .C2(new_n288), .ZN(new_n745));
  NOR2_X1   g559(.A1(new_n742), .A2(new_n745), .ZN(new_n746));
  NOR2_X1   g560(.A1(new_n577), .A2(new_n583), .ZN(new_n747));
  NOR2_X1   g561(.A1(new_n585), .A2(new_n652), .ZN(new_n748));
  NAND4_X1  g562(.A1(new_n620), .A2(new_n675), .A3(new_n747), .A4(new_n748), .ZN(new_n749));
  NAND4_X1  g563(.A1(new_n660), .A2(new_n588), .A3(new_n626), .A4(new_n749), .ZN(new_n750));
  INV_X1    g564(.A(KEYINPUT52), .ZN(new_n751));
  AND2_X1   g565(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  NOR2_X1   g566(.A1(new_n750), .A2(new_n751), .ZN(new_n753));
  OAI21_X1  g567(.A(new_n746), .B1(new_n752), .B2(new_n753), .ZN(new_n754));
  NOR3_X1   g568(.A1(new_n487), .A2(new_n530), .A3(new_n583), .ZN(new_n755));
  NAND3_X1  g569(.A1(new_n408), .A2(new_n581), .A3(new_n755), .ZN(new_n756));
  NOR2_X1   g570(.A1(new_n650), .A2(new_n539), .ZN(new_n757));
  NAND3_X1  g571(.A1(new_n675), .A2(new_n757), .A3(new_n625), .ZN(new_n758));
  NAND2_X1  g572(.A1(new_n756), .A2(new_n758), .ZN(new_n759));
  NAND3_X1  g573(.A1(new_n759), .A2(new_n577), .A3(new_n677), .ZN(new_n760));
  AOI21_X1  g574(.A(new_n663), .B1(new_n687), .B2(new_n680), .ZN(new_n761));
  NOR2_X1   g575(.A1(new_n679), .A2(new_n664), .ZN(new_n762));
  OAI211_X1 g576(.A(new_n691), .B(new_n760), .C1(new_n761), .C2(new_n762), .ZN(new_n763));
  OAI21_X1  g577(.A(new_n741), .B1(new_n754), .B2(new_n763), .ZN(new_n764));
  NAND2_X1  g578(.A1(new_n760), .A2(new_n691), .ZN(new_n765));
  AOI21_X1  g579(.A(new_n765), .B1(new_n688), .B2(new_n682), .ZN(new_n766));
  XNOR2_X1  g580(.A(new_n750), .B(new_n751), .ZN(new_n767));
  NAND4_X1  g581(.A1(new_n766), .A2(KEYINPUT53), .A3(new_n767), .A4(new_n746), .ZN(new_n768));
  NAND2_X1  g582(.A1(new_n764), .A2(new_n768), .ZN(new_n769));
  INV_X1    g583(.A(KEYINPUT54), .ZN(new_n770));
  NAND2_X1  g584(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  NAND3_X1  g585(.A1(new_n764), .A2(new_n768), .A3(KEYINPUT54), .ZN(new_n772));
  NAND2_X1  g586(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  AND3_X1   g587(.A1(new_n700), .A2(new_n491), .A3(new_n702), .ZN(new_n774));
  AND2_X1   g588(.A1(new_n774), .A2(new_n651), .ZN(new_n775));
  NAND2_X1  g589(.A1(new_n775), .A2(new_n645), .ZN(new_n776));
  NAND2_X1  g590(.A1(new_n737), .A2(new_n191), .ZN(new_n777));
  INV_X1    g591(.A(KEYINPUT46), .ZN(new_n778));
  AND2_X1   g592(.A1(new_n719), .A2(new_n720), .ZN(new_n779));
  OAI21_X1  g593(.A(new_n778), .B1(new_n779), .B2(new_n672), .ZN(new_n780));
  NAND3_X1  g594(.A1(new_n780), .A2(new_n593), .A3(new_n722), .ZN(new_n781));
  AOI21_X1  g595(.A(new_n730), .B1(new_n781), .B2(new_n595), .ZN(new_n782));
  INV_X1    g596(.A(new_n733), .ZN(new_n783));
  OAI21_X1  g597(.A(new_n777), .B1(new_n782), .B2(new_n783), .ZN(new_n784));
  NAND3_X1  g598(.A1(new_n784), .A2(new_n677), .A3(new_n775), .ZN(new_n785));
  NAND2_X1  g599(.A1(new_n609), .A2(new_n676), .ZN(new_n786));
  NAND3_X1  g600(.A1(new_n774), .A2(new_n632), .A3(new_n651), .ZN(new_n787));
  OAI21_X1  g601(.A(KEYINPUT113), .B1(new_n786), .B2(new_n787), .ZN(new_n788));
  NAND2_X1  g602(.A1(new_n788), .A2(KEYINPUT50), .ZN(new_n789));
  INV_X1    g603(.A(KEYINPUT50), .ZN(new_n790));
  OAI211_X1 g604(.A(KEYINPUT113), .B(new_n790), .C1(new_n786), .C2(new_n787), .ZN(new_n791));
  NAND2_X1  g605(.A1(new_n789), .A2(new_n791), .ZN(new_n792));
  NAND3_X1  g606(.A1(new_n632), .A2(new_n491), .A3(new_n677), .ZN(new_n793));
  NOR3_X1   g607(.A1(new_n793), .A2(new_n710), .A3(new_n711), .ZN(new_n794));
  INV_X1    g608(.A(KEYINPUT114), .ZN(new_n795));
  XNOR2_X1  g609(.A(new_n794), .B(new_n795), .ZN(new_n796));
  INV_X1    g610(.A(new_n657), .ZN(new_n797));
  OR2_X1    g611(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  OR3_X1    g612(.A1(new_n620), .A2(new_n448), .A3(new_n793), .ZN(new_n799));
  OR3_X1    g613(.A1(new_n799), .A2(new_n487), .A3(new_n553), .ZN(new_n800));
  NAND4_X1  g614(.A1(new_n785), .A2(new_n792), .A3(new_n798), .A4(new_n800), .ZN(new_n801));
  INV_X1    g615(.A(KEYINPUT115), .ZN(new_n802));
  AOI21_X1  g616(.A(KEYINPUT51), .B1(new_n785), .B2(new_n802), .ZN(new_n803));
  OAI21_X1  g617(.A(new_n488), .B1(new_n801), .B2(new_n803), .ZN(new_n804));
  AND2_X1   g618(.A1(new_n801), .A2(new_n803), .ZN(new_n805));
  NOR2_X1   g619(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  NAND3_X1  g620(.A1(new_n773), .A2(new_n776), .A3(new_n806), .ZN(new_n807));
  NOR2_X1   g621(.A1(new_n799), .A2(new_n554), .ZN(new_n808));
  INV_X1    g622(.A(new_n686), .ZN(new_n809));
  NOR2_X1   g623(.A1(new_n796), .A2(new_n809), .ZN(new_n810));
  XNOR2_X1  g624(.A(new_n810), .B(KEYINPUT48), .ZN(new_n811));
  NOR3_X1   g625(.A1(new_n807), .A2(new_n808), .A3(new_n811), .ZN(new_n812));
  NOR2_X1   g626(.A1(G952), .A2(G953), .ZN(new_n813));
  OAI21_X1  g627(.A(new_n740), .B1(new_n812), .B2(new_n813), .ZN(G75));
  NOR2_X1   g628(.A1(new_n334), .A2(G952), .ZN(new_n815));
  XOR2_X1   g629(.A(new_n815), .B(KEYINPUT116), .Z(new_n816));
  NAND2_X1  g630(.A1(new_n240), .A2(new_n269), .ZN(new_n817));
  XNOR2_X1  g631(.A(new_n817), .B(new_n267), .ZN(new_n818));
  XNOR2_X1  g632(.A(new_n818), .B(KEYINPUT55), .ZN(new_n819));
  AOI21_X1  g633(.A(new_n189), .B1(new_n764), .B2(new_n768), .ZN(new_n820));
  AOI211_X1 g634(.A(KEYINPUT56), .B(new_n819), .C1(new_n820), .C2(G210), .ZN(new_n821));
  INV_X1    g635(.A(new_n819), .ZN(new_n822));
  NAND3_X1  g636(.A1(new_n769), .A2(G210), .A3(G902), .ZN(new_n823));
  INV_X1    g637(.A(KEYINPUT56), .ZN(new_n824));
  AOI21_X1  g638(.A(new_n822), .B1(new_n823), .B2(new_n824), .ZN(new_n825));
  OAI21_X1  g639(.A(new_n816), .B1(new_n821), .B2(new_n825), .ZN(new_n826));
  INV_X1    g640(.A(KEYINPUT117), .ZN(new_n827));
  NAND2_X1  g641(.A1(new_n826), .A2(new_n827), .ZN(new_n828));
  OAI211_X1 g642(.A(KEYINPUT117), .B(new_n816), .C1(new_n821), .C2(new_n825), .ZN(new_n829));
  NAND2_X1  g643(.A1(new_n828), .A2(new_n829), .ZN(G51));
  XOR2_X1   g644(.A(new_n672), .B(KEYINPUT57), .Z(new_n831));
  OAI21_X1  g645(.A(new_n591), .B1(new_n773), .B2(new_n831), .ZN(new_n832));
  NAND2_X1  g646(.A1(new_n820), .A2(new_n779), .ZN(new_n833));
  AOI21_X1  g647(.A(new_n815), .B1(new_n832), .B2(new_n833), .ZN(G54));
  NAND2_X1  g648(.A1(new_n482), .A2(new_n466), .ZN(new_n835));
  INV_X1    g649(.A(new_n835), .ZN(new_n836));
  INV_X1    g650(.A(new_n820), .ZN(new_n837));
  INV_X1    g651(.A(KEYINPUT118), .ZN(new_n838));
  AND3_X1   g652(.A1(new_n838), .A2(KEYINPUT58), .A3(G475), .ZN(new_n839));
  OR2_X1    g653(.A1(new_n837), .A2(new_n839), .ZN(new_n840));
  AOI21_X1  g654(.A(new_n838), .B1(KEYINPUT58), .B2(G475), .ZN(new_n841));
  OAI21_X1  g655(.A(new_n836), .B1(new_n840), .B2(new_n841), .ZN(new_n842));
  OR4_X1    g656(.A1(new_n836), .A2(new_n837), .A3(new_n841), .A4(new_n839), .ZN(new_n843));
  INV_X1    g657(.A(new_n815), .ZN(new_n844));
  AND3_X1   g658(.A1(new_n842), .A2(new_n843), .A3(new_n844), .ZN(G60));
  NAND2_X1  g659(.A1(G478), .A2(G902), .ZN(new_n846));
  XNOR2_X1  g660(.A(new_n846), .B(KEYINPUT119), .ZN(new_n847));
  XNOR2_X1  g661(.A(new_n847), .B(KEYINPUT59), .ZN(new_n848));
  NAND3_X1  g662(.A1(new_n771), .A2(new_n772), .A3(new_n848), .ZN(new_n849));
  NAND2_X1  g663(.A1(new_n544), .A2(new_n545), .ZN(new_n850));
  NAND2_X1  g664(.A1(new_n849), .A2(new_n850), .ZN(new_n851));
  INV_X1    g665(.A(new_n850), .ZN(new_n852));
  NAND4_X1  g666(.A1(new_n771), .A2(new_n852), .A3(new_n772), .A4(new_n848), .ZN(new_n853));
  NAND3_X1  g667(.A1(new_n851), .A2(new_n816), .A3(new_n853), .ZN(new_n854));
  INV_X1    g668(.A(KEYINPUT120), .ZN(new_n855));
  NAND2_X1  g669(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  NAND4_X1  g670(.A1(new_n851), .A2(KEYINPUT120), .A3(new_n816), .A4(new_n853), .ZN(new_n857));
  NAND2_X1  g671(.A1(new_n856), .A2(new_n857), .ZN(G63));
  NAND2_X1  g672(.A1(G217), .A2(G902), .ZN(new_n859));
  XOR2_X1   g673(.A(new_n859), .B(KEYINPUT60), .Z(new_n860));
  NAND2_X1  g674(.A1(new_n769), .A2(new_n860), .ZN(new_n861));
  NAND2_X1  g675(.A1(new_n861), .A2(new_n438), .ZN(new_n862));
  NAND2_X1  g676(.A1(new_n574), .A2(new_n575), .ZN(new_n863));
  XOR2_X1   g677(.A(new_n863), .B(KEYINPUT121), .Z(new_n864));
  OAI211_X1 g678(.A(new_n862), .B(new_n816), .C1(new_n861), .C2(new_n864), .ZN(new_n865));
  INV_X1    g679(.A(KEYINPUT61), .ZN(new_n866));
  XNOR2_X1  g680(.A(new_n865), .B(new_n866), .ZN(G66));
  OAI21_X1  g681(.A(G953), .B1(new_n493), .B2(new_n264), .ZN(new_n868));
  OAI21_X1  g682(.A(new_n868), .B1(new_n746), .B2(G953), .ZN(new_n869));
  OAI21_X1  g683(.A(new_n817), .B1(G898), .B2(new_n334), .ZN(new_n870));
  XOR2_X1   g684(.A(new_n870), .B(KEYINPUT122), .Z(new_n871));
  XNOR2_X1  g685(.A(new_n869), .B(new_n871), .ZN(G69));
  AND2_X1   g686(.A1(new_n588), .A2(new_n626), .ZN(new_n873));
  NAND2_X1  g687(.A1(new_n873), .A2(new_n660), .ZN(new_n874));
  AOI21_X1  g688(.A(new_n874), .B1(new_n688), .B2(new_n682), .ZN(new_n875));
  NAND3_X1  g689(.A1(new_n726), .A2(new_n686), .A3(new_n748), .ZN(new_n876));
  NAND2_X1  g690(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  NAND3_X1  g691(.A1(new_n727), .A2(new_n691), .A3(new_n735), .ZN(new_n878));
  OAI21_X1  g692(.A(KEYINPUT123), .B1(new_n877), .B2(new_n878), .ZN(new_n879));
  AND3_X1   g693(.A1(new_n727), .A2(new_n691), .A3(new_n735), .ZN(new_n880));
  INV_X1    g694(.A(KEYINPUT123), .ZN(new_n881));
  NAND4_X1  g695(.A1(new_n880), .A2(new_n881), .A3(new_n875), .A4(new_n876), .ZN(new_n882));
  NAND3_X1  g696(.A1(new_n879), .A2(new_n882), .A3(new_n334), .ZN(new_n883));
  NAND2_X1  g697(.A1(new_n386), .A2(new_n387), .ZN(new_n884));
  XOR2_X1   g698(.A(new_n884), .B(new_n478), .Z(new_n885));
  NAND2_X1  g699(.A1(G900), .A2(G953), .ZN(new_n886));
  NAND3_X1  g700(.A1(new_n883), .A2(new_n885), .A3(new_n886), .ZN(new_n887));
  AOI21_X1  g701(.A(new_n334), .B1(G227), .B2(G900), .ZN(new_n888));
  NAND2_X1  g702(.A1(new_n888), .A2(KEYINPUT124), .ZN(new_n889));
  INV_X1    g703(.A(new_n885), .ZN(new_n890));
  INV_X1    g704(.A(KEYINPUT62), .ZN(new_n891));
  AND3_X1   g705(.A1(new_n602), .A2(new_n613), .A3(new_n620), .ZN(new_n892));
  OAI21_X1  g706(.A(new_n891), .B1(new_n892), .B2(new_n874), .ZN(new_n893));
  NAND4_X1  g707(.A1(new_n621), .A2(KEYINPUT62), .A3(new_n660), .A4(new_n873), .ZN(new_n894));
  NAND2_X1  g708(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  NAND4_X1  g709(.A1(new_n686), .A2(new_n598), .A3(new_n677), .A4(new_n743), .ZN(new_n896));
  AND2_X1   g710(.A1(new_n727), .A2(new_n735), .ZN(new_n897));
  AND3_X1   g711(.A1(new_n895), .A2(new_n896), .A3(new_n897), .ZN(new_n898));
  OAI21_X1  g712(.A(new_n890), .B1(new_n898), .B2(G953), .ZN(new_n899));
  NAND3_X1  g713(.A1(new_n887), .A2(new_n889), .A3(new_n899), .ZN(new_n900));
  NOR2_X1   g714(.A1(new_n888), .A2(KEYINPUT124), .ZN(new_n901));
  XOR2_X1   g715(.A(new_n900), .B(new_n901), .Z(G72));
  NAND3_X1  g716(.A1(new_n879), .A2(new_n882), .A3(new_n746), .ZN(new_n903));
  XNOR2_X1  g717(.A(KEYINPUT125), .B(KEYINPUT63), .ZN(new_n904));
  NAND2_X1  g718(.A1(G472), .A2(G902), .ZN(new_n905));
  XNOR2_X1  g719(.A(new_n904), .B(new_n905), .ZN(new_n906));
  AOI211_X1 g720(.A(new_n378), .B(new_n389), .C1(new_n903), .C2(new_n906), .ZN(new_n907));
  OAI21_X1  g721(.A(KEYINPUT127), .B1(new_n907), .B2(new_n815), .ZN(new_n908));
  INV_X1    g722(.A(new_n391), .ZN(new_n909));
  NAND2_X1  g723(.A1(new_n909), .A2(new_n398), .ZN(new_n910));
  AND3_X1   g724(.A1(new_n769), .A2(new_n906), .A3(new_n910), .ZN(new_n911));
  NAND4_X1  g725(.A1(new_n895), .A2(new_n746), .A3(new_n896), .A4(new_n897), .ZN(new_n912));
  AOI21_X1  g726(.A(KEYINPUT126), .B1(new_n912), .B2(new_n906), .ZN(new_n913));
  NOR3_X1   g727(.A1(new_n913), .A2(new_n379), .A3(new_n390), .ZN(new_n914));
  NAND3_X1  g728(.A1(new_n912), .A2(KEYINPUT126), .A3(new_n906), .ZN(new_n915));
  AOI21_X1  g729(.A(new_n911), .B1(new_n914), .B2(new_n915), .ZN(new_n916));
  NAND2_X1  g730(.A1(new_n903), .A2(new_n906), .ZN(new_n917));
  NAND3_X1  g731(.A1(new_n917), .A2(new_n379), .A3(new_n390), .ZN(new_n918));
  INV_X1    g732(.A(KEYINPUT127), .ZN(new_n919));
  NAND3_X1  g733(.A1(new_n918), .A2(new_n919), .A3(new_n844), .ZN(new_n920));
  AND3_X1   g734(.A1(new_n908), .A2(new_n916), .A3(new_n920), .ZN(G57));
endmodule


