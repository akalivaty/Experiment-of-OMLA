//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 1 1 0 0 1 1 0 0 0 1 1 1 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 0 1 0 0 0 1 1 1 1 0 0 0 0 0 1 0 1 0 0 0 0 0 0 1 0 1 1 1 1 0 0 1 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:20:17 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n634, new_n635, new_n636, new_n637,
    new_n639, new_n640, new_n641, new_n642, new_n643, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n675,
    new_n676, new_n677, new_n678, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n708, new_n709, new_n710, new_n712, new_n713, new_n714,
    new_n716, new_n717, new_n718, new_n719, new_n720, new_n722, new_n724,
    new_n725, new_n726, new_n727, new_n728, new_n729, new_n730, new_n731,
    new_n732, new_n733, new_n734, new_n735, new_n736, new_n737, new_n738,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n812, new_n813,
    new_n814, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n823, new_n824, new_n825, new_n826, new_n827, new_n828, new_n829,
    new_n830, new_n831, new_n832, new_n833, new_n834, new_n835, new_n836,
    new_n837, new_n838, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n877, new_n878, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n897, new_n898,
    new_n900, new_n901, new_n902, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n935, new_n936, new_n937, new_n938,
    new_n940, new_n941;
  XNOR2_X1  g000(.A(G57gat), .B(G64gat), .ZN(new_n202));
  AOI21_X1  g001(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n203));
  OR2_X1    g002(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  XOR2_X1   g003(.A(G71gat), .B(G78gat), .Z(new_n205));
  XNOR2_X1  g004(.A(new_n204), .B(new_n205), .ZN(new_n206));
  INV_X1    g005(.A(KEYINPUT21), .ZN(new_n207));
  NAND2_X1  g006(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  NAND2_X1  g007(.A1(G231gat), .A2(G233gat), .ZN(new_n209));
  XNOR2_X1  g008(.A(new_n208), .B(new_n209), .ZN(new_n210));
  XNOR2_X1  g009(.A(KEYINPUT91), .B(KEYINPUT19), .ZN(new_n211));
  XNOR2_X1  g010(.A(new_n210), .B(new_n211), .ZN(new_n212));
  XNOR2_X1  g011(.A(G127gat), .B(G155gat), .ZN(new_n213));
  XNOR2_X1  g012(.A(new_n212), .B(new_n213), .ZN(new_n214));
  XOR2_X1   g013(.A(G183gat), .B(G211gat), .Z(new_n215));
  NAND2_X1  g014(.A1(new_n214), .A2(new_n215), .ZN(new_n216));
  OR2_X1    g015(.A1(new_n212), .A2(new_n213), .ZN(new_n217));
  INV_X1    g016(.A(new_n215), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n212), .A2(new_n213), .ZN(new_n219));
  NAND3_X1  g018(.A1(new_n217), .A2(new_n218), .A3(new_n219), .ZN(new_n220));
  XNOR2_X1  g019(.A(G15gat), .B(G22gat), .ZN(new_n221));
  INV_X1    g020(.A(KEYINPUT88), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  XNOR2_X1  g022(.A(new_n223), .B(G8gat), .ZN(new_n224));
  INV_X1    g023(.A(KEYINPUT16), .ZN(new_n225));
  AOI21_X1  g024(.A(G1gat), .B1(new_n221), .B2(new_n225), .ZN(new_n226));
  XNOR2_X1  g025(.A(new_n224), .B(new_n226), .ZN(new_n227));
  INV_X1    g026(.A(new_n206), .ZN(new_n228));
  AOI21_X1  g027(.A(new_n227), .B1(KEYINPUT21), .B2(new_n228), .ZN(new_n229));
  XNOR2_X1  g028(.A(KEYINPUT92), .B(KEYINPUT20), .ZN(new_n230));
  XNOR2_X1  g029(.A(new_n229), .B(new_n230), .ZN(new_n231));
  AND3_X1   g030(.A1(new_n216), .A2(new_n220), .A3(new_n231), .ZN(new_n232));
  AOI21_X1  g031(.A(new_n231), .B1(new_n216), .B2(new_n220), .ZN(new_n233));
  NOR2_X1   g032(.A1(new_n232), .A2(new_n233), .ZN(new_n234));
  XNOR2_X1  g033(.A(G190gat), .B(G218gat), .ZN(new_n235));
  XNOR2_X1  g034(.A(new_n235), .B(KEYINPUT95), .ZN(new_n236));
  INV_X1    g035(.A(new_n236), .ZN(new_n237));
  NAND2_X1  g036(.A1(G85gat), .A2(G92gat), .ZN(new_n238));
  NAND2_X1  g037(.A1(KEYINPUT94), .A2(KEYINPUT7), .ZN(new_n239));
  XOR2_X1   g038(.A(new_n238), .B(new_n239), .Z(new_n240));
  NAND2_X1  g039(.A1(G99gat), .A2(G106gat), .ZN(new_n241));
  INV_X1    g040(.A(G85gat), .ZN(new_n242));
  INV_X1    g041(.A(G92gat), .ZN(new_n243));
  AOI22_X1  g042(.A1(KEYINPUT8), .A2(new_n241), .B1(new_n242), .B2(new_n243), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n240), .A2(new_n244), .ZN(new_n245));
  XNOR2_X1  g044(.A(G99gat), .B(G106gat), .ZN(new_n246));
  XNOR2_X1  g045(.A(new_n245), .B(new_n246), .ZN(new_n247));
  INV_X1    g046(.A(G29gat), .ZN(new_n248));
  NAND3_X1  g047(.A1(new_n248), .A2(KEYINPUT14), .A3(G36gat), .ZN(new_n249));
  XOR2_X1   g048(.A(KEYINPUT14), .B(G29gat), .Z(new_n250));
  OAI21_X1  g049(.A(new_n249), .B1(new_n250), .B2(G36gat), .ZN(new_n251));
  XNOR2_X1  g050(.A(G43gat), .B(G50gat), .ZN(new_n252));
  AOI22_X1  g051(.A1(new_n251), .A2(KEYINPUT87), .B1(KEYINPUT15), .B2(new_n252), .ZN(new_n253));
  OAI21_X1  g052(.A(new_n251), .B1(KEYINPUT15), .B2(new_n252), .ZN(new_n254));
  OR2_X1    g053(.A1(new_n253), .A2(new_n254), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n253), .A2(new_n254), .ZN(new_n256));
  NAND2_X1  g055(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  INV_X1    g056(.A(KEYINPUT17), .ZN(new_n258));
  NAND2_X1  g057(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  NAND3_X1  g058(.A1(new_n255), .A2(KEYINPUT17), .A3(new_n256), .ZN(new_n260));
  AOI21_X1  g059(.A(new_n247), .B1(new_n259), .B2(new_n260), .ZN(new_n261));
  AND2_X1   g060(.A1(G232gat), .A2(G233gat), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n262), .A2(KEYINPUT41), .ZN(new_n263));
  XOR2_X1   g062(.A(new_n245), .B(new_n246), .Z(new_n264));
  OAI21_X1  g063(.A(new_n263), .B1(new_n257), .B2(new_n264), .ZN(new_n265));
  OAI21_X1  g064(.A(new_n237), .B1(new_n261), .B2(new_n265), .ZN(new_n266));
  OR2_X1    g065(.A1(new_n266), .A2(KEYINPUT97), .ZN(new_n267));
  NOR2_X1   g066(.A1(new_n261), .A2(new_n265), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n268), .A2(new_n236), .ZN(new_n269));
  NOR2_X1   g068(.A1(new_n262), .A2(KEYINPUT41), .ZN(new_n270));
  XNOR2_X1  g069(.A(G134gat), .B(G162gat), .ZN(new_n271));
  XOR2_X1   g070(.A(new_n270), .B(new_n271), .Z(new_n272));
  INV_X1    g071(.A(new_n272), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n266), .A2(KEYINPUT97), .ZN(new_n274));
  NAND4_X1  g073(.A1(new_n267), .A2(new_n269), .A3(new_n273), .A4(new_n274), .ZN(new_n275));
  NAND2_X1  g074(.A1(new_n269), .A2(new_n266), .ZN(new_n276));
  XOR2_X1   g075(.A(new_n272), .B(KEYINPUT93), .Z(new_n277));
  AOI21_X1  g076(.A(KEYINPUT96), .B1(new_n276), .B2(new_n277), .ZN(new_n278));
  INV_X1    g077(.A(KEYINPUT96), .ZN(new_n279));
  INV_X1    g078(.A(new_n277), .ZN(new_n280));
  AOI211_X1 g079(.A(new_n279), .B(new_n280), .C1(new_n269), .C2(new_n266), .ZN(new_n281));
  OAI21_X1  g080(.A(new_n275), .B1(new_n278), .B2(new_n281), .ZN(new_n282));
  INV_X1    g081(.A(new_n282), .ZN(new_n283));
  XNOR2_X1  g082(.A(G113gat), .B(G141gat), .ZN(new_n284));
  XNOR2_X1  g083(.A(new_n284), .B(G197gat), .ZN(new_n285));
  XOR2_X1   g084(.A(KEYINPUT11), .B(G169gat), .Z(new_n286));
  XNOR2_X1  g085(.A(new_n285), .B(new_n286), .ZN(new_n287));
  XOR2_X1   g086(.A(new_n287), .B(KEYINPUT12), .Z(new_n288));
  INV_X1    g087(.A(new_n227), .ZN(new_n289));
  NOR2_X1   g088(.A1(new_n289), .A2(new_n257), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n259), .A2(new_n260), .ZN(new_n291));
  AOI21_X1  g090(.A(new_n290), .B1(new_n291), .B2(new_n289), .ZN(new_n292));
  NAND2_X1  g091(.A1(G229gat), .A2(G233gat), .ZN(new_n293));
  XOR2_X1   g092(.A(new_n293), .B(KEYINPUT89), .Z(new_n294));
  INV_X1    g093(.A(KEYINPUT18), .ZN(new_n295));
  NAND2_X1  g094(.A1(new_n295), .A2(KEYINPUT90), .ZN(new_n296));
  NAND3_X1  g095(.A1(new_n292), .A2(new_n294), .A3(new_n296), .ZN(new_n297));
  XNOR2_X1  g096(.A(new_n289), .B(new_n257), .ZN(new_n298));
  XOR2_X1   g097(.A(new_n294), .B(KEYINPUT13), .Z(new_n299));
  NAND2_X1  g098(.A1(new_n298), .A2(new_n299), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n297), .A2(new_n300), .ZN(new_n301));
  AOI21_X1  g100(.A(new_n296), .B1(new_n292), .B2(new_n294), .ZN(new_n302));
  OAI21_X1  g101(.A(new_n288), .B1(new_n301), .B2(new_n302), .ZN(new_n303));
  INV_X1    g102(.A(new_n302), .ZN(new_n304));
  INV_X1    g103(.A(new_n288), .ZN(new_n305));
  NAND4_X1  g104(.A1(new_n304), .A2(new_n305), .A3(new_n300), .A4(new_n297), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n303), .A2(new_n306), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n264), .A2(new_n206), .ZN(new_n308));
  INV_X1    g107(.A(KEYINPUT10), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n247), .A2(new_n228), .ZN(new_n310));
  NAND3_X1  g109(.A1(new_n308), .A2(new_n309), .A3(new_n310), .ZN(new_n311));
  NAND3_X1  g110(.A1(new_n247), .A2(new_n228), .A3(KEYINPUT10), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  NAND2_X1  g112(.A1(G230gat), .A2(G233gat), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n313), .A2(new_n314), .ZN(new_n315));
  XNOR2_X1  g114(.A(G120gat), .B(G148gat), .ZN(new_n316));
  XNOR2_X1  g115(.A(G176gat), .B(G204gat), .ZN(new_n317));
  XOR2_X1   g116(.A(new_n316), .B(new_n317), .Z(new_n318));
  INV_X1    g117(.A(new_n318), .ZN(new_n319));
  AOI21_X1  g118(.A(new_n314), .B1(new_n308), .B2(new_n310), .ZN(new_n320));
  AOI21_X1  g119(.A(new_n319), .B1(new_n320), .B2(KEYINPUT98), .ZN(new_n321));
  OAI211_X1 g120(.A(new_n315), .B(new_n321), .C1(KEYINPUT98), .C2(new_n320), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n315), .A2(KEYINPUT99), .ZN(new_n323));
  INV_X1    g122(.A(KEYINPUT99), .ZN(new_n324));
  NAND3_X1  g123(.A1(new_n313), .A2(new_n324), .A3(new_n314), .ZN(new_n325));
  AOI21_X1  g124(.A(new_n320), .B1(new_n323), .B2(new_n325), .ZN(new_n326));
  OAI21_X1  g125(.A(new_n322), .B1(new_n326), .B2(new_n318), .ZN(new_n327));
  INV_X1    g126(.A(new_n327), .ZN(new_n328));
  NAND4_X1  g127(.A1(new_n234), .A2(new_n283), .A3(new_n307), .A4(new_n328), .ZN(new_n329));
  INV_X1    g128(.A(G228gat), .ZN(new_n330));
  INV_X1    g129(.A(G233gat), .ZN(new_n331));
  NOR2_X1   g130(.A1(new_n330), .A2(new_n331), .ZN(new_n332));
  INV_X1    g131(.A(KEYINPUT3), .ZN(new_n333));
  OR2_X1    g132(.A1(G141gat), .A2(G148gat), .ZN(new_n334));
  INV_X1    g133(.A(KEYINPUT2), .ZN(new_n335));
  NAND2_X1  g134(.A1(G141gat), .A2(G148gat), .ZN(new_n336));
  NAND3_X1  g135(.A1(new_n334), .A2(new_n335), .A3(new_n336), .ZN(new_n337));
  INV_X1    g136(.A(G162gat), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n338), .A2(G155gat), .ZN(new_n339));
  INV_X1    g138(.A(G155gat), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n340), .A2(G162gat), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n339), .A2(new_n341), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n337), .A2(new_n342), .ZN(new_n343));
  XNOR2_X1  g142(.A(KEYINPUT75), .B(G162gat), .ZN(new_n344));
  AOI21_X1  g143(.A(new_n335), .B1(new_n344), .B2(G155gat), .ZN(new_n345));
  NAND4_X1  g144(.A1(new_n334), .A2(new_n339), .A3(new_n341), .A4(new_n336), .ZN(new_n346));
  OAI211_X1 g145(.A(new_n333), .B(new_n343), .C1(new_n345), .C2(new_n346), .ZN(new_n347));
  INV_X1    g146(.A(KEYINPUT29), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n347), .A2(new_n348), .ZN(new_n349));
  AND2_X1   g148(.A1(G211gat), .A2(G218gat), .ZN(new_n350));
  NOR2_X1   g149(.A1(G211gat), .A2(G218gat), .ZN(new_n351));
  NOR2_X1   g150(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  AND2_X1   g151(.A1(G197gat), .A2(G204gat), .ZN(new_n353));
  NOR2_X1   g152(.A1(G197gat), .A2(G204gat), .ZN(new_n354));
  NOR2_X1   g153(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  AOI21_X1  g154(.A(KEYINPUT22), .B1(G211gat), .B2(G218gat), .ZN(new_n356));
  OAI21_X1  g155(.A(new_n352), .B1(new_n355), .B2(new_n356), .ZN(new_n357));
  XNOR2_X1  g156(.A(G211gat), .B(G218gat), .ZN(new_n358));
  XNOR2_X1  g157(.A(G197gat), .B(G204gat), .ZN(new_n359));
  INV_X1    g158(.A(new_n356), .ZN(new_n360));
  NAND3_X1  g159(.A1(new_n358), .A2(new_n359), .A3(new_n360), .ZN(new_n361));
  NAND3_X1  g160(.A1(new_n357), .A2(new_n361), .A3(KEYINPUT71), .ZN(new_n362));
  INV_X1    g161(.A(KEYINPUT71), .ZN(new_n363));
  OAI211_X1 g162(.A(new_n363), .B(new_n352), .C1(new_n355), .C2(new_n356), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n362), .A2(new_n364), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n349), .A2(new_n365), .ZN(new_n366));
  OAI21_X1  g165(.A(new_n343), .B1(new_n345), .B2(new_n346), .ZN(new_n367));
  AOI21_X1  g166(.A(KEYINPUT29), .B1(new_n357), .B2(new_n361), .ZN(new_n368));
  OAI21_X1  g167(.A(new_n367), .B1(new_n368), .B2(KEYINPUT3), .ZN(new_n369));
  AOI21_X1  g168(.A(new_n332), .B1(new_n366), .B2(new_n369), .ZN(new_n370));
  INV_X1    g169(.A(KEYINPUT78), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n366), .A2(new_n332), .ZN(new_n372));
  AND2_X1   g171(.A1(KEYINPUT75), .A2(G162gat), .ZN(new_n373));
  NOR2_X1   g172(.A1(KEYINPUT75), .A2(G162gat), .ZN(new_n374));
  OAI21_X1  g173(.A(G155gat), .B1(new_n373), .B2(new_n374), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n375), .A2(KEYINPUT2), .ZN(new_n376));
  AND4_X1   g175(.A1(new_n339), .A2(new_n334), .A3(new_n341), .A4(new_n336), .ZN(new_n377));
  AOI22_X1  g176(.A1(new_n376), .A2(new_n377), .B1(new_n342), .B2(new_n337), .ZN(new_n378));
  NAND3_X1  g177(.A1(new_n362), .A2(new_n348), .A3(new_n364), .ZN(new_n379));
  AOI21_X1  g178(.A(new_n378), .B1(new_n379), .B2(new_n333), .ZN(new_n380));
  OAI21_X1  g179(.A(new_n371), .B1(new_n372), .B2(new_n380), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n379), .A2(new_n333), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n382), .A2(new_n367), .ZN(new_n383));
  INV_X1    g182(.A(new_n332), .ZN(new_n384));
  AOI21_X1  g183(.A(new_n384), .B1(new_n349), .B2(new_n365), .ZN(new_n385));
  NAND3_X1  g184(.A1(new_n383), .A2(KEYINPUT78), .A3(new_n385), .ZN(new_n386));
  AOI211_X1 g185(.A(G22gat), .B(new_n370), .C1(new_n381), .C2(new_n386), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n387), .A2(KEYINPUT80), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n381), .A2(new_n386), .ZN(new_n389));
  INV_X1    g188(.A(G22gat), .ZN(new_n390));
  INV_X1    g189(.A(new_n370), .ZN(new_n391));
  NAND3_X1  g190(.A1(new_n389), .A2(new_n390), .A3(new_n391), .ZN(new_n392));
  INV_X1    g191(.A(KEYINPUT80), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n392), .A2(new_n393), .ZN(new_n394));
  AOI22_X1  g193(.A1(new_n347), .A2(new_n348), .B1(new_n362), .B2(new_n364), .ZN(new_n395));
  NOR4_X1   g194(.A1(new_n380), .A2(new_n395), .A3(new_n371), .A4(new_n384), .ZN(new_n396));
  AOI21_X1  g195(.A(KEYINPUT78), .B1(new_n383), .B2(new_n385), .ZN(new_n397));
  OAI21_X1  g196(.A(new_n391), .B1(new_n396), .B2(new_n397), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n398), .A2(G22gat), .ZN(new_n399));
  XNOR2_X1  g198(.A(G78gat), .B(G106gat), .ZN(new_n400));
  XNOR2_X1  g199(.A(KEYINPUT31), .B(G50gat), .ZN(new_n401));
  XOR2_X1   g200(.A(new_n400), .B(new_n401), .Z(new_n402));
  INV_X1    g201(.A(new_n402), .ZN(new_n403));
  NAND4_X1  g202(.A1(new_n388), .A2(new_n394), .A3(new_n399), .A4(new_n403), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n399), .A2(new_n392), .ZN(new_n405));
  XOR2_X1   g204(.A(new_n402), .B(KEYINPUT77), .Z(new_n406));
  INV_X1    g205(.A(new_n406), .ZN(new_n407));
  AOI21_X1  g206(.A(KEYINPUT79), .B1(new_n405), .B2(new_n407), .ZN(new_n408));
  INV_X1    g207(.A(KEYINPUT79), .ZN(new_n409));
  AOI211_X1 g208(.A(new_n409), .B(new_n406), .C1(new_n399), .C2(new_n392), .ZN(new_n410));
  OAI21_X1  g209(.A(new_n404), .B1(new_n408), .B2(new_n410), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n411), .A2(KEYINPUT81), .ZN(new_n412));
  NOR2_X1   g211(.A1(G169gat), .A2(G176gat), .ZN(new_n413));
  INV_X1    g212(.A(new_n413), .ZN(new_n414));
  OR2_X1    g213(.A1(new_n414), .A2(KEYINPUT26), .ZN(new_n415));
  NAND2_X1  g214(.A1(G169gat), .A2(G176gat), .ZN(new_n416));
  INV_X1    g215(.A(new_n416), .ZN(new_n417));
  AOI21_X1  g216(.A(new_n417), .B1(new_n414), .B2(KEYINPUT26), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n415), .A2(new_n418), .ZN(new_n419));
  NAND2_X1  g218(.A1(G183gat), .A2(G190gat), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  INV_X1    g220(.A(KEYINPUT27), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n422), .A2(G183gat), .ZN(new_n423));
  NOR2_X1   g222(.A1(KEYINPUT28), .A2(G190gat), .ZN(new_n424));
  XNOR2_X1  g223(.A(KEYINPUT66), .B(G183gat), .ZN(new_n425));
  OAI211_X1 g224(.A(new_n423), .B(new_n424), .C1(new_n425), .C2(new_n422), .ZN(new_n426));
  INV_X1    g225(.A(G183gat), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n427), .A2(KEYINPUT27), .ZN(new_n428));
  INV_X1    g227(.A(G190gat), .ZN(new_n429));
  NAND3_X1  g228(.A1(new_n423), .A2(new_n428), .A3(new_n429), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n430), .A2(KEYINPUT28), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n426), .A2(new_n431), .ZN(new_n432));
  INV_X1    g231(.A(KEYINPUT67), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n432), .A2(new_n433), .ZN(new_n434));
  NAND3_X1  g233(.A1(new_n426), .A2(KEYINPUT67), .A3(new_n431), .ZN(new_n435));
  AOI21_X1  g234(.A(new_n421), .B1(new_n434), .B2(new_n435), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n420), .A2(KEYINPUT24), .ZN(new_n437));
  INV_X1    g236(.A(KEYINPUT24), .ZN(new_n438));
  NAND3_X1  g237(.A1(new_n438), .A2(G183gat), .A3(G190gat), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n437), .A2(new_n439), .ZN(new_n440));
  OAI21_X1  g239(.A(new_n440), .B1(new_n425), .B2(G190gat), .ZN(new_n441));
  XNOR2_X1  g240(.A(new_n416), .B(KEYINPUT65), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n413), .A2(KEYINPUT23), .ZN(new_n443));
  INV_X1    g242(.A(KEYINPUT23), .ZN(new_n444));
  OAI21_X1  g243(.A(new_n444), .B1(G169gat), .B2(G176gat), .ZN(new_n445));
  AND2_X1   g244(.A1(new_n443), .A2(new_n445), .ZN(new_n446));
  NAND3_X1  g245(.A1(new_n441), .A2(new_n442), .A3(new_n446), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n447), .A2(KEYINPUT25), .ZN(new_n448));
  NOR2_X1   g247(.A1(new_n443), .A2(KEYINPUT64), .ZN(new_n449));
  INV_X1    g248(.A(KEYINPUT25), .ZN(new_n450));
  NAND3_X1  g249(.A1(new_n445), .A2(new_n450), .A3(new_n416), .ZN(new_n451));
  INV_X1    g250(.A(KEYINPUT64), .ZN(new_n452));
  AOI21_X1  g251(.A(new_n452), .B1(new_n413), .B2(KEYINPUT23), .ZN(new_n453));
  NOR3_X1   g252(.A1(new_n449), .A2(new_n451), .A3(new_n453), .ZN(new_n454));
  OAI21_X1  g253(.A(new_n440), .B1(G183gat), .B2(G190gat), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n448), .A2(new_n456), .ZN(new_n457));
  INV_X1    g256(.A(G226gat), .ZN(new_n458));
  NOR2_X1   g257(.A1(new_n458), .A2(new_n331), .ZN(new_n459));
  NOR3_X1   g258(.A1(new_n436), .A2(new_n457), .A3(new_n459), .ZN(new_n460));
  NOR2_X1   g259(.A1(new_n459), .A2(KEYINPUT29), .ZN(new_n461));
  AND2_X1   g260(.A1(new_n419), .A2(new_n420), .ZN(new_n462));
  AND3_X1   g261(.A1(new_n426), .A2(KEYINPUT67), .A3(new_n431), .ZN(new_n463));
  AOI21_X1  g262(.A(KEYINPUT67), .B1(new_n426), .B2(new_n431), .ZN(new_n464));
  OAI21_X1  g263(.A(new_n462), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  AOI22_X1  g264(.A1(new_n447), .A2(KEYINPUT25), .B1(new_n454), .B2(new_n455), .ZN(new_n466));
  AOI21_X1  g265(.A(new_n461), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  OAI21_X1  g266(.A(new_n365), .B1(new_n460), .B2(new_n467), .ZN(new_n468));
  INV_X1    g267(.A(KEYINPUT72), .ZN(new_n469));
  OAI22_X1  g268(.A1(new_n436), .A2(new_n457), .B1(KEYINPUT29), .B2(new_n459), .ZN(new_n470));
  OAI211_X1 g269(.A(new_n465), .B(new_n466), .C1(new_n458), .C2(new_n331), .ZN(new_n471));
  INV_X1    g270(.A(new_n365), .ZN(new_n472));
  NAND3_X1  g271(.A1(new_n470), .A2(new_n471), .A3(new_n472), .ZN(new_n473));
  NAND3_X1  g272(.A1(new_n468), .A2(new_n469), .A3(new_n473), .ZN(new_n474));
  NAND4_X1  g273(.A1(new_n470), .A2(new_n471), .A3(KEYINPUT72), .A4(new_n472), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  XNOR2_X1  g275(.A(G8gat), .B(G36gat), .ZN(new_n477));
  XNOR2_X1  g276(.A(G64gat), .B(G92gat), .ZN(new_n478));
  XNOR2_X1  g277(.A(new_n477), .B(new_n478), .ZN(new_n479));
  XNOR2_X1  g278(.A(KEYINPUT73), .B(KEYINPUT74), .ZN(new_n480));
  XOR2_X1   g279(.A(new_n479), .B(new_n480), .Z(new_n481));
  NAND2_X1  g280(.A1(new_n476), .A2(new_n481), .ZN(new_n482));
  INV_X1    g281(.A(new_n481), .ZN(new_n483));
  NAND3_X1  g282(.A1(new_n474), .A2(new_n475), .A3(new_n483), .ZN(new_n484));
  NAND3_X1  g283(.A1(new_n482), .A2(KEYINPUT30), .A3(new_n484), .ZN(new_n485));
  INV_X1    g284(.A(KEYINPUT30), .ZN(new_n486));
  NAND3_X1  g285(.A1(new_n476), .A2(new_n486), .A3(new_n481), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n485), .A2(new_n487), .ZN(new_n488));
  NAND2_X1  g287(.A1(new_n367), .A2(KEYINPUT3), .ZN(new_n489));
  INV_X1    g288(.A(KEYINPUT68), .ZN(new_n490));
  INV_X1    g289(.A(KEYINPUT1), .ZN(new_n491));
  OAI21_X1  g290(.A(new_n491), .B1(G113gat), .B2(G120gat), .ZN(new_n492));
  AND2_X1   g291(.A1(G113gat), .A2(G120gat), .ZN(new_n493));
  OAI21_X1  g292(.A(new_n490), .B1(new_n492), .B2(new_n493), .ZN(new_n494));
  XNOR2_X1  g293(.A(G127gat), .B(G134gat), .ZN(new_n495));
  INV_X1    g294(.A(new_n495), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n494), .A2(new_n496), .ZN(new_n497));
  OAI211_X1 g296(.A(new_n495), .B(new_n490), .C1(new_n493), .C2(new_n492), .ZN(new_n498));
  AND2_X1   g297(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  NAND3_X1  g298(.A1(new_n489), .A2(new_n499), .A3(new_n347), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n497), .A2(new_n498), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n378), .A2(new_n501), .ZN(new_n502));
  INV_X1    g301(.A(KEYINPUT4), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  NAND3_X1  g303(.A1(new_n378), .A2(KEYINPUT4), .A3(new_n501), .ZN(new_n505));
  NAND3_X1  g304(.A1(new_n500), .A2(new_n504), .A3(new_n505), .ZN(new_n506));
  NAND2_X1  g305(.A1(G225gat), .A2(G233gat), .ZN(new_n507));
  INV_X1    g306(.A(new_n507), .ZN(new_n508));
  INV_X1    g307(.A(KEYINPUT5), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n499), .A2(new_n367), .ZN(new_n510));
  AOI21_X1  g309(.A(new_n507), .B1(new_n510), .B2(new_n502), .ZN(new_n511));
  OAI22_X1  g310(.A1(new_n506), .A2(new_n508), .B1(new_n509), .B2(new_n511), .ZN(new_n512));
  INV_X1    g311(.A(new_n505), .ZN(new_n513));
  AOI21_X1  g312(.A(KEYINPUT4), .B1(new_n378), .B2(new_n501), .ZN(new_n514));
  NOR2_X1   g313(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  NAND4_X1  g314(.A1(new_n515), .A2(KEYINPUT5), .A3(new_n507), .A4(new_n500), .ZN(new_n516));
  XOR2_X1   g315(.A(G1gat), .B(G29gat), .Z(new_n517));
  XNOR2_X1  g316(.A(KEYINPUT76), .B(KEYINPUT0), .ZN(new_n518));
  XNOR2_X1  g317(.A(new_n517), .B(new_n518), .ZN(new_n519));
  XNOR2_X1  g318(.A(G57gat), .B(G85gat), .ZN(new_n520));
  XNOR2_X1  g319(.A(new_n519), .B(new_n520), .ZN(new_n521));
  INV_X1    g320(.A(new_n521), .ZN(new_n522));
  NAND4_X1  g321(.A1(new_n512), .A2(new_n516), .A3(KEYINPUT6), .A4(new_n522), .ZN(new_n523));
  NAND3_X1  g322(.A1(new_n512), .A2(new_n522), .A3(new_n516), .ZN(new_n524));
  INV_X1    g323(.A(KEYINPUT6), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  AOI21_X1  g325(.A(new_n522), .B1(new_n512), .B2(new_n516), .ZN(new_n527));
  OAI21_X1  g326(.A(new_n523), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n488), .A2(new_n528), .ZN(new_n529));
  AOI21_X1  g328(.A(new_n390), .B1(new_n389), .B2(new_n391), .ZN(new_n530));
  OAI21_X1  g329(.A(new_n407), .B1(new_n530), .B2(new_n387), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n531), .A2(new_n409), .ZN(new_n532));
  NAND3_X1  g331(.A1(new_n405), .A2(KEYINPUT79), .A3(new_n407), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  INV_X1    g333(.A(KEYINPUT81), .ZN(new_n535));
  NAND3_X1  g334(.A1(new_n534), .A2(new_n535), .A3(new_n404), .ZN(new_n536));
  NAND3_X1  g335(.A1(new_n412), .A2(new_n529), .A3(new_n536), .ZN(new_n537));
  OAI21_X1  g336(.A(new_n501), .B1(new_n436), .B2(new_n457), .ZN(new_n538));
  NAND3_X1  g337(.A1(new_n465), .A2(new_n466), .A3(new_n499), .ZN(new_n539));
  NAND4_X1  g338(.A1(new_n538), .A2(G227gat), .A3(G233gat), .A4(new_n539), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n540), .A2(KEYINPUT32), .ZN(new_n541));
  INV_X1    g340(.A(KEYINPUT33), .ZN(new_n542));
  NAND2_X1  g341(.A1(new_n540), .A2(new_n542), .ZN(new_n543));
  XOR2_X1   g342(.A(G15gat), .B(G43gat), .Z(new_n544));
  XNOR2_X1  g343(.A(G71gat), .B(G99gat), .ZN(new_n545));
  XNOR2_X1  g344(.A(new_n544), .B(new_n545), .ZN(new_n546));
  NAND3_X1  g345(.A1(new_n541), .A2(new_n543), .A3(new_n546), .ZN(new_n547));
  INV_X1    g346(.A(new_n546), .ZN(new_n548));
  OAI211_X1 g347(.A(new_n540), .B(KEYINPUT32), .C1(new_n542), .C2(new_n548), .ZN(new_n549));
  NAND2_X1  g348(.A1(new_n547), .A2(new_n549), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n538), .A2(new_n539), .ZN(new_n551));
  INV_X1    g350(.A(KEYINPUT34), .ZN(new_n552));
  NAND2_X1  g351(.A1(G227gat), .A2(G233gat), .ZN(new_n553));
  NAND3_X1  g352(.A1(new_n551), .A2(new_n552), .A3(new_n553), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n554), .A2(KEYINPUT69), .ZN(new_n555));
  AOI21_X1  g354(.A(new_n552), .B1(new_n551), .B2(new_n553), .ZN(new_n556));
  INV_X1    g355(.A(new_n556), .ZN(new_n557));
  INV_X1    g356(.A(KEYINPUT69), .ZN(new_n558));
  NAND4_X1  g357(.A1(new_n551), .A2(new_n558), .A3(new_n552), .A4(new_n553), .ZN(new_n559));
  NAND3_X1  g358(.A1(new_n555), .A2(new_n557), .A3(new_n559), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n550), .A2(new_n560), .ZN(new_n561));
  AOI21_X1  g360(.A(new_n556), .B1(KEYINPUT69), .B2(new_n554), .ZN(new_n562));
  NAND4_X1  g361(.A1(new_n562), .A2(new_n547), .A3(new_n549), .A4(new_n559), .ZN(new_n563));
  AND2_X1   g362(.A1(new_n561), .A2(new_n563), .ZN(new_n564));
  XNOR2_X1  g363(.A(KEYINPUT70), .B(KEYINPUT36), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n561), .A2(new_n563), .ZN(new_n567));
  NAND2_X1  g366(.A1(KEYINPUT70), .A2(KEYINPUT36), .ZN(new_n568));
  NAND2_X1  g367(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n566), .A2(new_n569), .ZN(new_n570));
  NAND2_X1  g369(.A1(new_n537), .A2(new_n570), .ZN(new_n571));
  INV_X1    g370(.A(KEYINPUT82), .ZN(new_n572));
  NAND2_X1  g371(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  NAND3_X1  g372(.A1(new_n537), .A2(KEYINPUT82), .A3(new_n570), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n483), .A2(KEYINPUT37), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n484), .A2(new_n575), .ZN(new_n576));
  NAND3_X1  g375(.A1(new_n474), .A2(KEYINPUT37), .A3(new_n475), .ZN(new_n577));
  NAND2_X1  g376(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n578), .A2(KEYINPUT38), .ZN(new_n579));
  NAND2_X1  g378(.A1(new_n523), .A2(KEYINPUT85), .ZN(new_n580));
  INV_X1    g379(.A(new_n580), .ZN(new_n581));
  INV_X1    g380(.A(KEYINPUT85), .ZN(new_n582));
  AOI21_X1  g381(.A(new_n581), .B1(new_n528), .B2(new_n582), .ZN(new_n583));
  INV_X1    g382(.A(KEYINPUT37), .ZN(new_n584));
  AOI21_X1  g383(.A(new_n472), .B1(new_n470), .B2(new_n471), .ZN(new_n585));
  INV_X1    g384(.A(KEYINPUT84), .ZN(new_n586));
  AOI21_X1  g385(.A(new_n584), .B1(new_n585), .B2(new_n586), .ZN(new_n587));
  NAND3_X1  g386(.A1(new_n468), .A2(KEYINPUT84), .A3(new_n473), .ZN(new_n588));
  AOI21_X1  g387(.A(KEYINPUT38), .B1(new_n587), .B2(new_n588), .ZN(new_n589));
  AOI22_X1  g388(.A1(new_n576), .A2(new_n589), .B1(new_n476), .B2(new_n481), .ZN(new_n590));
  NAND3_X1  g389(.A1(new_n579), .A2(new_n583), .A3(new_n590), .ZN(new_n591));
  INV_X1    g390(.A(KEYINPUT40), .ZN(new_n592));
  XNOR2_X1  g391(.A(KEYINPUT83), .B(KEYINPUT39), .ZN(new_n593));
  NAND3_X1  g392(.A1(new_n506), .A2(new_n508), .A3(new_n593), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n594), .A2(new_n521), .ZN(new_n595));
  NAND3_X1  g394(.A1(new_n510), .A2(new_n507), .A3(new_n502), .ZN(new_n596));
  NAND2_X1  g395(.A1(new_n596), .A2(KEYINPUT39), .ZN(new_n597));
  AOI21_X1  g396(.A(new_n597), .B1(new_n508), .B2(new_n506), .ZN(new_n598));
  OAI21_X1  g397(.A(new_n592), .B1(new_n595), .B2(new_n598), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n599), .A2(new_n524), .ZN(new_n600));
  NOR3_X1   g399(.A1(new_n595), .A2(new_n598), .A3(new_n592), .ZN(new_n601));
  NOR2_X1   g400(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  NAND3_X1  g401(.A1(new_n485), .A2(new_n487), .A3(new_n602), .ZN(new_n603));
  NAND3_X1  g402(.A1(new_n591), .A2(new_n411), .A3(new_n603), .ZN(new_n604));
  NAND3_X1  g403(.A1(new_n573), .A2(new_n574), .A3(new_n604), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n528), .A2(new_n582), .ZN(new_n606));
  AOI21_X1  g405(.A(KEYINPUT35), .B1(new_n606), .B2(new_n580), .ZN(new_n607));
  NAND4_X1  g406(.A1(new_n411), .A2(new_n607), .A3(new_n564), .A4(new_n488), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n608), .A2(KEYINPUT86), .ZN(new_n609));
  NAND2_X1  g408(.A1(new_n411), .A2(new_n564), .ZN(new_n610));
  OAI21_X1  g409(.A(KEYINPUT35), .B1(new_n610), .B2(new_n529), .ZN(new_n611));
  AOI21_X1  g410(.A(new_n567), .B1(new_n534), .B2(new_n404), .ZN(new_n612));
  INV_X1    g411(.A(KEYINPUT86), .ZN(new_n613));
  NAND4_X1  g412(.A1(new_n612), .A2(new_n613), .A3(new_n488), .A4(new_n607), .ZN(new_n614));
  AND3_X1   g413(.A1(new_n609), .A2(new_n611), .A3(new_n614), .ZN(new_n615));
  INV_X1    g414(.A(new_n615), .ZN(new_n616));
  AOI21_X1  g415(.A(new_n329), .B1(new_n605), .B2(new_n616), .ZN(new_n617));
  OR2_X1    g416(.A1(new_n528), .A2(KEYINPUT100), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n528), .A2(KEYINPUT100), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  INV_X1    g419(.A(new_n620), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n617), .A2(new_n621), .ZN(new_n622));
  XNOR2_X1  g421(.A(KEYINPUT101), .B(G1gat), .ZN(new_n623));
  XNOR2_X1  g422(.A(new_n622), .B(new_n623), .ZN(G1324gat));
  INV_X1    g423(.A(KEYINPUT42), .ZN(new_n625));
  INV_X1    g424(.A(new_n488), .ZN(new_n626));
  NAND2_X1  g425(.A1(new_n617), .A2(new_n626), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n627), .A2(G8gat), .ZN(new_n628));
  XOR2_X1   g427(.A(KEYINPUT16), .B(G8gat), .Z(new_n629));
  NAND3_X1  g428(.A1(new_n617), .A2(new_n626), .A3(new_n629), .ZN(new_n630));
  AOI21_X1  g429(.A(new_n625), .B1(new_n628), .B2(new_n630), .ZN(new_n631));
  AOI21_X1  g430(.A(new_n631), .B1(new_n625), .B2(new_n630), .ZN(new_n632));
  XNOR2_X1  g431(.A(new_n632), .B(KEYINPUT102), .ZN(G1325gat));
  INV_X1    g432(.A(G15gat), .ZN(new_n634));
  NAND3_X1  g433(.A1(new_n617), .A2(new_n634), .A3(new_n564), .ZN(new_n635));
  INV_X1    g434(.A(new_n570), .ZN(new_n636));
  AND2_X1   g435(.A1(new_n617), .A2(new_n636), .ZN(new_n637));
  OAI21_X1  g436(.A(new_n635), .B1(new_n637), .B2(new_n634), .ZN(G1326gat));
  NAND2_X1  g437(.A1(new_n412), .A2(new_n536), .ZN(new_n639));
  INV_X1    g438(.A(new_n639), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n617), .A2(new_n640), .ZN(new_n641));
  XNOR2_X1  g440(.A(new_n641), .B(KEYINPUT103), .ZN(new_n642));
  XOR2_X1   g441(.A(KEYINPUT43), .B(G22gat), .Z(new_n643));
  XNOR2_X1  g442(.A(new_n642), .B(new_n643), .ZN(G1327gat));
  AND3_X1   g443(.A1(new_n537), .A2(KEYINPUT82), .A3(new_n570), .ZN(new_n645));
  AOI21_X1  g444(.A(KEYINPUT82), .B1(new_n537), .B2(new_n570), .ZN(new_n646));
  INV_X1    g445(.A(new_n604), .ZN(new_n647));
  NOR3_X1   g446(.A1(new_n645), .A2(new_n646), .A3(new_n647), .ZN(new_n648));
  OAI21_X1  g447(.A(new_n282), .B1(new_n648), .B2(new_n615), .ZN(new_n649));
  INV_X1    g448(.A(new_n307), .ZN(new_n650));
  NOR3_X1   g449(.A1(new_n234), .A2(new_n650), .A3(new_n327), .ZN(new_n651));
  INV_X1    g450(.A(new_n651), .ZN(new_n652));
  NOR2_X1   g451(.A1(new_n649), .A2(new_n652), .ZN(new_n653));
  NAND3_X1  g452(.A1(new_n653), .A2(new_n248), .A3(new_n621), .ZN(new_n654));
  XNOR2_X1  g453(.A(new_n654), .B(KEYINPUT45), .ZN(new_n655));
  AOI21_X1  g454(.A(KEYINPUT104), .B1(new_n649), .B2(KEYINPUT44), .ZN(new_n656));
  AOI21_X1  g455(.A(new_n283), .B1(new_n605), .B2(new_n616), .ZN(new_n657));
  INV_X1    g456(.A(KEYINPUT104), .ZN(new_n658));
  INV_X1    g457(.A(KEYINPUT44), .ZN(new_n659));
  NOR3_X1   g458(.A1(new_n657), .A2(new_n658), .A3(new_n659), .ZN(new_n660));
  NAND3_X1  g459(.A1(new_n537), .A2(new_n604), .A3(new_n570), .ZN(new_n661));
  INV_X1    g460(.A(KEYINPUT105), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  NAND4_X1  g462(.A1(new_n537), .A2(new_n604), .A3(KEYINPUT105), .A4(new_n570), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  AOI21_X1  g464(.A(new_n283), .B1(new_n665), .B2(new_n616), .ZN(new_n666));
  AOI21_X1  g465(.A(KEYINPUT106), .B1(new_n666), .B2(new_n659), .ZN(new_n667));
  AOI21_X1  g466(.A(new_n615), .B1(new_n663), .B2(new_n664), .ZN(new_n668));
  INV_X1    g467(.A(KEYINPUT106), .ZN(new_n669));
  NOR4_X1   g468(.A1(new_n668), .A2(new_n669), .A3(KEYINPUT44), .A4(new_n283), .ZN(new_n670));
  OAI22_X1  g469(.A1(new_n656), .A2(new_n660), .B1(new_n667), .B2(new_n670), .ZN(new_n671));
  INV_X1    g470(.A(new_n671), .ZN(new_n672));
  NOR3_X1   g471(.A1(new_n672), .A2(new_n620), .A3(new_n652), .ZN(new_n673));
  OAI21_X1  g472(.A(new_n655), .B1(new_n673), .B2(new_n248), .ZN(G1328gat));
  INV_X1    g473(.A(G36gat), .ZN(new_n675));
  NAND3_X1  g474(.A1(new_n653), .A2(new_n675), .A3(new_n626), .ZN(new_n676));
  XOR2_X1   g475(.A(new_n676), .B(KEYINPUT46), .Z(new_n677));
  NOR3_X1   g476(.A1(new_n672), .A2(new_n488), .A3(new_n652), .ZN(new_n678));
  OAI21_X1  g477(.A(new_n677), .B1(new_n678), .B2(new_n675), .ZN(G1329gat));
  NAND4_X1  g478(.A1(new_n671), .A2(G43gat), .A3(new_n636), .A4(new_n651), .ZN(new_n680));
  AOI21_X1  g479(.A(G43gat), .B1(new_n653), .B2(new_n564), .ZN(new_n681));
  INV_X1    g480(.A(new_n681), .ZN(new_n682));
  NAND2_X1  g481(.A1(new_n680), .A2(new_n682), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n683), .A2(KEYINPUT47), .ZN(new_n684));
  INV_X1    g483(.A(KEYINPUT47), .ZN(new_n685));
  NAND3_X1  g484(.A1(new_n680), .A2(new_n685), .A3(new_n682), .ZN(new_n686));
  NAND2_X1  g485(.A1(new_n684), .A2(new_n686), .ZN(G1330gat));
  INV_X1    g486(.A(G50gat), .ZN(new_n688));
  NAND3_X1  g487(.A1(new_n653), .A2(new_n688), .A3(new_n640), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n665), .A2(new_n616), .ZN(new_n690));
  NAND3_X1  g489(.A1(new_n690), .A2(new_n659), .A3(new_n282), .ZN(new_n691));
  NAND2_X1  g490(.A1(new_n691), .A2(new_n669), .ZN(new_n692));
  NAND3_X1  g491(.A1(new_n666), .A2(KEYINPUT106), .A3(new_n659), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  NAND3_X1  g493(.A1(new_n649), .A2(KEYINPUT104), .A3(KEYINPUT44), .ZN(new_n695));
  OAI21_X1  g494(.A(new_n658), .B1(new_n657), .B2(new_n659), .ZN(new_n696));
  NAND2_X1  g495(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  AOI211_X1 g496(.A(new_n411), .B(new_n652), .C1(new_n694), .C2(new_n697), .ZN(new_n698));
  OAI211_X1 g497(.A(KEYINPUT48), .B(new_n689), .C1(new_n698), .C2(new_n688), .ZN(new_n699));
  NAND3_X1  g498(.A1(new_n671), .A2(new_n640), .A3(new_n651), .ZN(new_n700));
  INV_X1    g499(.A(KEYINPUT107), .ZN(new_n701));
  NAND3_X1  g500(.A1(new_n700), .A2(new_n701), .A3(G50gat), .ZN(new_n702));
  INV_X1    g501(.A(KEYINPUT48), .ZN(new_n703));
  NAND2_X1  g502(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n689), .A2(KEYINPUT107), .ZN(new_n705));
  AOI21_X1  g504(.A(new_n705), .B1(new_n700), .B2(G50gat), .ZN(new_n706));
  OAI21_X1  g505(.A(new_n699), .B1(new_n704), .B2(new_n706), .ZN(G1331gat));
  NAND2_X1  g506(.A1(new_n234), .A2(new_n283), .ZN(new_n708));
  NOR4_X1   g507(.A1(new_n668), .A2(new_n307), .A3(new_n708), .A4(new_n328), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n709), .A2(new_n621), .ZN(new_n710));
  XNOR2_X1  g509(.A(new_n710), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g510(.A1(new_n709), .A2(new_n626), .ZN(new_n712));
  OAI21_X1  g511(.A(new_n712), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n713));
  XOR2_X1   g512(.A(KEYINPUT49), .B(G64gat), .Z(new_n714));
  OAI21_X1  g513(.A(new_n713), .B1(new_n712), .B2(new_n714), .ZN(G1333gat));
  INV_X1    g514(.A(G71gat), .ZN(new_n716));
  NAND3_X1  g515(.A1(new_n709), .A2(new_n716), .A3(new_n564), .ZN(new_n717));
  AND2_X1   g516(.A1(new_n709), .A2(new_n636), .ZN(new_n718));
  OAI21_X1  g517(.A(new_n717), .B1(new_n718), .B2(new_n716), .ZN(new_n719));
  XNOR2_X1  g518(.A(KEYINPUT108), .B(KEYINPUT50), .ZN(new_n720));
  XNOR2_X1  g519(.A(new_n719), .B(new_n720), .ZN(G1334gat));
  NAND2_X1  g520(.A1(new_n709), .A2(new_n640), .ZN(new_n722));
  XNOR2_X1  g521(.A(new_n722), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g522(.A1(new_n234), .A2(new_n307), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n724), .A2(new_n327), .ZN(new_n725));
  AOI21_X1  g524(.A(new_n725), .B1(new_n694), .B2(new_n697), .ZN(new_n726));
  AOI21_X1  g525(.A(new_n242), .B1(new_n726), .B2(new_n621), .ZN(new_n727));
  AOI21_X1  g526(.A(KEYINPUT51), .B1(new_n666), .B2(new_n724), .ZN(new_n728));
  INV_X1    g527(.A(new_n728), .ZN(new_n729));
  NAND3_X1  g528(.A1(new_n666), .A2(KEYINPUT51), .A3(new_n724), .ZN(new_n730));
  AOI21_X1  g529(.A(new_n328), .B1(new_n729), .B2(new_n730), .ZN(new_n731));
  NOR2_X1   g530(.A1(new_n620), .A2(G85gat), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  INV_X1    g532(.A(new_n733), .ZN(new_n734));
  OAI21_X1  g533(.A(KEYINPUT109), .B1(new_n727), .B2(new_n734), .ZN(new_n735));
  INV_X1    g534(.A(KEYINPUT109), .ZN(new_n736));
  AOI211_X1 g535(.A(new_n620), .B(new_n725), .C1(new_n694), .C2(new_n697), .ZN(new_n737));
  OAI211_X1 g536(.A(new_n736), .B(new_n733), .C1(new_n737), .C2(new_n242), .ZN(new_n738));
  NAND2_X1  g537(.A1(new_n735), .A2(new_n738), .ZN(G1336gat));
  AOI21_X1  g538(.A(new_n243), .B1(new_n726), .B2(new_n626), .ZN(new_n740));
  NOR2_X1   g539(.A1(new_n488), .A2(G92gat), .ZN(new_n741));
  NAND2_X1  g540(.A1(new_n731), .A2(new_n741), .ZN(new_n742));
  INV_X1    g541(.A(new_n742), .ZN(new_n743));
  OAI21_X1  g542(.A(KEYINPUT52), .B1(new_n740), .B2(new_n743), .ZN(new_n744));
  INV_X1    g543(.A(KEYINPUT52), .ZN(new_n745));
  AOI211_X1 g544(.A(new_n488), .B(new_n725), .C1(new_n694), .C2(new_n697), .ZN(new_n746));
  OAI211_X1 g545(.A(new_n745), .B(new_n742), .C1(new_n746), .C2(new_n243), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n744), .A2(new_n747), .ZN(G1337gat));
  XNOR2_X1  g547(.A(KEYINPUT110), .B(G99gat), .ZN(new_n749));
  INV_X1    g548(.A(new_n749), .ZN(new_n750));
  NAND3_X1  g549(.A1(new_n726), .A2(new_n636), .A3(new_n750), .ZN(new_n751));
  INV_X1    g550(.A(new_n730), .ZN(new_n752));
  OAI21_X1  g551(.A(new_n327), .B1(new_n752), .B2(new_n728), .ZN(new_n753));
  OAI21_X1  g552(.A(new_n749), .B1(new_n753), .B2(new_n567), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n751), .A2(new_n754), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n755), .A2(KEYINPUT111), .ZN(new_n756));
  INV_X1    g555(.A(KEYINPUT111), .ZN(new_n757));
  NAND3_X1  g556(.A1(new_n751), .A2(new_n757), .A3(new_n754), .ZN(new_n758));
  NAND2_X1  g557(.A1(new_n756), .A2(new_n758), .ZN(G1338gat));
  NAND2_X1  g558(.A1(new_n726), .A2(new_n640), .ZN(new_n760));
  INV_X1    g559(.A(new_n411), .ZN(new_n761));
  INV_X1    g560(.A(G106gat), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  INV_X1    g562(.A(new_n763), .ZN(new_n764));
  AOI22_X1  g563(.A1(new_n760), .A2(G106gat), .B1(new_n731), .B2(new_n764), .ZN(new_n765));
  INV_X1    g564(.A(KEYINPUT53), .ZN(new_n766));
  AOI21_X1  g565(.A(new_n762), .B1(new_n726), .B2(new_n761), .ZN(new_n767));
  OAI21_X1  g566(.A(new_n766), .B1(new_n753), .B2(new_n763), .ZN(new_n768));
  OAI22_X1  g567(.A1(new_n765), .A2(new_n766), .B1(new_n767), .B2(new_n768), .ZN(G1339gat));
  NOR2_X1   g568(.A1(new_n626), .A2(new_n620), .ZN(new_n770));
  INV_X1    g569(.A(new_n770), .ZN(new_n771));
  NOR2_X1   g570(.A1(new_n771), .A2(new_n567), .ZN(new_n772));
  INV_X1    g571(.A(new_n234), .ZN(new_n773));
  INV_X1    g572(.A(KEYINPUT112), .ZN(new_n774));
  OAI21_X1  g573(.A(new_n774), .B1(new_n313), .B2(new_n314), .ZN(new_n775));
  INV_X1    g574(.A(new_n314), .ZN(new_n776));
  NAND4_X1  g575(.A1(new_n311), .A2(new_n312), .A3(KEYINPUT112), .A4(new_n776), .ZN(new_n777));
  NAND2_X1  g576(.A1(new_n775), .A2(new_n777), .ZN(new_n778));
  NAND3_X1  g577(.A1(new_n778), .A2(KEYINPUT54), .A3(new_n315), .ZN(new_n779));
  INV_X1    g578(.A(KEYINPUT54), .ZN(new_n780));
  NAND3_X1  g579(.A1(new_n323), .A2(new_n780), .A3(new_n325), .ZN(new_n781));
  NAND3_X1  g580(.A1(new_n779), .A2(new_n319), .A3(new_n781), .ZN(new_n782));
  INV_X1    g581(.A(KEYINPUT55), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n782), .A2(new_n783), .ZN(new_n784));
  NAND4_X1  g583(.A1(new_n779), .A2(new_n781), .A3(KEYINPUT55), .A4(new_n319), .ZN(new_n785));
  NAND4_X1  g584(.A1(new_n784), .A2(new_n307), .A3(new_n322), .A4(new_n785), .ZN(new_n786));
  OAI22_X1  g585(.A1(new_n292), .A2(new_n294), .B1(new_n298), .B2(new_n299), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n787), .A2(new_n287), .ZN(new_n788));
  INV_X1    g587(.A(KEYINPUT113), .ZN(new_n789));
  XNOR2_X1  g588(.A(new_n788), .B(new_n789), .ZN(new_n790));
  NAND3_X1  g589(.A1(new_n790), .A2(new_n306), .A3(new_n327), .ZN(new_n791));
  AOI21_X1  g590(.A(new_n282), .B1(new_n786), .B2(new_n791), .ZN(new_n792));
  NAND4_X1  g591(.A1(new_n790), .A2(new_n306), .A3(new_n322), .A4(new_n785), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n282), .A2(new_n784), .ZN(new_n794));
  NOR2_X1   g593(.A1(new_n793), .A2(new_n794), .ZN(new_n795));
  OAI21_X1  g594(.A(new_n773), .B1(new_n792), .B2(new_n795), .ZN(new_n796));
  NAND4_X1  g595(.A1(new_n234), .A2(new_n283), .A3(new_n650), .A4(new_n328), .ZN(new_n797));
  AND3_X1   g596(.A1(new_n796), .A2(KEYINPUT114), .A3(new_n797), .ZN(new_n798));
  AOI21_X1  g597(.A(KEYINPUT114), .B1(new_n796), .B2(new_n797), .ZN(new_n799));
  OAI211_X1 g598(.A(new_n639), .B(new_n772), .C1(new_n798), .C2(new_n799), .ZN(new_n800));
  OAI21_X1  g599(.A(G113gat), .B1(new_n800), .B2(new_n650), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n796), .A2(new_n797), .ZN(new_n802));
  INV_X1    g601(.A(KEYINPUT114), .ZN(new_n803));
  NAND2_X1  g602(.A1(new_n802), .A2(new_n803), .ZN(new_n804));
  NAND3_X1  g603(.A1(new_n796), .A2(KEYINPUT114), .A3(new_n797), .ZN(new_n805));
  AOI21_X1  g604(.A(new_n620), .B1(new_n804), .B2(new_n805), .ZN(new_n806));
  NOR2_X1   g605(.A1(new_n610), .A2(new_n626), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n806), .A2(new_n807), .ZN(new_n808));
  NOR2_X1   g607(.A1(new_n650), .A2(G113gat), .ZN(new_n809));
  XNOR2_X1  g608(.A(new_n809), .B(KEYINPUT115), .ZN(new_n810));
  OAI21_X1  g609(.A(new_n801), .B1(new_n808), .B2(new_n810), .ZN(G1340gat));
  INV_X1    g610(.A(G120gat), .ZN(new_n812));
  NOR3_X1   g611(.A1(new_n800), .A2(new_n812), .A3(new_n328), .ZN(new_n813));
  NAND3_X1  g612(.A1(new_n806), .A2(new_n807), .A3(new_n327), .ZN(new_n814));
  AOI21_X1  g613(.A(new_n813), .B1(new_n812), .B2(new_n814), .ZN(G1341gat));
  INV_X1    g614(.A(KEYINPUT116), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n234), .A2(G127gat), .ZN(new_n817));
  OR3_X1    g616(.A1(new_n800), .A2(new_n816), .A3(new_n817), .ZN(new_n818));
  OAI21_X1  g617(.A(new_n816), .B1(new_n800), .B2(new_n817), .ZN(new_n819));
  NOR2_X1   g618(.A1(new_n808), .A2(new_n773), .ZN(new_n820));
  OAI211_X1 g619(.A(new_n818), .B(new_n819), .C1(new_n820), .C2(G127gat), .ZN(new_n821));
  XNOR2_X1  g620(.A(new_n821), .B(KEYINPUT117), .ZN(G1342gat));
  OAI21_X1  g621(.A(G134gat), .B1(new_n800), .B2(new_n283), .ZN(new_n823));
  AND2_X1   g622(.A1(new_n823), .A2(KEYINPUT118), .ZN(new_n824));
  INV_X1    g623(.A(KEYINPUT118), .ZN(new_n825));
  OAI211_X1 g624(.A(new_n825), .B(G134gat), .C1(new_n800), .C2(new_n283), .ZN(new_n826));
  INV_X1    g625(.A(new_n826), .ZN(new_n827));
  NOR2_X1   g626(.A1(new_n824), .A2(new_n827), .ZN(new_n828));
  NOR2_X1   g627(.A1(new_n283), .A2(G134gat), .ZN(new_n829));
  INV_X1    g628(.A(new_n829), .ZN(new_n830));
  OAI21_X1  g629(.A(KEYINPUT56), .B1(new_n808), .B2(new_n830), .ZN(new_n831));
  INV_X1    g630(.A(KEYINPUT56), .ZN(new_n832));
  NAND4_X1  g631(.A1(new_n806), .A2(new_n832), .A3(new_n807), .A4(new_n829), .ZN(new_n833));
  NAND2_X1  g632(.A1(new_n831), .A2(new_n833), .ZN(new_n834));
  OAI21_X1  g633(.A(KEYINPUT119), .B1(new_n828), .B2(new_n834), .ZN(new_n835));
  AND2_X1   g634(.A1(new_n831), .A2(new_n833), .ZN(new_n836));
  INV_X1    g635(.A(KEYINPUT119), .ZN(new_n837));
  OAI211_X1 g636(.A(new_n836), .B(new_n837), .C1(new_n824), .C2(new_n827), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n835), .A2(new_n838), .ZN(G1343gat));
  INV_X1    g638(.A(KEYINPUT58), .ZN(new_n840));
  NOR3_X1   g639(.A1(new_n636), .A2(new_n411), .A3(new_n626), .ZN(new_n841));
  NAND2_X1  g640(.A1(new_n806), .A2(new_n841), .ZN(new_n842));
  INV_X1    g641(.A(new_n842), .ZN(new_n843));
  INV_X1    g642(.A(G141gat), .ZN(new_n844));
  NAND3_X1  g643(.A1(new_n843), .A2(new_n844), .A3(new_n307), .ZN(new_n845));
  AOI21_X1  g644(.A(new_n840), .B1(new_n845), .B2(KEYINPUT122), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n570), .A2(new_n770), .ZN(new_n847));
  XOR2_X1   g646(.A(new_n847), .B(KEYINPUT120), .Z(new_n848));
  INV_X1    g647(.A(KEYINPUT121), .ZN(new_n849));
  OR2_X1    g648(.A1(new_n796), .A2(new_n849), .ZN(new_n850));
  INV_X1    g649(.A(new_n797), .ZN(new_n851));
  AOI21_X1  g650(.A(new_n851), .B1(new_n796), .B2(new_n849), .ZN(new_n852));
  AOI21_X1  g651(.A(new_n639), .B1(new_n850), .B2(new_n852), .ZN(new_n853));
  INV_X1    g652(.A(KEYINPUT57), .ZN(new_n854));
  OAI21_X1  g653(.A(new_n848), .B1(new_n853), .B2(new_n854), .ZN(new_n855));
  AOI211_X1 g654(.A(KEYINPUT57), .B(new_n411), .C1(new_n804), .C2(new_n805), .ZN(new_n856));
  NOR2_X1   g655(.A1(new_n855), .A2(new_n856), .ZN(new_n857));
  AOI21_X1  g656(.A(new_n844), .B1(new_n857), .B2(new_n307), .ZN(new_n858));
  INV_X1    g657(.A(new_n845), .ZN(new_n859));
  OAI21_X1  g658(.A(new_n846), .B1(new_n858), .B2(new_n859), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n804), .A2(new_n805), .ZN(new_n861));
  NAND3_X1  g660(.A1(new_n861), .A2(new_n854), .A3(new_n761), .ZN(new_n862));
  OAI211_X1 g661(.A(new_n862), .B(new_n848), .C1(new_n854), .C2(new_n853), .ZN(new_n863));
  OAI21_X1  g662(.A(G141gat), .B1(new_n863), .B2(new_n650), .ZN(new_n864));
  OAI211_X1 g663(.A(new_n864), .B(new_n845), .C1(KEYINPUT122), .C2(new_n840), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n860), .A2(new_n865), .ZN(G1344gat));
  INV_X1    g665(.A(KEYINPUT59), .ZN(new_n867));
  AOI211_X1 g666(.A(new_n867), .B(G148gat), .C1(new_n843), .C2(new_n327), .ZN(new_n868));
  OAI21_X1  g667(.A(new_n867), .B1(new_n863), .B2(new_n328), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n861), .A2(new_n761), .ZN(new_n870));
  NAND2_X1  g669(.A1(new_n870), .A2(KEYINPUT57), .ZN(new_n871));
  NAND3_X1  g670(.A1(new_n802), .A2(new_n854), .A3(new_n640), .ZN(new_n872));
  NAND2_X1  g671(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  NAND3_X1  g672(.A1(new_n848), .A2(KEYINPUT59), .A3(new_n327), .ZN(new_n874));
  OAI21_X1  g673(.A(new_n869), .B1(new_n873), .B2(new_n874), .ZN(new_n875));
  AOI21_X1  g674(.A(new_n868), .B1(new_n875), .B2(G148gat), .ZN(G1345gat));
  OAI21_X1  g675(.A(G155gat), .B1(new_n863), .B2(new_n773), .ZN(new_n877));
  NAND3_X1  g676(.A1(new_n843), .A2(new_n340), .A3(new_n234), .ZN(new_n878));
  NAND2_X1  g677(.A1(new_n877), .A2(new_n878), .ZN(G1346gat));
  OR3_X1    g678(.A1(new_n842), .A2(new_n344), .A3(new_n283), .ZN(new_n880));
  INV_X1    g679(.A(KEYINPUT123), .ZN(new_n881));
  NAND3_X1  g680(.A1(new_n857), .A2(new_n881), .A3(new_n282), .ZN(new_n882));
  NAND2_X1  g681(.A1(new_n882), .A2(new_n344), .ZN(new_n883));
  AOI21_X1  g682(.A(new_n881), .B1(new_n857), .B2(new_n282), .ZN(new_n884));
  OAI21_X1  g683(.A(new_n880), .B1(new_n883), .B2(new_n884), .ZN(G1347gat));
  NAND3_X1  g684(.A1(new_n626), .A2(new_n620), .A3(new_n564), .ZN(new_n886));
  XOR2_X1   g685(.A(new_n886), .B(KEYINPUT124), .Z(new_n887));
  OAI211_X1 g686(.A(new_n639), .B(new_n887), .C1(new_n798), .C2(new_n799), .ZN(new_n888));
  INV_X1    g687(.A(G169gat), .ZN(new_n889));
  NOR3_X1   g688(.A1(new_n888), .A2(new_n889), .A3(new_n650), .ZN(new_n890));
  AOI21_X1  g689(.A(new_n621), .B1(new_n804), .B2(new_n805), .ZN(new_n891));
  NOR2_X1   g690(.A1(new_n610), .A2(new_n488), .ZN(new_n892));
  NAND2_X1  g691(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  INV_X1    g692(.A(new_n893), .ZN(new_n894));
  NAND2_X1  g693(.A1(new_n894), .A2(new_n307), .ZN(new_n895));
  AOI21_X1  g694(.A(new_n890), .B1(new_n895), .B2(new_n889), .ZN(G1348gat));
  OAI21_X1  g695(.A(G176gat), .B1(new_n888), .B2(new_n328), .ZN(new_n897));
  OR2_X1    g696(.A1(new_n328), .A2(G176gat), .ZN(new_n898));
  OAI21_X1  g697(.A(new_n897), .B1(new_n893), .B2(new_n898), .ZN(G1349gat));
  OAI21_X1  g698(.A(new_n425), .B1(new_n888), .B2(new_n773), .ZN(new_n900));
  NAND3_X1  g699(.A1(new_n234), .A2(new_n423), .A3(new_n428), .ZN(new_n901));
  OAI21_X1  g700(.A(new_n900), .B1(new_n893), .B2(new_n901), .ZN(new_n902));
  XNOR2_X1  g701(.A(new_n902), .B(KEYINPUT60), .ZN(G1350gat));
  INV_X1    g702(.A(KEYINPUT126), .ZN(new_n904));
  OAI21_X1  g703(.A(G190gat), .B1(new_n888), .B2(new_n283), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n905), .A2(KEYINPUT125), .ZN(new_n906));
  INV_X1    g705(.A(KEYINPUT125), .ZN(new_n907));
  OAI211_X1 g706(.A(new_n907), .B(G190gat), .C1(new_n888), .C2(new_n283), .ZN(new_n908));
  AND3_X1   g707(.A1(new_n906), .A2(KEYINPUT61), .A3(new_n908), .ZN(new_n909));
  NAND3_X1  g708(.A1(new_n894), .A2(new_n429), .A3(new_n282), .ZN(new_n910));
  INV_X1    g709(.A(KEYINPUT61), .ZN(new_n911));
  NAND3_X1  g710(.A1(new_n905), .A2(KEYINPUT125), .A3(new_n911), .ZN(new_n912));
  NAND2_X1  g711(.A1(new_n910), .A2(new_n912), .ZN(new_n913));
  OAI21_X1  g712(.A(new_n904), .B1(new_n909), .B2(new_n913), .ZN(new_n914));
  NAND3_X1  g713(.A1(new_n906), .A2(KEYINPUT61), .A3(new_n908), .ZN(new_n915));
  NAND4_X1  g714(.A1(new_n915), .A2(KEYINPUT126), .A3(new_n912), .A4(new_n910), .ZN(new_n916));
  NAND2_X1  g715(.A1(new_n914), .A2(new_n916), .ZN(G1351gat));
  NOR3_X1   g716(.A1(new_n636), .A2(new_n488), .A3(new_n621), .ZN(new_n918));
  NAND3_X1  g717(.A1(new_n871), .A2(new_n872), .A3(new_n918), .ZN(new_n919));
  INV_X1    g718(.A(G197gat), .ZN(new_n920));
  NOR3_X1   g719(.A1(new_n919), .A2(new_n920), .A3(new_n650), .ZN(new_n921));
  NOR3_X1   g720(.A1(new_n636), .A2(new_n411), .A3(new_n488), .ZN(new_n922));
  NAND2_X1  g721(.A1(new_n891), .A2(new_n922), .ZN(new_n923));
  INV_X1    g722(.A(new_n923), .ZN(new_n924));
  AOI21_X1  g723(.A(G197gat), .B1(new_n924), .B2(new_n307), .ZN(new_n925));
  NOR2_X1   g724(.A1(new_n921), .A2(new_n925), .ZN(G1352gat));
  OAI21_X1  g725(.A(G204gat), .B1(new_n919), .B2(new_n328), .ZN(new_n927));
  INV_X1    g726(.A(G204gat), .ZN(new_n928));
  NAND2_X1  g727(.A1(KEYINPUT127), .A2(KEYINPUT62), .ZN(new_n929));
  NAND4_X1  g728(.A1(new_n924), .A2(new_n928), .A3(new_n327), .A4(new_n929), .ZN(new_n930));
  XNOR2_X1  g729(.A(KEYINPUT127), .B(KEYINPUT62), .ZN(new_n931));
  NAND2_X1  g730(.A1(new_n327), .A2(new_n928), .ZN(new_n932));
  OAI21_X1  g731(.A(new_n931), .B1(new_n923), .B2(new_n932), .ZN(new_n933));
  NAND3_X1  g732(.A1(new_n927), .A2(new_n930), .A3(new_n933), .ZN(G1353gat));
  OR3_X1    g733(.A1(new_n923), .A2(G211gat), .A3(new_n773), .ZN(new_n935));
  NAND4_X1  g734(.A1(new_n871), .A2(new_n234), .A3(new_n872), .A4(new_n918), .ZN(new_n936));
  AND3_X1   g735(.A1(new_n936), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n937));
  AOI21_X1  g736(.A(KEYINPUT63), .B1(new_n936), .B2(G211gat), .ZN(new_n938));
  OAI21_X1  g737(.A(new_n935), .B1(new_n937), .B2(new_n938), .ZN(G1354gat));
  OAI21_X1  g738(.A(G218gat), .B1(new_n919), .B2(new_n283), .ZN(new_n940));
  OR3_X1    g739(.A1(new_n923), .A2(G218gat), .A3(new_n283), .ZN(new_n941));
  NAND2_X1  g740(.A1(new_n940), .A2(new_n941), .ZN(G1355gat));
endmodule


