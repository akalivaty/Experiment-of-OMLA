

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599,
         n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610,
         n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621,
         n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632,
         n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643,
         n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654,
         n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665,
         n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676,
         n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687,
         n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698,
         n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709,
         n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720,
         n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731,
         n732, n733, n734, n735, n736, n737, n738, n739, n740, n741, n742,
         n743, n744, n745, n746, n747, n748, n749, n750, n751, n752, n753,
         n754, n755, n756, n757, n758, n759, n760, n761, n762, n763, n764,
         n765, n766, n767, n768, n769, n770, n771, n772, n773, n774, n775,
         n776, n777, n778, n779, n780, n781, n782, n783, n784, n785, n786,
         n787, n788, n789, n790, n791, n792, n793, n794, n795, n796, n797,
         n798, n799, n800, n801, n802, n803, n804, n805, n806, n807, n808,
         n809, n810, n811, n812, n813, n814, n815, n816, n817, n818, n819,
         n820, n821, n822, n823, n824, n825, n826, n827, n828, n829, n830,
         n831, n832, n833, n834, n835, n836, n837, n838, n839, n840, n841,
         n842, n843, n844, n845, n846, n847, n848, n849, n850, n851, n852,
         n853, n854, n855, n856, n857, n858, n859, n860, n861, n862, n863,
         n864, n865, n866, n867, n868, n869, n870, n871, n872, n873, n874,
         n875, n876, n877, n878, n879, n880, n881, n882, n883, n884, n885,
         n886, n887, n888, n889, n890, n891, n892, n893, n894, n895, n896,
         n897, n898, n899, n900, n901, n902, n903, n904, n905, n906, n907,
         n908, n909, n910, n911, n912, n913, n914, n915, n916, n917, n918,
         n919, n920, n921, n922, n923, n924, n925, n926, n927, n928, n929,
         n930, n931, n932, n933, n934, n935, n936, n937, n938, n939, n940,
         n941, n942, n943, n944, n945, n946, n947, n948, n949, n950, n951,
         n952, n953, n954, n955, n956, n957, n958, n959, n960, n961, n962,
         n963, n964, n965, n966, n967, n968, n969, n970, n971, n972, n973,
         n974, n975, n976, n977, n978, n979, n980, n981, n982, n983, n984,
         n985, n986, n987, n988, n989, n990, n991, n992, n993, n994, n995,
         n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005,
         n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015,
         n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025,
         n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035,
         n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045,
         n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055,
         n1056;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NOR2_X1 U563 ( .A1(G651), .A2(n677), .ZN(n681) );
  NAND2_X1 U564 ( .A1(n775), .A2(G8), .ZN(n776) );
  NOR2_X4 U565 ( .A1(n570), .A2(n569), .ZN(G160) );
  XNOR2_X1 U566 ( .A(KEYINPUT71), .B(n614), .ZN(n970) );
  NOR2_X1 U567 ( .A1(n719), .A2(G1384), .ZN(n734) );
  BUF_X2 U568 ( .A(n564), .Z(n530) );
  NOR2_X1 U569 ( .A1(G2105), .A2(n537), .ZN(n560) );
  INV_X2 U570 ( .A(n770), .ZN(n775) );
  OR2_X1 U571 ( .A1(n814), .A2(n813), .ZN(n824) );
  INV_X1 U572 ( .A(G2104), .ZN(n537) );
  NOR2_X1 U573 ( .A1(n740), .A2(n970), .ZN(n742) );
  AND2_X1 U574 ( .A1(n767), .A2(n766), .ZN(n768) );
  INV_X1 U575 ( .A(KEYINPUT110), .ZN(n827) );
  NAND2_X1 U576 ( .A1(n831), .A2(n804), .ZN(n531) );
  NOR2_X1 U577 ( .A1(n807), .A2(n819), .ZN(n532) );
  OR2_X1 U578 ( .A1(n814), .A2(n800), .ZN(n533) );
  INV_X1 U579 ( .A(KEYINPUT65), .ZN(n741) );
  XNOR2_X1 U580 ( .A(n742), .B(n741), .ZN(n757) );
  NOR2_X1 U581 ( .A1(n757), .A2(n960), .ZN(n758) );
  NAND2_X1 U582 ( .A1(n734), .A2(n733), .ZN(n736) );
  INV_X1 U583 ( .A(KEYINPUT32), .ZN(n793) );
  NOR2_X1 U584 ( .A1(G2104), .A2(G2105), .ZN(n534) );
  AND2_X2 U585 ( .A1(n537), .A2(G2105), .ZN(n912) );
  NOR2_X1 U586 ( .A1(n544), .A2(n543), .ZN(n719) );
  BUF_X1 U587 ( .A(n719), .Z(G164) );
  XOR2_X1 U588 ( .A(KEYINPUT17), .B(n534), .Z(n564) );
  NAND2_X1 U589 ( .A1(G138), .A2(n530), .ZN(n536) );
  BUF_X1 U590 ( .A(n560), .Z(n909) );
  NAND2_X1 U591 ( .A1(G102), .A2(n909), .ZN(n535) );
  NAND2_X1 U592 ( .A1(n536), .A2(n535), .ZN(n544) );
  INV_X1 U593 ( .A(KEYINPUT91), .ZN(n542) );
  NAND2_X1 U594 ( .A1(n912), .A2(G126), .ZN(n538) );
  XNOR2_X1 U595 ( .A(n538), .B(KEYINPUT90), .ZN(n540) );
  AND2_X1 U596 ( .A1(G2104), .A2(G2105), .ZN(n913) );
  NAND2_X1 U597 ( .A1(G114), .A2(n913), .ZN(n539) );
  NAND2_X1 U598 ( .A1(n540), .A2(n539), .ZN(n541) );
  XNOR2_X1 U599 ( .A(n542), .B(n541), .ZN(n543) );
  XOR2_X1 U600 ( .A(G543), .B(KEYINPUT0), .Z(n677) );
  NAND2_X1 U601 ( .A1(G51), .A2(n681), .ZN(n548) );
  INV_X1 U602 ( .A(G651), .ZN(n551) );
  NOR2_X1 U603 ( .A1(G543), .A2(n551), .ZN(n546) );
  XNOR2_X1 U604 ( .A(KEYINPUT67), .B(KEYINPUT1), .ZN(n545) );
  XNOR2_X1 U605 ( .A(n546), .B(n545), .ZN(n689) );
  NAND2_X1 U606 ( .A1(G63), .A2(n689), .ZN(n547) );
  NAND2_X1 U607 ( .A1(n548), .A2(n547), .ZN(n549) );
  XNOR2_X1 U608 ( .A(KEYINPUT6), .B(n549), .ZN(n557) );
  NOR2_X1 U609 ( .A1(G651), .A2(G543), .ZN(n680) );
  NAND2_X1 U610 ( .A1(n680), .A2(G89), .ZN(n550) );
  XNOR2_X1 U611 ( .A(n550), .B(KEYINPUT4), .ZN(n553) );
  NOR2_X2 U612 ( .A1(n677), .A2(n551), .ZN(n684) );
  NAND2_X1 U613 ( .A1(G76), .A2(n684), .ZN(n552) );
  NAND2_X1 U614 ( .A1(n553), .A2(n552), .ZN(n554) );
  XOR2_X1 U615 ( .A(KEYINPUT5), .B(n554), .Z(n555) );
  XNOR2_X1 U616 ( .A(KEYINPUT78), .B(n555), .ZN(n556) );
  NOR2_X1 U617 ( .A1(n557), .A2(n556), .ZN(n559) );
  XNOR2_X1 U618 ( .A(KEYINPUT79), .B(KEYINPUT7), .ZN(n558) );
  XNOR2_X1 U619 ( .A(n559), .B(n558), .ZN(G168) );
  XOR2_X1 U620 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U621 ( .A1(G101), .A2(n560), .ZN(n561) );
  XNOR2_X1 U622 ( .A(n561), .B(KEYINPUT23), .ZN(n563) );
  INV_X1 U623 ( .A(KEYINPUT66), .ZN(n562) );
  XNOR2_X1 U624 ( .A(n563), .B(n562), .ZN(n566) );
  NAND2_X1 U625 ( .A1(G137), .A2(n530), .ZN(n565) );
  NAND2_X1 U626 ( .A1(n566), .A2(n565), .ZN(n570) );
  NAND2_X1 U627 ( .A1(G125), .A2(n912), .ZN(n568) );
  NAND2_X1 U628 ( .A1(G113), .A2(n913), .ZN(n567) );
  NAND2_X1 U629 ( .A1(n568), .A2(n567), .ZN(n569) );
  NAND2_X1 U630 ( .A1(G91), .A2(n680), .ZN(n572) );
  NAND2_X1 U631 ( .A1(G78), .A2(n684), .ZN(n571) );
  NAND2_X1 U632 ( .A1(n572), .A2(n571), .ZN(n575) );
  NAND2_X1 U633 ( .A1(n689), .A2(G65), .ZN(n573) );
  XOR2_X1 U634 ( .A(KEYINPUT68), .B(n573), .Z(n574) );
  NOR2_X1 U635 ( .A1(n575), .A2(n574), .ZN(n577) );
  NAND2_X1 U636 ( .A1(n681), .A2(G53), .ZN(n576) );
  NAND2_X1 U637 ( .A1(n577), .A2(n576), .ZN(G299) );
  NAND2_X1 U638 ( .A1(G85), .A2(n680), .ZN(n579) );
  NAND2_X1 U639 ( .A1(G72), .A2(n684), .ZN(n578) );
  NAND2_X1 U640 ( .A1(n579), .A2(n578), .ZN(n583) );
  NAND2_X1 U641 ( .A1(G47), .A2(n681), .ZN(n581) );
  NAND2_X1 U642 ( .A1(G60), .A2(n689), .ZN(n580) );
  NAND2_X1 U643 ( .A1(n581), .A2(n580), .ZN(n582) );
  OR2_X1 U644 ( .A1(n583), .A2(n582), .ZN(G290) );
  XOR2_X1 U645 ( .A(G2443), .B(G2446), .Z(n585) );
  XNOR2_X1 U646 ( .A(G2427), .B(G2451), .ZN(n584) );
  XNOR2_X1 U647 ( .A(n585), .B(n584), .ZN(n591) );
  XOR2_X1 U648 ( .A(G2430), .B(G2454), .Z(n587) );
  XNOR2_X1 U649 ( .A(G1348), .B(G1341), .ZN(n586) );
  XNOR2_X1 U650 ( .A(n587), .B(n586), .ZN(n589) );
  XOR2_X1 U651 ( .A(G2435), .B(G2438), .Z(n588) );
  XNOR2_X1 U652 ( .A(n589), .B(n588), .ZN(n590) );
  XOR2_X1 U653 ( .A(n591), .B(n590), .Z(n592) );
  AND2_X1 U654 ( .A1(G14), .A2(n592), .ZN(G401) );
  NAND2_X1 U655 ( .A1(G52), .A2(n681), .ZN(n594) );
  NAND2_X1 U656 ( .A1(G64), .A2(n689), .ZN(n593) );
  NAND2_X1 U657 ( .A1(n594), .A2(n593), .ZN(n599) );
  NAND2_X1 U658 ( .A1(G90), .A2(n680), .ZN(n596) );
  NAND2_X1 U659 ( .A1(G77), .A2(n684), .ZN(n595) );
  NAND2_X1 U660 ( .A1(n596), .A2(n595), .ZN(n597) );
  XOR2_X1 U661 ( .A(KEYINPUT9), .B(n597), .Z(n598) );
  NOR2_X1 U662 ( .A1(n599), .A2(n598), .ZN(G171) );
  AND2_X1 U663 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U664 ( .A(G132), .ZN(G219) );
  INV_X1 U665 ( .A(G82), .ZN(G220) );
  INV_X1 U666 ( .A(G120), .ZN(G236) );
  INV_X1 U667 ( .A(G69), .ZN(G235) );
  INV_X1 U668 ( .A(G108), .ZN(G238) );
  NAND2_X1 U669 ( .A1(G7), .A2(G661), .ZN(n600) );
  XNOR2_X1 U670 ( .A(n600), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U671 ( .A(G223), .ZN(n601) );
  NAND2_X1 U672 ( .A1(n601), .A2(G567), .ZN(n602) );
  XNOR2_X1 U673 ( .A(n602), .B(KEYINPUT11), .ZN(n603) );
  XNOR2_X1 U674 ( .A(KEYINPUT69), .B(n603), .ZN(G234) );
  NAND2_X1 U675 ( .A1(n684), .A2(G68), .ZN(n604) );
  XNOR2_X1 U676 ( .A(KEYINPUT70), .B(n604), .ZN(n607) );
  NAND2_X1 U677 ( .A1(n680), .A2(G81), .ZN(n605) );
  XNOR2_X1 U678 ( .A(KEYINPUT12), .B(n605), .ZN(n606) );
  NAND2_X1 U679 ( .A1(n607), .A2(n606), .ZN(n608) );
  XNOR2_X1 U680 ( .A(n608), .B(KEYINPUT13), .ZN(n610) );
  NAND2_X1 U681 ( .A1(G43), .A2(n681), .ZN(n609) );
  NAND2_X1 U682 ( .A1(n610), .A2(n609), .ZN(n613) );
  NAND2_X1 U683 ( .A1(n689), .A2(G56), .ZN(n611) );
  XOR2_X1 U684 ( .A(KEYINPUT14), .B(n611), .Z(n612) );
  NOR2_X1 U685 ( .A1(n613), .A2(n612), .ZN(n614) );
  INV_X1 U686 ( .A(n970), .ZN(n615) );
  XNOR2_X1 U687 ( .A(G860), .B(KEYINPUT72), .ZN(n640) );
  NAND2_X1 U688 ( .A1(n615), .A2(n640), .ZN(G153) );
  INV_X1 U689 ( .A(G171), .ZN(G301) );
  INV_X1 U690 ( .A(G868), .ZN(n701) );
  NOR2_X1 U691 ( .A1(KEYINPUT73), .A2(G171), .ZN(n616) );
  NOR2_X1 U692 ( .A1(KEYINPUT77), .A2(n616), .ZN(n617) );
  NOR2_X1 U693 ( .A1(n701), .A2(n617), .ZN(n633) );
  NAND2_X1 U694 ( .A1(G301), .A2(G868), .ZN(n618) );
  NAND2_X1 U695 ( .A1(n618), .A2(KEYINPUT73), .ZN(n631) );
  NAND2_X1 U696 ( .A1(G66), .A2(n689), .ZN(n627) );
  NAND2_X1 U697 ( .A1(G54), .A2(n681), .ZN(n619) );
  XNOR2_X1 U698 ( .A(n619), .B(KEYINPUT76), .ZN(n622) );
  NAND2_X1 U699 ( .A1(G92), .A2(n680), .ZN(n620) );
  XNOR2_X1 U700 ( .A(n620), .B(KEYINPUT74), .ZN(n621) );
  NAND2_X1 U701 ( .A1(n622), .A2(n621), .ZN(n625) );
  NAND2_X1 U702 ( .A1(G79), .A2(n684), .ZN(n623) );
  XNOR2_X1 U703 ( .A(KEYINPUT75), .B(n623), .ZN(n624) );
  NOR2_X1 U704 ( .A1(n625), .A2(n624), .ZN(n626) );
  NAND2_X1 U705 ( .A1(n627), .A2(n626), .ZN(n628) );
  XNOR2_X1 U706 ( .A(n628), .B(KEYINPUT15), .ZN(n960) );
  NOR2_X1 U707 ( .A1(n960), .A2(KEYINPUT77), .ZN(n629) );
  NAND2_X1 U708 ( .A1(n701), .A2(n629), .ZN(n630) );
  NAND2_X1 U709 ( .A1(n631), .A2(n630), .ZN(n632) );
  NOR2_X1 U710 ( .A1(n633), .A2(n632), .ZN(n635) );
  NAND2_X1 U711 ( .A1(n960), .A2(KEYINPUT77), .ZN(n634) );
  NAND2_X1 U712 ( .A1(n635), .A2(n634), .ZN(G284) );
  XNOR2_X1 U713 ( .A(KEYINPUT80), .B(n701), .ZN(n636) );
  NOR2_X1 U714 ( .A1(G286), .A2(n636), .ZN(n639) );
  NOR2_X1 U715 ( .A1(G868), .A2(G299), .ZN(n637) );
  XOR2_X1 U716 ( .A(KEYINPUT81), .B(n637), .Z(n638) );
  NOR2_X1 U717 ( .A1(n639), .A2(n638), .ZN(G297) );
  INV_X1 U718 ( .A(n960), .ZN(n643) );
  INV_X1 U719 ( .A(G559), .ZN(n641) );
  NOR2_X1 U720 ( .A1(n641), .A2(n640), .ZN(n642) );
  NOR2_X1 U721 ( .A1(n643), .A2(n642), .ZN(n644) );
  XOR2_X1 U722 ( .A(n644), .B(KEYINPUT82), .Z(n645) );
  XNOR2_X1 U723 ( .A(KEYINPUT16), .B(n645), .ZN(G148) );
  NAND2_X1 U724 ( .A1(n960), .A2(G868), .ZN(n646) );
  XOR2_X1 U725 ( .A(KEYINPUT83), .B(n646), .Z(n647) );
  NOR2_X1 U726 ( .A1(G559), .A2(n647), .ZN(n648) );
  XNOR2_X1 U727 ( .A(n648), .B(KEYINPUT84), .ZN(n650) );
  NOR2_X1 U728 ( .A1(n970), .A2(G868), .ZN(n649) );
  NOR2_X1 U729 ( .A1(n650), .A2(n649), .ZN(G282) );
  NAND2_X1 U730 ( .A1(n912), .A2(G123), .ZN(n651) );
  XNOR2_X1 U731 ( .A(n651), .B(KEYINPUT18), .ZN(n653) );
  NAND2_X1 U732 ( .A1(G111), .A2(n913), .ZN(n652) );
  NAND2_X1 U733 ( .A1(n653), .A2(n652), .ZN(n657) );
  NAND2_X1 U734 ( .A1(G135), .A2(n530), .ZN(n655) );
  NAND2_X1 U735 ( .A1(G99), .A2(n909), .ZN(n654) );
  NAND2_X1 U736 ( .A1(n655), .A2(n654), .ZN(n656) );
  NOR2_X1 U737 ( .A1(n657), .A2(n656), .ZN(n1009) );
  XNOR2_X1 U738 ( .A(n1009), .B(G2096), .ZN(n659) );
  INV_X1 U739 ( .A(G2100), .ZN(n658) );
  NAND2_X1 U740 ( .A1(n659), .A2(n658), .ZN(G156) );
  NAND2_X1 U741 ( .A1(G559), .A2(n960), .ZN(n660) );
  XNOR2_X1 U742 ( .A(n660), .B(n970), .ZN(n698) );
  NOR2_X1 U743 ( .A1(n698), .A2(G860), .ZN(n667) );
  NAND2_X1 U744 ( .A1(G93), .A2(n680), .ZN(n662) );
  NAND2_X1 U745 ( .A1(G80), .A2(n684), .ZN(n661) );
  NAND2_X1 U746 ( .A1(n662), .A2(n661), .ZN(n666) );
  NAND2_X1 U747 ( .A1(G55), .A2(n681), .ZN(n664) );
  NAND2_X1 U748 ( .A1(G67), .A2(n689), .ZN(n663) );
  NAND2_X1 U749 ( .A1(n664), .A2(n663), .ZN(n665) );
  OR2_X1 U750 ( .A1(n666), .A2(n665), .ZN(n700) );
  XOR2_X1 U751 ( .A(n667), .B(n700), .Z(G145) );
  NAND2_X1 U752 ( .A1(G88), .A2(n680), .ZN(n669) );
  NAND2_X1 U753 ( .A1(G75), .A2(n684), .ZN(n668) );
  NAND2_X1 U754 ( .A1(n669), .A2(n668), .ZN(n673) );
  NAND2_X1 U755 ( .A1(G50), .A2(n681), .ZN(n671) );
  NAND2_X1 U756 ( .A1(G62), .A2(n689), .ZN(n670) );
  NAND2_X1 U757 ( .A1(n671), .A2(n670), .ZN(n672) );
  NOR2_X1 U758 ( .A1(n673), .A2(n672), .ZN(G166) );
  NAND2_X1 U759 ( .A1(G49), .A2(n681), .ZN(n675) );
  NAND2_X1 U760 ( .A1(G74), .A2(G651), .ZN(n674) );
  NAND2_X1 U761 ( .A1(n675), .A2(n674), .ZN(n676) );
  NOR2_X1 U762 ( .A1(n689), .A2(n676), .ZN(n679) );
  NAND2_X1 U763 ( .A1(n677), .A2(G87), .ZN(n678) );
  NAND2_X1 U764 ( .A1(n679), .A2(n678), .ZN(G288) );
  NAND2_X1 U765 ( .A1(G86), .A2(n680), .ZN(n683) );
  NAND2_X1 U766 ( .A1(G48), .A2(n681), .ZN(n682) );
  NAND2_X1 U767 ( .A1(n683), .A2(n682), .ZN(n688) );
  NAND2_X1 U768 ( .A1(G73), .A2(n684), .ZN(n685) );
  XNOR2_X1 U769 ( .A(n685), .B(KEYINPUT2), .ZN(n686) );
  XNOR2_X1 U770 ( .A(n686), .B(KEYINPUT85), .ZN(n687) );
  NOR2_X1 U771 ( .A1(n688), .A2(n687), .ZN(n691) );
  NAND2_X1 U772 ( .A1(n689), .A2(G61), .ZN(n690) );
  NAND2_X1 U773 ( .A1(n691), .A2(n690), .ZN(G305) );
  XNOR2_X1 U774 ( .A(G166), .B(G290), .ZN(n697) );
  XNOR2_X1 U775 ( .A(KEYINPUT19), .B(KEYINPUT86), .ZN(n693) );
  INV_X1 U776 ( .A(G299), .ZN(n763) );
  XNOR2_X1 U777 ( .A(G288), .B(n763), .ZN(n692) );
  XNOR2_X1 U778 ( .A(n693), .B(n692), .ZN(n694) );
  XOR2_X1 U779 ( .A(n700), .B(n694), .Z(n695) );
  XNOR2_X1 U780 ( .A(n695), .B(G305), .ZN(n696) );
  XNOR2_X1 U781 ( .A(n697), .B(n696), .ZN(n923) );
  XNOR2_X1 U782 ( .A(n698), .B(n923), .ZN(n699) );
  NAND2_X1 U783 ( .A1(n699), .A2(G868), .ZN(n703) );
  NAND2_X1 U784 ( .A1(n701), .A2(n700), .ZN(n702) );
  NAND2_X1 U785 ( .A1(n703), .A2(n702), .ZN(G295) );
  XOR2_X1 U786 ( .A(KEYINPUT87), .B(KEYINPUT21), .Z(n707) );
  NAND2_X1 U787 ( .A1(G2078), .A2(G2084), .ZN(n704) );
  XOR2_X1 U788 ( .A(KEYINPUT20), .B(n704), .Z(n705) );
  NAND2_X1 U789 ( .A1(n705), .A2(G2090), .ZN(n706) );
  XNOR2_X1 U790 ( .A(n707), .B(n706), .ZN(n708) );
  NAND2_X1 U791 ( .A1(G2072), .A2(n708), .ZN(G158) );
  XNOR2_X1 U792 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U793 ( .A1(G235), .A2(G236), .ZN(n709) );
  XOR2_X1 U794 ( .A(KEYINPUT88), .B(n709), .Z(n710) );
  NOR2_X1 U795 ( .A1(G238), .A2(n710), .ZN(n711) );
  NAND2_X1 U796 ( .A1(G57), .A2(n711), .ZN(n880) );
  NAND2_X1 U797 ( .A1(G567), .A2(n880), .ZN(n712) );
  XNOR2_X1 U798 ( .A(n712), .B(KEYINPUT89), .ZN(n717) );
  INV_X1 U799 ( .A(G2106), .ZN(n874) );
  NOR2_X1 U800 ( .A1(G220), .A2(G219), .ZN(n713) );
  XNOR2_X1 U801 ( .A(KEYINPUT22), .B(n713), .ZN(n714) );
  NAND2_X1 U802 ( .A1(n714), .A2(G96), .ZN(n715) );
  NOR2_X1 U803 ( .A1(G218), .A2(n715), .ZN(n882) );
  NOR2_X1 U804 ( .A1(n874), .A2(n882), .ZN(n716) );
  NOR2_X1 U805 ( .A1(n717), .A2(n716), .ZN(G319) );
  INV_X1 U806 ( .A(G319), .ZN(n947) );
  NAND2_X1 U807 ( .A1(G483), .A2(G661), .ZN(n718) );
  NOR2_X1 U808 ( .A1(n947), .A2(n718), .ZN(n878) );
  NAND2_X1 U809 ( .A1(n878), .A2(G36), .ZN(G176) );
  XOR2_X1 U810 ( .A(KEYINPUT92), .B(G166), .Z(G303) );
  NAND2_X1 U811 ( .A1(G160), .A2(G40), .ZN(n732) );
  NOR2_X1 U812 ( .A1(n734), .A2(n732), .ZN(n720) );
  XOR2_X1 U813 ( .A(KEYINPUT93), .B(n720), .Z(n869) );
  XNOR2_X1 U814 ( .A(G2067), .B(KEYINPUT37), .ZN(n867) );
  NAND2_X1 U815 ( .A1(G140), .A2(n530), .ZN(n722) );
  NAND2_X1 U816 ( .A1(G104), .A2(n909), .ZN(n721) );
  NAND2_X1 U817 ( .A1(n722), .A2(n721), .ZN(n723) );
  XNOR2_X1 U818 ( .A(KEYINPUT34), .B(n723), .ZN(n729) );
  NAND2_X1 U819 ( .A1(n913), .A2(G116), .ZN(n724) );
  XNOR2_X1 U820 ( .A(n724), .B(KEYINPUT94), .ZN(n726) );
  NAND2_X1 U821 ( .A1(G128), .A2(n912), .ZN(n725) );
  NAND2_X1 U822 ( .A1(n726), .A2(n725), .ZN(n727) );
  XOR2_X1 U823 ( .A(n727), .B(KEYINPUT35), .Z(n728) );
  NOR2_X1 U824 ( .A1(n729), .A2(n728), .ZN(n730) );
  XOR2_X1 U825 ( .A(KEYINPUT36), .B(n730), .Z(n731) );
  XNOR2_X1 U826 ( .A(KEYINPUT95), .B(n731), .ZN(n919) );
  NOR2_X1 U827 ( .A1(n867), .A2(n919), .ZN(n1016) );
  NAND2_X1 U828 ( .A1(n869), .A2(n1016), .ZN(n865) );
  INV_X1 U829 ( .A(n865), .ZN(n835) );
  INV_X1 U830 ( .A(n732), .ZN(n733) );
  INV_X1 U831 ( .A(KEYINPUT64), .ZN(n735) );
  XNOR2_X2 U832 ( .A(n736), .B(n735), .ZN(n770) );
  NAND2_X1 U833 ( .A1(n770), .A2(G1996), .ZN(n737) );
  XNOR2_X1 U834 ( .A(n737), .B(KEYINPUT26), .ZN(n739) );
  NAND2_X1 U835 ( .A1(n775), .A2(G1341), .ZN(n738) );
  NAND2_X1 U836 ( .A1(n739), .A2(n738), .ZN(n740) );
  NAND2_X1 U837 ( .A1(n757), .A2(n960), .ZN(n751) );
  NAND2_X1 U838 ( .A1(G2067), .A2(n770), .ZN(n743) );
  XNOR2_X1 U839 ( .A(KEYINPUT104), .B(n743), .ZN(n744) );
  NAND2_X1 U840 ( .A1(n775), .A2(G1348), .ZN(n746) );
  NAND2_X1 U841 ( .A1(n744), .A2(n746), .ZN(n745) );
  NOR2_X1 U842 ( .A1(KEYINPUT103), .A2(n745), .ZN(n749) );
  NAND2_X1 U843 ( .A1(KEYINPUT104), .A2(KEYINPUT103), .ZN(n747) );
  NOR2_X1 U844 ( .A1(n747), .A2(n746), .ZN(n748) );
  NOR2_X1 U845 ( .A1(n749), .A2(n748), .ZN(n750) );
  NAND2_X1 U846 ( .A1(n751), .A2(n750), .ZN(n756) );
  NAND2_X1 U847 ( .A1(G2072), .A2(n770), .ZN(n752) );
  XNOR2_X1 U848 ( .A(n752), .B(KEYINPUT27), .ZN(n754) );
  XOR2_X1 U849 ( .A(KEYINPUT102), .B(G1956), .Z(n981) );
  NOR2_X1 U850 ( .A1(n770), .A2(n981), .ZN(n753) );
  NOR2_X1 U851 ( .A1(n754), .A2(n753), .ZN(n762) );
  NOR2_X1 U852 ( .A1(n763), .A2(n762), .ZN(n755) );
  XOR2_X1 U853 ( .A(n755), .B(KEYINPUT28), .Z(n761) );
  AND2_X1 U854 ( .A1(n756), .A2(n761), .ZN(n760) );
  XNOR2_X1 U855 ( .A(n758), .B(KEYINPUT105), .ZN(n759) );
  NAND2_X1 U856 ( .A1(n760), .A2(n759), .ZN(n767) );
  INV_X1 U857 ( .A(n761), .ZN(n765) );
  NAND2_X1 U858 ( .A1(n763), .A2(n762), .ZN(n764) );
  OR2_X1 U859 ( .A1(n765), .A2(n764), .ZN(n766) );
  XOR2_X1 U860 ( .A(n768), .B(KEYINPUT29), .Z(n774) );
  XOR2_X1 U861 ( .A(G2078), .B(KEYINPUT25), .Z(n1036) );
  NOR2_X1 U862 ( .A1(n775), .A2(n1036), .ZN(n769) );
  XNOR2_X1 U863 ( .A(n769), .B(KEYINPUT101), .ZN(n772) );
  OR2_X1 U864 ( .A1(n770), .A2(G1961), .ZN(n771) );
  NAND2_X1 U865 ( .A1(n772), .A2(n771), .ZN(n780) );
  NAND2_X1 U866 ( .A1(G171), .A2(n780), .ZN(n773) );
  NAND2_X1 U867 ( .A1(n774), .A2(n773), .ZN(n785) );
  XNOR2_X2 U868 ( .A(KEYINPUT100), .B(n776), .ZN(n831) );
  NOR2_X1 U869 ( .A1(n831), .A2(G1966), .ZN(n797) );
  NOR2_X1 U870 ( .A1(n775), .A2(G2084), .ZN(n795) );
  NOR2_X1 U871 ( .A1(n797), .A2(n795), .ZN(n777) );
  NAND2_X1 U872 ( .A1(G8), .A2(n777), .ZN(n778) );
  XNOR2_X1 U873 ( .A(KEYINPUT30), .B(n778), .ZN(n779) );
  NOR2_X1 U874 ( .A1(G168), .A2(n779), .ZN(n782) );
  NOR2_X1 U875 ( .A1(G171), .A2(n780), .ZN(n781) );
  NOR2_X1 U876 ( .A1(n782), .A2(n781), .ZN(n783) );
  XOR2_X1 U877 ( .A(KEYINPUT31), .B(n783), .Z(n784) );
  NAND2_X1 U878 ( .A1(n785), .A2(n784), .ZN(n799) );
  NAND2_X1 U879 ( .A1(n799), .A2(G286), .ZN(n790) );
  NOR2_X1 U880 ( .A1(n831), .A2(G1971), .ZN(n787) );
  NOR2_X1 U881 ( .A1(n775), .A2(G2090), .ZN(n786) );
  NOR2_X1 U882 ( .A1(n787), .A2(n786), .ZN(n788) );
  NAND2_X1 U883 ( .A1(G303), .A2(n788), .ZN(n789) );
  NAND2_X1 U884 ( .A1(n790), .A2(n789), .ZN(n791) );
  XNOR2_X1 U885 ( .A(n791), .B(KEYINPUT106), .ZN(n792) );
  NAND2_X1 U886 ( .A1(n792), .A2(G8), .ZN(n794) );
  XNOR2_X1 U887 ( .A(n794), .B(n793), .ZN(n814) );
  AND2_X1 U888 ( .A1(G8), .A2(n795), .ZN(n796) );
  NOR2_X1 U889 ( .A1(n797), .A2(n796), .ZN(n798) );
  AND2_X1 U890 ( .A1(n799), .A2(n798), .ZN(n807) );
  INV_X1 U891 ( .A(n831), .ZN(n808) );
  OR2_X1 U892 ( .A1(n807), .A2(n808), .ZN(n800) );
  INV_X1 U893 ( .A(G8), .ZN(n803) );
  NOR2_X1 U894 ( .A1(G303), .A2(G2090), .ZN(n801) );
  XNOR2_X1 U895 ( .A(n801), .B(KEYINPUT109), .ZN(n802) );
  NOR2_X1 U896 ( .A1(n803), .A2(n802), .ZN(n804) );
  NAND2_X1 U897 ( .A1(n533), .A2(n531), .ZN(n826) );
  NAND2_X1 U898 ( .A1(G288), .A2(G1976), .ZN(n805) );
  XNOR2_X1 U899 ( .A(n805), .B(KEYINPUT107), .ZN(n956) );
  NOR2_X1 U900 ( .A1(n831), .A2(n956), .ZN(n806) );
  NOR2_X1 U901 ( .A1(KEYINPUT33), .A2(n806), .ZN(n819) );
  INV_X1 U902 ( .A(KEYINPUT33), .ZN(n816) );
  NOR2_X1 U903 ( .A1(G1976), .A2(G288), .ZN(n957) );
  NAND2_X1 U904 ( .A1(n957), .A2(n808), .ZN(n809) );
  NOR2_X1 U905 ( .A1(n816), .A2(n809), .ZN(n810) );
  XNOR2_X1 U906 ( .A(n810), .B(KEYINPUT108), .ZN(n821) );
  INV_X1 U907 ( .A(n821), .ZN(n811) );
  NAND2_X1 U908 ( .A1(n532), .A2(n811), .ZN(n812) );
  XNOR2_X1 U909 ( .A(G1981), .B(G305), .ZN(n972) );
  OR2_X1 U910 ( .A1(n812), .A2(n972), .ZN(n813) );
  NOR2_X1 U911 ( .A1(G1971), .A2(G303), .ZN(n815) );
  NOR2_X1 U912 ( .A1(n957), .A2(n815), .ZN(n817) );
  AND2_X1 U913 ( .A1(n817), .A2(n816), .ZN(n818) );
  OR2_X1 U914 ( .A1(n819), .A2(n818), .ZN(n820) );
  OR2_X1 U915 ( .A1(n821), .A2(n820), .ZN(n822) );
  OR2_X1 U916 ( .A1(n972), .A2(n822), .ZN(n823) );
  NAND2_X1 U917 ( .A1(n824), .A2(n823), .ZN(n825) );
  NOR2_X1 U918 ( .A1(n826), .A2(n825), .ZN(n828) );
  XNOR2_X1 U919 ( .A(n828), .B(n827), .ZN(n833) );
  NOR2_X1 U920 ( .A1(G1981), .A2(G305), .ZN(n829) );
  XOR2_X1 U921 ( .A(n829), .B(KEYINPUT24), .Z(n830) );
  NOR2_X1 U922 ( .A1(n831), .A2(n830), .ZN(n832) );
  NOR2_X1 U923 ( .A1(n833), .A2(n832), .ZN(n834) );
  NOR2_X1 U924 ( .A1(n835), .A2(n834), .ZN(n857) );
  NAND2_X1 U925 ( .A1(G129), .A2(n912), .ZN(n836) );
  XNOR2_X1 U926 ( .A(n836), .B(KEYINPUT96), .ZN(n845) );
  NAND2_X1 U927 ( .A1(G105), .A2(n909), .ZN(n837) );
  XNOR2_X1 U928 ( .A(n837), .B(KEYINPUT98), .ZN(n838) );
  XNOR2_X1 U929 ( .A(n838), .B(KEYINPUT38), .ZN(n840) );
  NAND2_X1 U930 ( .A1(G141), .A2(n530), .ZN(n839) );
  NAND2_X1 U931 ( .A1(n840), .A2(n839), .ZN(n843) );
  NAND2_X1 U932 ( .A1(G117), .A2(n913), .ZN(n841) );
  XNOR2_X1 U933 ( .A(KEYINPUT97), .B(n841), .ZN(n842) );
  NOR2_X1 U934 ( .A1(n843), .A2(n842), .ZN(n844) );
  NAND2_X1 U935 ( .A1(n845), .A2(n844), .ZN(n894) );
  NAND2_X1 U936 ( .A1(n894), .A2(G1996), .ZN(n853) );
  NAND2_X1 U937 ( .A1(G119), .A2(n912), .ZN(n847) );
  NAND2_X1 U938 ( .A1(G131), .A2(n530), .ZN(n846) );
  NAND2_X1 U939 ( .A1(n847), .A2(n846), .ZN(n851) );
  NAND2_X1 U940 ( .A1(G107), .A2(n913), .ZN(n849) );
  NAND2_X1 U941 ( .A1(G95), .A2(n909), .ZN(n848) );
  NAND2_X1 U942 ( .A1(n849), .A2(n848), .ZN(n850) );
  OR2_X1 U943 ( .A1(n851), .A2(n850), .ZN(n890) );
  NAND2_X1 U944 ( .A1(G1991), .A2(n890), .ZN(n852) );
  NAND2_X1 U945 ( .A1(n853), .A2(n852), .ZN(n854) );
  XNOR2_X1 U946 ( .A(n854), .B(KEYINPUT99), .ZN(n859) );
  XOR2_X1 U947 ( .A(G1986), .B(G290), .Z(n959) );
  NAND2_X1 U948 ( .A1(n859), .A2(n959), .ZN(n855) );
  NAND2_X1 U949 ( .A1(n855), .A2(n869), .ZN(n856) );
  NAND2_X1 U950 ( .A1(n857), .A2(n856), .ZN(n872) );
  NOR2_X1 U951 ( .A1(G1986), .A2(G290), .ZN(n858) );
  NOR2_X1 U952 ( .A1(G1991), .A2(n890), .ZN(n1010) );
  NOR2_X1 U953 ( .A1(n858), .A2(n1010), .ZN(n860) );
  INV_X1 U954 ( .A(n859), .ZN(n1012) );
  NOR2_X1 U955 ( .A1(n860), .A2(n1012), .ZN(n862) );
  NOR2_X1 U956 ( .A1(G1996), .A2(n894), .ZN(n861) );
  XOR2_X1 U957 ( .A(KEYINPUT111), .B(n861), .Z(n1007) );
  NOR2_X1 U958 ( .A1(n862), .A2(n1007), .ZN(n863) );
  XNOR2_X1 U959 ( .A(n863), .B(KEYINPUT39), .ZN(n864) );
  XNOR2_X1 U960 ( .A(n864), .B(KEYINPUT112), .ZN(n866) );
  NAND2_X1 U961 ( .A1(n866), .A2(n865), .ZN(n868) );
  NAND2_X1 U962 ( .A1(n867), .A2(n919), .ZN(n1023) );
  NAND2_X1 U963 ( .A1(n868), .A2(n1023), .ZN(n870) );
  NAND2_X1 U964 ( .A1(n870), .A2(n869), .ZN(n871) );
  NAND2_X1 U965 ( .A1(n872), .A2(n871), .ZN(n873) );
  XNOR2_X1 U966 ( .A(n873), .B(KEYINPUT40), .ZN(G329) );
  NOR2_X1 U967 ( .A1(n874), .A2(G223), .ZN(n875) );
  XNOR2_X1 U968 ( .A(n875), .B(KEYINPUT113), .ZN(G217) );
  AND2_X1 U969 ( .A1(G15), .A2(G2), .ZN(n876) );
  NAND2_X1 U970 ( .A1(G661), .A2(n876), .ZN(G259) );
  NAND2_X1 U971 ( .A1(G3), .A2(G1), .ZN(n877) );
  XNOR2_X1 U972 ( .A(KEYINPUT114), .B(n877), .ZN(n879) );
  NAND2_X1 U973 ( .A1(n879), .A2(n878), .ZN(G188) );
  INV_X1 U975 ( .A(G96), .ZN(G221) );
  INV_X1 U976 ( .A(n880), .ZN(n881) );
  NAND2_X1 U977 ( .A1(n882), .A2(n881), .ZN(G261) );
  INV_X1 U978 ( .A(G261), .ZN(G325) );
  NAND2_X1 U979 ( .A1(n912), .A2(G124), .ZN(n883) );
  XNOR2_X1 U980 ( .A(n883), .B(KEYINPUT44), .ZN(n885) );
  NAND2_X1 U981 ( .A1(G112), .A2(n913), .ZN(n884) );
  NAND2_X1 U982 ( .A1(n885), .A2(n884), .ZN(n889) );
  NAND2_X1 U983 ( .A1(G136), .A2(n530), .ZN(n887) );
  NAND2_X1 U984 ( .A1(G100), .A2(n909), .ZN(n886) );
  NAND2_X1 U985 ( .A1(n887), .A2(n886), .ZN(n888) );
  NOR2_X1 U986 ( .A1(n889), .A2(n888), .ZN(G162) );
  XNOR2_X1 U987 ( .A(KEYINPUT48), .B(KEYINPUT118), .ZN(n892) );
  XNOR2_X1 U988 ( .A(n890), .B(KEYINPUT46), .ZN(n891) );
  XNOR2_X1 U989 ( .A(n892), .B(n891), .ZN(n908) );
  XOR2_X1 U990 ( .A(G162), .B(n1009), .Z(n893) );
  XNOR2_X1 U991 ( .A(n894), .B(n893), .ZN(n904) );
  NAND2_X1 U992 ( .A1(G142), .A2(n530), .ZN(n896) );
  NAND2_X1 U993 ( .A1(G106), .A2(n909), .ZN(n895) );
  NAND2_X1 U994 ( .A1(n896), .A2(n895), .ZN(n897) );
  XNOR2_X1 U995 ( .A(n897), .B(KEYINPUT45), .ZN(n899) );
  NAND2_X1 U996 ( .A1(G118), .A2(n913), .ZN(n898) );
  NAND2_X1 U997 ( .A1(n899), .A2(n898), .ZN(n902) );
  NAND2_X1 U998 ( .A1(G130), .A2(n912), .ZN(n900) );
  XNOR2_X1 U999 ( .A(KEYINPUT117), .B(n900), .ZN(n901) );
  NOR2_X1 U1000 ( .A1(n902), .A2(n901), .ZN(n903) );
  XOR2_X1 U1001 ( .A(n904), .B(n903), .Z(n906) );
  XNOR2_X1 U1002 ( .A(G164), .B(G160), .ZN(n905) );
  XNOR2_X1 U1003 ( .A(n906), .B(n905), .ZN(n907) );
  XNOR2_X1 U1004 ( .A(n908), .B(n907), .ZN(n921) );
  NAND2_X1 U1005 ( .A1(G139), .A2(n530), .ZN(n911) );
  NAND2_X1 U1006 ( .A1(G103), .A2(n909), .ZN(n910) );
  NAND2_X1 U1007 ( .A1(n911), .A2(n910), .ZN(n918) );
  NAND2_X1 U1008 ( .A1(G127), .A2(n912), .ZN(n915) );
  NAND2_X1 U1009 ( .A1(G115), .A2(n913), .ZN(n914) );
  NAND2_X1 U1010 ( .A1(n915), .A2(n914), .ZN(n916) );
  XOR2_X1 U1011 ( .A(KEYINPUT47), .B(n916), .Z(n917) );
  NOR2_X1 U1012 ( .A1(n918), .A2(n917), .ZN(n1019) );
  XNOR2_X1 U1013 ( .A(n919), .B(n1019), .ZN(n920) );
  XNOR2_X1 U1014 ( .A(n921), .B(n920), .ZN(n922) );
  NOR2_X1 U1015 ( .A1(G37), .A2(n922), .ZN(G395) );
  XOR2_X1 U1016 ( .A(n923), .B(G286), .Z(n925) );
  XNOR2_X1 U1017 ( .A(G171), .B(n960), .ZN(n924) );
  XNOR2_X1 U1018 ( .A(n925), .B(n924), .ZN(n926) );
  XNOR2_X1 U1019 ( .A(n926), .B(n970), .ZN(n927) );
  NOR2_X1 U1020 ( .A1(G37), .A2(n927), .ZN(G397) );
  XOR2_X1 U1021 ( .A(KEYINPUT115), .B(G2090), .Z(n929) );
  XNOR2_X1 U1022 ( .A(G2067), .B(G2084), .ZN(n928) );
  XNOR2_X1 U1023 ( .A(n929), .B(n928), .ZN(n930) );
  XOR2_X1 U1024 ( .A(n930), .B(G2100), .Z(n932) );
  XNOR2_X1 U1025 ( .A(G2078), .B(G2072), .ZN(n931) );
  XNOR2_X1 U1026 ( .A(n932), .B(n931), .ZN(n936) );
  XOR2_X1 U1027 ( .A(G2096), .B(G2678), .Z(n934) );
  XNOR2_X1 U1028 ( .A(KEYINPUT42), .B(KEYINPUT43), .ZN(n933) );
  XNOR2_X1 U1029 ( .A(n934), .B(n933), .ZN(n935) );
  XOR2_X1 U1030 ( .A(n936), .B(n935), .Z(G227) );
  XNOR2_X1 U1031 ( .A(G1996), .B(KEYINPUT116), .ZN(n946) );
  XOR2_X1 U1032 ( .A(G1956), .B(G1961), .Z(n938) );
  XNOR2_X1 U1033 ( .A(G1991), .B(G1981), .ZN(n937) );
  XNOR2_X1 U1034 ( .A(n938), .B(n937), .ZN(n942) );
  XOR2_X1 U1035 ( .A(G1966), .B(G1971), .Z(n940) );
  XNOR2_X1 U1036 ( .A(G1986), .B(G1976), .ZN(n939) );
  XNOR2_X1 U1037 ( .A(n940), .B(n939), .ZN(n941) );
  XOR2_X1 U1038 ( .A(n942), .B(n941), .Z(n944) );
  XNOR2_X1 U1039 ( .A(G2474), .B(KEYINPUT41), .ZN(n943) );
  XNOR2_X1 U1040 ( .A(n944), .B(n943), .ZN(n945) );
  XNOR2_X1 U1041 ( .A(n946), .B(n945), .ZN(G229) );
  NOR2_X1 U1042 ( .A1(G401), .A2(n947), .ZN(n952) );
  NOR2_X1 U1043 ( .A1(G227), .A2(G229), .ZN(n948) );
  XOR2_X1 U1044 ( .A(KEYINPUT49), .B(n948), .Z(n949) );
  XNOR2_X1 U1045 ( .A(n949), .B(KEYINPUT119), .ZN(n950) );
  NOR2_X1 U1046 ( .A1(G397), .A2(n950), .ZN(n951) );
  NAND2_X1 U1047 ( .A1(n952), .A2(n951), .ZN(n953) );
  NOR2_X1 U1048 ( .A1(G395), .A2(n953), .ZN(n954) );
  XOR2_X1 U1049 ( .A(KEYINPUT120), .B(n954), .Z(G225) );
  XNOR2_X1 U1050 ( .A(KEYINPUT121), .B(G225), .ZN(G308) );
  INV_X1 U1051 ( .A(G57), .ZN(G237) );
  XNOR2_X1 U1052 ( .A(KEYINPUT56), .B(G16), .ZN(n979) );
  XNOR2_X1 U1053 ( .A(G1956), .B(G299), .ZN(n955) );
  NOR2_X1 U1054 ( .A1(n956), .A2(n955), .ZN(n966) );
  INV_X1 U1055 ( .A(n957), .ZN(n958) );
  NAND2_X1 U1056 ( .A1(n959), .A2(n958), .ZN(n964) );
  XNOR2_X1 U1057 ( .A(G1348), .B(n960), .ZN(n962) );
  XNOR2_X1 U1058 ( .A(G171), .B(G1961), .ZN(n961) );
  NAND2_X1 U1059 ( .A1(n962), .A2(n961), .ZN(n963) );
  NOR2_X1 U1060 ( .A1(n964), .A2(n963), .ZN(n965) );
  NAND2_X1 U1061 ( .A1(n966), .A2(n965), .ZN(n969) );
  XNOR2_X1 U1062 ( .A(G303), .B(G1971), .ZN(n967) );
  XNOR2_X1 U1063 ( .A(KEYINPUT124), .B(n967), .ZN(n968) );
  NOR2_X1 U1064 ( .A1(n969), .A2(n968), .ZN(n977) );
  XNOR2_X1 U1065 ( .A(n970), .B(G1341), .ZN(n975) );
  XOR2_X1 U1066 ( .A(G1966), .B(G168), .Z(n971) );
  NOR2_X1 U1067 ( .A1(n972), .A2(n971), .ZN(n973) );
  XNOR2_X1 U1068 ( .A(KEYINPUT57), .B(n973), .ZN(n974) );
  NOR2_X1 U1069 ( .A1(n975), .A2(n974), .ZN(n976) );
  NAND2_X1 U1070 ( .A1(n977), .A2(n976), .ZN(n978) );
  NAND2_X1 U1071 ( .A1(n979), .A2(n978), .ZN(n980) );
  XNOR2_X1 U1072 ( .A(n980), .B(KEYINPUT125), .ZN(n1005) );
  XNOR2_X1 U1073 ( .A(n981), .B(G20), .ZN(n985) );
  XNOR2_X1 U1074 ( .A(G1981), .B(G6), .ZN(n983) );
  XNOR2_X1 U1075 ( .A(G19), .B(G1341), .ZN(n982) );
  NOR2_X1 U1076 ( .A1(n983), .A2(n982), .ZN(n984) );
  NAND2_X1 U1077 ( .A1(n985), .A2(n984), .ZN(n988) );
  XOR2_X1 U1078 ( .A(KEYINPUT59), .B(G1348), .Z(n986) );
  XNOR2_X1 U1079 ( .A(G4), .B(n986), .ZN(n987) );
  NOR2_X1 U1080 ( .A1(n988), .A2(n987), .ZN(n989) );
  XOR2_X1 U1081 ( .A(KEYINPUT60), .B(n989), .Z(n991) );
  XNOR2_X1 U1082 ( .A(G1961), .B(G5), .ZN(n990) );
  NOR2_X1 U1083 ( .A1(n991), .A2(n990), .ZN(n1001) );
  XNOR2_X1 U1084 ( .A(G1976), .B(G23), .ZN(n993) );
  XNOR2_X1 U1085 ( .A(G22), .B(G1971), .ZN(n992) );
  NOR2_X1 U1086 ( .A1(n993), .A2(n992), .ZN(n994) );
  XOR2_X1 U1087 ( .A(KEYINPUT126), .B(n994), .Z(n996) );
  XNOR2_X1 U1088 ( .A(G1986), .B(G24), .ZN(n995) );
  NOR2_X1 U1089 ( .A1(n996), .A2(n995), .ZN(n997) );
  XOR2_X1 U1090 ( .A(KEYINPUT58), .B(n997), .Z(n999) );
  XNOR2_X1 U1091 ( .A(G1966), .B(G21), .ZN(n998) );
  NOR2_X1 U1092 ( .A1(n999), .A2(n998), .ZN(n1000) );
  NAND2_X1 U1093 ( .A1(n1001), .A2(n1000), .ZN(n1002) );
  XNOR2_X1 U1094 ( .A(KEYINPUT61), .B(n1002), .ZN(n1003) );
  NOR2_X1 U1095 ( .A1(n1003), .A2(G16), .ZN(n1004) );
  NOR2_X1 U1096 ( .A1(n1005), .A2(n1004), .ZN(n1032) );
  XOR2_X1 U1097 ( .A(G2090), .B(G162), .Z(n1006) );
  NOR2_X1 U1098 ( .A1(n1007), .A2(n1006), .ZN(n1008) );
  XOR2_X1 U1099 ( .A(KEYINPUT51), .B(n1008), .Z(n1018) );
  NOR2_X1 U1100 ( .A1(n1010), .A2(n1009), .ZN(n1014) );
  XOR2_X1 U1101 ( .A(G160), .B(G2084), .Z(n1011) );
  NOR2_X1 U1102 ( .A1(n1012), .A2(n1011), .ZN(n1013) );
  NAND2_X1 U1103 ( .A1(n1014), .A2(n1013), .ZN(n1015) );
  NOR2_X1 U1104 ( .A1(n1016), .A2(n1015), .ZN(n1017) );
  NAND2_X1 U1105 ( .A1(n1018), .A2(n1017), .ZN(n1026) );
  XOR2_X1 U1106 ( .A(G2072), .B(n1019), .Z(n1021) );
  XOR2_X1 U1107 ( .A(G164), .B(G2078), .Z(n1020) );
  NOR2_X1 U1108 ( .A1(n1021), .A2(n1020), .ZN(n1022) );
  XNOR2_X1 U1109 ( .A(n1022), .B(KEYINPUT50), .ZN(n1024) );
  NAND2_X1 U1110 ( .A1(n1024), .A2(n1023), .ZN(n1025) );
  NOR2_X1 U1111 ( .A1(n1026), .A2(n1025), .ZN(n1027) );
  XOR2_X1 U1112 ( .A(KEYINPUT52), .B(n1027), .Z(n1028) );
  NOR2_X1 U1113 ( .A1(KEYINPUT55), .A2(n1028), .ZN(n1029) );
  XOR2_X1 U1114 ( .A(KEYINPUT122), .B(n1029), .Z(n1030) );
  NAND2_X1 U1115 ( .A1(G29), .A2(n1030), .ZN(n1031) );
  NAND2_X1 U1116 ( .A1(n1032), .A2(n1031), .ZN(n1055) );
  XOR2_X1 U1117 ( .A(G1991), .B(G25), .Z(n1033) );
  NAND2_X1 U1118 ( .A1(n1033), .A2(G28), .ZN(n1042) );
  XNOR2_X1 U1119 ( .A(G2067), .B(G26), .ZN(n1035) );
  XNOR2_X1 U1120 ( .A(G33), .B(G2072), .ZN(n1034) );
  NOR2_X1 U1121 ( .A1(n1035), .A2(n1034), .ZN(n1040) );
  XNOR2_X1 U1122 ( .A(G1996), .B(G32), .ZN(n1038) );
  XNOR2_X1 U1123 ( .A(G27), .B(n1036), .ZN(n1037) );
  NOR2_X1 U1124 ( .A1(n1038), .A2(n1037), .ZN(n1039) );
  NAND2_X1 U1125 ( .A1(n1040), .A2(n1039), .ZN(n1041) );
  NOR2_X1 U1126 ( .A1(n1042), .A2(n1041), .ZN(n1043) );
  XOR2_X1 U1127 ( .A(KEYINPUT53), .B(n1043), .Z(n1046) );
  XOR2_X1 U1128 ( .A(KEYINPUT54), .B(G34), .Z(n1044) );
  XNOR2_X1 U1129 ( .A(G2084), .B(n1044), .ZN(n1045) );
  NAND2_X1 U1130 ( .A1(n1046), .A2(n1045), .ZN(n1049) );
  XOR2_X1 U1131 ( .A(KEYINPUT123), .B(G2090), .Z(n1047) );
  XNOR2_X1 U1132 ( .A(G35), .B(n1047), .ZN(n1048) );
  NOR2_X1 U1133 ( .A1(n1049), .A2(n1048), .ZN(n1050) );
  XNOR2_X1 U1134 ( .A(KEYINPUT55), .B(n1050), .ZN(n1052) );
  INV_X1 U1135 ( .A(G29), .ZN(n1051) );
  NAND2_X1 U1136 ( .A1(n1052), .A2(n1051), .ZN(n1053) );
  NAND2_X1 U1137 ( .A1(n1053), .A2(G11), .ZN(n1054) );
  NOR2_X1 U1138 ( .A1(n1055), .A2(n1054), .ZN(n1056) );
  XNOR2_X1 U1139 ( .A(n1056), .B(KEYINPUT62), .ZN(G311) );
  INV_X1 U1140 ( .A(G311), .ZN(G150) );
endmodule

