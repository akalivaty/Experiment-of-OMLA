//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 1 1 0 0 1 1 1 1 0 1 1 0 0 0 1 1 0 0 1 1 1 0 1 1 1 0 1 1 1 1 1 1 0 0 0 1 0 1 1 1 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 0 1 1 1 1 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:42:26 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n203, new_n204, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n237, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n245, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1195, new_n1196, new_n1197, new_n1198, new_n1199,
    new_n1200, new_n1201, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1217, new_n1218,
    new_n1219, new_n1220, new_n1222, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1273, new_n1274, new_n1275,
    new_n1276, new_n1277, new_n1278, new_n1279;
  NOR4_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .A4(G77), .ZN(G353));
  OAI21_X1  g0001(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0002(.A(G1), .ZN(new_n203));
  INV_X1    g0003(.A(G20), .ZN(new_n204));
  NOR2_X1   g0004(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  INV_X1    g0005(.A(new_n205), .ZN(new_n206));
  AOI22_X1  g0006(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n207));
  XOR2_X1   g0007(.A(new_n207), .B(KEYINPUT65), .Z(new_n208));
  NAND2_X1  g0008(.A1(G68), .A2(G238), .ZN(new_n209));
  NAND2_X1  g0009(.A1(G77), .A2(G244), .ZN(new_n210));
  NAND2_X1  g0010(.A1(G50), .A2(G226), .ZN(new_n211));
  NAND2_X1  g0011(.A1(G116), .A2(G270), .ZN(new_n212));
  NAND4_X1  g0012(.A1(new_n209), .A2(new_n210), .A3(new_n211), .A4(new_n212), .ZN(new_n213));
  INV_X1    g0013(.A(new_n213), .ZN(new_n214));
  OAI21_X1  g0014(.A(new_n208), .B1(KEYINPUT64), .B2(new_n214), .ZN(new_n215));
  AOI22_X1  g0015(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n216));
  INV_X1    g0016(.A(KEYINPUT64), .ZN(new_n217));
  OAI21_X1  g0017(.A(new_n216), .B1(new_n213), .B2(new_n217), .ZN(new_n218));
  OAI21_X1  g0018(.A(new_n206), .B1(new_n215), .B2(new_n218), .ZN(new_n219));
  NAND2_X1  g0019(.A1(new_n219), .A2(KEYINPUT1), .ZN(new_n220));
  XOR2_X1   g0020(.A(new_n220), .B(KEYINPUT66), .Z(new_n221));
  NOR2_X1   g0021(.A1(new_n206), .A2(G13), .ZN(new_n222));
  OAI211_X1 g0022(.A(new_n222), .B(G250), .C1(G257), .C2(G264), .ZN(new_n223));
  XNOR2_X1  g0023(.A(new_n223), .B(KEYINPUT0), .ZN(new_n224));
  NAND3_X1  g0024(.A1(G1), .A2(G13), .A3(G20), .ZN(new_n225));
  OAI21_X1  g0025(.A(G50), .B1(G58), .B2(G68), .ZN(new_n226));
  OAI221_X1 g0026(.A(new_n224), .B1(new_n225), .B2(new_n226), .C1(new_n219), .C2(KEYINPUT1), .ZN(new_n227));
  NOR2_X1   g0027(.A1(new_n221), .A2(new_n227), .ZN(G361));
  XNOR2_X1  g0028(.A(G238), .B(G244), .ZN(new_n229));
  XNOR2_X1  g0029(.A(new_n229), .B(G232), .ZN(new_n230));
  XNOR2_X1  g0030(.A(KEYINPUT2), .B(G226), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n230), .B(new_n231), .ZN(new_n232));
  XOR2_X1   g0032(.A(G264), .B(G270), .Z(new_n233));
  XNOR2_X1  g0033(.A(G250), .B(G257), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n232), .B(new_n235), .ZN(G358));
  XOR2_X1   g0036(.A(G107), .B(G116), .Z(new_n237));
  XNOR2_X1  g0037(.A(new_n237), .B(KEYINPUT69), .ZN(new_n238));
  XNOR2_X1  g0038(.A(G87), .B(G97), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XOR2_X1   g0040(.A(G68), .B(G77), .Z(new_n241));
  XNOR2_X1  g0041(.A(G50), .B(G58), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XNOR2_X1  g0043(.A(KEYINPUT67), .B(KEYINPUT68), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n240), .B(new_n245), .ZN(G351));
  XNOR2_X1  g0046(.A(KEYINPUT3), .B(G33), .ZN(new_n247));
  INV_X1    g0047(.A(G1698), .ZN(new_n248));
  NAND3_X1  g0048(.A1(new_n247), .A2(G222), .A3(new_n248), .ZN(new_n249));
  NAND3_X1  g0049(.A1(new_n247), .A2(G223), .A3(G1698), .ZN(new_n250));
  INV_X1    g0050(.A(G77), .ZN(new_n251));
  OAI211_X1 g0051(.A(new_n249), .B(new_n250), .C1(new_n251), .C2(new_n247), .ZN(new_n252));
  NAND2_X1  g0052(.A1(G1), .A2(G13), .ZN(new_n253));
  AOI21_X1  g0053(.A(new_n253), .B1(G33), .B2(G41), .ZN(new_n254));
  NAND2_X1  g0054(.A1(new_n252), .A2(new_n254), .ZN(new_n255));
  OAI21_X1  g0055(.A(new_n203), .B1(G41), .B2(G45), .ZN(new_n256));
  INV_X1    g0056(.A(G274), .ZN(new_n257));
  NOR2_X1   g0057(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  INV_X1    g0058(.A(G41), .ZN(new_n259));
  INV_X1    g0059(.A(G45), .ZN(new_n260));
  AOI21_X1  g0060(.A(G1), .B1(new_n259), .B2(new_n260), .ZN(new_n261));
  NOR2_X1   g0061(.A1(new_n254), .A2(new_n261), .ZN(new_n262));
  AOI21_X1  g0062(.A(new_n258), .B1(new_n262), .B2(G226), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n255), .A2(new_n263), .ZN(new_n264));
  INV_X1    g0064(.A(G190), .ZN(new_n265));
  NOR2_X1   g0065(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  NOR3_X1   g0066(.A1(G50), .A2(G58), .A3(G68), .ZN(new_n267));
  INV_X1    g0067(.A(G33), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n204), .A2(new_n268), .ZN(new_n269));
  INV_X1    g0069(.A(G150), .ZN(new_n270));
  OAI22_X1  g0070(.A1(new_n267), .A2(new_n204), .B1(new_n269), .B2(new_n270), .ZN(new_n271));
  INV_X1    g0071(.A(G58), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n272), .A2(KEYINPUT8), .ZN(new_n273));
  INV_X1    g0073(.A(KEYINPUT8), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n274), .A2(G58), .ZN(new_n275));
  NAND3_X1  g0075(.A1(new_n273), .A2(new_n275), .A3(KEYINPUT70), .ZN(new_n276));
  INV_X1    g0076(.A(new_n276), .ZN(new_n277));
  AOI21_X1  g0077(.A(KEYINPUT70), .B1(new_n273), .B2(new_n275), .ZN(new_n278));
  NOR2_X1   g0078(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  NOR2_X1   g0079(.A1(new_n268), .A2(G20), .ZN(new_n280));
  AOI21_X1  g0080(.A(new_n271), .B1(new_n279), .B2(new_n280), .ZN(new_n281));
  NAND3_X1  g0081(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n282), .A2(new_n253), .ZN(new_n283));
  INV_X1    g0083(.A(new_n283), .ZN(new_n284));
  NOR2_X1   g0084(.A1(new_n281), .A2(new_n284), .ZN(new_n285));
  NAND3_X1  g0085(.A1(new_n203), .A2(G13), .A3(G20), .ZN(new_n286));
  INV_X1    g0086(.A(new_n286), .ZN(new_n287));
  NOR2_X1   g0087(.A1(new_n287), .A2(new_n283), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n203), .A2(G20), .ZN(new_n289));
  NAND3_X1  g0089(.A1(new_n288), .A2(G50), .A3(new_n289), .ZN(new_n290));
  OAI21_X1  g0090(.A(new_n290), .B1(G50), .B2(new_n286), .ZN(new_n291));
  NOR2_X1   g0091(.A1(new_n285), .A2(new_n291), .ZN(new_n292));
  AOI21_X1  g0092(.A(new_n266), .B1(new_n292), .B2(KEYINPUT9), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n264), .A2(G200), .ZN(new_n294));
  OAI211_X1 g0094(.A(new_n293), .B(new_n294), .C1(KEYINPUT9), .C2(new_n292), .ZN(new_n295));
  XNOR2_X1  g0095(.A(new_n295), .B(KEYINPUT10), .ZN(new_n296));
  INV_X1    g0096(.A(G169), .ZN(new_n297));
  AOI21_X1  g0097(.A(new_n292), .B1(new_n297), .B2(new_n264), .ZN(new_n298));
  OAI21_X1  g0098(.A(new_n298), .B1(G179), .B2(new_n264), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n296), .A2(new_n299), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n204), .A2(G33), .ZN(new_n301));
  OAI22_X1  g0101(.A1(new_n301), .A2(new_n251), .B1(new_n204), .B2(G68), .ZN(new_n302));
  INV_X1    g0102(.A(G50), .ZN(new_n303));
  NOR2_X1   g0103(.A1(new_n269), .A2(new_n303), .ZN(new_n304));
  OAI21_X1  g0104(.A(new_n283), .B1(new_n302), .B2(new_n304), .ZN(new_n305));
  XNOR2_X1  g0105(.A(new_n305), .B(KEYINPUT11), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n286), .A2(KEYINPUT72), .ZN(new_n307));
  INV_X1    g0107(.A(KEYINPUT72), .ZN(new_n308));
  NAND4_X1  g0108(.A1(new_n308), .A2(new_n203), .A3(G13), .A4(G20), .ZN(new_n309));
  AND2_X1   g0109(.A1(new_n307), .A2(new_n309), .ZN(new_n310));
  INV_X1    g0110(.A(G68), .ZN(new_n311));
  NAND3_X1  g0111(.A1(new_n310), .A2(KEYINPUT12), .A3(new_n311), .ZN(new_n312));
  OAI211_X1 g0112(.A(new_n306), .B(new_n312), .C1(KEYINPUT12), .C2(new_n287), .ZN(new_n313));
  AOI21_X1  g0113(.A(new_n283), .B1(new_n307), .B2(new_n309), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n314), .A2(new_n289), .ZN(new_n315));
  AOI21_X1  g0115(.A(new_n311), .B1(new_n315), .B2(KEYINPUT12), .ZN(new_n316));
  NOR2_X1   g0116(.A1(new_n313), .A2(new_n316), .ZN(new_n317));
  INV_X1    g0117(.A(new_n317), .ZN(new_n318));
  NAND3_X1  g0118(.A1(new_n247), .A2(G226), .A3(new_n248), .ZN(new_n319));
  NAND3_X1  g0119(.A1(new_n247), .A2(G232), .A3(G1698), .ZN(new_n320));
  NAND2_X1  g0120(.A1(G33), .A2(G97), .ZN(new_n321));
  NAND3_X1  g0121(.A1(new_n319), .A2(new_n320), .A3(new_n321), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n322), .A2(new_n254), .ZN(new_n323));
  INV_X1    g0123(.A(new_n323), .ZN(new_n324));
  INV_X1    g0124(.A(new_n258), .ZN(new_n325));
  OAI211_X1 g0125(.A(G1), .B(G13), .C1(new_n268), .C2(new_n259), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n326), .A2(new_n256), .ZN(new_n327));
  AND2_X1   g0127(.A1(new_n327), .A2(KEYINPUT73), .ZN(new_n328));
  OAI21_X1  g0128(.A(G238), .B1(new_n327), .B2(KEYINPUT73), .ZN(new_n329));
  OAI21_X1  g0129(.A(new_n325), .B1(new_n328), .B2(new_n329), .ZN(new_n330));
  OAI21_X1  g0130(.A(KEYINPUT13), .B1(new_n324), .B2(new_n330), .ZN(new_n331));
  OR2_X1    g0131(.A1(new_n328), .A2(new_n329), .ZN(new_n332));
  INV_X1    g0132(.A(KEYINPUT13), .ZN(new_n333));
  NAND4_X1  g0133(.A1(new_n332), .A2(new_n333), .A3(new_n323), .A4(new_n325), .ZN(new_n334));
  AOI21_X1  g0134(.A(new_n297), .B1(new_n331), .B2(new_n334), .ZN(new_n335));
  INV_X1    g0135(.A(KEYINPUT14), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n331), .A2(new_n334), .ZN(new_n337));
  INV_X1    g0137(.A(G179), .ZN(new_n338));
  OAI22_X1  g0138(.A1(new_n335), .A2(new_n336), .B1(new_n337), .B2(new_n338), .ZN(new_n339));
  AND2_X1   g0139(.A1(new_n335), .A2(new_n336), .ZN(new_n340));
  OAI21_X1  g0140(.A(new_n318), .B1(new_n339), .B2(new_n340), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n337), .A2(G200), .ZN(new_n342));
  OAI211_X1 g0142(.A(new_n342), .B(new_n317), .C1(new_n265), .C2(new_n337), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n341), .A2(new_n343), .ZN(new_n344));
  INV_X1    g0144(.A(KEYINPUT3), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n345), .A2(new_n268), .ZN(new_n346));
  NAND2_X1  g0146(.A1(KEYINPUT3), .A2(G33), .ZN(new_n347));
  NAND3_X1  g0147(.A1(new_n346), .A2(new_n204), .A3(new_n347), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n348), .A2(KEYINPUT7), .ZN(new_n349));
  INV_X1    g0149(.A(KEYINPUT7), .ZN(new_n350));
  NAND4_X1  g0150(.A1(new_n346), .A2(new_n350), .A3(new_n204), .A4(new_n347), .ZN(new_n351));
  NAND3_X1  g0151(.A1(new_n349), .A2(G68), .A3(new_n351), .ZN(new_n352));
  INV_X1    g0152(.A(G159), .ZN(new_n353));
  NOR2_X1   g0153(.A1(new_n269), .A2(new_n353), .ZN(new_n354));
  XNOR2_X1  g0154(.A(G58), .B(G68), .ZN(new_n355));
  AOI21_X1  g0155(.A(new_n354), .B1(G20), .B2(new_n355), .ZN(new_n356));
  AND3_X1   g0156(.A1(new_n352), .A2(KEYINPUT16), .A3(new_n356), .ZN(new_n357));
  AOI21_X1  g0157(.A(KEYINPUT16), .B1(new_n352), .B2(new_n356), .ZN(new_n358));
  NOR3_X1   g0158(.A1(new_n357), .A2(new_n358), .A3(new_n284), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n273), .A2(new_n275), .ZN(new_n360));
  INV_X1    g0160(.A(KEYINPUT70), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  NAND4_X1  g0162(.A1(new_n288), .A2(new_n362), .A3(new_n289), .A4(new_n276), .ZN(new_n363));
  OAI21_X1  g0163(.A(new_n287), .B1(new_n277), .B2(new_n278), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n363), .A2(new_n364), .ZN(new_n365));
  INV_X1    g0165(.A(KEYINPUT74), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n365), .A2(new_n366), .ZN(new_n367));
  NAND3_X1  g0167(.A1(new_n363), .A2(new_n364), .A3(KEYINPUT74), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  NOR2_X1   g0169(.A1(new_n359), .A2(new_n369), .ZN(new_n370));
  AOI21_X1  g0170(.A(new_n258), .B1(new_n262), .B2(G232), .ZN(new_n371));
  INV_X1    g0171(.A(G223), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n372), .A2(new_n248), .ZN(new_n373));
  INV_X1    g0173(.A(G226), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n374), .A2(G1698), .ZN(new_n375));
  AND2_X1   g0175(.A1(KEYINPUT3), .A2(G33), .ZN(new_n376));
  NOR2_X1   g0176(.A1(KEYINPUT3), .A2(G33), .ZN(new_n377));
  OAI211_X1 g0177(.A(new_n373), .B(new_n375), .C1(new_n376), .C2(new_n377), .ZN(new_n378));
  NAND2_X1  g0178(.A1(G33), .A2(G87), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n378), .A2(new_n379), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n380), .A2(new_n254), .ZN(new_n381));
  NAND3_X1  g0181(.A1(new_n371), .A2(new_n381), .A3(new_n265), .ZN(new_n382));
  INV_X1    g0182(.A(G200), .ZN(new_n383));
  INV_X1    g0183(.A(G232), .ZN(new_n384));
  OAI21_X1  g0184(.A(new_n325), .B1(new_n327), .B2(new_n384), .ZN(new_n385));
  AOI21_X1  g0185(.A(new_n326), .B1(new_n378), .B2(new_n379), .ZN(new_n386));
  OAI21_X1  g0186(.A(new_n383), .B1(new_n385), .B2(new_n386), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n382), .A2(new_n387), .ZN(new_n388));
  INV_X1    g0188(.A(KEYINPUT75), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n388), .A2(new_n389), .ZN(new_n390));
  NAND3_X1  g0190(.A1(new_n382), .A2(new_n387), .A3(KEYINPUT75), .ZN(new_n391));
  NAND4_X1  g0191(.A1(new_n370), .A2(KEYINPUT17), .A3(new_n390), .A4(new_n391), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n352), .A2(new_n356), .ZN(new_n393));
  INV_X1    g0193(.A(KEYINPUT16), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n393), .A2(new_n394), .ZN(new_n395));
  NAND3_X1  g0195(.A1(new_n352), .A2(KEYINPUT16), .A3(new_n356), .ZN(new_n396));
  NAND3_X1  g0196(.A1(new_n395), .A2(new_n283), .A3(new_n396), .ZN(new_n397));
  AND3_X1   g0197(.A1(new_n363), .A2(new_n364), .A3(KEYINPUT74), .ZN(new_n398));
  AOI21_X1  g0198(.A(KEYINPUT74), .B1(new_n363), .B2(new_n364), .ZN(new_n399));
  NOR2_X1   g0199(.A1(new_n398), .A2(new_n399), .ZN(new_n400));
  NAND4_X1  g0200(.A1(new_n390), .A2(new_n397), .A3(new_n400), .A4(new_n391), .ZN(new_n401));
  INV_X1    g0201(.A(KEYINPUT17), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n401), .A2(new_n402), .ZN(new_n403));
  OAI21_X1  g0203(.A(new_n297), .B1(new_n385), .B2(new_n386), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n371), .A2(new_n381), .ZN(new_n405));
  OAI21_X1  g0205(.A(new_n404), .B1(new_n405), .B2(G179), .ZN(new_n406));
  INV_X1    g0206(.A(new_n406), .ZN(new_n407));
  OAI21_X1  g0207(.A(new_n407), .B1(new_n359), .B2(new_n369), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n408), .A2(KEYINPUT18), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n397), .A2(new_n400), .ZN(new_n410));
  INV_X1    g0210(.A(KEYINPUT18), .ZN(new_n411));
  NAND3_X1  g0211(.A1(new_n410), .A2(new_n411), .A3(new_n407), .ZN(new_n412));
  NAND4_X1  g0212(.A1(new_n392), .A2(new_n403), .A3(new_n409), .A4(new_n412), .ZN(new_n413));
  NAND3_X1  g0213(.A1(new_n247), .A2(G232), .A3(new_n248), .ZN(new_n414));
  NAND3_X1  g0214(.A1(new_n247), .A2(G238), .A3(G1698), .ZN(new_n415));
  INV_X1    g0215(.A(G107), .ZN(new_n416));
  OAI211_X1 g0216(.A(new_n414), .B(new_n415), .C1(new_n416), .C2(new_n247), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n417), .A2(new_n254), .ZN(new_n418));
  AOI21_X1  g0218(.A(new_n258), .B1(new_n262), .B2(G244), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n418), .A2(new_n419), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n420), .A2(G200), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n269), .A2(KEYINPUT71), .ZN(new_n422));
  INV_X1    g0222(.A(new_n422), .ZN(new_n423));
  XNOR2_X1  g0223(.A(KEYINPUT8), .B(G58), .ZN(new_n424));
  NOR2_X1   g0224(.A1(new_n269), .A2(KEYINPUT71), .ZN(new_n425));
  NOR3_X1   g0225(.A1(new_n423), .A2(new_n424), .A3(new_n425), .ZN(new_n426));
  XNOR2_X1  g0226(.A(KEYINPUT15), .B(G87), .ZN(new_n427));
  OAI22_X1  g0227(.A1(new_n427), .A2(new_n301), .B1(new_n204), .B2(new_n251), .ZN(new_n428));
  OAI21_X1  g0228(.A(new_n283), .B1(new_n426), .B2(new_n428), .ZN(new_n429));
  NAND3_X1  g0229(.A1(new_n314), .A2(G77), .A3(new_n289), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n310), .A2(new_n251), .ZN(new_n431));
  AND3_X1   g0231(.A1(new_n429), .A2(new_n430), .A3(new_n431), .ZN(new_n432));
  NAND3_X1  g0232(.A1(new_n418), .A2(G190), .A3(new_n419), .ZN(new_n433));
  NAND3_X1  g0233(.A1(new_n421), .A2(new_n432), .A3(new_n433), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n420), .A2(new_n297), .ZN(new_n435));
  NAND3_X1  g0235(.A1(new_n418), .A2(new_n338), .A3(new_n419), .ZN(new_n436));
  NAND3_X1  g0236(.A1(new_n429), .A2(new_n430), .A3(new_n431), .ZN(new_n437));
  NAND3_X1  g0237(.A1(new_n435), .A2(new_n436), .A3(new_n437), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n434), .A2(new_n438), .ZN(new_n439));
  NOR4_X1   g0239(.A1(new_n300), .A2(new_n344), .A3(new_n413), .A4(new_n439), .ZN(new_n440));
  INV_X1    g0240(.A(KEYINPUT21), .ZN(new_n441));
  INV_X1    g0241(.A(G116), .ZN(new_n442));
  NOR2_X1   g0242(.A1(new_n268), .A2(G1), .ZN(new_n443));
  NOR2_X1   g0243(.A1(new_n443), .A2(new_n442), .ZN(new_n444));
  AOI22_X1  g0244(.A1(new_n442), .A2(new_n310), .B1(new_n314), .B2(new_n444), .ZN(new_n445));
  INV_X1    g0245(.A(KEYINPUT81), .ZN(new_n446));
  NAND2_X1  g0246(.A1(G33), .A2(G283), .ZN(new_n447));
  INV_X1    g0247(.A(G97), .ZN(new_n448));
  OAI211_X1 g0248(.A(new_n447), .B(new_n204), .C1(G33), .C2(new_n448), .ZN(new_n449));
  INV_X1    g0249(.A(KEYINPUT80), .ZN(new_n450));
  INV_X1    g0250(.A(KEYINPUT20), .ZN(new_n451));
  AOI22_X1  g0251(.A1(new_n450), .A2(new_n451), .B1(new_n442), .B2(G20), .ZN(new_n452));
  NAND3_X1  g0252(.A1(new_n449), .A2(new_n452), .A3(new_n283), .ZN(new_n453));
  NAND2_X1  g0253(.A1(KEYINPUT80), .A2(KEYINPUT20), .ZN(new_n454));
  INV_X1    g0254(.A(new_n454), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n453), .A2(new_n455), .ZN(new_n456));
  NAND4_X1  g0256(.A1(new_n449), .A2(new_n452), .A3(new_n283), .A4(new_n454), .ZN(new_n457));
  NAND4_X1  g0257(.A1(new_n445), .A2(new_n446), .A3(new_n456), .A4(new_n457), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n314), .A2(new_n444), .ZN(new_n459));
  NAND3_X1  g0259(.A1(new_n307), .A2(new_n442), .A3(new_n309), .ZN(new_n460));
  NAND4_X1  g0260(.A1(new_n459), .A2(new_n460), .A3(new_n456), .A4(new_n457), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n461), .A2(KEYINPUT81), .ZN(new_n462));
  AND2_X1   g0262(.A1(new_n458), .A2(new_n462), .ZN(new_n463));
  NOR2_X1   g0263(.A1(new_n260), .A2(G1), .ZN(new_n464));
  AND2_X1   g0264(.A1(KEYINPUT5), .A2(G41), .ZN(new_n465));
  NOR2_X1   g0265(.A1(KEYINPUT5), .A2(G41), .ZN(new_n466));
  OAI21_X1  g0266(.A(new_n464), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  NAND3_X1  g0267(.A1(new_n467), .A2(G270), .A3(new_n326), .ZN(new_n468));
  XNOR2_X1  g0268(.A(KEYINPUT5), .B(G41), .ZN(new_n469));
  NAND4_X1  g0269(.A1(new_n469), .A2(new_n326), .A3(G274), .A4(new_n464), .ZN(new_n470));
  AND2_X1   g0270(.A1(new_n468), .A2(new_n470), .ZN(new_n471));
  OAI211_X1 g0271(.A(G264), .B(G1698), .C1(new_n376), .C2(new_n377), .ZN(new_n472));
  OAI211_X1 g0272(.A(G257), .B(new_n248), .C1(new_n376), .C2(new_n377), .ZN(new_n473));
  NAND3_X1  g0273(.A1(new_n346), .A2(G303), .A3(new_n347), .ZN(new_n474));
  NAND3_X1  g0274(.A1(new_n472), .A2(new_n473), .A3(new_n474), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n475), .A2(new_n254), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n471), .A2(new_n476), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n477), .A2(G169), .ZN(new_n478));
  OAI21_X1  g0278(.A(new_n441), .B1(new_n463), .B2(new_n478), .ZN(new_n479));
  NAND3_X1  g0279(.A1(new_n471), .A2(G179), .A3(new_n476), .ZN(new_n480));
  AOI21_X1  g0280(.A(new_n480), .B1(new_n458), .B2(new_n462), .ZN(new_n481));
  AOI21_X1  g0281(.A(new_n478), .B1(new_n458), .B2(new_n462), .ZN(new_n482));
  AOI21_X1  g0282(.A(new_n481), .B1(new_n482), .B2(KEYINPUT21), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n203), .A2(G33), .ZN(new_n484));
  NAND4_X1  g0284(.A1(new_n286), .A2(new_n484), .A3(new_n253), .A4(new_n282), .ZN(new_n485));
  INV_X1    g0285(.A(KEYINPUT78), .ZN(new_n486));
  OR3_X1    g0286(.A1(new_n485), .A2(new_n486), .A3(new_n427), .ZN(new_n487));
  OAI21_X1  g0287(.A(new_n486), .B1(new_n485), .B2(new_n427), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  INV_X1    g0289(.A(KEYINPUT19), .ZN(new_n490));
  OAI21_X1  g0290(.A(new_n204), .B1(new_n321), .B2(new_n490), .ZN(new_n491));
  NOR2_X1   g0291(.A1(G97), .A2(G107), .ZN(new_n492));
  INV_X1    g0292(.A(G87), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n491), .A2(new_n494), .ZN(new_n495));
  OAI211_X1 g0295(.A(new_n204), .B(G68), .C1(new_n376), .C2(new_n377), .ZN(new_n496));
  OAI21_X1  g0296(.A(new_n490), .B1(new_n301), .B2(new_n448), .ZN(new_n497));
  NAND3_X1  g0297(.A1(new_n495), .A2(new_n496), .A3(new_n497), .ZN(new_n498));
  AOI22_X1  g0298(.A1(new_n498), .A2(new_n283), .B1(new_n310), .B2(new_n427), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n489), .A2(new_n499), .ZN(new_n500));
  INV_X1    g0300(.A(KEYINPUT79), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  NAND3_X1  g0302(.A1(new_n489), .A2(new_n499), .A3(KEYINPUT79), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  OAI211_X1 g0304(.A(G238), .B(new_n248), .C1(new_n376), .C2(new_n377), .ZN(new_n505));
  OAI211_X1 g0305(.A(G244), .B(G1698), .C1(new_n376), .C2(new_n377), .ZN(new_n506));
  OAI211_X1 g0306(.A(new_n505), .B(new_n506), .C1(new_n268), .C2(new_n442), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n507), .A2(new_n254), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n203), .A2(G45), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n509), .A2(G250), .ZN(new_n510));
  OAI22_X1  g0310(.A1(new_n254), .A2(new_n510), .B1(new_n257), .B2(new_n509), .ZN(new_n511));
  INV_X1    g0311(.A(new_n511), .ZN(new_n512));
  AOI21_X1  g0312(.A(G169), .B1(new_n508), .B2(new_n512), .ZN(new_n513));
  AOI211_X1 g0313(.A(G179), .B(new_n511), .C1(new_n507), .C2(new_n254), .ZN(new_n514));
  NOR2_X1   g0314(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  AOI21_X1  g0315(.A(new_n511), .B1(new_n507), .B2(new_n254), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n516), .A2(G190), .ZN(new_n517));
  AOI21_X1  g0317(.A(new_n383), .B1(new_n508), .B2(new_n512), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n498), .A2(new_n283), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n310), .A2(new_n427), .ZN(new_n520));
  INV_X1    g0320(.A(new_n485), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n521), .A2(G87), .ZN(new_n522));
  NAND3_X1  g0322(.A1(new_n519), .A2(new_n520), .A3(new_n522), .ZN(new_n523));
  NOR2_X1   g0323(.A1(new_n518), .A2(new_n523), .ZN(new_n524));
  AOI22_X1  g0324(.A1(new_n504), .A2(new_n515), .B1(new_n517), .B2(new_n524), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n477), .A2(G200), .ZN(new_n526));
  OAI211_X1 g0326(.A(new_n463), .B(new_n526), .C1(new_n265), .C2(new_n477), .ZN(new_n527));
  AND4_X1   g0327(.A1(new_n479), .A2(new_n483), .A3(new_n525), .A4(new_n527), .ZN(new_n528));
  NAND3_X1  g0328(.A1(new_n247), .A2(new_n204), .A3(G87), .ZN(new_n529));
  XNOR2_X1  g0329(.A(KEYINPUT82), .B(KEYINPUT22), .ZN(new_n530));
  INV_X1    g0330(.A(new_n530), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n529), .A2(new_n531), .ZN(new_n532));
  NAND4_X1  g0332(.A1(new_n247), .A2(new_n530), .A3(new_n204), .A4(G87), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  INV_X1    g0334(.A(KEYINPUT24), .ZN(new_n535));
  NOR3_X1   g0335(.A1(new_n268), .A2(new_n442), .A3(G20), .ZN(new_n536));
  INV_X1    g0336(.A(KEYINPUT23), .ZN(new_n537));
  OAI21_X1  g0337(.A(new_n537), .B1(new_n204), .B2(G107), .ZN(new_n538));
  NAND3_X1  g0338(.A1(new_n416), .A2(KEYINPUT23), .A3(G20), .ZN(new_n539));
  AOI21_X1  g0339(.A(new_n536), .B1(new_n538), .B2(new_n539), .ZN(new_n540));
  AND3_X1   g0340(.A1(new_n534), .A2(new_n535), .A3(new_n540), .ZN(new_n541));
  AOI21_X1  g0341(.A(new_n535), .B1(new_n534), .B2(new_n540), .ZN(new_n542));
  OAI21_X1  g0342(.A(new_n283), .B1(new_n541), .B2(new_n542), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n287), .A2(new_n416), .ZN(new_n544));
  INV_X1    g0344(.A(KEYINPUT25), .ZN(new_n545));
  NOR2_X1   g0345(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  XNOR2_X1  g0346(.A(new_n546), .B(KEYINPUT83), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n544), .A2(new_n545), .ZN(new_n548));
  XNOR2_X1  g0348(.A(new_n548), .B(KEYINPUT84), .ZN(new_n549));
  AOI22_X1  g0349(.A1(new_n547), .A2(new_n549), .B1(G107), .B2(new_n521), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n543), .A2(new_n550), .ZN(new_n551));
  INV_X1    g0351(.A(KEYINPUT85), .ZN(new_n552));
  OAI211_X1 g0352(.A(G250), .B(new_n248), .C1(new_n376), .C2(new_n377), .ZN(new_n553));
  OAI211_X1 g0353(.A(G257), .B(G1698), .C1(new_n376), .C2(new_n377), .ZN(new_n554));
  INV_X1    g0354(.A(G294), .ZN(new_n555));
  OAI211_X1 g0355(.A(new_n553), .B(new_n554), .C1(new_n268), .C2(new_n555), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n556), .A2(new_n254), .ZN(new_n557));
  AOI21_X1  g0357(.A(new_n254), .B1(new_n464), .B2(new_n469), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n558), .A2(G264), .ZN(new_n559));
  NAND3_X1  g0359(.A1(new_n557), .A2(new_n470), .A3(new_n559), .ZN(new_n560));
  AOI21_X1  g0360(.A(new_n552), .B1(new_n560), .B2(G169), .ZN(new_n561));
  NOR2_X1   g0361(.A1(new_n560), .A2(new_n338), .ZN(new_n562));
  NOR2_X1   g0362(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  NOR3_X1   g0363(.A1(new_n560), .A2(new_n552), .A3(new_n338), .ZN(new_n564));
  OAI21_X1  g0364(.A(new_n551), .B1(new_n563), .B2(new_n564), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n560), .A2(new_n383), .ZN(new_n566));
  OAI21_X1  g0366(.A(new_n566), .B1(G190), .B2(new_n560), .ZN(new_n567));
  NAND3_X1  g0367(.A1(new_n567), .A2(new_n543), .A3(new_n550), .ZN(new_n568));
  AND2_X1   g0368(.A1(new_n565), .A2(new_n568), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n287), .A2(new_n448), .ZN(new_n570));
  OAI21_X1  g0370(.A(new_n570), .B1(new_n485), .B2(new_n448), .ZN(new_n571));
  NOR2_X1   g0371(.A1(new_n269), .A2(new_n251), .ZN(new_n572));
  INV_X1    g0372(.A(KEYINPUT6), .ZN(new_n573));
  AND2_X1   g0373(.A1(G97), .A2(G107), .ZN(new_n574));
  OAI21_X1  g0374(.A(new_n573), .B1(new_n574), .B2(new_n492), .ZN(new_n575));
  NAND3_X1  g0375(.A1(new_n416), .A2(KEYINPUT6), .A3(G97), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  AOI21_X1  g0377(.A(new_n572), .B1(new_n577), .B2(G20), .ZN(new_n578));
  NAND3_X1  g0378(.A1(new_n349), .A2(G107), .A3(new_n351), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n580), .A2(new_n283), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n581), .A2(KEYINPUT76), .ZN(new_n582));
  INV_X1    g0382(.A(KEYINPUT76), .ZN(new_n583));
  NAND3_X1  g0383(.A1(new_n580), .A2(new_n583), .A3(new_n283), .ZN(new_n584));
  AOI21_X1  g0384(.A(new_n571), .B1(new_n582), .B2(new_n584), .ZN(new_n585));
  NAND3_X1  g0385(.A1(new_n467), .A2(G257), .A3(new_n326), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n586), .A2(new_n470), .ZN(new_n587));
  OAI211_X1 g0387(.A(G244), .B(new_n248), .C1(new_n376), .C2(new_n377), .ZN(new_n588));
  INV_X1    g0388(.A(KEYINPUT4), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  NAND4_X1  g0390(.A1(new_n247), .A2(KEYINPUT4), .A3(G244), .A4(new_n248), .ZN(new_n591));
  NAND3_X1  g0391(.A1(new_n247), .A2(G250), .A3(G1698), .ZN(new_n592));
  NAND4_X1  g0392(.A1(new_n590), .A2(new_n591), .A3(new_n447), .A4(new_n592), .ZN(new_n593));
  AOI21_X1  g0393(.A(new_n587), .B1(new_n593), .B2(new_n254), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n594), .A2(new_n338), .ZN(new_n595));
  OAI21_X1  g0395(.A(new_n595), .B1(G169), .B2(new_n594), .ZN(new_n596));
  NOR2_X1   g0396(.A1(new_n585), .A2(new_n596), .ZN(new_n597));
  AOI211_X1 g0397(.A(G190), .B(new_n587), .C1(new_n593), .C2(new_n254), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n593), .A2(new_n254), .ZN(new_n599));
  INV_X1    g0399(.A(new_n587), .ZN(new_n600));
  AOI21_X1  g0400(.A(G200), .B1(new_n599), .B2(new_n600), .ZN(new_n601));
  NOR2_X1   g0401(.A1(new_n598), .A2(new_n601), .ZN(new_n602));
  INV_X1    g0402(.A(new_n571), .ZN(new_n603));
  AOI21_X1  g0403(.A(new_n583), .B1(new_n580), .B2(new_n283), .ZN(new_n604));
  AOI211_X1 g0404(.A(KEYINPUT76), .B(new_n284), .C1(new_n578), .C2(new_n579), .ZN(new_n605));
  OAI21_X1  g0405(.A(new_n603), .B1(new_n604), .B2(new_n605), .ZN(new_n606));
  NOR2_X1   g0406(.A1(new_n602), .A2(new_n606), .ZN(new_n607));
  OAI21_X1  g0407(.A(KEYINPUT77), .B1(new_n597), .B2(new_n607), .ZN(new_n608));
  OAI221_X1 g0408(.A(new_n603), .B1(new_n604), .B2(new_n605), .C1(new_n598), .C2(new_n601), .ZN(new_n609));
  NOR2_X1   g0409(.A1(new_n594), .A2(G169), .ZN(new_n610));
  AOI211_X1 g0410(.A(G179), .B(new_n587), .C1(new_n593), .C2(new_n254), .ZN(new_n611));
  NOR2_X1   g0411(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n612), .A2(new_n606), .ZN(new_n613));
  INV_X1    g0413(.A(KEYINPUT77), .ZN(new_n614));
  NAND3_X1  g0414(.A1(new_n609), .A2(new_n613), .A3(new_n614), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n608), .A2(new_n615), .ZN(new_n616));
  AND4_X1   g0416(.A1(new_n440), .A2(new_n528), .A3(new_n569), .A4(new_n616), .ZN(G372));
  INV_X1    g0417(.A(new_n299), .ZN(new_n618));
  INV_X1    g0418(.A(new_n296), .ZN(new_n619));
  INV_X1    g0419(.A(KEYINPUT88), .ZN(new_n620));
  AOI211_X1 g0420(.A(KEYINPUT18), .B(new_n406), .C1(new_n397), .C2(new_n400), .ZN(new_n621));
  AOI21_X1  g0421(.A(new_n411), .B1(new_n410), .B2(new_n407), .ZN(new_n622));
  OAI21_X1  g0422(.A(new_n620), .B1(new_n621), .B2(new_n622), .ZN(new_n623));
  NAND3_X1  g0423(.A1(new_n409), .A2(KEYINPUT88), .A3(new_n412), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  INV_X1    g0425(.A(new_n438), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n343), .A2(new_n626), .ZN(new_n627));
  AND2_X1   g0427(.A1(new_n341), .A2(new_n627), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n392), .A2(new_n403), .ZN(new_n629));
  OAI21_X1  g0429(.A(new_n625), .B1(new_n628), .B2(new_n629), .ZN(new_n630));
  INV_X1    g0430(.A(KEYINPUT89), .ZN(new_n631));
  AOI21_X1  g0431(.A(new_n619), .B1(new_n630), .B2(new_n631), .ZN(new_n632));
  OAI211_X1 g0432(.A(KEYINPUT89), .B(new_n625), .C1(new_n628), .C2(new_n629), .ZN(new_n633));
  AOI21_X1  g0433(.A(new_n618), .B1(new_n632), .B2(new_n633), .ZN(new_n634));
  INV_X1    g0434(.A(new_n503), .ZN(new_n635));
  AOI21_X1  g0435(.A(KEYINPUT79), .B1(new_n489), .B2(new_n499), .ZN(new_n636));
  OAI21_X1  g0436(.A(new_n515), .B1(new_n635), .B2(new_n636), .ZN(new_n637));
  INV_X1    g0437(.A(new_n637), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n508), .A2(new_n512), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n639), .A2(G200), .ZN(new_n640));
  INV_X1    g0440(.A(KEYINPUT86), .ZN(new_n641));
  INV_X1    g0441(.A(new_n523), .ZN(new_n642));
  NAND3_X1  g0442(.A1(new_n640), .A2(new_n641), .A3(new_n642), .ZN(new_n643));
  OAI21_X1  g0443(.A(KEYINPUT86), .B1(new_n518), .B2(new_n523), .ZN(new_n644));
  NAND3_X1  g0444(.A1(new_n643), .A2(new_n517), .A3(new_n644), .ZN(new_n645));
  AND4_X1   g0445(.A1(new_n568), .A2(new_n609), .A3(new_n613), .A4(new_n645), .ZN(new_n646));
  NAND3_X1  g0446(.A1(new_n565), .A2(new_n479), .A3(new_n483), .ZN(new_n647));
  AOI21_X1  g0447(.A(new_n638), .B1(new_n646), .B2(new_n647), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n524), .A2(new_n517), .ZN(new_n649));
  NAND4_X1  g0449(.A1(new_n637), .A2(new_n612), .A3(new_n649), .A4(new_n606), .ZN(new_n650));
  INV_X1    g0450(.A(KEYINPUT26), .ZN(new_n651));
  OAI21_X1  g0451(.A(KEYINPUT87), .B1(new_n650), .B2(new_n651), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n645), .A2(new_n637), .ZN(new_n653));
  OAI21_X1  g0453(.A(new_n651), .B1(new_n653), .B2(new_n613), .ZN(new_n654));
  INV_X1    g0454(.A(KEYINPUT87), .ZN(new_n655));
  NAND4_X1  g0455(.A1(new_n597), .A2(new_n525), .A3(new_n655), .A4(KEYINPUT26), .ZN(new_n656));
  NAND3_X1  g0456(.A1(new_n652), .A2(new_n654), .A3(new_n656), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n648), .A2(new_n657), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n440), .A2(new_n658), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n634), .A2(new_n659), .ZN(G369));
  NAND3_X1  g0460(.A1(new_n203), .A2(new_n204), .A3(G13), .ZN(new_n661));
  OR2_X1    g0461(.A1(new_n661), .A2(KEYINPUT27), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n661), .A2(KEYINPUT27), .ZN(new_n663));
  NAND3_X1  g0463(.A1(new_n662), .A2(G213), .A3(new_n663), .ZN(new_n664));
  INV_X1    g0464(.A(G343), .ZN(new_n665));
  NOR2_X1   g0465(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  INV_X1    g0466(.A(new_n666), .ZN(new_n667));
  AOI21_X1  g0467(.A(new_n667), .B1(new_n543), .B2(new_n550), .ZN(new_n668));
  XNOR2_X1  g0468(.A(new_n668), .B(KEYINPUT91), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n669), .A2(new_n569), .ZN(new_n670));
  OAI21_X1  g0470(.A(new_n670), .B1(new_n565), .B2(new_n667), .ZN(new_n671));
  XOR2_X1   g0471(.A(KEYINPUT90), .B(G330), .Z(new_n672));
  NAND2_X1  g0472(.A1(new_n483), .A2(new_n479), .ZN(new_n673));
  NOR2_X1   g0473(.A1(new_n463), .A2(new_n667), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  INV_X1    g0475(.A(new_n674), .ZN(new_n676));
  NAND4_X1  g0476(.A1(new_n676), .A2(new_n483), .A3(new_n479), .A4(new_n527), .ZN(new_n677));
  AOI21_X1  g0477(.A(new_n672), .B1(new_n675), .B2(new_n677), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n671), .A2(new_n678), .ZN(new_n679));
  OR2_X1    g0479(.A1(new_n565), .A2(new_n666), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n673), .A2(new_n667), .ZN(new_n681));
  INV_X1    g0481(.A(new_n681), .ZN(new_n682));
  NAND3_X1  g0482(.A1(new_n682), .A2(new_n569), .A3(new_n669), .ZN(new_n683));
  NAND3_X1  g0483(.A1(new_n679), .A2(new_n680), .A3(new_n683), .ZN(G399));
  INV_X1    g0484(.A(new_n222), .ZN(new_n685));
  NOR2_X1   g0485(.A1(new_n685), .A2(G41), .ZN(new_n686));
  INV_X1    g0486(.A(new_n686), .ZN(new_n687));
  NOR2_X1   g0487(.A1(new_n494), .A2(G116), .ZN(new_n688));
  NAND3_X1  g0488(.A1(new_n687), .A2(G1), .A3(new_n688), .ZN(new_n689));
  OAI21_X1  g0489(.A(new_n689), .B1(new_n226), .B2(new_n687), .ZN(new_n690));
  XNOR2_X1  g0490(.A(new_n690), .B(KEYINPUT28), .ZN(new_n691));
  AOI21_X1  g0491(.A(new_n666), .B1(new_n648), .B2(new_n657), .ZN(new_n692));
  INV_X1    g0492(.A(KEYINPUT29), .ZN(new_n693));
  AND2_X1   g0493(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n650), .A2(new_n651), .ZN(new_n695));
  INV_X1    g0495(.A(KEYINPUT93), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  NAND4_X1  g0497(.A1(new_n597), .A2(KEYINPUT26), .A3(new_n637), .A4(new_n645), .ZN(new_n698));
  NAND3_X1  g0498(.A1(new_n650), .A2(KEYINPUT93), .A3(new_n651), .ZN(new_n699));
  NAND3_X1  g0499(.A1(new_n697), .A2(new_n698), .A3(new_n699), .ZN(new_n700));
  AOI21_X1  g0500(.A(new_n666), .B1(new_n700), .B2(new_n648), .ZN(new_n701));
  NOR2_X1   g0501(.A1(new_n701), .A2(new_n693), .ZN(new_n702));
  NAND4_X1  g0502(.A1(new_n616), .A2(new_n528), .A3(new_n569), .A4(new_n667), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n480), .A2(KEYINPUT92), .ZN(new_n704));
  AOI22_X1  g0504(.A1(new_n556), .A2(new_n254), .B1(new_n558), .B2(G264), .ZN(new_n705));
  AND2_X1   g0505(.A1(new_n705), .A2(new_n516), .ZN(new_n706));
  INV_X1    g0506(.A(KEYINPUT92), .ZN(new_n707));
  NAND4_X1  g0507(.A1(new_n471), .A2(new_n707), .A3(new_n476), .A4(G179), .ZN(new_n708));
  NAND4_X1  g0508(.A1(new_n704), .A2(new_n706), .A3(new_n594), .A4(new_n708), .ZN(new_n709));
  INV_X1    g0509(.A(KEYINPUT30), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  AND3_X1   g0511(.A1(new_n594), .A2(new_n516), .A3(new_n705), .ZN(new_n712));
  NAND4_X1  g0512(.A1(new_n712), .A2(KEYINPUT30), .A3(new_n708), .A4(new_n704), .ZN(new_n713));
  AOI21_X1  g0513(.A(new_n594), .B1(new_n470), .B2(new_n705), .ZN(new_n714));
  NAND4_X1  g0514(.A1(new_n714), .A2(new_n338), .A3(new_n477), .A4(new_n639), .ZN(new_n715));
  NAND3_X1  g0515(.A1(new_n711), .A2(new_n713), .A3(new_n715), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n716), .A2(new_n666), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n717), .A2(KEYINPUT31), .ZN(new_n718));
  INV_X1    g0518(.A(KEYINPUT31), .ZN(new_n719));
  NAND3_X1  g0519(.A1(new_n716), .A2(new_n719), .A3(new_n666), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n718), .A2(new_n720), .ZN(new_n721));
  AOI21_X1  g0521(.A(new_n672), .B1(new_n703), .B2(new_n721), .ZN(new_n722));
  NOR3_X1   g0522(.A1(new_n694), .A2(new_n702), .A3(new_n722), .ZN(new_n723));
  OAI21_X1  g0523(.A(new_n691), .B1(new_n723), .B2(G1), .ZN(G364));
  INV_X1    g0524(.A(G13), .ZN(new_n725));
  NOR3_X1   g0525(.A1(new_n725), .A2(new_n260), .A3(G20), .ZN(new_n726));
  OR2_X1    g0526(.A1(new_n726), .A2(KEYINPUT94), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n726), .A2(KEYINPUT94), .ZN(new_n728));
  NAND3_X1  g0528(.A1(new_n727), .A2(G1), .A3(new_n728), .ZN(new_n729));
  OR3_X1    g0529(.A1(new_n686), .A2(new_n729), .A3(KEYINPUT95), .ZN(new_n730));
  OAI21_X1  g0530(.A(KEYINPUT95), .B1(new_n686), .B2(new_n729), .ZN(new_n731));
  NAND2_X1  g0531(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  INV_X1    g0532(.A(new_n732), .ZN(new_n733));
  NAND2_X1  g0533(.A1(new_n245), .A2(G45), .ZN(new_n734));
  NOR2_X1   g0534(.A1(new_n685), .A2(new_n247), .ZN(new_n735));
  OAI211_X1 g0535(.A(new_n734), .B(new_n735), .C1(G45), .C2(new_n226), .ZN(new_n736));
  INV_X1    g0536(.A(new_n247), .ZN(new_n737));
  NOR2_X1   g0537(.A1(new_n685), .A2(new_n737), .ZN(new_n738));
  XNOR2_X1  g0538(.A(G355), .B(KEYINPUT96), .ZN(new_n739));
  AOI22_X1  g0539(.A1(new_n738), .A2(new_n739), .B1(new_n442), .B2(new_n685), .ZN(new_n740));
  AND2_X1   g0540(.A1(new_n736), .A2(new_n740), .ZN(new_n741));
  NOR2_X1   g0541(.A1(G13), .A2(G33), .ZN(new_n742));
  INV_X1    g0542(.A(new_n742), .ZN(new_n743));
  NOR2_X1   g0543(.A1(new_n743), .A2(G20), .ZN(new_n744));
  XOR2_X1   g0544(.A(new_n744), .B(KEYINPUT97), .Z(new_n745));
  INV_X1    g0545(.A(new_n745), .ZN(new_n746));
  NOR2_X1   g0546(.A1(new_n297), .A2(KEYINPUT98), .ZN(new_n747));
  INV_X1    g0547(.A(new_n747), .ZN(new_n748));
  AOI21_X1  g0548(.A(new_n204), .B1(KEYINPUT98), .B2(new_n297), .ZN(new_n749));
  AOI21_X1  g0549(.A(new_n253), .B1(new_n748), .B2(new_n749), .ZN(new_n750));
  NOR2_X1   g0550(.A1(new_n746), .A2(new_n750), .ZN(new_n751));
  INV_X1    g0551(.A(new_n751), .ZN(new_n752));
  OAI21_X1  g0552(.A(new_n733), .B1(new_n741), .B2(new_n752), .ZN(new_n753));
  NOR2_X1   g0553(.A1(new_n204), .A2(G190), .ZN(new_n754));
  NOR2_X1   g0554(.A1(G179), .A2(G200), .ZN(new_n755));
  XNOR2_X1  g0555(.A(new_n755), .B(KEYINPUT100), .ZN(new_n756));
  AOI21_X1  g0556(.A(new_n754), .B1(new_n756), .B2(G20), .ZN(new_n757));
  XNOR2_X1  g0557(.A(new_n757), .B(KEYINPUT101), .ZN(new_n758));
  OR2_X1    g0558(.A1(new_n758), .A2(KEYINPUT102), .ZN(new_n759));
  NAND2_X1  g0559(.A1(new_n758), .A2(KEYINPUT102), .ZN(new_n760));
  NAND2_X1  g0560(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  INV_X1    g0561(.A(new_n761), .ZN(new_n762));
  NAND2_X1  g0562(.A1(new_n762), .A2(G97), .ZN(new_n763));
  INV_X1    g0563(.A(new_n754), .ZN(new_n764));
  NOR2_X1   g0564(.A1(new_n756), .A2(new_n764), .ZN(new_n765));
  NAND2_X1  g0565(.A1(new_n765), .A2(G159), .ZN(new_n766));
  XOR2_X1   g0566(.A(new_n766), .B(KEYINPUT32), .Z(new_n767));
  NOR3_X1   g0567(.A1(new_n764), .A2(new_n338), .A3(new_n383), .ZN(new_n768));
  NOR2_X1   g0568(.A1(new_n204), .A2(new_n265), .ZN(new_n769));
  NOR2_X1   g0569(.A1(new_n338), .A2(G200), .ZN(new_n770));
  NAND2_X1  g0570(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  INV_X1    g0571(.A(new_n771), .ZN(new_n772));
  AOI22_X1  g0572(.A1(new_n768), .A2(G68), .B1(new_n772), .B2(G58), .ZN(new_n773));
  NOR2_X1   g0573(.A1(new_n383), .A2(G179), .ZN(new_n774));
  NAND2_X1  g0574(.A1(new_n769), .A2(new_n774), .ZN(new_n775));
  INV_X1    g0575(.A(new_n775), .ZN(new_n776));
  NAND2_X1  g0576(.A1(new_n754), .A2(new_n770), .ZN(new_n777));
  INV_X1    g0577(.A(new_n777), .ZN(new_n778));
  AOI22_X1  g0578(.A1(G87), .A2(new_n776), .B1(new_n778), .B2(G77), .ZN(new_n779));
  NAND2_X1  g0579(.A1(new_n754), .A2(new_n774), .ZN(new_n780));
  INV_X1    g0580(.A(new_n780), .ZN(new_n781));
  AOI21_X1  g0581(.A(new_n737), .B1(new_n781), .B2(G107), .ZN(new_n782));
  NAND3_X1  g0582(.A1(new_n773), .A2(new_n779), .A3(new_n782), .ZN(new_n783));
  NAND3_X1  g0583(.A1(new_n769), .A2(G179), .A3(G200), .ZN(new_n784));
  NAND2_X1  g0584(.A1(new_n784), .A2(KEYINPUT99), .ZN(new_n785));
  INV_X1    g0585(.A(new_n785), .ZN(new_n786));
  NOR2_X1   g0586(.A1(new_n784), .A2(KEYINPUT99), .ZN(new_n787));
  OR2_X1    g0587(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  AOI21_X1  g0588(.A(new_n783), .B1(G50), .B2(new_n788), .ZN(new_n789));
  NAND3_X1  g0589(.A1(new_n763), .A2(new_n767), .A3(new_n789), .ZN(new_n790));
  XNOR2_X1  g0590(.A(new_n790), .B(KEYINPUT103), .ZN(new_n791));
  AOI22_X1  g0591(.A1(G283), .A2(new_n781), .B1(new_n778), .B2(G311), .ZN(new_n792));
  INV_X1    g0592(.A(G303), .ZN(new_n793));
  INV_X1    g0593(.A(new_n768), .ZN(new_n794));
  XOR2_X1   g0594(.A(KEYINPUT33), .B(G317), .Z(new_n795));
  OAI221_X1 g0595(.A(new_n792), .B1(new_n793), .B2(new_n775), .C1(new_n794), .C2(new_n795), .ZN(new_n796));
  AOI211_X1 g0596(.A(new_n247), .B(new_n796), .C1(G322), .C2(new_n772), .ZN(new_n797));
  AOI22_X1  g0597(.A1(new_n788), .A2(G326), .B1(new_n765), .B2(G329), .ZN(new_n798));
  INV_X1    g0598(.A(new_n758), .ZN(new_n799));
  OAI211_X1 g0599(.A(new_n797), .B(new_n798), .C1(new_n799), .C2(new_n555), .ZN(new_n800));
  AOI21_X1  g0600(.A(KEYINPUT104), .B1(new_n791), .B2(new_n800), .ZN(new_n801));
  INV_X1    g0601(.A(new_n750), .ZN(new_n802));
  NOR2_X1   g0602(.A1(new_n801), .A2(new_n802), .ZN(new_n803));
  NAND3_X1  g0603(.A1(new_n791), .A2(KEYINPUT104), .A3(new_n800), .ZN(new_n804));
  AOI21_X1  g0604(.A(new_n753), .B1(new_n803), .B2(new_n804), .ZN(new_n805));
  NAND3_X1  g0605(.A1(new_n675), .A2(new_n677), .A3(new_n746), .ZN(new_n806));
  NAND2_X1  g0606(.A1(new_n805), .A2(new_n806), .ZN(new_n807));
  NOR2_X1   g0607(.A1(new_n678), .A2(new_n733), .ZN(new_n808));
  NAND3_X1  g0608(.A1(new_n675), .A2(new_n672), .A3(new_n677), .ZN(new_n809));
  NAND2_X1  g0609(.A1(new_n808), .A2(new_n809), .ZN(new_n810));
  AND2_X1   g0610(.A1(new_n807), .A2(new_n810), .ZN(new_n811));
  INV_X1    g0611(.A(new_n811), .ZN(G396));
  NAND2_X1  g0612(.A1(new_n802), .A2(new_n743), .ZN(new_n813));
  OAI21_X1  g0613(.A(new_n733), .B1(G77), .B2(new_n813), .ZN(new_n814));
  XOR2_X1   g0614(.A(new_n814), .B(KEYINPUT105), .Z(new_n815));
  OAI211_X1 g0615(.A(new_n434), .B(new_n438), .C1(new_n432), .C2(new_n667), .ZN(new_n816));
  XNOR2_X1  g0616(.A(new_n816), .B(KEYINPUT107), .ZN(new_n817));
  OAI21_X1  g0617(.A(new_n817), .B1(new_n438), .B2(new_n667), .ZN(new_n818));
  AOI22_X1  g0618(.A1(new_n768), .A2(G283), .B1(new_n772), .B2(G294), .ZN(new_n819));
  NAND2_X1  g0619(.A1(new_n781), .A2(G87), .ZN(new_n820));
  NAND2_X1  g0620(.A1(new_n778), .A2(G116), .ZN(new_n821));
  NAND3_X1  g0621(.A1(new_n819), .A2(new_n820), .A3(new_n821), .ZN(new_n822));
  AOI211_X1 g0622(.A(new_n247), .B(new_n822), .C1(G107), .C2(new_n776), .ZN(new_n823));
  AOI22_X1  g0623(.A1(new_n788), .A2(G303), .B1(new_n765), .B2(G311), .ZN(new_n824));
  NAND3_X1  g0624(.A1(new_n763), .A2(new_n823), .A3(new_n824), .ZN(new_n825));
  OR2_X1    g0625(.A1(new_n825), .A2(KEYINPUT106), .ZN(new_n826));
  NAND2_X1  g0626(.A1(new_n825), .A2(KEYINPUT106), .ZN(new_n827));
  INV_X1    g0627(.A(new_n765), .ZN(new_n828));
  INV_X1    g0628(.A(G132), .ZN(new_n829));
  NOR2_X1   g0629(.A1(new_n828), .A2(new_n829), .ZN(new_n830));
  NAND2_X1  g0630(.A1(new_n781), .A2(G68), .ZN(new_n831));
  OAI211_X1 g0631(.A(new_n831), .B(new_n247), .C1(new_n303), .C2(new_n775), .ZN(new_n832));
  AOI22_X1  g0632(.A1(G143), .A2(new_n772), .B1(new_n778), .B2(G159), .ZN(new_n833));
  INV_X1    g0633(.A(new_n788), .ZN(new_n834));
  INV_X1    g0634(.A(G137), .ZN(new_n835));
  OAI221_X1 g0635(.A(new_n833), .B1(new_n270), .B2(new_n794), .C1(new_n834), .C2(new_n835), .ZN(new_n836));
  INV_X1    g0636(.A(KEYINPUT34), .ZN(new_n837));
  AOI211_X1 g0637(.A(new_n830), .B(new_n832), .C1(new_n836), .C2(new_n837), .ZN(new_n838));
  OAI221_X1 g0638(.A(new_n838), .B1(new_n837), .B2(new_n836), .C1(new_n272), .C2(new_n799), .ZN(new_n839));
  AND3_X1   g0639(.A1(new_n826), .A2(new_n827), .A3(new_n839), .ZN(new_n840));
  OAI221_X1 g0640(.A(new_n815), .B1(new_n743), .B2(new_n818), .C1(new_n840), .C2(new_n802), .ZN(new_n841));
  INV_X1    g0641(.A(new_n722), .ZN(new_n842));
  NOR2_X1   g0642(.A1(new_n692), .A2(new_n818), .ZN(new_n843));
  AOI211_X1 g0643(.A(new_n666), .B(new_n817), .C1(new_n648), .C2(new_n657), .ZN(new_n844));
  OAI21_X1  g0644(.A(new_n842), .B1(new_n843), .B2(new_n844), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n845), .A2(new_n732), .ZN(new_n846));
  NOR3_X1   g0646(.A1(new_n842), .A2(new_n843), .A3(new_n844), .ZN(new_n847));
  OAI21_X1  g0647(.A(new_n841), .B1(new_n846), .B2(new_n847), .ZN(new_n848));
  XOR2_X1   g0648(.A(new_n848), .B(KEYINPUT108), .Z(new_n849));
  INV_X1    g0649(.A(new_n849), .ZN(G384));
  NAND2_X1  g0650(.A1(new_n703), .A2(new_n721), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n318), .A2(new_n666), .ZN(new_n852));
  NAND3_X1  g0652(.A1(new_n341), .A2(new_n343), .A3(new_n852), .ZN(new_n853));
  OAI211_X1 g0653(.A(new_n318), .B(new_n666), .C1(new_n339), .C2(new_n340), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  NAND3_X1  g0655(.A1(new_n851), .A2(new_n818), .A3(new_n855), .ZN(new_n856));
  INV_X1    g0656(.A(new_n856), .ZN(new_n857));
  NOR2_X1   g0657(.A1(new_n370), .A2(new_n664), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n413), .A2(new_n858), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n401), .A2(new_n408), .ZN(new_n860));
  OAI21_X1  g0660(.A(KEYINPUT37), .B1(new_n860), .B2(new_n858), .ZN(new_n861));
  XOR2_X1   g0661(.A(new_n664), .B(KEYINPUT111), .Z(new_n862));
  OAI21_X1  g0662(.A(new_n862), .B1(new_n359), .B2(new_n369), .ZN(new_n863));
  INV_X1    g0663(.A(KEYINPUT37), .ZN(new_n864));
  NAND4_X1  g0664(.A1(new_n401), .A2(new_n408), .A3(new_n863), .A4(new_n864), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n861), .A2(new_n865), .ZN(new_n866));
  NAND3_X1  g0666(.A1(new_n859), .A2(new_n866), .A3(KEYINPUT38), .ZN(new_n867));
  INV_X1    g0667(.A(new_n867), .ZN(new_n868));
  AOI21_X1  g0668(.A(KEYINPUT38), .B1(new_n859), .B2(new_n866), .ZN(new_n869));
  OR2_X1    g0669(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  AOI21_X1  g0670(.A(KEYINPUT40), .B1(new_n857), .B2(new_n870), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n856), .A2(KEYINPUT113), .ZN(new_n872));
  INV_X1    g0672(.A(KEYINPUT113), .ZN(new_n873));
  NAND4_X1  g0673(.A1(new_n851), .A2(new_n873), .A3(new_n818), .A4(new_n855), .ZN(new_n874));
  INV_X1    g0674(.A(KEYINPUT40), .ZN(new_n875));
  INV_X1    g0675(.A(KEYINPUT38), .ZN(new_n876));
  INV_X1    g0676(.A(new_n629), .ZN(new_n877));
  AOI21_X1  g0677(.A(new_n863), .B1(new_n625), .B2(new_n877), .ZN(new_n878));
  NAND3_X1  g0678(.A1(new_n401), .A2(new_n408), .A3(new_n863), .ZN(new_n879));
  XNOR2_X1  g0679(.A(new_n879), .B(new_n864), .ZN(new_n880));
  OAI21_X1  g0680(.A(new_n876), .B1(new_n878), .B2(new_n880), .ZN(new_n881));
  AOI21_X1  g0681(.A(new_n875), .B1(new_n881), .B2(new_n867), .ZN(new_n882));
  NAND3_X1  g0682(.A1(new_n872), .A2(new_n874), .A3(new_n882), .ZN(new_n883));
  INV_X1    g0683(.A(KEYINPUT114), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  NAND4_X1  g0685(.A1(new_n872), .A2(new_n882), .A3(KEYINPUT114), .A4(new_n874), .ZN(new_n886));
  AOI21_X1  g0686(.A(new_n871), .B1(new_n885), .B2(new_n886), .ZN(new_n887));
  AND3_X1   g0687(.A1(new_n887), .A2(new_n440), .A3(new_n851), .ZN(new_n888));
  AOI21_X1  g0688(.A(new_n887), .B1(new_n440), .B2(new_n851), .ZN(new_n889));
  NOR3_X1   g0689(.A1(new_n888), .A2(new_n889), .A3(new_n672), .ZN(new_n890));
  INV_X1    g0690(.A(KEYINPUT112), .ZN(new_n891));
  INV_X1    g0691(.A(KEYINPUT39), .ZN(new_n892));
  NOR3_X1   g0692(.A1(new_n621), .A2(new_n622), .A3(new_n620), .ZN(new_n893));
  AOI21_X1  g0693(.A(KEYINPUT88), .B1(new_n409), .B2(new_n412), .ZN(new_n894));
  OAI21_X1  g0694(.A(new_n877), .B1(new_n893), .B2(new_n894), .ZN(new_n895));
  INV_X1    g0695(.A(new_n863), .ZN(new_n896));
  AOI21_X1  g0696(.A(new_n880), .B1(new_n895), .B2(new_n896), .ZN(new_n897));
  OAI211_X1 g0697(.A(new_n892), .B(new_n867), .C1(new_n897), .C2(KEYINPUT38), .ZN(new_n898));
  OAI21_X1  g0698(.A(KEYINPUT39), .B1(new_n868), .B2(new_n869), .ZN(new_n899));
  AOI21_X1  g0699(.A(new_n891), .B1(new_n898), .B2(new_n899), .ZN(new_n900));
  INV_X1    g0700(.A(new_n900), .ZN(new_n901));
  INV_X1    g0701(.A(new_n341), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n902), .A2(new_n667), .ZN(new_n903));
  INV_X1    g0703(.A(new_n903), .ZN(new_n904));
  NAND3_X1  g0704(.A1(new_n898), .A2(new_n899), .A3(new_n891), .ZN(new_n905));
  NAND3_X1  g0705(.A1(new_n901), .A2(new_n904), .A3(new_n905), .ZN(new_n906));
  INV_X1    g0706(.A(new_n855), .ZN(new_n907));
  NOR2_X1   g0707(.A1(new_n438), .A2(new_n666), .ZN(new_n908));
  OAI21_X1  g0708(.A(KEYINPUT110), .B1(new_n844), .B2(new_n908), .ZN(new_n909));
  INV_X1    g0709(.A(new_n817), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n692), .A2(new_n910), .ZN(new_n911));
  INV_X1    g0711(.A(KEYINPUT110), .ZN(new_n912));
  INV_X1    g0712(.A(new_n908), .ZN(new_n913));
  NAND3_X1  g0713(.A1(new_n911), .A2(new_n912), .A3(new_n913), .ZN(new_n914));
  AOI21_X1  g0714(.A(new_n907), .B1(new_n909), .B2(new_n914), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n915), .A2(new_n870), .ZN(new_n916));
  OR2_X1    g0716(.A1(new_n625), .A2(new_n862), .ZN(new_n917));
  NAND3_X1  g0717(.A1(new_n906), .A2(new_n916), .A3(new_n917), .ZN(new_n918));
  OAI21_X1  g0718(.A(new_n440), .B1(new_n694), .B2(new_n702), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n634), .A2(new_n919), .ZN(new_n920));
  XOR2_X1   g0720(.A(new_n918), .B(new_n920), .Z(new_n921));
  OR2_X1    g0721(.A1(new_n890), .A2(new_n921), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n890), .A2(new_n921), .ZN(new_n923));
  OAI21_X1  g0723(.A(G1), .B1(new_n725), .B2(G20), .ZN(new_n924));
  NAND3_X1  g0724(.A1(new_n922), .A2(new_n923), .A3(new_n924), .ZN(new_n925));
  INV_X1    g0725(.A(new_n577), .ZN(new_n926));
  INV_X1    g0726(.A(KEYINPUT35), .ZN(new_n927));
  AOI211_X1 g0727(.A(new_n442), .B(new_n225), .C1(new_n926), .C2(new_n927), .ZN(new_n928));
  OAI22_X1  g0728(.A1(new_n928), .A2(KEYINPUT109), .B1(new_n927), .B2(new_n926), .ZN(new_n929));
  AOI21_X1  g0729(.A(new_n929), .B1(KEYINPUT109), .B2(new_n928), .ZN(new_n930));
  XOR2_X1   g0730(.A(new_n930), .B(KEYINPUT36), .Z(new_n931));
  INV_X1    g0731(.A(new_n226), .ZN(new_n932));
  OAI211_X1 g0732(.A(new_n932), .B(G77), .C1(new_n272), .C2(new_n311), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n303), .A2(G68), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n933), .A2(new_n934), .ZN(new_n935));
  NAND3_X1  g0735(.A1(new_n935), .A2(G1), .A3(new_n725), .ZN(new_n936));
  NAND3_X1  g0736(.A1(new_n925), .A2(new_n931), .A3(new_n936), .ZN(G367));
  INV_X1    g0737(.A(new_n735), .ZN(new_n938));
  OAI221_X1 g0738(.A(new_n751), .B1(new_n222), .B2(new_n427), .C1(new_n235), .C2(new_n938), .ZN(new_n939));
  AND2_X1   g0739(.A1(new_n939), .A2(new_n733), .ZN(new_n940));
  NOR2_X1   g0740(.A1(new_n642), .A2(new_n667), .ZN(new_n941));
  OR2_X1    g0741(.A1(new_n653), .A2(new_n941), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n638), .A2(new_n941), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n762), .A2(G68), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n788), .A2(G143), .ZN(new_n946));
  AOI21_X1  g0746(.A(new_n737), .B1(new_n768), .B2(G159), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n772), .A2(G150), .ZN(new_n948));
  AOI22_X1  g0748(.A1(G50), .A2(new_n778), .B1(new_n781), .B2(G77), .ZN(new_n949));
  NAND4_X1  g0749(.A1(new_n946), .A2(new_n947), .A3(new_n948), .A4(new_n949), .ZN(new_n950));
  AOI22_X1  g0750(.A1(new_n765), .A2(G137), .B1(G58), .B2(new_n776), .ZN(new_n951));
  AOI21_X1  g0751(.A(new_n950), .B1(KEYINPUT116), .B2(new_n951), .ZN(new_n952));
  OAI211_X1 g0752(.A(new_n945), .B(new_n952), .C1(KEYINPUT116), .C2(new_n951), .ZN(new_n953));
  NOR2_X1   g0753(.A1(new_n775), .A2(new_n442), .ZN(new_n954));
  XNOR2_X1  g0754(.A(new_n954), .B(KEYINPUT46), .ZN(new_n955));
  AOI22_X1  g0755(.A1(new_n768), .A2(G294), .B1(new_n772), .B2(G303), .ZN(new_n956));
  INV_X1    g0756(.A(G283), .ZN(new_n957));
  OAI21_X1  g0757(.A(new_n956), .B1(new_n957), .B2(new_n777), .ZN(new_n958));
  AOI211_X1 g0758(.A(new_n955), .B(new_n958), .C1(G311), .C2(new_n788), .ZN(new_n959));
  INV_X1    g0759(.A(G317), .ZN(new_n960));
  OAI221_X1 g0760(.A(new_n737), .B1(new_n448), .B2(new_n780), .C1(new_n828), .C2(new_n960), .ZN(new_n961));
  INV_X1    g0761(.A(KEYINPUT115), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n961), .A2(new_n962), .ZN(new_n963));
  AND2_X1   g0763(.A1(new_n959), .A2(new_n963), .ZN(new_n964));
  OAI221_X1 g0764(.A(new_n964), .B1(new_n962), .B2(new_n961), .C1(new_n416), .C2(new_n799), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n953), .A2(new_n965), .ZN(new_n966));
  XOR2_X1   g0766(.A(new_n966), .B(KEYINPUT47), .Z(new_n967));
  OAI221_X1 g0767(.A(new_n940), .B1(new_n745), .B2(new_n944), .C1(new_n967), .C2(new_n802), .ZN(new_n968));
  OAI211_X1 g0768(.A(new_n609), .B(new_n613), .C1(new_n585), .C2(new_n667), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n597), .A2(new_n666), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n969), .A2(new_n970), .ZN(new_n971));
  NAND3_X1  g0771(.A1(new_n683), .A2(new_n680), .A3(new_n971), .ZN(new_n972));
  INV_X1    g0772(.A(KEYINPUT45), .ZN(new_n973));
  NOR2_X1   g0773(.A1(new_n972), .A2(new_n973), .ZN(new_n974));
  AND2_X1   g0774(.A1(new_n972), .A2(new_n973), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n683), .A2(new_n680), .ZN(new_n976));
  INV_X1    g0776(.A(new_n971), .ZN(new_n977));
  AND3_X1   g0777(.A1(new_n976), .A2(KEYINPUT44), .A3(new_n977), .ZN(new_n978));
  AOI21_X1  g0778(.A(KEYINPUT44), .B1(new_n976), .B2(new_n977), .ZN(new_n979));
  OAI22_X1  g0779(.A1(new_n974), .A2(new_n975), .B1(new_n978), .B2(new_n979), .ZN(new_n980));
  NAND3_X1  g0780(.A1(new_n980), .A2(new_n678), .A3(new_n671), .ZN(new_n981));
  OAI221_X1 g0781(.A(new_n679), .B1(new_n978), .B2(new_n979), .C1(new_n974), .C2(new_n975), .ZN(new_n982));
  OAI21_X1  g0782(.A(new_n683), .B1(new_n671), .B2(new_n682), .ZN(new_n983));
  XNOR2_X1  g0783(.A(new_n983), .B(new_n678), .ZN(new_n984));
  NAND4_X1  g0784(.A1(new_n981), .A2(new_n982), .A3(new_n723), .A4(new_n984), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n985), .A2(new_n723), .ZN(new_n986));
  XOR2_X1   g0786(.A(new_n686), .B(KEYINPUT41), .Z(new_n987));
  INV_X1    g0787(.A(new_n987), .ZN(new_n988));
  AOI21_X1  g0788(.A(new_n729), .B1(new_n986), .B2(new_n988), .ZN(new_n989));
  OR2_X1    g0789(.A1(new_n683), .A2(new_n977), .ZN(new_n990));
  OR2_X1    g0790(.A1(new_n990), .A2(KEYINPUT42), .ZN(new_n991));
  OR2_X1    g0791(.A1(new_n969), .A2(new_n565), .ZN(new_n992));
  AOI21_X1  g0792(.A(new_n666), .B1(new_n992), .B2(new_n613), .ZN(new_n993));
  AOI21_X1  g0793(.A(new_n993), .B1(new_n990), .B2(KEYINPUT42), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n991), .A2(new_n994), .ZN(new_n995));
  INV_X1    g0795(.A(new_n944), .ZN(new_n996));
  INV_X1    g0796(.A(KEYINPUT43), .ZN(new_n997));
  NAND2_X1  g0797(.A1(new_n996), .A2(new_n997), .ZN(new_n998));
  NAND2_X1  g0798(.A1(new_n944), .A2(KEYINPUT43), .ZN(new_n999));
  NAND3_X1  g0799(.A1(new_n995), .A2(new_n998), .A3(new_n999), .ZN(new_n1000));
  NAND4_X1  g0800(.A1(new_n991), .A2(new_n994), .A3(new_n997), .A4(new_n996), .ZN(new_n1001));
  NAND2_X1  g0801(.A1(new_n1000), .A2(new_n1001), .ZN(new_n1002));
  OAI21_X1  g0802(.A(new_n1002), .B1(new_n679), .B2(new_n977), .ZN(new_n1003));
  NOR2_X1   g0803(.A1(new_n679), .A2(new_n977), .ZN(new_n1004));
  NAND3_X1  g0804(.A1(new_n1000), .A2(new_n1001), .A3(new_n1004), .ZN(new_n1005));
  NAND2_X1  g0805(.A1(new_n1003), .A2(new_n1005), .ZN(new_n1006));
  OAI21_X1  g0806(.A(new_n968), .B1(new_n989), .B2(new_n1006), .ZN(new_n1007));
  NAND2_X1  g0807(.A1(new_n1007), .A2(KEYINPUT117), .ZN(new_n1008));
  AOI21_X1  g0808(.A(new_n987), .B1(new_n985), .B2(new_n723), .ZN(new_n1009));
  OAI211_X1 g0809(.A(new_n1005), .B(new_n1003), .C1(new_n1009), .C2(new_n729), .ZN(new_n1010));
  INV_X1    g0810(.A(KEYINPUT117), .ZN(new_n1011));
  NAND3_X1  g0811(.A1(new_n1010), .A2(new_n1011), .A3(new_n968), .ZN(new_n1012));
  NAND2_X1  g0812(.A1(new_n1008), .A2(new_n1012), .ZN(new_n1013));
  INV_X1    g0813(.A(new_n1013), .ZN(G387));
  AOI22_X1  g0814(.A1(new_n768), .A2(G311), .B1(new_n778), .B2(G303), .ZN(new_n1015));
  OAI21_X1  g0815(.A(new_n1015), .B1(new_n960), .B2(new_n771), .ZN(new_n1016));
  AOI21_X1  g0816(.A(new_n1016), .B1(G322), .B2(new_n788), .ZN(new_n1017));
  XOR2_X1   g0817(.A(new_n1017), .B(KEYINPUT48), .Z(new_n1018));
  OAI221_X1 g0818(.A(new_n1018), .B1(new_n957), .B2(new_n799), .C1(new_n555), .C2(new_n775), .ZN(new_n1019));
  XOR2_X1   g0819(.A(new_n1019), .B(KEYINPUT49), .Z(new_n1020));
  NAND2_X1  g0820(.A1(new_n765), .A2(G326), .ZN(new_n1021));
  OAI211_X1 g0821(.A(new_n1021), .B(new_n737), .C1(new_n442), .C2(new_n780), .ZN(new_n1022));
  NOR2_X1   g0822(.A1(new_n1020), .A2(new_n1022), .ZN(new_n1023));
  NOR2_X1   g0823(.A1(new_n761), .A2(new_n427), .ZN(new_n1024));
  AOI22_X1  g0824(.A1(G50), .A2(new_n772), .B1(new_n776), .B2(G77), .ZN(new_n1025));
  AOI21_X1  g0825(.A(new_n737), .B1(new_n781), .B2(G97), .ZN(new_n1026));
  OAI211_X1 g0826(.A(new_n1025), .B(new_n1026), .C1(new_n311), .C2(new_n777), .ZN(new_n1027));
  XNOR2_X1  g0827(.A(KEYINPUT119), .B(G150), .ZN(new_n1028));
  AOI22_X1  g0828(.A1(new_n788), .A2(G159), .B1(new_n765), .B2(new_n1028), .ZN(new_n1029));
  INV_X1    g0829(.A(new_n279), .ZN(new_n1030));
  OAI21_X1  g0830(.A(new_n1029), .B1(new_n1030), .B2(new_n794), .ZN(new_n1031));
  NOR3_X1   g0831(.A1(new_n1024), .A2(new_n1027), .A3(new_n1031), .ZN(new_n1032));
  OAI21_X1  g0832(.A(new_n750), .B1(new_n1023), .B2(new_n1032), .ZN(new_n1033));
  INV_X1    g0833(.A(new_n688), .ZN(new_n1034));
  AOI22_X1  g0834(.A1(new_n738), .A2(new_n1034), .B1(new_n416), .B2(new_n685), .ZN(new_n1035));
  XOR2_X1   g0835(.A(new_n1035), .B(KEYINPUT118), .Z(new_n1036));
  NOR2_X1   g0836(.A1(new_n232), .A2(new_n260), .ZN(new_n1037));
  NAND2_X1  g0837(.A1(new_n360), .A2(new_n303), .ZN(new_n1038));
  XNOR2_X1  g0838(.A(new_n1038), .B(KEYINPUT50), .ZN(new_n1039));
  OAI211_X1 g0839(.A(new_n688), .B(new_n260), .C1(new_n311), .C2(new_n251), .ZN(new_n1040));
  OAI21_X1  g0840(.A(new_n735), .B1(new_n1039), .B2(new_n1040), .ZN(new_n1041));
  OAI21_X1  g0841(.A(new_n1036), .B1(new_n1037), .B2(new_n1041), .ZN(new_n1042));
  AOI21_X1  g0842(.A(new_n732), .B1(new_n1042), .B2(new_n751), .ZN(new_n1043));
  OAI211_X1 g0843(.A(new_n1033), .B(new_n1043), .C1(new_n671), .C2(new_n745), .ZN(new_n1044));
  NAND2_X1  g0844(.A1(new_n984), .A2(new_n729), .ZN(new_n1045));
  AND2_X1   g0845(.A1(new_n1044), .A2(new_n1045), .ZN(new_n1046));
  NAND2_X1  g0846(.A1(new_n984), .A2(new_n723), .ZN(new_n1047));
  XNOR2_X1  g0847(.A(new_n686), .B(KEYINPUT120), .ZN(new_n1048));
  NAND3_X1  g0848(.A1(new_n1047), .A2(KEYINPUT121), .A3(new_n1048), .ZN(new_n1049));
  OAI21_X1  g0849(.A(new_n1049), .B1(new_n723), .B2(new_n984), .ZN(new_n1050));
  AOI21_X1  g0850(.A(KEYINPUT121), .B1(new_n1047), .B2(new_n1048), .ZN(new_n1051));
  OAI21_X1  g0851(.A(new_n1046), .B1(new_n1050), .B2(new_n1051), .ZN(G393));
  NAND2_X1  g0852(.A1(new_n981), .A2(new_n982), .ZN(new_n1053));
  INV_X1    g0853(.A(new_n729), .ZN(new_n1054));
  NOR2_X1   g0854(.A1(new_n1053), .A2(new_n1054), .ZN(new_n1055));
  NAND2_X1  g0855(.A1(new_n977), .A2(new_n746), .ZN(new_n1056));
  OAI21_X1  g0856(.A(new_n751), .B1(new_n448), .B2(new_n222), .ZN(new_n1057));
  AOI21_X1  g0857(.A(new_n1057), .B1(new_n240), .B2(new_n735), .ZN(new_n1058));
  NOR2_X1   g0858(.A1(new_n761), .A2(new_n251), .ZN(new_n1059));
  INV_X1    g0859(.A(new_n1059), .ZN(new_n1060));
  AOI22_X1  g0860(.A1(new_n788), .A2(G150), .B1(G159), .B2(new_n772), .ZN(new_n1061));
  XOR2_X1   g0861(.A(new_n1061), .B(KEYINPUT51), .Z(new_n1062));
  NAND2_X1  g0862(.A1(new_n820), .A2(new_n247), .ZN(new_n1063));
  AOI22_X1  g0863(.A1(new_n768), .A2(G50), .B1(new_n776), .B2(G68), .ZN(new_n1064));
  OAI21_X1  g0864(.A(new_n1064), .B1(new_n424), .B2(new_n777), .ZN(new_n1065));
  AOI211_X1 g0865(.A(new_n1063), .B(new_n1065), .C1(G143), .C2(new_n765), .ZN(new_n1066));
  NAND3_X1  g0866(.A1(new_n1060), .A2(new_n1062), .A3(new_n1066), .ZN(new_n1067));
  AOI22_X1  g0867(.A1(new_n788), .A2(G317), .B1(G311), .B2(new_n772), .ZN(new_n1068));
  XNOR2_X1  g0868(.A(new_n1068), .B(KEYINPUT52), .ZN(new_n1069));
  OAI21_X1  g0869(.A(new_n737), .B1(new_n780), .B2(new_n416), .ZN(new_n1070));
  AOI22_X1  g0870(.A1(G283), .A2(new_n776), .B1(new_n778), .B2(G294), .ZN(new_n1071));
  OAI21_X1  g0871(.A(new_n1071), .B1(new_n793), .B2(new_n794), .ZN(new_n1072));
  AOI211_X1 g0872(.A(new_n1070), .B(new_n1072), .C1(G322), .C2(new_n765), .ZN(new_n1073));
  OAI21_X1  g0873(.A(new_n1073), .B1(new_n442), .B2(new_n799), .ZN(new_n1074));
  OAI21_X1  g0874(.A(new_n1067), .B1(new_n1069), .B2(new_n1074), .ZN(new_n1075));
  AOI211_X1 g0875(.A(new_n732), .B(new_n1058), .C1(new_n1075), .C2(new_n750), .ZN(new_n1076));
  AOI21_X1  g0876(.A(new_n1055), .B1(new_n1056), .B2(new_n1076), .ZN(new_n1077));
  NAND2_X1  g0877(.A1(new_n1053), .A2(new_n1047), .ZN(new_n1078));
  NAND3_X1  g0878(.A1(new_n1078), .A2(new_n985), .A3(new_n1048), .ZN(new_n1079));
  NAND2_X1  g0879(.A1(new_n1077), .A2(new_n1079), .ZN(G390));
  AND3_X1   g0880(.A1(new_n851), .A2(G330), .A3(new_n818), .ZN(new_n1081));
  NAND2_X1  g0881(.A1(new_n1081), .A2(new_n855), .ZN(new_n1082));
  AND2_X1   g0882(.A1(new_n722), .A2(new_n818), .ZN(new_n1083));
  OAI21_X1  g0883(.A(new_n1082), .B1(new_n1083), .B2(new_n855), .ZN(new_n1084));
  NAND2_X1  g0884(.A1(new_n909), .A2(new_n914), .ZN(new_n1085));
  NAND2_X1  g0885(.A1(new_n1084), .A2(new_n1085), .ZN(new_n1086));
  NAND2_X1  g0886(.A1(new_n1083), .A2(new_n855), .ZN(new_n1087));
  AOI21_X1  g0887(.A(new_n908), .B1(new_n701), .B2(new_n910), .ZN(new_n1088));
  OAI211_X1 g0888(.A(new_n1087), .B(new_n1088), .C1(new_n855), .C2(new_n1081), .ZN(new_n1089));
  NAND2_X1  g0889(.A1(new_n1086), .A2(new_n1089), .ZN(new_n1090));
  NAND3_X1  g0890(.A1(new_n440), .A2(G330), .A3(new_n851), .ZN(new_n1091));
  NAND3_X1  g0891(.A1(new_n634), .A2(new_n919), .A3(new_n1091), .ZN(new_n1092));
  INV_X1    g0892(.A(new_n1092), .ZN(new_n1093));
  NAND2_X1  g0893(.A1(new_n1090), .A2(new_n1093), .ZN(new_n1094));
  AND3_X1   g0894(.A1(new_n898), .A2(new_n899), .A3(new_n891), .ZN(new_n1095));
  OAI22_X1  g0895(.A1(new_n915), .A2(new_n904), .B1(new_n1095), .B2(new_n900), .ZN(new_n1096));
  NOR2_X1   g0896(.A1(new_n1088), .A2(new_n907), .ZN(new_n1097));
  NAND2_X1  g0897(.A1(new_n881), .A2(new_n867), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n1098), .A2(new_n903), .ZN(new_n1099));
  NOR2_X1   g0899(.A1(new_n1097), .A2(new_n1099), .ZN(new_n1100));
  INV_X1    g0900(.A(new_n1100), .ZN(new_n1101));
  AND3_X1   g0901(.A1(new_n1096), .A2(new_n1101), .A3(new_n1087), .ZN(new_n1102));
  AOI21_X1  g0902(.A(new_n1082), .B1(new_n1096), .B2(new_n1101), .ZN(new_n1103));
  OAI21_X1  g0903(.A(new_n1094), .B1(new_n1102), .B2(new_n1103), .ZN(new_n1104));
  NAND3_X1  g0904(.A1(new_n1096), .A2(new_n1101), .A3(new_n1087), .ZN(new_n1105));
  AOI21_X1  g0905(.A(new_n1092), .B1(new_n1086), .B2(new_n1089), .ZN(new_n1106));
  NOR3_X1   g0906(.A1(new_n844), .A2(KEYINPUT110), .A3(new_n908), .ZN(new_n1107));
  AOI21_X1  g0907(.A(new_n912), .B1(new_n911), .B2(new_n913), .ZN(new_n1108));
  OAI21_X1  g0908(.A(new_n855), .B1(new_n1107), .B2(new_n1108), .ZN(new_n1109));
  NAND2_X1  g0909(.A1(new_n1109), .A2(new_n903), .ZN(new_n1110));
  NAND2_X1  g0910(.A1(new_n901), .A2(new_n905), .ZN(new_n1111));
  AOI21_X1  g0911(.A(new_n1100), .B1(new_n1110), .B2(new_n1111), .ZN(new_n1112));
  OAI211_X1 g0912(.A(new_n1105), .B(new_n1106), .C1(new_n1112), .C2(new_n1082), .ZN(new_n1113));
  NAND3_X1  g0913(.A1(new_n1104), .A2(new_n1113), .A3(new_n1048), .ZN(new_n1114));
  OAI211_X1 g0914(.A(new_n1105), .B(new_n729), .C1(new_n1112), .C2(new_n1082), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n1111), .A2(new_n742), .ZN(new_n1116));
  AOI22_X1  g0916(.A1(new_n768), .A2(G107), .B1(new_n778), .B2(G97), .ZN(new_n1117));
  OAI21_X1  g0917(.A(new_n1117), .B1(new_n834), .B2(new_n957), .ZN(new_n1118));
  AND2_X1   g0918(.A1(new_n1118), .A2(KEYINPUT122), .ZN(new_n1119));
  NOR2_X1   g0919(.A1(new_n1118), .A2(KEYINPUT122), .ZN(new_n1120));
  NOR2_X1   g0920(.A1(new_n828), .A2(new_n555), .ZN(new_n1121));
  AOI21_X1  g0921(.A(new_n247), .B1(new_n776), .B2(G87), .ZN(new_n1122));
  OAI211_X1 g0922(.A(new_n1122), .B(new_n831), .C1(new_n442), .C2(new_n771), .ZN(new_n1123));
  NOR4_X1   g0923(.A1(new_n1119), .A2(new_n1120), .A3(new_n1121), .A4(new_n1123), .ZN(new_n1124));
  NAND2_X1  g0924(.A1(new_n762), .A2(G159), .ZN(new_n1125));
  AOI21_X1  g0925(.A(new_n737), .B1(new_n768), .B2(G137), .ZN(new_n1126));
  XNOR2_X1  g0926(.A(KEYINPUT54), .B(G143), .ZN(new_n1127));
  INV_X1    g0927(.A(new_n1127), .ZN(new_n1128));
  AOI22_X1  g0928(.A1(new_n778), .A2(new_n1128), .B1(new_n781), .B2(G50), .ZN(new_n1129));
  OAI211_X1 g0929(.A(new_n1126), .B(new_n1129), .C1(new_n829), .C2(new_n771), .ZN(new_n1130));
  NAND2_X1  g0930(.A1(new_n776), .A2(new_n1028), .ZN(new_n1131));
  XOR2_X1   g0931(.A(new_n1131), .B(KEYINPUT53), .Z(new_n1132));
  INV_X1    g0932(.A(G128), .ZN(new_n1133));
  OAI21_X1  g0933(.A(new_n1132), .B1(new_n1133), .B2(new_n834), .ZN(new_n1134));
  AOI211_X1 g0934(.A(new_n1130), .B(new_n1134), .C1(G125), .C2(new_n765), .ZN(new_n1135));
  AOI22_X1  g0935(.A1(new_n1124), .A2(new_n1060), .B1(new_n1125), .B2(new_n1135), .ZN(new_n1136));
  OAI221_X1 g0936(.A(new_n733), .B1(new_n279), .B2(new_n813), .C1(new_n1136), .C2(new_n802), .ZN(new_n1137));
  XOR2_X1   g0937(.A(new_n1137), .B(KEYINPUT123), .Z(new_n1138));
  NAND2_X1  g0938(.A1(new_n1116), .A2(new_n1138), .ZN(new_n1139));
  AND2_X1   g0939(.A1(new_n1115), .A2(new_n1139), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n1114), .A2(new_n1140), .ZN(G378));
  INV_X1    g0941(.A(new_n1048), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n885), .A2(new_n886), .ZN(new_n1143));
  INV_X1    g0943(.A(new_n871), .ZN(new_n1144));
  NOR2_X1   g0944(.A1(new_n292), .A2(new_n664), .ZN(new_n1145));
  XNOR2_X1  g0945(.A(new_n300), .B(new_n1145), .ZN(new_n1146));
  XNOR2_X1  g0946(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1147));
  XOR2_X1   g0947(.A(new_n1146), .B(new_n1147), .Z(new_n1148));
  AND4_X1   g0948(.A1(G330), .A2(new_n1143), .A3(new_n1144), .A4(new_n1148), .ZN(new_n1149));
  AOI21_X1  g0949(.A(new_n1148), .B1(new_n887), .B2(G330), .ZN(new_n1150));
  OAI21_X1  g0950(.A(new_n918), .B1(new_n1149), .B2(new_n1150), .ZN(new_n1151));
  NAND3_X1  g0951(.A1(new_n1143), .A2(G330), .A3(new_n1144), .ZN(new_n1152));
  INV_X1    g0952(.A(new_n1148), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n1152), .A2(new_n1153), .ZN(new_n1154));
  INV_X1    g0954(.A(new_n918), .ZN(new_n1155));
  NAND3_X1  g0955(.A1(new_n887), .A2(G330), .A3(new_n1148), .ZN(new_n1156));
  NAND3_X1  g0956(.A1(new_n1154), .A2(new_n1155), .A3(new_n1156), .ZN(new_n1157));
  AOI22_X1  g0957(.A1(new_n1151), .A2(new_n1157), .B1(new_n1093), .B2(new_n1113), .ZN(new_n1158));
  AOI21_X1  g0958(.A(new_n1142), .B1(new_n1158), .B2(KEYINPUT57), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n1113), .A2(new_n1093), .ZN(new_n1160));
  NOR3_X1   g0960(.A1(new_n1149), .A2(new_n1150), .A3(new_n918), .ZN(new_n1161));
  AOI21_X1  g0961(.A(new_n1155), .B1(new_n1154), .B2(new_n1156), .ZN(new_n1162));
  OAI21_X1  g0962(.A(new_n1160), .B1(new_n1161), .B2(new_n1162), .ZN(new_n1163));
  INV_X1    g0963(.A(KEYINPUT57), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n1163), .A2(new_n1164), .ZN(new_n1165));
  NAND2_X1  g0965(.A1(new_n1159), .A2(new_n1165), .ZN(new_n1166));
  OAI21_X1  g0966(.A(new_n729), .B1(new_n1161), .B2(new_n1162), .ZN(new_n1167));
  NAND2_X1  g0967(.A1(new_n1153), .A2(new_n742), .ZN(new_n1168));
  OAI21_X1  g0968(.A(new_n733), .B1(G50), .B2(new_n813), .ZN(new_n1169));
  AOI21_X1  g0969(.A(G50), .B1(new_n347), .B2(new_n259), .ZN(new_n1170));
  OAI22_X1  g0970(.A1(new_n794), .A2(new_n448), .B1(new_n780), .B2(new_n272), .ZN(new_n1171));
  OAI211_X1 g0971(.A(new_n737), .B(new_n259), .C1(new_n251), .C2(new_n775), .ZN(new_n1172));
  OAI22_X1  g0972(.A1(new_n771), .A2(new_n416), .B1(new_n777), .B2(new_n427), .ZN(new_n1173));
  NOR3_X1   g0973(.A1(new_n1171), .A2(new_n1172), .A3(new_n1173), .ZN(new_n1174));
  AOI22_X1  g0974(.A1(new_n788), .A2(G116), .B1(new_n765), .B2(G283), .ZN(new_n1175));
  NAND3_X1  g0975(.A1(new_n945), .A2(new_n1174), .A3(new_n1175), .ZN(new_n1176));
  INV_X1    g0976(.A(KEYINPUT58), .ZN(new_n1177));
  AOI21_X1  g0977(.A(new_n1170), .B1(new_n1176), .B2(new_n1177), .ZN(new_n1178));
  XNOR2_X1  g0978(.A(new_n1178), .B(KEYINPUT124), .ZN(new_n1179));
  OAI22_X1  g0979(.A1(new_n1133), .A2(new_n771), .B1(new_n775), .B2(new_n1127), .ZN(new_n1180));
  OAI22_X1  g0980(.A1(new_n794), .A2(new_n829), .B1(new_n835), .B2(new_n777), .ZN(new_n1181));
  AOI211_X1 g0981(.A(new_n1180), .B(new_n1181), .C1(new_n788), .C2(G125), .ZN(new_n1182));
  OAI21_X1  g0982(.A(new_n1182), .B1(new_n761), .B2(new_n270), .ZN(new_n1183));
  NOR2_X1   g0983(.A1(new_n1183), .A2(KEYINPUT59), .ZN(new_n1184));
  NAND2_X1  g0984(.A1(new_n1183), .A2(KEYINPUT59), .ZN(new_n1185));
  OAI211_X1 g0985(.A(new_n268), .B(new_n259), .C1(new_n780), .C2(new_n353), .ZN(new_n1186));
  AOI21_X1  g0986(.A(new_n1186), .B1(new_n765), .B2(G124), .ZN(new_n1187));
  NAND2_X1  g0987(.A1(new_n1185), .A2(new_n1187), .ZN(new_n1188));
  OAI221_X1 g0988(.A(new_n1179), .B1(new_n1177), .B2(new_n1176), .C1(new_n1184), .C2(new_n1188), .ZN(new_n1189));
  AOI21_X1  g0989(.A(new_n1169), .B1(new_n1189), .B2(new_n750), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n1168), .A2(new_n1190), .ZN(new_n1191));
  NAND2_X1  g0991(.A1(new_n1167), .A2(new_n1191), .ZN(new_n1192));
  INV_X1    g0992(.A(new_n1192), .ZN(new_n1193));
  NAND2_X1  g0993(.A1(new_n1166), .A2(new_n1193), .ZN(G375));
  INV_X1    g0994(.A(KEYINPUT125), .ZN(new_n1195));
  OAI21_X1  g0995(.A(new_n1195), .B1(new_n1090), .B2(new_n1093), .ZN(new_n1196));
  NAND4_X1  g0996(.A1(new_n1086), .A2(KEYINPUT125), .A3(new_n1092), .A4(new_n1089), .ZN(new_n1197));
  NAND4_X1  g0997(.A1(new_n1196), .A2(new_n988), .A3(new_n1094), .A4(new_n1197), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(new_n907), .A2(new_n742), .ZN(new_n1199));
  OAI21_X1  g0999(.A(new_n733), .B1(G68), .B2(new_n813), .ZN(new_n1200));
  OAI21_X1  g1000(.A(new_n247), .B1(new_n780), .B2(new_n272), .ZN(new_n1201));
  OAI22_X1  g1001(.A1(new_n775), .A2(new_n353), .B1(new_n777), .B2(new_n270), .ZN(new_n1202));
  AOI211_X1 g1002(.A(new_n1201), .B(new_n1202), .C1(G128), .C2(new_n765), .ZN(new_n1203));
  OAI21_X1  g1003(.A(new_n1203), .B1(new_n761), .B2(new_n303), .ZN(new_n1204));
  XOR2_X1   g1004(.A(new_n1204), .B(KEYINPUT126), .Z(new_n1205));
  AOI22_X1  g1005(.A1(new_n768), .A2(new_n1128), .B1(new_n772), .B2(G137), .ZN(new_n1206));
  OAI21_X1  g1006(.A(new_n1206), .B1(new_n834), .B2(new_n829), .ZN(new_n1207));
  AOI22_X1  g1007(.A1(new_n788), .A2(G294), .B1(new_n765), .B2(G303), .ZN(new_n1208));
  AOI21_X1  g1008(.A(new_n247), .B1(new_n781), .B2(G77), .ZN(new_n1209));
  AOI22_X1  g1009(.A1(G97), .A2(new_n776), .B1(new_n772), .B2(G283), .ZN(new_n1210));
  AOI22_X1  g1010(.A1(new_n768), .A2(G116), .B1(new_n778), .B2(G107), .ZN(new_n1211));
  NAND4_X1  g1011(.A1(new_n1208), .A2(new_n1209), .A3(new_n1210), .A4(new_n1211), .ZN(new_n1212));
  OAI22_X1  g1012(.A1(new_n1205), .A2(new_n1207), .B1(new_n1024), .B2(new_n1212), .ZN(new_n1213));
  AOI21_X1  g1013(.A(new_n1200), .B1(new_n1213), .B2(new_n750), .ZN(new_n1214));
  AOI22_X1  g1014(.A1(new_n1090), .A2(new_n729), .B1(new_n1199), .B2(new_n1214), .ZN(new_n1215));
  NAND2_X1  g1015(.A1(new_n1198), .A2(new_n1215), .ZN(G381));
  AOI21_X1  g1016(.A(new_n1192), .B1(new_n1159), .B2(new_n1165), .ZN(new_n1217));
  INV_X1    g1017(.A(G378), .ZN(new_n1218));
  OR2_X1    g1018(.A1(G393), .A2(G396), .ZN(new_n1219));
  NOR4_X1   g1019(.A1(new_n1219), .A2(G381), .A3(G390), .A4(G384), .ZN(new_n1220));
  NAND4_X1  g1020(.A1(new_n1217), .A2(new_n1013), .A3(new_n1218), .A4(new_n1220), .ZN(G407));
  NAND2_X1  g1021(.A1(new_n1217), .A2(new_n1218), .ZN(new_n1222));
  OAI211_X1 g1022(.A(G407), .B(G213), .C1(G343), .C2(new_n1222), .ZN(G409));
  AND2_X1   g1023(.A1(new_n665), .A2(G213), .ZN(new_n1224));
  AOI21_X1  g1024(.A(new_n1054), .B1(new_n1151), .B2(new_n1157), .ZN(new_n1225));
  INV_X1    g1025(.A(new_n1191), .ZN(new_n1226));
  NOR3_X1   g1026(.A1(G378), .A2(new_n1225), .A3(new_n1226), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(new_n1158), .A2(new_n988), .ZN(new_n1228));
  AOI21_X1  g1028(.A(new_n1224), .B1(new_n1227), .B2(new_n1228), .ZN(new_n1229));
  OAI21_X1  g1029(.A(new_n1229), .B1(new_n1218), .B2(new_n1217), .ZN(new_n1230));
  NAND2_X1  g1030(.A1(new_n1224), .A2(G2897), .ZN(new_n1231));
  INV_X1    g1031(.A(KEYINPUT60), .ZN(new_n1232));
  OAI211_X1 g1032(.A(new_n1196), .B(new_n1197), .C1(new_n1232), .C2(new_n1106), .ZN(new_n1233));
  NOR2_X1   g1033(.A1(new_n1090), .A2(new_n1093), .ZN(new_n1234));
  AOI21_X1  g1034(.A(new_n1142), .B1(new_n1234), .B2(KEYINPUT60), .ZN(new_n1235));
  NAND2_X1  g1035(.A1(new_n1233), .A2(new_n1235), .ZN(new_n1236));
  NAND3_X1  g1036(.A1(new_n1236), .A2(new_n849), .A3(new_n1215), .ZN(new_n1237));
  INV_X1    g1037(.A(new_n1237), .ZN(new_n1238));
  AOI21_X1  g1038(.A(new_n849), .B1(new_n1236), .B2(new_n1215), .ZN(new_n1239));
  OAI21_X1  g1039(.A(new_n1231), .B1(new_n1238), .B2(new_n1239), .ZN(new_n1240));
  NAND2_X1  g1040(.A1(new_n1236), .A2(new_n1215), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(new_n1241), .A2(G384), .ZN(new_n1242));
  INV_X1    g1042(.A(new_n1231), .ZN(new_n1243));
  NAND3_X1  g1043(.A1(new_n1242), .A2(new_n1237), .A3(new_n1243), .ZN(new_n1244));
  AND2_X1   g1044(.A1(new_n1240), .A2(new_n1244), .ZN(new_n1245));
  AOI21_X1  g1045(.A(KEYINPUT61), .B1(new_n1230), .B2(new_n1245), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(new_n1242), .A2(new_n1237), .ZN(new_n1247));
  OAI211_X1 g1047(.A(new_n1229), .B(new_n1247), .C1(new_n1218), .C2(new_n1217), .ZN(new_n1248));
  NAND2_X1  g1048(.A1(new_n1248), .A2(KEYINPUT62), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(G375), .A2(G378), .ZN(new_n1250));
  INV_X1    g1050(.A(KEYINPUT62), .ZN(new_n1251));
  NAND4_X1  g1051(.A1(new_n1250), .A2(new_n1251), .A3(new_n1229), .A4(new_n1247), .ZN(new_n1252));
  NAND3_X1  g1052(.A1(new_n1246), .A2(new_n1249), .A3(new_n1252), .ZN(new_n1253));
  INV_X1    g1053(.A(G390), .ZN(new_n1254));
  NAND3_X1  g1054(.A1(new_n1008), .A2(new_n1012), .A3(new_n1254), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(new_n1255), .A2(KEYINPUT127), .ZN(new_n1256));
  INV_X1    g1056(.A(KEYINPUT127), .ZN(new_n1257));
  NAND4_X1  g1057(.A1(new_n1008), .A2(new_n1257), .A3(new_n1012), .A4(new_n1254), .ZN(new_n1258));
  NOR2_X1   g1058(.A1(new_n1254), .A2(new_n1007), .ZN(new_n1259));
  XNOR2_X1  g1059(.A(G393), .B(new_n811), .ZN(new_n1260));
  NOR2_X1   g1060(.A1(new_n1259), .A2(new_n1260), .ZN(new_n1261));
  NAND3_X1  g1061(.A1(new_n1256), .A2(new_n1258), .A3(new_n1261), .ZN(new_n1262));
  AOI21_X1  g1062(.A(G390), .B1(new_n1010), .B2(new_n968), .ZN(new_n1263));
  OAI21_X1  g1063(.A(new_n1260), .B1(new_n1259), .B2(new_n1263), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(new_n1262), .A2(new_n1264), .ZN(new_n1265));
  INV_X1    g1065(.A(new_n1265), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(new_n1253), .A2(new_n1266), .ZN(new_n1267));
  INV_X1    g1067(.A(KEYINPUT63), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1248), .A2(new_n1268), .ZN(new_n1269));
  NAND4_X1  g1069(.A1(new_n1250), .A2(KEYINPUT63), .A3(new_n1229), .A4(new_n1247), .ZN(new_n1270));
  NAND4_X1  g1070(.A1(new_n1246), .A2(new_n1269), .A3(new_n1270), .A4(new_n1265), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(new_n1267), .A2(new_n1271), .ZN(G405));
  AOI21_X1  g1072(.A(new_n1247), .B1(new_n1262), .B2(new_n1264), .ZN(new_n1273));
  INV_X1    g1073(.A(new_n1273), .ZN(new_n1274));
  NAND3_X1  g1074(.A1(new_n1262), .A2(new_n1264), .A3(new_n1247), .ZN(new_n1275));
  AOI22_X1  g1075(.A1(new_n1274), .A2(new_n1275), .B1(new_n1222), .B2(new_n1250), .ZN(new_n1276));
  INV_X1    g1076(.A(new_n1275), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(new_n1250), .A2(new_n1222), .ZN(new_n1278));
  NOR3_X1   g1078(.A1(new_n1277), .A2(new_n1278), .A3(new_n1273), .ZN(new_n1279));
  NOR2_X1   g1079(.A1(new_n1276), .A2(new_n1279), .ZN(G402));
endmodule


