//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 0 1 0 0 1 0 1 1 0 1 0 1 0 0 0 0 1 0 0 1 1 1 1 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 1 0 0 0 1 0 1 1 1 1 0 0 1 0 1 1 1 0 0 1 0 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:24:44 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n709, new_n710,
    new_n711, new_n712, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n731, new_n732, new_n734, new_n735,
    new_n736, new_n737, new_n738, new_n739, new_n740, new_n741, new_n742,
    new_n743, new_n744, new_n745, new_n747, new_n748, new_n749, new_n750,
    new_n751, new_n752, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n771, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n790, new_n791, new_n792, new_n793, new_n794, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n908, new_n909, new_n910,
    new_n911, new_n912, new_n913, new_n914, new_n915, new_n916, new_n917,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n935, new_n936, new_n937, new_n938, new_n939, new_n940, new_n941,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n951, new_n952, new_n953, new_n954, new_n955, new_n956,
    new_n957, new_n958, new_n960, new_n961, new_n962, new_n963, new_n964,
    new_n965, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1021, new_n1022, new_n1023, new_n1024;
  OAI21_X1  g000(.A(G214), .B1(G237), .B2(G902), .ZN(new_n187));
  INV_X1    g001(.A(G146), .ZN(new_n188));
  NOR2_X1   g002(.A1(new_n188), .A2(G143), .ZN(new_n189));
  INV_X1    g003(.A(G143), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n190), .A2(KEYINPUT65), .ZN(new_n191));
  INV_X1    g005(.A(KEYINPUT65), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n192), .A2(G143), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n191), .A2(new_n193), .ZN(new_n194));
  AOI21_X1  g008(.A(new_n189), .B1(new_n194), .B2(new_n188), .ZN(new_n195));
  INV_X1    g009(.A(G128), .ZN(new_n196));
  NOR2_X1   g010(.A1(new_n190), .A2(G146), .ZN(new_n197));
  INV_X1    g011(.A(new_n197), .ZN(new_n198));
  AOI21_X1  g012(.A(new_n196), .B1(new_n198), .B2(KEYINPUT1), .ZN(new_n199));
  NOR2_X1   g013(.A1(new_n195), .A2(new_n199), .ZN(new_n200));
  INV_X1    g014(.A(KEYINPUT1), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n201), .A2(G128), .ZN(new_n202));
  XNOR2_X1  g016(.A(KEYINPUT65), .B(G143), .ZN(new_n203));
  AOI211_X1 g017(.A(new_n197), .B(new_n202), .C1(new_n203), .C2(G146), .ZN(new_n204));
  NOR2_X1   g018(.A1(new_n200), .A2(new_n204), .ZN(new_n205));
  INV_X1    g019(.A(G125), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  OAI21_X1  g021(.A(KEYINPUT64), .B1(KEYINPUT0), .B2(G128), .ZN(new_n208));
  INV_X1    g022(.A(new_n208), .ZN(new_n209));
  NOR3_X1   g023(.A1(KEYINPUT64), .A2(KEYINPUT0), .A3(G128), .ZN(new_n210));
  INV_X1    g024(.A(KEYINPUT0), .ZN(new_n211));
  OAI22_X1  g025(.A1(new_n209), .A2(new_n210), .B1(new_n211), .B2(new_n196), .ZN(new_n212));
  OAI21_X1  g026(.A(KEYINPUT66), .B1(new_n195), .B2(new_n212), .ZN(new_n213));
  INV_X1    g027(.A(new_n189), .ZN(new_n214));
  OAI21_X1  g028(.A(new_n214), .B1(new_n203), .B2(G146), .ZN(new_n215));
  NOR2_X1   g029(.A1(new_n211), .A2(new_n196), .ZN(new_n216));
  OR3_X1    g030(.A1(KEYINPUT64), .A2(KEYINPUT0), .A3(G128), .ZN(new_n217));
  AOI21_X1  g031(.A(new_n216), .B1(new_n217), .B2(new_n208), .ZN(new_n218));
  INV_X1    g032(.A(KEYINPUT66), .ZN(new_n219));
  NAND3_X1  g033(.A1(new_n215), .A2(new_n218), .A3(new_n219), .ZN(new_n220));
  AOI21_X1  g034(.A(new_n197), .B1(new_n203), .B2(G146), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n221), .A2(new_n216), .ZN(new_n222));
  NAND3_X1  g036(.A1(new_n213), .A2(new_n220), .A3(new_n222), .ZN(new_n223));
  INV_X1    g037(.A(new_n223), .ZN(new_n224));
  OAI21_X1  g038(.A(new_n207), .B1(new_n224), .B2(new_n206), .ZN(new_n225));
  INV_X1    g039(.A(G953), .ZN(new_n226));
  AND2_X1   g040(.A1(new_n226), .A2(G224), .ZN(new_n227));
  XOR2_X1   g041(.A(new_n225), .B(new_n227), .Z(new_n228));
  INV_X1    g042(.A(KEYINPUT6), .ZN(new_n229));
  XNOR2_X1  g043(.A(G110), .B(G122), .ZN(new_n230));
  INV_X1    g044(.A(new_n230), .ZN(new_n231));
  INV_X1    g045(.A(G119), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n232), .A2(G116), .ZN(new_n233));
  INV_X1    g047(.A(G116), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n234), .A2(G119), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n233), .A2(new_n235), .ZN(new_n236));
  XNOR2_X1  g050(.A(KEYINPUT2), .B(G113), .ZN(new_n237));
  OR2_X1    g051(.A1(new_n236), .A2(new_n237), .ZN(new_n238));
  INV_X1    g052(.A(KEYINPUT69), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n236), .A2(new_n237), .ZN(new_n240));
  NAND3_X1  g054(.A1(new_n238), .A2(new_n239), .A3(new_n240), .ZN(new_n241));
  NAND3_X1  g055(.A1(new_n236), .A2(new_n237), .A3(KEYINPUT69), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n241), .A2(new_n242), .ZN(new_n243));
  INV_X1    g057(.A(new_n243), .ZN(new_n244));
  INV_X1    g058(.A(KEYINPUT4), .ZN(new_n245));
  XNOR2_X1  g059(.A(KEYINPUT79), .B(G104), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n246), .A2(G107), .ZN(new_n247));
  INV_X1    g061(.A(KEYINPUT3), .ZN(new_n248));
  INV_X1    g062(.A(G107), .ZN(new_n249));
  NAND3_X1  g063(.A1(new_n248), .A2(new_n249), .A3(G104), .ZN(new_n250));
  INV_X1    g064(.A(G104), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n251), .A2(KEYINPUT79), .ZN(new_n252));
  INV_X1    g066(.A(KEYINPUT79), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n253), .A2(G104), .ZN(new_n254));
  AOI21_X1  g068(.A(G107), .B1(new_n252), .B2(new_n254), .ZN(new_n255));
  OAI211_X1 g069(.A(new_n247), .B(new_n250), .C1(new_n248), .C2(new_n255), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n256), .A2(G101), .ZN(new_n257));
  OAI21_X1  g071(.A(KEYINPUT3), .B1(new_n246), .B2(G107), .ZN(new_n258));
  INV_X1    g072(.A(G101), .ZN(new_n259));
  NAND4_X1  g073(.A1(new_n258), .A2(new_n259), .A3(new_n250), .A4(new_n247), .ZN(new_n260));
  AOI21_X1  g074(.A(new_n245), .B1(new_n257), .B2(new_n260), .ZN(new_n261));
  AOI21_X1  g075(.A(KEYINPUT4), .B1(new_n256), .B2(G101), .ZN(new_n262));
  OAI21_X1  g076(.A(new_n244), .B1(new_n261), .B2(new_n262), .ZN(new_n263));
  INV_X1    g077(.A(KEYINPUT81), .ZN(new_n264));
  NAND3_X1  g078(.A1(new_n233), .A2(new_n235), .A3(KEYINPUT5), .ZN(new_n265));
  OAI211_X1 g079(.A(new_n265), .B(G113), .C1(KEYINPUT5), .C2(new_n233), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n266), .A2(new_n238), .ZN(new_n267));
  INV_X1    g081(.A(new_n267), .ZN(new_n268));
  INV_X1    g082(.A(KEYINPUT80), .ZN(new_n269));
  NOR2_X1   g083(.A1(new_n249), .A2(G104), .ZN(new_n270));
  OAI21_X1  g084(.A(G101), .B1(new_n255), .B2(new_n270), .ZN(new_n271));
  OAI21_X1  g085(.A(new_n250), .B1(new_n255), .B2(new_n248), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n247), .A2(new_n259), .ZN(new_n273));
  OAI211_X1 g087(.A(new_n269), .B(new_n271), .C1(new_n272), .C2(new_n273), .ZN(new_n274));
  INV_X1    g088(.A(new_n274), .ZN(new_n275));
  AOI21_X1  g089(.A(new_n269), .B1(new_n260), .B2(new_n271), .ZN(new_n276));
  OAI211_X1 g090(.A(new_n264), .B(new_n268), .C1(new_n275), .C2(new_n276), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n263), .A2(new_n277), .ZN(new_n278));
  OAI21_X1  g092(.A(new_n271), .B1(new_n272), .B2(new_n273), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n279), .A2(KEYINPUT80), .ZN(new_n280));
  AOI21_X1  g094(.A(new_n267), .B1(new_n280), .B2(new_n274), .ZN(new_n281));
  NOR2_X1   g095(.A1(new_n281), .A2(new_n264), .ZN(new_n282));
  OAI211_X1 g096(.A(new_n229), .B(new_n231), .C1(new_n278), .C2(new_n282), .ZN(new_n283));
  INV_X1    g097(.A(new_n283), .ZN(new_n284));
  OAI21_X1  g098(.A(new_n268), .B1(new_n275), .B2(new_n276), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n285), .A2(KEYINPUT81), .ZN(new_n286));
  NAND4_X1  g100(.A1(new_n286), .A2(new_n230), .A3(new_n277), .A4(new_n263), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n287), .A2(KEYINPUT82), .ZN(new_n288));
  AND2_X1   g102(.A1(new_n263), .A2(new_n277), .ZN(new_n289));
  INV_X1    g103(.A(KEYINPUT82), .ZN(new_n290));
  NAND4_X1  g104(.A1(new_n289), .A2(new_n290), .A3(new_n230), .A4(new_n286), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n288), .A2(new_n291), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n289), .A2(new_n286), .ZN(new_n293));
  AOI21_X1  g107(.A(new_n229), .B1(new_n293), .B2(new_n231), .ZN(new_n294));
  AOI211_X1 g108(.A(new_n228), .B(new_n284), .C1(new_n292), .C2(new_n294), .ZN(new_n295));
  XNOR2_X1  g109(.A(new_n230), .B(KEYINPUT8), .ZN(new_n296));
  AND2_X1   g110(.A1(new_n279), .A2(new_n267), .ZN(new_n297));
  OAI21_X1  g111(.A(new_n296), .B1(new_n281), .B2(new_n297), .ZN(new_n298));
  INV_X1    g112(.A(KEYINPUT7), .ZN(new_n299));
  INV_X1    g113(.A(KEYINPUT84), .ZN(new_n300));
  AOI21_X1  g114(.A(new_n299), .B1(new_n227), .B2(new_n300), .ZN(new_n301));
  OAI21_X1  g115(.A(new_n301), .B1(new_n300), .B2(new_n227), .ZN(new_n302));
  OAI21_X1  g116(.A(new_n298), .B1(new_n225), .B2(new_n302), .ZN(new_n303));
  OAI21_X1  g117(.A(new_n225), .B1(new_n299), .B2(new_n227), .ZN(new_n304));
  INV_X1    g118(.A(KEYINPUT83), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  OAI211_X1 g120(.A(new_n225), .B(KEYINPUT83), .C1(new_n299), .C2(new_n227), .ZN(new_n307));
  AOI21_X1  g121(.A(new_n303), .B1(new_n306), .B2(new_n307), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n292), .A2(new_n308), .ZN(new_n309));
  INV_X1    g123(.A(G902), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  OAI21_X1  g125(.A(G210), .B1(G237), .B2(G902), .ZN(new_n312));
  INV_X1    g126(.A(new_n312), .ZN(new_n313));
  NOR3_X1   g127(.A1(new_n295), .A2(new_n311), .A3(new_n313), .ZN(new_n314));
  AOI21_X1  g128(.A(new_n284), .B1(new_n292), .B2(new_n294), .ZN(new_n315));
  INV_X1    g129(.A(new_n228), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n315), .A2(new_n316), .ZN(new_n317));
  AOI21_X1  g131(.A(G902), .B1(new_n292), .B2(new_n308), .ZN(new_n318));
  AOI21_X1  g132(.A(new_n312), .B1(new_n317), .B2(new_n318), .ZN(new_n319));
  OAI21_X1  g133(.A(new_n187), .B1(new_n314), .B2(new_n319), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n320), .A2(KEYINPUT85), .ZN(new_n321));
  INV_X1    g135(.A(new_n187), .ZN(new_n322));
  OAI21_X1  g136(.A(new_n313), .B1(new_n295), .B2(new_n311), .ZN(new_n323));
  NAND3_X1  g137(.A1(new_n317), .A2(new_n318), .A3(new_n312), .ZN(new_n324));
  AOI21_X1  g138(.A(new_n322), .B1(new_n323), .B2(new_n324), .ZN(new_n325));
  INV_X1    g139(.A(KEYINPUT85), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  XNOR2_X1  g141(.A(KEYINPUT9), .B(G234), .ZN(new_n328));
  OAI21_X1  g142(.A(G221), .B1(new_n328), .B2(G902), .ZN(new_n329));
  XOR2_X1   g143(.A(new_n329), .B(KEYINPUT77), .Z(new_n330));
  INV_X1    g144(.A(G469), .ZN(new_n331));
  NOR2_X1   g145(.A1(new_n331), .A2(new_n310), .ZN(new_n332));
  OAI21_X1  g146(.A(KEYINPUT1), .B1(new_n203), .B2(G146), .ZN(new_n333));
  AOI21_X1  g147(.A(new_n221), .B1(G128), .B2(new_n333), .ZN(new_n334));
  OAI211_X1 g148(.A(new_n260), .B(new_n271), .C1(new_n334), .C2(new_n204), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n280), .A2(new_n274), .ZN(new_n336));
  INV_X1    g150(.A(new_n205), .ZN(new_n337));
  OAI21_X1  g151(.A(new_n335), .B1(new_n336), .B2(new_n337), .ZN(new_n338));
  INV_X1    g152(.A(KEYINPUT67), .ZN(new_n339));
  INV_X1    g153(.A(G137), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  AND2_X1   g155(.A1(KEYINPUT11), .A2(G134), .ZN(new_n342));
  NAND2_X1  g156(.A1(KEYINPUT67), .A2(G137), .ZN(new_n343));
  NAND3_X1  g157(.A1(new_n341), .A2(new_n342), .A3(new_n343), .ZN(new_n344));
  NAND2_X1  g158(.A1(KEYINPUT11), .A2(G134), .ZN(new_n345));
  NOR2_X1   g159(.A1(KEYINPUT11), .A2(G134), .ZN(new_n346));
  OAI21_X1  g160(.A(new_n345), .B1(new_n346), .B2(G137), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n344), .A2(new_n347), .ZN(new_n348));
  INV_X1    g162(.A(G131), .ZN(new_n349));
  NOR2_X1   g163(.A1(new_n349), .A2(KEYINPUT68), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n348), .A2(new_n350), .ZN(new_n351));
  INV_X1    g165(.A(new_n350), .ZN(new_n352));
  NAND3_X1  g166(.A1(new_n344), .A2(new_n347), .A3(new_n352), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n351), .A2(new_n353), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n338), .A2(new_n354), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n355), .A2(KEYINPUT12), .ZN(new_n356));
  INV_X1    g170(.A(KEYINPUT10), .ZN(new_n357));
  NOR2_X1   g171(.A1(new_n205), .A2(new_n357), .ZN(new_n358));
  AOI22_X1  g172(.A1(new_n336), .A2(new_n358), .B1(new_n357), .B2(new_n335), .ZN(new_n359));
  INV_X1    g173(.A(KEYINPUT70), .ZN(new_n360));
  AND3_X1   g174(.A1(new_n344), .A2(new_n352), .A3(new_n347), .ZN(new_n361));
  AOI21_X1  g175(.A(new_n352), .B1(new_n344), .B2(new_n347), .ZN(new_n362));
  OAI21_X1  g176(.A(new_n360), .B1(new_n361), .B2(new_n362), .ZN(new_n363));
  NAND3_X1  g177(.A1(new_n351), .A2(KEYINPUT70), .A3(new_n353), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n363), .A2(new_n364), .ZN(new_n365));
  OAI21_X1  g179(.A(new_n224), .B1(new_n261), .B2(new_n262), .ZN(new_n366));
  NAND3_X1  g180(.A1(new_n359), .A2(new_n365), .A3(new_n366), .ZN(new_n367));
  XNOR2_X1  g181(.A(G110), .B(G140), .ZN(new_n368));
  XNOR2_X1  g182(.A(new_n368), .B(KEYINPUT78), .ZN(new_n369));
  INV_X1    g183(.A(G227), .ZN(new_n370));
  NOR2_X1   g184(.A1(new_n370), .A2(G953), .ZN(new_n371));
  XOR2_X1   g185(.A(new_n369), .B(new_n371), .Z(new_n372));
  INV_X1    g186(.A(new_n372), .ZN(new_n373));
  INV_X1    g187(.A(KEYINPUT12), .ZN(new_n374));
  INV_X1    g188(.A(new_n365), .ZN(new_n375));
  NAND3_X1  g189(.A1(new_n338), .A2(new_n374), .A3(new_n375), .ZN(new_n376));
  NAND4_X1  g190(.A1(new_n356), .A2(new_n367), .A3(new_n373), .A4(new_n376), .ZN(new_n377));
  AND3_X1   g191(.A1(new_n359), .A2(new_n365), .A3(new_n366), .ZN(new_n378));
  AOI21_X1  g192(.A(new_n365), .B1(new_n359), .B2(new_n366), .ZN(new_n379));
  OAI21_X1  g193(.A(new_n372), .B1(new_n378), .B2(new_n379), .ZN(new_n380));
  AOI21_X1  g194(.A(G902), .B1(new_n377), .B2(new_n380), .ZN(new_n381));
  AOI21_X1  g195(.A(new_n332), .B1(new_n381), .B2(new_n331), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n367), .A2(new_n376), .ZN(new_n383));
  AOI21_X1  g197(.A(new_n374), .B1(new_n338), .B2(new_n354), .ZN(new_n384));
  OAI21_X1  g198(.A(new_n372), .B1(new_n383), .B2(new_n384), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n359), .A2(new_n366), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n386), .A2(new_n375), .ZN(new_n387));
  NAND3_X1  g201(.A1(new_n387), .A2(new_n367), .A3(new_n373), .ZN(new_n388));
  NAND3_X1  g202(.A1(new_n385), .A2(G469), .A3(new_n388), .ZN(new_n389));
  AOI21_X1  g203(.A(new_n330), .B1(new_n382), .B2(new_n389), .ZN(new_n390));
  INV_X1    g204(.A(new_n390), .ZN(new_n391));
  INV_X1    g205(.A(G237), .ZN(new_n392));
  NAND3_X1  g206(.A1(new_n392), .A2(new_n226), .A3(G214), .ZN(new_n393));
  NAND3_X1  g207(.A1(new_n393), .A2(new_n191), .A3(new_n193), .ZN(new_n394));
  NAND4_X1  g208(.A1(new_n392), .A2(new_n226), .A3(G143), .A4(G214), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n394), .A2(new_n395), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n396), .A2(G131), .ZN(new_n397));
  INV_X1    g211(.A(KEYINPUT86), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n397), .A2(new_n398), .ZN(new_n399));
  INV_X1    g213(.A(KEYINPUT17), .ZN(new_n400));
  NAND3_X1  g214(.A1(new_n396), .A2(KEYINPUT86), .A3(G131), .ZN(new_n401));
  NAND3_X1  g215(.A1(new_n394), .A2(new_n349), .A3(new_n395), .ZN(new_n402));
  NAND4_X1  g216(.A1(new_n399), .A2(new_n400), .A3(new_n401), .A4(new_n402), .ZN(new_n403));
  INV_X1    g217(.A(G140), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n404), .A2(G125), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n206), .A2(G140), .ZN(new_n406));
  NAND3_X1  g220(.A1(new_n405), .A2(new_n406), .A3(KEYINPUT16), .ZN(new_n407));
  OR3_X1    g221(.A1(new_n206), .A2(KEYINPUT16), .A3(G140), .ZN(new_n408));
  NAND3_X1  g222(.A1(new_n407), .A2(new_n408), .A3(G146), .ZN(new_n409));
  INV_X1    g223(.A(new_n409), .ZN(new_n410));
  AOI21_X1  g224(.A(G146), .B1(new_n407), .B2(new_n408), .ZN(new_n411));
  NOR2_X1   g225(.A1(new_n410), .A2(new_n411), .ZN(new_n412));
  AOI21_X1  g226(.A(KEYINPUT86), .B1(new_n396), .B2(G131), .ZN(new_n413));
  AOI211_X1 g227(.A(new_n398), .B(new_n349), .C1(new_n394), .C2(new_n395), .ZN(new_n414));
  OAI21_X1  g228(.A(KEYINPUT17), .B1(new_n413), .B2(new_n414), .ZN(new_n415));
  NAND3_X1  g229(.A1(new_n403), .A2(new_n412), .A3(new_n415), .ZN(new_n416));
  XNOR2_X1  g230(.A(G113), .B(G122), .ZN(new_n417));
  XNOR2_X1  g231(.A(new_n417), .B(new_n251), .ZN(new_n418));
  NAND2_X1  g232(.A1(KEYINPUT18), .A2(G131), .ZN(new_n419));
  XNOR2_X1  g233(.A(new_n396), .B(new_n419), .ZN(new_n420));
  AOI21_X1  g234(.A(KEYINPUT74), .B1(new_n405), .B2(new_n406), .ZN(new_n421));
  INV_X1    g235(.A(new_n421), .ZN(new_n422));
  XNOR2_X1  g236(.A(G125), .B(G140), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n423), .A2(KEYINPUT74), .ZN(new_n424));
  NAND3_X1  g238(.A1(new_n422), .A2(new_n424), .A3(new_n188), .ZN(new_n425));
  OAI21_X1  g239(.A(new_n425), .B1(new_n188), .B2(new_n423), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n420), .A2(new_n426), .ZN(new_n427));
  AND3_X1   g241(.A1(new_n416), .A2(new_n418), .A3(new_n427), .ZN(new_n428));
  AOI21_X1  g242(.A(new_n418), .B1(new_n416), .B2(new_n427), .ZN(new_n429));
  OAI21_X1  g243(.A(new_n310), .B1(new_n428), .B2(new_n429), .ZN(new_n430));
  INV_X1    g244(.A(KEYINPUT89), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  INV_X1    g246(.A(G475), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n416), .A2(new_n427), .ZN(new_n434));
  INV_X1    g248(.A(new_n418), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  NAND3_X1  g250(.A1(new_n416), .A2(new_n418), .A3(new_n427), .ZN(new_n437));
  AOI21_X1  g251(.A(G902), .B1(new_n436), .B2(new_n437), .ZN(new_n438));
  AOI21_X1  g252(.A(new_n433), .B1(new_n438), .B2(KEYINPUT89), .ZN(new_n439));
  NOR2_X1   g253(.A1(G475), .A2(G902), .ZN(new_n440));
  NAND3_X1  g254(.A1(new_n399), .A2(new_n401), .A3(new_n402), .ZN(new_n441));
  INV_X1    g255(.A(KEYINPUT87), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n441), .A2(new_n442), .ZN(new_n443));
  INV_X1    g257(.A(KEYINPUT88), .ZN(new_n444));
  INV_X1    g258(.A(KEYINPUT19), .ZN(new_n445));
  NAND4_X1  g259(.A1(new_n422), .A2(new_n424), .A3(new_n444), .A4(new_n445), .ZN(new_n446));
  AND3_X1   g260(.A1(new_n405), .A2(new_n406), .A3(KEYINPUT74), .ZN(new_n447));
  NOR3_X1   g261(.A1(new_n447), .A2(new_n421), .A3(KEYINPUT19), .ZN(new_n448));
  OAI21_X1  g262(.A(KEYINPUT88), .B1(new_n423), .B2(new_n445), .ZN(new_n449));
  OAI21_X1  g263(.A(new_n446), .B1(new_n448), .B2(new_n449), .ZN(new_n450));
  AOI21_X1  g264(.A(new_n410), .B1(new_n450), .B2(new_n188), .ZN(new_n451));
  NAND4_X1  g265(.A1(new_n399), .A2(KEYINPUT87), .A3(new_n401), .A4(new_n402), .ZN(new_n452));
  NAND3_X1  g266(.A1(new_n443), .A2(new_n451), .A3(new_n452), .ZN(new_n453));
  AOI21_X1  g267(.A(new_n418), .B1(new_n453), .B2(new_n427), .ZN(new_n454));
  OAI21_X1  g268(.A(new_n440), .B1(new_n454), .B2(new_n428), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n455), .A2(KEYINPUT20), .ZN(new_n456));
  INV_X1    g270(.A(KEYINPUT20), .ZN(new_n457));
  OAI211_X1 g271(.A(new_n457), .B(new_n440), .C1(new_n454), .C2(new_n428), .ZN(new_n458));
  AOI22_X1  g272(.A1(new_n432), .A2(new_n439), .B1(new_n456), .B2(new_n458), .ZN(new_n459));
  XOR2_X1   g273(.A(KEYINPUT21), .B(G898), .Z(new_n460));
  XNOR2_X1  g274(.A(new_n460), .B(KEYINPUT92), .ZN(new_n461));
  NAND2_X1  g275(.A1(G234), .A2(G237), .ZN(new_n462));
  AND3_X1   g276(.A1(new_n462), .A2(G902), .A3(G953), .ZN(new_n463));
  INV_X1    g277(.A(new_n463), .ZN(new_n464));
  NOR2_X1   g278(.A1(new_n461), .A2(new_n464), .ZN(new_n465));
  AND3_X1   g279(.A1(new_n462), .A2(G952), .A3(new_n226), .ZN(new_n466));
  NOR2_X1   g280(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  XNOR2_X1  g281(.A(new_n467), .B(KEYINPUT93), .ZN(new_n468));
  INV_X1    g282(.A(G122), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n469), .A2(G116), .ZN(new_n470));
  AOI21_X1  g284(.A(new_n249), .B1(new_n470), .B2(KEYINPUT14), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n234), .A2(G122), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n470), .A2(new_n472), .ZN(new_n473));
  OR2_X1    g287(.A1(new_n471), .A2(new_n473), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n471), .A2(new_n473), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  NOR2_X1   g290(.A1(new_n190), .A2(G128), .ZN(new_n477));
  AOI21_X1  g291(.A(new_n477), .B1(new_n203), .B2(G128), .ZN(new_n478));
  INV_X1    g292(.A(G134), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  OR2_X1    g294(.A1(new_n478), .A2(new_n479), .ZN(new_n481));
  AOI21_X1  g295(.A(new_n476), .B1(new_n480), .B2(new_n481), .ZN(new_n482));
  INV_X1    g296(.A(new_n482), .ZN(new_n483));
  INV_X1    g297(.A(KEYINPUT13), .ZN(new_n484));
  NAND4_X1  g298(.A1(new_n191), .A2(new_n193), .A3(new_n484), .A4(G128), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n485), .A2(G134), .ZN(new_n486));
  INV_X1    g300(.A(new_n486), .ZN(new_n487));
  NAND3_X1  g301(.A1(new_n191), .A2(new_n193), .A3(G128), .ZN(new_n488));
  INV_X1    g302(.A(new_n477), .ZN(new_n489));
  NAND3_X1  g303(.A1(new_n488), .A2(KEYINPUT13), .A3(new_n489), .ZN(new_n490));
  AOI22_X1  g304(.A1(new_n487), .A2(new_n490), .B1(new_n479), .B2(new_n478), .ZN(new_n491));
  INV_X1    g305(.A(KEYINPUT90), .ZN(new_n492));
  AND3_X1   g306(.A1(new_n470), .A2(new_n472), .A3(new_n492), .ZN(new_n493));
  AOI21_X1  g307(.A(new_n492), .B1(new_n470), .B2(new_n472), .ZN(new_n494));
  OAI21_X1  g308(.A(G107), .B1(new_n493), .B2(new_n494), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n473), .A2(KEYINPUT90), .ZN(new_n496));
  NAND3_X1  g310(.A1(new_n470), .A2(new_n472), .A3(new_n492), .ZN(new_n497));
  NAND3_X1  g311(.A1(new_n496), .A2(new_n497), .A3(new_n249), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n495), .A2(new_n498), .ZN(new_n499));
  AND3_X1   g313(.A1(new_n491), .A2(KEYINPUT91), .A3(new_n499), .ZN(new_n500));
  AOI21_X1  g314(.A(KEYINPUT91), .B1(new_n491), .B2(new_n499), .ZN(new_n501));
  OAI21_X1  g315(.A(new_n483), .B1(new_n500), .B2(new_n501), .ZN(new_n502));
  INV_X1    g316(.A(G217), .ZN(new_n503));
  NOR3_X1   g317(.A1(new_n328), .A2(new_n503), .A3(G953), .ZN(new_n504));
  INV_X1    g318(.A(new_n504), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n502), .A2(new_n505), .ZN(new_n506));
  INV_X1    g320(.A(KEYINPUT91), .ZN(new_n507));
  AND2_X1   g321(.A1(new_n495), .A2(new_n498), .ZN(new_n508));
  INV_X1    g322(.A(new_n490), .ZN(new_n509));
  OAI21_X1  g323(.A(new_n480), .B1(new_n509), .B2(new_n486), .ZN(new_n510));
  OAI21_X1  g324(.A(new_n507), .B1(new_n508), .B2(new_n510), .ZN(new_n511));
  NAND3_X1  g325(.A1(new_n491), .A2(KEYINPUT91), .A3(new_n499), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  NAND3_X1  g327(.A1(new_n513), .A2(new_n483), .A3(new_n504), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n506), .A2(new_n514), .ZN(new_n515));
  INV_X1    g329(.A(G478), .ZN(new_n516));
  OAI211_X1 g330(.A(new_n515), .B(new_n310), .C1(KEYINPUT15), .C2(new_n516), .ZN(new_n517));
  AOI21_X1  g331(.A(new_n504), .B1(new_n513), .B2(new_n483), .ZN(new_n518));
  AOI211_X1 g332(.A(new_n505), .B(new_n482), .C1(new_n511), .C2(new_n512), .ZN(new_n519));
  OAI21_X1  g333(.A(new_n310), .B1(new_n518), .B2(new_n519), .ZN(new_n520));
  NOR2_X1   g334(.A1(new_n516), .A2(KEYINPUT15), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n517), .A2(new_n522), .ZN(new_n523));
  INV_X1    g337(.A(new_n523), .ZN(new_n524));
  NAND3_X1  g338(.A1(new_n459), .A2(new_n468), .A3(new_n524), .ZN(new_n525));
  NOR2_X1   g339(.A1(new_n391), .A2(new_n525), .ZN(new_n526));
  INV_X1    g340(.A(KEYINPUT75), .ZN(new_n527));
  NOR2_X1   g341(.A1(new_n232), .A2(G128), .ZN(new_n528));
  AND2_X1   g342(.A1(KEYINPUT73), .A2(KEYINPUT23), .ZN(new_n529));
  NOR2_X1   g343(.A1(KEYINPUT73), .A2(KEYINPUT23), .ZN(new_n530));
  OAI21_X1  g344(.A(new_n528), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  INV_X1    g345(.A(G110), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n232), .A2(G128), .ZN(new_n533));
  NAND2_X1  g347(.A1(KEYINPUT73), .A2(KEYINPUT23), .ZN(new_n534));
  OAI21_X1  g348(.A(new_n534), .B1(new_n232), .B2(G128), .ZN(new_n535));
  NAND4_X1  g349(.A1(new_n531), .A2(new_n532), .A3(new_n533), .A4(new_n535), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n196), .A2(G119), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n537), .A2(new_n533), .ZN(new_n538));
  XNOR2_X1  g352(.A(KEYINPUT24), .B(G110), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n536), .A2(new_n540), .ZN(new_n541));
  NAND3_X1  g355(.A1(new_n541), .A2(new_n409), .A3(new_n425), .ZN(new_n542));
  INV_X1    g356(.A(new_n530), .ZN(new_n543));
  AOI21_X1  g357(.A(new_n537), .B1(new_n543), .B2(new_n534), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n535), .A2(new_n533), .ZN(new_n545));
  OAI21_X1  g359(.A(G110), .B1(new_n544), .B2(new_n545), .ZN(new_n546));
  OR2_X1    g360(.A1(new_n538), .A2(new_n539), .ZN(new_n547));
  OAI211_X1 g361(.A(new_n546), .B(new_n547), .C1(new_n410), .C2(new_n411), .ZN(new_n548));
  XNOR2_X1  g362(.A(KEYINPUT22), .B(G137), .ZN(new_n549));
  NAND3_X1  g363(.A1(new_n226), .A2(G221), .A3(G234), .ZN(new_n550));
  XNOR2_X1  g364(.A(new_n549), .B(new_n550), .ZN(new_n551));
  AND3_X1   g365(.A1(new_n542), .A2(new_n548), .A3(new_n551), .ZN(new_n552));
  AOI21_X1  g366(.A(new_n551), .B1(new_n542), .B2(new_n548), .ZN(new_n553));
  NOR3_X1   g367(.A1(new_n552), .A2(new_n553), .A3(G902), .ZN(new_n554));
  OAI21_X1  g368(.A(new_n527), .B1(new_n554), .B2(KEYINPUT25), .ZN(new_n555));
  INV_X1    g369(.A(KEYINPUT76), .ZN(new_n556));
  NAND3_X1  g370(.A1(new_n554), .A2(new_n556), .A3(KEYINPUT25), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n542), .A2(new_n548), .ZN(new_n558));
  INV_X1    g372(.A(new_n551), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  NAND3_X1  g374(.A1(new_n542), .A2(new_n548), .A3(new_n551), .ZN(new_n561));
  NAND4_X1  g375(.A1(new_n560), .A2(KEYINPUT25), .A3(new_n310), .A4(new_n561), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n562), .A2(KEYINPUT76), .ZN(new_n563));
  NAND3_X1  g377(.A1(new_n560), .A2(new_n310), .A3(new_n561), .ZN(new_n564));
  INV_X1    g378(.A(KEYINPUT25), .ZN(new_n565));
  NAND3_X1  g379(.A1(new_n564), .A2(KEYINPUT75), .A3(new_n565), .ZN(new_n566));
  NAND4_X1  g380(.A1(new_n555), .A2(new_n557), .A3(new_n563), .A4(new_n566), .ZN(new_n567));
  AOI21_X1  g381(.A(new_n503), .B1(G234), .B2(new_n310), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  NOR2_X1   g383(.A1(new_n552), .A2(new_n553), .ZN(new_n570));
  NOR2_X1   g384(.A1(new_n568), .A2(G902), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  AND2_X1   g386(.A1(new_n569), .A2(new_n572), .ZN(new_n573));
  INV_X1    g387(.A(new_n573), .ZN(new_n574));
  NAND3_X1  g388(.A1(new_n344), .A2(new_n347), .A3(new_n349), .ZN(new_n575));
  NAND3_X1  g389(.A1(new_n341), .A2(new_n479), .A3(new_n343), .ZN(new_n576));
  OAI211_X1 g390(.A(new_n576), .B(G131), .C1(new_n479), .C2(new_n340), .ZN(new_n577));
  OAI211_X1 g391(.A(new_n575), .B(new_n577), .C1(new_n200), .C2(new_n204), .ZN(new_n578));
  OAI211_X1 g392(.A(new_n578), .B(new_n243), .C1(new_n365), .C2(new_n223), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n579), .A2(KEYINPUT28), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n215), .A2(new_n218), .ZN(new_n581));
  AOI22_X1  g395(.A1(new_n581), .A2(KEYINPUT66), .B1(new_n216), .B2(new_n221), .ZN(new_n582));
  NAND4_X1  g396(.A1(new_n582), .A2(new_n220), .A3(new_n364), .A4(new_n363), .ZN(new_n583));
  INV_X1    g397(.A(KEYINPUT28), .ZN(new_n584));
  NAND4_X1  g398(.A1(new_n583), .A2(new_n584), .A3(new_n578), .A4(new_n243), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n580), .A2(new_n585), .ZN(new_n586));
  NAND4_X1  g400(.A1(new_n354), .A2(new_n213), .A3(new_n220), .A4(new_n222), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n587), .A2(new_n578), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n588), .A2(new_n244), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n586), .A2(new_n589), .ZN(new_n590));
  XNOR2_X1  g404(.A(KEYINPUT71), .B(KEYINPUT27), .ZN(new_n591));
  INV_X1    g405(.A(G210), .ZN(new_n592));
  NOR3_X1   g406(.A1(new_n592), .A2(G237), .A3(G953), .ZN(new_n593));
  XNOR2_X1  g407(.A(new_n591), .B(new_n593), .ZN(new_n594));
  XNOR2_X1  g408(.A(KEYINPUT26), .B(G101), .ZN(new_n595));
  XNOR2_X1  g409(.A(new_n594), .B(new_n595), .ZN(new_n596));
  INV_X1    g410(.A(new_n596), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n590), .A2(new_n597), .ZN(new_n598));
  INV_X1    g412(.A(KEYINPUT30), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n588), .A2(new_n599), .ZN(new_n600));
  OAI211_X1 g414(.A(KEYINPUT30), .B(new_n578), .C1(new_n365), .C2(new_n223), .ZN(new_n601));
  NAND3_X1  g415(.A1(new_n600), .A2(new_n244), .A3(new_n601), .ZN(new_n602));
  NAND3_X1  g416(.A1(new_n602), .A2(new_n579), .A3(new_n596), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n603), .A2(KEYINPUT31), .ZN(new_n604));
  XOR2_X1   g418(.A(KEYINPUT72), .B(KEYINPUT31), .Z(new_n605));
  NAND4_X1  g419(.A1(new_n602), .A2(new_n579), .A3(new_n596), .A4(new_n605), .ZN(new_n606));
  NAND3_X1  g420(.A1(new_n598), .A2(new_n604), .A3(new_n606), .ZN(new_n607));
  NOR2_X1   g421(.A1(G472), .A2(G902), .ZN(new_n608));
  AND3_X1   g422(.A1(new_n607), .A2(KEYINPUT32), .A3(new_n608), .ZN(new_n609));
  AOI21_X1  g423(.A(KEYINPUT32), .B1(new_n607), .B2(new_n608), .ZN(new_n610));
  NOR2_X1   g424(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  NOR2_X1   g425(.A1(new_n590), .A2(new_n597), .ZN(new_n612));
  AOI21_X1  g426(.A(new_n596), .B1(new_n602), .B2(new_n579), .ZN(new_n613));
  NOR3_X1   g427(.A1(new_n612), .A2(KEYINPUT29), .A3(new_n613), .ZN(new_n614));
  AOI21_X1  g428(.A(new_n243), .B1(new_n583), .B2(new_n578), .ZN(new_n615));
  AOI21_X1  g429(.A(new_n615), .B1(new_n580), .B2(new_n585), .ZN(new_n616));
  NAND3_X1  g430(.A1(new_n616), .A2(KEYINPUT29), .A3(new_n596), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n617), .A2(new_n310), .ZN(new_n618));
  OAI21_X1  g432(.A(G472), .B1(new_n614), .B2(new_n618), .ZN(new_n619));
  AOI21_X1  g433(.A(new_n574), .B1(new_n611), .B2(new_n619), .ZN(new_n620));
  NAND4_X1  g434(.A1(new_n321), .A2(new_n327), .A3(new_n526), .A4(new_n620), .ZN(new_n621));
  XNOR2_X1  g435(.A(new_n621), .B(G101), .ZN(G3));
  INV_X1    g436(.A(new_n468), .ZN(new_n623));
  NOR2_X1   g437(.A1(new_n320), .A2(new_n623), .ZN(new_n624));
  OAI21_X1  g438(.A(KEYINPUT33), .B1(new_n518), .B2(new_n519), .ZN(new_n625));
  INV_X1    g439(.A(KEYINPUT33), .ZN(new_n626));
  NAND3_X1  g440(.A1(new_n506), .A2(new_n626), .A3(new_n514), .ZN(new_n627));
  NAND3_X1  g441(.A1(new_n625), .A2(new_n627), .A3(G478), .ZN(new_n628));
  NAND3_X1  g442(.A1(new_n515), .A2(new_n516), .A3(new_n310), .ZN(new_n629));
  NAND2_X1  g443(.A1(G478), .A2(G902), .ZN(new_n630));
  NAND3_X1  g444(.A1(new_n628), .A2(new_n629), .A3(new_n630), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n438), .A2(KEYINPUT89), .ZN(new_n632));
  NAND3_X1  g446(.A1(new_n632), .A2(new_n432), .A3(G475), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n456), .A2(new_n458), .ZN(new_n634));
  AOI21_X1  g448(.A(new_n631), .B1(new_n633), .B2(new_n634), .ZN(new_n635));
  NAND2_X1  g449(.A1(new_n607), .A2(new_n310), .ZN(new_n636));
  NAND2_X1  g450(.A1(KEYINPUT94), .A2(G472), .ZN(new_n637));
  XNOR2_X1  g451(.A(new_n636), .B(new_n637), .ZN(new_n638));
  AND3_X1   g452(.A1(new_n638), .A2(new_n390), .A3(new_n573), .ZN(new_n639));
  NAND3_X1  g453(.A1(new_n624), .A2(new_n635), .A3(new_n639), .ZN(new_n640));
  XOR2_X1   g454(.A(KEYINPUT34), .B(G104), .Z(new_n641));
  XNOR2_X1  g455(.A(new_n640), .B(new_n641), .ZN(G6));
  NAND2_X1  g456(.A1(new_n634), .A2(new_n633), .ZN(new_n643));
  NOR2_X1   g457(.A1(new_n643), .A2(new_n524), .ZN(new_n644));
  NAND3_X1  g458(.A1(new_n624), .A2(new_n639), .A3(new_n644), .ZN(new_n645));
  XNOR2_X1  g459(.A(new_n645), .B(G107), .ZN(new_n646));
  XOR2_X1   g460(.A(KEYINPUT95), .B(KEYINPUT35), .Z(new_n647));
  XNOR2_X1  g461(.A(new_n646), .B(new_n647), .ZN(G9));
  INV_X1    g462(.A(new_n637), .ZN(new_n649));
  XNOR2_X1  g463(.A(new_n636), .B(new_n649), .ZN(new_n650));
  INV_X1    g464(.A(KEYINPUT97), .ZN(new_n651));
  NOR2_X1   g465(.A1(new_n559), .A2(KEYINPUT36), .ZN(new_n652));
  XNOR2_X1  g466(.A(new_n558), .B(new_n652), .ZN(new_n653));
  NAND2_X1  g467(.A1(new_n653), .A2(new_n571), .ZN(new_n654));
  AOI21_X1  g468(.A(KEYINPUT96), .B1(new_n569), .B2(new_n654), .ZN(new_n655));
  INV_X1    g469(.A(KEYINPUT96), .ZN(new_n656));
  INV_X1    g470(.A(new_n654), .ZN(new_n657));
  AOI211_X1 g471(.A(new_n656), .B(new_n657), .C1(new_n567), .C2(new_n568), .ZN(new_n658));
  OAI21_X1  g472(.A(new_n651), .B1(new_n655), .B2(new_n658), .ZN(new_n659));
  INV_X1    g473(.A(new_n568), .ZN(new_n660));
  AND3_X1   g474(.A1(new_n564), .A2(KEYINPUT75), .A3(new_n565), .ZN(new_n661));
  AOI21_X1  g475(.A(KEYINPUT75), .B1(new_n564), .B2(new_n565), .ZN(new_n662));
  NOR2_X1   g476(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  XNOR2_X1  g477(.A(new_n562), .B(new_n556), .ZN(new_n664));
  AOI21_X1  g478(.A(new_n660), .B1(new_n663), .B2(new_n664), .ZN(new_n665));
  OAI21_X1  g479(.A(new_n656), .B1(new_n665), .B2(new_n657), .ZN(new_n666));
  NAND3_X1  g480(.A1(new_n569), .A2(KEYINPUT96), .A3(new_n654), .ZN(new_n667));
  NAND3_X1  g481(.A1(new_n666), .A2(KEYINPUT97), .A3(new_n667), .ZN(new_n668));
  AOI21_X1  g482(.A(new_n650), .B1(new_n659), .B2(new_n668), .ZN(new_n669));
  NAND4_X1  g483(.A1(new_n321), .A2(new_n327), .A3(new_n526), .A4(new_n669), .ZN(new_n670));
  XOR2_X1   g484(.A(KEYINPUT37), .B(G110), .Z(new_n671));
  XNOR2_X1  g485(.A(new_n670), .B(new_n671), .ZN(G12));
  AOI22_X1  g486(.A1(new_n659), .A2(new_n668), .B1(new_n611), .B2(new_n619), .ZN(new_n673));
  INV_X1    g487(.A(G900), .ZN(new_n674));
  AOI21_X1  g488(.A(new_n466), .B1(new_n463), .B2(new_n674), .ZN(new_n675));
  INV_X1    g489(.A(new_n675), .ZN(new_n676));
  NAND4_X1  g490(.A1(new_n634), .A2(new_n633), .A3(new_n523), .A4(new_n676), .ZN(new_n677));
  INV_X1    g491(.A(KEYINPUT98), .ZN(new_n678));
  NAND2_X1  g492(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  NAND4_X1  g493(.A1(new_n459), .A2(KEYINPUT98), .A3(new_n523), .A4(new_n676), .ZN(new_n680));
  AND2_X1   g494(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  NAND4_X1  g495(.A1(new_n673), .A2(new_n325), .A3(new_n390), .A4(new_n681), .ZN(new_n682));
  XNOR2_X1  g496(.A(new_n682), .B(G128), .ZN(G30));
  XOR2_X1   g497(.A(new_n675), .B(KEYINPUT39), .Z(new_n684));
  NAND2_X1  g498(.A1(new_n390), .A2(new_n684), .ZN(new_n685));
  XNOR2_X1  g499(.A(new_n685), .B(KEYINPUT40), .ZN(new_n686));
  NAND2_X1  g500(.A1(new_n323), .A2(new_n324), .ZN(new_n687));
  XNOR2_X1  g501(.A(KEYINPUT99), .B(KEYINPUT38), .ZN(new_n688));
  XNOR2_X1  g502(.A(new_n687), .B(new_n688), .ZN(new_n689));
  NAND2_X1  g503(.A1(new_n666), .A2(new_n667), .ZN(new_n690));
  NAND2_X1  g504(.A1(new_n643), .A2(new_n523), .ZN(new_n691));
  OR3_X1    g505(.A1(new_n690), .A2(new_n691), .A3(new_n322), .ZN(new_n692));
  NAND2_X1  g506(.A1(new_n607), .A2(new_n608), .ZN(new_n693));
  INV_X1    g507(.A(KEYINPUT32), .ZN(new_n694));
  NAND2_X1  g508(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  NAND3_X1  g509(.A1(new_n607), .A2(KEYINPUT32), .A3(new_n608), .ZN(new_n696));
  AOI21_X1  g510(.A(new_n597), .B1(new_n602), .B2(new_n579), .ZN(new_n697));
  NAND2_X1  g511(.A1(new_n579), .A2(new_n597), .ZN(new_n698));
  OAI21_X1  g512(.A(new_n310), .B1(new_n698), .B2(new_n615), .ZN(new_n699));
  OAI21_X1  g513(.A(G472), .B1(new_n697), .B2(new_n699), .ZN(new_n700));
  NAND3_X1  g514(.A1(new_n695), .A2(new_n696), .A3(new_n700), .ZN(new_n701));
  NAND2_X1  g515(.A1(new_n701), .A2(KEYINPUT100), .ZN(new_n702));
  INV_X1    g516(.A(KEYINPUT100), .ZN(new_n703));
  NAND4_X1  g517(.A1(new_n695), .A2(new_n703), .A3(new_n696), .A4(new_n700), .ZN(new_n704));
  NAND2_X1  g518(.A1(new_n702), .A2(new_n704), .ZN(new_n705));
  INV_X1    g519(.A(new_n705), .ZN(new_n706));
  NOR4_X1   g520(.A1(new_n686), .A2(new_n689), .A3(new_n692), .A4(new_n706), .ZN(new_n707));
  XNOR2_X1  g521(.A(new_n707), .B(new_n203), .ZN(G45));
  INV_X1    g522(.A(new_n631), .ZN(new_n709));
  NAND3_X1  g523(.A1(new_n643), .A2(new_n709), .A3(new_n676), .ZN(new_n710));
  INV_X1    g524(.A(new_n710), .ZN(new_n711));
  NAND4_X1  g525(.A1(new_n673), .A2(new_n325), .A3(new_n390), .A4(new_n711), .ZN(new_n712));
  XNOR2_X1  g526(.A(new_n712), .B(G146), .ZN(G48));
  NOR2_X1   g527(.A1(new_n381), .A2(new_n331), .ZN(new_n714));
  AOI211_X1 g528(.A(G469), .B(G902), .C1(new_n377), .C2(new_n380), .ZN(new_n715));
  INV_X1    g529(.A(new_n329), .ZN(new_n716));
  NOR3_X1   g530(.A1(new_n714), .A2(new_n715), .A3(new_n716), .ZN(new_n717));
  NAND3_X1  g531(.A1(new_n619), .A2(new_n695), .A3(new_n696), .ZN(new_n718));
  AND3_X1   g532(.A1(new_n717), .A2(new_n718), .A3(new_n573), .ZN(new_n719));
  NAND4_X1  g533(.A1(new_n719), .A2(new_n325), .A3(new_n468), .A4(new_n635), .ZN(new_n720));
  XNOR2_X1  g534(.A(KEYINPUT41), .B(G113), .ZN(new_n721));
  XNOR2_X1  g535(.A(new_n721), .B(KEYINPUT101), .ZN(new_n722));
  XNOR2_X1  g536(.A(new_n720), .B(new_n722), .ZN(G15));
  INV_X1    g537(.A(KEYINPUT102), .ZN(new_n724));
  NAND4_X1  g538(.A1(new_n624), .A2(new_n719), .A3(new_n724), .A4(new_n644), .ZN(new_n725));
  NAND3_X1  g539(.A1(new_n325), .A2(new_n468), .A3(new_n644), .ZN(new_n726));
  NAND2_X1  g540(.A1(new_n620), .A2(new_n717), .ZN(new_n727));
  OAI21_X1  g541(.A(KEYINPUT102), .B1(new_n726), .B2(new_n727), .ZN(new_n728));
  NAND2_X1  g542(.A1(new_n725), .A2(new_n728), .ZN(new_n729));
  XNOR2_X1  g543(.A(new_n729), .B(G116), .ZN(G18));
  AOI21_X1  g544(.A(new_n525), .B1(new_n659), .B2(new_n668), .ZN(new_n731));
  NAND4_X1  g545(.A1(new_n731), .A2(new_n325), .A3(new_n718), .A4(new_n717), .ZN(new_n732));
  XNOR2_X1  g546(.A(new_n732), .B(G119), .ZN(G21));
  INV_X1    g547(.A(new_n714), .ZN(new_n734));
  NAND2_X1  g548(.A1(new_n377), .A2(new_n380), .ZN(new_n735));
  NAND3_X1  g549(.A1(new_n735), .A2(new_n331), .A3(new_n310), .ZN(new_n736));
  NAND4_X1  g550(.A1(new_n734), .A2(new_n468), .A3(new_n736), .A4(new_n329), .ZN(new_n737));
  NAND2_X1  g551(.A1(new_n636), .A2(G472), .ZN(new_n738));
  OAI211_X1 g552(.A(new_n604), .B(new_n606), .C1(new_n616), .C2(new_n596), .ZN(new_n739));
  NAND2_X1  g553(.A1(new_n739), .A2(new_n608), .ZN(new_n740));
  NAND3_X1  g554(.A1(new_n738), .A2(new_n573), .A3(new_n740), .ZN(new_n741));
  NOR2_X1   g555(.A1(new_n737), .A2(new_n741), .ZN(new_n742));
  INV_X1    g556(.A(KEYINPUT103), .ZN(new_n743));
  XNOR2_X1  g557(.A(new_n691), .B(new_n743), .ZN(new_n744));
  NAND3_X1  g558(.A1(new_n742), .A2(new_n744), .A3(new_n325), .ZN(new_n745));
  XNOR2_X1  g559(.A(new_n745), .B(G122), .ZN(G24));
  INV_X1    g560(.A(KEYINPUT104), .ZN(new_n747));
  AOI21_X1  g561(.A(new_n747), .B1(new_n635), .B2(new_n676), .ZN(new_n748));
  NOR4_X1   g562(.A1(new_n459), .A2(KEYINPUT104), .A3(new_n631), .A4(new_n675), .ZN(new_n749));
  NOR2_X1   g563(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  AND3_X1   g564(.A1(new_n690), .A2(new_n740), .A3(new_n738), .ZN(new_n751));
  NAND4_X1  g565(.A1(new_n750), .A2(new_n325), .A3(new_n751), .A4(new_n717), .ZN(new_n752));
  XNOR2_X1  g566(.A(new_n752), .B(G125), .ZN(G27));
  AND3_X1   g567(.A1(new_n323), .A2(new_n324), .A3(new_n187), .ZN(new_n754));
  NAND2_X1  g568(.A1(new_n388), .A2(KEYINPUT105), .ZN(new_n755));
  INV_X1    g569(.A(KEYINPUT105), .ZN(new_n756));
  NAND4_X1  g570(.A1(new_n387), .A2(new_n756), .A3(new_n367), .A4(new_n373), .ZN(new_n757));
  NAND4_X1  g571(.A1(new_n755), .A2(G469), .A3(new_n385), .A4(new_n757), .ZN(new_n758));
  INV_X1    g572(.A(new_n332), .ZN(new_n759));
  NAND3_X1  g573(.A1(new_n758), .A2(new_n736), .A3(new_n759), .ZN(new_n760));
  NAND2_X1  g574(.A1(new_n760), .A2(new_n329), .ZN(new_n761));
  INV_X1    g575(.A(new_n761), .ZN(new_n762));
  NAND4_X1  g576(.A1(new_n750), .A2(new_n754), .A3(new_n620), .A4(new_n762), .ZN(new_n763));
  INV_X1    g577(.A(KEYINPUT42), .ZN(new_n764));
  NAND2_X1  g578(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  NAND3_X1  g579(.A1(new_n323), .A2(new_n324), .A3(new_n187), .ZN(new_n766));
  NOR2_X1   g580(.A1(new_n766), .A2(new_n761), .ZN(new_n767));
  NAND4_X1  g581(.A1(new_n767), .A2(KEYINPUT42), .A3(new_n620), .A4(new_n750), .ZN(new_n768));
  NAND2_X1  g582(.A1(new_n765), .A2(new_n768), .ZN(new_n769));
  XNOR2_X1  g583(.A(new_n769), .B(G131), .ZN(G33));
  NAND3_X1  g584(.A1(new_n767), .A2(new_n620), .A3(new_n681), .ZN(new_n771));
  XNOR2_X1  g585(.A(new_n771), .B(G134), .ZN(G36));
  NAND2_X1  g586(.A1(new_n459), .A2(new_n709), .ZN(new_n773));
  XNOR2_X1  g587(.A(new_n773), .B(KEYINPUT43), .ZN(new_n774));
  NAND2_X1  g588(.A1(new_n650), .A2(new_n690), .ZN(new_n775));
  NOR2_X1   g589(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  OR2_X1    g590(.A1(new_n776), .A2(KEYINPUT44), .ZN(new_n777));
  NAND2_X1  g591(.A1(new_n776), .A2(KEYINPUT44), .ZN(new_n778));
  AND3_X1   g592(.A1(new_n777), .A2(new_n754), .A3(new_n778), .ZN(new_n779));
  NAND4_X1  g593(.A1(new_n755), .A2(KEYINPUT45), .A3(new_n385), .A4(new_n757), .ZN(new_n780));
  AND2_X1   g594(.A1(new_n385), .A2(new_n388), .ZN(new_n781));
  OAI211_X1 g595(.A(new_n780), .B(G469), .C1(KEYINPUT45), .C2(new_n781), .ZN(new_n782));
  NAND3_X1  g596(.A1(new_n782), .A2(KEYINPUT46), .A3(new_n759), .ZN(new_n783));
  XOR2_X1   g597(.A(new_n783), .B(KEYINPUT106), .Z(new_n784));
  AOI21_X1  g598(.A(KEYINPUT46), .B1(new_n782), .B2(new_n759), .ZN(new_n785));
  NOR2_X1   g599(.A1(new_n785), .A2(new_n715), .ZN(new_n786));
  AOI21_X1  g600(.A(new_n716), .B1(new_n784), .B2(new_n786), .ZN(new_n787));
  NAND3_X1  g601(.A1(new_n779), .A2(new_n684), .A3(new_n787), .ZN(new_n788));
  XNOR2_X1  g602(.A(new_n788), .B(G137), .ZN(G39));
  NOR4_X1   g603(.A1(new_n766), .A2(new_n718), .A3(new_n573), .A4(new_n710), .ZN(new_n790));
  NOR2_X1   g604(.A1(new_n787), .A2(KEYINPUT47), .ZN(new_n791));
  INV_X1    g605(.A(KEYINPUT47), .ZN(new_n792));
  AOI211_X1 g606(.A(new_n792), .B(new_n716), .C1(new_n784), .C2(new_n786), .ZN(new_n793));
  OAI21_X1  g607(.A(new_n790), .B1(new_n791), .B2(new_n793), .ZN(new_n794));
  XNOR2_X1  g608(.A(new_n794), .B(G140), .ZN(G42));
  NAND3_X1  g609(.A1(new_n569), .A2(new_n654), .A3(new_n676), .ZN(new_n796));
  NOR2_X1   g610(.A1(new_n761), .A2(new_n796), .ZN(new_n797));
  NAND4_X1  g611(.A1(new_n705), .A2(new_n744), .A3(new_n797), .A4(new_n325), .ZN(new_n798));
  NAND4_X1  g612(.A1(new_n798), .A2(new_n682), .A3(new_n712), .A4(new_n752), .ZN(new_n799));
  INV_X1    g613(.A(KEYINPUT110), .ZN(new_n800));
  NAND2_X1  g614(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  NOR3_X1   g615(.A1(new_n655), .A2(new_n658), .A3(new_n651), .ZN(new_n802));
  AOI21_X1  g616(.A(KEYINPUT97), .B1(new_n666), .B2(new_n667), .ZN(new_n803));
  OAI211_X1 g617(.A(new_n718), .B(new_n390), .C1(new_n802), .C2(new_n803), .ZN(new_n804));
  INV_X1    g618(.A(new_n804), .ZN(new_n805));
  OAI211_X1 g619(.A(new_n805), .B(new_n325), .C1(new_n681), .C2(new_n711), .ZN(new_n806));
  NAND4_X1  g620(.A1(new_n806), .A2(KEYINPUT110), .A3(new_n752), .A4(new_n798), .ZN(new_n807));
  AND3_X1   g621(.A1(new_n801), .A2(new_n807), .A3(KEYINPUT52), .ZN(new_n808));
  AOI21_X1  g622(.A(KEYINPUT52), .B1(new_n801), .B2(new_n807), .ZN(new_n809));
  OAI21_X1  g623(.A(KEYINPUT111), .B1(new_n808), .B2(new_n809), .ZN(new_n810));
  INV_X1    g624(.A(KEYINPUT52), .ZN(new_n811));
  NAND4_X1  g625(.A1(new_n687), .A2(new_n187), .A3(new_n679), .A4(new_n680), .ZN(new_n812));
  NAND3_X1  g626(.A1(new_n687), .A2(new_n187), .A3(new_n711), .ZN(new_n813));
  AOI21_X1  g627(.A(new_n804), .B1(new_n812), .B2(new_n813), .ZN(new_n814));
  NAND2_X1  g628(.A1(new_n325), .A2(new_n717), .ZN(new_n815));
  NAND2_X1  g629(.A1(new_n710), .A2(KEYINPUT104), .ZN(new_n816));
  AND2_X1   g630(.A1(new_n738), .A2(new_n740), .ZN(new_n817));
  NAND3_X1  g631(.A1(new_n635), .A2(new_n747), .A3(new_n676), .ZN(new_n818));
  NAND4_X1  g632(.A1(new_n816), .A2(new_n817), .A3(new_n818), .A4(new_n690), .ZN(new_n819));
  NOR2_X1   g633(.A1(new_n815), .A2(new_n819), .ZN(new_n820));
  NOR2_X1   g634(.A1(new_n814), .A2(new_n820), .ZN(new_n821));
  AOI21_X1  g635(.A(KEYINPUT110), .B1(new_n821), .B2(new_n798), .ZN(new_n822));
  NOR2_X1   g636(.A1(new_n799), .A2(new_n800), .ZN(new_n823));
  OAI21_X1  g637(.A(new_n811), .B1(new_n822), .B2(new_n823), .ZN(new_n824));
  INV_X1    g638(.A(KEYINPUT111), .ZN(new_n825));
  NAND3_X1  g639(.A1(new_n801), .A2(new_n807), .A3(KEYINPUT52), .ZN(new_n826));
  NAND3_X1  g640(.A1(new_n824), .A2(new_n825), .A3(new_n826), .ZN(new_n827));
  AND3_X1   g641(.A1(new_n720), .A2(new_n732), .A3(new_n745), .ZN(new_n828));
  NAND3_X1  g642(.A1(new_n828), .A2(new_n729), .A3(new_n769), .ZN(new_n829));
  INV_X1    g643(.A(KEYINPUT107), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n523), .A2(new_n830), .ZN(new_n831));
  NAND3_X1  g645(.A1(new_n517), .A2(new_n522), .A3(KEYINPUT107), .ZN(new_n832));
  NAND2_X1  g646(.A1(new_n831), .A2(new_n832), .ZN(new_n833));
  NAND2_X1  g647(.A1(new_n833), .A2(new_n459), .ZN(new_n834));
  NAND2_X1  g648(.A1(new_n643), .A2(new_n709), .ZN(new_n835));
  AOI21_X1  g649(.A(new_n623), .B1(new_n834), .B2(new_n835), .ZN(new_n836));
  NAND4_X1  g650(.A1(new_n321), .A2(new_n327), .A3(new_n639), .A4(new_n836), .ZN(new_n837));
  NAND3_X1  g651(.A1(new_n621), .A2(new_n670), .A3(new_n837), .ZN(new_n838));
  INV_X1    g652(.A(KEYINPUT108), .ZN(new_n839));
  AND4_X1   g653(.A1(new_n459), .A2(new_n831), .A3(new_n676), .A4(new_n832), .ZN(new_n840));
  NAND3_X1  g654(.A1(new_n754), .A2(new_n839), .A3(new_n840), .ZN(new_n841));
  NAND4_X1  g655(.A1(new_n840), .A2(new_n323), .A3(new_n187), .A4(new_n324), .ZN(new_n842));
  NAND2_X1  g656(.A1(new_n842), .A2(KEYINPUT108), .ZN(new_n843));
  NAND3_X1  g657(.A1(new_n841), .A2(new_n805), .A3(new_n843), .ZN(new_n844));
  NAND3_X1  g658(.A1(new_n767), .A2(new_n751), .A3(new_n750), .ZN(new_n845));
  NAND3_X1  g659(.A1(new_n844), .A2(new_n771), .A3(new_n845), .ZN(new_n846));
  NOR3_X1   g660(.A1(new_n829), .A2(new_n838), .A3(new_n846), .ZN(new_n847));
  NAND3_X1  g661(.A1(new_n810), .A2(new_n827), .A3(new_n847), .ZN(new_n848));
  NAND2_X1  g662(.A1(new_n848), .A2(KEYINPUT53), .ZN(new_n849));
  AOI21_X1  g663(.A(KEYINPUT53), .B1(new_n847), .B2(KEYINPUT109), .ZN(new_n850));
  NAND2_X1  g664(.A1(new_n799), .A2(KEYINPUT52), .ZN(new_n851));
  NAND2_X1  g665(.A1(new_n824), .A2(new_n851), .ZN(new_n852));
  INV_X1    g666(.A(new_n852), .ZN(new_n853));
  OAI211_X1 g667(.A(new_n850), .B(new_n853), .C1(KEYINPUT109), .C2(new_n847), .ZN(new_n854));
  AND2_X1   g668(.A1(new_n849), .A2(new_n854), .ZN(new_n855));
  NAND2_X1  g669(.A1(new_n855), .A2(KEYINPUT54), .ZN(new_n856));
  AND4_X1   g670(.A1(KEYINPUT53), .A2(new_n828), .A3(new_n729), .A4(new_n769), .ZN(new_n857));
  INV_X1    g671(.A(new_n846), .ZN(new_n858));
  AND3_X1   g672(.A1(new_n621), .A2(new_n670), .A3(new_n837), .ZN(new_n859));
  INV_X1    g673(.A(KEYINPUT112), .ZN(new_n860));
  NAND3_X1  g674(.A1(new_n858), .A2(new_n859), .A3(new_n860), .ZN(new_n861));
  OAI21_X1  g675(.A(KEYINPUT112), .B1(new_n838), .B2(new_n846), .ZN(new_n862));
  NAND3_X1  g676(.A1(new_n857), .A2(new_n861), .A3(new_n862), .ZN(new_n863));
  NOR2_X1   g677(.A1(new_n852), .A2(new_n863), .ZN(new_n864));
  INV_X1    g678(.A(KEYINPUT53), .ZN(new_n865));
  AOI21_X1  g679(.A(new_n864), .B1(new_n848), .B2(new_n865), .ZN(new_n866));
  INV_X1    g680(.A(new_n866), .ZN(new_n867));
  OAI21_X1  g681(.A(new_n856), .B1(KEYINPUT54), .B2(new_n867), .ZN(new_n868));
  INV_X1    g682(.A(KEYINPUT51), .ZN(new_n869));
  NOR2_X1   g683(.A1(new_n714), .A2(new_n715), .ZN(new_n870));
  AOI211_X1 g684(.A(new_n793), .B(new_n791), .C1(new_n330), .C2(new_n870), .ZN(new_n871));
  INV_X1    g685(.A(new_n466), .ZN(new_n872));
  OR2_X1    g686(.A1(new_n774), .A2(new_n872), .ZN(new_n873));
  NOR4_X1   g687(.A1(new_n871), .A2(new_n741), .A3(new_n766), .A4(new_n873), .ZN(new_n874));
  INV_X1    g688(.A(KEYINPUT50), .ZN(new_n875));
  NOR2_X1   g689(.A1(new_n873), .A2(new_n741), .ZN(new_n876));
  NAND4_X1  g690(.A1(new_n876), .A2(new_n322), .A3(new_n689), .A4(new_n717), .ZN(new_n877));
  INV_X1    g691(.A(KEYINPUT113), .ZN(new_n878));
  NOR2_X1   g692(.A1(new_n877), .A2(new_n878), .ZN(new_n879));
  OAI21_X1  g693(.A(new_n875), .B1(new_n879), .B2(KEYINPUT114), .ZN(new_n880));
  NAND2_X1  g694(.A1(new_n754), .A2(new_n717), .ZN(new_n881));
  OR4_X1    g695(.A1(new_n574), .A2(new_n881), .A3(new_n872), .A4(new_n705), .ZN(new_n882));
  OR3_X1    g696(.A1(new_n882), .A2(new_n643), .A3(new_n709), .ZN(new_n883));
  NOR2_X1   g697(.A1(new_n873), .A2(new_n881), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n884), .A2(new_n751), .ZN(new_n885));
  OAI21_X1  g699(.A(KEYINPUT113), .B1(new_n875), .B2(KEYINPUT114), .ZN(new_n886));
  NAND2_X1  g700(.A1(new_n877), .A2(new_n886), .ZN(new_n887));
  NAND4_X1  g701(.A1(new_n880), .A2(new_n883), .A3(new_n885), .A4(new_n887), .ZN(new_n888));
  OAI21_X1  g702(.A(new_n869), .B1(new_n874), .B2(new_n888), .ZN(new_n889));
  NAND2_X1  g703(.A1(new_n884), .A2(new_n620), .ZN(new_n890));
  XOR2_X1   g704(.A(new_n890), .B(KEYINPUT48), .Z(new_n891));
  INV_X1    g705(.A(G952), .ZN(new_n892));
  INV_X1    g706(.A(new_n815), .ZN(new_n893));
  AOI211_X1 g707(.A(new_n892), .B(G953), .C1(new_n876), .C2(new_n893), .ZN(new_n894));
  OAI21_X1  g708(.A(new_n894), .B1(new_n835), .B2(new_n882), .ZN(new_n895));
  NOR2_X1   g709(.A1(new_n891), .A2(new_n895), .ZN(new_n896));
  OR2_X1    g710(.A1(new_n874), .A2(new_n869), .ZN(new_n897));
  XOR2_X1   g711(.A(new_n888), .B(KEYINPUT115), .Z(new_n898));
  OAI211_X1 g712(.A(new_n889), .B(new_n896), .C1(new_n897), .C2(new_n898), .ZN(new_n899));
  OAI22_X1  g713(.A1(new_n868), .A2(new_n899), .B1(G952), .B2(G953), .ZN(new_n900));
  INV_X1    g714(.A(new_n870), .ZN(new_n901));
  AND2_X1   g715(.A1(new_n901), .A2(KEYINPUT49), .ZN(new_n902));
  NOR2_X1   g716(.A1(new_n901), .A2(KEYINPUT49), .ZN(new_n903));
  OR3_X1    g717(.A1(new_n574), .A2(new_n322), .A3(new_n330), .ZN(new_n904));
  NOR4_X1   g718(.A1(new_n902), .A2(new_n903), .A3(new_n904), .A4(new_n773), .ZN(new_n905));
  NAND3_X1  g719(.A1(new_n905), .A2(new_n689), .A3(new_n706), .ZN(new_n906));
  NAND2_X1  g720(.A1(new_n900), .A2(new_n906), .ZN(G75));
  INV_X1    g721(.A(KEYINPUT56), .ZN(new_n908));
  NAND2_X1  g722(.A1(new_n867), .A2(G902), .ZN(new_n909));
  OAI21_X1  g723(.A(new_n908), .B1(new_n909), .B2(new_n592), .ZN(new_n910));
  NOR2_X1   g724(.A1(new_n315), .A2(new_n316), .ZN(new_n911));
  NOR2_X1   g725(.A1(new_n911), .A2(new_n295), .ZN(new_n912));
  XNOR2_X1  g726(.A(KEYINPUT116), .B(KEYINPUT55), .ZN(new_n913));
  XOR2_X1   g727(.A(new_n912), .B(new_n913), .Z(new_n914));
  AND2_X1   g728(.A1(new_n910), .A2(new_n914), .ZN(new_n915));
  NOR2_X1   g729(.A1(new_n910), .A2(new_n914), .ZN(new_n916));
  NOR2_X1   g730(.A1(new_n226), .A2(G952), .ZN(new_n917));
  NOR3_X1   g731(.A1(new_n915), .A2(new_n916), .A3(new_n917), .ZN(G51));
  XNOR2_X1  g732(.A(new_n332), .B(KEYINPUT57), .ZN(new_n919));
  NOR2_X1   g733(.A1(new_n867), .A2(KEYINPUT54), .ZN(new_n920));
  INV_X1    g734(.A(KEYINPUT54), .ZN(new_n921));
  NOR2_X1   g735(.A1(new_n866), .A2(new_n921), .ZN(new_n922));
  OAI21_X1  g736(.A(new_n919), .B1(new_n920), .B2(new_n922), .ZN(new_n923));
  XOR2_X1   g737(.A(new_n735), .B(KEYINPUT117), .Z(new_n924));
  NAND2_X1  g738(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  OR2_X1    g739(.A1(new_n909), .A2(new_n782), .ZN(new_n926));
  AOI21_X1  g740(.A(new_n917), .B1(new_n925), .B2(new_n926), .ZN(G54));
  INV_X1    g741(.A(new_n909), .ZN(new_n928));
  NOR2_X1   g742(.A1(new_n454), .A2(new_n428), .ZN(new_n929));
  INV_X1    g743(.A(new_n929), .ZN(new_n930));
  AND2_X1   g744(.A1(KEYINPUT58), .A2(G475), .ZN(new_n931));
  AND3_X1   g745(.A1(new_n928), .A2(new_n930), .A3(new_n931), .ZN(new_n932));
  AOI21_X1  g746(.A(new_n930), .B1(new_n928), .B2(new_n931), .ZN(new_n933));
  NOR3_X1   g747(.A1(new_n932), .A2(new_n933), .A3(new_n917), .ZN(G60));
  AND2_X1   g748(.A1(new_n625), .A2(new_n627), .ZN(new_n935));
  INV_X1    g749(.A(new_n935), .ZN(new_n936));
  XNOR2_X1  g750(.A(new_n630), .B(KEYINPUT59), .ZN(new_n937));
  AOI21_X1  g751(.A(new_n936), .B1(new_n868), .B2(new_n937), .ZN(new_n938));
  OAI211_X1 g752(.A(new_n936), .B(new_n937), .C1(new_n920), .C2(new_n922), .ZN(new_n939));
  INV_X1    g753(.A(new_n917), .ZN(new_n940));
  NAND2_X1  g754(.A1(new_n939), .A2(new_n940), .ZN(new_n941));
  NOR2_X1   g755(.A1(new_n938), .A2(new_n941), .ZN(G63));
  XOR2_X1   g756(.A(new_n570), .B(KEYINPUT119), .Z(new_n943));
  XNOR2_X1  g757(.A(KEYINPUT118), .B(KEYINPUT60), .ZN(new_n944));
  NAND2_X1  g758(.A1(G217), .A2(G902), .ZN(new_n945));
  XNOR2_X1  g759(.A(new_n944), .B(new_n945), .ZN(new_n946));
  OAI21_X1  g760(.A(new_n943), .B1(new_n866), .B2(new_n946), .ZN(new_n947));
  OR2_X1    g761(.A1(new_n947), .A2(KEYINPUT121), .ZN(new_n948));
  NOR2_X1   g762(.A1(new_n866), .A2(new_n946), .ZN(new_n949));
  NAND2_X1  g763(.A1(new_n949), .A2(new_n653), .ZN(new_n950));
  NAND2_X1  g764(.A1(new_n947), .A2(KEYINPUT121), .ZN(new_n951));
  AND2_X1   g765(.A1(new_n940), .A2(KEYINPUT61), .ZN(new_n952));
  NAND4_X1  g766(.A1(new_n948), .A2(new_n950), .A3(new_n951), .A4(new_n952), .ZN(new_n953));
  INV_X1    g767(.A(KEYINPUT120), .ZN(new_n954));
  AND3_X1   g768(.A1(new_n947), .A2(new_n954), .A3(new_n940), .ZN(new_n955));
  AOI21_X1  g769(.A(new_n954), .B1(new_n947), .B2(new_n940), .ZN(new_n956));
  AND2_X1   g770(.A1(new_n949), .A2(new_n653), .ZN(new_n957));
  NOR3_X1   g771(.A1(new_n955), .A2(new_n956), .A3(new_n957), .ZN(new_n958));
  OAI21_X1  g772(.A(new_n953), .B1(new_n958), .B2(KEYINPUT61), .ZN(G66));
  AOI21_X1  g773(.A(new_n226), .B1(new_n461), .B2(G224), .ZN(new_n960));
  NAND3_X1  g774(.A1(new_n859), .A2(new_n729), .A3(new_n828), .ZN(new_n961));
  AOI21_X1  g775(.A(new_n960), .B1(new_n961), .B2(new_n226), .ZN(new_n962));
  INV_X1    g776(.A(G898), .ZN(new_n963));
  AOI21_X1  g777(.A(new_n315), .B1(new_n963), .B2(G953), .ZN(new_n964));
  XOR2_X1   g778(.A(new_n964), .B(KEYINPUT122), .Z(new_n965));
  XNOR2_X1  g779(.A(new_n962), .B(new_n965), .ZN(G69));
  OAI21_X1  g780(.A(G953), .B1(new_n370), .B2(new_n674), .ZN(new_n967));
  INV_X1    g781(.A(new_n967), .ZN(new_n968));
  NAND2_X1  g782(.A1(new_n784), .A2(new_n786), .ZN(new_n969));
  NAND2_X1  g783(.A1(new_n969), .A2(new_n329), .ZN(new_n970));
  NAND3_X1  g784(.A1(new_n777), .A2(new_n754), .A3(new_n778), .ZN(new_n971));
  INV_X1    g785(.A(new_n684), .ZN(new_n972));
  NOR3_X1   g786(.A1(new_n970), .A2(new_n971), .A3(new_n972), .ZN(new_n973));
  NAND2_X1  g787(.A1(new_n834), .A2(new_n835), .ZN(new_n974));
  NAND2_X1  g788(.A1(new_n620), .A2(new_n974), .ZN(new_n975));
  NOR3_X1   g789(.A1(new_n975), .A2(new_n685), .A3(new_n766), .ZN(new_n976));
  OR2_X1    g790(.A1(new_n976), .A2(KEYINPUT123), .ZN(new_n977));
  NAND2_X1  g791(.A1(new_n976), .A2(KEYINPUT123), .ZN(new_n978));
  NAND2_X1  g792(.A1(new_n977), .A2(new_n978), .ZN(new_n979));
  OAI21_X1  g793(.A(KEYINPUT124), .B1(new_n973), .B2(new_n979), .ZN(new_n980));
  INV_X1    g794(.A(KEYINPUT124), .ZN(new_n981));
  NAND4_X1  g795(.A1(new_n788), .A2(new_n981), .A3(new_n977), .A4(new_n978), .ZN(new_n982));
  NAND2_X1  g796(.A1(new_n980), .A2(new_n982), .ZN(new_n983));
  INV_X1    g797(.A(new_n821), .ZN(new_n984));
  NOR2_X1   g798(.A1(new_n707), .A2(new_n984), .ZN(new_n985));
  XNOR2_X1  g799(.A(new_n985), .B(KEYINPUT62), .ZN(new_n986));
  NAND3_X1  g800(.A1(new_n983), .A2(new_n794), .A3(new_n986), .ZN(new_n987));
  NAND2_X1  g801(.A1(new_n987), .A2(new_n226), .ZN(new_n988));
  NAND2_X1  g802(.A1(new_n600), .A2(new_n601), .ZN(new_n989));
  XNOR2_X1  g803(.A(new_n989), .B(new_n450), .ZN(new_n990));
  NAND2_X1  g804(.A1(new_n988), .A2(new_n990), .ZN(new_n991));
  INV_X1    g805(.A(KEYINPUT126), .ZN(new_n992));
  NOR2_X1   g806(.A1(new_n226), .A2(G900), .ZN(new_n993));
  AND3_X1   g807(.A1(new_n744), .A2(new_n620), .A3(new_n325), .ZN(new_n994));
  OAI211_X1 g808(.A(new_n684), .B(new_n787), .C1(new_n779), .C2(new_n994), .ZN(new_n995));
  AND2_X1   g809(.A1(new_n821), .A2(new_n771), .ZN(new_n996));
  NAND4_X1  g810(.A1(new_n794), .A2(new_n995), .A3(new_n769), .A4(new_n996), .ZN(new_n997));
  AOI21_X1  g811(.A(new_n993), .B1(new_n997), .B2(new_n226), .ZN(new_n998));
  INV_X1    g812(.A(KEYINPUT125), .ZN(new_n999));
  NAND2_X1  g813(.A1(new_n998), .A2(new_n999), .ZN(new_n1000));
  INV_X1    g814(.A(new_n1000), .ZN(new_n1001));
  INV_X1    g815(.A(new_n990), .ZN(new_n1002));
  OAI21_X1  g816(.A(new_n1002), .B1(new_n998), .B2(new_n999), .ZN(new_n1003));
  OAI211_X1 g817(.A(new_n991), .B(new_n992), .C1(new_n1001), .C2(new_n1003), .ZN(new_n1004));
  INV_X1    g818(.A(new_n1004), .ZN(new_n1005));
  AND2_X1   g819(.A1(new_n997), .A2(new_n226), .ZN(new_n1006));
  OAI21_X1  g820(.A(KEYINPUT125), .B1(new_n1006), .B2(new_n993), .ZN(new_n1007));
  NAND3_X1  g821(.A1(new_n1007), .A2(new_n1002), .A3(new_n1000), .ZN(new_n1008));
  AOI21_X1  g822(.A(new_n992), .B1(new_n1008), .B2(new_n991), .ZN(new_n1009));
  OAI21_X1  g823(.A(new_n968), .B1(new_n1005), .B2(new_n1009), .ZN(new_n1010));
  NAND2_X1  g824(.A1(new_n1008), .A2(new_n991), .ZN(new_n1011));
  NAND2_X1  g825(.A1(new_n1011), .A2(KEYINPUT126), .ZN(new_n1012));
  NAND3_X1  g826(.A1(new_n1012), .A2(new_n967), .A3(new_n1004), .ZN(new_n1013));
  NAND2_X1  g827(.A1(new_n1010), .A2(new_n1013), .ZN(G72));
  NAND2_X1  g828(.A1(G472), .A2(G902), .ZN(new_n1015));
  XOR2_X1   g829(.A(new_n1015), .B(KEYINPUT63), .Z(new_n1016));
  OAI21_X1  g830(.A(new_n1016), .B1(new_n987), .B2(new_n961), .ZN(new_n1017));
  NAND2_X1  g831(.A1(new_n1017), .A2(new_n697), .ZN(new_n1018));
  OAI21_X1  g832(.A(new_n1016), .B1(new_n997), .B2(new_n961), .ZN(new_n1019));
  AND3_X1   g833(.A1(new_n602), .A2(new_n579), .A3(new_n597), .ZN(new_n1020));
  AOI21_X1  g834(.A(new_n917), .B1(new_n1019), .B2(new_n1020), .ZN(new_n1021));
  NAND2_X1  g835(.A1(new_n1018), .A2(new_n1021), .ZN(new_n1022));
  INV_X1    g836(.A(new_n1016), .ZN(new_n1023));
  NOR3_X1   g837(.A1(new_n1020), .A2(new_n697), .A3(new_n1023), .ZN(new_n1024));
  AOI21_X1  g838(.A(new_n1022), .B1(new_n855), .B2(new_n1024), .ZN(G57));
endmodule


