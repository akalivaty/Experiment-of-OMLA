//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 1 1 0 0 1 1 0 0 1 1 0 1 1 1 1 1 1 1 0 0 1 0 0 0 0 0 1 1 0 0 1 1 1 0 0 1 0 1 0 1 0 1 1 1 0 1 0 1 0 0 1 0 0 1 0 1 0 1 1 0 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:33:53 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n456, new_n457,
    new_n458, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n535, new_n536, new_n537, new_n538, new_n539, new_n540,
    new_n541, new_n542, new_n545, new_n546, new_n547, new_n548, new_n549,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n559,
    new_n560, new_n562, new_n563, new_n564, new_n565, new_n566, new_n567,
    new_n568, new_n569, new_n570, new_n571, new_n572, new_n573, new_n574,
    new_n575, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n586, new_n587, new_n588, new_n589, new_n590, new_n591,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n614, new_n617, new_n619,
    new_n620, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1182, new_n1183, new_n1184,
    new_n1185, new_n1186, new_n1187;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  XOR2_X1   g002(.A(KEYINPUT64), .B(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  XNOR2_X1  g005(.A(KEYINPUT65), .B(G2066), .ZN(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  XOR2_X1   g008(.A(KEYINPUT66), .B(G44), .Z(G218));
  XOR2_X1   g009(.A(KEYINPUT67), .B(G132), .Z(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G218), .A2(G219), .A3(G220), .A4(G221), .ZN(new_n450));
  XOR2_X1   g025(.A(new_n450), .B(KEYINPUT2), .Z(new_n451));
  NOR4_X1   g026(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n452));
  INV_X1    g027(.A(new_n452), .ZN(new_n453));
  NOR2_X1   g028(.A1(new_n451), .A2(new_n453), .ZN(G325));
  INV_X1    g029(.A(G325), .ZN(G261));
  NAND2_X1  g030(.A1(new_n451), .A2(G2106), .ZN(new_n456));
  NAND2_X1  g031(.A1(new_n453), .A2(G567), .ZN(new_n457));
  NAND2_X1  g032(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  INV_X1    g033(.A(new_n458), .ZN(G319));
  INV_X1    g034(.A(G2105), .ZN(new_n460));
  AND2_X1   g035(.A1(new_n460), .A2(G2104), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n461), .A2(G101), .ZN(new_n462));
  OR2_X1    g037(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n463));
  NAND2_X1  g038(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n465), .A2(new_n460), .ZN(new_n466));
  INV_X1    g041(.A(G137), .ZN(new_n467));
  OAI21_X1  g042(.A(new_n462), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n465), .A2(G125), .ZN(new_n469));
  NAND2_X1  g044(.A1(G113), .A2(G2104), .ZN(new_n470));
  AOI21_X1  g045(.A(new_n460), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  NOR2_X1   g046(.A1(new_n468), .A2(new_n471), .ZN(G160));
  AND2_X1   g047(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n473));
  NOR2_X1   g048(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n474));
  NOR2_X1   g049(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  NOR2_X1   g050(.A1(new_n475), .A2(G2105), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n476), .A2(G136), .ZN(new_n477));
  NOR2_X1   g052(.A1(new_n475), .A2(new_n460), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n478), .A2(G124), .ZN(new_n479));
  OR2_X1    g054(.A1(G100), .A2(G2105), .ZN(new_n480));
  OAI211_X1 g055(.A(new_n480), .B(G2104), .C1(G112), .C2(new_n460), .ZN(new_n481));
  NAND3_X1  g056(.A1(new_n477), .A2(new_n479), .A3(new_n481), .ZN(new_n482));
  INV_X1    g057(.A(new_n482), .ZN(G162));
  NAND2_X1  g058(.A1(G126), .A2(G2105), .ZN(new_n484));
  AOI21_X1  g059(.A(new_n484), .B1(new_n463), .B2(new_n464), .ZN(new_n485));
  NOR2_X1   g060(.A1(new_n460), .A2(G114), .ZN(new_n486));
  OAI21_X1  g061(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n487));
  NOR2_X1   g062(.A1(new_n486), .A2(new_n487), .ZN(new_n488));
  OAI21_X1  g063(.A(KEYINPUT68), .B1(new_n485), .B2(new_n488), .ZN(new_n489));
  OAI211_X1 g064(.A(G126), .B(G2105), .C1(new_n473), .C2(new_n474), .ZN(new_n490));
  INV_X1    g065(.A(KEYINPUT68), .ZN(new_n491));
  OR2_X1    g066(.A1(G102), .A2(G2105), .ZN(new_n492));
  INV_X1    g067(.A(G114), .ZN(new_n493));
  NAND2_X1  g068(.A1(new_n493), .A2(G2105), .ZN(new_n494));
  NAND3_X1  g069(.A1(new_n492), .A2(new_n494), .A3(G2104), .ZN(new_n495));
  NAND3_X1  g070(.A1(new_n490), .A2(new_n491), .A3(new_n495), .ZN(new_n496));
  NAND2_X1  g071(.A1(new_n489), .A2(new_n496), .ZN(new_n497));
  OAI211_X1 g072(.A(G138), .B(new_n460), .C1(new_n473), .C2(new_n474), .ZN(new_n498));
  NAND2_X1  g073(.A1(new_n498), .A2(KEYINPUT4), .ZN(new_n499));
  INV_X1    g074(.A(KEYINPUT4), .ZN(new_n500));
  NAND4_X1  g075(.A1(new_n465), .A2(new_n500), .A3(G138), .A4(new_n460), .ZN(new_n501));
  NAND2_X1  g076(.A1(new_n499), .A2(new_n501), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n497), .A2(new_n502), .ZN(new_n503));
  NAND2_X1  g078(.A1(new_n503), .A2(KEYINPUT69), .ZN(new_n504));
  INV_X1    g079(.A(KEYINPUT69), .ZN(new_n505));
  NAND3_X1  g080(.A1(new_n497), .A2(new_n505), .A3(new_n502), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n504), .A2(new_n506), .ZN(G164));
  INV_X1    g082(.A(G543), .ZN(new_n508));
  INV_X1    g083(.A(KEYINPUT5), .ZN(new_n509));
  OAI21_X1  g084(.A(new_n508), .B1(new_n509), .B2(KEYINPUT72), .ZN(new_n510));
  INV_X1    g085(.A(KEYINPUT72), .ZN(new_n511));
  NAND3_X1  g086(.A1(new_n511), .A2(KEYINPUT5), .A3(G543), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n510), .A2(new_n512), .ZN(new_n513));
  AOI22_X1  g088(.A1(new_n513), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n514));
  XNOR2_X1  g089(.A(KEYINPUT70), .B(G651), .ZN(new_n515));
  INV_X1    g090(.A(new_n515), .ZN(new_n516));
  OR2_X1    g091(.A1(new_n514), .A2(new_n516), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n515), .A2(KEYINPUT6), .ZN(new_n518));
  NOR2_X1   g093(.A1(KEYINPUT6), .A2(G651), .ZN(new_n519));
  INV_X1    g094(.A(new_n519), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n518), .A2(new_n520), .ZN(new_n521));
  NAND3_X1  g096(.A1(new_n521), .A2(KEYINPUT73), .A3(new_n513), .ZN(new_n522));
  INV_X1    g097(.A(KEYINPUT73), .ZN(new_n523));
  AOI21_X1  g098(.A(new_n519), .B1(new_n515), .B2(KEYINPUT6), .ZN(new_n524));
  INV_X1    g099(.A(new_n513), .ZN(new_n525));
  OAI21_X1  g100(.A(new_n523), .B1(new_n524), .B2(new_n525), .ZN(new_n526));
  NAND2_X1  g101(.A1(new_n522), .A2(new_n526), .ZN(new_n527));
  INV_X1    g102(.A(G88), .ZN(new_n528));
  AND2_X1   g103(.A1(G50), .A2(G543), .ZN(new_n529));
  NAND2_X1  g104(.A1(new_n521), .A2(new_n529), .ZN(new_n530));
  AND2_X1   g105(.A1(new_n530), .A2(KEYINPUT71), .ZN(new_n531));
  NOR2_X1   g106(.A1(new_n530), .A2(KEYINPUT71), .ZN(new_n532));
  OAI221_X1 g107(.A(new_n517), .B1(new_n527), .B2(new_n528), .C1(new_n531), .C2(new_n532), .ZN(G303));
  INV_X1    g108(.A(G303), .ZN(G166));
  AND3_X1   g109(.A1(new_n513), .A2(G63), .A3(G651), .ZN(new_n535));
  XOR2_X1   g110(.A(KEYINPUT74), .B(KEYINPUT7), .Z(new_n536));
  NAND3_X1  g111(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n537));
  XNOR2_X1  g112(.A(new_n536), .B(new_n537), .ZN(new_n538));
  NOR2_X1   g113(.A1(new_n524), .A2(new_n508), .ZN(new_n539));
  AOI211_X1 g114(.A(new_n535), .B(new_n538), .C1(G51), .C2(new_n539), .ZN(new_n540));
  INV_X1    g115(.A(new_n527), .ZN(new_n541));
  NAND2_X1  g116(.A1(new_n541), .A2(G89), .ZN(new_n542));
  NAND2_X1  g117(.A1(new_n540), .A2(new_n542), .ZN(G286));
  INV_X1    g118(.A(G286), .ZN(G168));
  NAND2_X1  g119(.A1(new_n541), .A2(G90), .ZN(new_n545));
  NAND2_X1  g120(.A1(G77), .A2(G543), .ZN(new_n546));
  INV_X1    g121(.A(G64), .ZN(new_n547));
  OAI21_X1  g122(.A(new_n546), .B1(new_n525), .B2(new_n547), .ZN(new_n548));
  AOI22_X1  g123(.A1(G52), .A2(new_n539), .B1(new_n548), .B2(new_n515), .ZN(new_n549));
  AND2_X1   g124(.A1(new_n545), .A2(new_n549), .ZN(G171));
  AOI22_X1  g125(.A1(new_n513), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n551));
  OR2_X1    g126(.A1(new_n551), .A2(new_n516), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n539), .A2(G43), .ZN(new_n553));
  INV_X1    g128(.A(G81), .ZN(new_n554));
  OAI211_X1 g129(.A(new_n552), .B(new_n553), .C1(new_n527), .C2(new_n554), .ZN(new_n555));
  INV_X1    g130(.A(new_n555), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n556), .A2(G860), .ZN(G153));
  NAND4_X1  g132(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g133(.A1(G1), .A2(G3), .ZN(new_n559));
  XNOR2_X1  g134(.A(new_n559), .B(KEYINPUT8), .ZN(new_n560));
  NAND4_X1  g135(.A1(G319), .A2(G483), .A3(G661), .A4(new_n560), .ZN(G188));
  INV_X1    g136(.A(G91), .ZN(new_n562));
  OAI21_X1  g137(.A(KEYINPUT75), .B1(new_n527), .B2(new_n562), .ZN(new_n563));
  INV_X1    g138(.A(KEYINPUT75), .ZN(new_n564));
  NAND4_X1  g139(.A1(new_n522), .A2(new_n526), .A3(new_n564), .A4(G91), .ZN(new_n565));
  NAND2_X1  g140(.A1(new_n563), .A2(new_n565), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n539), .A2(G53), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n567), .A2(KEYINPUT9), .ZN(new_n568));
  INV_X1    g143(.A(KEYINPUT9), .ZN(new_n569));
  NAND3_X1  g144(.A1(new_n539), .A2(new_n569), .A3(G53), .ZN(new_n570));
  NAND2_X1  g145(.A1(G78), .A2(G543), .ZN(new_n571));
  XNOR2_X1  g146(.A(new_n513), .B(KEYINPUT76), .ZN(new_n572));
  INV_X1    g147(.A(G65), .ZN(new_n573));
  OAI21_X1  g148(.A(new_n571), .B1(new_n572), .B2(new_n573), .ZN(new_n574));
  AOI22_X1  g149(.A1(new_n568), .A2(new_n570), .B1(new_n574), .B2(G651), .ZN(new_n575));
  NAND2_X1  g150(.A1(new_n566), .A2(new_n575), .ZN(G299));
  INV_X1    g151(.A(G171), .ZN(G301));
  INV_X1    g152(.A(G87), .ZN(new_n578));
  OAI21_X1  g153(.A(KEYINPUT77), .B1(new_n527), .B2(new_n578), .ZN(new_n579));
  INV_X1    g154(.A(KEYINPUT77), .ZN(new_n580));
  NAND4_X1  g155(.A1(new_n522), .A2(new_n526), .A3(new_n580), .A4(G87), .ZN(new_n581));
  NAND2_X1  g156(.A1(new_n579), .A2(new_n581), .ZN(new_n582));
  OR2_X1    g157(.A1(new_n513), .A2(G74), .ZN(new_n583));
  AOI22_X1  g158(.A1(new_n539), .A2(G49), .B1(new_n583), .B2(G651), .ZN(new_n584));
  NAND2_X1  g159(.A1(new_n582), .A2(new_n584), .ZN(G288));
  NAND2_X1  g160(.A1(new_n513), .A2(G61), .ZN(new_n586));
  NAND2_X1  g161(.A1(G73), .A2(G543), .ZN(new_n587));
  XNOR2_X1  g162(.A(new_n587), .B(KEYINPUT78), .ZN(new_n588));
  AOI21_X1  g163(.A(new_n516), .B1(new_n586), .B2(new_n588), .ZN(new_n589));
  AOI21_X1  g164(.A(new_n589), .B1(G48), .B2(new_n539), .ZN(new_n590));
  NAND3_X1  g165(.A1(new_n522), .A2(G86), .A3(new_n526), .ZN(new_n591));
  NAND2_X1  g166(.A1(new_n590), .A2(new_n591), .ZN(G305));
  AND2_X1   g167(.A1(new_n513), .A2(G60), .ZN(new_n593));
  AND2_X1   g168(.A1(G72), .A2(G543), .ZN(new_n594));
  OAI21_X1  g169(.A(new_n515), .B1(new_n593), .B2(new_n594), .ZN(new_n595));
  XNOR2_X1  g170(.A(new_n595), .B(KEYINPUT79), .ZN(new_n596));
  NAND2_X1  g171(.A1(new_n541), .A2(G85), .ZN(new_n597));
  NAND2_X1  g172(.A1(new_n539), .A2(G47), .ZN(new_n598));
  NAND3_X1  g173(.A1(new_n596), .A2(new_n597), .A3(new_n598), .ZN(G290));
  INV_X1    g174(.A(G868), .ZN(new_n600));
  NOR2_X1   g175(.A1(G301), .A2(new_n600), .ZN(new_n601));
  NAND3_X1  g176(.A1(new_n522), .A2(G92), .A3(new_n526), .ZN(new_n602));
  XOR2_X1   g177(.A(KEYINPUT80), .B(KEYINPUT10), .Z(new_n603));
  XNOR2_X1  g178(.A(new_n602), .B(new_n603), .ZN(new_n604));
  NAND2_X1  g179(.A1(G79), .A2(G543), .ZN(new_n605));
  INV_X1    g180(.A(G66), .ZN(new_n606));
  OAI21_X1  g181(.A(new_n605), .B1(new_n572), .B2(new_n606), .ZN(new_n607));
  AOI22_X1  g182(.A1(new_n607), .A2(G651), .B1(G54), .B2(new_n539), .ZN(new_n608));
  NAND2_X1  g183(.A1(new_n604), .A2(new_n608), .ZN(new_n609));
  INV_X1    g184(.A(KEYINPUT81), .ZN(new_n610));
  XNOR2_X1  g185(.A(new_n609), .B(new_n610), .ZN(new_n611));
  AOI21_X1  g186(.A(new_n601), .B1(new_n611), .B2(new_n600), .ZN(G284));
  AOI21_X1  g187(.A(new_n601), .B1(new_n611), .B2(new_n600), .ZN(G321));
  NAND2_X1  g188(.A1(G299), .A2(new_n600), .ZN(new_n614));
  OAI21_X1  g189(.A(new_n614), .B1(new_n600), .B2(G168), .ZN(G297));
  XNOR2_X1  g190(.A(G297), .B(KEYINPUT82), .ZN(G280));
  INV_X1    g191(.A(G559), .ZN(new_n617));
  OAI21_X1  g192(.A(new_n611), .B1(new_n617), .B2(G860), .ZN(G148));
  NAND2_X1  g193(.A1(new_n555), .A2(new_n600), .ZN(new_n619));
  AND2_X1   g194(.A1(new_n611), .A2(new_n617), .ZN(new_n620));
  OAI21_X1  g195(.A(new_n619), .B1(new_n620), .B2(new_n600), .ZN(G323));
  XNOR2_X1  g196(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g197(.A1(new_n465), .A2(new_n461), .ZN(new_n623));
  XNOR2_X1  g198(.A(new_n623), .B(KEYINPUT12), .ZN(new_n624));
  XNOR2_X1  g199(.A(new_n624), .B(KEYINPUT13), .ZN(new_n625));
  INV_X1    g200(.A(G2100), .ZN(new_n626));
  OR2_X1    g201(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  NAND2_X1  g202(.A1(new_n625), .A2(new_n626), .ZN(new_n628));
  NAND2_X1  g203(.A1(new_n476), .A2(G135), .ZN(new_n629));
  NAND2_X1  g204(.A1(new_n478), .A2(G123), .ZN(new_n630));
  NOR2_X1   g205(.A1(new_n460), .A2(G111), .ZN(new_n631));
  OAI21_X1  g206(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n632));
  OAI211_X1 g207(.A(new_n629), .B(new_n630), .C1(new_n631), .C2(new_n632), .ZN(new_n633));
  INV_X1    g208(.A(G2096), .ZN(new_n634));
  XNOR2_X1  g209(.A(new_n633), .B(new_n634), .ZN(new_n635));
  NAND3_X1  g210(.A1(new_n627), .A2(new_n628), .A3(new_n635), .ZN(new_n636));
  XNOR2_X1  g211(.A(new_n636), .B(KEYINPUT83), .ZN(G156));
  XNOR2_X1  g212(.A(G2427), .B(G2438), .ZN(new_n638));
  XNOR2_X1  g213(.A(new_n638), .B(G2430), .ZN(new_n639));
  XNOR2_X1  g214(.A(KEYINPUT15), .B(G2435), .ZN(new_n640));
  OR2_X1    g215(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  NAND2_X1  g216(.A1(new_n639), .A2(new_n640), .ZN(new_n642));
  NAND3_X1  g217(.A1(new_n641), .A2(KEYINPUT14), .A3(new_n642), .ZN(new_n643));
  XNOR2_X1  g218(.A(new_n643), .B(KEYINPUT84), .ZN(new_n644));
  INV_X1    g219(.A(G1341), .ZN(new_n645));
  XNOR2_X1  g220(.A(new_n644), .B(new_n645), .ZN(new_n646));
  XNOR2_X1  g221(.A(new_n646), .B(G1348), .ZN(new_n647));
  XOR2_X1   g222(.A(G2451), .B(G2454), .Z(new_n648));
  XNOR2_X1  g223(.A(new_n648), .B(KEYINPUT16), .ZN(new_n649));
  XOR2_X1   g224(.A(G2443), .B(G2446), .Z(new_n650));
  XNOR2_X1  g225(.A(new_n649), .B(new_n650), .ZN(new_n651));
  NAND2_X1  g226(.A1(new_n647), .A2(new_n651), .ZN(new_n652));
  NAND2_X1  g227(.A1(new_n652), .A2(G14), .ZN(new_n653));
  NOR2_X1   g228(.A1(new_n647), .A2(new_n651), .ZN(new_n654));
  OR2_X1    g229(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  INV_X1    g230(.A(new_n655), .ZN(G401));
  INV_X1    g231(.A(KEYINPUT18), .ZN(new_n657));
  XOR2_X1   g232(.A(G2084), .B(G2090), .Z(new_n658));
  XNOR2_X1  g233(.A(G2067), .B(G2678), .ZN(new_n659));
  NAND2_X1  g234(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  NAND2_X1  g235(.A1(new_n660), .A2(KEYINPUT17), .ZN(new_n661));
  NOR2_X1   g236(.A1(new_n658), .A2(new_n659), .ZN(new_n662));
  OAI21_X1  g237(.A(new_n657), .B1(new_n661), .B2(new_n662), .ZN(new_n663));
  XNOR2_X1  g238(.A(new_n663), .B(new_n626), .ZN(new_n664));
  XOR2_X1   g239(.A(G2072), .B(G2078), .Z(new_n665));
  AOI21_X1  g240(.A(new_n665), .B1(new_n660), .B2(KEYINPUT18), .ZN(new_n666));
  XNOR2_X1  g241(.A(new_n666), .B(new_n634), .ZN(new_n667));
  XNOR2_X1  g242(.A(new_n664), .B(new_n667), .ZN(G227));
  XOR2_X1   g243(.A(G1971), .B(G1976), .Z(new_n669));
  XNOR2_X1  g244(.A(KEYINPUT85), .B(KEYINPUT19), .ZN(new_n670));
  XNOR2_X1  g245(.A(new_n669), .B(new_n670), .ZN(new_n671));
  XNOR2_X1  g246(.A(G1956), .B(G2474), .ZN(new_n672));
  XNOR2_X1  g247(.A(G1961), .B(G1966), .ZN(new_n673));
  NOR2_X1   g248(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  INV_X1    g249(.A(new_n674), .ZN(new_n675));
  NOR2_X1   g250(.A1(new_n671), .A2(new_n675), .ZN(new_n676));
  XOR2_X1   g251(.A(new_n676), .B(KEYINPUT20), .Z(new_n677));
  NAND2_X1  g252(.A1(new_n672), .A2(new_n673), .ZN(new_n678));
  NAND3_X1  g253(.A1(new_n671), .A2(new_n675), .A3(new_n678), .ZN(new_n679));
  OAI211_X1 g254(.A(new_n677), .B(new_n679), .C1(new_n671), .C2(new_n678), .ZN(new_n680));
  XNOR2_X1  g255(.A(G1991), .B(G1996), .ZN(new_n681));
  XNOR2_X1  g256(.A(new_n680), .B(new_n681), .ZN(new_n682));
  XOR2_X1   g257(.A(G1981), .B(G1986), .Z(new_n683));
  XNOR2_X1  g258(.A(new_n683), .B(KEYINPUT86), .ZN(new_n684));
  XOR2_X1   g259(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n685));
  XNOR2_X1  g260(.A(new_n684), .B(new_n685), .ZN(new_n686));
  XNOR2_X1  g261(.A(new_n682), .B(new_n686), .ZN(G229));
  INV_X1    g262(.A(G16), .ZN(new_n688));
  NAND2_X1  g263(.A1(new_n688), .A2(G23), .ZN(new_n689));
  AND2_X1   g264(.A1(new_n582), .A2(new_n584), .ZN(new_n690));
  OAI21_X1  g265(.A(new_n689), .B1(new_n690), .B2(new_n688), .ZN(new_n691));
  XNOR2_X1  g266(.A(KEYINPUT33), .B(G1976), .ZN(new_n692));
  INV_X1    g267(.A(new_n692), .ZN(new_n693));
  XNOR2_X1  g268(.A(new_n691), .B(new_n693), .ZN(new_n694));
  INV_X1    g269(.A(KEYINPUT87), .ZN(new_n695));
  NAND2_X1  g270(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  XNOR2_X1  g271(.A(new_n691), .B(new_n692), .ZN(new_n697));
  NAND2_X1  g272(.A1(new_n697), .A2(KEYINPUT87), .ZN(new_n698));
  NAND2_X1  g273(.A1(new_n688), .A2(G22), .ZN(new_n699));
  OAI21_X1  g274(.A(new_n699), .B1(G166), .B2(new_n688), .ZN(new_n700));
  XNOR2_X1  g275(.A(new_n700), .B(G1971), .ZN(new_n701));
  NOR2_X1   g276(.A1(G6), .A2(G16), .ZN(new_n702));
  INV_X1    g277(.A(G305), .ZN(new_n703));
  AOI21_X1  g278(.A(new_n702), .B1(new_n703), .B2(G16), .ZN(new_n704));
  XNOR2_X1  g279(.A(KEYINPUT32), .B(G1981), .ZN(new_n705));
  XNOR2_X1  g280(.A(new_n704), .B(new_n705), .ZN(new_n706));
  NOR2_X1   g281(.A1(new_n701), .A2(new_n706), .ZN(new_n707));
  NAND3_X1  g282(.A1(new_n696), .A2(new_n698), .A3(new_n707), .ZN(new_n708));
  NAND2_X1  g283(.A1(new_n708), .A2(KEYINPUT34), .ZN(new_n709));
  INV_X1    g284(.A(KEYINPUT34), .ZN(new_n710));
  NAND4_X1  g285(.A1(new_n696), .A2(new_n698), .A3(new_n710), .A4(new_n707), .ZN(new_n711));
  INV_X1    g286(.A(G29), .ZN(new_n712));
  NAND2_X1  g287(.A1(new_n712), .A2(G25), .ZN(new_n713));
  NAND2_X1  g288(.A1(new_n476), .A2(G131), .ZN(new_n714));
  NAND2_X1  g289(.A1(new_n478), .A2(G119), .ZN(new_n715));
  OR2_X1    g290(.A1(G95), .A2(G2105), .ZN(new_n716));
  OAI211_X1 g291(.A(new_n716), .B(G2104), .C1(G107), .C2(new_n460), .ZN(new_n717));
  NAND3_X1  g292(.A1(new_n714), .A2(new_n715), .A3(new_n717), .ZN(new_n718));
  INV_X1    g293(.A(new_n718), .ZN(new_n719));
  OAI21_X1  g294(.A(new_n713), .B1(new_n719), .B2(new_n712), .ZN(new_n720));
  XOR2_X1   g295(.A(KEYINPUT35), .B(G1991), .Z(new_n721));
  XNOR2_X1  g296(.A(new_n720), .B(new_n721), .ZN(new_n722));
  AND2_X1   g297(.A1(new_n688), .A2(G24), .ZN(new_n723));
  AOI21_X1  g298(.A(new_n723), .B1(G290), .B2(G16), .ZN(new_n724));
  INV_X1    g299(.A(G1986), .ZN(new_n725));
  OAI21_X1  g300(.A(new_n722), .B1(new_n724), .B2(new_n725), .ZN(new_n726));
  AOI21_X1  g301(.A(new_n726), .B1(new_n725), .B2(new_n724), .ZN(new_n727));
  NAND3_X1  g302(.A1(new_n709), .A2(new_n711), .A3(new_n727), .ZN(new_n728));
  NAND2_X1  g303(.A1(new_n728), .A2(KEYINPUT36), .ZN(new_n729));
  INV_X1    g304(.A(KEYINPUT36), .ZN(new_n730));
  NAND4_X1  g305(.A1(new_n709), .A2(new_n730), .A3(new_n711), .A4(new_n727), .ZN(new_n731));
  NAND2_X1  g306(.A1(new_n729), .A2(new_n731), .ZN(new_n732));
  INV_X1    g307(.A(KEYINPUT25), .ZN(new_n733));
  NAND2_X1  g308(.A1(G103), .A2(G2104), .ZN(new_n734));
  OAI21_X1  g309(.A(new_n733), .B1(new_n734), .B2(G2105), .ZN(new_n735));
  NAND4_X1  g310(.A1(new_n460), .A2(KEYINPUT25), .A3(G103), .A4(G2104), .ZN(new_n736));
  AOI22_X1  g311(.A1(new_n476), .A2(G139), .B1(new_n735), .B2(new_n736), .ZN(new_n737));
  AOI22_X1  g312(.A1(new_n465), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n738));
  OAI21_X1  g313(.A(new_n737), .B1(new_n460), .B2(new_n738), .ZN(new_n739));
  MUX2_X1   g314(.A(G33), .B(new_n739), .S(G29), .Z(new_n740));
  XNOR2_X1  g315(.A(new_n740), .B(KEYINPUT89), .ZN(new_n741));
  INV_X1    g316(.A(G2072), .ZN(new_n742));
  NAND2_X1  g317(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  INV_X1    g318(.A(KEYINPUT90), .ZN(new_n744));
  XNOR2_X1  g319(.A(new_n743), .B(new_n744), .ZN(new_n745));
  NAND2_X1  g320(.A1(new_n688), .A2(G5), .ZN(new_n746));
  OAI21_X1  g321(.A(new_n746), .B1(G171), .B2(new_n688), .ZN(new_n747));
  XNOR2_X1  g322(.A(KEYINPUT94), .B(G1961), .ZN(new_n748));
  INV_X1    g323(.A(new_n748), .ZN(new_n749));
  NAND2_X1  g324(.A1(new_n747), .A2(new_n749), .ZN(new_n750));
  NAND2_X1  g325(.A1(new_n712), .A2(G27), .ZN(new_n751));
  OAI21_X1  g326(.A(new_n751), .B1(G164), .B2(new_n712), .ZN(new_n752));
  XNOR2_X1  g327(.A(KEYINPUT95), .B(G2078), .ZN(new_n753));
  INV_X1    g328(.A(new_n753), .ZN(new_n754));
  NAND2_X1  g329(.A1(new_n752), .A2(new_n754), .ZN(new_n755));
  OR2_X1    g330(.A1(new_n752), .A2(new_n754), .ZN(new_n756));
  NAND3_X1  g331(.A1(new_n750), .A2(new_n755), .A3(new_n756), .ZN(new_n757));
  INV_X1    g332(.A(new_n757), .ZN(new_n758));
  NOR2_X1   g333(.A1(new_n747), .A2(new_n749), .ZN(new_n759));
  INV_X1    g334(.A(G34), .ZN(new_n760));
  AND2_X1   g335(.A1(new_n760), .A2(KEYINPUT24), .ZN(new_n761));
  NOR2_X1   g336(.A1(new_n760), .A2(KEYINPUT24), .ZN(new_n762));
  OAI21_X1  g337(.A(new_n712), .B1(new_n761), .B2(new_n762), .ZN(new_n763));
  OAI21_X1  g338(.A(new_n763), .B1(G160), .B2(new_n712), .ZN(new_n764));
  XNOR2_X1  g339(.A(new_n764), .B(G2084), .ZN(new_n765));
  XNOR2_X1  g340(.A(KEYINPUT30), .B(G28), .ZN(new_n766));
  OR2_X1    g341(.A1(KEYINPUT31), .A2(G11), .ZN(new_n767));
  NAND2_X1  g342(.A1(KEYINPUT31), .A2(G11), .ZN(new_n768));
  AOI22_X1  g343(.A1(new_n766), .A2(new_n712), .B1(new_n767), .B2(new_n768), .ZN(new_n769));
  OAI21_X1  g344(.A(new_n769), .B1(new_n633), .B2(new_n712), .ZN(new_n770));
  AND2_X1   g345(.A1(new_n712), .A2(G32), .ZN(new_n771));
  AOI22_X1  g346(.A1(new_n476), .A2(G141), .B1(G105), .B2(new_n461), .ZN(new_n772));
  NAND2_X1  g347(.A1(new_n478), .A2(G129), .ZN(new_n773));
  NAND3_X1  g348(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n774));
  XOR2_X1   g349(.A(new_n774), .B(KEYINPUT26), .Z(new_n775));
  NAND3_X1  g350(.A1(new_n772), .A2(new_n773), .A3(new_n775), .ZN(new_n776));
  AOI21_X1  g351(.A(new_n771), .B1(new_n776), .B2(G29), .ZN(new_n777));
  XNOR2_X1  g352(.A(KEYINPUT27), .B(G1996), .ZN(new_n778));
  AOI21_X1  g353(.A(new_n770), .B1(new_n777), .B2(new_n778), .ZN(new_n779));
  OAI21_X1  g354(.A(new_n779), .B1(new_n777), .B2(new_n778), .ZN(new_n780));
  NOR3_X1   g355(.A1(new_n759), .A2(new_n765), .A3(new_n780), .ZN(new_n781));
  AND3_X1   g356(.A1(new_n745), .A2(new_n758), .A3(new_n781), .ZN(new_n782));
  INV_X1    g357(.A(KEYINPUT91), .ZN(new_n783));
  OR3_X1    g358(.A1(new_n741), .A2(new_n783), .A3(new_n742), .ZN(new_n784));
  OAI21_X1  g359(.A(new_n783), .B1(new_n741), .B2(new_n742), .ZN(new_n785));
  NAND2_X1  g360(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  AND2_X1   g361(.A1(new_n688), .A2(G21), .ZN(new_n787));
  AOI21_X1  g362(.A(new_n787), .B1(G286), .B2(G16), .ZN(new_n788));
  INV_X1    g363(.A(G1966), .ZN(new_n789));
  OR2_X1    g364(.A1(new_n788), .A2(new_n789), .ZN(new_n790));
  INV_X1    g365(.A(KEYINPUT92), .ZN(new_n791));
  OR2_X1    g366(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  NAND2_X1  g367(.A1(new_n790), .A2(new_n791), .ZN(new_n793));
  NAND3_X1  g368(.A1(new_n786), .A2(new_n792), .A3(new_n793), .ZN(new_n794));
  INV_X1    g369(.A(new_n794), .ZN(new_n795));
  INV_X1    g370(.A(KEYINPUT96), .ZN(new_n796));
  NAND2_X1  g371(.A1(new_n788), .A2(new_n789), .ZN(new_n797));
  XNOR2_X1  g372(.A(new_n797), .B(KEYINPUT93), .ZN(new_n798));
  NAND4_X1  g373(.A1(new_n782), .A2(new_n795), .A3(new_n796), .A4(new_n798), .ZN(new_n799));
  NAND4_X1  g374(.A1(new_n745), .A2(new_n798), .A3(new_n758), .A4(new_n781), .ZN(new_n800));
  OAI21_X1  g375(.A(KEYINPUT96), .B1(new_n800), .B2(new_n794), .ZN(new_n801));
  OR2_X1    g376(.A1(G16), .A2(G19), .ZN(new_n802));
  OAI21_X1  g377(.A(new_n802), .B1(new_n555), .B2(new_n688), .ZN(new_n803));
  OR2_X1    g378(.A1(new_n803), .A2(new_n645), .ZN(new_n804));
  NAND2_X1  g379(.A1(new_n712), .A2(G26), .ZN(new_n805));
  XOR2_X1   g380(.A(new_n805), .B(KEYINPUT28), .Z(new_n806));
  NAND2_X1  g381(.A1(new_n476), .A2(G140), .ZN(new_n807));
  INV_X1    g382(.A(KEYINPUT88), .ZN(new_n808));
  XNOR2_X1  g383(.A(new_n807), .B(new_n808), .ZN(new_n809));
  OAI21_X1  g384(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n810));
  INV_X1    g385(.A(G116), .ZN(new_n811));
  AOI21_X1  g386(.A(new_n810), .B1(new_n811), .B2(G2105), .ZN(new_n812));
  AOI21_X1  g387(.A(new_n812), .B1(new_n478), .B2(G128), .ZN(new_n813));
  NAND2_X1  g388(.A1(new_n809), .A2(new_n813), .ZN(new_n814));
  AOI21_X1  g389(.A(new_n806), .B1(new_n814), .B2(G29), .ZN(new_n815));
  XNOR2_X1  g390(.A(new_n815), .B(G2067), .ZN(new_n816));
  NAND2_X1  g391(.A1(new_n803), .A2(new_n645), .ZN(new_n817));
  NAND2_X1  g392(.A1(new_n712), .A2(G35), .ZN(new_n818));
  OAI21_X1  g393(.A(new_n818), .B1(G162), .B2(new_n712), .ZN(new_n819));
  XNOR2_X1  g394(.A(new_n819), .B(KEYINPUT29), .ZN(new_n820));
  NAND2_X1  g395(.A1(new_n820), .A2(G2090), .ZN(new_n821));
  AND4_X1   g396(.A1(new_n804), .A2(new_n816), .A3(new_n817), .A4(new_n821), .ZN(new_n822));
  NAND2_X1  g397(.A1(new_n688), .A2(G20), .ZN(new_n823));
  XOR2_X1   g398(.A(new_n823), .B(KEYINPUT23), .Z(new_n824));
  AOI21_X1  g399(.A(new_n824), .B1(G299), .B2(G16), .ZN(new_n825));
  XNOR2_X1  g400(.A(KEYINPUT98), .B(G1956), .ZN(new_n826));
  XNOR2_X1  g401(.A(new_n825), .B(new_n826), .ZN(new_n827));
  INV_X1    g402(.A(KEYINPUT97), .ZN(new_n828));
  INV_X1    g403(.A(new_n820), .ZN(new_n829));
  INV_X1    g404(.A(G2090), .ZN(new_n830));
  AOI21_X1  g405(.A(new_n828), .B1(new_n829), .B2(new_n830), .ZN(new_n831));
  NOR3_X1   g406(.A1(new_n820), .A2(KEYINPUT97), .A3(G2090), .ZN(new_n832));
  OAI211_X1 g407(.A(new_n822), .B(new_n827), .C1(new_n831), .C2(new_n832), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n688), .A2(G4), .ZN(new_n834));
  OAI21_X1  g409(.A(new_n834), .B1(new_n611), .B2(new_n688), .ZN(new_n835));
  AOI21_X1  g410(.A(new_n833), .B1(G1348), .B2(new_n835), .ZN(new_n836));
  OR2_X1    g411(.A1(new_n835), .A2(G1348), .ZN(new_n837));
  NAND4_X1  g412(.A1(new_n799), .A2(new_n801), .A3(new_n836), .A4(new_n837), .ZN(new_n838));
  INV_X1    g413(.A(new_n838), .ZN(new_n839));
  AOI21_X1  g414(.A(KEYINPUT99), .B1(new_n732), .B2(new_n839), .ZN(new_n840));
  INV_X1    g415(.A(KEYINPUT99), .ZN(new_n841));
  AOI211_X1 g416(.A(new_n841), .B(new_n838), .C1(new_n729), .C2(new_n731), .ZN(new_n842));
  NOR2_X1   g417(.A1(new_n840), .A2(new_n842), .ZN(G311));
  NAND2_X1  g418(.A1(new_n732), .A2(new_n839), .ZN(G150));
  AOI22_X1  g419(.A1(new_n513), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n845));
  OR2_X1    g420(.A1(new_n845), .A2(new_n516), .ZN(new_n846));
  XOR2_X1   g421(.A(KEYINPUT100), .B(G93), .Z(new_n847));
  NAND3_X1  g422(.A1(new_n522), .A2(new_n526), .A3(new_n847), .ZN(new_n848));
  NAND2_X1  g423(.A1(new_n539), .A2(G55), .ZN(new_n849));
  AND3_X1   g424(.A1(new_n848), .A2(KEYINPUT101), .A3(new_n849), .ZN(new_n850));
  AOI21_X1  g425(.A(KEYINPUT101), .B1(new_n848), .B2(new_n849), .ZN(new_n851));
  OAI21_X1  g426(.A(new_n846), .B1(new_n850), .B2(new_n851), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n852), .A2(G860), .ZN(new_n853));
  XNOR2_X1  g428(.A(new_n853), .B(KEYINPUT102), .ZN(new_n854));
  XNOR2_X1  g429(.A(new_n854), .B(KEYINPUT37), .ZN(new_n855));
  INV_X1    g430(.A(G860), .ZN(new_n856));
  NAND2_X1  g431(.A1(new_n611), .A2(G559), .ZN(new_n857));
  XNOR2_X1  g432(.A(new_n857), .B(KEYINPUT38), .ZN(new_n858));
  NAND2_X1  g433(.A1(new_n852), .A2(new_n555), .ZN(new_n859));
  OAI211_X1 g434(.A(new_n556), .B(new_n846), .C1(new_n850), .C2(new_n851), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  INV_X1    g436(.A(new_n861), .ZN(new_n862));
  XNOR2_X1  g437(.A(new_n858), .B(new_n862), .ZN(new_n863));
  OAI21_X1  g438(.A(new_n856), .B1(new_n863), .B2(KEYINPUT39), .ZN(new_n864));
  XNOR2_X1  g439(.A(new_n858), .B(new_n861), .ZN(new_n865));
  INV_X1    g440(.A(KEYINPUT39), .ZN(new_n866));
  NOR2_X1   g441(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  OAI21_X1  g442(.A(new_n855), .B1(new_n864), .B2(new_n867), .ZN(new_n868));
  NAND2_X1  g443(.A1(new_n868), .A2(KEYINPUT103), .ZN(new_n869));
  INV_X1    g444(.A(KEYINPUT103), .ZN(new_n870));
  OAI211_X1 g445(.A(new_n870), .B(new_n855), .C1(new_n864), .C2(new_n867), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n869), .A2(new_n871), .ZN(G145));
  INV_X1    g447(.A(KEYINPUT106), .ZN(new_n873));
  XNOR2_X1  g448(.A(new_n814), .B(new_n739), .ZN(new_n874));
  NOR2_X1   g449(.A1(new_n485), .A2(new_n488), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n502), .A2(new_n875), .ZN(new_n876));
  XOR2_X1   g451(.A(new_n874), .B(new_n876), .Z(new_n877));
  NAND2_X1  g452(.A1(new_n877), .A2(new_n776), .ZN(new_n878));
  XNOR2_X1  g453(.A(new_n874), .B(new_n876), .ZN(new_n879));
  INV_X1    g454(.A(new_n776), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n878), .A2(new_n881), .ZN(new_n882));
  XNOR2_X1  g457(.A(new_n718), .B(new_n624), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n476), .A2(G142), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n478), .A2(G130), .ZN(new_n885));
  OAI21_X1  g460(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n886));
  INV_X1    g461(.A(KEYINPUT104), .ZN(new_n887));
  INV_X1    g462(.A(G118), .ZN(new_n888));
  AOI22_X1  g463(.A1(new_n886), .A2(new_n887), .B1(new_n888), .B2(G2105), .ZN(new_n889));
  OAI21_X1  g464(.A(new_n889), .B1(new_n887), .B2(new_n886), .ZN(new_n890));
  NAND3_X1  g465(.A1(new_n884), .A2(new_n885), .A3(new_n890), .ZN(new_n891));
  XNOR2_X1  g466(.A(new_n883), .B(new_n891), .ZN(new_n892));
  XOR2_X1   g467(.A(new_n892), .B(KEYINPUT105), .Z(new_n893));
  NAND2_X1  g468(.A1(new_n882), .A2(new_n893), .ZN(new_n894));
  XOR2_X1   g469(.A(G160), .B(new_n633), .Z(new_n895));
  XNOR2_X1  g470(.A(new_n895), .B(new_n482), .ZN(new_n896));
  INV_X1    g471(.A(new_n896), .ZN(new_n897));
  NAND3_X1  g472(.A1(new_n878), .A2(new_n881), .A3(new_n892), .ZN(new_n898));
  NAND3_X1  g473(.A1(new_n894), .A2(new_n897), .A3(new_n898), .ZN(new_n899));
  INV_X1    g474(.A(G37), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  INV_X1    g476(.A(new_n893), .ZN(new_n902));
  NAND3_X1  g477(.A1(new_n878), .A2(new_n881), .A3(new_n902), .ZN(new_n903));
  AOI21_X1  g478(.A(new_n897), .B1(new_n894), .B2(new_n903), .ZN(new_n904));
  OAI21_X1  g479(.A(new_n873), .B1(new_n901), .B2(new_n904), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n894), .A2(new_n903), .ZN(new_n906));
  NAND2_X1  g481(.A1(new_n906), .A2(new_n896), .ZN(new_n907));
  NAND4_X1  g482(.A1(new_n907), .A2(KEYINPUT106), .A3(new_n900), .A4(new_n899), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n905), .A2(new_n908), .ZN(new_n909));
  XNOR2_X1  g484(.A(new_n909), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g485(.A1(new_n852), .A2(new_n600), .ZN(new_n911));
  XNOR2_X1  g486(.A(new_n620), .B(new_n861), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n609), .A2(G299), .ZN(new_n913));
  NAND4_X1  g488(.A1(new_n604), .A2(new_n566), .A3(new_n575), .A4(new_n608), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n915), .A2(KEYINPUT41), .ZN(new_n916));
  INV_X1    g491(.A(KEYINPUT108), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  NAND3_X1  g493(.A1(new_n915), .A2(KEYINPUT108), .A3(KEYINPUT41), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  INV_X1    g495(.A(KEYINPUT41), .ZN(new_n921));
  NAND3_X1  g496(.A1(new_n913), .A2(new_n921), .A3(new_n914), .ZN(new_n922));
  INV_X1    g497(.A(KEYINPUT107), .ZN(new_n923));
  XNOR2_X1  g498(.A(new_n922), .B(new_n923), .ZN(new_n924));
  NOR2_X1   g499(.A1(new_n920), .A2(new_n924), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n912), .A2(new_n925), .ZN(new_n926));
  INV_X1    g501(.A(new_n915), .ZN(new_n927));
  OAI21_X1  g502(.A(new_n926), .B1(new_n912), .B2(new_n927), .ZN(new_n928));
  XNOR2_X1  g503(.A(G303), .B(new_n703), .ZN(new_n929));
  AND2_X1   g504(.A1(new_n690), .A2(G290), .ZN(new_n930));
  NOR2_X1   g505(.A1(new_n690), .A2(G290), .ZN(new_n931));
  OAI21_X1  g506(.A(new_n929), .B1(new_n930), .B2(new_n931), .ZN(new_n932));
  XNOR2_X1  g507(.A(G288), .B(G290), .ZN(new_n933));
  XNOR2_X1  g508(.A(G303), .B(G305), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n933), .A2(new_n934), .ZN(new_n935));
  AOI21_X1  g510(.A(KEYINPUT42), .B1(new_n932), .B2(new_n935), .ZN(new_n936));
  AND3_X1   g511(.A1(new_n932), .A2(new_n935), .A3(KEYINPUT109), .ZN(new_n937));
  AOI21_X1  g512(.A(KEYINPUT109), .B1(new_n932), .B2(new_n935), .ZN(new_n938));
  NOR2_X1   g513(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  INV_X1    g514(.A(new_n939), .ZN(new_n940));
  AOI21_X1  g515(.A(new_n936), .B1(new_n940), .B2(KEYINPUT42), .ZN(new_n941));
  XOR2_X1   g516(.A(new_n928), .B(new_n941), .Z(new_n942));
  OAI21_X1  g517(.A(new_n911), .B1(new_n942), .B2(new_n600), .ZN(G295));
  OAI21_X1  g518(.A(new_n911), .B1(new_n942), .B2(new_n600), .ZN(G331));
  NAND3_X1  g519(.A1(new_n859), .A2(G301), .A3(new_n860), .ZN(new_n945));
  INV_X1    g520(.A(new_n945), .ZN(new_n946));
  AOI21_X1  g521(.A(G301), .B1(new_n859), .B2(new_n860), .ZN(new_n947));
  NOR3_X1   g522(.A1(new_n946), .A2(new_n947), .A3(G286), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n861), .A2(G171), .ZN(new_n949));
  AOI21_X1  g524(.A(G168), .B1(new_n949), .B2(new_n945), .ZN(new_n950));
  OAI21_X1  g525(.A(new_n927), .B1(new_n948), .B2(new_n950), .ZN(new_n951));
  INV_X1    g526(.A(KEYINPUT111), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n951), .A2(new_n952), .ZN(new_n953));
  OAI21_X1  g528(.A(G286), .B1(new_n946), .B2(new_n947), .ZN(new_n954));
  NAND3_X1  g529(.A1(new_n949), .A2(G168), .A3(new_n945), .ZN(new_n955));
  AOI21_X1  g530(.A(new_n915), .B1(new_n954), .B2(new_n955), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n956), .A2(KEYINPUT111), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n916), .A2(new_n922), .ZN(new_n958));
  INV_X1    g533(.A(KEYINPUT110), .ZN(new_n959));
  NAND4_X1  g534(.A1(new_n954), .A2(new_n958), .A3(new_n955), .A4(new_n959), .ZN(new_n960));
  NAND3_X1  g535(.A1(new_n954), .A2(new_n958), .A3(new_n955), .ZN(new_n961));
  NAND2_X1  g536(.A1(new_n961), .A2(KEYINPUT110), .ZN(new_n962));
  NAND4_X1  g537(.A1(new_n953), .A2(new_n957), .A3(new_n960), .A4(new_n962), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n963), .A2(new_n940), .ZN(new_n964));
  XNOR2_X1  g539(.A(new_n922), .B(KEYINPUT107), .ZN(new_n965));
  NAND3_X1  g540(.A1(new_n965), .A2(new_n918), .A3(new_n919), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n954), .A2(new_n955), .ZN(new_n967));
  INV_X1    g542(.A(new_n967), .ZN(new_n968));
  AOI21_X1  g543(.A(new_n956), .B1(new_n966), .B2(new_n968), .ZN(new_n969));
  AOI21_X1  g544(.A(G37), .B1(new_n969), .B2(new_n939), .ZN(new_n970));
  NAND3_X1  g545(.A1(new_n964), .A2(KEYINPUT43), .A3(new_n970), .ZN(new_n971));
  INV_X1    g546(.A(KEYINPUT43), .ZN(new_n972));
  OAI211_X1 g547(.A(new_n939), .B(new_n951), .C1(new_n925), .C2(new_n967), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n973), .A2(new_n900), .ZN(new_n974));
  NOR2_X1   g549(.A1(new_n969), .A2(new_n939), .ZN(new_n975));
  OAI21_X1  g550(.A(new_n972), .B1(new_n974), .B2(new_n975), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n971), .A2(new_n976), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n977), .A2(KEYINPUT44), .ZN(new_n978));
  NAND3_X1  g553(.A1(new_n964), .A2(new_n972), .A3(new_n970), .ZN(new_n979));
  OAI21_X1  g554(.A(KEYINPUT43), .B1(new_n974), .B2(new_n975), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n979), .A2(new_n980), .ZN(new_n981));
  INV_X1    g556(.A(KEYINPUT44), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n981), .A2(new_n982), .ZN(new_n983));
  NAND2_X1  g558(.A1(new_n978), .A2(new_n983), .ZN(G397));
  NOR2_X1   g559(.A1(G290), .A2(G1986), .ZN(new_n985));
  XOR2_X1   g560(.A(new_n985), .B(KEYINPUT112), .Z(new_n986));
  AOI22_X1  g561(.A1(new_n476), .A2(G137), .B1(G101), .B2(new_n461), .ZN(new_n987));
  AND2_X1   g562(.A1(new_n469), .A2(new_n470), .ZN(new_n988));
  OAI211_X1 g563(.A(new_n987), .B(G40), .C1(new_n988), .C2(new_n460), .ZN(new_n989));
  AOI21_X1  g564(.A(G1384), .B1(new_n502), .B2(new_n875), .ZN(new_n990));
  NOR3_X1   g565(.A1(new_n989), .A2(new_n990), .A3(KEYINPUT45), .ZN(new_n991));
  AND2_X1   g566(.A1(new_n986), .A2(new_n991), .ZN(new_n992));
  OR2_X1    g567(.A1(new_n992), .A2(KEYINPUT48), .ZN(new_n993));
  INV_X1    g568(.A(new_n991), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n814), .A2(G2067), .ZN(new_n995));
  INV_X1    g570(.A(G2067), .ZN(new_n996));
  NAND3_X1  g571(.A1(new_n809), .A2(new_n996), .A3(new_n813), .ZN(new_n997));
  AOI21_X1  g572(.A(new_n994), .B1(new_n995), .B2(new_n997), .ZN(new_n998));
  OR2_X1    g573(.A1(new_n998), .A2(KEYINPUT113), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n998), .A2(KEYINPUT113), .ZN(new_n1000));
  XOR2_X1   g575(.A(new_n776), .B(G1996), .Z(new_n1001));
  OAI211_X1 g576(.A(new_n999), .B(new_n1000), .C1(new_n994), .C2(new_n1001), .ZN(new_n1002));
  XNOR2_X1  g577(.A(new_n718), .B(new_n721), .ZN(new_n1003));
  XNOR2_X1  g578(.A(new_n1003), .B(KEYINPUT114), .ZN(new_n1004));
  AOI21_X1  g579(.A(new_n1002), .B1(new_n991), .B2(new_n1004), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n992), .A2(KEYINPUT48), .ZN(new_n1006));
  AND3_X1   g581(.A1(new_n993), .A2(new_n1005), .A3(new_n1006), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n719), .A2(new_n721), .ZN(new_n1008));
  OAI21_X1  g583(.A(new_n997), .B1(new_n1002), .B2(new_n1008), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n1009), .A2(new_n991), .ZN(new_n1010));
  NAND3_X1  g585(.A1(new_n995), .A2(new_n880), .A3(new_n997), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n1011), .A2(new_n991), .ZN(new_n1012));
  XOR2_X1   g587(.A(new_n1012), .B(KEYINPUT125), .Z(new_n1013));
  NOR2_X1   g588(.A1(new_n994), .A2(G1996), .ZN(new_n1014));
  XOR2_X1   g589(.A(new_n1014), .B(KEYINPUT46), .Z(new_n1015));
  NAND2_X1  g590(.A1(new_n1013), .A2(new_n1015), .ZN(new_n1016));
  INV_X1    g591(.A(KEYINPUT126), .ZN(new_n1017));
  XNOR2_X1  g592(.A(new_n1016), .B(new_n1017), .ZN(new_n1018));
  INV_X1    g593(.A(KEYINPUT47), .ZN(new_n1019));
  OAI21_X1  g594(.A(new_n1010), .B1(new_n1018), .B2(new_n1019), .ZN(new_n1020));
  AOI211_X1 g595(.A(new_n1007), .B(new_n1020), .C1(new_n1019), .C2(new_n1018), .ZN(new_n1021));
  INV_X1    g596(.A(KEYINPUT124), .ZN(new_n1022));
  INV_X1    g597(.A(G8), .ZN(new_n1023));
  INV_X1    g598(.A(G2084), .ZN(new_n1024));
  INV_X1    g599(.A(G40), .ZN(new_n1025));
  NOR3_X1   g600(.A1(new_n468), .A2(new_n471), .A3(new_n1025), .ZN(new_n1026));
  INV_X1    g601(.A(G1384), .ZN(new_n1027));
  NAND2_X1  g602(.A1(new_n876), .A2(new_n1027), .ZN(new_n1028));
  OAI21_X1  g603(.A(new_n1026), .B1(new_n1028), .B2(KEYINPUT50), .ZN(new_n1029));
  NAND3_X1  g604(.A1(new_n504), .A2(new_n1027), .A3(new_n506), .ZN(new_n1030));
  AOI21_X1  g605(.A(new_n1029), .B1(new_n1030), .B2(KEYINPUT50), .ZN(new_n1031));
  INV_X1    g606(.A(KEYINPUT45), .ZN(new_n1032));
  AOI21_X1  g607(.A(new_n989), .B1(new_n1028), .B2(new_n1032), .ZN(new_n1033));
  OAI21_X1  g608(.A(new_n1033), .B1(new_n1030), .B2(new_n1032), .ZN(new_n1034));
  AOI22_X1  g609(.A1(new_n1024), .A2(new_n1031), .B1(new_n1034), .B2(new_n789), .ZN(new_n1035));
  AOI21_X1  g610(.A(new_n1023), .B1(new_n1035), .B2(G168), .ZN(new_n1036));
  INV_X1    g611(.A(KEYINPUT51), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n1036), .A2(new_n1037), .ZN(new_n1038));
  INV_X1    g613(.A(new_n1038), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n1034), .A2(new_n789), .ZN(new_n1040));
  INV_X1    g615(.A(new_n1031), .ZN(new_n1041));
  OAI21_X1  g616(.A(new_n1040), .B1(new_n1041), .B2(G2084), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n1042), .A2(G286), .ZN(new_n1043));
  AOI21_X1  g618(.A(new_n1037), .B1(new_n1036), .B2(new_n1043), .ZN(new_n1044));
  OAI21_X1  g619(.A(KEYINPUT62), .B1(new_n1039), .B2(new_n1044), .ZN(new_n1045));
  OAI21_X1  g620(.A(G8), .B1(new_n1042), .B2(G286), .ZN(new_n1046));
  NOR2_X1   g621(.A1(new_n1035), .A2(G168), .ZN(new_n1047));
  OAI21_X1  g622(.A(KEYINPUT51), .B1(new_n1046), .B2(new_n1047), .ZN(new_n1048));
  INV_X1    g623(.A(KEYINPUT62), .ZN(new_n1049));
  NAND3_X1  g624(.A1(new_n1048), .A2(new_n1049), .A3(new_n1038), .ZN(new_n1050));
  NAND2_X1  g625(.A1(new_n1045), .A2(new_n1050), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n1026), .A2(new_n990), .ZN(new_n1052));
  NAND2_X1  g627(.A1(new_n1052), .A2(G8), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n1053), .A2(KEYINPUT115), .ZN(new_n1054));
  INV_X1    g629(.A(KEYINPUT115), .ZN(new_n1055));
  NAND3_X1  g630(.A1(new_n1052), .A2(new_n1055), .A3(G8), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n1054), .A2(new_n1056), .ZN(new_n1057));
  NAND3_X1  g632(.A1(new_n582), .A2(G1976), .A3(new_n584), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n1057), .A2(new_n1058), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n1059), .A2(KEYINPUT52), .ZN(new_n1060));
  INV_X1    g635(.A(G1976), .ZN(new_n1061));
  AOI21_X1  g636(.A(KEYINPUT52), .B1(G288), .B2(new_n1061), .ZN(new_n1062));
  NAND3_X1  g637(.A1(new_n1062), .A2(new_n1057), .A3(new_n1058), .ZN(new_n1063));
  OAI21_X1  g638(.A(G1981), .B1(new_n589), .B2(KEYINPUT116), .ZN(new_n1064));
  INV_X1    g639(.A(new_n1064), .ZN(new_n1065));
  NOR2_X1   g640(.A1(G305), .A2(new_n1065), .ZN(new_n1066));
  INV_X1    g641(.A(KEYINPUT49), .ZN(new_n1067));
  AOI21_X1  g642(.A(new_n1064), .B1(new_n590), .B2(new_n591), .ZN(new_n1068));
  OR3_X1    g643(.A1(new_n1066), .A2(new_n1067), .A3(new_n1068), .ZN(new_n1069));
  OAI21_X1  g644(.A(new_n1067), .B1(new_n1066), .B2(new_n1068), .ZN(new_n1070));
  NAND3_X1  g645(.A1(new_n1069), .A2(new_n1057), .A3(new_n1070), .ZN(new_n1071));
  NAND3_X1  g646(.A1(new_n1060), .A2(new_n1063), .A3(new_n1071), .ZN(new_n1072));
  NAND2_X1  g647(.A1(G303), .A2(G8), .ZN(new_n1073));
  XNOR2_X1  g648(.A(new_n1073), .B(KEYINPUT55), .ZN(new_n1074));
  INV_X1    g649(.A(new_n1074), .ZN(new_n1075));
  NOR2_X1   g650(.A1(new_n1028), .A2(new_n1032), .ZN(new_n1076));
  AOI21_X1  g651(.A(new_n1076), .B1(new_n1030), .B2(new_n1032), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n1077), .A2(new_n1026), .ZN(new_n1078));
  INV_X1    g653(.A(G1971), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n1078), .A2(new_n1079), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1031), .A2(new_n830), .ZN(new_n1081));
  AOI21_X1  g656(.A(new_n1023), .B1(new_n1080), .B2(new_n1081), .ZN(new_n1082));
  AOI21_X1  g657(.A(new_n1072), .B1(new_n1075), .B2(new_n1082), .ZN(new_n1083));
  AOI21_X1  g658(.A(G1971), .B1(new_n1077), .B2(new_n1026), .ZN(new_n1084));
  AOI21_X1  g659(.A(new_n989), .B1(new_n1028), .B2(KEYINPUT50), .ZN(new_n1085));
  OAI21_X1  g660(.A(new_n1085), .B1(new_n1030), .B2(KEYINPUT50), .ZN(new_n1086));
  NOR2_X1   g661(.A1(new_n1086), .A2(G2090), .ZN(new_n1087));
  OAI21_X1  g662(.A(KEYINPUT118), .B1(new_n1084), .B2(new_n1087), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n1088), .A2(G8), .ZN(new_n1089));
  NOR3_X1   g664(.A1(new_n1084), .A2(new_n1087), .A3(KEYINPUT118), .ZN(new_n1090));
  OAI21_X1  g665(.A(new_n1074), .B1(new_n1089), .B2(new_n1090), .ZN(new_n1091));
  INV_X1    g666(.A(KEYINPUT53), .ZN(new_n1092));
  OAI21_X1  g667(.A(new_n1092), .B1(new_n1078), .B2(G2078), .ZN(new_n1093));
  OR2_X1    g668(.A1(new_n1031), .A2(G1961), .ZN(new_n1094));
  NOR2_X1   g669(.A1(new_n1092), .A2(G2078), .ZN(new_n1095));
  OAI211_X1 g670(.A(new_n1095), .B(new_n1033), .C1(new_n1030), .C2(new_n1032), .ZN(new_n1096));
  NAND3_X1  g671(.A1(new_n1093), .A2(new_n1094), .A3(new_n1096), .ZN(new_n1097));
  AND2_X1   g672(.A1(new_n1097), .A2(G171), .ZN(new_n1098));
  NAND3_X1  g673(.A1(new_n1083), .A2(new_n1091), .A3(new_n1098), .ZN(new_n1099));
  OAI21_X1  g674(.A(new_n1022), .B1(new_n1051), .B2(new_n1099), .ZN(new_n1100));
  AND3_X1   g675(.A1(new_n1083), .A2(new_n1091), .A3(new_n1098), .ZN(new_n1101));
  NAND4_X1  g676(.A1(new_n1101), .A2(KEYINPUT124), .A3(new_n1050), .A4(new_n1045), .ZN(new_n1102));
  NOR3_X1   g677(.A1(new_n1035), .A2(new_n1023), .A3(G286), .ZN(new_n1103));
  NAND3_X1  g678(.A1(new_n1083), .A2(new_n1091), .A3(new_n1103), .ZN(new_n1104));
  INV_X1    g679(.A(KEYINPUT63), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n1104), .A2(new_n1105), .ZN(new_n1106));
  XNOR2_X1  g681(.A(new_n1072), .B(KEYINPUT117), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n1075), .A2(new_n1082), .ZN(new_n1108));
  AND3_X1   g683(.A1(new_n1108), .A2(new_n1103), .A3(KEYINPUT63), .ZN(new_n1109));
  OR2_X1    g684(.A1(new_n1075), .A2(new_n1082), .ZN(new_n1110));
  NAND3_X1  g685(.A1(new_n1107), .A2(new_n1109), .A3(new_n1110), .ZN(new_n1111));
  NAND2_X1  g686(.A1(new_n1106), .A2(new_n1111), .ZN(new_n1112));
  INV_X1    g687(.A(new_n1108), .ZN(new_n1113));
  NAND3_X1  g688(.A1(new_n1071), .A2(new_n1061), .A3(new_n690), .ZN(new_n1114));
  OAI21_X1  g689(.A(new_n1114), .B1(G1981), .B2(G305), .ZN(new_n1115));
  AOI22_X1  g690(.A1(new_n1107), .A2(new_n1113), .B1(new_n1057), .B2(new_n1115), .ZN(new_n1116));
  NAND4_X1  g691(.A1(new_n1100), .A2(new_n1102), .A3(new_n1112), .A4(new_n1116), .ZN(new_n1117));
  XNOR2_X1  g692(.A(KEYINPUT56), .B(G2072), .ZN(new_n1118));
  NAND3_X1  g693(.A1(new_n1077), .A2(new_n1026), .A3(new_n1118), .ZN(new_n1119));
  INV_X1    g694(.A(G1956), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n1086), .A2(new_n1120), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n1119), .A2(new_n1121), .ZN(new_n1122));
  XNOR2_X1  g697(.A(KEYINPUT119), .B(KEYINPUT57), .ZN(new_n1123));
  AND3_X1   g698(.A1(new_n566), .A2(new_n575), .A3(new_n1123), .ZN(new_n1124));
  AOI21_X1  g699(.A(new_n1123), .B1(new_n566), .B2(new_n575), .ZN(new_n1125));
  NOR2_X1   g700(.A1(new_n1124), .A2(new_n1125), .ZN(new_n1126));
  NAND2_X1  g701(.A1(new_n1122), .A2(new_n1126), .ZN(new_n1127));
  OAI22_X1  g702(.A1(new_n1031), .A2(G1348), .B1(G2067), .B2(new_n1052), .ZN(new_n1128));
  INV_X1    g703(.A(new_n1128), .ZN(new_n1129));
  OAI21_X1  g704(.A(new_n1127), .B1(new_n1129), .B2(new_n609), .ZN(new_n1130));
  OAI211_X1 g705(.A(new_n1119), .B(new_n1121), .C1(new_n1124), .C2(new_n1125), .ZN(new_n1131));
  NAND2_X1  g706(.A1(new_n1130), .A2(new_n1131), .ZN(new_n1132));
  NAND2_X1  g707(.A1(new_n1129), .A2(KEYINPUT60), .ZN(new_n1133));
  XOR2_X1   g708(.A(new_n1133), .B(new_n609), .Z(new_n1134));
  OAI21_X1  g709(.A(new_n1134), .B1(KEYINPUT60), .B2(new_n1129), .ZN(new_n1135));
  INV_X1    g710(.A(KEYINPUT61), .ZN(new_n1136));
  AND3_X1   g711(.A1(new_n1127), .A2(new_n1136), .A3(new_n1131), .ZN(new_n1137));
  AOI21_X1  g712(.A(new_n1136), .B1(new_n1127), .B2(new_n1131), .ZN(new_n1138));
  NOR2_X1   g713(.A1(new_n1137), .A2(new_n1138), .ZN(new_n1139));
  INV_X1    g714(.A(KEYINPUT121), .ZN(new_n1140));
  INV_X1    g715(.A(new_n1076), .ZN(new_n1141));
  NOR2_X1   g716(.A1(new_n989), .A2(G1996), .ZN(new_n1142));
  AND3_X1   g717(.A1(new_n497), .A2(new_n505), .A3(new_n502), .ZN(new_n1143));
  AOI21_X1  g718(.A(new_n505), .B1(new_n497), .B2(new_n502), .ZN(new_n1144));
  NOR3_X1   g719(.A1(new_n1143), .A2(new_n1144), .A3(G1384), .ZN(new_n1145));
  OAI211_X1 g720(.A(new_n1141), .B(new_n1142), .C1(new_n1145), .C2(KEYINPUT45), .ZN(new_n1146));
  INV_X1    g721(.A(KEYINPUT120), .ZN(new_n1147));
  NAND2_X1  g722(.A1(new_n1146), .A2(new_n1147), .ZN(new_n1148));
  NAND3_X1  g723(.A1(new_n1077), .A2(KEYINPUT120), .A3(new_n1142), .ZN(new_n1149));
  NAND2_X1  g724(.A1(new_n1148), .A2(new_n1149), .ZN(new_n1150));
  XOR2_X1   g725(.A(KEYINPUT58), .B(G1341), .Z(new_n1151));
  AND2_X1   g726(.A1(new_n1052), .A2(new_n1151), .ZN(new_n1152));
  INV_X1    g727(.A(new_n1152), .ZN(new_n1153));
  AOI21_X1  g728(.A(new_n1140), .B1(new_n1150), .B2(new_n1153), .ZN(new_n1154));
  AOI211_X1 g729(.A(KEYINPUT121), .B(new_n1152), .C1(new_n1148), .C2(new_n1149), .ZN(new_n1155));
  OAI21_X1  g730(.A(new_n556), .B1(new_n1154), .B2(new_n1155), .ZN(new_n1156));
  NAND2_X1  g731(.A1(new_n1156), .A2(KEYINPUT59), .ZN(new_n1157));
  INV_X1    g732(.A(KEYINPUT59), .ZN(new_n1158));
  OAI211_X1 g733(.A(new_n1158), .B(new_n556), .C1(new_n1154), .C2(new_n1155), .ZN(new_n1159));
  AOI21_X1  g734(.A(new_n1139), .B1(new_n1157), .B2(new_n1159), .ZN(new_n1160));
  OAI21_X1  g735(.A(new_n1135), .B1(new_n1160), .B2(KEYINPUT122), .ZN(new_n1161));
  INV_X1    g736(.A(KEYINPUT122), .ZN(new_n1162));
  AOI211_X1 g737(.A(new_n1162), .B(new_n1139), .C1(new_n1157), .C2(new_n1159), .ZN(new_n1163));
  OAI21_X1  g738(.A(new_n1132), .B1(new_n1161), .B2(new_n1163), .ZN(new_n1164));
  INV_X1    g739(.A(KEYINPUT54), .ZN(new_n1165));
  NAND3_X1  g740(.A1(new_n1141), .A2(new_n1095), .A3(new_n1033), .ZN(new_n1166));
  NAND3_X1  g741(.A1(new_n1093), .A2(new_n1094), .A3(new_n1166), .ZN(new_n1167));
  AOI21_X1  g742(.A(new_n1165), .B1(new_n1167), .B2(G171), .ZN(new_n1168));
  OAI21_X1  g743(.A(new_n1168), .B1(G171), .B2(new_n1097), .ZN(new_n1169));
  NAND2_X1  g744(.A1(new_n1048), .A2(new_n1038), .ZN(new_n1170));
  NAND4_X1  g745(.A1(new_n1169), .A2(new_n1170), .A3(new_n1091), .A4(new_n1083), .ZN(new_n1171));
  NOR2_X1   g746(.A1(new_n1167), .A2(G171), .ZN(new_n1172));
  OAI21_X1  g747(.A(new_n1165), .B1(new_n1098), .B2(new_n1172), .ZN(new_n1173));
  OR2_X1    g748(.A1(new_n1173), .A2(KEYINPUT123), .ZN(new_n1174));
  NAND2_X1  g749(.A1(new_n1173), .A2(KEYINPUT123), .ZN(new_n1175));
  AOI21_X1  g750(.A(new_n1171), .B1(new_n1174), .B2(new_n1175), .ZN(new_n1176));
  AOI21_X1  g751(.A(new_n1117), .B1(new_n1164), .B2(new_n1176), .ZN(new_n1177));
  AOI21_X1  g752(.A(new_n986), .B1(G1986), .B2(G290), .ZN(new_n1178));
  OAI21_X1  g753(.A(new_n1005), .B1(new_n1178), .B2(new_n994), .ZN(new_n1179));
  OAI21_X1  g754(.A(new_n1021), .B1(new_n1177), .B2(new_n1179), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g755(.A(KEYINPUT127), .ZN(new_n1182));
  NOR3_X1   g756(.A1(G229), .A2(new_n458), .A3(G227), .ZN(new_n1183));
  AOI21_X1  g757(.A(new_n1182), .B1(new_n655), .B2(new_n1183), .ZN(new_n1184));
  OAI211_X1 g758(.A(new_n1183), .B(new_n1182), .C1(new_n654), .C2(new_n653), .ZN(new_n1185));
  INV_X1    g759(.A(new_n1185), .ZN(new_n1186));
  NOR2_X1   g760(.A1(new_n1184), .A2(new_n1186), .ZN(new_n1187));
  AND3_X1   g761(.A1(new_n981), .A2(new_n1187), .A3(new_n909), .ZN(G308));
  NAND3_X1  g762(.A1(new_n981), .A2(new_n1187), .A3(new_n909), .ZN(G225));
endmodule


