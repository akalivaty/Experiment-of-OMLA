//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 0 1 0 1 0 0 0 1 0 1 1 0 1 0 1 0 1 1 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 0 0 1 1 1 1 1 0 0 0 0 0 0 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:19:05 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n636, new_n637,
    new_n638, new_n640, new_n641, new_n642, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n729, new_n730, new_n731, new_n732, new_n733, new_n734, new_n735,
    new_n737, new_n738, new_n739, new_n740, new_n741, new_n743, new_n744,
    new_n746, new_n747, new_n748, new_n749, new_n750, new_n751, new_n752,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n772, new_n773, new_n774, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n814, new_n815, new_n817, new_n818, new_n819, new_n821, new_n822,
    new_n823, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n872, new_n873, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n888, new_n889, new_n891, new_n892,
    new_n893, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n911, new_n912, new_n913, new_n914, new_n916, new_n917,
    new_n918, new_n919, new_n920, new_n921, new_n923, new_n924;
  XNOR2_X1  g000(.A(KEYINPUT27), .B(G183gat), .ZN(new_n202));
  INV_X1    g001(.A(G190gat), .ZN(new_n203));
  NAND2_X1  g002(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  NAND2_X1  g003(.A1(new_n204), .A2(KEYINPUT28), .ZN(new_n205));
  NOR2_X1   g004(.A1(G169gat), .A2(G176gat), .ZN(new_n206));
  INV_X1    g005(.A(KEYINPUT26), .ZN(new_n207));
  OAI21_X1  g006(.A(KEYINPUT65), .B1(new_n206), .B2(new_n207), .ZN(new_n208));
  NAND2_X1  g007(.A1(G169gat), .A2(G176gat), .ZN(new_n209));
  NAND2_X1  g008(.A1(new_n206), .A2(new_n207), .ZN(new_n210));
  INV_X1    g009(.A(KEYINPUT65), .ZN(new_n211));
  OAI211_X1 g010(.A(new_n211), .B(KEYINPUT26), .C1(G169gat), .C2(G176gat), .ZN(new_n212));
  NAND4_X1  g011(.A1(new_n208), .A2(new_n209), .A3(new_n210), .A4(new_n212), .ZN(new_n213));
  NAND2_X1  g012(.A1(G183gat), .A2(G190gat), .ZN(new_n214));
  INV_X1    g013(.A(KEYINPUT28), .ZN(new_n215));
  NAND3_X1  g014(.A1(new_n202), .A2(new_n215), .A3(new_n203), .ZN(new_n216));
  NAND4_X1  g015(.A1(new_n205), .A2(new_n213), .A3(new_n214), .A4(new_n216), .ZN(new_n217));
  INV_X1    g016(.A(G169gat), .ZN(new_n218));
  INV_X1    g017(.A(G176gat), .ZN(new_n219));
  NAND3_X1  g018(.A1(new_n218), .A2(new_n219), .A3(KEYINPUT23), .ZN(new_n220));
  INV_X1    g019(.A(KEYINPUT23), .ZN(new_n221));
  OAI21_X1  g020(.A(new_n221), .B1(G169gat), .B2(G176gat), .ZN(new_n222));
  NAND3_X1  g021(.A1(new_n220), .A2(new_n222), .A3(new_n209), .ZN(new_n223));
  INV_X1    g022(.A(new_n223), .ZN(new_n224));
  INV_X1    g023(.A(KEYINPUT24), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n214), .A2(new_n225), .ZN(new_n226));
  NAND3_X1  g025(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n227));
  OAI211_X1 g026(.A(new_n226), .B(new_n227), .C1(G183gat), .C2(G190gat), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n224), .A2(new_n228), .ZN(new_n229));
  INV_X1    g028(.A(KEYINPUT25), .ZN(new_n230));
  OAI21_X1  g029(.A(new_n230), .B1(new_n223), .B2(KEYINPUT64), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n229), .A2(new_n231), .ZN(new_n232));
  NAND4_X1  g031(.A1(new_n224), .A2(new_n228), .A3(KEYINPUT64), .A4(new_n230), .ZN(new_n233));
  NAND3_X1  g032(.A1(new_n217), .A2(new_n232), .A3(new_n233), .ZN(new_n234));
  INV_X1    g033(.A(KEYINPUT29), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n234), .A2(new_n235), .ZN(new_n236));
  INV_X1    g035(.A(G226gat), .ZN(new_n237));
  INV_X1    g036(.A(G233gat), .ZN(new_n238));
  OAI21_X1  g037(.A(new_n236), .B1(new_n237), .B2(new_n238), .ZN(new_n239));
  NOR2_X1   g038(.A1(new_n237), .A2(new_n238), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n234), .A2(new_n240), .ZN(new_n241));
  NAND2_X1  g040(.A1(G211gat), .A2(G218gat), .ZN(new_n242));
  INV_X1    g041(.A(KEYINPUT22), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n242), .A2(new_n243), .ZN(new_n244));
  NOR2_X1   g043(.A1(G197gat), .A2(G204gat), .ZN(new_n245));
  AND2_X1   g044(.A1(G197gat), .A2(G204gat), .ZN(new_n246));
  OAI21_X1  g045(.A(new_n244), .B1(new_n245), .B2(new_n246), .ZN(new_n247));
  XOR2_X1   g046(.A(G211gat), .B(G218gat), .Z(new_n248));
  NAND2_X1  g047(.A1(new_n247), .A2(new_n248), .ZN(new_n249));
  XNOR2_X1  g048(.A(G211gat), .B(G218gat), .ZN(new_n250));
  XNOR2_X1  g049(.A(G197gat), .B(G204gat), .ZN(new_n251));
  NAND3_X1  g050(.A1(new_n250), .A2(new_n251), .A3(new_n244), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n249), .A2(new_n252), .ZN(new_n253));
  NAND3_X1  g052(.A1(new_n239), .A2(new_n241), .A3(new_n253), .ZN(new_n254));
  INV_X1    g053(.A(KEYINPUT68), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n253), .A2(new_n255), .ZN(new_n256));
  NAND3_X1  g055(.A1(new_n249), .A2(KEYINPUT68), .A3(new_n252), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  INV_X1    g057(.A(new_n258), .ZN(new_n259));
  INV_X1    g058(.A(new_n241), .ZN(new_n260));
  XOR2_X1   g059(.A(KEYINPUT69), .B(KEYINPUT29), .Z(new_n261));
  AOI21_X1  g060(.A(new_n240), .B1(new_n234), .B2(new_n261), .ZN(new_n262));
  OAI21_X1  g061(.A(new_n259), .B1(new_n260), .B2(new_n262), .ZN(new_n263));
  NAND2_X1  g062(.A1(new_n254), .A2(new_n263), .ZN(new_n264));
  XNOR2_X1  g063(.A(KEYINPUT70), .B(G8gat), .ZN(new_n265));
  XNOR2_X1  g064(.A(new_n265), .B(G36gat), .ZN(new_n266));
  XOR2_X1   g065(.A(G64gat), .B(G92gat), .Z(new_n267));
  XNOR2_X1  g066(.A(new_n266), .B(new_n267), .ZN(new_n268));
  OR2_X1    g067(.A1(new_n264), .A2(new_n268), .ZN(new_n269));
  INV_X1    g068(.A(KEYINPUT30), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n264), .A2(new_n268), .ZN(new_n272));
  OR3_X1    g071(.A1(new_n264), .A2(new_n270), .A3(new_n268), .ZN(new_n273));
  NAND3_X1  g072(.A1(new_n271), .A2(new_n272), .A3(new_n273), .ZN(new_n274));
  XNOR2_X1  g073(.A(G127gat), .B(G134gat), .ZN(new_n275));
  INV_X1    g074(.A(KEYINPUT1), .ZN(new_n276));
  INV_X1    g075(.A(G113gat), .ZN(new_n277));
  NOR2_X1   g076(.A1(new_n277), .A2(G120gat), .ZN(new_n278));
  INV_X1    g077(.A(G120gat), .ZN(new_n279));
  NOR2_X1   g078(.A1(new_n279), .A2(G113gat), .ZN(new_n280));
  OAI211_X1 g079(.A(new_n275), .B(new_n276), .C1(new_n278), .C2(new_n280), .ZN(new_n281));
  XNOR2_X1  g080(.A(G113gat), .B(G120gat), .ZN(new_n282));
  INV_X1    g081(.A(G134gat), .ZN(new_n283));
  AND2_X1   g082(.A1(new_n283), .A2(G127gat), .ZN(new_n284));
  NOR2_X1   g083(.A1(new_n283), .A2(G127gat), .ZN(new_n285));
  OAI22_X1  g084(.A1(new_n282), .A2(KEYINPUT1), .B1(new_n284), .B2(new_n285), .ZN(new_n286));
  AND2_X1   g085(.A1(new_n281), .A2(new_n286), .ZN(new_n287));
  INV_X1    g086(.A(KEYINPUT73), .ZN(new_n288));
  INV_X1    g087(.A(G148gat), .ZN(new_n289));
  INV_X1    g088(.A(KEYINPUT72), .ZN(new_n290));
  INV_X1    g089(.A(G141gat), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  NAND2_X1  g091(.A1(KEYINPUT72), .A2(G141gat), .ZN(new_n293));
  AOI21_X1  g092(.A(new_n289), .B1(new_n292), .B2(new_n293), .ZN(new_n294));
  NOR2_X1   g093(.A1(new_n291), .A2(G148gat), .ZN(new_n295));
  OAI21_X1  g094(.A(new_n288), .B1(new_n294), .B2(new_n295), .ZN(new_n296));
  INV_X1    g095(.A(G155gat), .ZN(new_n297));
  NOR2_X1   g096(.A1(new_n297), .A2(G162gat), .ZN(new_n298));
  INV_X1    g097(.A(G162gat), .ZN(new_n299));
  NOR2_X1   g098(.A1(new_n299), .A2(G155gat), .ZN(new_n300));
  OAI21_X1  g099(.A(KEYINPUT74), .B1(new_n298), .B2(new_n300), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n299), .A2(G155gat), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n297), .A2(G162gat), .ZN(new_n303));
  INV_X1    g102(.A(KEYINPUT74), .ZN(new_n304));
  NAND3_X1  g103(.A1(new_n302), .A2(new_n303), .A3(new_n304), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n301), .A2(new_n305), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n297), .A2(KEYINPUT75), .ZN(new_n307));
  INV_X1    g106(.A(KEYINPUT75), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n308), .A2(G155gat), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n307), .A2(new_n309), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n299), .A2(KEYINPUT76), .ZN(new_n311));
  INV_X1    g110(.A(KEYINPUT76), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n312), .A2(G162gat), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n311), .A2(new_n313), .ZN(new_n314));
  OAI21_X1  g113(.A(KEYINPUT2), .B1(new_n310), .B2(new_n314), .ZN(new_n315));
  AND2_X1   g114(.A1(KEYINPUT72), .A2(G141gat), .ZN(new_n316));
  NOR2_X1   g115(.A1(KEYINPUT72), .A2(G141gat), .ZN(new_n317));
  OAI21_X1  g116(.A(G148gat), .B1(new_n316), .B2(new_n317), .ZN(new_n318));
  INV_X1    g117(.A(new_n295), .ZN(new_n319));
  NAND3_X1  g118(.A1(new_n318), .A2(KEYINPUT73), .A3(new_n319), .ZN(new_n320));
  NAND4_X1  g119(.A1(new_n296), .A2(new_n306), .A3(new_n315), .A4(new_n320), .ZN(new_n321));
  XOR2_X1   g120(.A(KEYINPUT71), .B(KEYINPUT2), .Z(new_n322));
  XNOR2_X1  g121(.A(G141gat), .B(G148gat), .ZN(new_n323));
  OAI22_X1  g122(.A1(new_n322), .A2(new_n323), .B1(new_n298), .B2(new_n300), .ZN(new_n324));
  AOI21_X1  g123(.A(new_n287), .B1(new_n321), .B2(new_n324), .ZN(new_n325));
  NAND3_X1  g124(.A1(new_n321), .A2(new_n324), .A3(new_n287), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n326), .A2(KEYINPUT78), .ZN(new_n327));
  INV_X1    g126(.A(KEYINPUT78), .ZN(new_n328));
  NAND4_X1  g127(.A1(new_n321), .A2(new_n328), .A3(new_n287), .A4(new_n324), .ZN(new_n329));
  AOI21_X1  g128(.A(new_n325), .B1(new_n327), .B2(new_n329), .ZN(new_n330));
  NAND2_X1  g129(.A1(G225gat), .A2(G233gat), .ZN(new_n331));
  XNOR2_X1  g130(.A(new_n331), .B(KEYINPUT77), .ZN(new_n332));
  INV_X1    g131(.A(new_n332), .ZN(new_n333));
  OAI21_X1  g132(.A(KEYINPUT5), .B1(new_n330), .B2(new_n333), .ZN(new_n334));
  NAND2_X1  g133(.A1(new_n334), .A2(KEYINPUT79), .ZN(new_n335));
  INV_X1    g134(.A(KEYINPUT79), .ZN(new_n336));
  OAI211_X1 g135(.A(new_n336), .B(KEYINPUT5), .C1(new_n330), .C2(new_n333), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n335), .A2(new_n337), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n321), .A2(new_n324), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n339), .A2(KEYINPUT3), .ZN(new_n340));
  INV_X1    g139(.A(new_n287), .ZN(new_n341));
  INV_X1    g140(.A(KEYINPUT3), .ZN(new_n342));
  NAND3_X1  g141(.A1(new_n321), .A2(new_n342), .A3(new_n324), .ZN(new_n343));
  NAND3_X1  g142(.A1(new_n340), .A2(new_n341), .A3(new_n343), .ZN(new_n344));
  INV_X1    g143(.A(new_n326), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n345), .A2(KEYINPUT4), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n344), .A2(new_n346), .ZN(new_n347));
  AOI21_X1  g146(.A(KEYINPUT4), .B1(new_n327), .B2(new_n329), .ZN(new_n348));
  NOR3_X1   g147(.A1(new_n347), .A2(new_n332), .A3(new_n348), .ZN(new_n349));
  INV_X1    g148(.A(new_n349), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n338), .A2(new_n350), .ZN(new_n351));
  AOI21_X1  g150(.A(new_n345), .B1(new_n344), .B2(KEYINPUT4), .ZN(new_n352));
  AND3_X1   g151(.A1(new_n327), .A2(KEYINPUT4), .A3(new_n329), .ZN(new_n353));
  NOR4_X1   g152(.A1(new_n352), .A2(new_n353), .A3(KEYINPUT5), .A4(new_n332), .ZN(new_n354));
  INV_X1    g153(.A(new_n354), .ZN(new_n355));
  XNOR2_X1  g154(.A(G1gat), .B(G29gat), .ZN(new_n356));
  INV_X1    g155(.A(G85gat), .ZN(new_n357));
  XNOR2_X1  g156(.A(new_n356), .B(new_n357), .ZN(new_n358));
  XNOR2_X1  g157(.A(KEYINPUT0), .B(G57gat), .ZN(new_n359));
  XOR2_X1   g158(.A(new_n358), .B(new_n359), .Z(new_n360));
  INV_X1    g159(.A(new_n360), .ZN(new_n361));
  NAND3_X1  g160(.A1(new_n351), .A2(new_n355), .A3(new_n361), .ZN(new_n362));
  AOI21_X1  g161(.A(new_n349), .B1(new_n335), .B2(new_n337), .ZN(new_n363));
  OAI21_X1  g162(.A(new_n360), .B1(new_n363), .B2(new_n354), .ZN(new_n364));
  XNOR2_X1  g163(.A(KEYINPUT80), .B(KEYINPUT6), .ZN(new_n365));
  INV_X1    g164(.A(new_n365), .ZN(new_n366));
  NAND3_X1  g165(.A1(new_n362), .A2(new_n364), .A3(new_n366), .ZN(new_n367));
  OAI211_X1 g166(.A(new_n360), .B(new_n365), .C1(new_n363), .C2(new_n354), .ZN(new_n368));
  AOI21_X1  g167(.A(new_n274), .B1(new_n367), .B2(new_n368), .ZN(new_n369));
  XOR2_X1   g168(.A(G15gat), .B(G43gat), .Z(new_n370));
  XNOR2_X1  g169(.A(G71gat), .B(G99gat), .ZN(new_n371));
  XNOR2_X1  g170(.A(new_n370), .B(new_n371), .ZN(new_n372));
  NAND2_X1  g171(.A1(G227gat), .A2(G233gat), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n234), .A2(new_n341), .ZN(new_n374));
  NAND4_X1  g173(.A1(new_n217), .A2(new_n232), .A3(new_n287), .A4(new_n233), .ZN(new_n375));
  AOI21_X1  g174(.A(new_n373), .B1(new_n374), .B2(new_n375), .ZN(new_n376));
  OAI21_X1  g175(.A(new_n372), .B1(new_n376), .B2(KEYINPUT33), .ZN(new_n377));
  INV_X1    g176(.A(KEYINPUT32), .ZN(new_n378));
  OAI22_X1  g177(.A1(new_n377), .A2(KEYINPUT66), .B1(new_n378), .B2(new_n376), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n372), .A2(KEYINPUT33), .ZN(new_n380));
  NOR3_X1   g179(.A1(new_n376), .A2(new_n378), .A3(new_n380), .ZN(new_n381));
  INV_X1    g180(.A(KEYINPUT66), .ZN(new_n382));
  OAI21_X1  g181(.A(new_n381), .B1(new_n377), .B2(new_n382), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n379), .A2(new_n383), .ZN(new_n384));
  NAND3_X1  g183(.A1(new_n374), .A2(new_n373), .A3(new_n375), .ZN(new_n385));
  XNOR2_X1  g184(.A(new_n385), .B(KEYINPUT34), .ZN(new_n386));
  INV_X1    g185(.A(new_n386), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n384), .A2(new_n387), .ZN(new_n388));
  NAND3_X1  g187(.A1(new_n379), .A2(new_n383), .A3(new_n386), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n388), .A2(new_n389), .ZN(new_n390));
  NAND2_X1  g189(.A1(G228gat), .A2(G233gat), .ZN(new_n391));
  XOR2_X1   g190(.A(new_n391), .B(KEYINPUT81), .Z(new_n392));
  INV_X1    g191(.A(new_n392), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n343), .A2(new_n261), .ZN(new_n394));
  INV_X1    g193(.A(new_n253), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n394), .A2(new_n395), .ZN(new_n396));
  AOI21_X1  g195(.A(KEYINPUT3), .B1(new_n253), .B2(new_n261), .ZN(new_n397));
  AOI21_X1  g196(.A(new_n397), .B1(new_n324), .B2(new_n321), .ZN(new_n398));
  INV_X1    g197(.A(new_n398), .ZN(new_n399));
  AOI21_X1  g198(.A(new_n393), .B1(new_n396), .B2(new_n399), .ZN(new_n400));
  AOI21_X1  g199(.A(new_n258), .B1(new_n343), .B2(new_n261), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n253), .A2(new_n235), .ZN(new_n402));
  AOI22_X1  g201(.A1(new_n342), .A2(new_n402), .B1(new_n321), .B2(new_n324), .ZN(new_n403));
  NOR3_X1   g202(.A1(new_n401), .A2(new_n403), .A3(new_n391), .ZN(new_n404));
  OAI21_X1  g203(.A(G22gat), .B1(new_n400), .B2(new_n404), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n394), .A2(new_n259), .ZN(new_n406));
  INV_X1    g205(.A(new_n403), .ZN(new_n407));
  NAND4_X1  g206(.A1(new_n406), .A2(G228gat), .A3(G233gat), .A4(new_n407), .ZN(new_n408));
  AOI21_X1  g207(.A(new_n253), .B1(new_n343), .B2(new_n261), .ZN(new_n409));
  OAI21_X1  g208(.A(new_n392), .B1(new_n409), .B2(new_n398), .ZN(new_n410));
  INV_X1    g209(.A(G22gat), .ZN(new_n411));
  NAND3_X1  g210(.A1(new_n408), .A2(new_n410), .A3(new_n411), .ZN(new_n412));
  NAND3_X1  g211(.A1(new_n405), .A2(KEYINPUT82), .A3(new_n412), .ZN(new_n413));
  XOR2_X1   g212(.A(KEYINPUT31), .B(G50gat), .Z(new_n414));
  XNOR2_X1  g213(.A(G78gat), .B(G106gat), .ZN(new_n415));
  XNOR2_X1  g214(.A(new_n414), .B(new_n415), .ZN(new_n416));
  INV_X1    g215(.A(KEYINPUT82), .ZN(new_n417));
  NAND4_X1  g216(.A1(new_n408), .A2(new_n410), .A3(new_n417), .A4(new_n411), .ZN(new_n418));
  NAND3_X1  g217(.A1(new_n413), .A2(new_n416), .A3(new_n418), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n419), .A2(KEYINPUT83), .ZN(new_n420));
  INV_X1    g219(.A(KEYINPUT83), .ZN(new_n421));
  NAND4_X1  g220(.A1(new_n413), .A2(new_n421), .A3(new_n416), .A4(new_n418), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n420), .A2(new_n422), .ZN(new_n423));
  INV_X1    g222(.A(new_n412), .ZN(new_n424));
  NOR2_X1   g223(.A1(new_n424), .A2(new_n416), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n425), .A2(new_n405), .ZN(new_n426));
  AOI21_X1  g225(.A(new_n390), .B1(new_n423), .B2(new_n426), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n369), .A2(new_n427), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n428), .A2(KEYINPUT35), .ZN(new_n429));
  INV_X1    g228(.A(KEYINPUT67), .ZN(new_n430));
  NAND3_X1  g229(.A1(new_n384), .A2(new_n387), .A3(new_n430), .ZN(new_n431));
  NAND3_X1  g230(.A1(new_n388), .A2(KEYINPUT67), .A3(new_n389), .ZN(new_n432));
  AOI22_X1  g231(.A1(new_n423), .A2(new_n426), .B1(new_n431), .B2(new_n432), .ZN(new_n433));
  INV_X1    g232(.A(KEYINPUT35), .ZN(new_n434));
  NAND3_X1  g233(.A1(new_n433), .A2(new_n369), .A3(new_n434), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n429), .A2(new_n435), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n367), .A2(new_n368), .ZN(new_n437));
  INV_X1    g236(.A(new_n274), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n437), .A2(new_n438), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n423), .A2(new_n426), .ZN(new_n440));
  INV_X1    g239(.A(new_n440), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n439), .A2(new_n441), .ZN(new_n442));
  OAI21_X1  g241(.A(new_n332), .B1(new_n352), .B2(new_n353), .ZN(new_n443));
  INV_X1    g242(.A(KEYINPUT84), .ZN(new_n444));
  AOI211_X1 g243(.A(new_n332), .B(new_n325), .C1(new_n327), .C2(new_n329), .ZN(new_n445));
  INV_X1    g244(.A(KEYINPUT39), .ZN(new_n446));
  OAI21_X1  g245(.A(new_n444), .B1(new_n445), .B2(new_n446), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n330), .A2(new_n333), .ZN(new_n448));
  NAND3_X1  g247(.A1(new_n448), .A2(KEYINPUT84), .A3(KEYINPUT39), .ZN(new_n449));
  NAND3_X1  g248(.A1(new_n443), .A2(new_n447), .A3(new_n449), .ZN(new_n450));
  OAI211_X1 g249(.A(new_n446), .B(new_n332), .C1(new_n352), .C2(new_n353), .ZN(new_n451));
  NAND4_X1  g250(.A1(new_n450), .A2(KEYINPUT40), .A3(new_n361), .A4(new_n451), .ZN(new_n452));
  AND2_X1   g251(.A1(new_n364), .A2(new_n452), .ZN(new_n453));
  INV_X1    g252(.A(KEYINPUT40), .ZN(new_n454));
  AND3_X1   g253(.A1(new_n443), .A2(new_n447), .A3(new_n449), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n451), .A2(new_n361), .ZN(new_n456));
  OAI21_X1  g255(.A(new_n454), .B1(new_n455), .B2(new_n456), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n457), .A2(KEYINPUT85), .ZN(new_n458));
  INV_X1    g257(.A(KEYINPUT85), .ZN(new_n459));
  OAI211_X1 g258(.A(new_n459), .B(new_n454), .C1(new_n455), .C2(new_n456), .ZN(new_n460));
  NAND4_X1  g259(.A1(new_n453), .A2(new_n458), .A3(new_n274), .A4(new_n460), .ZN(new_n461));
  INV_X1    g260(.A(KEYINPUT37), .ZN(new_n462));
  NAND3_X1  g261(.A1(new_n254), .A2(new_n462), .A3(new_n263), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n463), .A2(new_n268), .ZN(new_n464));
  AOI21_X1  g263(.A(new_n462), .B1(new_n254), .B2(new_n263), .ZN(new_n465));
  OAI21_X1  g264(.A(KEYINPUT38), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  AOI21_X1  g265(.A(new_n253), .B1(new_n239), .B2(new_n241), .ZN(new_n467));
  NOR3_X1   g266(.A1(new_n260), .A2(new_n262), .A3(new_n259), .ZN(new_n468));
  OAI21_X1  g267(.A(KEYINPUT37), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  INV_X1    g268(.A(KEYINPUT38), .ZN(new_n470));
  NAND4_X1  g269(.A1(new_n469), .A2(new_n470), .A3(new_n268), .A4(new_n463), .ZN(new_n471));
  AND3_X1   g270(.A1(new_n466), .A2(new_n269), .A3(new_n471), .ZN(new_n472));
  NAND3_X1  g271(.A1(new_n367), .A2(new_n472), .A3(new_n368), .ZN(new_n473));
  NAND3_X1  g272(.A1(new_n461), .A2(new_n473), .A3(new_n440), .ZN(new_n474));
  INV_X1    g273(.A(new_n390), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n475), .A2(KEYINPUT36), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n432), .A2(new_n431), .ZN(new_n477));
  OAI21_X1  g276(.A(new_n476), .B1(new_n477), .B2(KEYINPUT36), .ZN(new_n478));
  NAND3_X1  g277(.A1(new_n442), .A2(new_n474), .A3(new_n478), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n436), .A2(new_n479), .ZN(new_n480));
  XNOR2_X1  g279(.A(G43gat), .B(G50gat), .ZN(new_n481));
  XNOR2_X1  g280(.A(new_n481), .B(KEYINPUT87), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n482), .A2(KEYINPUT15), .ZN(new_n483));
  OAI21_X1  g282(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n484));
  INV_X1    g283(.A(new_n484), .ZN(new_n485));
  NOR3_X1   g284(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n486));
  INV_X1    g285(.A(G29gat), .ZN(new_n487));
  INV_X1    g286(.A(G36gat), .ZN(new_n488));
  OAI22_X1  g287(.A1(new_n485), .A2(new_n486), .B1(new_n487), .B2(new_n488), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n483), .A2(new_n489), .ZN(new_n490));
  INV_X1    g289(.A(new_n490), .ZN(new_n491));
  OR2_X1    g290(.A1(new_n481), .A2(KEYINPUT15), .ZN(new_n492));
  AOI21_X1  g291(.A(new_n489), .B1(new_n483), .B2(new_n492), .ZN(new_n493));
  NOR2_X1   g292(.A1(new_n491), .A2(new_n493), .ZN(new_n494));
  XNOR2_X1  g293(.A(G15gat), .B(G22gat), .ZN(new_n495));
  INV_X1    g294(.A(G1gat), .ZN(new_n496));
  NAND3_X1  g295(.A1(new_n495), .A2(KEYINPUT16), .A3(new_n496), .ZN(new_n497));
  OAI221_X1 g296(.A(new_n497), .B1(KEYINPUT88), .B2(G8gat), .C1(new_n496), .C2(new_n495), .ZN(new_n498));
  NAND2_X1  g297(.A1(KEYINPUT88), .A2(G8gat), .ZN(new_n499));
  XNOR2_X1  g298(.A(new_n498), .B(new_n499), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n500), .A2(KEYINPUT89), .ZN(new_n501));
  INV_X1    g300(.A(new_n501), .ZN(new_n502));
  NOR2_X1   g301(.A1(new_n500), .A2(KEYINPUT89), .ZN(new_n503));
  OAI21_X1  g302(.A(new_n494), .B1(new_n502), .B2(new_n503), .ZN(new_n504));
  INV_X1    g303(.A(new_n493), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n505), .A2(new_n490), .ZN(new_n506));
  NAND2_X1  g305(.A1(new_n506), .A2(KEYINPUT17), .ZN(new_n507));
  XOR2_X1   g306(.A(new_n498), .B(new_n499), .Z(new_n508));
  INV_X1    g307(.A(KEYINPUT17), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n494), .A2(new_n509), .ZN(new_n510));
  NAND3_X1  g309(.A1(new_n507), .A2(new_n508), .A3(new_n510), .ZN(new_n511));
  NAND2_X1  g310(.A1(G229gat), .A2(G233gat), .ZN(new_n512));
  NAND3_X1  g311(.A1(new_n504), .A2(new_n511), .A3(new_n512), .ZN(new_n513));
  INV_X1    g312(.A(KEYINPUT18), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  INV_X1    g314(.A(new_n503), .ZN(new_n516));
  NAND3_X1  g315(.A1(new_n516), .A2(new_n506), .A3(new_n501), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n504), .A2(new_n517), .ZN(new_n518));
  XOR2_X1   g317(.A(new_n512), .B(KEYINPUT13), .Z(new_n519));
  NAND2_X1  g318(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  NAND4_X1  g319(.A1(new_n504), .A2(new_n511), .A3(KEYINPUT18), .A4(new_n512), .ZN(new_n521));
  NAND3_X1  g320(.A1(new_n515), .A2(new_n520), .A3(new_n521), .ZN(new_n522));
  XOR2_X1   g321(.A(KEYINPUT86), .B(KEYINPUT11), .Z(new_n523));
  XNOR2_X1  g322(.A(G113gat), .B(G141gat), .ZN(new_n524));
  XNOR2_X1  g323(.A(new_n523), .B(new_n524), .ZN(new_n525));
  XNOR2_X1  g324(.A(G169gat), .B(G197gat), .ZN(new_n526));
  XNOR2_X1  g325(.A(new_n525), .B(new_n526), .ZN(new_n527));
  XOR2_X1   g326(.A(new_n527), .B(KEYINPUT12), .Z(new_n528));
  NAND2_X1  g327(.A1(new_n522), .A2(new_n528), .ZN(new_n529));
  INV_X1    g328(.A(new_n528), .ZN(new_n530));
  NAND4_X1  g329(.A1(new_n515), .A2(new_n520), .A3(new_n521), .A4(new_n530), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n529), .A2(new_n531), .ZN(new_n532));
  AND3_X1   g331(.A1(new_n480), .A2(KEYINPUT90), .A3(new_n532), .ZN(new_n533));
  AOI21_X1  g332(.A(KEYINPUT90), .B1(new_n480), .B2(new_n532), .ZN(new_n534));
  OR2_X1    g333(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  INV_X1    g334(.A(KEYINPUT21), .ZN(new_n536));
  XNOR2_X1  g335(.A(G71gat), .B(G78gat), .ZN(new_n537));
  XNOR2_X1  g336(.A(new_n537), .B(KEYINPUT91), .ZN(new_n538));
  AOI21_X1  g337(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n539));
  XNOR2_X1  g338(.A(G57gat), .B(G64gat), .ZN(new_n540));
  OAI21_X1  g339(.A(new_n538), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  AOI21_X1  g340(.A(new_n539), .B1(new_n540), .B2(KEYINPUT92), .ZN(new_n542));
  OAI211_X1 g341(.A(new_n542), .B(new_n537), .C1(KEYINPUT92), .C2(new_n540), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n541), .A2(new_n543), .ZN(new_n544));
  OAI211_X1 g343(.A(new_n516), .B(new_n501), .C1(new_n536), .C2(new_n544), .ZN(new_n545));
  XOR2_X1   g344(.A(new_n545), .B(G183gat), .Z(new_n546));
  XNOR2_X1  g345(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  XNOR2_X1  g347(.A(new_n545), .B(G183gat), .ZN(new_n549));
  INV_X1    g348(.A(new_n547), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n544), .A2(new_n536), .ZN(new_n552));
  INV_X1    g351(.A(G211gat), .ZN(new_n553));
  XNOR2_X1  g352(.A(new_n552), .B(new_n553), .ZN(new_n554));
  INV_X1    g353(.A(new_n554), .ZN(new_n555));
  AND3_X1   g354(.A1(new_n548), .A2(new_n551), .A3(new_n555), .ZN(new_n556));
  AOI21_X1  g355(.A(new_n555), .B1(new_n548), .B2(new_n551), .ZN(new_n557));
  XNOR2_X1  g356(.A(G127gat), .B(G155gat), .ZN(new_n558));
  NAND2_X1  g357(.A1(G231gat), .A2(G233gat), .ZN(new_n559));
  XNOR2_X1  g358(.A(new_n558), .B(new_n559), .ZN(new_n560));
  INV_X1    g359(.A(new_n560), .ZN(new_n561));
  OR3_X1    g360(.A1(new_n556), .A2(new_n557), .A3(new_n561), .ZN(new_n562));
  OAI21_X1  g361(.A(new_n561), .B1(new_n556), .B2(new_n557), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  INV_X1    g363(.A(new_n564), .ZN(new_n565));
  XNOR2_X1  g364(.A(KEYINPUT93), .B(KEYINPUT94), .ZN(new_n566));
  NAND2_X1  g365(.A1(G85gat), .A2(G92gat), .ZN(new_n567));
  XNOR2_X1  g366(.A(new_n567), .B(KEYINPUT7), .ZN(new_n568));
  NAND2_X1  g367(.A1(G99gat), .A2(G106gat), .ZN(new_n569));
  INV_X1    g368(.A(G92gat), .ZN(new_n570));
  AOI22_X1  g369(.A1(KEYINPUT8), .A2(new_n569), .B1(new_n357), .B2(new_n570), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n568), .A2(new_n571), .ZN(new_n572));
  XNOR2_X1  g371(.A(G99gat), .B(G106gat), .ZN(new_n573));
  XNOR2_X1  g372(.A(new_n572), .B(new_n573), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n574), .A2(KEYINPUT95), .ZN(new_n575));
  INV_X1    g374(.A(KEYINPUT95), .ZN(new_n576));
  NAND4_X1  g375(.A1(new_n568), .A2(new_n576), .A3(new_n573), .A4(new_n571), .ZN(new_n577));
  NAND2_X1  g376(.A1(new_n575), .A2(new_n577), .ZN(new_n578));
  AND2_X1   g377(.A1(G232gat), .A2(G233gat), .ZN(new_n579));
  AOI22_X1  g378(.A1(new_n494), .A2(new_n578), .B1(KEYINPUT41), .B2(new_n579), .ZN(new_n580));
  NAND2_X1  g379(.A1(new_n507), .A2(new_n510), .ZN(new_n581));
  OAI21_X1  g380(.A(new_n580), .B1(new_n581), .B2(new_n578), .ZN(new_n582));
  XOR2_X1   g381(.A(G190gat), .B(G218gat), .Z(new_n583));
  INV_X1    g382(.A(new_n583), .ZN(new_n584));
  NOR2_X1   g383(.A1(new_n584), .A2(KEYINPUT96), .ZN(new_n585));
  INV_X1    g384(.A(new_n585), .ZN(new_n586));
  XNOR2_X1  g385(.A(G134gat), .B(G162gat), .ZN(new_n587));
  NAND3_X1  g386(.A1(new_n582), .A2(new_n586), .A3(new_n587), .ZN(new_n588));
  INV_X1    g387(.A(new_n588), .ZN(new_n589));
  AOI21_X1  g388(.A(new_n587), .B1(new_n582), .B2(new_n586), .ZN(new_n590));
  OAI21_X1  g389(.A(new_n566), .B1(new_n589), .B2(new_n590), .ZN(new_n591));
  INV_X1    g390(.A(new_n590), .ZN(new_n592));
  INV_X1    g391(.A(new_n566), .ZN(new_n593));
  NAND3_X1  g392(.A1(new_n592), .A2(new_n588), .A3(new_n593), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n584), .A2(KEYINPUT96), .ZN(new_n595));
  NOR2_X1   g394(.A1(new_n579), .A2(KEYINPUT41), .ZN(new_n596));
  XOR2_X1   g395(.A(new_n595), .B(new_n596), .Z(new_n597));
  AND3_X1   g396(.A1(new_n591), .A2(new_n594), .A3(new_n597), .ZN(new_n598));
  AOI21_X1  g397(.A(new_n597), .B1(new_n591), .B2(new_n594), .ZN(new_n599));
  NOR2_X1   g398(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  INV_X1    g399(.A(new_n600), .ZN(new_n601));
  XNOR2_X1  g400(.A(G120gat), .B(G148gat), .ZN(new_n602));
  XNOR2_X1  g401(.A(G176gat), .B(G204gat), .ZN(new_n603));
  XNOR2_X1  g402(.A(new_n602), .B(new_n603), .ZN(new_n604));
  INV_X1    g403(.A(new_n604), .ZN(new_n605));
  NAND2_X1  g404(.A1(G230gat), .A2(G233gat), .ZN(new_n606));
  AND2_X1   g405(.A1(new_n541), .A2(new_n543), .ZN(new_n607));
  AOI21_X1  g406(.A(new_n607), .B1(new_n577), .B2(new_n575), .ZN(new_n608));
  NOR2_X1   g407(.A1(new_n544), .A2(new_n574), .ZN(new_n609));
  OR2_X1    g408(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  INV_X1    g409(.A(KEYINPUT10), .ZN(new_n611));
  OAI21_X1  g410(.A(new_n611), .B1(new_n608), .B2(new_n609), .ZN(new_n612));
  NAND3_X1  g411(.A1(new_n578), .A2(KEYINPUT10), .A3(new_n607), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  AND2_X1   g413(.A1(new_n614), .A2(new_n606), .ZN(new_n615));
  NOR2_X1   g414(.A1(new_n615), .A2(KEYINPUT97), .ZN(new_n616));
  AND3_X1   g415(.A1(new_n614), .A2(KEYINPUT97), .A3(new_n606), .ZN(new_n617));
  OAI221_X1 g416(.A(new_n605), .B1(new_n606), .B2(new_n610), .C1(new_n616), .C2(new_n617), .ZN(new_n618));
  NOR2_X1   g417(.A1(new_n610), .A2(new_n606), .ZN(new_n619));
  OAI21_X1  g418(.A(new_n604), .B1(new_n615), .B2(new_n619), .ZN(new_n620));
  NAND2_X1  g419(.A1(new_n618), .A2(new_n620), .ZN(new_n621));
  NOR3_X1   g420(.A1(new_n565), .A2(new_n601), .A3(new_n621), .ZN(new_n622));
  NAND2_X1  g421(.A1(new_n535), .A2(new_n622), .ZN(new_n623));
  NOR2_X1   g422(.A1(new_n623), .A2(new_n437), .ZN(new_n624));
  XNOR2_X1  g423(.A(KEYINPUT98), .B(G1gat), .ZN(new_n625));
  XNOR2_X1  g424(.A(new_n624), .B(new_n625), .ZN(G1324gat));
  INV_X1    g425(.A(KEYINPUT99), .ZN(new_n627));
  INV_X1    g426(.A(new_n623), .ZN(new_n628));
  NAND2_X1  g427(.A1(new_n628), .A2(new_n274), .ZN(new_n629));
  XNOR2_X1  g428(.A(KEYINPUT16), .B(G8gat), .ZN(new_n630));
  OAI21_X1  g429(.A(new_n627), .B1(new_n629), .B2(new_n630), .ZN(new_n631));
  OR2_X1    g430(.A1(new_n631), .A2(KEYINPUT42), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n629), .A2(G8gat), .ZN(new_n633));
  NAND2_X1  g432(.A1(new_n631), .A2(KEYINPUT42), .ZN(new_n634));
  NAND3_X1  g433(.A1(new_n632), .A2(new_n633), .A3(new_n634), .ZN(G1325gat));
  INV_X1    g434(.A(G15gat), .ZN(new_n636));
  NOR3_X1   g435(.A1(new_n623), .A2(new_n636), .A3(new_n478), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n628), .A2(new_n477), .ZN(new_n638));
  AOI21_X1  g437(.A(new_n637), .B1(new_n636), .B2(new_n638), .ZN(G1326gat));
  NOR2_X1   g438(.A1(new_n623), .A2(new_n440), .ZN(new_n640));
  XNOR2_X1  g439(.A(new_n640), .B(KEYINPUT100), .ZN(new_n641));
  XNOR2_X1  g440(.A(KEYINPUT43), .B(G22gat), .ZN(new_n642));
  XNOR2_X1  g441(.A(new_n641), .B(new_n642), .ZN(G1327gat));
  INV_X1    g442(.A(new_n621), .ZN(new_n644));
  NAND3_X1  g443(.A1(new_n565), .A2(new_n601), .A3(new_n644), .ZN(new_n645));
  XNOR2_X1  g444(.A(new_n645), .B(KEYINPUT101), .ZN(new_n646));
  AND2_X1   g445(.A1(new_n535), .A2(new_n646), .ZN(new_n647));
  INV_X1    g446(.A(new_n437), .ZN(new_n648));
  NAND3_X1  g447(.A1(new_n647), .A2(new_n487), .A3(new_n648), .ZN(new_n649));
  XNOR2_X1  g448(.A(new_n649), .B(KEYINPUT45), .ZN(new_n650));
  INV_X1    g449(.A(KEYINPUT102), .ZN(new_n651));
  XNOR2_X1  g450(.A(new_n532), .B(new_n651), .ZN(new_n652));
  NOR3_X1   g451(.A1(new_n564), .A2(new_n621), .A3(new_n652), .ZN(new_n653));
  NAND3_X1  g452(.A1(new_n480), .A2(KEYINPUT44), .A3(new_n601), .ZN(new_n654));
  INV_X1    g453(.A(KEYINPUT104), .ZN(new_n655));
  AND3_X1   g454(.A1(new_n433), .A2(new_n369), .A3(new_n434), .ZN(new_n656));
  AOI21_X1  g455(.A(new_n434), .B1(new_n369), .B2(new_n427), .ZN(new_n657));
  OAI21_X1  g456(.A(new_n655), .B1(new_n656), .B2(new_n657), .ZN(new_n658));
  NAND3_X1  g457(.A1(new_n429), .A2(KEYINPUT104), .A3(new_n435), .ZN(new_n659));
  AND2_X1   g458(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  NAND2_X1  g459(.A1(new_n479), .A2(KEYINPUT103), .ZN(new_n661));
  INV_X1    g460(.A(KEYINPUT103), .ZN(new_n662));
  NAND4_X1  g461(.A1(new_n442), .A2(new_n474), .A3(new_n662), .A4(new_n478), .ZN(new_n663));
  NAND2_X1  g462(.A1(new_n661), .A2(new_n663), .ZN(new_n664));
  AOI21_X1  g463(.A(new_n600), .B1(new_n660), .B2(new_n664), .ZN(new_n665));
  OAI211_X1 g464(.A(new_n653), .B(new_n654), .C1(new_n665), .C2(KEYINPUT44), .ZN(new_n666));
  OAI21_X1  g465(.A(G29gat), .B1(new_n666), .B2(new_n437), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n650), .A2(new_n667), .ZN(G1328gat));
  NAND3_X1  g467(.A1(new_n647), .A2(new_n488), .A3(new_n274), .ZN(new_n669));
  AND2_X1   g468(.A1(KEYINPUT105), .A2(KEYINPUT46), .ZN(new_n670));
  OR2_X1    g469(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  NOR2_X1   g470(.A1(KEYINPUT105), .A2(KEYINPUT46), .ZN(new_n672));
  OAI21_X1  g471(.A(new_n669), .B1(new_n670), .B2(new_n672), .ZN(new_n673));
  INV_X1    g472(.A(new_n654), .ZN(new_n674));
  AND2_X1   g473(.A1(new_n661), .A2(new_n663), .ZN(new_n675));
  NAND2_X1  g474(.A1(new_n658), .A2(new_n659), .ZN(new_n676));
  OAI21_X1  g475(.A(new_n601), .B1(new_n675), .B2(new_n676), .ZN(new_n677));
  INV_X1    g476(.A(KEYINPUT44), .ZN(new_n678));
  AOI21_X1  g477(.A(new_n674), .B1(new_n677), .B2(new_n678), .ZN(new_n679));
  NAND4_X1  g478(.A1(new_n679), .A2(KEYINPUT106), .A3(new_n274), .A4(new_n653), .ZN(new_n680));
  INV_X1    g479(.A(KEYINPUT106), .ZN(new_n681));
  OAI21_X1  g480(.A(new_n681), .B1(new_n666), .B2(new_n438), .ZN(new_n682));
  NAND3_X1  g481(.A1(new_n680), .A2(new_n682), .A3(G36gat), .ZN(new_n683));
  NAND3_X1  g482(.A1(new_n671), .A2(new_n673), .A3(new_n683), .ZN(new_n684));
  NAND2_X1  g483(.A1(new_n684), .A2(KEYINPUT107), .ZN(new_n685));
  INV_X1    g484(.A(KEYINPUT107), .ZN(new_n686));
  NAND4_X1  g485(.A1(new_n671), .A2(new_n686), .A3(new_n673), .A4(new_n683), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n685), .A2(new_n687), .ZN(G1329gat));
  OR3_X1    g487(.A1(new_n666), .A2(KEYINPUT109), .A3(new_n478), .ZN(new_n689));
  OAI21_X1  g488(.A(KEYINPUT109), .B1(new_n666), .B2(new_n478), .ZN(new_n690));
  NAND3_X1  g489(.A1(new_n689), .A2(G43gat), .A3(new_n690), .ZN(new_n691));
  INV_X1    g490(.A(G43gat), .ZN(new_n692));
  NAND3_X1  g491(.A1(new_n647), .A2(new_n692), .A3(new_n477), .ZN(new_n693));
  NAND3_X1  g492(.A1(new_n691), .A2(KEYINPUT47), .A3(new_n693), .ZN(new_n694));
  OAI21_X1  g493(.A(G43gat), .B1(new_n666), .B2(new_n478), .ZN(new_n695));
  OR2_X1    g494(.A1(new_n695), .A2(KEYINPUT108), .ZN(new_n696));
  NAND2_X1  g495(.A1(new_n695), .A2(KEYINPUT108), .ZN(new_n697));
  AND3_X1   g496(.A1(new_n696), .A2(new_n693), .A3(new_n697), .ZN(new_n698));
  OAI21_X1  g497(.A(new_n694), .B1(new_n698), .B2(KEYINPUT47), .ZN(G1330gat));
  INV_X1    g498(.A(KEYINPUT48), .ZN(new_n700));
  INV_X1    g499(.A(KEYINPUT110), .ZN(new_n701));
  NAND4_X1  g500(.A1(new_n679), .A2(new_n701), .A3(new_n441), .A4(new_n653), .ZN(new_n702));
  OAI21_X1  g501(.A(KEYINPUT110), .B1(new_n666), .B2(new_n440), .ZN(new_n703));
  NAND3_X1  g502(.A1(new_n702), .A2(new_n703), .A3(G50gat), .ZN(new_n704));
  INV_X1    g503(.A(G50gat), .ZN(new_n705));
  NAND3_X1  g504(.A1(new_n647), .A2(new_n705), .A3(new_n441), .ZN(new_n706));
  AOI21_X1  g505(.A(new_n700), .B1(new_n704), .B2(new_n706), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n677), .A2(new_n678), .ZN(new_n708));
  NAND4_X1  g507(.A1(new_n708), .A2(new_n441), .A3(new_n653), .A4(new_n654), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n709), .A2(G50gat), .ZN(new_n710));
  AND3_X1   g509(.A1(new_n706), .A2(new_n700), .A3(new_n710), .ZN(new_n711));
  OAI21_X1  g510(.A(KEYINPUT111), .B1(new_n707), .B2(new_n711), .ZN(new_n712));
  INV_X1    g511(.A(KEYINPUT111), .ZN(new_n713));
  NAND3_X1  g512(.A1(new_n706), .A2(new_n710), .A3(new_n700), .ZN(new_n714));
  AND4_X1   g513(.A1(new_n705), .A2(new_n535), .A3(new_n646), .A4(new_n441), .ZN(new_n715));
  AOI21_X1  g514(.A(new_n705), .B1(new_n709), .B2(KEYINPUT110), .ZN(new_n716));
  AOI21_X1  g515(.A(new_n715), .B1(new_n716), .B2(new_n702), .ZN(new_n717));
  OAI211_X1 g516(.A(new_n713), .B(new_n714), .C1(new_n717), .C2(new_n700), .ZN(new_n718));
  AND2_X1   g517(.A1(new_n712), .A2(new_n718), .ZN(G1331gat));
  AOI211_X1 g518(.A(new_n565), .B(new_n601), .C1(new_n660), .C2(new_n664), .ZN(new_n720));
  NOR2_X1   g519(.A1(new_n532), .A2(new_n651), .ZN(new_n721));
  AOI21_X1  g520(.A(KEYINPUT102), .B1(new_n529), .B2(new_n531), .ZN(new_n722));
  NOR2_X1   g521(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  NOR2_X1   g522(.A1(new_n723), .A2(new_n644), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n720), .A2(new_n724), .ZN(new_n725));
  NOR2_X1   g524(.A1(new_n725), .A2(new_n437), .ZN(new_n726));
  XNOR2_X1  g525(.A(KEYINPUT112), .B(G57gat), .ZN(new_n727));
  XNOR2_X1  g526(.A(new_n726), .B(new_n727), .ZN(G1332gat));
  INV_X1    g527(.A(new_n725), .ZN(new_n729));
  INV_X1    g528(.A(KEYINPUT49), .ZN(new_n730));
  INV_X1    g529(.A(G64gat), .ZN(new_n731));
  OAI21_X1  g530(.A(new_n274), .B1(new_n730), .B2(new_n731), .ZN(new_n732));
  XNOR2_X1  g531(.A(new_n732), .B(KEYINPUT113), .ZN(new_n733));
  NAND2_X1  g532(.A1(new_n729), .A2(new_n733), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n730), .A2(new_n731), .ZN(new_n735));
  XNOR2_X1  g534(.A(new_n734), .B(new_n735), .ZN(G1333gat));
  OAI21_X1  g535(.A(G71gat), .B1(new_n725), .B2(new_n478), .ZN(new_n737));
  XNOR2_X1  g536(.A(new_n477), .B(KEYINPUT114), .ZN(new_n738));
  INV_X1    g537(.A(G71gat), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  OAI21_X1  g539(.A(new_n737), .B1(new_n725), .B2(new_n740), .ZN(new_n741));
  XOR2_X1   g540(.A(new_n741), .B(KEYINPUT50), .Z(G1334gat));
  NOR2_X1   g541(.A1(new_n725), .A2(new_n440), .ZN(new_n743));
  XOR2_X1   g542(.A(KEYINPUT115), .B(G78gat), .Z(new_n744));
  XNOR2_X1  g543(.A(new_n743), .B(new_n744), .ZN(G1335gat));
  NOR2_X1   g544(.A1(new_n564), .A2(new_n723), .ZN(new_n746));
  NAND3_X1  g545(.A1(new_n679), .A2(new_n621), .A3(new_n746), .ZN(new_n747));
  NOR3_X1   g546(.A1(new_n747), .A2(new_n357), .A3(new_n437), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n665), .A2(new_n746), .ZN(new_n749));
  INV_X1    g548(.A(KEYINPUT51), .ZN(new_n750));
  XNOR2_X1  g549(.A(new_n749), .B(new_n750), .ZN(new_n751));
  NAND3_X1  g550(.A1(new_n751), .A2(new_n648), .A3(new_n621), .ZN(new_n752));
  AOI21_X1  g551(.A(new_n748), .B1(new_n752), .B2(new_n357), .ZN(G1336gat));
  OAI21_X1  g552(.A(G92gat), .B1(new_n747), .B2(new_n438), .ZN(new_n754));
  INV_X1    g553(.A(KEYINPUT52), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n751), .A2(new_n621), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n274), .A2(new_n570), .ZN(new_n757));
  OAI211_X1 g556(.A(new_n754), .B(new_n755), .C1(new_n756), .C2(new_n757), .ZN(new_n758));
  INV_X1    g557(.A(KEYINPUT116), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n754), .A2(new_n759), .ZN(new_n760));
  INV_X1    g559(.A(KEYINPUT117), .ZN(new_n761));
  OAI21_X1  g560(.A(KEYINPUT118), .B1(new_n749), .B2(new_n761), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n762), .A2(new_n750), .ZN(new_n763));
  INV_X1    g562(.A(KEYINPUT118), .ZN(new_n764));
  OAI21_X1  g563(.A(KEYINPUT117), .B1(new_n764), .B2(new_n750), .ZN(new_n765));
  NAND2_X1  g564(.A1(new_n749), .A2(new_n765), .ZN(new_n766));
  NOR2_X1   g565(.A1(new_n644), .A2(new_n757), .ZN(new_n767));
  NAND3_X1  g566(.A1(new_n763), .A2(new_n766), .A3(new_n767), .ZN(new_n768));
  OAI211_X1 g567(.A(KEYINPUT116), .B(G92gat), .C1(new_n747), .C2(new_n438), .ZN(new_n769));
  AND3_X1   g568(.A1(new_n760), .A2(new_n768), .A3(new_n769), .ZN(new_n770));
  OAI21_X1  g569(.A(new_n758), .B1(new_n770), .B2(new_n755), .ZN(G1337gat));
  OAI21_X1  g570(.A(G99gat), .B1(new_n747), .B2(new_n478), .ZN(new_n772));
  INV_X1    g571(.A(G99gat), .ZN(new_n773));
  NAND2_X1  g572(.A1(new_n477), .A2(new_n773), .ZN(new_n774));
  OAI21_X1  g573(.A(new_n772), .B1(new_n756), .B2(new_n774), .ZN(G1338gat));
  NOR3_X1   g574(.A1(new_n644), .A2(G106gat), .A3(new_n440), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n751), .A2(new_n776), .ZN(new_n777));
  OAI21_X1  g576(.A(G106gat), .B1(new_n747), .B2(new_n440), .ZN(new_n778));
  INV_X1    g577(.A(KEYINPUT53), .ZN(new_n779));
  NAND3_X1  g578(.A1(new_n777), .A2(new_n778), .A3(new_n779), .ZN(new_n780));
  NAND3_X1  g579(.A1(new_n763), .A2(new_n766), .A3(new_n776), .ZN(new_n781));
  AND2_X1   g580(.A1(new_n781), .A2(new_n778), .ZN(new_n782));
  OAI21_X1  g581(.A(new_n780), .B1(new_n782), .B2(new_n779), .ZN(G1339gat));
  NAND4_X1  g582(.A1(new_n564), .A2(new_n600), .A3(new_n644), .A4(new_n652), .ZN(new_n784));
  NOR3_X1   g583(.A1(new_n614), .A2(KEYINPUT119), .A3(new_n606), .ZN(new_n785));
  INV_X1    g584(.A(KEYINPUT54), .ZN(new_n786));
  NOR2_X1   g585(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  OAI21_X1  g586(.A(KEYINPUT119), .B1(new_n614), .B2(new_n606), .ZN(new_n788));
  OAI211_X1 g587(.A(new_n787), .B(new_n788), .C1(new_n616), .C2(new_n617), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n615), .A2(new_n786), .ZN(new_n790));
  NAND3_X1  g589(.A1(new_n789), .A2(new_n604), .A3(new_n790), .ZN(new_n791));
  INV_X1    g590(.A(KEYINPUT55), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n791), .A2(new_n792), .ZN(new_n793));
  NAND4_X1  g592(.A1(new_n789), .A2(KEYINPUT55), .A3(new_n604), .A4(new_n790), .ZN(new_n794));
  NOR2_X1   g593(.A1(new_n518), .A2(new_n519), .ZN(new_n795));
  AOI21_X1  g594(.A(new_n512), .B1(new_n504), .B2(new_n511), .ZN(new_n796));
  OAI21_X1  g595(.A(new_n527), .B1(new_n795), .B2(new_n796), .ZN(new_n797));
  AND2_X1   g596(.A1(new_n797), .A2(new_n531), .ZN(new_n798));
  NAND4_X1  g597(.A1(new_n793), .A2(new_n618), .A3(new_n794), .A4(new_n798), .ZN(new_n799));
  NOR2_X1   g598(.A1(new_n799), .A2(new_n600), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n621), .A2(new_n798), .ZN(new_n801));
  NAND3_X1  g600(.A1(new_n793), .A2(new_n618), .A3(new_n794), .ZN(new_n802));
  OAI21_X1  g601(.A(new_n801), .B1(new_n802), .B2(new_n652), .ZN(new_n803));
  AOI21_X1  g602(.A(new_n800), .B1(new_n600), .B2(new_n803), .ZN(new_n804));
  OAI21_X1  g603(.A(new_n784), .B1(new_n804), .B2(new_n564), .ZN(new_n805));
  NOR2_X1   g604(.A1(new_n437), .A2(new_n274), .ZN(new_n806));
  AND3_X1   g605(.A1(new_n805), .A2(new_n433), .A3(new_n806), .ZN(new_n807));
  INV_X1    g606(.A(new_n807), .ZN(new_n808));
  INV_X1    g607(.A(new_n532), .ZN(new_n809));
  OAI21_X1  g608(.A(G113gat), .B1(new_n808), .B2(new_n809), .ZN(new_n810));
  AND3_X1   g609(.A1(new_n805), .A2(new_n427), .A3(new_n806), .ZN(new_n811));
  NAND3_X1  g610(.A1(new_n811), .A2(new_n277), .A3(new_n723), .ZN(new_n812));
  NAND2_X1  g611(.A1(new_n810), .A2(new_n812), .ZN(G1340gat));
  OAI21_X1  g612(.A(G120gat), .B1(new_n808), .B2(new_n644), .ZN(new_n814));
  NAND3_X1  g613(.A1(new_n811), .A2(new_n279), .A3(new_n621), .ZN(new_n815));
  NAND2_X1  g614(.A1(new_n814), .A2(new_n815), .ZN(G1341gat));
  NAND3_X1  g615(.A1(new_n807), .A2(G127gat), .A3(new_n564), .ZN(new_n817));
  AND2_X1   g616(.A1(new_n811), .A2(new_n564), .ZN(new_n818));
  OAI21_X1  g617(.A(new_n817), .B1(new_n818), .B2(G127gat), .ZN(new_n819));
  XNOR2_X1  g618(.A(new_n819), .B(KEYINPUT120), .ZN(G1342gat));
  NAND3_X1  g619(.A1(new_n811), .A2(new_n283), .A3(new_n601), .ZN(new_n821));
  XOR2_X1   g620(.A(new_n821), .B(KEYINPUT56), .Z(new_n822));
  OAI21_X1  g621(.A(G134gat), .B1(new_n808), .B2(new_n600), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n822), .A2(new_n823), .ZN(G1343gat));
  NAND4_X1  g623(.A1(new_n723), .A2(new_n618), .A3(new_n793), .A4(new_n794), .ZN(new_n825));
  AOI21_X1  g624(.A(new_n601), .B1(new_n825), .B2(new_n801), .ZN(new_n826));
  OAI21_X1  g625(.A(new_n565), .B1(new_n826), .B2(new_n800), .ZN(new_n827));
  AOI21_X1  g626(.A(new_n440), .B1(new_n827), .B2(new_n784), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n478), .A2(new_n806), .ZN(new_n829));
  INV_X1    g628(.A(new_n829), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n828), .A2(new_n830), .ZN(new_n831));
  NOR3_X1   g630(.A1(new_n831), .A2(G141gat), .A3(new_n809), .ZN(new_n832));
  INV_X1    g631(.A(KEYINPUT122), .ZN(new_n833));
  AOI21_X1  g632(.A(new_n832), .B1(new_n833), .B2(KEYINPUT58), .ZN(new_n834));
  NAND4_X1  g633(.A1(new_n793), .A2(new_n532), .A3(new_n618), .A4(new_n794), .ZN(new_n835));
  AOI21_X1  g634(.A(new_n601), .B1(new_n835), .B2(new_n801), .ZN(new_n836));
  OAI21_X1  g635(.A(new_n565), .B1(new_n836), .B2(new_n800), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n837), .A2(new_n784), .ZN(new_n838));
  NAND3_X1  g637(.A1(new_n838), .A2(KEYINPUT57), .A3(new_n441), .ZN(new_n839));
  OAI21_X1  g638(.A(new_n839), .B1(new_n828), .B2(KEYINPUT57), .ZN(new_n840));
  NAND3_X1  g639(.A1(new_n840), .A2(new_n532), .A3(new_n830), .ZN(new_n841));
  INV_X1    g640(.A(KEYINPUT58), .ZN(new_n842));
  NOR2_X1   g641(.A1(new_n316), .A2(new_n317), .ZN(new_n843));
  NAND3_X1  g642(.A1(new_n841), .A2(new_n842), .A3(new_n843), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n834), .A2(new_n844), .ZN(new_n845));
  INV_X1    g644(.A(KEYINPUT121), .ZN(new_n846));
  AOI21_X1  g645(.A(KEYINPUT57), .B1(new_n805), .B2(new_n441), .ZN(new_n847));
  INV_X1    g646(.A(KEYINPUT57), .ZN(new_n848));
  AOI211_X1 g647(.A(new_n848), .B(new_n440), .C1(new_n837), .C2(new_n784), .ZN(new_n849));
  OAI211_X1 g648(.A(new_n846), .B(new_n830), .C1(new_n847), .C2(new_n849), .ZN(new_n850));
  INV_X1    g649(.A(new_n850), .ZN(new_n851));
  AOI21_X1  g650(.A(new_n846), .B1(new_n840), .B2(new_n830), .ZN(new_n852));
  OAI21_X1  g651(.A(new_n723), .B1(new_n851), .B2(new_n852), .ZN(new_n853));
  AOI22_X1  g652(.A1(new_n853), .A2(new_n843), .B1(new_n833), .B2(new_n832), .ZN(new_n854));
  OAI21_X1  g653(.A(new_n845), .B1(new_n854), .B2(new_n842), .ZN(G1344gat));
  INV_X1    g654(.A(KEYINPUT59), .ZN(new_n856));
  OAI211_X1 g655(.A(new_n856), .B(new_n621), .C1(new_n851), .C2(new_n852), .ZN(new_n857));
  OAI21_X1  g656(.A(KEYINPUT59), .B1(new_n831), .B2(new_n644), .ZN(new_n858));
  NAND2_X1  g657(.A1(new_n858), .A2(new_n289), .ZN(new_n859));
  INV_X1    g658(.A(new_n828), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n860), .A2(KEYINPUT57), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n622), .A2(new_n809), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n862), .A2(new_n837), .ZN(new_n863));
  NAND3_X1  g662(.A1(new_n863), .A2(new_n848), .A3(new_n441), .ZN(new_n864));
  NAND3_X1  g663(.A1(new_n861), .A2(new_n621), .A3(new_n864), .ZN(new_n865));
  OAI211_X1 g664(.A(KEYINPUT59), .B(G148gat), .C1(new_n865), .C2(new_n829), .ZN(new_n866));
  NAND3_X1  g665(.A1(new_n857), .A2(new_n859), .A3(new_n866), .ZN(new_n867));
  INV_X1    g666(.A(KEYINPUT123), .ZN(new_n868));
  NAND2_X1  g667(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  NAND4_X1  g668(.A1(new_n857), .A2(new_n866), .A3(KEYINPUT123), .A4(new_n859), .ZN(new_n870));
  NAND2_X1  g669(.A1(new_n869), .A2(new_n870), .ZN(G1345gat));
  OAI21_X1  g670(.A(new_n564), .B1(new_n851), .B2(new_n852), .ZN(new_n872));
  NOR2_X1   g671(.A1(new_n831), .A2(new_n565), .ZN(new_n873));
  MUX2_X1   g672(.A(new_n872), .B(new_n873), .S(new_n310), .Z(G1346gat));
  NAND4_X1  g673(.A1(new_n828), .A2(new_n314), .A3(new_n601), .A4(new_n830), .ZN(new_n875));
  OAI21_X1  g674(.A(new_n601), .B1(new_n851), .B2(new_n852), .ZN(new_n876));
  NAND2_X1  g675(.A1(new_n876), .A2(KEYINPUT124), .ZN(new_n877));
  INV_X1    g676(.A(KEYINPUT124), .ZN(new_n878));
  OAI211_X1 g677(.A(new_n878), .B(new_n601), .C1(new_n851), .C2(new_n852), .ZN(new_n879));
  NAND2_X1  g678(.A1(new_n877), .A2(new_n879), .ZN(new_n880));
  OAI21_X1  g679(.A(new_n875), .B1(new_n880), .B2(new_n314), .ZN(G1347gat));
  AND4_X1   g680(.A1(new_n437), .A2(new_n805), .A3(new_n274), .A4(new_n440), .ZN(new_n882));
  AND2_X1   g681(.A1(new_n882), .A2(new_n475), .ZN(new_n883));
  NAND3_X1  g682(.A1(new_n883), .A2(new_n218), .A3(new_n723), .ZN(new_n884));
  NAND2_X1  g683(.A1(new_n882), .A2(new_n738), .ZN(new_n885));
  OAI21_X1  g684(.A(G169gat), .B1(new_n885), .B2(new_n809), .ZN(new_n886));
  NAND2_X1  g685(.A1(new_n884), .A2(new_n886), .ZN(G1348gat));
  AOI21_X1  g686(.A(G176gat), .B1(new_n883), .B2(new_n621), .ZN(new_n888));
  NOR3_X1   g687(.A1(new_n885), .A2(new_n219), .A3(new_n644), .ZN(new_n889));
  NOR2_X1   g688(.A1(new_n888), .A2(new_n889), .ZN(G1349gat));
  NAND3_X1  g689(.A1(new_n883), .A2(new_n202), .A3(new_n564), .ZN(new_n891));
  OAI21_X1  g690(.A(G183gat), .B1(new_n885), .B2(new_n565), .ZN(new_n892));
  NAND2_X1  g691(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  XNOR2_X1  g692(.A(new_n893), .B(KEYINPUT60), .ZN(G1350gat));
  NAND3_X1  g693(.A1(new_n883), .A2(new_n203), .A3(new_n601), .ZN(new_n895));
  NAND3_X1  g694(.A1(new_n882), .A2(new_n601), .A3(new_n738), .ZN(new_n896));
  INV_X1    g695(.A(KEYINPUT61), .ZN(new_n897));
  NAND3_X1  g696(.A1(new_n896), .A2(new_n897), .A3(G190gat), .ZN(new_n898));
  INV_X1    g697(.A(new_n898), .ZN(new_n899));
  AOI21_X1  g698(.A(new_n897), .B1(new_n896), .B2(G190gat), .ZN(new_n900));
  OAI21_X1  g699(.A(new_n895), .B1(new_n899), .B2(new_n900), .ZN(G1351gat));
  NAND3_X1  g700(.A1(new_n478), .A2(new_n437), .A3(new_n274), .ZN(new_n902));
  NOR2_X1   g701(.A1(new_n860), .A2(new_n902), .ZN(new_n903));
  INV_X1    g702(.A(G197gat), .ZN(new_n904));
  NAND3_X1  g703(.A1(new_n903), .A2(new_n904), .A3(new_n723), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n861), .A2(new_n864), .ZN(new_n906));
  XOR2_X1   g705(.A(new_n902), .B(KEYINPUT125), .Z(new_n907));
  XNOR2_X1  g706(.A(new_n907), .B(KEYINPUT126), .ZN(new_n908));
  NOR3_X1   g707(.A1(new_n906), .A2(new_n809), .A3(new_n908), .ZN(new_n909));
  OAI21_X1  g708(.A(new_n905), .B1(new_n909), .B2(new_n904), .ZN(G1352gat));
  INV_X1    g709(.A(G204gat), .ZN(new_n911));
  NAND3_X1  g710(.A1(new_n903), .A2(new_n911), .A3(new_n621), .ZN(new_n912));
  XOR2_X1   g711(.A(new_n912), .B(KEYINPUT62), .Z(new_n913));
  NOR3_X1   g712(.A1(new_n906), .A2(new_n644), .A3(new_n908), .ZN(new_n914));
  OAI21_X1  g713(.A(new_n913), .B1(new_n914), .B2(new_n911), .ZN(G1353gat));
  NAND3_X1  g714(.A1(new_n861), .A2(new_n564), .A3(new_n864), .ZN(new_n916));
  OAI21_X1  g715(.A(G211gat), .B1(new_n916), .B2(new_n907), .ZN(new_n917));
  OR2_X1    g716(.A1(new_n917), .A2(KEYINPUT63), .ZN(new_n918));
  NAND2_X1  g717(.A1(new_n917), .A2(KEYINPUT63), .ZN(new_n919));
  NAND3_X1  g718(.A1(new_n903), .A2(new_n553), .A3(new_n564), .ZN(new_n920));
  XNOR2_X1  g719(.A(new_n920), .B(KEYINPUT127), .ZN(new_n921));
  NAND3_X1  g720(.A1(new_n918), .A2(new_n919), .A3(new_n921), .ZN(G1354gat));
  AOI21_X1  g721(.A(G218gat), .B1(new_n903), .B2(new_n601), .ZN(new_n923));
  NOR3_X1   g722(.A1(new_n906), .A2(new_n600), .A3(new_n908), .ZN(new_n924));
  AOI21_X1  g723(.A(new_n923), .B1(new_n924), .B2(G218gat), .ZN(G1355gat));
endmodule


