//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 0 1 1 1 0 1 0 1 0 1 1 0 1 1 1 1 1 0 1 0 1 0 1 0 0 0 1 1 1 1 0 1 0 1 1 0 1 0 0 1 0 0 0 1 1 1 1 1 1 1 0 1 1 0 0 0 1 1 0 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:19:24 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n712, new_n713, new_n714,
    new_n715, new_n717, new_n718, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n754, new_n755, new_n756, new_n757, new_n758, new_n759,
    new_n760, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n772, new_n773, new_n774, new_n775,
    new_n776, new_n777, new_n778, new_n779, new_n780, new_n782, new_n783,
    new_n784, new_n785, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n793, new_n794, new_n795, new_n797, new_n798, new_n800, new_n801,
    new_n802, new_n803, new_n804, new_n805, new_n806, new_n807, new_n808,
    new_n809, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n821, new_n822, new_n823, new_n824,
    new_n825, new_n826, new_n827, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n866, new_n867, new_n869, new_n870,
    new_n872, new_n873, new_n874, new_n875, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n920, new_n921, new_n923, new_n924,
    new_n925, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n937, new_n938, new_n940, new_n941,
    new_n942, new_n944, new_n945, new_n946, new_n947, new_n949, new_n950,
    new_n951, new_n952, new_n953, new_n954, new_n955, new_n956, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n968, new_n969, new_n970, new_n971, new_n973, new_n974;
  XNOR2_X1  g000(.A(G15gat), .B(G43gat), .ZN(new_n202));
  XNOR2_X1  g001(.A(G71gat), .B(G99gat), .ZN(new_n203));
  XNOR2_X1  g002(.A(new_n202), .B(new_n203), .ZN(new_n204));
  INV_X1    g003(.A(KEYINPUT71), .ZN(new_n205));
  INV_X1    g004(.A(G113gat), .ZN(new_n206));
  NAND2_X1  g005(.A1(new_n206), .A2(KEYINPUT70), .ZN(new_n207));
  INV_X1    g006(.A(KEYINPUT70), .ZN(new_n208));
  NAND2_X1  g007(.A1(new_n208), .A2(G113gat), .ZN(new_n209));
  NAND3_X1  g008(.A1(new_n207), .A2(new_n209), .A3(G120gat), .ZN(new_n210));
  NOR2_X1   g009(.A1(new_n206), .A2(G120gat), .ZN(new_n211));
  INV_X1    g010(.A(new_n211), .ZN(new_n212));
  AOI21_X1  g011(.A(new_n205), .B1(new_n210), .B2(new_n212), .ZN(new_n213));
  INV_X1    g012(.A(new_n213), .ZN(new_n214));
  NAND3_X1  g013(.A1(new_n210), .A2(new_n205), .A3(new_n212), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n214), .A2(new_n215), .ZN(new_n216));
  INV_X1    g015(.A(G127gat), .ZN(new_n217));
  NAND2_X1  g016(.A1(new_n217), .A2(G134gat), .ZN(new_n218));
  INV_X1    g017(.A(G134gat), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n219), .A2(G127gat), .ZN(new_n220));
  INV_X1    g019(.A(KEYINPUT1), .ZN(new_n221));
  AND3_X1   g020(.A1(new_n218), .A2(new_n220), .A3(new_n221), .ZN(new_n222));
  INV_X1    g021(.A(G120gat), .ZN(new_n223));
  NOR2_X1   g022(.A1(new_n223), .A2(G113gat), .ZN(new_n224));
  OAI21_X1  g023(.A(new_n221), .B1(new_n211), .B2(new_n224), .ZN(new_n225));
  INV_X1    g024(.A(KEYINPUT69), .ZN(new_n226));
  NAND3_X1  g025(.A1(new_n218), .A2(new_n220), .A3(KEYINPUT68), .ZN(new_n227));
  OR3_X1    g026(.A1(new_n219), .A2(KEYINPUT68), .A3(G127gat), .ZN(new_n228));
  NAND4_X1  g027(.A1(new_n225), .A2(new_n226), .A3(new_n227), .A4(new_n228), .ZN(new_n229));
  XNOR2_X1  g028(.A(G113gat), .B(G120gat), .ZN(new_n230));
  OAI21_X1  g029(.A(new_n228), .B1(new_n230), .B2(KEYINPUT1), .ZN(new_n231));
  INV_X1    g030(.A(new_n227), .ZN(new_n232));
  OAI21_X1  g031(.A(KEYINPUT69), .B1(new_n231), .B2(new_n232), .ZN(new_n233));
  AOI22_X1  g032(.A1(new_n216), .A2(new_n222), .B1(new_n229), .B2(new_n233), .ZN(new_n234));
  OAI21_X1  g033(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n235));
  NAND2_X1  g034(.A1(G183gat), .A2(G190gat), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n235), .A2(new_n236), .ZN(new_n237));
  INV_X1    g036(.A(new_n237), .ZN(new_n238));
  NAND3_X1  g037(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n239));
  INV_X1    g038(.A(new_n239), .ZN(new_n240));
  NOR2_X1   g039(.A1(new_n238), .A2(new_n240), .ZN(new_n241));
  INV_X1    g040(.A(KEYINPUT23), .ZN(new_n242));
  INV_X1    g041(.A(G169gat), .ZN(new_n243));
  INV_X1    g042(.A(G176gat), .ZN(new_n244));
  NAND3_X1  g043(.A1(new_n242), .A2(new_n243), .A3(new_n244), .ZN(new_n245));
  OAI21_X1  g044(.A(KEYINPUT23), .B1(G169gat), .B2(G176gat), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n245), .A2(new_n246), .ZN(new_n247));
  NAND2_X1  g046(.A1(G169gat), .A2(G176gat), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n248), .A2(KEYINPUT67), .ZN(new_n249));
  INV_X1    g048(.A(KEYINPUT67), .ZN(new_n250));
  NAND3_X1  g049(.A1(new_n250), .A2(G169gat), .A3(G176gat), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n249), .A2(new_n251), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n247), .A2(new_n252), .ZN(new_n253));
  INV_X1    g052(.A(KEYINPUT25), .ZN(new_n254));
  NOR3_X1   g053(.A1(new_n241), .A2(new_n253), .A3(new_n254), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n239), .A2(KEYINPUT65), .ZN(new_n256));
  INV_X1    g055(.A(KEYINPUT65), .ZN(new_n257));
  NAND4_X1  g056(.A1(new_n257), .A2(KEYINPUT24), .A3(G183gat), .A4(G190gat), .ZN(new_n258));
  NAND2_X1  g057(.A1(new_n256), .A2(new_n258), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n259), .A2(new_n237), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n260), .A2(KEYINPUT66), .ZN(new_n261));
  AOI22_X1  g060(.A1(new_n256), .A2(new_n258), .B1(new_n236), .B2(new_n235), .ZN(new_n262));
  INV_X1    g061(.A(KEYINPUT66), .ZN(new_n263));
  NAND2_X1  g062(.A1(new_n262), .A2(new_n263), .ZN(new_n264));
  AOI22_X1  g063(.A1(new_n246), .A2(new_n245), .B1(new_n249), .B2(new_n251), .ZN(new_n265));
  NAND3_X1  g064(.A1(new_n261), .A2(new_n264), .A3(new_n265), .ZN(new_n266));
  AOI21_X1  g065(.A(new_n255), .B1(new_n266), .B2(new_n254), .ZN(new_n267));
  XNOR2_X1  g066(.A(KEYINPUT27), .B(G183gat), .ZN(new_n268));
  INV_X1    g067(.A(G190gat), .ZN(new_n269));
  AOI21_X1  g068(.A(KEYINPUT28), .B1(new_n268), .B2(new_n269), .ZN(new_n270));
  INV_X1    g069(.A(G183gat), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n271), .A2(KEYINPUT27), .ZN(new_n272));
  INV_X1    g071(.A(KEYINPUT27), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n273), .A2(G183gat), .ZN(new_n274));
  AND4_X1   g073(.A1(KEYINPUT28), .A2(new_n272), .A3(new_n274), .A4(new_n269), .ZN(new_n275));
  NOR2_X1   g074(.A1(new_n270), .A2(new_n275), .ZN(new_n276));
  OAI21_X1  g075(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n277));
  OR3_X1    g076(.A1(KEYINPUT26), .A2(G169gat), .A3(G176gat), .ZN(new_n278));
  NAND3_X1  g077(.A1(new_n252), .A2(new_n277), .A3(new_n278), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n279), .A2(new_n236), .ZN(new_n280));
  NOR2_X1   g079(.A1(new_n276), .A2(new_n280), .ZN(new_n281));
  OAI21_X1  g080(.A(new_n234), .B1(new_n267), .B2(new_n281), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n233), .A2(new_n229), .ZN(new_n283));
  INV_X1    g082(.A(new_n215), .ZN(new_n284));
  OAI21_X1  g083(.A(new_n222), .B1(new_n284), .B2(new_n213), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n283), .A2(new_n285), .ZN(new_n286));
  INV_X1    g085(.A(new_n281), .ZN(new_n287));
  AOI21_X1  g086(.A(new_n253), .B1(new_n260), .B2(KEYINPUT66), .ZN(new_n288));
  AOI21_X1  g087(.A(KEYINPUT25), .B1(new_n288), .B2(new_n264), .ZN(new_n289));
  OAI211_X1 g088(.A(new_n286), .B(new_n287), .C1(new_n289), .C2(new_n255), .ZN(new_n290));
  NAND2_X1  g089(.A1(G227gat), .A2(G233gat), .ZN(new_n291));
  XOR2_X1   g090(.A(new_n291), .B(KEYINPUT64), .Z(new_n292));
  NAND3_X1  g091(.A1(new_n282), .A2(new_n290), .A3(new_n292), .ZN(new_n293));
  AOI21_X1  g092(.A(new_n204), .B1(new_n293), .B2(KEYINPUT32), .ZN(new_n294));
  INV_X1    g093(.A(KEYINPUT72), .ZN(new_n295));
  INV_X1    g094(.A(KEYINPUT33), .ZN(new_n296));
  NAND3_X1  g095(.A1(new_n293), .A2(new_n295), .A3(new_n296), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n294), .A2(new_n297), .ZN(new_n298));
  AOI21_X1  g097(.A(new_n295), .B1(new_n293), .B2(new_n296), .ZN(new_n299));
  OAI21_X1  g098(.A(KEYINPUT73), .B1(new_n298), .B2(new_n299), .ZN(new_n300));
  INV_X1    g099(.A(new_n299), .ZN(new_n301));
  INV_X1    g100(.A(KEYINPUT73), .ZN(new_n302));
  NAND4_X1  g101(.A1(new_n301), .A2(new_n302), .A3(new_n297), .A4(new_n294), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n300), .A2(new_n303), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n293), .A2(KEYINPUT32), .ZN(new_n305));
  NOR2_X1   g104(.A1(new_n204), .A2(new_n296), .ZN(new_n306));
  NOR2_X1   g105(.A1(new_n305), .A2(new_n306), .ZN(new_n307));
  INV_X1    g106(.A(new_n307), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n304), .A2(new_n308), .ZN(new_n309));
  INV_X1    g108(.A(KEYINPUT34), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n282), .A2(new_n290), .ZN(new_n311));
  AOI21_X1  g110(.A(new_n310), .B1(new_n311), .B2(new_n291), .ZN(new_n312));
  AOI211_X1 g111(.A(KEYINPUT34), .B(new_n292), .C1(new_n282), .C2(new_n290), .ZN(new_n313));
  NOR2_X1   g112(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  INV_X1    g113(.A(new_n314), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n309), .A2(new_n315), .ZN(new_n316));
  INV_X1    g115(.A(KEYINPUT75), .ZN(new_n317));
  AOI21_X1  g116(.A(new_n307), .B1(new_n300), .B2(new_n303), .ZN(new_n318));
  AOI21_X1  g117(.A(new_n317), .B1(new_n318), .B2(new_n314), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n316), .A2(new_n319), .ZN(new_n320));
  INV_X1    g119(.A(KEYINPUT36), .ZN(new_n321));
  NAND3_X1  g120(.A1(new_n309), .A2(new_n317), .A3(new_n315), .ZN(new_n322));
  NAND3_X1  g121(.A1(new_n320), .A2(new_n321), .A3(new_n322), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n318), .A2(new_n314), .ZN(new_n324));
  INV_X1    g123(.A(KEYINPUT74), .ZN(new_n325));
  OAI21_X1  g124(.A(new_n315), .B1(new_n318), .B2(new_n325), .ZN(new_n326));
  AOI211_X1 g125(.A(KEYINPUT74), .B(new_n307), .C1(new_n300), .C2(new_n303), .ZN(new_n327));
  OAI211_X1 g126(.A(KEYINPUT36), .B(new_n324), .C1(new_n326), .C2(new_n327), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n323), .A2(new_n328), .ZN(new_n329));
  XNOR2_X1  g128(.A(G78gat), .B(G106gat), .ZN(new_n330));
  INV_X1    g129(.A(G50gat), .ZN(new_n331));
  XNOR2_X1  g130(.A(new_n330), .B(new_n331), .ZN(new_n332));
  AND2_X1   g131(.A1(G228gat), .A2(G233gat), .ZN(new_n333));
  OR2_X1    g132(.A1(KEYINPUT76), .A2(KEYINPUT22), .ZN(new_n334));
  NAND2_X1  g133(.A1(G211gat), .A2(G218gat), .ZN(new_n335));
  NAND2_X1  g134(.A1(KEYINPUT76), .A2(KEYINPUT22), .ZN(new_n336));
  NAND3_X1  g135(.A1(new_n334), .A2(new_n335), .A3(new_n336), .ZN(new_n337));
  INV_X1    g136(.A(G211gat), .ZN(new_n338));
  INV_X1    g137(.A(G218gat), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n338), .A2(new_n339), .ZN(new_n340));
  NAND3_X1  g139(.A1(new_n340), .A2(KEYINPUT77), .A3(new_n335), .ZN(new_n341));
  XNOR2_X1  g140(.A(G197gat), .B(G204gat), .ZN(new_n342));
  NAND3_X1  g141(.A1(new_n337), .A2(new_n341), .A3(new_n342), .ZN(new_n343));
  AOI21_X1  g142(.A(KEYINPUT77), .B1(new_n340), .B2(new_n335), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n340), .A2(new_n335), .ZN(new_n346));
  INV_X1    g145(.A(KEYINPUT77), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n346), .A2(new_n347), .ZN(new_n348));
  NAND4_X1  g147(.A1(new_n348), .A2(new_n337), .A3(new_n341), .A4(new_n342), .ZN(new_n349));
  INV_X1    g148(.A(KEYINPUT29), .ZN(new_n350));
  NAND3_X1  g149(.A1(new_n345), .A2(new_n349), .A3(new_n350), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n351), .A2(KEYINPUT85), .ZN(new_n352));
  INV_X1    g151(.A(KEYINPUT3), .ZN(new_n353));
  INV_X1    g152(.A(KEYINPUT85), .ZN(new_n354));
  NAND4_X1  g153(.A1(new_n345), .A2(new_n349), .A3(new_n354), .A4(new_n350), .ZN(new_n355));
  NAND3_X1  g154(.A1(new_n352), .A2(new_n353), .A3(new_n355), .ZN(new_n356));
  INV_X1    g155(.A(G141gat), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n357), .A2(G148gat), .ZN(new_n358));
  INV_X1    g157(.A(G148gat), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n359), .A2(G141gat), .ZN(new_n360));
  NAND2_X1  g159(.A1(G155gat), .A2(G162gat), .ZN(new_n361));
  AOI22_X1  g160(.A1(new_n358), .A2(new_n360), .B1(KEYINPUT2), .B2(new_n361), .ZN(new_n362));
  OAI21_X1  g161(.A(KEYINPUT79), .B1(G155gat), .B2(G162gat), .ZN(new_n363));
  INV_X1    g162(.A(new_n363), .ZN(new_n364));
  NOR3_X1   g163(.A1(KEYINPUT79), .A2(G155gat), .A3(G162gat), .ZN(new_n365));
  OAI21_X1  g164(.A(new_n361), .B1(new_n364), .B2(new_n365), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n366), .A2(KEYINPUT80), .ZN(new_n367));
  INV_X1    g166(.A(KEYINPUT79), .ZN(new_n368));
  INV_X1    g167(.A(G155gat), .ZN(new_n369));
  INV_X1    g168(.A(G162gat), .ZN(new_n370));
  NAND3_X1  g169(.A1(new_n368), .A2(new_n369), .A3(new_n370), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n371), .A2(new_n363), .ZN(new_n372));
  INV_X1    g171(.A(KEYINPUT80), .ZN(new_n373));
  NAND3_X1  g172(.A1(new_n372), .A2(new_n373), .A3(new_n361), .ZN(new_n374));
  AOI21_X1  g173(.A(new_n362), .B1(new_n367), .B2(new_n374), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n369), .A2(new_n370), .ZN(new_n376));
  NAND3_X1  g175(.A1(new_n362), .A2(new_n361), .A3(new_n376), .ZN(new_n377));
  INV_X1    g176(.A(new_n377), .ZN(new_n378));
  NOR2_X1   g177(.A1(new_n375), .A2(new_n378), .ZN(new_n379));
  AOI21_X1  g178(.A(new_n333), .B1(new_n356), .B2(new_n379), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n345), .A2(new_n349), .ZN(new_n381));
  INV_X1    g180(.A(new_n362), .ZN(new_n382));
  AOI21_X1  g181(.A(new_n373), .B1(new_n372), .B2(new_n361), .ZN(new_n383));
  AND2_X1   g182(.A1(G155gat), .A2(G162gat), .ZN(new_n384));
  AOI211_X1 g183(.A(KEYINPUT80), .B(new_n384), .C1(new_n371), .C2(new_n363), .ZN(new_n385));
  OAI21_X1  g184(.A(new_n382), .B1(new_n383), .B2(new_n385), .ZN(new_n386));
  AOI21_X1  g185(.A(KEYINPUT3), .B1(new_n386), .B2(new_n377), .ZN(new_n387));
  OAI21_X1  g186(.A(new_n381), .B1(new_n387), .B2(KEYINPUT29), .ZN(new_n388));
  INV_X1    g187(.A(KEYINPUT86), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n388), .A2(new_n389), .ZN(new_n390));
  OAI211_X1 g189(.A(KEYINPUT86), .B(new_n381), .C1(new_n387), .C2(KEYINPUT29), .ZN(new_n391));
  NAND3_X1  g190(.A1(new_n380), .A2(new_n390), .A3(new_n391), .ZN(new_n392));
  INV_X1    g191(.A(new_n388), .ZN(new_n393));
  OAI21_X1  g192(.A(KEYINPUT81), .B1(new_n375), .B2(new_n378), .ZN(new_n394));
  INV_X1    g193(.A(KEYINPUT81), .ZN(new_n395));
  NAND3_X1  g194(.A1(new_n386), .A2(new_n395), .A3(new_n377), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n351), .A2(new_n353), .ZN(new_n397));
  AND3_X1   g196(.A1(new_n394), .A2(new_n396), .A3(new_n397), .ZN(new_n398));
  OAI21_X1  g197(.A(new_n333), .B1(new_n393), .B2(new_n398), .ZN(new_n399));
  INV_X1    g198(.A(G22gat), .ZN(new_n400));
  NAND3_X1  g199(.A1(new_n392), .A2(new_n399), .A3(new_n400), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n401), .A2(KEYINPUT84), .ZN(new_n402));
  AOI21_X1  g201(.A(new_n400), .B1(new_n392), .B2(new_n399), .ZN(new_n403));
  OAI21_X1  g202(.A(new_n332), .B1(new_n402), .B2(new_n403), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n392), .A2(new_n399), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n405), .A2(G22gat), .ZN(new_n406));
  INV_X1    g205(.A(new_n332), .ZN(new_n407));
  NAND4_X1  g206(.A1(new_n406), .A2(KEYINPUT84), .A3(new_n407), .A4(new_n401), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n404), .A2(new_n408), .ZN(new_n409));
  XNOR2_X1  g208(.A(KEYINPUT83), .B(KEYINPUT31), .ZN(new_n410));
  INV_X1    g209(.A(new_n410), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n409), .A2(new_n411), .ZN(new_n412));
  NAND3_X1  g211(.A1(new_n404), .A2(new_n410), .A3(new_n408), .ZN(new_n413));
  AND2_X1   g212(.A1(new_n412), .A2(new_n413), .ZN(new_n414));
  INV_X1    g213(.A(new_n414), .ZN(new_n415));
  XOR2_X1   g214(.A(G8gat), .B(G36gat), .Z(new_n416));
  XNOR2_X1  g215(.A(new_n416), .B(KEYINPUT78), .ZN(new_n417));
  XNOR2_X1  g216(.A(G64gat), .B(G92gat), .ZN(new_n418));
  XNOR2_X1  g217(.A(new_n417), .B(new_n418), .ZN(new_n419));
  INV_X1    g218(.A(G226gat), .ZN(new_n420));
  INV_X1    g219(.A(G233gat), .ZN(new_n421));
  NOR2_X1   g220(.A1(new_n420), .A2(new_n421), .ZN(new_n422));
  INV_X1    g221(.A(new_n422), .ZN(new_n423));
  OAI21_X1  g222(.A(new_n265), .B1(new_n262), .B2(new_n263), .ZN(new_n424));
  AND3_X1   g223(.A1(new_n259), .A2(new_n263), .A3(new_n237), .ZN(new_n425));
  OAI21_X1  g224(.A(new_n254), .B1(new_n424), .B2(new_n425), .ZN(new_n426));
  OAI211_X1 g225(.A(new_n265), .B(KEYINPUT25), .C1(new_n238), .C2(new_n240), .ZN(new_n427));
  AOI21_X1  g226(.A(new_n281), .B1(new_n426), .B2(new_n427), .ZN(new_n428));
  OAI21_X1  g227(.A(new_n423), .B1(new_n428), .B2(KEYINPUT29), .ZN(new_n429));
  OAI21_X1  g228(.A(new_n422), .B1(new_n267), .B2(new_n281), .ZN(new_n430));
  AND3_X1   g229(.A1(new_n429), .A2(new_n381), .A3(new_n430), .ZN(new_n431));
  AOI21_X1  g230(.A(new_n381), .B1(new_n429), .B2(new_n430), .ZN(new_n432));
  OAI21_X1  g231(.A(new_n419), .B1(new_n431), .B2(new_n432), .ZN(new_n433));
  INV_X1    g232(.A(new_n381), .ZN(new_n434));
  OAI21_X1  g233(.A(new_n287), .B1(new_n289), .B2(new_n255), .ZN(new_n435));
  AOI21_X1  g234(.A(new_n422), .B1(new_n435), .B2(new_n350), .ZN(new_n436));
  NOR2_X1   g235(.A1(new_n428), .A2(new_n423), .ZN(new_n437));
  OAI21_X1  g236(.A(new_n434), .B1(new_n436), .B2(new_n437), .ZN(new_n438));
  INV_X1    g237(.A(new_n419), .ZN(new_n439));
  NAND3_X1  g238(.A1(new_n429), .A2(new_n381), .A3(new_n430), .ZN(new_n440));
  NAND3_X1  g239(.A1(new_n438), .A2(new_n439), .A3(new_n440), .ZN(new_n441));
  NAND3_X1  g240(.A1(new_n433), .A2(new_n441), .A3(KEYINPUT30), .ZN(new_n442));
  INV_X1    g241(.A(KEYINPUT30), .ZN(new_n443));
  OAI211_X1 g242(.A(new_n443), .B(new_n419), .C1(new_n431), .C2(new_n432), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n442), .A2(new_n444), .ZN(new_n445));
  INV_X1    g244(.A(KEYINPUT4), .ZN(new_n446));
  NOR3_X1   g245(.A1(new_n286), .A2(new_n379), .A3(new_n446), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n386), .A2(new_n377), .ZN(new_n448));
  AOI21_X1  g247(.A(KEYINPUT4), .B1(new_n234), .B2(new_n448), .ZN(new_n449));
  NOR2_X1   g248(.A1(new_n447), .A2(new_n449), .ZN(new_n450));
  NAND2_X1  g249(.A1(G225gat), .A2(G233gat), .ZN(new_n451));
  NAND3_X1  g250(.A1(new_n394), .A2(KEYINPUT3), .A3(new_n396), .ZN(new_n452));
  AOI22_X1  g251(.A1(new_n448), .A2(new_n353), .B1(new_n283), .B2(new_n285), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  NAND4_X1  g253(.A1(new_n450), .A2(KEYINPUT5), .A3(new_n451), .A4(new_n454), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n234), .A2(new_n448), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n456), .A2(new_n446), .ZN(new_n457));
  NAND3_X1  g256(.A1(new_n234), .A2(KEYINPUT4), .A3(new_n448), .ZN(new_n458));
  NAND4_X1  g257(.A1(new_n454), .A2(new_n457), .A3(new_n451), .A4(new_n458), .ZN(new_n459));
  INV_X1    g258(.A(new_n459), .ZN(new_n460));
  NAND3_X1  g259(.A1(new_n394), .A2(new_n286), .A3(new_n396), .ZN(new_n461));
  AOI21_X1  g260(.A(new_n451), .B1(new_n461), .B2(new_n456), .ZN(new_n462));
  INV_X1    g261(.A(KEYINPUT5), .ZN(new_n463));
  NOR2_X1   g262(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  OAI21_X1  g263(.A(new_n455), .B1(new_n460), .B2(new_n464), .ZN(new_n465));
  XOR2_X1   g264(.A(G1gat), .B(G29gat), .Z(new_n466));
  XNOR2_X1  g265(.A(G57gat), .B(G85gat), .ZN(new_n467));
  XNOR2_X1  g266(.A(new_n466), .B(new_n467), .ZN(new_n468));
  XNOR2_X1  g267(.A(KEYINPUT82), .B(KEYINPUT0), .ZN(new_n469));
  XOR2_X1   g268(.A(new_n468), .B(new_n469), .Z(new_n470));
  INV_X1    g269(.A(new_n470), .ZN(new_n471));
  AOI21_X1  g270(.A(KEYINPUT6), .B1(new_n465), .B2(new_n471), .ZN(new_n472));
  OAI21_X1  g271(.A(new_n459), .B1(new_n463), .B2(new_n462), .ZN(new_n473));
  NAND3_X1  g272(.A1(new_n473), .A2(new_n470), .A3(new_n455), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n472), .A2(new_n474), .ZN(new_n475));
  INV_X1    g274(.A(new_n475), .ZN(new_n476));
  INV_X1    g275(.A(KEYINPUT6), .ZN(new_n477));
  NOR2_X1   g276(.A1(new_n474), .A2(new_n477), .ZN(new_n478));
  OAI21_X1  g277(.A(new_n445), .B1(new_n476), .B2(new_n478), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n415), .A2(new_n479), .ZN(new_n480));
  NAND3_X1  g279(.A1(new_n461), .A2(new_n456), .A3(new_n451), .ZN(new_n481));
  NAND2_X1  g280(.A1(new_n481), .A2(KEYINPUT39), .ZN(new_n482));
  INV_X1    g281(.A(KEYINPUT89), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  NAND3_X1  g283(.A1(new_n481), .A2(KEYINPUT89), .A3(KEYINPUT39), .ZN(new_n485));
  AND2_X1   g284(.A1(new_n450), .A2(new_n454), .ZN(new_n486));
  OAI211_X1 g285(.A(new_n484), .B(new_n485), .C1(new_n486), .C2(new_n451), .ZN(new_n487));
  XNOR2_X1  g286(.A(new_n470), .B(KEYINPUT88), .ZN(new_n488));
  AOI21_X1  g287(.A(new_n451), .B1(new_n450), .B2(new_n454), .ZN(new_n489));
  INV_X1    g288(.A(KEYINPUT39), .ZN(new_n490));
  AOI21_X1  g289(.A(new_n488), .B1(new_n489), .B2(new_n490), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n487), .A2(new_n491), .ZN(new_n492));
  INV_X1    g291(.A(KEYINPUT40), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  NAND3_X1  g293(.A1(new_n473), .A2(new_n455), .A3(new_n488), .ZN(new_n495));
  NAND3_X1  g294(.A1(new_n487), .A2(new_n491), .A3(KEYINPUT40), .ZN(new_n496));
  AND3_X1   g295(.A1(new_n494), .A2(new_n495), .A3(new_n496), .ZN(new_n497));
  INV_X1    g296(.A(KEYINPUT90), .ZN(new_n498));
  NAND3_X1  g297(.A1(new_n442), .A2(KEYINPUT87), .A3(new_n444), .ZN(new_n499));
  INV_X1    g298(.A(KEYINPUT87), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n445), .A2(new_n500), .ZN(new_n501));
  NAND4_X1  g300(.A1(new_n497), .A2(new_n498), .A3(new_n499), .A4(new_n501), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n501), .A2(new_n499), .ZN(new_n503));
  NAND3_X1  g302(.A1(new_n494), .A2(new_n495), .A3(new_n496), .ZN(new_n504));
  OAI21_X1  g303(.A(KEYINPUT90), .B1(new_n503), .B2(new_n504), .ZN(new_n505));
  OAI21_X1  g304(.A(KEYINPUT37), .B1(new_n431), .B2(new_n432), .ZN(new_n506));
  INV_X1    g305(.A(KEYINPUT37), .ZN(new_n507));
  NAND3_X1  g306(.A1(new_n438), .A2(new_n507), .A3(new_n440), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n506), .A2(new_n508), .ZN(new_n509));
  INV_X1    g308(.A(KEYINPUT38), .ZN(new_n510));
  NAND3_X1  g309(.A1(new_n509), .A2(new_n510), .A3(new_n439), .ZN(new_n511));
  INV_X1    g310(.A(KEYINPUT91), .ZN(new_n512));
  NAND2_X1  g311(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  NAND4_X1  g312(.A1(new_n509), .A2(KEYINPUT91), .A3(new_n510), .A4(new_n439), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  AOI21_X1  g314(.A(new_n478), .B1(new_n472), .B2(new_n495), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n509), .A2(new_n439), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n517), .A2(KEYINPUT38), .ZN(new_n518));
  NAND4_X1  g317(.A1(new_n515), .A2(new_n516), .A3(new_n433), .A4(new_n518), .ZN(new_n519));
  NAND4_X1  g318(.A1(new_n502), .A2(new_n505), .A3(new_n519), .A4(new_n414), .ZN(new_n520));
  NAND3_X1  g319(.A1(new_n329), .A2(new_n480), .A3(new_n520), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n320), .A2(new_n322), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n465), .A2(new_n471), .ZN(new_n523));
  NAND3_X1  g322(.A1(new_n523), .A2(new_n477), .A3(new_n495), .ZN(new_n524));
  OR2_X1    g323(.A1(new_n474), .A2(new_n477), .ZN(new_n525));
  AOI21_X1  g324(.A(KEYINPUT35), .B1(new_n524), .B2(new_n525), .ZN(new_n526));
  AND4_X1   g325(.A1(new_n413), .A2(new_n526), .A3(new_n503), .A4(new_n412), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n522), .A2(new_n527), .ZN(new_n528));
  NOR2_X1   g327(.A1(new_n326), .A2(new_n327), .ZN(new_n529));
  NAND3_X1  g328(.A1(new_n412), .A2(new_n324), .A3(new_n413), .ZN(new_n530));
  NOR3_X1   g329(.A1(new_n529), .A2(new_n530), .A3(new_n479), .ZN(new_n531));
  INV_X1    g330(.A(KEYINPUT35), .ZN(new_n532));
  OAI21_X1  g331(.A(new_n528), .B1(new_n531), .B2(new_n532), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n521), .A2(new_n533), .ZN(new_n534));
  AND2_X1   g333(.A1(G232gat), .A2(G233gat), .ZN(new_n535));
  NOR2_X1   g334(.A1(new_n535), .A2(KEYINPUT41), .ZN(new_n536));
  XNOR2_X1  g335(.A(new_n536), .B(KEYINPUT106), .ZN(new_n537));
  XNOR2_X1  g336(.A(G134gat), .B(G162gat), .ZN(new_n538));
  XNOR2_X1  g337(.A(new_n537), .B(new_n538), .ZN(new_n539));
  INV_X1    g338(.A(new_n539), .ZN(new_n540));
  INV_X1    g339(.A(KEYINPUT96), .ZN(new_n541));
  XNOR2_X1  g340(.A(G43gat), .B(G50gat), .ZN(new_n542));
  NAND2_X1  g341(.A1(new_n542), .A2(KEYINPUT15), .ZN(new_n543));
  INV_X1    g342(.A(KEYINPUT95), .ZN(new_n544));
  XNOR2_X1  g343(.A(new_n543), .B(new_n544), .ZN(new_n545));
  NOR2_X1   g344(.A1(new_n542), .A2(KEYINPUT15), .ZN(new_n546));
  NAND2_X1  g345(.A1(G29gat), .A2(G36gat), .ZN(new_n547));
  INV_X1    g346(.A(KEYINPUT94), .ZN(new_n548));
  XNOR2_X1  g347(.A(new_n547), .B(new_n548), .ZN(new_n549));
  NOR2_X1   g348(.A1(new_n546), .A2(new_n549), .ZN(new_n550));
  NOR2_X1   g349(.A1(G29gat), .A2(G36gat), .ZN(new_n551));
  XOR2_X1   g350(.A(new_n551), .B(KEYINPUT14), .Z(new_n552));
  NAND2_X1  g351(.A1(new_n550), .A2(new_n552), .ZN(new_n553));
  OAI21_X1  g352(.A(new_n541), .B1(new_n545), .B2(new_n553), .ZN(new_n554));
  XNOR2_X1  g353(.A(new_n543), .B(KEYINPUT95), .ZN(new_n555));
  NAND4_X1  g354(.A1(new_n555), .A2(KEYINPUT96), .A3(new_n552), .A4(new_n550), .ZN(new_n556));
  INV_X1    g355(.A(new_n543), .ZN(new_n557));
  XNOR2_X1  g356(.A(new_n551), .B(KEYINPUT14), .ZN(new_n558));
  AOI21_X1  g357(.A(new_n549), .B1(new_n558), .B2(KEYINPUT93), .ZN(new_n559));
  OAI21_X1  g358(.A(new_n559), .B1(KEYINPUT93), .B2(new_n558), .ZN(new_n560));
  AOI22_X1  g359(.A1(new_n554), .A2(new_n556), .B1(new_n557), .B2(new_n560), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n561), .A2(KEYINPUT17), .ZN(new_n562));
  XNOR2_X1  g361(.A(new_n562), .B(KEYINPUT99), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n554), .A2(new_n556), .ZN(new_n564));
  NAND2_X1  g363(.A1(new_n560), .A2(new_n557), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  INV_X1    g365(.A(KEYINPUT97), .ZN(new_n567));
  INV_X1    g366(.A(KEYINPUT17), .ZN(new_n568));
  NAND3_X1  g367(.A1(new_n566), .A2(new_n567), .A3(new_n568), .ZN(new_n569));
  OAI21_X1  g368(.A(KEYINPUT97), .B1(new_n561), .B2(KEYINPUT17), .ZN(new_n570));
  NAND2_X1  g369(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  NAND2_X1  g370(.A1(G85gat), .A2(G92gat), .ZN(new_n572));
  XNOR2_X1  g371(.A(new_n572), .B(KEYINPUT7), .ZN(new_n573));
  NAND2_X1  g372(.A1(G99gat), .A2(G106gat), .ZN(new_n574));
  INV_X1    g373(.A(G85gat), .ZN(new_n575));
  INV_X1    g374(.A(G92gat), .ZN(new_n576));
  AOI22_X1  g375(.A1(KEYINPUT8), .A2(new_n574), .B1(new_n575), .B2(new_n576), .ZN(new_n577));
  NAND2_X1  g376(.A1(new_n573), .A2(new_n577), .ZN(new_n578));
  XNOR2_X1  g377(.A(G99gat), .B(G106gat), .ZN(new_n579));
  XNOR2_X1  g378(.A(new_n578), .B(new_n579), .ZN(new_n580));
  INV_X1    g379(.A(new_n580), .ZN(new_n581));
  NAND3_X1  g380(.A1(new_n563), .A2(new_n571), .A3(new_n581), .ZN(new_n582));
  XOR2_X1   g381(.A(G190gat), .B(G218gat), .Z(new_n583));
  INV_X1    g382(.A(new_n583), .ZN(new_n584));
  AOI22_X1  g383(.A1(new_n566), .A2(new_n580), .B1(KEYINPUT41), .B2(new_n535), .ZN(new_n585));
  NAND3_X1  g384(.A1(new_n582), .A2(new_n584), .A3(new_n585), .ZN(new_n586));
  INV_X1    g385(.A(new_n586), .ZN(new_n587));
  AOI21_X1  g386(.A(new_n584), .B1(new_n582), .B2(new_n585), .ZN(new_n588));
  OAI21_X1  g387(.A(new_n540), .B1(new_n587), .B2(new_n588), .ZN(new_n589));
  INV_X1    g388(.A(new_n588), .ZN(new_n590));
  NAND3_X1  g389(.A1(new_n590), .A2(new_n586), .A3(new_n539), .ZN(new_n591));
  AND2_X1   g390(.A1(new_n589), .A2(new_n591), .ZN(new_n592));
  XOR2_X1   g391(.A(G183gat), .B(G211gat), .Z(new_n593));
  XOR2_X1   g392(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n594));
  OR2_X1    g393(.A1(G57gat), .A2(G64gat), .ZN(new_n595));
  NAND2_X1  g394(.A1(G57gat), .A2(G64gat), .ZN(new_n596));
  AND2_X1   g395(.A1(G71gat), .A2(G78gat), .ZN(new_n597));
  OAI211_X1 g396(.A(new_n595), .B(new_n596), .C1(new_n597), .C2(KEYINPUT9), .ZN(new_n598));
  INV_X1    g397(.A(KEYINPUT101), .ZN(new_n599));
  OAI21_X1  g398(.A(new_n598), .B1(new_n599), .B2(new_n597), .ZN(new_n600));
  NOR2_X1   g399(.A1(G71gat), .A2(G78gat), .ZN(new_n601));
  NOR2_X1   g400(.A1(new_n597), .A2(new_n601), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n600), .A2(new_n602), .ZN(new_n603));
  INV_X1    g402(.A(new_n602), .ZN(new_n604));
  OAI211_X1 g403(.A(new_n604), .B(new_n598), .C1(new_n599), .C2(new_n597), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n603), .A2(new_n605), .ZN(new_n606));
  INV_X1    g405(.A(KEYINPUT102), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  NAND3_X1  g407(.A1(new_n603), .A2(KEYINPUT102), .A3(new_n605), .ZN(new_n609));
  NAND2_X1  g408(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  XNOR2_X1  g409(.A(KEYINPUT103), .B(KEYINPUT21), .ZN(new_n611));
  NAND2_X1  g410(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  INV_X1    g411(.A(G231gat), .ZN(new_n613));
  NOR2_X1   g412(.A1(new_n613), .A2(new_n421), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n612), .A2(new_n614), .ZN(new_n615));
  INV_X1    g414(.A(new_n615), .ZN(new_n616));
  OAI211_X1 g415(.A(new_n610), .B(new_n611), .C1(new_n613), .C2(new_n421), .ZN(new_n617));
  INV_X1    g416(.A(new_n617), .ZN(new_n618));
  OAI21_X1  g417(.A(new_n594), .B1(new_n616), .B2(new_n618), .ZN(new_n619));
  INV_X1    g418(.A(new_n619), .ZN(new_n620));
  NOR3_X1   g419(.A1(new_n616), .A2(new_n618), .A3(new_n594), .ZN(new_n621));
  OAI21_X1  g420(.A(new_n593), .B1(new_n620), .B2(new_n621), .ZN(new_n622));
  INV_X1    g421(.A(new_n621), .ZN(new_n623));
  INV_X1    g422(.A(new_n593), .ZN(new_n624));
  NAND3_X1  g423(.A1(new_n623), .A2(new_n624), .A3(new_n619), .ZN(new_n625));
  XNOR2_X1  g424(.A(G15gat), .B(G22gat), .ZN(new_n626));
  INV_X1    g425(.A(KEYINPUT98), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  XNOR2_X1  g427(.A(new_n628), .B(G8gat), .ZN(new_n629));
  INV_X1    g428(.A(KEYINPUT16), .ZN(new_n630));
  AOI21_X1  g429(.A(G1gat), .B1(new_n626), .B2(new_n630), .ZN(new_n631));
  XNOR2_X1  g430(.A(new_n629), .B(new_n631), .ZN(new_n632));
  INV_X1    g431(.A(new_n632), .ZN(new_n633));
  INV_X1    g432(.A(KEYINPUT21), .ZN(new_n634));
  OAI21_X1  g433(.A(new_n633), .B1(new_n634), .B2(new_n610), .ZN(new_n635));
  XOR2_X1   g434(.A(G127gat), .B(G155gat), .Z(new_n636));
  XNOR2_X1  g435(.A(KEYINPUT104), .B(KEYINPUT105), .ZN(new_n637));
  XNOR2_X1  g436(.A(new_n636), .B(new_n637), .ZN(new_n638));
  XNOR2_X1  g437(.A(new_n635), .B(new_n638), .ZN(new_n639));
  AND3_X1   g438(.A1(new_n622), .A2(new_n625), .A3(new_n639), .ZN(new_n640));
  AOI21_X1  g439(.A(new_n639), .B1(new_n622), .B2(new_n625), .ZN(new_n641));
  NOR2_X1   g440(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n592), .A2(new_n642), .ZN(new_n643));
  NAND2_X1  g442(.A1(new_n566), .A2(new_n632), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n633), .A2(new_n561), .ZN(new_n645));
  NAND3_X1  g444(.A1(new_n644), .A2(new_n645), .A3(KEYINPUT100), .ZN(new_n646));
  NAND2_X1  g445(.A1(G229gat), .A2(G233gat), .ZN(new_n647));
  XOR2_X1   g446(.A(new_n647), .B(KEYINPUT13), .Z(new_n648));
  INV_X1    g447(.A(KEYINPUT100), .ZN(new_n649));
  NAND3_X1  g448(.A1(new_n566), .A2(new_n649), .A3(new_n632), .ZN(new_n650));
  AND3_X1   g449(.A1(new_n646), .A2(new_n648), .A3(new_n650), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n571), .A2(new_n633), .ZN(new_n652));
  INV_X1    g451(.A(KEYINPUT99), .ZN(new_n653));
  XNOR2_X1  g452(.A(new_n562), .B(new_n653), .ZN(new_n654));
  OAI211_X1 g453(.A(new_n647), .B(new_n644), .C1(new_n652), .C2(new_n654), .ZN(new_n655));
  INV_X1    g454(.A(KEYINPUT18), .ZN(new_n656));
  AOI21_X1  g455(.A(new_n651), .B1(new_n655), .B2(new_n656), .ZN(new_n657));
  NAND3_X1  g456(.A1(new_n563), .A2(new_n633), .A3(new_n571), .ZN(new_n658));
  NAND4_X1  g457(.A1(new_n658), .A2(KEYINPUT18), .A3(new_n647), .A4(new_n644), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n657), .A2(new_n659), .ZN(new_n660));
  XNOR2_X1  g459(.A(G113gat), .B(G141gat), .ZN(new_n661));
  XNOR2_X1  g460(.A(KEYINPUT92), .B(KEYINPUT11), .ZN(new_n662));
  XNOR2_X1  g461(.A(new_n661), .B(new_n662), .ZN(new_n663));
  XOR2_X1   g462(.A(G169gat), .B(G197gat), .Z(new_n664));
  XNOR2_X1  g463(.A(new_n663), .B(new_n664), .ZN(new_n665));
  XNOR2_X1  g464(.A(new_n665), .B(KEYINPUT12), .ZN(new_n666));
  INV_X1    g465(.A(new_n666), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n660), .A2(new_n667), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n655), .A2(new_n656), .ZN(new_n669));
  INV_X1    g468(.A(new_n651), .ZN(new_n670));
  NAND4_X1  g469(.A1(new_n669), .A2(new_n659), .A3(new_n670), .A4(new_n666), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n668), .A2(new_n671), .ZN(new_n672));
  INV_X1    g471(.A(new_n672), .ZN(new_n673));
  NAND2_X1  g472(.A1(G230gat), .A2(G233gat), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n580), .A2(KEYINPUT10), .ZN(new_n675));
  INV_X1    g474(.A(new_n675), .ZN(new_n676));
  INV_X1    g475(.A(KEYINPUT107), .ZN(new_n677));
  NAND4_X1  g476(.A1(new_n676), .A2(new_n608), .A3(new_n677), .A4(new_n609), .ZN(new_n678));
  OAI21_X1  g477(.A(KEYINPUT107), .B1(new_n610), .B2(new_n675), .ZN(new_n679));
  NAND2_X1  g478(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  NAND3_X1  g479(.A1(new_n581), .A2(new_n608), .A3(new_n609), .ZN(new_n681));
  NAND3_X1  g480(.A1(new_n580), .A2(new_n603), .A3(new_n605), .ZN(new_n682));
  AOI21_X1  g481(.A(KEYINPUT10), .B1(new_n681), .B2(new_n682), .ZN(new_n683));
  OAI21_X1  g482(.A(new_n674), .B1(new_n680), .B2(new_n683), .ZN(new_n684));
  INV_X1    g483(.A(new_n674), .ZN(new_n685));
  NAND3_X1  g484(.A1(new_n681), .A2(new_n685), .A3(new_n682), .ZN(new_n686));
  AND2_X1   g485(.A1(new_n684), .A2(new_n686), .ZN(new_n687));
  XNOR2_X1  g486(.A(G120gat), .B(G148gat), .ZN(new_n688));
  XNOR2_X1  g487(.A(G176gat), .B(G204gat), .ZN(new_n689));
  XOR2_X1   g488(.A(new_n688), .B(new_n689), .Z(new_n690));
  OR2_X1    g489(.A1(new_n687), .A2(new_n690), .ZN(new_n691));
  NAND2_X1  g490(.A1(new_n684), .A2(KEYINPUT108), .ZN(new_n692));
  INV_X1    g491(.A(KEYINPUT108), .ZN(new_n693));
  OAI211_X1 g492(.A(new_n693), .B(new_n674), .C1(new_n680), .C2(new_n683), .ZN(new_n694));
  AND2_X1   g493(.A1(new_n686), .A2(new_n690), .ZN(new_n695));
  NAND3_X1  g494(.A1(new_n692), .A2(new_n694), .A3(new_n695), .ZN(new_n696));
  NAND2_X1  g495(.A1(new_n691), .A2(new_n696), .ZN(new_n697));
  NOR3_X1   g496(.A1(new_n643), .A2(new_n673), .A3(new_n697), .ZN(new_n698));
  AND2_X1   g497(.A1(new_n534), .A2(new_n698), .ZN(new_n699));
  NOR2_X1   g498(.A1(new_n476), .A2(new_n478), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  XNOR2_X1  g500(.A(new_n701), .B(G1gat), .ZN(G1324gat));
  INV_X1    g501(.A(KEYINPUT42), .ZN(new_n703));
  INV_X1    g502(.A(new_n503), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n699), .A2(new_n704), .ZN(new_n705));
  XNOR2_X1  g504(.A(new_n705), .B(KEYINPUT109), .ZN(new_n706));
  XNOR2_X1  g505(.A(KEYINPUT16), .B(G8gat), .ZN(new_n707));
  OAI21_X1  g506(.A(new_n703), .B1(new_n706), .B2(new_n707), .ZN(new_n708));
  NAND2_X1  g507(.A1(new_n706), .A2(G8gat), .ZN(new_n709));
  OR3_X1    g508(.A1(new_n705), .A2(new_n703), .A3(new_n707), .ZN(new_n710));
  NAND3_X1  g509(.A1(new_n708), .A2(new_n709), .A3(new_n710), .ZN(G1325gat));
  INV_X1    g510(.A(G15gat), .ZN(new_n712));
  NAND3_X1  g511(.A1(new_n699), .A2(new_n712), .A3(new_n522), .ZN(new_n713));
  INV_X1    g512(.A(new_n329), .ZN(new_n714));
  AND2_X1   g513(.A1(new_n699), .A2(new_n714), .ZN(new_n715));
  OAI21_X1  g514(.A(new_n713), .B1(new_n715), .B2(new_n712), .ZN(G1326gat));
  NAND2_X1  g515(.A1(new_n699), .A2(new_n415), .ZN(new_n717));
  XNOR2_X1  g516(.A(KEYINPUT43), .B(G22gat), .ZN(new_n718));
  XNOR2_X1  g517(.A(new_n717), .B(new_n718), .ZN(G1327gat));
  AND3_X1   g518(.A1(new_n412), .A2(new_n324), .A3(new_n413), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n309), .A2(KEYINPUT74), .ZN(new_n721));
  NAND2_X1  g520(.A1(new_n318), .A2(new_n325), .ZN(new_n722));
  NAND3_X1  g521(.A1(new_n721), .A2(new_n722), .A3(new_n315), .ZN(new_n723));
  AOI22_X1  g522(.A1(new_n475), .A2(new_n525), .B1(new_n444), .B2(new_n442), .ZN(new_n724));
  NAND3_X1  g523(.A1(new_n720), .A2(new_n723), .A3(new_n724), .ZN(new_n725));
  NAND2_X1  g524(.A1(new_n725), .A2(KEYINPUT35), .ZN(new_n726));
  INV_X1    g525(.A(KEYINPUT110), .ZN(new_n727));
  AND3_X1   g526(.A1(new_n726), .A2(new_n727), .A3(new_n528), .ZN(new_n728));
  AOI21_X1  g527(.A(new_n727), .B1(new_n726), .B2(new_n528), .ZN(new_n729));
  OAI21_X1  g528(.A(new_n521), .B1(new_n728), .B2(new_n729), .ZN(new_n730));
  NOR2_X1   g529(.A1(new_n592), .A2(KEYINPUT44), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n589), .A2(new_n591), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n534), .A2(new_n732), .ZN(new_n733));
  AOI22_X1  g532(.A1(new_n730), .A2(new_n731), .B1(new_n733), .B2(KEYINPUT44), .ZN(new_n734));
  NOR3_X1   g533(.A1(new_n673), .A2(new_n642), .A3(new_n697), .ZN(new_n735));
  INV_X1    g534(.A(new_n735), .ZN(new_n736));
  OAI21_X1  g535(.A(KEYINPUT111), .B1(new_n734), .B2(new_n736), .ZN(new_n737));
  INV_X1    g536(.A(KEYINPUT111), .ZN(new_n738));
  INV_X1    g537(.A(new_n731), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n533), .A2(KEYINPUT110), .ZN(new_n740));
  NAND3_X1  g539(.A1(new_n726), .A2(new_n727), .A3(new_n528), .ZN(new_n741));
  NAND2_X1  g540(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  AOI21_X1  g541(.A(new_n739), .B1(new_n742), .B2(new_n521), .ZN(new_n743));
  AOI21_X1  g542(.A(new_n592), .B1(new_n521), .B2(new_n533), .ZN(new_n744));
  INV_X1    g543(.A(KEYINPUT44), .ZN(new_n745));
  NOR2_X1   g544(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  OAI211_X1 g545(.A(new_n738), .B(new_n735), .C1(new_n743), .C2(new_n746), .ZN(new_n747));
  NAND3_X1  g546(.A1(new_n737), .A2(new_n700), .A3(new_n747), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n748), .A2(G29gat), .ZN(new_n749));
  INV_X1    g548(.A(new_n700), .ZN(new_n750));
  NOR4_X1   g549(.A1(new_n733), .A2(G29gat), .A3(new_n750), .A4(new_n736), .ZN(new_n751));
  XOR2_X1   g550(.A(new_n751), .B(KEYINPUT45), .Z(new_n752));
  NAND2_X1  g551(.A1(new_n749), .A2(new_n752), .ZN(G1328gat));
  NAND3_X1  g552(.A1(new_n737), .A2(new_n704), .A3(new_n747), .ZN(new_n754));
  INV_X1    g553(.A(KEYINPUT112), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  NAND4_X1  g555(.A1(new_n737), .A2(KEYINPUT112), .A3(new_n704), .A4(new_n747), .ZN(new_n757));
  NAND3_X1  g556(.A1(new_n756), .A2(G36gat), .A3(new_n757), .ZN(new_n758));
  NOR4_X1   g557(.A1(new_n733), .A2(G36gat), .A3(new_n503), .A4(new_n736), .ZN(new_n759));
  XNOR2_X1  g558(.A(new_n759), .B(KEYINPUT46), .ZN(new_n760));
  NAND2_X1  g559(.A1(new_n758), .A2(new_n760), .ZN(G1329gat));
  NOR2_X1   g560(.A1(new_n734), .A2(new_n736), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n762), .A2(new_n714), .ZN(new_n763));
  NAND2_X1  g562(.A1(new_n763), .A2(G43gat), .ZN(new_n764));
  INV_X1    g563(.A(new_n522), .ZN(new_n765));
  NOR4_X1   g564(.A1(new_n733), .A2(G43gat), .A3(new_n765), .A4(new_n736), .ZN(new_n766));
  INV_X1    g565(.A(new_n766), .ZN(new_n767));
  NAND3_X1  g566(.A1(new_n764), .A2(KEYINPUT47), .A3(new_n767), .ZN(new_n768));
  NAND3_X1  g567(.A1(new_n737), .A2(new_n714), .A3(new_n747), .ZN(new_n769));
  AOI21_X1  g568(.A(new_n766), .B1(new_n769), .B2(G43gat), .ZN(new_n770));
  OAI21_X1  g569(.A(new_n768), .B1(new_n770), .B2(KEYINPUT47), .ZN(G1330gat));
  NAND4_X1  g570(.A1(new_n744), .A2(new_n331), .A3(new_n415), .A4(new_n735), .ZN(new_n772));
  INV_X1    g571(.A(new_n772), .ZN(new_n773));
  NAND3_X1  g572(.A1(new_n737), .A2(new_n415), .A3(new_n747), .ZN(new_n774));
  AOI21_X1  g573(.A(new_n773), .B1(new_n774), .B2(G50gat), .ZN(new_n775));
  XNOR2_X1  g574(.A(KEYINPUT113), .B(KEYINPUT48), .ZN(new_n776));
  AOI21_X1  g575(.A(new_n331), .B1(new_n762), .B2(new_n415), .ZN(new_n777));
  OR2_X1    g576(.A1(new_n773), .A2(KEYINPUT114), .ZN(new_n778));
  NAND2_X1  g577(.A1(new_n773), .A2(KEYINPUT114), .ZN(new_n779));
  NAND3_X1  g578(.A1(new_n778), .A2(KEYINPUT48), .A3(new_n779), .ZN(new_n780));
  OAI22_X1  g579(.A1(new_n775), .A2(new_n776), .B1(new_n777), .B2(new_n780), .ZN(G1331gat));
  INV_X1    g580(.A(new_n697), .ZN(new_n782));
  NOR3_X1   g581(.A1(new_n643), .A2(new_n672), .A3(new_n782), .ZN(new_n783));
  AND2_X1   g582(.A1(new_n730), .A2(new_n783), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n784), .A2(new_n700), .ZN(new_n785));
  XNOR2_X1  g584(.A(new_n785), .B(G57gat), .ZN(G1332gat));
  NOR2_X1   g585(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n787));
  AND2_X1   g586(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n788));
  OAI211_X1 g587(.A(new_n784), .B(new_n704), .C1(new_n787), .C2(new_n788), .ZN(new_n789));
  AND2_X1   g588(.A1(new_n784), .A2(new_n704), .ZN(new_n790));
  OAI21_X1  g589(.A(new_n789), .B1(new_n790), .B2(new_n787), .ZN(new_n791));
  XNOR2_X1  g590(.A(new_n791), .B(KEYINPUT115), .ZN(G1333gat));
  NAND2_X1  g591(.A1(new_n784), .A2(new_n714), .ZN(new_n793));
  NOR2_X1   g592(.A1(new_n765), .A2(G71gat), .ZN(new_n794));
  AOI22_X1  g593(.A1(new_n793), .A2(G71gat), .B1(new_n784), .B2(new_n794), .ZN(new_n795));
  XNOR2_X1  g594(.A(new_n795), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g595(.A1(new_n784), .A2(new_n415), .ZN(new_n797));
  XOR2_X1   g596(.A(KEYINPUT116), .B(G78gat), .Z(new_n798));
  XNOR2_X1  g597(.A(new_n797), .B(new_n798), .ZN(G1335gat));
  INV_X1    g598(.A(new_n642), .ZN(new_n800));
  NAND3_X1  g599(.A1(new_n673), .A2(new_n800), .A3(new_n697), .ZN(new_n801));
  XOR2_X1   g600(.A(new_n801), .B(KEYINPUT117), .Z(new_n802));
  OAI21_X1  g601(.A(new_n802), .B1(new_n743), .B2(new_n746), .ZN(new_n803));
  OAI21_X1  g602(.A(G85gat), .B1(new_n803), .B2(new_n750), .ZN(new_n804));
  NOR3_X1   g603(.A1(new_n672), .A2(new_n592), .A3(new_n642), .ZN(new_n805));
  AND3_X1   g604(.A1(new_n730), .A2(KEYINPUT51), .A3(new_n805), .ZN(new_n806));
  AOI21_X1  g605(.A(KEYINPUT51), .B1(new_n730), .B2(new_n805), .ZN(new_n807));
  NOR2_X1   g606(.A1(new_n806), .A2(new_n807), .ZN(new_n808));
  NAND3_X1  g607(.A1(new_n700), .A2(new_n575), .A3(new_n697), .ZN(new_n809));
  OAI21_X1  g608(.A(new_n804), .B1(new_n808), .B2(new_n809), .ZN(G1336gat));
  OAI21_X1  g609(.A(G92gat), .B1(new_n803), .B2(new_n503), .ZN(new_n811));
  NOR3_X1   g610(.A1(new_n782), .A2(new_n503), .A3(G92gat), .ZN(new_n812));
  XNOR2_X1  g611(.A(new_n812), .B(KEYINPUT119), .ZN(new_n813));
  INV_X1    g612(.A(new_n813), .ZN(new_n814));
  OAI21_X1  g613(.A(new_n814), .B1(new_n806), .B2(new_n807), .ZN(new_n815));
  NAND2_X1  g614(.A1(new_n811), .A2(new_n815), .ZN(new_n816));
  INV_X1    g615(.A(KEYINPUT52), .ZN(new_n817));
  INV_X1    g616(.A(KEYINPUT118), .ZN(new_n818));
  AOI21_X1  g617(.A(new_n817), .B1(new_n815), .B2(new_n818), .ZN(new_n819));
  XNOR2_X1  g618(.A(new_n816), .B(new_n819), .ZN(G1337gat));
  OAI21_X1  g619(.A(G99gat), .B1(new_n803), .B2(new_n329), .ZN(new_n821));
  INV_X1    g620(.A(G99gat), .ZN(new_n822));
  NAND3_X1  g621(.A1(new_n522), .A2(new_n822), .A3(new_n697), .ZN(new_n823));
  OAI21_X1  g622(.A(new_n821), .B1(new_n808), .B2(new_n823), .ZN(new_n824));
  INV_X1    g623(.A(KEYINPUT120), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n824), .A2(new_n825), .ZN(new_n826));
  OAI211_X1 g625(.A(new_n821), .B(KEYINPUT120), .C1(new_n808), .C2(new_n823), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n826), .A2(new_n827), .ZN(G1338gat));
  OAI21_X1  g627(.A(G106gat), .B1(new_n803), .B2(new_n414), .ZN(new_n829));
  OR3_X1    g628(.A1(new_n414), .A2(G106gat), .A3(new_n782), .ZN(new_n830));
  OAI21_X1  g629(.A(new_n829), .B1(new_n808), .B2(new_n830), .ZN(new_n831));
  XNOR2_X1  g630(.A(KEYINPUT121), .B(KEYINPUT53), .ZN(new_n832));
  INV_X1    g631(.A(new_n832), .ZN(new_n833));
  NAND2_X1  g632(.A1(new_n831), .A2(new_n833), .ZN(new_n834));
  OAI211_X1 g633(.A(new_n829), .B(new_n832), .C1(new_n808), .C2(new_n830), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n834), .A2(new_n835), .ZN(G1339gat));
  NOR3_X1   g635(.A1(new_n643), .A2(new_n672), .A3(new_n697), .ZN(new_n837));
  INV_X1    g636(.A(new_n696), .ZN(new_n838));
  OR3_X1    g637(.A1(new_n680), .A2(new_n674), .A3(new_n683), .ZN(new_n839));
  NAND4_X1  g638(.A1(new_n692), .A2(KEYINPUT54), .A3(new_n839), .A4(new_n694), .ZN(new_n840));
  INV_X1    g639(.A(new_n684), .ZN(new_n841));
  XOR2_X1   g640(.A(KEYINPUT122), .B(KEYINPUT54), .Z(new_n842));
  AOI21_X1  g641(.A(new_n690), .B1(new_n841), .B2(new_n842), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n840), .A2(new_n843), .ZN(new_n844));
  INV_X1    g643(.A(KEYINPUT55), .ZN(new_n845));
  AOI21_X1  g644(.A(new_n838), .B1(new_n844), .B2(new_n845), .ZN(new_n846));
  NAND3_X1  g645(.A1(new_n840), .A2(new_n843), .A3(KEYINPUT55), .ZN(new_n847));
  AND2_X1   g646(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  AOI21_X1  g647(.A(new_n647), .B1(new_n658), .B2(new_n644), .ZN(new_n849));
  AOI21_X1  g648(.A(new_n648), .B1(new_n646), .B2(new_n650), .ZN(new_n850));
  OAI21_X1  g649(.A(new_n665), .B1(new_n849), .B2(new_n850), .ZN(new_n851));
  AND2_X1   g650(.A1(new_n671), .A2(new_n851), .ZN(new_n852));
  NAND3_X1  g651(.A1(new_n848), .A2(new_n852), .A3(new_n732), .ZN(new_n853));
  AOI22_X1  g652(.A1(new_n672), .A2(new_n848), .B1(new_n852), .B2(new_n697), .ZN(new_n854));
  OAI21_X1  g653(.A(new_n853), .B1(new_n854), .B2(new_n732), .ZN(new_n855));
  AOI21_X1  g654(.A(new_n837), .B1(new_n855), .B2(new_n800), .ZN(new_n856));
  NOR2_X1   g655(.A1(new_n856), .A2(new_n415), .ZN(new_n857));
  NOR2_X1   g656(.A1(new_n750), .A2(new_n704), .ZN(new_n858));
  NAND3_X1  g657(.A1(new_n857), .A2(new_n522), .A3(new_n858), .ZN(new_n859));
  OAI21_X1  g658(.A(G113gat), .B1(new_n859), .B2(new_n673), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n720), .A2(new_n723), .ZN(new_n861));
  INV_X1    g660(.A(new_n858), .ZN(new_n862));
  NOR3_X1   g661(.A1(new_n856), .A2(new_n861), .A3(new_n862), .ZN(new_n863));
  NAND4_X1  g662(.A1(new_n863), .A2(new_n207), .A3(new_n209), .A4(new_n672), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n860), .A2(new_n864), .ZN(G1340gat));
  NOR3_X1   g664(.A1(new_n859), .A2(new_n223), .A3(new_n782), .ZN(new_n866));
  AOI21_X1  g665(.A(G120gat), .B1(new_n863), .B2(new_n697), .ZN(new_n867));
  NOR2_X1   g666(.A1(new_n866), .A2(new_n867), .ZN(G1341gat));
  OAI21_X1  g667(.A(G127gat), .B1(new_n859), .B2(new_n800), .ZN(new_n869));
  NAND3_X1  g668(.A1(new_n863), .A2(new_n217), .A3(new_n642), .ZN(new_n870));
  NAND2_X1  g669(.A1(new_n869), .A2(new_n870), .ZN(G1342gat));
  NAND3_X1  g670(.A1(new_n863), .A2(new_n219), .A3(new_n732), .ZN(new_n872));
  XOR2_X1   g671(.A(KEYINPUT123), .B(KEYINPUT56), .Z(new_n873));
  XNOR2_X1  g672(.A(new_n872), .B(new_n873), .ZN(new_n874));
  OAI21_X1  g673(.A(G134gat), .B1(new_n859), .B2(new_n592), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n874), .A2(new_n875), .ZN(G1343gat));
  NOR2_X1   g675(.A1(new_n714), .A2(new_n862), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n415), .A2(KEYINPUT57), .ZN(new_n878));
  INV_X1    g677(.A(new_n671), .ZN(new_n879));
  AOI21_X1  g678(.A(new_n666), .B1(new_n657), .B2(new_n659), .ZN(new_n880));
  OAI211_X1 g679(.A(new_n847), .B(new_n846), .C1(new_n879), .C2(new_n880), .ZN(new_n881));
  NAND3_X1  g680(.A1(new_n671), .A2(new_n697), .A3(new_n851), .ZN(new_n882));
  AOI21_X1  g681(.A(new_n732), .B1(new_n881), .B2(new_n882), .ZN(new_n883));
  INV_X1    g682(.A(KEYINPUT124), .ZN(new_n884));
  OAI21_X1  g683(.A(new_n853), .B1(new_n883), .B2(new_n884), .ZN(new_n885));
  NOR3_X1   g684(.A1(new_n854), .A2(KEYINPUT124), .A3(new_n732), .ZN(new_n886));
  OAI21_X1  g685(.A(new_n800), .B1(new_n885), .B2(new_n886), .ZN(new_n887));
  NAND4_X1  g686(.A1(new_n673), .A2(new_n642), .A3(new_n592), .A4(new_n782), .ZN(new_n888));
  AOI21_X1  g687(.A(new_n878), .B1(new_n887), .B2(new_n888), .ZN(new_n889));
  AND3_X1   g688(.A1(new_n848), .A2(new_n852), .A3(new_n732), .ZN(new_n890));
  OAI21_X1  g689(.A(new_n800), .B1(new_n883), .B2(new_n890), .ZN(new_n891));
  NAND2_X1  g690(.A1(new_n891), .A2(new_n888), .ZN(new_n892));
  AOI21_X1  g691(.A(KEYINPUT57), .B1(new_n892), .B2(new_n415), .ZN(new_n893));
  OAI21_X1  g692(.A(new_n877), .B1(new_n889), .B2(new_n893), .ZN(new_n894));
  OAI21_X1  g693(.A(G141gat), .B1(new_n894), .B2(new_n673), .ZN(new_n895));
  NOR3_X1   g694(.A1(new_n856), .A2(new_n414), .A3(new_n714), .ZN(new_n896));
  NAND2_X1  g695(.A1(new_n896), .A2(new_n858), .ZN(new_n897));
  NAND2_X1  g696(.A1(new_n672), .A2(new_n357), .ZN(new_n898));
  OAI21_X1  g697(.A(new_n895), .B1(new_n897), .B2(new_n898), .ZN(new_n899));
  NAND2_X1  g698(.A1(new_n899), .A2(KEYINPUT58), .ZN(new_n900));
  INV_X1    g699(.A(KEYINPUT58), .ZN(new_n901));
  OAI211_X1 g700(.A(new_n895), .B(new_n901), .C1(new_n897), .C2(new_n898), .ZN(new_n902));
  NAND2_X1  g701(.A1(new_n900), .A2(new_n902), .ZN(G1344gat));
  INV_X1    g702(.A(KEYINPUT57), .ZN(new_n904));
  AOI211_X1 g703(.A(new_n904), .B(new_n414), .C1(new_n891), .C2(new_n888), .ZN(new_n905));
  OAI211_X1 g704(.A(new_n697), .B(new_n877), .C1(new_n893), .C2(new_n905), .ZN(new_n906));
  INV_X1    g705(.A(KEYINPUT126), .ZN(new_n907));
  OAI21_X1  g706(.A(G148gat), .B1(new_n906), .B2(new_n907), .ZN(new_n908));
  OAI21_X1  g707(.A(new_n904), .B1(new_n856), .B2(new_n414), .ZN(new_n909));
  NAND3_X1  g708(.A1(new_n892), .A2(KEYINPUT57), .A3(new_n415), .ZN(new_n910));
  AOI21_X1  g709(.A(new_n782), .B1(new_n909), .B2(new_n910), .ZN(new_n911));
  AOI21_X1  g710(.A(KEYINPUT126), .B1(new_n911), .B2(new_n877), .ZN(new_n912));
  OAI21_X1  g711(.A(KEYINPUT59), .B1(new_n908), .B2(new_n912), .ZN(new_n913));
  NOR2_X1   g712(.A1(new_n359), .A2(KEYINPUT59), .ZN(new_n914));
  OAI21_X1  g713(.A(new_n914), .B1(new_n894), .B2(new_n782), .ZN(new_n915));
  NAND2_X1  g714(.A1(new_n913), .A2(new_n915), .ZN(new_n916));
  AND4_X1   g715(.A1(new_n359), .A2(new_n896), .A3(new_n697), .A4(new_n858), .ZN(new_n917));
  XOR2_X1   g716(.A(new_n917), .B(KEYINPUT125), .Z(new_n918));
  NAND2_X1  g717(.A1(new_n916), .A2(new_n918), .ZN(G1345gat));
  OAI21_X1  g718(.A(G155gat), .B1(new_n894), .B2(new_n800), .ZN(new_n920));
  NAND2_X1  g719(.A1(new_n642), .A2(new_n369), .ZN(new_n921));
  OAI21_X1  g720(.A(new_n920), .B1(new_n897), .B2(new_n921), .ZN(G1346gat));
  OAI21_X1  g721(.A(G162gat), .B1(new_n894), .B2(new_n592), .ZN(new_n923));
  NOR3_X1   g722(.A1(new_n592), .A2(new_n750), .A3(G162gat), .ZN(new_n924));
  NAND3_X1  g723(.A1(new_n896), .A2(new_n503), .A3(new_n924), .ZN(new_n925));
  NAND2_X1  g724(.A1(new_n923), .A2(new_n925), .ZN(G1347gat));
  NAND2_X1  g725(.A1(new_n750), .A2(new_n704), .ZN(new_n927));
  NOR2_X1   g726(.A1(new_n861), .A2(new_n927), .ZN(new_n928));
  NAND2_X1  g727(.A1(new_n892), .A2(new_n928), .ZN(new_n929));
  INV_X1    g728(.A(new_n929), .ZN(new_n930));
  AOI21_X1  g729(.A(G169gat), .B1(new_n930), .B2(new_n672), .ZN(new_n931));
  NOR2_X1   g730(.A1(new_n765), .A2(new_n927), .ZN(new_n932));
  NAND2_X1  g731(.A1(new_n857), .A2(new_n932), .ZN(new_n933));
  INV_X1    g732(.A(new_n933), .ZN(new_n934));
  NOR2_X1   g733(.A1(new_n673), .A2(new_n243), .ZN(new_n935));
  AOI21_X1  g734(.A(new_n931), .B1(new_n934), .B2(new_n935), .ZN(G1348gat));
  OAI21_X1  g735(.A(G176gat), .B1(new_n933), .B2(new_n782), .ZN(new_n937));
  NAND3_X1  g736(.A1(new_n930), .A2(new_n244), .A3(new_n697), .ZN(new_n938));
  NAND2_X1  g737(.A1(new_n937), .A2(new_n938), .ZN(G1349gat));
  OAI21_X1  g738(.A(G183gat), .B1(new_n933), .B2(new_n800), .ZN(new_n940));
  NAND2_X1  g739(.A1(new_n642), .A2(new_n268), .ZN(new_n941));
  OAI21_X1  g740(.A(new_n940), .B1(new_n929), .B2(new_n941), .ZN(new_n942));
  XNOR2_X1  g741(.A(new_n942), .B(KEYINPUT60), .ZN(G1350gat));
  NAND3_X1  g742(.A1(new_n930), .A2(new_n269), .A3(new_n732), .ZN(new_n944));
  OAI21_X1  g743(.A(G190gat), .B1(new_n933), .B2(new_n592), .ZN(new_n945));
  AND2_X1   g744(.A1(new_n945), .A2(KEYINPUT61), .ZN(new_n946));
  NOR2_X1   g745(.A1(new_n945), .A2(KEYINPUT61), .ZN(new_n947));
  OAI21_X1  g746(.A(new_n944), .B1(new_n946), .B2(new_n947), .ZN(G1351gat));
  NAND2_X1  g747(.A1(new_n909), .A2(new_n910), .ZN(new_n949));
  NOR2_X1   g748(.A1(new_n714), .A2(new_n927), .ZN(new_n950));
  NAND2_X1  g749(.A1(new_n949), .A2(new_n950), .ZN(new_n951));
  INV_X1    g750(.A(G197gat), .ZN(new_n952));
  NOR3_X1   g751(.A1(new_n951), .A2(new_n952), .A3(new_n673), .ZN(new_n953));
  NOR2_X1   g752(.A1(new_n856), .A2(new_n414), .ZN(new_n954));
  AND2_X1   g753(.A1(new_n954), .A2(new_n950), .ZN(new_n955));
  AOI21_X1  g754(.A(G197gat), .B1(new_n955), .B2(new_n672), .ZN(new_n956));
  NOR2_X1   g755(.A1(new_n953), .A2(new_n956), .ZN(G1352gat));
  INV_X1    g756(.A(G204gat), .ZN(new_n958));
  NAND4_X1  g757(.A1(new_n954), .A2(new_n958), .A3(new_n697), .A4(new_n950), .ZN(new_n959));
  XOR2_X1   g758(.A(new_n959), .B(KEYINPUT62), .Z(new_n960));
  AOI21_X1  g759(.A(new_n958), .B1(new_n911), .B2(new_n950), .ZN(new_n961));
  INV_X1    g760(.A(new_n961), .ZN(new_n962));
  NAND3_X1  g761(.A1(new_n960), .A2(KEYINPUT127), .A3(new_n962), .ZN(new_n963));
  INV_X1    g762(.A(KEYINPUT127), .ZN(new_n964));
  XNOR2_X1  g763(.A(new_n959), .B(KEYINPUT62), .ZN(new_n965));
  OAI21_X1  g764(.A(new_n964), .B1(new_n965), .B2(new_n961), .ZN(new_n966));
  NAND2_X1  g765(.A1(new_n963), .A2(new_n966), .ZN(G1353gat));
  NAND3_X1  g766(.A1(new_n955), .A2(new_n338), .A3(new_n642), .ZN(new_n968));
  NAND3_X1  g767(.A1(new_n949), .A2(new_n642), .A3(new_n950), .ZN(new_n969));
  AND3_X1   g768(.A1(new_n969), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n970));
  AOI21_X1  g769(.A(KEYINPUT63), .B1(new_n969), .B2(G211gat), .ZN(new_n971));
  OAI21_X1  g770(.A(new_n968), .B1(new_n970), .B2(new_n971), .ZN(G1354gat));
  OAI21_X1  g771(.A(G218gat), .B1(new_n951), .B2(new_n592), .ZN(new_n973));
  NAND3_X1  g772(.A1(new_n955), .A2(new_n339), .A3(new_n732), .ZN(new_n974));
  NAND2_X1  g773(.A1(new_n973), .A2(new_n974), .ZN(G1355gat));
endmodule


