

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n351, n352, n354, n355, n356, n357, n358, n359, n360, n361, n362,
         n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373,
         n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, n384,
         n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395,
         n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406,
         n407, n408, n409, n410, n411, n412, n413, n414, n415, n416, n417,
         n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, n428,
         n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, n439,
         n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450,
         n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461,
         n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472,
         n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483,
         n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494,
         n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505,
         n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516,
         n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527,
         n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538,
         n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549,
         n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560,
         n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571,
         n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582,
         n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593,
         n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604,
         n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615,
         n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n627,
         n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638,
         n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649,
         n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660,
         n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671,
         n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682,
         n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693,
         n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704,
         n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715,
         n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726,
         n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737,
         n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748,
         n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759,
         n760, n761, n762, n763, n764, n765, n766, n767, n768, n769, n770;

  AND2_X1 U373 ( .A1(n692), .A2(n689), .ZN(n716) );
  OR2_X1 U374 ( .A1(n557), .A2(n556), .ZN(n555) );
  NOR2_X1 U375 ( .A1(n596), .A2(n700), .ZN(n580) );
  OR2_X1 U376 ( .A1(n578), .A2(n697), .ZN(n586) );
  INV_X2 U377 ( .A(G953), .ZN(n765) );
  INV_X1 U378 ( .A(n351), .ZN(n452) );
  NAND2_X1 U379 ( .A1(n453), .A2(n688), .ZN(n351) );
  XNOR2_X2 U380 ( .A(n352), .B(n451), .ZN(n388) );
  NAND2_X1 U381 ( .A1(n625), .A2(n624), .ZN(n352) );
  XNOR2_X1 U382 ( .A(n490), .B(n523), .ZN(n495) );
  XNOR2_X2 U383 ( .A(n489), .B(n488), .ZN(n523) );
  XNOR2_X2 U384 ( .A(G113), .B(G122), .ZN(n397) );
  INV_X1 U385 ( .A(n586), .ZN(n702) );
  NOR2_X1 U386 ( .A1(n602), .A2(n601), .ZN(n694) );
  INV_X1 U387 ( .A(G146), .ZN(n653) );
  XNOR2_X2 U388 ( .A(n614), .B(KEYINPUT1), .ZN(n408) );
  XNOR2_X1 U389 ( .A(n371), .B(KEYINPUT90), .ZN(n566) );
  NAND2_X1 U390 ( .A1(n654), .A2(n647), .ZN(n371) );
  NOR2_X1 U391 ( .A1(n770), .A2(n651), .ZN(n623) );
  XNOR2_X1 U392 ( .A(n555), .B(KEYINPUT104), .ZN(n692) );
  XNOR2_X1 U393 ( .A(n396), .B(G119), .ZN(n536) );
  NOR2_X1 U394 ( .A1(n383), .A2(n648), .ZN(n382) );
  AND2_X1 U395 ( .A1(G217), .A2(n516), .ZN(n517) );
  XNOR2_X1 U396 ( .A(n397), .B(G104), .ZN(n479) );
  OR2_X2 U397 ( .A1(n611), .A2(n584), .ZN(n683) );
  XNOR2_X1 U398 ( .A(n539), .B(n538), .ZN(n661) );
  NOR2_X1 U399 ( .A1(G953), .A2(G237), .ZN(n531) );
  NAND2_X2 U400 ( .A1(n425), .A2(n422), .ZN(n553) );
  NAND2_X1 U401 ( .A1(n424), .A2(n423), .ZN(n422) );
  AND2_X1 U402 ( .A1(n427), .A2(n426), .ZN(n425) );
  NOR2_X1 U403 ( .A1(n471), .A2(n359), .ZN(n423) );
  INV_X1 U404 ( .A(KEYINPUT44), .ZN(n414) );
  AND2_X1 U405 ( .A1(n691), .A2(n679), .ZN(n558) );
  XOR2_X1 U406 ( .A(KEYINPUT100), .B(KEYINPUT101), .Z(n475) );
  XNOR2_X1 U407 ( .A(n632), .B(n392), .ZN(n712) );
  INV_X1 U408 ( .A(KEYINPUT38), .ZN(n392) );
  INV_X1 U409 ( .A(KEYINPUT48), .ZN(n451) );
  XNOR2_X1 U410 ( .A(n523), .B(n448), .ZN(n760) );
  XNOR2_X1 U411 ( .A(n521), .B(n522), .ZN(n448) );
  XNOR2_X1 U412 ( .A(n431), .B(KEYINPUT17), .ZN(n430) );
  XNOR2_X1 U413 ( .A(KEYINPUT4), .B(KEYINPUT18), .ZN(n431) );
  XNOR2_X1 U414 ( .A(KEYINPUT75), .B(KEYINPUT91), .ZN(n429) );
  NAND2_X1 U415 ( .A1(n712), .A2(n711), .ZN(n715) );
  OR2_X1 U416 ( .A1(n661), .A2(n440), .ZN(n439) );
  AND2_X1 U417 ( .A1(n380), .A2(n444), .ZN(n443) );
  NAND2_X1 U418 ( .A1(n442), .A2(n441), .ZN(n440) );
  XNOR2_X1 U419 ( .A(n393), .B(n464), .ZN(n587) );
  XNOR2_X1 U420 ( .A(n463), .B(KEYINPUT93), .ZN(n464) );
  XNOR2_X1 U421 ( .A(G116), .B(G113), .ZN(n532) );
  XNOR2_X1 U422 ( .A(n421), .B(n459), .ZN(n752) );
  XNOR2_X1 U423 ( .A(n479), .B(n536), .ZN(n421) );
  XNOR2_X1 U424 ( .A(KEYINPUT16), .B(G110), .ZN(n458) );
  XNOR2_X1 U425 ( .A(n760), .B(n653), .ZN(n539) );
  INV_X1 U426 ( .A(KEYINPUT32), .ZN(n405) );
  NAND2_X1 U427 ( .A1(n553), .A2(n500), .ZN(n503) );
  BUF_X1 U428 ( .A(n545), .Z(n628) );
  NAND2_X1 U429 ( .A1(n667), .A2(G475), .ZN(n370) );
  BUF_X1 U430 ( .A(n667), .Z(n670) );
  XNOR2_X1 U431 ( .A(n694), .B(n377), .ZN(n604) );
  INV_X1 U432 ( .A(KEYINPUT85), .ZN(n377) );
  NOR2_X1 U433 ( .A1(n683), .A2(n394), .ZN(n603) );
  NAND2_X1 U434 ( .A1(n456), .A2(n395), .ZN(n394) );
  INV_X1 U435 ( .A(KEYINPUT47), .ZN(n395) );
  INV_X1 U436 ( .A(n716), .ZN(n456) );
  AND2_X1 U437 ( .A1(n563), .A2(n413), .ZN(n412) );
  INV_X1 U438 ( .A(KEYINPUT88), .ZN(n564) );
  XNOR2_X1 U439 ( .A(KEYINPUT20), .B(n497), .ZN(n516) );
  INV_X1 U440 ( .A(n540), .ZN(n442) );
  NAND2_X1 U441 ( .A1(n540), .A2(G902), .ZN(n444) );
  NOR2_X1 U442 ( .A1(n650), .A2(n386), .ZN(n385) );
  INV_X1 U443 ( .A(KEYINPUT83), .ZN(n386) );
  XNOR2_X1 U444 ( .A(KEYINPUT77), .B(KEYINPUT8), .ZN(n486) );
  XNOR2_X1 U445 ( .A(G116), .B(G107), .ZN(n491) );
  XNOR2_X1 U446 ( .A(n476), .B(n457), .ZN(n477) );
  XNOR2_X1 U447 ( .A(n475), .B(n474), .ZN(n476) );
  XNOR2_X1 U448 ( .A(G143), .B(KEYINPUT11), .ZN(n474) );
  NAND2_X1 U449 ( .A1(n354), .A2(n637), .ZN(n449) );
  AND2_X1 U450 ( .A1(n545), .A2(n702), .ZN(n378) );
  NAND2_X1 U451 ( .A1(G237), .A2(G234), .ZN(n467) );
  XOR2_X1 U452 ( .A(KEYINPUT71), .B(KEYINPUT14), .Z(n468) );
  NAND2_X1 U453 ( .A1(n471), .A2(n359), .ZN(n426) );
  BUF_X1 U454 ( .A(n700), .Z(n379) );
  XNOR2_X1 U455 ( .A(n700), .B(KEYINPUT6), .ZN(n545) );
  BUF_X1 U456 ( .A(n737), .Z(n747) );
  XNOR2_X1 U457 ( .A(G128), .B(G119), .ZN(n510) );
  XNOR2_X1 U458 ( .A(n505), .B(KEYINPUT74), .ZN(n506) );
  INV_X1 U459 ( .A(KEYINPUT96), .ZN(n505) );
  INV_X1 U460 ( .A(G134), .ZN(n488) );
  XNOR2_X1 U461 ( .A(G107), .B(G101), .ZN(n524) );
  XNOR2_X1 U462 ( .A(n752), .B(n419), .ZN(n657) );
  XNOR2_X1 U463 ( .A(n430), .B(n429), .ZN(n462) );
  BUF_X1 U464 ( .A(n587), .Z(n632) );
  XNOR2_X1 U465 ( .A(n610), .B(n609), .ZN(n732) );
  XNOR2_X1 U466 ( .A(n608), .B(KEYINPUT41), .ZN(n609) );
  NOR2_X1 U467 ( .A1(n715), .A2(n714), .ZN(n610) );
  OR2_X1 U468 ( .A1(n596), .A2(n391), .ZN(n627) );
  XNOR2_X1 U469 ( .A(n390), .B(n389), .ZN(n618) );
  INV_X1 U470 ( .A(KEYINPUT30), .ZN(n389) );
  OR2_X1 U471 ( .A1(n700), .A2(n391), .ZN(n390) );
  NAND2_X1 U472 ( .A1(n587), .A2(n711), .ZN(n416) );
  XNOR2_X1 U473 ( .A(n583), .B(KEYINPUT108), .ZN(n611) );
  XNOR2_X1 U474 ( .A(n485), .B(n484), .ZN(n557) );
  INV_X1 U475 ( .A(n379), .ZN(n590) );
  BUF_X1 U476 ( .A(n408), .Z(n406) );
  XNOR2_X1 U477 ( .A(KEYINPUT98), .B(KEYINPUT5), .ZN(n534) );
  AND2_X1 U478 ( .A1(n541), .A2(n358), .ZN(n404) );
  XOR2_X1 U479 ( .A(KEYINPUT31), .B(n550), .Z(n691) );
  XNOR2_X1 U480 ( .A(n374), .B(n373), .ZN(n669) );
  NAND2_X1 U481 ( .A1(n670), .A2(G217), .ZN(n374) );
  INV_X1 U482 ( .A(KEYINPUT60), .ZN(n367) );
  XNOR2_X1 U483 ( .A(n370), .B(n363), .ZN(n369) );
  NAND2_X1 U484 ( .A1(n641), .A2(n640), .ZN(n354) );
  INV_X1 U485 ( .A(n650), .ZN(n450) );
  OR2_X1 U486 ( .A1(G902), .A2(G237), .ZN(n355) );
  NAND2_X1 U487 ( .A1(n465), .A2(G214), .ZN(n711) );
  INV_X1 U488 ( .A(n711), .ZN(n391) );
  AND2_X1 U489 ( .A1(n541), .A2(n696), .ZN(n356) );
  XOR2_X1 U490 ( .A(KEYINPUT24), .B(KEYINPUT94), .Z(n357) );
  AND2_X1 U491 ( .A1(n696), .A2(n405), .ZN(n358) );
  INV_X1 U492 ( .A(G902), .ZN(n441) );
  XNOR2_X1 U493 ( .A(KEYINPUT65), .B(KEYINPUT0), .ZN(n359) );
  XNOR2_X1 U494 ( .A(KEYINPUT82), .B(KEYINPUT35), .ZN(n360) );
  XOR2_X1 U495 ( .A(KEYINPUT107), .B(KEYINPUT28), .Z(n361) );
  XOR2_X1 U496 ( .A(n657), .B(n656), .Z(n362) );
  XOR2_X1 U497 ( .A(n655), .B(KEYINPUT59), .Z(n363) );
  INV_X1 U498 ( .A(KEYINPUT79), .ZN(n436) );
  NAND2_X1 U499 ( .A1(n548), .A2(KEYINPUT44), .ZN(n364) );
  AND2_X1 U500 ( .A1(n354), .A2(n436), .ZN(n365) );
  NOR2_X1 U501 ( .A1(n765), .A2(G952), .ZN(n675) );
  XOR2_X1 U502 ( .A(KEYINPUT84), .B(KEYINPUT56), .Z(n366) );
  XNOR2_X1 U503 ( .A(n368), .B(n367), .ZN(G60) );
  NAND2_X1 U504 ( .A1(n369), .A2(n664), .ZN(n368) );
  XNOR2_X1 U505 ( .A(n372), .B(KEYINPUT87), .ZN(n418) );
  NAND2_X1 U506 ( .A1(n438), .A2(n428), .ZN(n372) );
  INV_X1 U507 ( .A(n668), .ZN(n373) );
  XNOR2_X1 U508 ( .A(n375), .B(n366), .ZN(G51) );
  NAND2_X1 U509 ( .A1(n376), .A2(n664), .ZN(n375) );
  NAND2_X1 U510 ( .A1(n403), .A2(n402), .ZN(n654) );
  NAND2_X1 U511 ( .A1(n388), .A2(n385), .ZN(n384) );
  NAND2_X1 U512 ( .A1(n384), .A2(n382), .ZN(n381) );
  XNOR2_X1 U513 ( .A(n658), .B(n362), .ZN(n376) );
  AND2_X2 U514 ( .A1(n761), .A2(n365), .ZN(n399) );
  NAND2_X1 U515 ( .A1(n434), .A2(n449), .ZN(n433) );
  NOR2_X4 U516 ( .A1(n381), .A2(n387), .ZN(n761) );
  NAND2_X1 U517 ( .A1(n378), .A2(n408), .ZN(n546) );
  NAND2_X1 U518 ( .A1(n661), .A2(n540), .ZN(n380) );
  AND2_X1 U519 ( .A1(n400), .A2(KEYINPUT79), .ZN(n435) );
  NAND2_X1 U520 ( .A1(n418), .A2(n570), .ZN(n417) );
  NOR2_X1 U521 ( .A1(n450), .A2(KEYINPUT83), .ZN(n383) );
  NOR2_X2 U522 ( .A1(n388), .A2(KEYINPUT83), .ZN(n387) );
  NAND2_X1 U523 ( .A1(n591), .A2(n618), .ZN(n592) );
  INV_X1 U524 ( .A(n712), .ZN(n616) );
  NAND2_X1 U525 ( .A1(n657), .A2(n641), .ZN(n393) );
  XNOR2_X2 U526 ( .A(G101), .B(KEYINPUT3), .ZN(n396) );
  NAND2_X1 U527 ( .A1(n398), .A2(n737), .ZN(n437) );
  AND2_X2 U528 ( .A1(n761), .A2(KEYINPUT2), .ZN(n398) );
  NAND2_X1 U529 ( .A1(n737), .A2(n761), .ZN(n400) );
  NAND2_X1 U530 ( .A1(n399), .A2(n737), .ZN(n434) );
  NAND2_X1 U531 ( .A1(n401), .A2(KEYINPUT32), .ZN(n403) );
  NAND2_X1 U532 ( .A1(n356), .A2(n561), .ZN(n401) );
  NAND2_X1 U533 ( .A1(n404), .A2(n561), .ZN(n402) );
  AND2_X1 U534 ( .A1(n561), .A2(n696), .ZN(n543) );
  XNOR2_X1 U535 ( .A(n758), .B(n477), .ZN(n481) );
  NAND2_X1 U536 ( .A1(n716), .A2(KEYINPUT47), .ZN(n453) );
  NOR2_X1 U537 ( .A1(n406), .A2(n590), .ZN(n542) );
  NOR2_X1 U538 ( .A1(n702), .A2(n406), .ZN(n704) );
  AND2_X1 U539 ( .A1(n549), .A2(n408), .ZN(n707) );
  XNOR2_X1 U540 ( .A(n408), .B(n407), .ZN(n601) );
  INV_X1 U541 ( .A(KEYINPUT92), .ZN(n407) );
  NOR2_X1 U542 ( .A1(n559), .A2(n406), .ZN(n560) );
  NOR2_X1 U543 ( .A1(n630), .A2(n406), .ZN(n631) );
  NAND2_X1 U544 ( .A1(n410), .A2(n409), .ZN(n415) );
  NAND2_X1 U545 ( .A1(n567), .A2(n364), .ZN(n409) );
  NAND2_X1 U546 ( .A1(n411), .A2(n548), .ZN(n410) );
  INV_X1 U547 ( .A(n567), .ZN(n411) );
  NAND2_X1 U548 ( .A1(n415), .A2(n412), .ZN(n565) );
  NAND2_X1 U549 ( .A1(KEYINPUT89), .A2(n414), .ZN(n413) );
  XNOR2_X2 U550 ( .A(n445), .B(n360), .ZN(n567) );
  XNOR2_X2 U551 ( .A(n416), .B(n466), .ZN(n584) );
  XNOR2_X2 U552 ( .A(n417), .B(n571), .ZN(n737) );
  XNOR2_X1 U553 ( .A(n420), .B(n462), .ZN(n419) );
  XNOR2_X1 U554 ( .A(n461), .B(n473), .ZN(n420) );
  INV_X1 U555 ( .A(n584), .ZN(n424) );
  NAND2_X1 U556 ( .A1(n584), .A2(n359), .ZN(n427) );
  XNOR2_X1 U557 ( .A(n544), .B(KEYINPUT64), .ZN(n428) );
  NOR2_X4 U558 ( .A1(n741), .A2(n432), .ZN(n667) );
  NOR2_X2 U559 ( .A1(n435), .A2(n433), .ZN(n432) );
  XNOR2_X2 U560 ( .A(n437), .B(KEYINPUT73), .ZN(n741) );
  XNOR2_X1 U561 ( .A(n565), .B(n564), .ZN(n438) );
  NAND2_X4 U562 ( .A1(n443), .A2(n439), .ZN(n700) );
  NAND2_X1 U563 ( .A1(n446), .A2(n593), .ZN(n445) );
  XNOR2_X1 U564 ( .A(n547), .B(n447), .ZN(n446) );
  INV_X1 U565 ( .A(KEYINPUT34), .ZN(n447) );
  XNOR2_X2 U566 ( .A(KEYINPUT66), .B(G131), .ZN(n522) );
  XNOR2_X2 U567 ( .A(G143), .B(G128), .ZN(n489) );
  NAND2_X1 U568 ( .A1(n455), .A2(n452), .ZN(n454) );
  XNOR2_X1 U569 ( .A(n454), .B(n595), .ZN(n606) );
  NAND2_X1 U570 ( .A1(n683), .A2(KEYINPUT47), .ZN(n455) );
  XNOR2_X1 U571 ( .A(n507), .B(n506), .ZN(n508) );
  XNOR2_X2 U572 ( .A(G902), .B(KEYINPUT15), .ZN(n641) );
  AND2_X1 U573 ( .A1(n531), .A2(G214), .ZN(n457) );
  INV_X1 U574 ( .A(KEYINPUT89), .ZN(n548) );
  XNOR2_X1 U575 ( .A(G140), .B(KEYINPUT10), .ZN(n472) );
  INV_X1 U576 ( .A(KEYINPUT109), .ZN(n608) );
  INV_X1 U577 ( .A(KEYINPUT122), .ZN(n645) );
  BUF_X1 U578 ( .A(n567), .Z(n659) );
  XNOR2_X1 U579 ( .A(n491), .B(n458), .ZN(n459) );
  XNOR2_X2 U580 ( .A(n653), .B(G125), .ZN(n473) );
  NAND2_X1 U581 ( .A1(G224), .A2(n765), .ZN(n460) );
  XNOR2_X1 U582 ( .A(n489), .B(n460), .ZN(n461) );
  XNOR2_X1 U583 ( .A(KEYINPUT72), .B(n355), .ZN(n465) );
  NAND2_X1 U584 ( .A1(n465), .A2(G210), .ZN(n463) );
  INV_X1 U585 ( .A(KEYINPUT19), .ZN(n466) );
  XNOR2_X1 U586 ( .A(n468), .B(n467), .ZN(n727) );
  NOR2_X1 U587 ( .A1(G898), .A2(n765), .ZN(n753) );
  NAND2_X1 U588 ( .A1(n753), .A2(G902), .ZN(n469) );
  NAND2_X1 U589 ( .A1(G952), .A2(n765), .ZN(n574) );
  NAND2_X1 U590 ( .A1(n469), .A2(n574), .ZN(n470) );
  NAND2_X1 U591 ( .A1(n727), .A2(n470), .ZN(n471) );
  XNOR2_X2 U592 ( .A(n473), .B(n472), .ZN(n758) );
  XNOR2_X1 U593 ( .A(n522), .B(KEYINPUT12), .ZN(n478) );
  XNOR2_X1 U594 ( .A(n479), .B(n478), .ZN(n480) );
  XNOR2_X1 U595 ( .A(n481), .B(n480), .ZN(n655) );
  NAND2_X1 U596 ( .A1(n655), .A2(n441), .ZN(n485) );
  XOR2_X1 U597 ( .A(KEYINPUT103), .B(KEYINPUT13), .Z(n483) );
  XNOR2_X1 U598 ( .A(KEYINPUT102), .B(G475), .ZN(n482) );
  XOR2_X1 U599 ( .A(n483), .B(n482), .Z(n484) );
  NAND2_X1 U600 ( .A1(n765), .A2(G234), .ZN(n487) );
  XNOR2_X1 U601 ( .A(n487), .B(n486), .ZN(n509) );
  NAND2_X1 U602 ( .A1(n509), .A2(G217), .ZN(n490) );
  XNOR2_X1 U603 ( .A(KEYINPUT9), .B(n491), .ZN(n493) );
  XNOR2_X1 U604 ( .A(G122), .B(KEYINPUT7), .ZN(n492) );
  XNOR2_X1 U605 ( .A(n493), .B(n492), .ZN(n494) );
  XNOR2_X1 U606 ( .A(n495), .B(n494), .ZN(n642) );
  NAND2_X1 U607 ( .A1(n642), .A2(n441), .ZN(n496) );
  XNOR2_X1 U608 ( .A(n496), .B(G478), .ZN(n554) );
  OR2_X1 U609 ( .A1(n557), .A2(n554), .ZN(n714) );
  NAND2_X1 U610 ( .A1(G234), .A2(n641), .ZN(n497) );
  AND2_X1 U611 ( .A1(n516), .A2(G221), .ZN(n499) );
  INV_X1 U612 ( .A(KEYINPUT21), .ZN(n498) );
  XNOR2_X1 U613 ( .A(n499), .B(n498), .ZN(n697) );
  NOR2_X1 U614 ( .A1(n714), .A2(n697), .ZN(n500) );
  INV_X1 U615 ( .A(KEYINPUT70), .ZN(n501) );
  XNOR2_X1 U616 ( .A(n501), .B(KEYINPUT22), .ZN(n502) );
  XNOR2_X2 U617 ( .A(n503), .B(n502), .ZN(n561) );
  XNOR2_X1 U618 ( .A(KEYINPUT23), .B(KEYINPUT95), .ZN(n504) );
  XNOR2_X1 U619 ( .A(n357), .B(n504), .ZN(n507) );
  XNOR2_X1 U620 ( .A(n508), .B(n758), .ZN(n515) );
  NAND2_X1 U621 ( .A1(n509), .A2(G221), .ZN(n513) );
  XOR2_X1 U622 ( .A(G137), .B(G110), .Z(n511) );
  XNOR2_X1 U623 ( .A(n511), .B(n510), .ZN(n512) );
  XNOR2_X1 U624 ( .A(n513), .B(n512), .ZN(n514) );
  XNOR2_X1 U625 ( .A(n515), .B(n514), .ZN(n668) );
  NAND2_X1 U626 ( .A1(n668), .A2(n441), .ZN(n520) );
  XNOR2_X1 U627 ( .A(KEYINPUT97), .B(n517), .ZN(n518) );
  XNOR2_X1 U628 ( .A(n518), .B(KEYINPUT25), .ZN(n519) );
  XNOR2_X2 U629 ( .A(n520), .B(n519), .ZN(n578) );
  BUF_X1 U630 ( .A(n578), .Z(n696) );
  XNOR2_X1 U631 ( .A(KEYINPUT4), .B(G137), .ZN(n521) );
  XOR2_X1 U632 ( .A(G140), .B(G110), .Z(n525) );
  XNOR2_X1 U633 ( .A(n525), .B(n524), .ZN(n526) );
  XOR2_X1 U634 ( .A(G104), .B(n526), .Z(n528) );
  NAND2_X1 U635 ( .A1(G227), .A2(n765), .ZN(n527) );
  XNOR2_X1 U636 ( .A(n528), .B(n527), .ZN(n529) );
  XNOR2_X1 U637 ( .A(n539), .B(n529), .ZN(n672) );
  NAND2_X1 U638 ( .A1(n672), .A2(n441), .ZN(n530) );
  XNOR2_X2 U639 ( .A(n530), .B(G469), .ZN(n614) );
  NAND2_X1 U640 ( .A1(n531), .A2(G210), .ZN(n533) );
  XNOR2_X1 U641 ( .A(n533), .B(n532), .ZN(n535) );
  XNOR2_X1 U642 ( .A(n535), .B(n534), .ZN(n537) );
  XNOR2_X1 U643 ( .A(n536), .B(n537), .ZN(n538) );
  XNOR2_X1 U644 ( .A(G472), .B(KEYINPUT99), .ZN(n540) );
  NOR2_X1 U645 ( .A1(n601), .A2(n628), .ZN(n541) );
  NAND2_X1 U646 ( .A1(n543), .A2(n542), .ZN(n647) );
  NAND2_X1 U647 ( .A1(n566), .A2(KEYINPUT44), .ZN(n544) );
  XNOR2_X2 U648 ( .A(n546), .B(KEYINPUT33), .ZN(n719) );
  NAND2_X1 U649 ( .A1(n719), .A2(n553), .ZN(n547) );
  AND2_X1 U650 ( .A1(n557), .A2(n554), .ZN(n593) );
  NOR2_X1 U651 ( .A1(n586), .A2(n379), .ZN(n549) );
  NAND2_X1 U652 ( .A1(n553), .A2(n707), .ZN(n550) );
  NAND2_X1 U653 ( .A1(n702), .A2(n614), .ZN(n551) );
  NOR2_X1 U654 ( .A1(n551), .A2(n590), .ZN(n552) );
  NAND2_X1 U655 ( .A1(n553), .A2(n552), .ZN(n679) );
  INV_X1 U656 ( .A(n554), .ZN(n556) );
  NAND2_X1 U657 ( .A1(n557), .A2(n556), .ZN(n689) );
  NOR2_X1 U658 ( .A1(n558), .A2(n716), .ZN(n562) );
  OR2_X1 U659 ( .A1(n628), .A2(n696), .ZN(n559) );
  AND2_X1 U660 ( .A1(n561), .A2(n560), .ZN(n677) );
  NOR2_X1 U661 ( .A1(n562), .A2(n677), .ZN(n563) );
  INV_X1 U662 ( .A(n566), .ZN(n569) );
  NOR2_X1 U663 ( .A1(n659), .A2(KEYINPUT44), .ZN(n568) );
  NAND2_X1 U664 ( .A1(n569), .A2(n568), .ZN(n570) );
  XOR2_X1 U665 ( .A(KEYINPUT81), .B(KEYINPUT45), .Z(n571) );
  NOR2_X1 U666 ( .A1(G900), .A2(n765), .ZN(n572) );
  NAND2_X1 U667 ( .A1(G902), .A2(n572), .ZN(n573) );
  NAND2_X1 U668 ( .A1(n574), .A2(n573), .ZN(n575) );
  NAND2_X1 U669 ( .A1(n727), .A2(n575), .ZN(n585) );
  NOR2_X1 U670 ( .A1(n697), .A2(n585), .ZN(n576) );
  XOR2_X1 U671 ( .A(n576), .B(KEYINPUT69), .Z(n577) );
  NAND2_X1 U672 ( .A1(n578), .A2(n577), .ZN(n579) );
  XNOR2_X1 U673 ( .A(n579), .B(KEYINPUT68), .ZN(n596) );
  XNOR2_X1 U674 ( .A(n580), .B(n361), .ZN(n582) );
  XNOR2_X1 U675 ( .A(n614), .B(KEYINPUT106), .ZN(n581) );
  NAND2_X1 U676 ( .A1(n582), .A2(n581), .ZN(n583) );
  NOR2_X1 U677 ( .A1(n586), .A2(n585), .ZN(n615) );
  NAND2_X1 U678 ( .A1(n615), .A2(n632), .ZN(n589) );
  INV_X1 U679 ( .A(n614), .ZN(n588) );
  NOR2_X1 U680 ( .A1(n589), .A2(n588), .ZN(n591) );
  XNOR2_X1 U681 ( .A(n592), .B(KEYINPUT105), .ZN(n594) );
  NAND2_X1 U682 ( .A1(n594), .A2(n593), .ZN(n688) );
  INV_X1 U683 ( .A(KEYINPUT76), .ZN(n595) );
  INV_X1 U684 ( .A(n689), .ZN(n597) );
  NAND2_X1 U685 ( .A1(n597), .A2(n632), .ZN(n598) );
  NOR2_X1 U686 ( .A1(n627), .A2(n598), .ZN(n599) );
  NAND2_X1 U687 ( .A1(n599), .A2(n628), .ZN(n600) );
  XNOR2_X1 U688 ( .A(n600), .B(KEYINPUT36), .ZN(n602) );
  NOR2_X1 U689 ( .A1(n604), .A2(n603), .ZN(n605) );
  NAND2_X1 U690 ( .A1(n606), .A2(n605), .ZN(n607) );
  XNOR2_X1 U691 ( .A(n607), .B(KEYINPUT67), .ZN(n625) );
  NOR2_X1 U692 ( .A1(n732), .A2(n611), .ZN(n613) );
  XNOR2_X1 U693 ( .A(KEYINPUT110), .B(KEYINPUT42), .ZN(n612) );
  XNOR2_X1 U694 ( .A(n613), .B(n612), .ZN(n770) );
  NAND2_X1 U695 ( .A1(n615), .A2(n614), .ZN(n617) );
  NOR2_X1 U696 ( .A1(n617), .A2(n616), .ZN(n619) );
  NAND2_X1 U697 ( .A1(n619), .A2(n618), .ZN(n621) );
  XOR2_X1 U698 ( .A(KEYINPUT86), .B(KEYINPUT39), .Z(n620) );
  XNOR2_X1 U699 ( .A(n621), .B(n620), .ZN(n634) );
  NOR2_X1 U700 ( .A1(n634), .A2(n689), .ZN(n622) );
  XNOR2_X1 U701 ( .A(n622), .B(KEYINPUT40), .ZN(n651) );
  XNOR2_X1 U702 ( .A(n623), .B(KEYINPUT46), .ZN(n624) );
  NOR2_X1 U703 ( .A1(n627), .A2(n689), .ZN(n629) );
  NAND2_X1 U704 ( .A1(n629), .A2(n628), .ZN(n630) );
  XNOR2_X1 U705 ( .A(n631), .B(KEYINPUT43), .ZN(n633) );
  NOR2_X1 U706 ( .A1(n633), .A2(n632), .ZN(n650) );
  NOR2_X1 U707 ( .A1(n634), .A2(n692), .ZN(n648) );
  INV_X1 U708 ( .A(n641), .ZN(n636) );
  NAND2_X1 U709 ( .A1(KEYINPUT2), .A2(KEYINPUT80), .ZN(n635) );
  NAND2_X1 U710 ( .A1(n636), .A2(n635), .ZN(n637) );
  INV_X1 U711 ( .A(KEYINPUT2), .ZN(n638) );
  NOR2_X1 U712 ( .A1(n638), .A2(KEYINPUT80), .ZN(n639) );
  NOR2_X1 U713 ( .A1(n639), .A2(KEYINPUT79), .ZN(n640) );
  NAND2_X1 U714 ( .A1(n667), .A2(G478), .ZN(n643) );
  XNOR2_X1 U715 ( .A(n643), .B(n642), .ZN(n644) );
  INV_X1 U716 ( .A(n675), .ZN(n664) );
  NAND2_X1 U717 ( .A1(n644), .A2(n664), .ZN(n646) );
  XNOR2_X1 U718 ( .A(n646), .B(n645), .ZN(G63) );
  XNOR2_X1 U719 ( .A(n647), .B(G110), .ZN(G12) );
  XNOR2_X1 U720 ( .A(G134), .B(KEYINPUT114), .ZN(n649) );
  XOR2_X1 U721 ( .A(n649), .B(n648), .Z(G36) );
  XOR2_X1 U722 ( .A(G140), .B(n650), .Z(G42) );
  XOR2_X1 U723 ( .A(n651), .B(G131), .Z(G33) );
  NOR2_X1 U724 ( .A1(n683), .A2(n689), .ZN(n652) );
  XNOR2_X1 U725 ( .A(n653), .B(n652), .ZN(G48) );
  XNOR2_X1 U726 ( .A(n654), .B(G119), .ZN(G21) );
  NAND2_X1 U727 ( .A1(n667), .A2(G210), .ZN(n658) );
  XNOR2_X1 U728 ( .A(KEYINPUT54), .B(KEYINPUT55), .ZN(n656) );
  XOR2_X1 U729 ( .A(n659), .B(G122), .Z(G24) );
  NAND2_X1 U730 ( .A1(n667), .A2(G472), .ZN(n663) );
  XNOR2_X1 U731 ( .A(KEYINPUT111), .B(KEYINPUT62), .ZN(n660) );
  XNOR2_X1 U732 ( .A(n661), .B(n660), .ZN(n662) );
  XNOR2_X1 U733 ( .A(n663), .B(n662), .ZN(n665) );
  NAND2_X1 U734 ( .A1(n665), .A2(n664), .ZN(n666) );
  XNOR2_X1 U735 ( .A(n666), .B(KEYINPUT63), .ZN(G57) );
  NOR2_X1 U736 ( .A1(n669), .A2(n675), .ZN(G66) );
  NAND2_X1 U737 ( .A1(n670), .A2(G469), .ZN(n674) );
  XNOR2_X1 U738 ( .A(KEYINPUT57), .B(KEYINPUT58), .ZN(n671) );
  XNOR2_X1 U739 ( .A(n672), .B(n671), .ZN(n673) );
  XNOR2_X1 U740 ( .A(n674), .B(n673), .ZN(n676) );
  NOR2_X1 U741 ( .A1(n676), .A2(n675), .ZN(G54) );
  XOR2_X1 U742 ( .A(G101), .B(n677), .Z(G3) );
  NOR2_X1 U743 ( .A1(n689), .A2(n679), .ZN(n678) );
  XOR2_X1 U744 ( .A(G104), .B(n678), .Z(G6) );
  NOR2_X1 U745 ( .A1(n692), .A2(n679), .ZN(n681) );
  XNOR2_X1 U746 ( .A(KEYINPUT27), .B(KEYINPUT26), .ZN(n680) );
  XNOR2_X1 U747 ( .A(n681), .B(n680), .ZN(n682) );
  XNOR2_X1 U748 ( .A(G107), .B(n682), .ZN(G9) );
  XOR2_X1 U749 ( .A(KEYINPUT112), .B(KEYINPUT29), .Z(n685) );
  NOR2_X1 U750 ( .A1(n683), .A2(n692), .ZN(n684) );
  XOR2_X1 U751 ( .A(n685), .B(n684), .Z(n686) );
  XNOR2_X1 U752 ( .A(G128), .B(n686), .ZN(G30) );
  XOR2_X1 U753 ( .A(G143), .B(KEYINPUT113), .Z(n687) );
  XNOR2_X1 U754 ( .A(n688), .B(n687), .ZN(G45) );
  NOR2_X1 U755 ( .A1(n689), .A2(n691), .ZN(n690) );
  XOR2_X1 U756 ( .A(G113), .B(n690), .Z(G15) );
  NOR2_X1 U757 ( .A1(n692), .A2(n691), .ZN(n693) );
  XOR2_X1 U758 ( .A(G116), .B(n693), .Z(G18) );
  XNOR2_X1 U759 ( .A(G125), .B(n694), .ZN(n695) );
  XNOR2_X1 U760 ( .A(n695), .B(KEYINPUT37), .ZN(G27) );
  XNOR2_X1 U761 ( .A(KEYINPUT53), .B(KEYINPUT121), .ZN(n746) );
  XOR2_X1 U762 ( .A(KEYINPUT117), .B(KEYINPUT118), .Z(n726) );
  NAND2_X1 U763 ( .A1(n697), .A2(n696), .ZN(n698) );
  XNOR2_X1 U764 ( .A(n698), .B(KEYINPUT49), .ZN(n699) );
  XNOR2_X1 U765 ( .A(KEYINPUT115), .B(n699), .ZN(n701) );
  NAND2_X1 U766 ( .A1(n701), .A2(n379), .ZN(n706) );
  XNOR2_X1 U767 ( .A(KEYINPUT50), .B(KEYINPUT116), .ZN(n703) );
  XNOR2_X1 U768 ( .A(n704), .B(n703), .ZN(n705) );
  NOR2_X1 U769 ( .A1(n706), .A2(n705), .ZN(n708) );
  OR2_X1 U770 ( .A1(n708), .A2(n707), .ZN(n709) );
  XNOR2_X1 U771 ( .A(KEYINPUT51), .B(n709), .ZN(n710) );
  NOR2_X1 U772 ( .A1(n710), .A2(n732), .ZN(n723) );
  NOR2_X1 U773 ( .A1(n712), .A2(n711), .ZN(n713) );
  NOR2_X1 U774 ( .A1(n714), .A2(n713), .ZN(n718) );
  NOR2_X1 U775 ( .A1(n716), .A2(n715), .ZN(n717) );
  NOR2_X1 U776 ( .A1(n718), .A2(n717), .ZN(n721) );
  BUF_X1 U777 ( .A(n719), .Z(n720) );
  INV_X1 U778 ( .A(n720), .ZN(n731) );
  NOR2_X1 U779 ( .A1(n721), .A2(n731), .ZN(n722) );
  NOR2_X1 U780 ( .A1(n723), .A2(n722), .ZN(n724) );
  XNOR2_X1 U781 ( .A(n724), .B(KEYINPUT52), .ZN(n725) );
  XNOR2_X1 U782 ( .A(n726), .B(n725), .ZN(n729) );
  NAND2_X1 U783 ( .A1(G952), .A2(n727), .ZN(n728) );
  NOR2_X1 U784 ( .A1(n729), .A2(n728), .ZN(n730) );
  XOR2_X1 U785 ( .A(KEYINPUT119), .B(n730), .Z(n734) );
  NOR2_X1 U786 ( .A1(n732), .A2(n731), .ZN(n733) );
  NOR2_X1 U787 ( .A1(n734), .A2(n733), .ZN(n735) );
  XNOR2_X1 U788 ( .A(KEYINPUT120), .B(n735), .ZN(n744) );
  NOR2_X1 U789 ( .A1(n761), .A2(KEYINPUT2), .ZN(n736) );
  XNOR2_X1 U790 ( .A(n736), .B(KEYINPUT78), .ZN(n739) );
  NOR2_X1 U791 ( .A1(n747), .A2(KEYINPUT2), .ZN(n738) );
  OR2_X1 U792 ( .A1(n739), .A2(n738), .ZN(n740) );
  NOR2_X1 U793 ( .A1(n741), .A2(n740), .ZN(n742) );
  NOR2_X1 U794 ( .A1(n742), .A2(G953), .ZN(n743) );
  NAND2_X1 U795 ( .A1(n744), .A2(n743), .ZN(n745) );
  XNOR2_X1 U796 ( .A(n746), .B(n745), .ZN(G75) );
  NAND2_X1 U797 ( .A1(n747), .A2(n765), .ZN(n751) );
  NAND2_X1 U798 ( .A1(G953), .A2(G224), .ZN(n748) );
  XNOR2_X1 U799 ( .A(KEYINPUT61), .B(n748), .ZN(n749) );
  NAND2_X1 U800 ( .A1(n749), .A2(G898), .ZN(n750) );
  NAND2_X1 U801 ( .A1(n751), .A2(n750), .ZN(n756) );
  XOR2_X1 U802 ( .A(KEYINPUT123), .B(n752), .Z(n754) );
  NOR2_X1 U803 ( .A1(n754), .A2(n753), .ZN(n755) );
  XNOR2_X1 U804 ( .A(n756), .B(n755), .ZN(n757) );
  XNOR2_X1 U805 ( .A(KEYINPUT124), .B(n757), .ZN(G69) );
  XNOR2_X1 U806 ( .A(n758), .B(KEYINPUT125), .ZN(n759) );
  XOR2_X1 U807 ( .A(n760), .B(n759), .Z(n763) );
  XOR2_X1 U808 ( .A(n763), .B(n761), .Z(n762) );
  NAND2_X1 U809 ( .A1(n762), .A2(n765), .ZN(n768) );
  XNOR2_X1 U810 ( .A(n763), .B(G227), .ZN(n764) );
  NOR2_X1 U811 ( .A1(n765), .A2(n764), .ZN(n766) );
  NAND2_X1 U812 ( .A1(G900), .A2(n766), .ZN(n767) );
  NAND2_X1 U813 ( .A1(n768), .A2(n767), .ZN(n769) );
  XOR2_X1 U814 ( .A(KEYINPUT126), .B(n769), .Z(G72) );
  XOR2_X1 U815 ( .A(G137), .B(n770), .Z(G39) );
endmodule

