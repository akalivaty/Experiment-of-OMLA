//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 1 0 1 1 0 0 0 1 0 1 1 1 1 0 1 1 0 0 0 1 1 1 1 1 1 1 0 0 1 0 0 0 0 1 0 0 1 1 1 1 1 1 0 1 1 1 0 1 1 0 1 1 1 0 1 1 1 1 0 1 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:34:44 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n443, new_n447, new_n449, new_n452, new_n453, new_n454, new_n455,
    new_n456, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n517, new_n518,
    new_n519, new_n520, new_n521, new_n522, new_n523, new_n524, new_n526,
    new_n527, new_n528, new_n529, new_n530, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n543,
    new_n544, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n556, new_n557, new_n558, new_n559, new_n561, new_n562, new_n563,
    new_n564, new_n565, new_n566, new_n567, new_n568, new_n569, new_n571,
    new_n572, new_n573, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n586, new_n587, new_n590,
    new_n591, new_n593, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n609, new_n610, new_n611, new_n612, new_n613, new_n614, new_n615,
    new_n616, new_n617, new_n618, new_n619, new_n620, new_n621, new_n622,
    new_n623, new_n624, new_n626, new_n627, new_n628, new_n629, new_n630,
    new_n631, new_n632, new_n633, new_n634, new_n635, new_n636, new_n637,
    new_n639, new_n640, new_n641, new_n642, new_n643, new_n644, new_n645,
    new_n646, new_n647, new_n648, new_n649, new_n650, new_n651, new_n652,
    new_n653, new_n654, new_n655, new_n656, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n814, new_n815, new_n816, new_n817,
    new_n818, new_n819, new_n820, new_n821, new_n822, new_n823, new_n824,
    new_n825, new_n826, new_n827, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1142,
    new_n1143, new_n1144, new_n1145, new_n1146, new_n1147, new_n1148,
    new_n1149;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  XOR2_X1   g006(.A(KEYINPUT64), .B(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(new_n443));
  XOR2_X1   g018(.A(new_n443), .B(KEYINPUT65), .Z(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(new_n449));
  XNOR2_X1  g024(.A(new_n449), .B(KEYINPUT66), .ZN(G234));
  NAND3_X1  g025(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g026(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n452));
  XNOR2_X1  g027(.A(new_n452), .B(KEYINPUT2), .ZN(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NOR4_X1   g029(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n455));
  INV_X1    g030(.A(new_n455), .ZN(new_n456));
  NOR2_X1   g031(.A1(new_n454), .A2(new_n456), .ZN(G325));
  INV_X1    g032(.A(G325), .ZN(G261));
  AOI22_X1  g033(.A1(new_n454), .A2(G2106), .B1(G567), .B2(new_n456), .ZN(G319));
  INV_X1    g034(.A(G2105), .ZN(new_n460));
  NAND3_X1  g035(.A1(new_n460), .A2(G101), .A3(G2104), .ZN(new_n461));
  XNOR2_X1  g036(.A(new_n461), .B(KEYINPUT68), .ZN(new_n462));
  INV_X1    g037(.A(KEYINPUT3), .ZN(new_n463));
  OAI21_X1  g038(.A(KEYINPUT67), .B1(new_n463), .B2(G2104), .ZN(new_n464));
  INV_X1    g039(.A(KEYINPUT67), .ZN(new_n465));
  INV_X1    g040(.A(G2104), .ZN(new_n466));
  NAND3_X1  g041(.A1(new_n465), .A2(new_n466), .A3(KEYINPUT3), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n463), .A2(G2104), .ZN(new_n468));
  NAND3_X1  g043(.A1(new_n464), .A2(new_n467), .A3(new_n468), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n460), .A2(G137), .ZN(new_n470));
  OAI21_X1  g045(.A(new_n462), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  XNOR2_X1  g046(.A(KEYINPUT3), .B(G2104), .ZN(new_n472));
  AOI22_X1  g047(.A1(new_n472), .A2(G125), .B1(G113), .B2(G2104), .ZN(new_n473));
  NOR2_X1   g048(.A1(new_n473), .A2(new_n460), .ZN(new_n474));
  NOR2_X1   g049(.A1(new_n471), .A2(new_n474), .ZN(G160));
  OR2_X1    g050(.A1(G100), .A2(G2105), .ZN(new_n476));
  OAI211_X1 g051(.A(new_n476), .B(G2104), .C1(G112), .C2(new_n460), .ZN(new_n477));
  XNOR2_X1  g052(.A(new_n477), .B(KEYINPUT70), .ZN(new_n478));
  INV_X1    g053(.A(KEYINPUT69), .ZN(new_n479));
  XNOR2_X1  g054(.A(new_n469), .B(new_n479), .ZN(new_n480));
  AND2_X1   g055(.A1(new_n480), .A2(new_n460), .ZN(new_n481));
  AND2_X1   g056(.A1(new_n481), .A2(G136), .ZN(new_n482));
  AND2_X1   g057(.A1(new_n480), .A2(G2105), .ZN(new_n483));
  AOI211_X1 g058(.A(new_n478), .B(new_n482), .C1(G124), .C2(new_n483), .ZN(G162));
  AND2_X1   g059(.A1(new_n467), .A2(new_n468), .ZN(new_n485));
  NAND4_X1  g060(.A1(new_n485), .A2(G126), .A3(G2105), .A4(new_n464), .ZN(new_n486));
  OR2_X1    g061(.A1(G102), .A2(G2105), .ZN(new_n487));
  OAI211_X1 g062(.A(new_n487), .B(G2104), .C1(G114), .C2(new_n460), .ZN(new_n488));
  NAND2_X1  g063(.A1(new_n486), .A2(new_n488), .ZN(new_n489));
  INV_X1    g064(.A(KEYINPUT4), .ZN(new_n490));
  INV_X1    g065(.A(G138), .ZN(new_n491));
  NOR2_X1   g066(.A1(new_n491), .A2(G2105), .ZN(new_n492));
  NAND3_X1  g067(.A1(new_n472), .A2(new_n490), .A3(new_n492), .ZN(new_n493));
  INV_X1    g068(.A(new_n493), .ZN(new_n494));
  INV_X1    g069(.A(KEYINPUT71), .ZN(new_n495));
  NAND4_X1  g070(.A1(new_n485), .A2(new_n495), .A3(new_n464), .A4(new_n492), .ZN(new_n496));
  NAND4_X1  g071(.A1(new_n464), .A2(new_n467), .A3(new_n468), .A4(new_n492), .ZN(new_n497));
  NAND2_X1  g072(.A1(new_n497), .A2(KEYINPUT71), .ZN(new_n498));
  NAND3_X1  g073(.A1(new_n496), .A2(KEYINPUT4), .A3(new_n498), .ZN(new_n499));
  AOI21_X1  g074(.A(new_n494), .B1(new_n499), .B2(KEYINPUT72), .ZN(new_n500));
  INV_X1    g075(.A(KEYINPUT72), .ZN(new_n501));
  NAND4_X1  g076(.A1(new_n496), .A2(new_n501), .A3(KEYINPUT4), .A4(new_n498), .ZN(new_n502));
  AOI21_X1  g077(.A(new_n489), .B1(new_n500), .B2(new_n502), .ZN(G164));
  INV_X1    g078(.A(G651), .ZN(new_n504));
  XNOR2_X1  g079(.A(KEYINPUT5), .B(G543), .ZN(new_n505));
  AOI21_X1  g080(.A(KEYINPUT73), .B1(new_n505), .B2(G62), .ZN(new_n506));
  AOI21_X1  g081(.A(new_n506), .B1(G75), .B2(G543), .ZN(new_n507));
  NAND3_X1  g082(.A1(new_n505), .A2(KEYINPUT73), .A3(G62), .ZN(new_n508));
  AOI21_X1  g083(.A(new_n504), .B1(new_n507), .B2(new_n508), .ZN(new_n509));
  XNOR2_X1  g084(.A(KEYINPUT6), .B(G651), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n505), .A2(new_n510), .ZN(new_n511));
  INV_X1    g086(.A(G88), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n510), .A2(G543), .ZN(new_n513));
  INV_X1    g088(.A(G50), .ZN(new_n514));
  OAI22_X1  g089(.A1(new_n511), .A2(new_n512), .B1(new_n513), .B2(new_n514), .ZN(new_n515));
  NOR2_X1   g090(.A1(new_n509), .A2(new_n515), .ZN(G166));
  NAND3_X1  g091(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n517));
  XNOR2_X1  g092(.A(new_n517), .B(KEYINPUT7), .ZN(new_n518));
  INV_X1    g093(.A(G51), .ZN(new_n519));
  OAI21_X1  g094(.A(new_n518), .B1(new_n513), .B2(new_n519), .ZN(new_n520));
  INV_X1    g095(.A(new_n505), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n510), .A2(G89), .ZN(new_n522));
  NAND2_X1  g097(.A1(G63), .A2(G651), .ZN(new_n523));
  AOI21_X1  g098(.A(new_n521), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  NOR2_X1   g099(.A1(new_n520), .A2(new_n524), .ZN(G168));
  INV_X1    g100(.A(G90), .ZN(new_n526));
  XNOR2_X1  g101(.A(KEYINPUT74), .B(G52), .ZN(new_n527));
  OAI22_X1  g102(.A1(new_n511), .A2(new_n526), .B1(new_n513), .B2(new_n527), .ZN(new_n528));
  AOI22_X1  g103(.A1(new_n505), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n529));
  NOR2_X1   g104(.A1(new_n529), .A2(new_n504), .ZN(new_n530));
  NOR2_X1   g105(.A1(new_n528), .A2(new_n530), .ZN(G171));
  INV_X1    g106(.A(G81), .ZN(new_n532));
  INV_X1    g107(.A(G43), .ZN(new_n533));
  OAI22_X1  g108(.A1(new_n511), .A2(new_n532), .B1(new_n513), .B2(new_n533), .ZN(new_n534));
  INV_X1    g109(.A(KEYINPUT75), .ZN(new_n535));
  XNOR2_X1  g110(.A(new_n534), .B(new_n535), .ZN(new_n536));
  AOI22_X1  g111(.A1(new_n505), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n537));
  OR2_X1    g112(.A1(new_n537), .A2(new_n504), .ZN(new_n538));
  NAND2_X1  g113(.A1(new_n536), .A2(new_n538), .ZN(new_n539));
  INV_X1    g114(.A(new_n539), .ZN(new_n540));
  NAND2_X1  g115(.A1(new_n540), .A2(G860), .ZN(G153));
  NAND4_X1  g116(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g117(.A1(G1), .A2(G3), .ZN(new_n543));
  XNOR2_X1  g118(.A(new_n543), .B(KEYINPUT8), .ZN(new_n544));
  NAND4_X1  g119(.A1(G319), .A2(G483), .A3(G661), .A4(new_n544), .ZN(G188));
  INV_X1    g120(.A(new_n513), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n546), .A2(G53), .ZN(new_n547));
  XNOR2_X1  g122(.A(new_n547), .B(KEYINPUT9), .ZN(new_n548));
  AND3_X1   g123(.A1(new_n505), .A2(new_n510), .A3(G91), .ZN(new_n549));
  XOR2_X1   g124(.A(new_n549), .B(KEYINPUT76), .Z(new_n550));
  AOI22_X1  g125(.A1(new_n505), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n551));
  OAI211_X1 g126(.A(new_n548), .B(new_n550), .C1(new_n504), .C2(new_n551), .ZN(G299));
  INV_X1    g127(.A(G171), .ZN(G301));
  INV_X1    g128(.A(G168), .ZN(G286));
  INV_X1    g129(.A(G166), .ZN(G303));
  OAI21_X1  g130(.A(G651), .B1(new_n505), .B2(G74), .ZN(new_n556));
  XNOR2_X1  g131(.A(new_n556), .B(KEYINPUT77), .ZN(new_n557));
  INV_X1    g132(.A(new_n511), .ZN(new_n558));
  AOI22_X1  g133(.A1(G87), .A2(new_n558), .B1(new_n546), .B2(G49), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n557), .A2(new_n559), .ZN(G288));
  AOI22_X1  g135(.A1(new_n505), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n561));
  INV_X1    g136(.A(G86), .ZN(new_n562));
  OAI22_X1  g137(.A1(new_n561), .A2(new_n504), .B1(new_n511), .B2(new_n562), .ZN(new_n563));
  INV_X1    g138(.A(new_n563), .ZN(new_n564));
  INV_X1    g139(.A(G48), .ZN(new_n565));
  OAI21_X1  g140(.A(KEYINPUT78), .B1(new_n513), .B2(new_n565), .ZN(new_n566));
  INV_X1    g141(.A(KEYINPUT78), .ZN(new_n567));
  NAND4_X1  g142(.A1(new_n510), .A2(new_n567), .A3(G48), .A4(G543), .ZN(new_n568));
  NAND2_X1  g143(.A1(new_n566), .A2(new_n568), .ZN(new_n569));
  NAND2_X1  g144(.A1(new_n564), .A2(new_n569), .ZN(G305));
  XOR2_X1   g145(.A(KEYINPUT79), .B(G85), .Z(new_n571));
  AOI22_X1  g146(.A1(new_n558), .A2(new_n571), .B1(new_n546), .B2(G47), .ZN(new_n572));
  AOI22_X1  g147(.A1(new_n505), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n573));
  OAI21_X1  g148(.A(new_n572), .B1(new_n504), .B2(new_n573), .ZN(G290));
  NAND2_X1  g149(.A1(G301), .A2(G868), .ZN(new_n575));
  NAND2_X1  g150(.A1(new_n558), .A2(G92), .ZN(new_n576));
  XOR2_X1   g151(.A(new_n576), .B(KEYINPUT10), .Z(new_n577));
  NAND2_X1  g152(.A1(G79), .A2(G543), .ZN(new_n578));
  INV_X1    g153(.A(G66), .ZN(new_n579));
  OAI21_X1  g154(.A(new_n578), .B1(new_n521), .B2(new_n579), .ZN(new_n580));
  AOI22_X1  g155(.A1(new_n580), .A2(G651), .B1(new_n546), .B2(G54), .ZN(new_n581));
  NAND2_X1  g156(.A1(new_n577), .A2(new_n581), .ZN(new_n582));
  INV_X1    g157(.A(new_n582), .ZN(new_n583));
  OAI21_X1  g158(.A(new_n575), .B1(new_n583), .B2(G868), .ZN(G321));
  XNOR2_X1  g159(.A(G321), .B(KEYINPUT80), .ZN(G284));
  INV_X1    g160(.A(G868), .ZN(new_n586));
  NAND2_X1  g161(.A1(G299), .A2(new_n586), .ZN(new_n587));
  OAI21_X1  g162(.A(new_n587), .B1(new_n586), .B2(G168), .ZN(G297));
  OAI21_X1  g163(.A(new_n587), .B1(new_n586), .B2(G168), .ZN(G280));
  NOR2_X1   g164(.A1(new_n582), .A2(G559), .ZN(new_n590));
  AOI21_X1  g165(.A(new_n590), .B1(G860), .B2(new_n583), .ZN(new_n591));
  XNOR2_X1  g166(.A(new_n591), .B(KEYINPUT81), .ZN(G148));
  NAND2_X1  g167(.A1(new_n539), .A2(new_n586), .ZN(new_n593));
  OAI21_X1  g168(.A(new_n593), .B1(new_n590), .B2(new_n586), .ZN(G323));
  XNOR2_X1  g169(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g170(.A1(new_n481), .A2(G135), .ZN(new_n596));
  NAND2_X1  g171(.A1(new_n483), .A2(G123), .ZN(new_n597));
  OR2_X1    g172(.A1(G99), .A2(G2105), .ZN(new_n598));
  OAI211_X1 g173(.A(new_n598), .B(G2104), .C1(G111), .C2(new_n460), .ZN(new_n599));
  NAND3_X1  g174(.A1(new_n596), .A2(new_n597), .A3(new_n599), .ZN(new_n600));
  OR2_X1    g175(.A1(new_n600), .A2(G2096), .ZN(new_n601));
  NAND2_X1  g176(.A1(new_n600), .A2(G2096), .ZN(new_n602));
  NOR2_X1   g177(.A1(new_n466), .A2(G2105), .ZN(new_n603));
  NAND2_X1  g178(.A1(new_n472), .A2(new_n603), .ZN(new_n604));
  XNOR2_X1  g179(.A(new_n604), .B(KEYINPUT12), .ZN(new_n605));
  XNOR2_X1  g180(.A(new_n605), .B(KEYINPUT13), .ZN(new_n606));
  XNOR2_X1  g181(.A(new_n606), .B(G2100), .ZN(new_n607));
  NAND3_X1  g182(.A1(new_n601), .A2(new_n602), .A3(new_n607), .ZN(G156));
  XNOR2_X1  g183(.A(G2427), .B(G2438), .ZN(new_n609));
  XNOR2_X1  g184(.A(new_n609), .B(G2430), .ZN(new_n610));
  XNOR2_X1  g185(.A(KEYINPUT15), .B(G2435), .ZN(new_n611));
  OR2_X1    g186(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  NAND2_X1  g187(.A1(new_n610), .A2(new_n611), .ZN(new_n613));
  NAND3_X1  g188(.A1(new_n612), .A2(KEYINPUT14), .A3(new_n613), .ZN(new_n614));
  XOR2_X1   g189(.A(G2443), .B(G2446), .Z(new_n615));
  XNOR2_X1  g190(.A(new_n614), .B(new_n615), .ZN(new_n616));
  XOR2_X1   g191(.A(G2451), .B(G2454), .Z(new_n617));
  XNOR2_X1  g192(.A(KEYINPUT82), .B(KEYINPUT16), .ZN(new_n618));
  XNOR2_X1  g193(.A(new_n617), .B(new_n618), .ZN(new_n619));
  XNOR2_X1  g194(.A(new_n616), .B(new_n619), .ZN(new_n620));
  XOR2_X1   g195(.A(G1341), .B(G1348), .Z(new_n621));
  NOR2_X1   g196(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  XNOR2_X1  g197(.A(new_n622), .B(KEYINPUT83), .ZN(new_n623));
  NAND2_X1  g198(.A1(new_n620), .A2(new_n621), .ZN(new_n624));
  AND3_X1   g199(.A1(new_n623), .A2(G14), .A3(new_n624), .ZN(G401));
  XOR2_X1   g200(.A(KEYINPUT84), .B(KEYINPUT18), .Z(new_n626));
  INV_X1    g201(.A(new_n626), .ZN(new_n627));
  XOR2_X1   g202(.A(G2084), .B(G2090), .Z(new_n628));
  XNOR2_X1  g203(.A(G2067), .B(G2678), .ZN(new_n629));
  NAND2_X1  g204(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  NAND2_X1  g205(.A1(new_n630), .A2(KEYINPUT17), .ZN(new_n631));
  NOR2_X1   g206(.A1(new_n628), .A2(new_n629), .ZN(new_n632));
  OAI21_X1  g207(.A(new_n627), .B1(new_n631), .B2(new_n632), .ZN(new_n633));
  XOR2_X1   g208(.A(G2072), .B(G2078), .Z(new_n634));
  AOI21_X1  g209(.A(new_n634), .B1(new_n630), .B2(new_n626), .ZN(new_n635));
  XNOR2_X1  g210(.A(new_n633), .B(new_n635), .ZN(new_n636));
  XNOR2_X1  g211(.A(G2096), .B(G2100), .ZN(new_n637));
  XNOR2_X1  g212(.A(new_n636), .B(new_n637), .ZN(G227));
  XOR2_X1   g213(.A(G1961), .B(G1966), .Z(new_n639));
  XNOR2_X1  g214(.A(new_n639), .B(KEYINPUT85), .ZN(new_n640));
  XNOR2_X1  g215(.A(G1956), .B(G2474), .ZN(new_n641));
  INV_X1    g216(.A(new_n641), .ZN(new_n642));
  NAND2_X1  g217(.A1(new_n640), .A2(new_n642), .ZN(new_n643));
  XNOR2_X1  g218(.A(G1971), .B(G1976), .ZN(new_n644));
  XNOR2_X1  g219(.A(new_n644), .B(KEYINPUT19), .ZN(new_n645));
  NOR2_X1   g220(.A1(new_n643), .A2(new_n645), .ZN(new_n646));
  XOR2_X1   g221(.A(new_n646), .B(KEYINPUT20), .Z(new_n647));
  OR2_X1    g222(.A1(new_n640), .A2(new_n642), .ZN(new_n648));
  NAND3_X1  g223(.A1(new_n648), .A2(new_n645), .A3(new_n643), .ZN(new_n649));
  OAI211_X1 g224(.A(new_n647), .B(new_n649), .C1(new_n645), .C2(new_n648), .ZN(new_n650));
  XNOR2_X1  g225(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n651));
  XNOR2_X1  g226(.A(new_n650), .B(new_n651), .ZN(new_n652));
  XNOR2_X1  g227(.A(G1991), .B(G1996), .ZN(new_n653));
  XNOR2_X1  g228(.A(new_n652), .B(new_n653), .ZN(new_n654));
  XNOR2_X1  g229(.A(G1981), .B(G1986), .ZN(new_n655));
  XOR2_X1   g230(.A(new_n654), .B(new_n655), .Z(new_n656));
  INV_X1    g231(.A(new_n656), .ZN(G229));
  INV_X1    g232(.A(G16), .ZN(new_n658));
  NAND2_X1  g233(.A1(new_n658), .A2(G23), .ZN(new_n659));
  INV_X1    g234(.A(G288), .ZN(new_n660));
  OAI21_X1  g235(.A(new_n659), .B1(new_n660), .B2(new_n658), .ZN(new_n661));
  XNOR2_X1  g236(.A(new_n661), .B(KEYINPUT33), .ZN(new_n662));
  INV_X1    g237(.A(G1976), .ZN(new_n663));
  XNOR2_X1  g238(.A(new_n662), .B(new_n663), .ZN(new_n664));
  NOR2_X1   g239(.A1(G166), .A2(new_n658), .ZN(new_n665));
  AOI21_X1  g240(.A(new_n665), .B1(new_n658), .B2(G22), .ZN(new_n666));
  INV_X1    g241(.A(G1971), .ZN(new_n667));
  NOR2_X1   g242(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  MUX2_X1   g243(.A(G6), .B(G305), .S(G16), .Z(new_n669));
  XNOR2_X1  g244(.A(KEYINPUT32), .B(G1981), .ZN(new_n670));
  XNOR2_X1  g245(.A(new_n669), .B(new_n670), .ZN(new_n671));
  NOR2_X1   g246(.A1(new_n668), .A2(new_n671), .ZN(new_n672));
  NAND2_X1  g247(.A1(new_n666), .A2(new_n667), .ZN(new_n673));
  NAND2_X1  g248(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  NOR2_X1   g249(.A1(new_n664), .A2(new_n674), .ZN(new_n675));
  INV_X1    g250(.A(new_n675), .ZN(new_n676));
  XOR2_X1   g251(.A(KEYINPUT35), .B(G1991), .Z(new_n677));
  NAND2_X1  g252(.A1(new_n481), .A2(G131), .ZN(new_n678));
  NAND2_X1  g253(.A1(new_n483), .A2(G119), .ZN(new_n679));
  NOR2_X1   g254(.A1(new_n460), .A2(G107), .ZN(new_n680));
  OAI21_X1  g255(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n681));
  OAI211_X1 g256(.A(new_n678), .B(new_n679), .C1(new_n680), .C2(new_n681), .ZN(new_n682));
  MUX2_X1   g257(.A(G25), .B(new_n682), .S(G29), .Z(new_n683));
  XOR2_X1   g258(.A(new_n683), .B(KEYINPUT86), .Z(new_n684));
  AOI22_X1  g259(.A1(new_n676), .A2(KEYINPUT34), .B1(new_n677), .B2(new_n684), .ZN(new_n685));
  NAND2_X1  g260(.A1(new_n658), .A2(G24), .ZN(new_n686));
  XOR2_X1   g261(.A(new_n686), .B(KEYINPUT87), .Z(new_n687));
  AOI21_X1  g262(.A(new_n687), .B1(G290), .B2(G16), .ZN(new_n688));
  XOR2_X1   g263(.A(new_n688), .B(G1986), .Z(new_n689));
  INV_X1    g264(.A(KEYINPUT34), .ZN(new_n690));
  AOI21_X1  g265(.A(new_n689), .B1(new_n675), .B2(new_n690), .ZN(new_n691));
  OAI211_X1 g266(.A(new_n685), .B(new_n691), .C1(new_n677), .C2(new_n684), .ZN(new_n692));
  AND2_X1   g267(.A1(KEYINPUT88), .A2(KEYINPUT36), .ZN(new_n693));
  XNOR2_X1  g268(.A(new_n692), .B(new_n693), .ZN(new_n694));
  INV_X1    g269(.A(G29), .ZN(new_n695));
  INV_X1    g270(.A(KEYINPUT24), .ZN(new_n696));
  OAI21_X1  g271(.A(new_n695), .B1(new_n696), .B2(G34), .ZN(new_n697));
  AOI21_X1  g272(.A(new_n697), .B1(new_n696), .B2(G34), .ZN(new_n698));
  AOI21_X1  g273(.A(new_n698), .B1(G160), .B2(G29), .ZN(new_n699));
  NOR2_X1   g274(.A1(new_n699), .A2(G2084), .ZN(new_n700));
  NAND2_X1  g275(.A1(new_n658), .A2(G4), .ZN(new_n701));
  OAI21_X1  g276(.A(new_n701), .B1(new_n583), .B2(new_n658), .ZN(new_n702));
  XNOR2_X1  g277(.A(KEYINPUT89), .B(G1348), .ZN(new_n703));
  XNOR2_X1  g278(.A(new_n703), .B(KEYINPUT90), .ZN(new_n704));
  XNOR2_X1  g279(.A(new_n702), .B(new_n704), .ZN(new_n705));
  INV_X1    g280(.A(G1961), .ZN(new_n706));
  NOR2_X1   g281(.A1(G171), .A2(new_n658), .ZN(new_n707));
  AOI21_X1  g282(.A(new_n707), .B1(G5), .B2(new_n658), .ZN(new_n708));
  AOI211_X1 g283(.A(new_n700), .B(new_n705), .C1(new_n706), .C2(new_n708), .ZN(new_n709));
  NAND2_X1  g284(.A1(G162), .A2(G29), .ZN(new_n710));
  OAI21_X1  g285(.A(new_n710), .B1(G29), .B2(G35), .ZN(new_n711));
  XOR2_X1   g286(.A(KEYINPUT29), .B(G2090), .Z(new_n712));
  OR2_X1    g287(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  NAND2_X1  g288(.A1(new_n658), .A2(G19), .ZN(new_n714));
  OAI21_X1  g289(.A(new_n714), .B1(new_n540), .B2(new_n658), .ZN(new_n715));
  XOR2_X1   g290(.A(new_n715), .B(G1341), .Z(new_n716));
  NAND2_X1  g291(.A1(new_n481), .A2(G140), .ZN(new_n717));
  NAND2_X1  g292(.A1(new_n483), .A2(G128), .ZN(new_n718));
  NOR2_X1   g293(.A1(new_n460), .A2(G116), .ZN(new_n719));
  OAI21_X1  g294(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n720));
  OAI211_X1 g295(.A(new_n717), .B(new_n718), .C1(new_n719), .C2(new_n720), .ZN(new_n721));
  NAND2_X1  g296(.A1(new_n721), .A2(G29), .ZN(new_n722));
  NAND2_X1  g297(.A1(new_n695), .A2(G26), .ZN(new_n723));
  XNOR2_X1  g298(.A(new_n723), .B(KEYINPUT28), .ZN(new_n724));
  NAND2_X1  g299(.A1(new_n722), .A2(new_n724), .ZN(new_n725));
  AOI22_X1  g300(.A1(new_n711), .A2(new_n712), .B1(G2067), .B2(new_n725), .ZN(new_n726));
  NAND4_X1  g301(.A1(new_n709), .A2(new_n713), .A3(new_n716), .A4(new_n726), .ZN(new_n727));
  NAND2_X1  g302(.A1(new_n481), .A2(G141), .ZN(new_n728));
  NAND2_X1  g303(.A1(new_n483), .A2(G129), .ZN(new_n729));
  NAND3_X1  g304(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n730));
  INV_X1    g305(.A(KEYINPUT26), .ZN(new_n731));
  OR2_X1    g306(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  NAND2_X1  g307(.A1(new_n730), .A2(new_n731), .ZN(new_n733));
  AOI22_X1  g308(.A1(new_n732), .A2(new_n733), .B1(G105), .B2(new_n603), .ZN(new_n734));
  NAND3_X1  g309(.A1(new_n728), .A2(new_n729), .A3(new_n734), .ZN(new_n735));
  INV_X1    g310(.A(new_n735), .ZN(new_n736));
  NOR2_X1   g311(.A1(new_n736), .A2(new_n695), .ZN(new_n737));
  AOI21_X1  g312(.A(new_n737), .B1(new_n695), .B2(G32), .ZN(new_n738));
  XNOR2_X1  g313(.A(KEYINPUT27), .B(G1996), .ZN(new_n739));
  NOR2_X1   g314(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  INV_X1    g315(.A(G1956), .ZN(new_n741));
  NAND2_X1  g316(.A1(new_n658), .A2(G20), .ZN(new_n742));
  XOR2_X1   g317(.A(new_n742), .B(KEYINPUT23), .Z(new_n743));
  AOI21_X1  g318(.A(new_n743), .B1(G299), .B2(G16), .ZN(new_n744));
  XOR2_X1   g319(.A(new_n744), .B(KEYINPUT98), .Z(new_n745));
  AOI21_X1  g320(.A(new_n740), .B1(new_n741), .B2(new_n745), .ZN(new_n746));
  OAI221_X1 g321(.A(new_n746), .B1(new_n741), .B2(new_n745), .C1(G2067), .C2(new_n725), .ZN(new_n747));
  NAND2_X1  g322(.A1(new_n695), .A2(G27), .ZN(new_n748));
  XNOR2_X1  g323(.A(new_n748), .B(KEYINPUT97), .ZN(new_n749));
  AND2_X1   g324(.A1(new_n497), .A2(KEYINPUT71), .ZN(new_n750));
  OAI21_X1  g325(.A(KEYINPUT4), .B1(new_n497), .B2(KEYINPUT71), .ZN(new_n751));
  OAI21_X1  g326(.A(KEYINPUT72), .B1(new_n750), .B2(new_n751), .ZN(new_n752));
  NAND3_X1  g327(.A1(new_n752), .A2(new_n502), .A3(new_n493), .ZN(new_n753));
  INV_X1    g328(.A(new_n489), .ZN(new_n754));
  NAND2_X1  g329(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  AOI21_X1  g330(.A(new_n749), .B1(new_n755), .B2(G29), .ZN(new_n756));
  INV_X1    g331(.A(G2078), .ZN(new_n757));
  XNOR2_X1  g332(.A(new_n756), .B(new_n757), .ZN(new_n758));
  NOR3_X1   g333(.A1(new_n727), .A2(new_n747), .A3(new_n758), .ZN(new_n759));
  XOR2_X1   g334(.A(KEYINPUT31), .B(G11), .Z(new_n760));
  INV_X1    g335(.A(G28), .ZN(new_n761));
  NOR2_X1   g336(.A1(new_n761), .A2(KEYINPUT30), .ZN(new_n762));
  XNOR2_X1  g337(.A(new_n762), .B(KEYINPUT93), .ZN(new_n763));
  AOI21_X1  g338(.A(G29), .B1(new_n761), .B2(KEYINPUT30), .ZN(new_n764));
  AOI21_X1  g339(.A(new_n760), .B1(new_n763), .B2(new_n764), .ZN(new_n765));
  OAI21_X1  g340(.A(new_n765), .B1(new_n600), .B2(new_n695), .ZN(new_n766));
  XOR2_X1   g341(.A(new_n766), .B(KEYINPUT94), .Z(new_n767));
  NAND2_X1  g342(.A1(new_n658), .A2(G21), .ZN(new_n768));
  OAI21_X1  g343(.A(new_n768), .B1(G168), .B2(new_n658), .ZN(new_n769));
  INV_X1    g344(.A(G1966), .ZN(new_n770));
  XNOR2_X1  g345(.A(new_n769), .B(new_n770), .ZN(new_n771));
  NOR2_X1   g346(.A1(new_n708), .A2(new_n706), .ZN(new_n772));
  XNOR2_X1  g347(.A(new_n772), .B(KEYINPUT95), .ZN(new_n773));
  NAND3_X1  g348(.A1(new_n767), .A2(new_n771), .A3(new_n773), .ZN(new_n774));
  XNOR2_X1  g349(.A(new_n774), .B(KEYINPUT96), .ZN(new_n775));
  NAND2_X1  g350(.A1(new_n695), .A2(G33), .ZN(new_n776));
  NAND3_X1  g351(.A1(new_n460), .A2(G103), .A3(G2104), .ZN(new_n777));
  XOR2_X1   g352(.A(new_n777), .B(KEYINPUT25), .Z(new_n778));
  AOI22_X1  g353(.A1(new_n472), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n779));
  OAI21_X1  g354(.A(new_n778), .B1(new_n779), .B2(new_n460), .ZN(new_n780));
  AOI21_X1  g355(.A(new_n780), .B1(new_n481), .B2(G139), .ZN(new_n781));
  OAI21_X1  g356(.A(new_n776), .B1(new_n781), .B2(new_n695), .ZN(new_n782));
  XOR2_X1   g357(.A(new_n782), .B(KEYINPUT91), .Z(new_n783));
  INV_X1    g358(.A(G2072), .ZN(new_n784));
  OR2_X1    g359(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  AOI22_X1  g360(.A1(new_n738), .A2(new_n739), .B1(G2084), .B2(new_n699), .ZN(new_n786));
  NAND2_X1  g361(.A1(new_n783), .A2(new_n784), .ZN(new_n787));
  NAND3_X1  g362(.A1(new_n785), .A2(new_n786), .A3(new_n787), .ZN(new_n788));
  XNOR2_X1  g363(.A(new_n788), .B(KEYINPUT92), .ZN(new_n789));
  AND3_X1   g364(.A1(new_n759), .A2(new_n775), .A3(new_n789), .ZN(new_n790));
  NAND2_X1  g365(.A1(new_n694), .A2(new_n790), .ZN(G150));
  INV_X1    g366(.A(G150), .ZN(G311));
  AND2_X1   g367(.A1(new_n505), .A2(G67), .ZN(new_n793));
  AND2_X1   g368(.A1(G80), .A2(G543), .ZN(new_n794));
  OAI21_X1  g369(.A(G651), .B1(new_n793), .B2(new_n794), .ZN(new_n795));
  INV_X1    g370(.A(KEYINPUT99), .ZN(new_n796));
  OR2_X1    g371(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  NAND2_X1  g372(.A1(new_n795), .A2(new_n796), .ZN(new_n798));
  AOI22_X1  g373(.A1(G93), .A2(new_n558), .B1(new_n546), .B2(G55), .ZN(new_n799));
  NAND3_X1  g374(.A1(new_n797), .A2(new_n798), .A3(new_n799), .ZN(new_n800));
  XOR2_X1   g375(.A(KEYINPUT101), .B(G860), .Z(new_n801));
  NAND2_X1  g376(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  XOR2_X1   g377(.A(KEYINPUT102), .B(KEYINPUT37), .Z(new_n803));
  XNOR2_X1  g378(.A(new_n802), .B(new_n803), .ZN(new_n804));
  NAND2_X1  g379(.A1(new_n583), .A2(G559), .ZN(new_n805));
  XNOR2_X1  g380(.A(new_n805), .B(KEYINPUT100), .ZN(new_n806));
  XNOR2_X1  g381(.A(new_n806), .B(KEYINPUT38), .ZN(new_n807));
  OR2_X1    g382(.A1(new_n539), .A2(new_n800), .ZN(new_n808));
  NAND2_X1  g383(.A1(new_n539), .A2(new_n800), .ZN(new_n809));
  NAND2_X1  g384(.A1(new_n808), .A2(new_n809), .ZN(new_n810));
  XNOR2_X1  g385(.A(new_n807), .B(new_n810), .ZN(new_n811));
  XNOR2_X1  g386(.A(new_n811), .B(KEYINPUT39), .ZN(new_n812));
  OAI21_X1  g387(.A(new_n804), .B1(new_n812), .B2(new_n801), .ZN(G145));
  INV_X1    g388(.A(KEYINPUT103), .ZN(new_n814));
  NAND2_X1  g389(.A1(new_n755), .A2(new_n814), .ZN(new_n815));
  NAND3_X1  g390(.A1(new_n753), .A2(KEYINPUT103), .A3(new_n754), .ZN(new_n816));
  AND2_X1   g391(.A1(new_n815), .A2(new_n816), .ZN(new_n817));
  INV_X1    g392(.A(new_n817), .ZN(new_n818));
  INV_X1    g393(.A(KEYINPUT104), .ZN(new_n819));
  NOR2_X1   g394(.A1(new_n781), .A2(new_n819), .ZN(new_n820));
  XNOR2_X1  g395(.A(new_n736), .B(new_n820), .ZN(new_n821));
  AND2_X1   g396(.A1(new_n821), .A2(new_n721), .ZN(new_n822));
  NOR2_X1   g397(.A1(new_n821), .A2(new_n721), .ZN(new_n823));
  OAI21_X1  g398(.A(new_n818), .B1(new_n822), .B2(new_n823), .ZN(new_n824));
  OR2_X1    g399(.A1(new_n821), .A2(new_n721), .ZN(new_n825));
  NAND2_X1  g400(.A1(new_n821), .A2(new_n721), .ZN(new_n826));
  NAND3_X1  g401(.A1(new_n825), .A2(new_n817), .A3(new_n826), .ZN(new_n827));
  NAND2_X1  g402(.A1(new_n824), .A2(new_n827), .ZN(new_n828));
  XNOR2_X1  g403(.A(new_n682), .B(KEYINPUT105), .ZN(new_n829));
  XNOR2_X1  g404(.A(new_n829), .B(new_n605), .ZN(new_n830));
  NAND2_X1  g405(.A1(new_n481), .A2(G142), .ZN(new_n831));
  NAND2_X1  g406(.A1(new_n483), .A2(G130), .ZN(new_n832));
  OR2_X1    g407(.A1(G106), .A2(G2105), .ZN(new_n833));
  OAI211_X1 g408(.A(new_n833), .B(G2104), .C1(G118), .C2(new_n460), .ZN(new_n834));
  NAND3_X1  g409(.A1(new_n831), .A2(new_n832), .A3(new_n834), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n830), .A2(new_n835), .ZN(new_n836));
  OR2_X1    g411(.A1(new_n829), .A2(new_n605), .ZN(new_n837));
  INV_X1    g412(.A(new_n835), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n829), .A2(new_n605), .ZN(new_n839));
  NAND3_X1  g414(.A1(new_n837), .A2(new_n838), .A3(new_n839), .ZN(new_n840));
  NAND2_X1  g415(.A1(new_n836), .A2(new_n840), .ZN(new_n841));
  INV_X1    g416(.A(KEYINPUT106), .ZN(new_n842));
  AND3_X1   g417(.A1(new_n828), .A2(new_n841), .A3(new_n842), .ZN(new_n843));
  AOI21_X1  g418(.A(new_n842), .B1(new_n828), .B2(new_n841), .ZN(new_n844));
  OAI22_X1  g419(.A1(new_n843), .A2(new_n844), .B1(new_n841), .B2(new_n828), .ZN(new_n845));
  XOR2_X1   g420(.A(new_n600), .B(G160), .Z(new_n846));
  XOR2_X1   g421(.A(new_n846), .B(G162), .Z(new_n847));
  NAND2_X1  g422(.A1(new_n845), .A2(new_n847), .ZN(new_n848));
  INV_X1    g423(.A(new_n828), .ZN(new_n849));
  INV_X1    g424(.A(new_n841), .ZN(new_n850));
  AOI21_X1  g425(.A(new_n847), .B1(new_n849), .B2(new_n850), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n828), .A2(new_n841), .ZN(new_n852));
  AOI21_X1  g427(.A(G37), .B1(new_n851), .B2(new_n852), .ZN(new_n853));
  AND3_X1   g428(.A1(new_n848), .A2(KEYINPUT40), .A3(new_n853), .ZN(new_n854));
  AOI21_X1  g429(.A(KEYINPUT40), .B1(new_n848), .B2(new_n853), .ZN(new_n855));
  NOR2_X1   g430(.A1(new_n854), .A2(new_n855), .ZN(G395));
  NAND2_X1  g431(.A1(new_n800), .A2(new_n586), .ZN(new_n857));
  XNOR2_X1  g432(.A(G290), .B(G288), .ZN(new_n858));
  AND2_X1   g433(.A1(new_n858), .A2(KEYINPUT107), .ZN(new_n859));
  XNOR2_X1  g434(.A(G166), .B(G305), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  NOR2_X1   g436(.A1(new_n858), .A2(KEYINPUT107), .ZN(new_n862));
  OR2_X1    g437(.A1(new_n859), .A2(new_n862), .ZN(new_n863));
  OAI21_X1  g438(.A(new_n861), .B1(new_n863), .B2(new_n860), .ZN(new_n864));
  INV_X1    g439(.A(KEYINPUT108), .ZN(new_n865));
  XNOR2_X1  g440(.A(new_n864), .B(new_n865), .ZN(new_n866));
  INV_X1    g441(.A(new_n866), .ZN(new_n867));
  MUX2_X1   g442(.A(new_n864), .B(new_n867), .S(KEYINPUT42), .Z(new_n868));
  AND2_X1   g443(.A1(new_n808), .A2(new_n809), .ZN(new_n869));
  XNOR2_X1  g444(.A(new_n869), .B(new_n590), .ZN(new_n870));
  OR2_X1    g445(.A1(new_n582), .A2(G299), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n582), .A2(G299), .ZN(new_n872));
  AND3_X1   g447(.A1(new_n871), .A2(KEYINPUT41), .A3(new_n872), .ZN(new_n873));
  AOI21_X1  g448(.A(KEYINPUT41), .B1(new_n871), .B2(new_n872), .ZN(new_n874));
  NOR2_X1   g449(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  NOR2_X1   g450(.A1(new_n870), .A2(new_n875), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n871), .A2(new_n872), .ZN(new_n877));
  AOI21_X1  g452(.A(new_n876), .B1(new_n877), .B2(new_n870), .ZN(new_n878));
  XNOR2_X1  g453(.A(new_n868), .B(new_n878), .ZN(new_n879));
  OAI21_X1  g454(.A(new_n857), .B1(new_n879), .B2(new_n586), .ZN(G295));
  OAI21_X1  g455(.A(new_n857), .B1(new_n879), .B2(new_n586), .ZN(G331));
  XOR2_X1   g456(.A(KEYINPUT109), .B(KEYINPUT44), .Z(new_n882));
  INV_X1    g457(.A(KEYINPUT43), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n869), .A2(G301), .ZN(new_n884));
  AOI21_X1  g459(.A(G301), .B1(new_n808), .B2(new_n809), .ZN(new_n885));
  INV_X1    g460(.A(new_n885), .ZN(new_n886));
  NAND3_X1  g461(.A1(new_n884), .A2(G168), .A3(new_n886), .ZN(new_n887));
  NOR2_X1   g462(.A1(new_n810), .A2(G171), .ZN(new_n888));
  OAI21_X1  g463(.A(G286), .B1(new_n888), .B2(new_n885), .ZN(new_n889));
  AND3_X1   g464(.A1(new_n887), .A2(new_n889), .A3(new_n875), .ZN(new_n890));
  AOI21_X1  g465(.A(new_n877), .B1(new_n887), .B2(new_n889), .ZN(new_n891));
  OAI21_X1  g466(.A(KEYINPUT110), .B1(new_n890), .B2(new_n891), .ZN(new_n892));
  NAND3_X1  g467(.A1(new_n887), .A2(new_n889), .A3(new_n875), .ZN(new_n893));
  INV_X1    g468(.A(KEYINPUT110), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n892), .A2(new_n895), .ZN(new_n896));
  AOI21_X1  g471(.A(G37), .B1(new_n896), .B2(new_n866), .ZN(new_n897));
  NAND3_X1  g472(.A1(new_n867), .A2(new_n892), .A3(new_n895), .ZN(new_n898));
  AOI21_X1  g473(.A(new_n883), .B1(new_n897), .B2(new_n898), .ZN(new_n899));
  NOR2_X1   g474(.A1(new_n896), .A2(new_n866), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n887), .A2(new_n889), .ZN(new_n901));
  INV_X1    g476(.A(new_n877), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n903), .A2(new_n893), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n866), .A2(new_n904), .ZN(new_n905));
  INV_X1    g480(.A(G37), .ZN(new_n906));
  NAND2_X1  g481(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  NOR3_X1   g482(.A1(new_n900), .A2(new_n907), .A3(KEYINPUT43), .ZN(new_n908));
  OAI21_X1  g483(.A(new_n882), .B1(new_n899), .B2(new_n908), .ZN(new_n909));
  INV_X1    g484(.A(KEYINPUT111), .ZN(new_n910));
  OAI21_X1  g485(.A(new_n910), .B1(new_n900), .B2(new_n907), .ZN(new_n911));
  AOI21_X1  g486(.A(G37), .B1(new_n866), .B2(new_n904), .ZN(new_n912));
  NAND3_X1  g487(.A1(new_n898), .A2(KEYINPUT111), .A3(new_n912), .ZN(new_n913));
  AND3_X1   g488(.A1(new_n911), .A2(KEYINPUT43), .A3(new_n913), .ZN(new_n914));
  NAND3_X1  g489(.A1(new_n897), .A2(new_n883), .A3(new_n898), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n915), .A2(KEYINPUT44), .ZN(new_n916));
  OAI21_X1  g491(.A(new_n909), .B1(new_n914), .B2(new_n916), .ZN(G397));
  INV_X1    g492(.A(G1384), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n817), .A2(new_n918), .ZN(new_n919));
  INV_X1    g494(.A(KEYINPUT45), .ZN(new_n920));
  NAND2_X1  g495(.A1(G160), .A2(G40), .ZN(new_n921));
  INV_X1    g496(.A(new_n921), .ZN(new_n922));
  NAND3_X1  g497(.A1(new_n919), .A2(new_n920), .A3(new_n922), .ZN(new_n923));
  INV_X1    g498(.A(KEYINPUT113), .ZN(new_n924));
  XNOR2_X1  g499(.A(new_n923), .B(new_n924), .ZN(new_n925));
  INV_X1    g500(.A(G2067), .ZN(new_n926));
  XNOR2_X1  g501(.A(new_n721), .B(new_n926), .ZN(new_n927));
  INV_X1    g502(.A(G1996), .ZN(new_n928));
  OAI21_X1  g503(.A(new_n927), .B1(new_n928), .B2(new_n736), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n925), .A2(new_n929), .ZN(new_n930));
  NOR2_X1   g505(.A1(new_n923), .A2(G1996), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n931), .A2(new_n736), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n930), .A2(new_n932), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n933), .A2(KEYINPUT114), .ZN(new_n934));
  OR3_X1    g509(.A1(new_n923), .A2(G1986), .A3(G290), .ZN(new_n935));
  NAND2_X1  g510(.A1(G290), .A2(G1986), .ZN(new_n936));
  OAI21_X1  g511(.A(new_n935), .B1(new_n923), .B2(new_n936), .ZN(new_n937));
  XNOR2_X1  g512(.A(new_n937), .B(KEYINPUT112), .ZN(new_n938));
  INV_X1    g513(.A(KEYINPUT114), .ZN(new_n939));
  NAND3_X1  g514(.A1(new_n930), .A2(new_n939), .A3(new_n932), .ZN(new_n940));
  INV_X1    g515(.A(new_n677), .ZN(new_n941));
  AND2_X1   g516(.A1(new_n682), .A2(new_n941), .ZN(new_n942));
  NOR2_X1   g517(.A1(new_n682), .A2(new_n941), .ZN(new_n943));
  OAI21_X1  g518(.A(new_n925), .B1(new_n942), .B2(new_n943), .ZN(new_n944));
  AND4_X1   g519(.A1(new_n934), .A2(new_n938), .A3(new_n940), .A4(new_n944), .ZN(new_n945));
  INV_X1    g520(.A(KEYINPUT54), .ZN(new_n946));
  NOR2_X1   g521(.A1(new_n920), .A2(G1384), .ZN(new_n947));
  AOI21_X1  g522(.A(KEYINPUT118), .B1(new_n755), .B2(new_n947), .ZN(new_n948));
  INV_X1    g523(.A(KEYINPUT118), .ZN(new_n949));
  INV_X1    g524(.A(new_n947), .ZN(new_n950));
  AOI211_X1 g525(.A(new_n949), .B(new_n950), .C1(new_n753), .C2(new_n754), .ZN(new_n951));
  NOR2_X1   g526(.A1(new_n948), .A2(new_n951), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n755), .A2(new_n918), .ZN(new_n953));
  AOI21_X1  g528(.A(new_n921), .B1(new_n953), .B2(new_n920), .ZN(new_n954));
  NAND4_X1  g529(.A1(new_n952), .A2(KEYINPUT53), .A3(new_n954), .A4(new_n757), .ZN(new_n955));
  AOI21_X1  g530(.A(G1384), .B1(new_n753), .B2(new_n754), .ZN(new_n956));
  INV_X1    g531(.A(KEYINPUT50), .ZN(new_n957));
  OAI21_X1  g532(.A(new_n922), .B1(new_n956), .B2(new_n957), .ZN(new_n958));
  AOI211_X1 g533(.A(KEYINPUT50), .B(G1384), .C1(new_n753), .C2(new_n754), .ZN(new_n959));
  OAI21_X1  g534(.A(new_n706), .B1(new_n958), .B2(new_n959), .ZN(new_n960));
  NAND3_X1  g535(.A1(new_n815), .A2(new_n816), .A3(new_n947), .ZN(new_n961));
  NAND3_X1  g536(.A1(new_n954), .A2(new_n757), .A3(new_n961), .ZN(new_n962));
  INV_X1    g537(.A(KEYINPUT125), .ZN(new_n963));
  INV_X1    g538(.A(KEYINPUT53), .ZN(new_n964));
  AND3_X1   g539(.A1(new_n962), .A2(new_n963), .A3(new_n964), .ZN(new_n965));
  AOI21_X1  g540(.A(new_n963), .B1(new_n962), .B2(new_n964), .ZN(new_n966));
  OAI211_X1 g541(.A(new_n955), .B(new_n960), .C1(new_n965), .C2(new_n966), .ZN(new_n967));
  AND2_X1   g542(.A1(new_n967), .A2(G171), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n919), .A2(new_n920), .ZN(new_n969));
  AND4_X1   g544(.A1(KEYINPUT53), .A2(new_n961), .A3(new_n757), .A4(new_n922), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n969), .A2(new_n970), .ZN(new_n971));
  OAI211_X1 g546(.A(new_n960), .B(new_n971), .C1(new_n965), .C2(new_n966), .ZN(new_n972));
  NOR2_X1   g547(.A1(new_n972), .A2(G171), .ZN(new_n973));
  OAI21_X1  g548(.A(new_n946), .B1(new_n968), .B2(new_n973), .ZN(new_n974));
  INV_X1    g549(.A(G8), .ZN(new_n975));
  NOR2_X1   g550(.A1(G168), .A2(new_n975), .ZN(new_n976));
  INV_X1    g551(.A(new_n976), .ZN(new_n977));
  OAI21_X1  g552(.A(new_n920), .B1(G164), .B2(G1384), .ZN(new_n978));
  OAI21_X1  g553(.A(new_n949), .B1(G164), .B2(new_n950), .ZN(new_n979));
  NAND3_X1  g554(.A1(new_n755), .A2(KEYINPUT118), .A3(new_n947), .ZN(new_n980));
  NAND4_X1  g555(.A1(new_n978), .A2(new_n979), .A3(new_n980), .A4(new_n922), .ZN(new_n981));
  NOR2_X1   g556(.A1(new_n958), .A2(new_n959), .ZN(new_n982));
  INV_X1    g557(.A(G2084), .ZN(new_n983));
  AOI22_X1  g558(.A1(new_n770), .A2(new_n981), .B1(new_n982), .B2(new_n983), .ZN(new_n984));
  OAI211_X1 g559(.A(KEYINPUT51), .B(new_n977), .C1(new_n984), .C2(new_n975), .ZN(new_n985));
  INV_X1    g560(.A(KEYINPUT51), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n979), .A2(new_n980), .ZN(new_n987));
  OAI21_X1  g562(.A(new_n922), .B1(new_n956), .B2(KEYINPUT45), .ZN(new_n988));
  OAI21_X1  g563(.A(new_n770), .B1(new_n987), .B2(new_n988), .ZN(new_n989));
  AOI21_X1  g564(.A(new_n921), .B1(new_n953), .B2(KEYINPUT50), .ZN(new_n990));
  INV_X1    g565(.A(new_n959), .ZN(new_n991));
  NAND3_X1  g566(.A1(new_n990), .A2(new_n983), .A3(new_n991), .ZN(new_n992));
  NAND2_X1  g567(.A1(new_n989), .A2(new_n992), .ZN(new_n993));
  OAI211_X1 g568(.A(new_n986), .B(G8), .C1(new_n993), .C2(G286), .ZN(new_n994));
  AOI21_X1  g569(.A(KEYINPUT124), .B1(new_n993), .B2(new_n976), .ZN(new_n995));
  INV_X1    g570(.A(KEYINPUT124), .ZN(new_n996));
  AOI211_X1 g571(.A(new_n996), .B(new_n977), .C1(new_n989), .C2(new_n992), .ZN(new_n997));
  OAI211_X1 g572(.A(new_n985), .B(new_n994), .C1(new_n995), .C2(new_n997), .ZN(new_n998));
  AOI21_X1  g573(.A(G1971), .B1(new_n954), .B2(new_n961), .ZN(new_n999));
  XOR2_X1   g574(.A(KEYINPUT115), .B(G2090), .Z(new_n1000));
  NOR3_X1   g575(.A1(new_n958), .A2(new_n959), .A3(new_n1000), .ZN(new_n1001));
  OAI21_X1  g576(.A(G8), .B1(new_n999), .B2(new_n1001), .ZN(new_n1002));
  NOR2_X1   g577(.A1(G166), .A2(new_n975), .ZN(new_n1003));
  XOR2_X1   g578(.A(new_n1003), .B(KEYINPUT55), .Z(new_n1004));
  NAND2_X1  g579(.A1(new_n1002), .A2(new_n1004), .ZN(new_n1005));
  INV_X1    g580(.A(KEYINPUT116), .ZN(new_n1006));
  NOR2_X1   g581(.A1(new_n1006), .A2(KEYINPUT49), .ZN(new_n1007));
  INV_X1    g582(.A(new_n1007), .ZN(new_n1008));
  AND2_X1   g583(.A1(new_n566), .A2(new_n568), .ZN(new_n1009));
  OAI21_X1  g584(.A(G1981), .B1(new_n1009), .B2(new_n563), .ZN(new_n1010));
  INV_X1    g585(.A(G1981), .ZN(new_n1011));
  NAND3_X1  g586(.A1(new_n564), .A2(new_n1011), .A3(new_n569), .ZN(new_n1012));
  AOI21_X1  g587(.A(new_n1008), .B1(new_n1010), .B2(new_n1012), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n1006), .A2(KEYINPUT49), .ZN(new_n1014));
  NOR3_X1   g589(.A1(new_n1009), .A2(G1981), .A3(new_n563), .ZN(new_n1015));
  AOI21_X1  g590(.A(new_n1011), .B1(new_n564), .B2(new_n569), .ZN(new_n1016));
  OAI21_X1  g591(.A(new_n1014), .B1(new_n1015), .B2(new_n1016), .ZN(new_n1017));
  AOI21_X1  g592(.A(new_n1013), .B1(new_n1017), .B2(new_n1008), .ZN(new_n1018));
  AOI21_X1  g593(.A(new_n975), .B1(new_n956), .B2(new_n922), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n1018), .A2(new_n1019), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n660), .A2(G1976), .ZN(new_n1021));
  AOI21_X1  g596(.A(KEYINPUT52), .B1(G288), .B2(new_n663), .ZN(new_n1022));
  NAND3_X1  g597(.A1(new_n1019), .A2(new_n1021), .A3(new_n1022), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n1020), .A2(new_n1023), .ZN(new_n1024));
  INV_X1    g599(.A(KEYINPUT52), .ZN(new_n1025));
  AOI21_X1  g600(.A(new_n1025), .B1(new_n1019), .B2(new_n1021), .ZN(new_n1026));
  NOR2_X1   g601(.A1(new_n1024), .A2(new_n1026), .ZN(new_n1027));
  INV_X1    g602(.A(new_n1004), .ZN(new_n1028));
  OAI211_X1 g603(.A(new_n1028), .B(G8), .C1(new_n999), .C2(new_n1001), .ZN(new_n1029));
  NAND3_X1  g604(.A1(new_n1005), .A2(new_n1027), .A3(new_n1029), .ZN(new_n1030));
  INV_X1    g605(.A(new_n1030), .ZN(new_n1031));
  AND2_X1   g606(.A1(new_n998), .A2(new_n1031), .ZN(new_n1032));
  AOI21_X1  g607(.A(new_n946), .B1(new_n972), .B2(G171), .ZN(new_n1033));
  OAI21_X1  g608(.A(new_n1033), .B1(G171), .B2(new_n967), .ZN(new_n1034));
  NAND3_X1  g609(.A1(new_n974), .A2(new_n1032), .A3(new_n1034), .ZN(new_n1035));
  INV_X1    g610(.A(KEYINPUT121), .ZN(new_n1036));
  NOR2_X1   g611(.A1(new_n1036), .A2(KEYINPUT59), .ZN(new_n1037));
  INV_X1    g612(.A(new_n1037), .ZN(new_n1038));
  AOI21_X1  g613(.A(new_n539), .B1(new_n1036), .B2(KEYINPUT59), .ZN(new_n1039));
  INV_X1    g614(.A(new_n1039), .ZN(new_n1040));
  NAND3_X1  g615(.A1(new_n954), .A2(new_n928), .A3(new_n961), .ZN(new_n1041));
  INV_X1    g616(.A(KEYINPUT120), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n956), .A2(new_n922), .ZN(new_n1043));
  XOR2_X1   g618(.A(KEYINPUT58), .B(G1341), .Z(new_n1044));
  AOI22_X1  g619(.A1(new_n1041), .A2(new_n1042), .B1(new_n1043), .B2(new_n1044), .ZN(new_n1045));
  NAND4_X1  g620(.A1(new_n954), .A2(new_n961), .A3(KEYINPUT120), .A4(new_n928), .ZN(new_n1046));
  AOI211_X1 g621(.A(new_n1038), .B(new_n1040), .C1(new_n1045), .C2(new_n1046), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n1041), .A2(new_n1042), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n1043), .A2(new_n1044), .ZN(new_n1049));
  NAND3_X1  g624(.A1(new_n1048), .A2(new_n1046), .A3(new_n1049), .ZN(new_n1050));
  AOI21_X1  g625(.A(new_n1037), .B1(new_n1050), .B2(new_n1039), .ZN(new_n1051));
  NOR2_X1   g626(.A1(new_n1047), .A2(new_n1051), .ZN(new_n1052));
  INV_X1    g627(.A(KEYINPUT61), .ZN(new_n1053));
  XNOR2_X1  g628(.A(KEYINPUT56), .B(G2072), .ZN(new_n1054));
  NAND3_X1  g629(.A1(new_n954), .A2(new_n961), .A3(new_n1054), .ZN(new_n1055));
  XOR2_X1   g630(.A(G299), .B(KEYINPUT57), .Z(new_n1056));
  OAI21_X1  g631(.A(new_n741), .B1(new_n958), .B2(new_n959), .ZN(new_n1057));
  AND3_X1   g632(.A1(new_n1055), .A2(new_n1056), .A3(new_n1057), .ZN(new_n1058));
  AOI21_X1  g633(.A(new_n1056), .B1(new_n1055), .B2(new_n1057), .ZN(new_n1059));
  OAI21_X1  g634(.A(new_n1053), .B1(new_n1058), .B2(new_n1059), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n1055), .A2(new_n1057), .ZN(new_n1061));
  INV_X1    g636(.A(new_n1056), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n1061), .A2(new_n1062), .ZN(new_n1063));
  NAND3_X1  g638(.A1(new_n1055), .A2(new_n1056), .A3(new_n1057), .ZN(new_n1064));
  NAND3_X1  g639(.A1(new_n1063), .A2(KEYINPUT61), .A3(new_n1064), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n1060), .A2(new_n1065), .ZN(new_n1066));
  OAI21_X1  g641(.A(KEYINPUT122), .B1(new_n1052), .B2(new_n1066), .ZN(new_n1067));
  AND2_X1   g642(.A1(new_n1060), .A2(new_n1065), .ZN(new_n1068));
  INV_X1    g643(.A(KEYINPUT122), .ZN(new_n1069));
  OAI211_X1 g644(.A(new_n1068), .B(new_n1069), .C1(new_n1051), .C2(new_n1047), .ZN(new_n1070));
  INV_X1    g645(.A(G1348), .ZN(new_n1071));
  OAI21_X1  g646(.A(new_n1071), .B1(new_n958), .B2(new_n959), .ZN(new_n1072));
  NAND3_X1  g647(.A1(new_n956), .A2(new_n926), .A3(new_n922), .ZN(new_n1073));
  AND2_X1   g648(.A1(new_n1072), .A2(new_n1073), .ZN(new_n1074));
  OAI211_X1 g649(.A(KEYINPUT123), .B(new_n583), .C1(new_n1074), .C2(KEYINPUT60), .ZN(new_n1075));
  AND2_X1   g650(.A1(new_n1074), .A2(KEYINPUT60), .ZN(new_n1076));
  INV_X1    g651(.A(KEYINPUT123), .ZN(new_n1077));
  AOI21_X1  g652(.A(KEYINPUT60), .B1(new_n1072), .B2(new_n1073), .ZN(new_n1078));
  OAI21_X1  g653(.A(new_n1077), .B1(new_n1078), .B2(new_n582), .ZN(new_n1079));
  AND3_X1   g654(.A1(new_n1075), .A2(new_n1076), .A3(new_n1079), .ZN(new_n1080));
  AOI21_X1  g655(.A(new_n1076), .B1(new_n1075), .B2(new_n1079), .ZN(new_n1081));
  NOR2_X1   g656(.A1(new_n1080), .A2(new_n1081), .ZN(new_n1082));
  NAND3_X1  g657(.A1(new_n1067), .A2(new_n1070), .A3(new_n1082), .ZN(new_n1083));
  NOR2_X1   g658(.A1(new_n1074), .A2(new_n582), .ZN(new_n1084));
  OAI21_X1  g659(.A(new_n1064), .B1(new_n1084), .B2(new_n1059), .ZN(new_n1085));
  AOI21_X1  g660(.A(new_n1035), .B1(new_n1083), .B2(new_n1085), .ZN(new_n1086));
  AOI211_X1 g661(.A(G1976), .B(G288), .C1(new_n1018), .C2(new_n1019), .ZN(new_n1087));
  OAI21_X1  g662(.A(new_n1019), .B1(new_n1087), .B2(new_n1015), .ZN(new_n1088));
  INV_X1    g663(.A(KEYINPUT117), .ZN(new_n1089));
  OAI21_X1  g664(.A(new_n1089), .B1(new_n1024), .B2(new_n1026), .ZN(new_n1090));
  INV_X1    g665(.A(new_n1026), .ZN(new_n1091));
  NAND4_X1  g666(.A1(new_n1091), .A2(KEYINPUT117), .A3(new_n1023), .A4(new_n1020), .ZN(new_n1092));
  NAND2_X1  g667(.A1(new_n1090), .A2(new_n1092), .ZN(new_n1093));
  INV_X1    g668(.A(new_n1093), .ZN(new_n1094));
  OAI21_X1  g669(.A(new_n1088), .B1(new_n1094), .B2(new_n1029), .ZN(new_n1095));
  AOI21_X1  g670(.A(G1966), .B1(new_n952), .B2(new_n954), .ZN(new_n1096));
  NOR3_X1   g671(.A1(new_n958), .A2(G2084), .A3(new_n959), .ZN(new_n1097));
  OAI211_X1 g672(.A(G8), .B(G168), .C1(new_n1096), .C2(new_n1097), .ZN(new_n1098));
  INV_X1    g673(.A(KEYINPUT63), .ZN(new_n1099));
  NOR2_X1   g674(.A1(new_n1098), .A2(new_n1099), .ZN(new_n1100));
  NAND4_X1  g675(.A1(new_n1100), .A2(new_n1005), .A3(new_n1029), .A4(new_n1093), .ZN(new_n1101));
  AOI211_X1 g676(.A(new_n975), .B(G286), .C1(new_n989), .C2(new_n992), .ZN(new_n1102));
  NAND4_X1  g677(.A1(new_n1005), .A2(new_n1102), .A3(new_n1027), .A4(new_n1029), .ZN(new_n1103));
  AOI22_X1  g678(.A1(new_n1101), .A2(KEYINPUT119), .B1(new_n1099), .B2(new_n1103), .ZN(new_n1104));
  AND2_X1   g679(.A1(new_n1005), .A2(new_n1029), .ZN(new_n1105));
  INV_X1    g680(.A(KEYINPUT119), .ZN(new_n1106));
  NAND4_X1  g681(.A1(new_n1105), .A2(new_n1106), .A3(new_n1093), .A4(new_n1100), .ZN(new_n1107));
  AOI21_X1  g682(.A(new_n1095), .B1(new_n1104), .B2(new_n1107), .ZN(new_n1108));
  OAI21_X1  g683(.A(new_n996), .B1(new_n984), .B2(new_n977), .ZN(new_n1109));
  NAND3_X1  g684(.A1(new_n993), .A2(KEYINPUT124), .A3(new_n976), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n1109), .A2(new_n1110), .ZN(new_n1111));
  INV_X1    g686(.A(KEYINPUT62), .ZN(new_n1112));
  NAND4_X1  g687(.A1(new_n1111), .A2(new_n1112), .A3(new_n985), .A4(new_n994), .ZN(new_n1113));
  NAND4_X1  g688(.A1(new_n1113), .A2(KEYINPUT126), .A3(new_n968), .A4(new_n1031), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n998), .A2(KEYINPUT62), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n1114), .A2(new_n1115), .ZN(new_n1116));
  NAND2_X1  g691(.A1(new_n967), .A2(G171), .ZN(new_n1117));
  NOR2_X1   g692(.A1(new_n1117), .A2(new_n1030), .ZN(new_n1118));
  AOI21_X1  g693(.A(KEYINPUT126), .B1(new_n1118), .B2(new_n1113), .ZN(new_n1119));
  OAI21_X1  g694(.A(new_n1108), .B1(new_n1116), .B2(new_n1119), .ZN(new_n1120));
  OAI21_X1  g695(.A(new_n945), .B1(new_n1086), .B2(new_n1120), .ZN(new_n1121));
  XNOR2_X1  g696(.A(new_n935), .B(KEYINPUT48), .ZN(new_n1122));
  NAND4_X1  g697(.A1(new_n934), .A2(new_n940), .A3(new_n944), .A4(new_n1122), .ZN(new_n1123));
  INV_X1    g698(.A(KEYINPUT47), .ZN(new_n1124));
  NAND2_X1  g699(.A1(new_n931), .A2(KEYINPUT46), .ZN(new_n1125));
  INV_X1    g700(.A(KEYINPUT127), .ZN(new_n1126));
  XNOR2_X1  g701(.A(new_n1125), .B(new_n1126), .ZN(new_n1127));
  OR2_X1    g702(.A1(new_n931), .A2(KEYINPUT46), .ZN(new_n1128));
  INV_X1    g703(.A(new_n927), .ZN(new_n1129));
  OAI21_X1  g704(.A(new_n925), .B1(new_n735), .B2(new_n1129), .ZN(new_n1130));
  AND4_X1   g705(.A1(new_n1124), .A2(new_n1127), .A3(new_n1128), .A4(new_n1130), .ZN(new_n1131));
  AND2_X1   g706(.A1(new_n1130), .A2(new_n1128), .ZN(new_n1132));
  AOI21_X1  g707(.A(new_n1124), .B1(new_n1132), .B2(new_n1127), .ZN(new_n1133));
  OAI21_X1  g708(.A(new_n1123), .B1(new_n1131), .B2(new_n1133), .ZN(new_n1134));
  INV_X1    g709(.A(new_n925), .ZN(new_n1135));
  NAND3_X1  g710(.A1(new_n934), .A2(new_n940), .A3(new_n943), .ZN(new_n1136));
  OR2_X1    g711(.A1(new_n721), .A2(G2067), .ZN(new_n1137));
  AOI21_X1  g712(.A(new_n1135), .B1(new_n1136), .B2(new_n1137), .ZN(new_n1138));
  NOR2_X1   g713(.A1(new_n1134), .A2(new_n1138), .ZN(new_n1139));
  NAND2_X1  g714(.A1(new_n1121), .A2(new_n1139), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g715(.A(G319), .ZN(new_n1142));
  NOR3_X1   g716(.A1(G401), .A2(new_n1142), .A3(G227), .ZN(new_n1143));
  AND2_X1   g717(.A1(new_n656), .A2(new_n1143), .ZN(new_n1144));
  NAND2_X1  g718(.A1(new_n852), .A2(KEYINPUT106), .ZN(new_n1145));
  NAND3_X1  g719(.A1(new_n828), .A2(new_n841), .A3(new_n842), .ZN(new_n1146));
  AOI22_X1  g720(.A1(new_n1145), .A2(new_n1146), .B1(new_n850), .B2(new_n849), .ZN(new_n1147));
  INV_X1    g721(.A(new_n847), .ZN(new_n1148));
  OAI21_X1  g722(.A(new_n853), .B1(new_n1147), .B2(new_n1148), .ZN(new_n1149));
  OAI211_X1 g723(.A(new_n1144), .B(new_n1149), .C1(new_n899), .C2(new_n908), .ZN(G225));
  INV_X1    g724(.A(G225), .ZN(G308));
endmodule


