//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 0 1 1 0 1 0 0 0 0 0 1 1 1 1 0 1 0 0 1 0 1 0 0 1 0 1 1 0 0 1 0 1 1 1 1 0 1 1 0 0 0 1 1 1 1 0 0 1 1 1 0 1 1 1 0 1 1 1 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:14:50 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n617, new_n618, new_n619, new_n620, new_n621, new_n622,
    new_n624, new_n625, new_n626, new_n627, new_n629, new_n630, new_n631,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n688, new_n689, new_n690, new_n691, new_n692,
    new_n693, new_n695, new_n696, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n707, new_n709, new_n710,
    new_n711, new_n712, new_n713, new_n714, new_n715, new_n716, new_n717,
    new_n718, new_n719, new_n720, new_n721, new_n722, new_n723, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n735, new_n736, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n749,
    new_n750, new_n751, new_n752, new_n753, new_n754, new_n755, new_n756,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n789, new_n790, new_n791, new_n793,
    new_n794, new_n795, new_n796, new_n798, new_n799, new_n800, new_n801,
    new_n802, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n823, new_n824,
    new_n825, new_n826, new_n827, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n859, new_n860, new_n862, new_n863, new_n864,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n883, new_n884, new_n885, new_n886, new_n887, new_n889,
    new_n890, new_n891, new_n892, new_n894, new_n895;
  NAND2_X1  g000(.A1(G229gat), .A2(G233gat), .ZN(new_n202));
  XNOR2_X1  g001(.A(G15gat), .B(G22gat), .ZN(new_n203));
  AND2_X1   g002(.A1(new_n203), .A2(KEYINPUT91), .ZN(new_n204));
  NOR2_X1   g003(.A1(new_n203), .A2(KEYINPUT91), .ZN(new_n205));
  OR3_X1    g004(.A1(new_n204), .A2(new_n205), .A3(G1gat), .ZN(new_n206));
  INV_X1    g005(.A(KEYINPUT16), .ZN(new_n207));
  OAI22_X1  g006(.A1(new_n204), .A2(new_n205), .B1(new_n207), .B2(G1gat), .ZN(new_n208));
  INV_X1    g007(.A(KEYINPUT92), .ZN(new_n209));
  NAND2_X1  g008(.A1(new_n209), .A2(G8gat), .ZN(new_n210));
  NAND3_X1  g009(.A1(new_n206), .A2(new_n208), .A3(new_n210), .ZN(new_n211));
  NOR2_X1   g010(.A1(new_n209), .A2(G8gat), .ZN(new_n212));
  XNOR2_X1  g011(.A(new_n211), .B(new_n212), .ZN(new_n213));
  XOR2_X1   g012(.A(G43gat), .B(G50gat), .Z(new_n214));
  INV_X1    g013(.A(KEYINPUT15), .ZN(new_n215));
  OR2_X1    g014(.A1(new_n214), .A2(new_n215), .ZN(new_n216));
  NAND2_X1  g015(.A1(G29gat), .A2(G36gat), .ZN(new_n217));
  INV_X1    g016(.A(KEYINPUT14), .ZN(new_n218));
  INV_X1    g017(.A(G29gat), .ZN(new_n219));
  INV_X1    g018(.A(G36gat), .ZN(new_n220));
  NAND3_X1  g019(.A1(new_n218), .A2(new_n219), .A3(new_n220), .ZN(new_n221));
  OAI21_X1  g020(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n214), .A2(new_n215), .ZN(new_n224));
  NAND4_X1  g023(.A1(new_n216), .A2(new_n217), .A3(new_n223), .A4(new_n224), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n222), .A2(KEYINPUT89), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n226), .A2(new_n221), .ZN(new_n227));
  NAND4_X1  g026(.A1(new_n218), .A2(new_n219), .A3(new_n220), .A4(KEYINPUT89), .ZN(new_n228));
  AOI22_X1  g027(.A1(new_n227), .A2(new_n228), .B1(G29gat), .B2(G36gat), .ZN(new_n229));
  OAI21_X1  g028(.A(new_n225), .B1(new_n229), .B2(new_n216), .ZN(new_n230));
  OR2_X1    g029(.A1(new_n230), .A2(KEYINPUT90), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n230), .A2(KEYINPUT90), .ZN(new_n232));
  AOI21_X1  g031(.A(KEYINPUT17), .B1(new_n231), .B2(new_n232), .ZN(new_n233));
  AND2_X1   g032(.A1(new_n230), .A2(KEYINPUT17), .ZN(new_n234));
  OAI21_X1  g033(.A(new_n213), .B1(new_n233), .B2(new_n234), .ZN(new_n235));
  AND2_X1   g034(.A1(new_n231), .A2(new_n232), .ZN(new_n236));
  INV_X1    g035(.A(new_n213), .ZN(new_n237));
  AND3_X1   g036(.A1(new_n236), .A2(new_n237), .A3(KEYINPUT93), .ZN(new_n238));
  AOI21_X1  g037(.A(KEYINPUT93), .B1(new_n236), .B2(new_n237), .ZN(new_n239));
  OAI211_X1 g038(.A(new_n202), .B(new_n235), .C1(new_n238), .C2(new_n239), .ZN(new_n240));
  NOR2_X1   g039(.A1(KEYINPUT94), .A2(KEYINPUT18), .ZN(new_n241));
  OR2_X1    g040(.A1(new_n240), .A2(new_n241), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n240), .A2(new_n241), .ZN(new_n243));
  OAI22_X1  g042(.A1(new_n238), .A2(new_n239), .B1(new_n237), .B2(new_n236), .ZN(new_n244));
  XOR2_X1   g043(.A(new_n202), .B(KEYINPUT13), .Z(new_n245));
  NAND2_X1  g044(.A1(new_n244), .A2(new_n245), .ZN(new_n246));
  NAND3_X1  g045(.A1(new_n242), .A2(new_n243), .A3(new_n246), .ZN(new_n247));
  XNOR2_X1  g046(.A(G113gat), .B(G141gat), .ZN(new_n248));
  XNOR2_X1  g047(.A(new_n248), .B(KEYINPUT11), .ZN(new_n249));
  INV_X1    g048(.A(G169gat), .ZN(new_n250));
  XNOR2_X1  g049(.A(new_n249), .B(new_n250), .ZN(new_n251));
  XNOR2_X1  g050(.A(new_n251), .B(G197gat), .ZN(new_n252));
  XOR2_X1   g051(.A(KEYINPUT88), .B(KEYINPUT12), .Z(new_n253));
  XNOR2_X1  g052(.A(new_n252), .B(new_n253), .ZN(new_n254));
  INV_X1    g053(.A(new_n254), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n247), .A2(new_n255), .ZN(new_n256));
  NAND4_X1  g055(.A1(new_n242), .A2(new_n243), .A3(new_n254), .A4(new_n246), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  INV_X1    g057(.A(new_n258), .ZN(new_n259));
  INV_X1    g058(.A(KEYINPUT32), .ZN(new_n260));
  XNOR2_X1  g059(.A(G113gat), .B(G120gat), .ZN(new_n261));
  NOR2_X1   g060(.A1(new_n261), .A2(KEYINPUT1), .ZN(new_n262));
  XOR2_X1   g061(.A(G127gat), .B(G134gat), .Z(new_n263));
  XNOR2_X1  g062(.A(new_n262), .B(new_n263), .ZN(new_n264));
  NOR2_X1   g063(.A1(G183gat), .A2(G190gat), .ZN(new_n265));
  INV_X1    g064(.A(new_n265), .ZN(new_n266));
  NAND2_X1  g065(.A1(G183gat), .A2(G190gat), .ZN(new_n267));
  INV_X1    g066(.A(KEYINPUT24), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  NAND3_X1  g068(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n270));
  NAND3_X1  g069(.A1(new_n266), .A2(new_n269), .A3(new_n270), .ZN(new_n271));
  INV_X1    g070(.A(G176gat), .ZN(new_n272));
  NAND3_X1  g071(.A1(new_n250), .A2(new_n272), .A3(KEYINPUT23), .ZN(new_n273));
  INV_X1    g072(.A(KEYINPUT23), .ZN(new_n274));
  OAI21_X1  g073(.A(new_n274), .B1(G169gat), .B2(G176gat), .ZN(new_n275));
  NAND2_X1  g074(.A1(G169gat), .A2(G176gat), .ZN(new_n276));
  NAND4_X1  g075(.A1(new_n271), .A2(new_n273), .A3(new_n275), .A4(new_n276), .ZN(new_n277));
  XNOR2_X1  g076(.A(KEYINPUT64), .B(KEYINPUT25), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n269), .A2(KEYINPUT65), .ZN(new_n279));
  INV_X1    g078(.A(KEYINPUT65), .ZN(new_n280));
  NAND3_X1  g079(.A1(new_n267), .A2(new_n280), .A3(new_n268), .ZN(new_n281));
  NAND4_X1  g080(.A1(new_n279), .A2(new_n266), .A3(new_n270), .A4(new_n281), .ZN(new_n282));
  AND4_X1   g081(.A1(KEYINPUT25), .A2(new_n273), .A3(new_n275), .A4(new_n276), .ZN(new_n283));
  AOI22_X1  g082(.A1(new_n277), .A2(new_n278), .B1(new_n282), .B2(new_n283), .ZN(new_n284));
  NOR2_X1   g083(.A1(G169gat), .A2(G176gat), .ZN(new_n285));
  INV_X1    g084(.A(KEYINPUT26), .ZN(new_n286));
  AOI22_X1  g085(.A1(new_n285), .A2(KEYINPUT67), .B1(new_n276), .B2(new_n286), .ZN(new_n287));
  INV_X1    g086(.A(KEYINPUT67), .ZN(new_n288));
  NOR4_X1   g087(.A1(new_n288), .A2(KEYINPUT26), .A3(G169gat), .A4(G176gat), .ZN(new_n289));
  OAI21_X1  g088(.A(new_n267), .B1(new_n287), .B2(new_n289), .ZN(new_n290));
  NOR2_X1   g089(.A1(KEYINPUT66), .A2(KEYINPUT28), .ZN(new_n291));
  INV_X1    g090(.A(new_n291), .ZN(new_n292));
  XNOR2_X1  g091(.A(KEYINPUT27), .B(G183gat), .ZN(new_n293));
  INV_X1    g092(.A(G190gat), .ZN(new_n294));
  AOI21_X1  g093(.A(new_n292), .B1(new_n293), .B2(new_n294), .ZN(new_n295));
  INV_X1    g094(.A(new_n295), .ZN(new_n296));
  NAND3_X1  g095(.A1(new_n293), .A2(new_n294), .A3(new_n292), .ZN(new_n297));
  AOI21_X1  g096(.A(new_n290), .B1(new_n296), .B2(new_n297), .ZN(new_n298));
  OAI21_X1  g097(.A(new_n264), .B1(new_n284), .B2(new_n298), .ZN(new_n299));
  NAND2_X1  g098(.A1(G227gat), .A2(G233gat), .ZN(new_n300));
  INV_X1    g099(.A(new_n300), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n282), .A2(new_n283), .ZN(new_n302));
  AND3_X1   g101(.A1(new_n266), .A2(new_n269), .A3(new_n270), .ZN(new_n303));
  NAND3_X1  g102(.A1(new_n273), .A2(new_n275), .A3(new_n276), .ZN(new_n304));
  OAI21_X1  g103(.A(new_n278), .B1(new_n303), .B2(new_n304), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n302), .A2(new_n305), .ZN(new_n306));
  INV_X1    g105(.A(new_n287), .ZN(new_n307));
  NAND3_X1  g106(.A1(new_n285), .A2(KEYINPUT67), .A3(new_n286), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  INV_X1    g108(.A(new_n297), .ZN(new_n310));
  OAI211_X1 g109(.A(new_n309), .B(new_n267), .C1(new_n310), .C2(new_n295), .ZN(new_n311));
  OR3_X1    g110(.A1(new_n263), .A2(KEYINPUT1), .A3(new_n261), .ZN(new_n312));
  OAI21_X1  g111(.A(new_n263), .B1(KEYINPUT1), .B2(new_n261), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  NAND3_X1  g113(.A1(new_n306), .A2(new_n311), .A3(new_n314), .ZN(new_n315));
  NAND3_X1  g114(.A1(new_n299), .A2(new_n301), .A3(new_n315), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n316), .A2(KEYINPUT68), .ZN(new_n317));
  INV_X1    g116(.A(KEYINPUT68), .ZN(new_n318));
  NAND4_X1  g117(.A1(new_n299), .A2(new_n318), .A3(new_n315), .A4(new_n301), .ZN(new_n319));
  AOI21_X1  g118(.A(new_n260), .B1(new_n317), .B2(new_n319), .ZN(new_n320));
  XNOR2_X1  g119(.A(G15gat), .B(G43gat), .ZN(new_n321));
  XNOR2_X1  g120(.A(G71gat), .B(G99gat), .ZN(new_n322));
  XNOR2_X1  g121(.A(new_n321), .B(new_n322), .ZN(new_n323));
  INV_X1    g122(.A(KEYINPUT33), .ZN(new_n324));
  OR2_X1    g123(.A1(new_n323), .A2(new_n324), .ZN(new_n325));
  AND3_X1   g124(.A1(new_n320), .A2(KEYINPUT71), .A3(new_n325), .ZN(new_n326));
  AOI21_X1  g125(.A(KEYINPUT71), .B1(new_n320), .B2(new_n325), .ZN(new_n327));
  NOR2_X1   g126(.A1(new_n326), .A2(new_n327), .ZN(new_n328));
  NOR2_X1   g127(.A1(new_n320), .A2(new_n323), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n317), .A2(new_n319), .ZN(new_n330));
  AOI21_X1  g129(.A(KEYINPUT69), .B1(new_n330), .B2(new_n324), .ZN(new_n331));
  INV_X1    g130(.A(KEYINPUT69), .ZN(new_n332));
  AOI211_X1 g131(.A(new_n332), .B(KEYINPUT33), .C1(new_n317), .C2(new_n319), .ZN(new_n333));
  OAI21_X1  g132(.A(new_n329), .B1(new_n331), .B2(new_n333), .ZN(new_n334));
  NAND2_X1  g133(.A1(new_n334), .A2(KEYINPUT70), .ZN(new_n335));
  INV_X1    g134(.A(KEYINPUT70), .ZN(new_n336));
  OAI211_X1 g135(.A(new_n329), .B(new_n336), .C1(new_n331), .C2(new_n333), .ZN(new_n337));
  AOI21_X1  g136(.A(new_n328), .B1(new_n335), .B2(new_n337), .ZN(new_n338));
  AOI21_X1  g137(.A(new_n301), .B1(new_n299), .B2(new_n315), .ZN(new_n339));
  INV_X1    g138(.A(KEYINPUT34), .ZN(new_n340));
  AOI21_X1  g139(.A(new_n340), .B1(new_n300), .B2(KEYINPUT72), .ZN(new_n341));
  XNOR2_X1  g140(.A(new_n341), .B(KEYINPUT73), .ZN(new_n342));
  XOR2_X1   g141(.A(new_n339), .B(new_n342), .Z(new_n343));
  OR2_X1    g142(.A1(new_n338), .A2(new_n343), .ZN(new_n344));
  XNOR2_X1  g143(.A(G78gat), .B(G106gat), .ZN(new_n345));
  INV_X1    g144(.A(new_n345), .ZN(new_n346));
  INV_X1    g145(.A(G22gat), .ZN(new_n347));
  NAND2_X1  g146(.A1(G228gat), .A2(G233gat), .ZN(new_n348));
  XOR2_X1   g147(.A(G197gat), .B(G204gat), .Z(new_n349));
  AOI21_X1  g148(.A(KEYINPUT22), .B1(G211gat), .B2(G218gat), .ZN(new_n350));
  NOR2_X1   g149(.A1(new_n349), .A2(new_n350), .ZN(new_n351));
  XNOR2_X1  g150(.A(G211gat), .B(G218gat), .ZN(new_n352));
  XNOR2_X1  g151(.A(new_n351), .B(new_n352), .ZN(new_n353));
  INV_X1    g152(.A(KEYINPUT29), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  INV_X1    g154(.A(KEYINPUT3), .ZN(new_n356));
  INV_X1    g155(.A(G155gat), .ZN(new_n357));
  INV_X1    g156(.A(G162gat), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n357), .A2(new_n358), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n359), .A2(KEYINPUT76), .ZN(new_n360));
  NAND2_X1  g159(.A1(G155gat), .A2(G162gat), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  INV_X1    g161(.A(KEYINPUT76), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n361), .A2(KEYINPUT2), .ZN(new_n364));
  INV_X1    g163(.A(new_n364), .ZN(new_n365));
  XNOR2_X1  g164(.A(G141gat), .B(G148gat), .ZN(new_n366));
  OAI221_X1 g165(.A(new_n362), .B1(new_n363), .B2(new_n361), .C1(new_n365), .C2(new_n366), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n359), .A2(new_n361), .ZN(new_n368));
  XNOR2_X1  g167(.A(new_n368), .B(KEYINPUT78), .ZN(new_n369));
  INV_X1    g168(.A(G148gat), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n370), .A2(G141gat), .ZN(new_n371));
  XNOR2_X1  g170(.A(KEYINPUT77), .B(G141gat), .ZN(new_n372));
  OAI21_X1  g171(.A(new_n371), .B1(new_n372), .B2(new_n370), .ZN(new_n373));
  NAND3_X1  g172(.A1(new_n369), .A2(new_n364), .A3(new_n373), .ZN(new_n374));
  AOI22_X1  g173(.A1(new_n355), .A2(new_n356), .B1(new_n367), .B2(new_n374), .ZN(new_n375));
  NAND3_X1  g174(.A1(new_n374), .A2(new_n356), .A3(new_n367), .ZN(new_n376));
  AOI21_X1  g175(.A(new_n353), .B1(new_n376), .B2(new_n354), .ZN(new_n377));
  OAI21_X1  g176(.A(new_n348), .B1(new_n375), .B2(new_n377), .ZN(new_n378));
  NOR2_X1   g177(.A1(new_n375), .A2(new_n348), .ZN(new_n379));
  INV_X1    g178(.A(new_n379), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n376), .A2(new_n354), .ZN(new_n381));
  INV_X1    g180(.A(KEYINPUT80), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n381), .A2(new_n382), .ZN(new_n383));
  NAND3_X1  g182(.A1(new_n376), .A2(KEYINPUT80), .A3(new_n354), .ZN(new_n384));
  AOI21_X1  g183(.A(new_n353), .B1(new_n383), .B2(new_n384), .ZN(new_n385));
  OAI211_X1 g184(.A(new_n347), .B(new_n378), .C1(new_n380), .C2(new_n385), .ZN(new_n386));
  INV_X1    g185(.A(new_n386), .ZN(new_n387));
  INV_X1    g186(.A(new_n353), .ZN(new_n388));
  INV_X1    g187(.A(new_n384), .ZN(new_n389));
  AOI21_X1  g188(.A(KEYINPUT80), .B1(new_n376), .B2(new_n354), .ZN(new_n390));
  OAI21_X1  g189(.A(new_n388), .B1(new_n389), .B2(new_n390), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n391), .A2(new_n379), .ZN(new_n392));
  AOI21_X1  g191(.A(new_n347), .B1(new_n392), .B2(new_n378), .ZN(new_n393));
  OAI21_X1  g192(.A(new_n346), .B1(new_n387), .B2(new_n393), .ZN(new_n394));
  OAI21_X1  g193(.A(new_n378), .B1(new_n380), .B2(new_n385), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n395), .A2(G22gat), .ZN(new_n396));
  NAND3_X1  g195(.A1(new_n396), .A2(new_n386), .A3(new_n345), .ZN(new_n397));
  XOR2_X1   g196(.A(KEYINPUT31), .B(G50gat), .Z(new_n398));
  INV_X1    g197(.A(new_n398), .ZN(new_n399));
  NAND3_X1  g198(.A1(new_n394), .A2(new_n397), .A3(new_n399), .ZN(new_n400));
  INV_X1    g199(.A(new_n400), .ZN(new_n401));
  AOI21_X1  g200(.A(new_n399), .B1(new_n394), .B2(new_n397), .ZN(new_n402));
  NOR2_X1   g201(.A1(new_n401), .A2(new_n402), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n335), .A2(new_n337), .ZN(new_n404));
  INV_X1    g203(.A(new_n328), .ZN(new_n405));
  AND4_X1   g204(.A1(KEYINPUT74), .A2(new_n404), .A3(new_n405), .A4(new_n343), .ZN(new_n406));
  AOI21_X1  g205(.A(KEYINPUT74), .B1(new_n338), .B2(new_n343), .ZN(new_n407));
  OAI211_X1 g206(.A(new_n344), .B(new_n403), .C1(new_n406), .C2(new_n407), .ZN(new_n408));
  INV_X1    g207(.A(KEYINPUT6), .ZN(new_n409));
  XNOR2_X1  g208(.A(G1gat), .B(G29gat), .ZN(new_n410));
  XNOR2_X1  g209(.A(new_n410), .B(KEYINPUT0), .ZN(new_n411));
  XNOR2_X1  g210(.A(G57gat), .B(G85gat), .ZN(new_n412));
  XOR2_X1   g211(.A(new_n411), .B(new_n412), .Z(new_n413));
  NAND2_X1  g212(.A1(new_n374), .A2(new_n367), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n414), .A2(KEYINPUT3), .ZN(new_n415));
  NAND3_X1  g214(.A1(new_n415), .A2(new_n376), .A3(new_n314), .ZN(new_n416));
  NAND2_X1  g215(.A1(G225gat), .A2(G233gat), .ZN(new_n417));
  NAND3_X1  g216(.A1(new_n374), .A2(new_n264), .A3(new_n367), .ZN(new_n418));
  AND2_X1   g217(.A1(new_n418), .A2(KEYINPUT4), .ZN(new_n419));
  NOR2_X1   g218(.A1(new_n418), .A2(KEYINPUT4), .ZN(new_n420));
  OAI211_X1 g219(.A(new_n416), .B(new_n417), .C1(new_n419), .C2(new_n420), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n414), .A2(new_n314), .ZN(new_n422));
  AND2_X1   g221(.A1(new_n422), .A2(new_n418), .ZN(new_n423));
  OAI211_X1 g222(.A(new_n421), .B(KEYINPUT5), .C1(new_n417), .C2(new_n423), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n420), .A2(KEYINPUT79), .ZN(new_n425));
  INV_X1    g224(.A(KEYINPUT79), .ZN(new_n426));
  AOI21_X1  g225(.A(new_n426), .B1(new_n418), .B2(KEYINPUT4), .ZN(new_n427));
  OAI21_X1  g226(.A(new_n425), .B1(new_n420), .B2(new_n427), .ZN(new_n428));
  INV_X1    g227(.A(KEYINPUT5), .ZN(new_n429));
  NAND4_X1  g228(.A1(new_n428), .A2(new_n429), .A3(new_n416), .A4(new_n417), .ZN(new_n430));
  AOI211_X1 g229(.A(new_n409), .B(new_n413), .C1(new_n424), .C2(new_n430), .ZN(new_n431));
  AOI21_X1  g230(.A(new_n413), .B1(new_n424), .B2(new_n430), .ZN(new_n432));
  NOR2_X1   g231(.A1(new_n432), .A2(KEYINPUT6), .ZN(new_n433));
  NAND3_X1  g232(.A1(new_n424), .A2(new_n413), .A3(new_n430), .ZN(new_n434));
  AOI21_X1  g233(.A(new_n431), .B1(new_n433), .B2(new_n434), .ZN(new_n435));
  INV_X1    g234(.A(new_n435), .ZN(new_n436));
  XNOR2_X1  g235(.A(G8gat), .B(G36gat), .ZN(new_n437));
  XNOR2_X1  g236(.A(G64gat), .B(G92gat), .ZN(new_n438));
  XNOR2_X1  g237(.A(new_n437), .B(new_n438), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n306), .A2(new_n311), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n440), .A2(new_n354), .ZN(new_n441));
  NAND2_X1  g240(.A1(G226gat), .A2(G233gat), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n441), .A2(new_n442), .ZN(new_n443));
  NAND3_X1  g242(.A1(new_n440), .A2(G226gat), .A3(G233gat), .ZN(new_n444));
  AOI21_X1  g243(.A(new_n388), .B1(new_n443), .B2(new_n444), .ZN(new_n445));
  INV_X1    g244(.A(new_n445), .ZN(new_n446));
  NAND3_X1  g245(.A1(new_n443), .A2(new_n388), .A3(new_n444), .ZN(new_n447));
  AOI21_X1  g246(.A(new_n439), .B1(new_n446), .B2(new_n447), .ZN(new_n448));
  INV_X1    g247(.A(new_n448), .ZN(new_n449));
  INV_X1    g248(.A(KEYINPUT75), .ZN(new_n450));
  INV_X1    g249(.A(KEYINPUT30), .ZN(new_n451));
  NAND3_X1  g250(.A1(new_n449), .A2(new_n450), .A3(new_n451), .ZN(new_n452));
  OAI21_X1  g251(.A(KEYINPUT30), .B1(new_n448), .B2(KEYINPUT75), .ZN(new_n453));
  NAND3_X1  g252(.A1(new_n446), .A2(new_n439), .A3(new_n447), .ZN(new_n454));
  NAND3_X1  g253(.A1(new_n452), .A2(new_n453), .A3(new_n454), .ZN(new_n455));
  INV_X1    g254(.A(new_n455), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n436), .A2(new_n456), .ZN(new_n457));
  OAI21_X1  g256(.A(KEYINPUT35), .B1(new_n408), .B2(new_n457), .ZN(new_n458));
  INV_X1    g257(.A(KEYINPUT86), .ZN(new_n459));
  AOI22_X1  g258(.A1(new_n433), .A2(new_n434), .B1(new_n431), .B2(KEYINPUT84), .ZN(new_n460));
  OR2_X1    g259(.A1(new_n431), .A2(KEYINPUT84), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  INV_X1    g261(.A(KEYINPUT35), .ZN(new_n463));
  NAND3_X1  g262(.A1(new_n462), .A2(new_n463), .A3(new_n456), .ZN(new_n464));
  OAI21_X1  g263(.A(new_n459), .B1(new_n408), .B2(new_n464), .ZN(new_n465));
  NOR2_X1   g264(.A1(new_n338), .A2(new_n343), .ZN(new_n466));
  NAND3_X1  g265(.A1(new_n404), .A2(new_n405), .A3(new_n343), .ZN(new_n467));
  INV_X1    g266(.A(KEYINPUT74), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  NAND3_X1  g268(.A1(new_n338), .A2(KEYINPUT74), .A3(new_n343), .ZN(new_n470));
  AOI21_X1  g269(.A(new_n466), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  AOI211_X1 g270(.A(KEYINPUT35), .B(new_n455), .C1(new_n460), .C2(new_n461), .ZN(new_n472));
  NAND4_X1  g271(.A1(new_n471), .A2(KEYINPUT86), .A3(new_n403), .A4(new_n472), .ZN(new_n473));
  NAND3_X1  g272(.A1(new_n458), .A2(new_n465), .A3(new_n473), .ZN(new_n474));
  OAI21_X1  g273(.A(KEYINPUT81), .B1(new_n401), .B2(new_n402), .ZN(new_n475));
  INV_X1    g274(.A(new_n402), .ZN(new_n476));
  INV_X1    g275(.A(KEYINPUT81), .ZN(new_n477));
  NAND3_X1  g276(.A1(new_n476), .A2(new_n477), .A3(new_n400), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n475), .A2(new_n478), .ZN(new_n479));
  INV_X1    g278(.A(KEYINPUT40), .ZN(new_n480));
  AOI21_X1  g279(.A(new_n417), .B1(new_n428), .B2(new_n416), .ZN(new_n481));
  INV_X1    g280(.A(KEYINPUT39), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  INV_X1    g282(.A(new_n483), .ZN(new_n484));
  NAND3_X1  g283(.A1(new_n422), .A2(new_n418), .A3(new_n417), .ZN(new_n485));
  AOI21_X1  g284(.A(new_n482), .B1(new_n485), .B2(KEYINPUT82), .ZN(new_n486));
  OAI21_X1  g285(.A(new_n486), .B1(KEYINPUT82), .B2(new_n485), .ZN(new_n487));
  OAI21_X1  g286(.A(new_n413), .B1(new_n481), .B2(new_n487), .ZN(new_n488));
  OAI21_X1  g287(.A(new_n480), .B1(new_n484), .B2(new_n488), .ZN(new_n489));
  OR2_X1    g288(.A1(new_n481), .A2(new_n487), .ZN(new_n490));
  NAND4_X1  g289(.A1(new_n490), .A2(new_n483), .A3(KEYINPUT40), .A4(new_n413), .ZN(new_n491));
  INV_X1    g290(.A(new_n432), .ZN(new_n492));
  NAND4_X1  g291(.A1(new_n455), .A2(new_n489), .A3(new_n491), .A4(new_n492), .ZN(new_n493));
  AND3_X1   g292(.A1(new_n493), .A2(new_n476), .A3(new_n400), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n446), .A2(new_n447), .ZN(new_n495));
  INV_X1    g294(.A(KEYINPUT37), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  INV_X1    g296(.A(KEYINPUT38), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  NAND3_X1  g298(.A1(new_n446), .A2(KEYINPUT37), .A3(new_n447), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n500), .A2(new_n439), .ZN(new_n501));
  OAI21_X1  g300(.A(KEYINPUT83), .B1(new_n499), .B2(new_n501), .ZN(new_n502));
  AOI21_X1  g301(.A(KEYINPUT38), .B1(new_n495), .B2(new_n496), .ZN(new_n503));
  INV_X1    g302(.A(KEYINPUT83), .ZN(new_n504));
  NAND4_X1  g303(.A1(new_n503), .A2(new_n504), .A3(new_n439), .A4(new_n500), .ZN(new_n505));
  AND3_X1   g304(.A1(new_n502), .A2(new_n505), .A3(new_n449), .ZN(new_n506));
  INV_X1    g305(.A(KEYINPUT85), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n501), .A2(new_n507), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n508), .A2(new_n497), .ZN(new_n509));
  NOR2_X1   g308(.A1(new_n501), .A2(new_n507), .ZN(new_n510));
  OAI21_X1  g309(.A(KEYINPUT38), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  NAND4_X1  g310(.A1(new_n506), .A2(new_n461), .A3(new_n460), .A4(new_n511), .ZN(new_n512));
  AOI22_X1  g311(.A1(new_n479), .A2(new_n457), .B1(new_n494), .B2(new_n512), .ZN(new_n513));
  NOR2_X1   g312(.A1(new_n471), .A2(KEYINPUT36), .ZN(new_n514));
  OAI21_X1  g313(.A(new_n344), .B1(new_n406), .B2(new_n407), .ZN(new_n515));
  INV_X1    g314(.A(KEYINPUT36), .ZN(new_n516));
  NOR2_X1   g315(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  OAI21_X1  g316(.A(new_n513), .B1(new_n514), .B2(new_n517), .ZN(new_n518));
  NAND2_X1  g317(.A1(new_n474), .A2(new_n518), .ZN(new_n519));
  INV_X1    g318(.A(KEYINPUT87), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  NAND3_X1  g320(.A1(new_n474), .A2(new_n518), .A3(KEYINPUT87), .ZN(new_n522));
  AOI21_X1  g321(.A(new_n259), .B1(new_n521), .B2(new_n522), .ZN(new_n523));
  XOR2_X1   g322(.A(G183gat), .B(G211gat), .Z(new_n524));
  INV_X1    g323(.A(new_n524), .ZN(new_n525));
  INV_X1    g324(.A(KEYINPUT21), .ZN(new_n526));
  NAND2_X1  g325(.A1(G71gat), .A2(G78gat), .ZN(new_n527));
  INV_X1    g326(.A(new_n527), .ZN(new_n528));
  NOR2_X1   g327(.A1(new_n528), .A2(KEYINPUT9), .ZN(new_n529));
  XNOR2_X1  g328(.A(G57gat), .B(G64gat), .ZN(new_n530));
  NOR2_X1   g329(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  NOR2_X1   g330(.A1(G71gat), .A2(G78gat), .ZN(new_n532));
  NOR2_X1   g331(.A1(new_n528), .A2(new_n532), .ZN(new_n533));
  NOR2_X1   g332(.A1(new_n528), .A2(KEYINPUT95), .ZN(new_n534));
  OR3_X1    g333(.A1(new_n531), .A2(new_n533), .A3(new_n534), .ZN(new_n535));
  OAI21_X1  g334(.A(new_n533), .B1(new_n531), .B2(new_n534), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  INV_X1    g336(.A(new_n537), .ZN(new_n538));
  OAI21_X1  g337(.A(new_n213), .B1(new_n526), .B2(new_n538), .ZN(new_n539));
  XNOR2_X1  g338(.A(G127gat), .B(G155gat), .ZN(new_n540));
  XOR2_X1   g339(.A(new_n540), .B(KEYINPUT20), .Z(new_n541));
  INV_X1    g340(.A(new_n541), .ZN(new_n542));
  NAND2_X1  g341(.A1(new_n538), .A2(new_n526), .ZN(new_n543));
  NAND2_X1  g342(.A1(G231gat), .A2(G233gat), .ZN(new_n544));
  XNOR2_X1  g343(.A(new_n543), .B(new_n544), .ZN(new_n545));
  XOR2_X1   g344(.A(KEYINPUT96), .B(KEYINPUT19), .Z(new_n546));
  NAND2_X1  g345(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  INV_X1    g346(.A(new_n547), .ZN(new_n548));
  NOR2_X1   g347(.A1(new_n545), .A2(new_n546), .ZN(new_n549));
  OAI21_X1  g348(.A(new_n542), .B1(new_n548), .B2(new_n549), .ZN(new_n550));
  OR2_X1    g349(.A1(new_n545), .A2(new_n546), .ZN(new_n551));
  NAND3_X1  g350(.A1(new_n551), .A2(new_n541), .A3(new_n547), .ZN(new_n552));
  AOI21_X1  g351(.A(new_n539), .B1(new_n550), .B2(new_n552), .ZN(new_n553));
  INV_X1    g352(.A(new_n553), .ZN(new_n554));
  NAND3_X1  g353(.A1(new_n550), .A2(new_n539), .A3(new_n552), .ZN(new_n555));
  AOI21_X1  g354(.A(new_n525), .B1(new_n554), .B2(new_n555), .ZN(new_n556));
  INV_X1    g355(.A(new_n555), .ZN(new_n557));
  NOR3_X1   g356(.A1(new_n557), .A2(new_n553), .A3(new_n524), .ZN(new_n558));
  NOR2_X1   g357(.A1(new_n556), .A2(new_n558), .ZN(new_n559));
  NAND2_X1  g358(.A1(G99gat), .A2(G106gat), .ZN(new_n560));
  INV_X1    g359(.A(G85gat), .ZN(new_n561));
  INV_X1    g360(.A(G92gat), .ZN(new_n562));
  AOI22_X1  g361(.A1(KEYINPUT8), .A2(new_n560), .B1(new_n561), .B2(new_n562), .ZN(new_n563));
  XNOR2_X1  g362(.A(new_n563), .B(KEYINPUT98), .ZN(new_n564));
  NAND2_X1  g363(.A1(G85gat), .A2(G92gat), .ZN(new_n565));
  XNOR2_X1  g364(.A(new_n565), .B(KEYINPUT7), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n564), .A2(new_n566), .ZN(new_n567));
  XOR2_X1   g366(.A(G99gat), .B(G106gat), .Z(new_n568));
  NAND2_X1  g367(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  INV_X1    g368(.A(KEYINPUT99), .ZN(new_n570));
  NAND2_X1  g369(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  NAND3_X1  g370(.A1(new_n567), .A2(KEYINPUT99), .A3(new_n568), .ZN(new_n572));
  OR2_X1    g371(.A1(new_n567), .A2(new_n568), .ZN(new_n573));
  NAND3_X1  g372(.A1(new_n571), .A2(new_n572), .A3(new_n573), .ZN(new_n574));
  INV_X1    g373(.A(new_n574), .ZN(new_n575));
  AND2_X1   g374(.A1(G232gat), .A2(G233gat), .ZN(new_n576));
  AOI22_X1  g375(.A1(new_n236), .A2(new_n575), .B1(KEYINPUT41), .B2(new_n576), .ZN(new_n577));
  OAI21_X1  g376(.A(new_n574), .B1(new_n233), .B2(new_n234), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  XNOR2_X1  g378(.A(G190gat), .B(G218gat), .ZN(new_n580));
  XNOR2_X1  g379(.A(new_n580), .B(KEYINPUT100), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n579), .A2(new_n581), .ZN(new_n582));
  INV_X1    g381(.A(new_n581), .ZN(new_n583));
  NAND3_X1  g382(.A1(new_n577), .A2(new_n578), .A3(new_n583), .ZN(new_n584));
  NAND3_X1  g383(.A1(new_n582), .A2(KEYINPUT101), .A3(new_n584), .ZN(new_n585));
  NOR2_X1   g384(.A1(new_n576), .A2(KEYINPUT41), .ZN(new_n586));
  XOR2_X1   g385(.A(new_n586), .B(KEYINPUT97), .Z(new_n587));
  XOR2_X1   g386(.A(G134gat), .B(G162gat), .Z(new_n588));
  XNOR2_X1  g387(.A(new_n587), .B(new_n588), .ZN(new_n589));
  INV_X1    g388(.A(new_n589), .ZN(new_n590));
  NAND2_X1  g389(.A1(new_n585), .A2(new_n590), .ZN(new_n591));
  AOI21_X1  g390(.A(KEYINPUT101), .B1(new_n582), .B2(new_n584), .ZN(new_n592));
  XNOR2_X1  g391(.A(new_n591), .B(new_n592), .ZN(new_n593));
  XNOR2_X1  g392(.A(G120gat), .B(G148gat), .ZN(new_n594));
  XNOR2_X1  g393(.A(G176gat), .B(G204gat), .ZN(new_n595));
  XNOR2_X1  g394(.A(new_n594), .B(new_n595), .ZN(new_n596));
  NAND2_X1  g395(.A1(G230gat), .A2(G233gat), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n574), .A2(new_n538), .ZN(new_n598));
  INV_X1    g397(.A(KEYINPUT10), .ZN(new_n599));
  NAND3_X1  g398(.A1(new_n573), .A2(new_n537), .A3(new_n569), .ZN(new_n600));
  AND3_X1   g399(.A1(new_n598), .A2(new_n599), .A3(new_n600), .ZN(new_n601));
  NOR3_X1   g400(.A1(new_n574), .A2(new_n599), .A3(new_n538), .ZN(new_n602));
  OAI21_X1  g401(.A(new_n597), .B1(new_n601), .B2(new_n602), .ZN(new_n603));
  INV_X1    g402(.A(new_n603), .ZN(new_n604));
  AND2_X1   g403(.A1(new_n598), .A2(new_n600), .ZN(new_n605));
  NOR2_X1   g404(.A1(new_n605), .A2(new_n597), .ZN(new_n606));
  OAI21_X1  g405(.A(new_n596), .B1(new_n604), .B2(new_n606), .ZN(new_n607));
  INV_X1    g406(.A(new_n596), .ZN(new_n608));
  OAI211_X1 g407(.A(new_n603), .B(new_n608), .C1(new_n605), .C2(new_n597), .ZN(new_n609));
  NAND2_X1  g408(.A1(new_n607), .A2(new_n609), .ZN(new_n610));
  INV_X1    g409(.A(new_n610), .ZN(new_n611));
  NAND3_X1  g410(.A1(new_n559), .A2(new_n593), .A3(new_n611), .ZN(new_n612));
  INV_X1    g411(.A(new_n612), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n523), .A2(new_n613), .ZN(new_n614));
  NOR2_X1   g413(.A1(new_n614), .A2(new_n436), .ZN(new_n615));
  XOR2_X1   g414(.A(new_n615), .B(G1gat), .Z(G1324gat));
  NAND3_X1  g415(.A1(new_n523), .A2(new_n455), .A3(new_n613), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n617), .A2(G8gat), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n618), .A2(KEYINPUT42), .ZN(new_n619));
  XOR2_X1   g418(.A(KEYINPUT16), .B(G8gat), .Z(new_n620));
  INV_X1    g419(.A(new_n620), .ZN(new_n621));
  NOR2_X1   g420(.A1(new_n617), .A2(new_n621), .ZN(new_n622));
  MUX2_X1   g421(.A(new_n619), .B(KEYINPUT42), .S(new_n622), .Z(G1325gat));
  NOR2_X1   g422(.A1(new_n514), .A2(new_n517), .ZN(new_n624));
  INV_X1    g423(.A(new_n624), .ZN(new_n625));
  OAI21_X1  g424(.A(G15gat), .B1(new_n614), .B2(new_n625), .ZN(new_n626));
  OR2_X1    g425(.A1(new_n515), .A2(G15gat), .ZN(new_n627));
  OAI21_X1  g426(.A(new_n626), .B1(new_n614), .B2(new_n627), .ZN(G1326gat));
  INV_X1    g427(.A(new_n479), .ZN(new_n629));
  NOR2_X1   g428(.A1(new_n614), .A2(new_n629), .ZN(new_n630));
  XOR2_X1   g429(.A(KEYINPUT43), .B(G22gat), .Z(new_n631));
  XNOR2_X1  g430(.A(new_n630), .B(new_n631), .ZN(G1327gat));
  INV_X1    g431(.A(new_n559), .ZN(new_n633));
  NAND2_X1  g432(.A1(new_n633), .A2(new_n611), .ZN(new_n634));
  NOR2_X1   g433(.A1(new_n634), .A2(new_n593), .ZN(new_n635));
  AND3_X1   g434(.A1(new_n474), .A2(KEYINPUT87), .A3(new_n518), .ZN(new_n636));
  AOI21_X1  g435(.A(KEYINPUT87), .B1(new_n474), .B2(new_n518), .ZN(new_n637));
  OAI211_X1 g436(.A(new_n258), .B(new_n635), .C1(new_n636), .C2(new_n637), .ZN(new_n638));
  NOR3_X1   g437(.A1(new_n638), .A2(G29gat), .A3(new_n436), .ZN(new_n639));
  OR2_X1    g438(.A1(new_n639), .A2(KEYINPUT45), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n639), .A2(KEYINPUT45), .ZN(new_n641));
  INV_X1    g440(.A(KEYINPUT44), .ZN(new_n642));
  NOR2_X1   g441(.A1(new_n593), .A2(new_n642), .ZN(new_n643));
  OAI21_X1  g442(.A(new_n643), .B1(new_n636), .B2(new_n637), .ZN(new_n644));
  INV_X1    g443(.A(new_n593), .ZN(new_n645));
  NAND2_X1  g444(.A1(new_n519), .A2(new_n645), .ZN(new_n646));
  NAND2_X1  g445(.A1(new_n646), .A2(new_n642), .ZN(new_n647));
  AND2_X1   g446(.A1(new_n644), .A2(new_n647), .ZN(new_n648));
  NOR2_X1   g447(.A1(new_n634), .A2(new_n259), .ZN(new_n649));
  AND3_X1   g448(.A1(new_n648), .A2(new_n435), .A3(new_n649), .ZN(new_n650));
  OAI211_X1 g449(.A(new_n640), .B(new_n641), .C1(new_n650), .C2(new_n219), .ZN(G1328gat));
  NOR2_X1   g450(.A1(new_n456), .A2(G36gat), .ZN(new_n652));
  INV_X1    g451(.A(new_n652), .ZN(new_n653));
  OAI21_X1  g452(.A(KEYINPUT102), .B1(new_n638), .B2(new_n653), .ZN(new_n654));
  INV_X1    g453(.A(KEYINPUT102), .ZN(new_n655));
  NAND4_X1  g454(.A1(new_n523), .A2(new_n655), .A3(new_n635), .A4(new_n652), .ZN(new_n656));
  INV_X1    g455(.A(KEYINPUT46), .ZN(new_n657));
  NAND3_X1  g456(.A1(new_n654), .A2(new_n656), .A3(new_n657), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n658), .A2(KEYINPUT103), .ZN(new_n659));
  INV_X1    g458(.A(KEYINPUT103), .ZN(new_n660));
  NAND4_X1  g459(.A1(new_n654), .A2(new_n656), .A3(new_n660), .A4(new_n657), .ZN(new_n661));
  NAND2_X1  g460(.A1(new_n659), .A2(new_n661), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n654), .A2(new_n656), .ZN(new_n663));
  NAND4_X1  g462(.A1(new_n644), .A2(new_n455), .A3(new_n647), .A4(new_n649), .ZN(new_n664));
  AOI22_X1  g463(.A1(new_n663), .A2(KEYINPUT46), .B1(G36gat), .B2(new_n664), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n662), .A2(new_n665), .ZN(G1329gat));
  NAND4_X1  g465(.A1(new_n644), .A2(new_n624), .A3(new_n647), .A4(new_n649), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n667), .A2(G43gat), .ZN(new_n668));
  NOR2_X1   g467(.A1(new_n515), .A2(G43gat), .ZN(new_n669));
  NAND3_X1  g468(.A1(new_n523), .A2(new_n635), .A3(new_n669), .ZN(new_n670));
  NAND3_X1  g469(.A1(new_n668), .A2(KEYINPUT47), .A3(new_n670), .ZN(new_n671));
  INV_X1    g470(.A(KEYINPUT105), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n670), .A2(new_n672), .ZN(new_n673));
  INV_X1    g472(.A(new_n638), .ZN(new_n674));
  NAND3_X1  g473(.A1(new_n674), .A2(KEYINPUT105), .A3(new_n669), .ZN(new_n675));
  AOI22_X1  g474(.A1(new_n673), .A2(new_n675), .B1(G43gat), .B2(new_n667), .ZN(new_n676));
  XOR2_X1   g475(.A(KEYINPUT104), .B(KEYINPUT47), .Z(new_n677));
  OAI21_X1  g476(.A(new_n671), .B1(new_n676), .B2(new_n677), .ZN(G1330gat));
  INV_X1    g477(.A(new_n403), .ZN(new_n679));
  NAND4_X1  g478(.A1(new_n644), .A2(new_n679), .A3(new_n647), .A4(new_n649), .ZN(new_n680));
  NAND2_X1  g479(.A1(new_n680), .A2(G50gat), .ZN(new_n681));
  NOR2_X1   g480(.A1(new_n629), .A2(G50gat), .ZN(new_n682));
  NAND2_X1  g481(.A1(new_n674), .A2(new_n682), .ZN(new_n683));
  NAND3_X1  g482(.A1(new_n681), .A2(KEYINPUT48), .A3(new_n683), .ZN(new_n684));
  NAND3_X1  g483(.A1(new_n648), .A2(new_n479), .A3(new_n649), .ZN(new_n685));
  AOI22_X1  g484(.A1(new_n685), .A2(G50gat), .B1(new_n674), .B2(new_n682), .ZN(new_n686));
  OAI21_X1  g485(.A(new_n684), .B1(new_n686), .B2(KEYINPUT48), .ZN(G1331gat));
  NOR4_X1   g486(.A1(new_n633), .A2(new_n645), .A3(new_n258), .A4(new_n611), .ZN(new_n688));
  NAND2_X1  g487(.A1(new_n519), .A2(new_n688), .ZN(new_n689));
  INV_X1    g488(.A(new_n689), .ZN(new_n690));
  INV_X1    g489(.A(KEYINPUT106), .ZN(new_n691));
  XNOR2_X1  g490(.A(new_n435), .B(new_n691), .ZN(new_n692));
  NAND2_X1  g491(.A1(new_n690), .A2(new_n692), .ZN(new_n693));
  XNOR2_X1  g492(.A(new_n693), .B(G57gat), .ZN(G1332gat));
  AOI211_X1 g493(.A(new_n456), .B(new_n689), .C1(KEYINPUT49), .C2(G64gat), .ZN(new_n695));
  NOR2_X1   g494(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n696));
  XNOR2_X1  g495(.A(new_n695), .B(new_n696), .ZN(G1333gat));
  NAND3_X1  g496(.A1(new_n690), .A2(KEYINPUT108), .A3(new_n471), .ZN(new_n698));
  INV_X1    g497(.A(G71gat), .ZN(new_n699));
  INV_X1    g498(.A(KEYINPUT108), .ZN(new_n700));
  OAI21_X1  g499(.A(new_n700), .B1(new_n689), .B2(new_n515), .ZN(new_n701));
  NAND3_X1  g500(.A1(new_n698), .A2(new_n699), .A3(new_n701), .ZN(new_n702));
  NAND4_X1  g501(.A1(new_n519), .A2(G71gat), .A3(new_n624), .A4(new_n688), .ZN(new_n703));
  XNOR2_X1  g502(.A(new_n703), .B(KEYINPUT107), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n702), .A2(new_n704), .ZN(new_n705));
  XNOR2_X1  g504(.A(new_n705), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g505(.A1(new_n690), .A2(new_n479), .ZN(new_n707));
  XNOR2_X1  g506(.A(new_n707), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g507(.A1(new_n559), .A2(new_n258), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n709), .A2(new_n610), .ZN(new_n710));
  XOR2_X1   g509(.A(new_n710), .B(KEYINPUT109), .Z(new_n711));
  NAND2_X1  g510(.A1(new_n648), .A2(new_n711), .ZN(new_n712));
  OAI21_X1  g511(.A(G85gat), .B1(new_n712), .B2(new_n436), .ZN(new_n713));
  AOI21_X1  g512(.A(new_n593), .B1(new_n474), .B2(new_n518), .ZN(new_n714));
  NAND2_X1  g513(.A1(new_n714), .A2(new_n709), .ZN(new_n715));
  INV_X1    g514(.A(KEYINPUT51), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  INV_X1    g516(.A(KEYINPUT110), .ZN(new_n718));
  NAND3_X1  g517(.A1(new_n714), .A2(KEYINPUT51), .A3(new_n709), .ZN(new_n719));
  AND3_X1   g518(.A1(new_n717), .A2(new_n718), .A3(new_n719), .ZN(new_n720));
  AOI21_X1  g519(.A(new_n718), .B1(new_n717), .B2(new_n719), .ZN(new_n721));
  OAI21_X1  g520(.A(new_n610), .B1(new_n720), .B2(new_n721), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n435), .A2(new_n561), .ZN(new_n723));
  OAI21_X1  g522(.A(new_n713), .B1(new_n722), .B2(new_n723), .ZN(G1336gat));
  AOI21_X1  g523(.A(new_n611), .B1(new_n717), .B2(new_n719), .ZN(new_n725));
  NAND3_X1  g524(.A1(new_n725), .A2(new_n562), .A3(new_n455), .ZN(new_n726));
  NAND4_X1  g525(.A1(new_n644), .A2(new_n455), .A3(new_n647), .A4(new_n711), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n727), .A2(G92gat), .ZN(new_n728));
  NAND2_X1  g527(.A1(new_n726), .A2(new_n728), .ZN(new_n729));
  XOR2_X1   g528(.A(KEYINPUT111), .B(KEYINPUT52), .Z(new_n730));
  NAND2_X1  g529(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  INV_X1    g530(.A(new_n730), .ZN(new_n732));
  NAND3_X1  g531(.A1(new_n726), .A2(new_n728), .A3(new_n732), .ZN(new_n733));
  NAND2_X1  g532(.A1(new_n731), .A2(new_n733), .ZN(G1337gat));
  OAI21_X1  g533(.A(G99gat), .B1(new_n712), .B2(new_n625), .ZN(new_n735));
  OR2_X1    g534(.A1(new_n515), .A2(G99gat), .ZN(new_n736));
  OAI21_X1  g535(.A(new_n735), .B1(new_n722), .B2(new_n736), .ZN(G1338gat));
  NAND4_X1  g536(.A1(new_n644), .A2(new_n679), .A3(new_n647), .A4(new_n711), .ZN(new_n738));
  AOI21_X1  g537(.A(KEYINPUT53), .B1(new_n738), .B2(G106gat), .ZN(new_n739));
  NOR2_X1   g538(.A1(new_n403), .A2(G106gat), .ZN(new_n740));
  AND3_X1   g539(.A1(new_n725), .A2(KEYINPUT112), .A3(new_n740), .ZN(new_n741));
  AOI21_X1  g540(.A(KEYINPUT112), .B1(new_n725), .B2(new_n740), .ZN(new_n742));
  OAI21_X1  g541(.A(new_n739), .B1(new_n741), .B2(new_n742), .ZN(new_n743));
  AND2_X1   g542(.A1(new_n725), .A2(new_n740), .ZN(new_n744));
  NAND4_X1  g543(.A1(new_n644), .A2(new_n479), .A3(new_n647), .A4(new_n711), .ZN(new_n745));
  AND2_X1   g544(.A1(new_n745), .A2(G106gat), .ZN(new_n746));
  OAI21_X1  g545(.A(KEYINPUT53), .B1(new_n744), .B2(new_n746), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n743), .A2(new_n747), .ZN(G1339gat));
  INV_X1    g547(.A(KEYINPUT54), .ZN(new_n749));
  AOI21_X1  g548(.A(new_n608), .B1(new_n604), .B2(new_n749), .ZN(new_n750));
  OR3_X1    g549(.A1(new_n601), .A2(new_n602), .A3(new_n597), .ZN(new_n751));
  NAND4_X1  g550(.A1(new_n751), .A2(new_n603), .A3(KEYINPUT113), .A4(KEYINPUT54), .ZN(new_n752));
  AND2_X1   g551(.A1(new_n750), .A2(new_n752), .ZN(new_n753));
  NOR2_X1   g552(.A1(new_n604), .A2(new_n749), .ZN(new_n754));
  AND2_X1   g553(.A1(new_n754), .A2(new_n751), .ZN(new_n755));
  OAI211_X1 g554(.A(new_n753), .B(KEYINPUT55), .C1(new_n755), .C2(KEYINPUT113), .ZN(new_n756));
  INV_X1    g555(.A(KEYINPUT55), .ZN(new_n757));
  AOI21_X1  g556(.A(KEYINPUT113), .B1(new_n754), .B2(new_n751), .ZN(new_n758));
  NAND2_X1  g557(.A1(new_n750), .A2(new_n752), .ZN(new_n759));
  OAI21_X1  g558(.A(new_n757), .B1(new_n758), .B2(new_n759), .ZN(new_n760));
  NAND4_X1  g559(.A1(new_n258), .A2(new_n756), .A3(new_n609), .A4(new_n760), .ZN(new_n761));
  OR2_X1    g560(.A1(new_n238), .A2(new_n239), .ZN(new_n762));
  AOI21_X1  g561(.A(new_n202), .B1(new_n762), .B2(new_n235), .ZN(new_n763));
  NOR2_X1   g562(.A1(new_n244), .A2(new_n245), .ZN(new_n764));
  OAI21_X1  g563(.A(new_n252), .B1(new_n763), .B2(new_n764), .ZN(new_n765));
  NAND3_X1  g564(.A1(new_n257), .A2(new_n765), .A3(new_n610), .ZN(new_n766));
  AND2_X1   g565(.A1(new_n593), .A2(new_n766), .ZN(new_n767));
  AOI21_X1  g566(.A(new_n559), .B1(new_n761), .B2(new_n767), .ZN(new_n768));
  NAND2_X1  g567(.A1(new_n257), .A2(new_n765), .ZN(new_n769));
  NAND2_X1  g568(.A1(new_n769), .A2(KEYINPUT114), .ZN(new_n770));
  INV_X1    g569(.A(KEYINPUT114), .ZN(new_n771));
  NAND3_X1  g570(.A1(new_n257), .A2(new_n765), .A3(new_n771), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n770), .A2(new_n772), .ZN(new_n773));
  NAND3_X1  g572(.A1(new_n756), .A2(new_n609), .A3(new_n760), .ZN(new_n774));
  OAI21_X1  g573(.A(new_n645), .B1(new_n773), .B2(new_n774), .ZN(new_n775));
  AOI22_X1  g574(.A1(new_n768), .A2(new_n775), .B1(new_n259), .B2(new_n613), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n692), .A2(new_n456), .ZN(new_n777));
  NOR2_X1   g576(.A1(new_n776), .A2(new_n777), .ZN(new_n778));
  INV_X1    g577(.A(new_n408), .ZN(new_n779));
  NAND2_X1  g578(.A1(new_n778), .A2(new_n779), .ZN(new_n780));
  XOR2_X1   g579(.A(new_n780), .B(KEYINPUT115), .Z(new_n781));
  INV_X1    g580(.A(G113gat), .ZN(new_n782));
  NAND3_X1  g581(.A1(new_n781), .A2(new_n782), .A3(new_n258), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n629), .A2(new_n471), .ZN(new_n784));
  NOR2_X1   g583(.A1(new_n776), .A2(new_n784), .ZN(new_n785));
  NAND3_X1  g584(.A1(new_n785), .A2(new_n435), .A3(new_n456), .ZN(new_n786));
  OAI21_X1  g585(.A(G113gat), .B1(new_n786), .B2(new_n259), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n783), .A2(new_n787), .ZN(G1340gat));
  INV_X1    g587(.A(G120gat), .ZN(new_n789));
  NAND3_X1  g588(.A1(new_n781), .A2(new_n789), .A3(new_n610), .ZN(new_n790));
  OAI21_X1  g589(.A(G120gat), .B1(new_n786), .B2(new_n611), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n790), .A2(new_n791), .ZN(G1341gat));
  OAI21_X1  g591(.A(G127gat), .B1(new_n786), .B2(new_n633), .ZN(new_n793));
  INV_X1    g592(.A(G127gat), .ZN(new_n794));
  NAND4_X1  g593(.A1(new_n778), .A2(new_n794), .A3(new_n779), .A4(new_n559), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n793), .A2(new_n795), .ZN(new_n796));
  XOR2_X1   g595(.A(new_n796), .B(KEYINPUT116), .Z(G1342gat));
  NOR3_X1   g596(.A1(new_n776), .A2(new_n593), .A3(new_n777), .ZN(new_n798));
  INV_X1    g597(.A(G134gat), .ZN(new_n799));
  NAND3_X1  g598(.A1(new_n798), .A2(new_n799), .A3(new_n779), .ZN(new_n800));
  XOR2_X1   g599(.A(new_n800), .B(KEYINPUT56), .Z(new_n801));
  OAI21_X1  g600(.A(G134gat), .B1(new_n786), .B2(new_n593), .ZN(new_n802));
  NAND2_X1  g601(.A1(new_n801), .A2(new_n802), .ZN(G1343gat));
  NAND2_X1  g602(.A1(new_n768), .A2(new_n775), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n613), .A2(new_n259), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  INV_X1    g605(.A(KEYINPUT57), .ZN(new_n807));
  NAND3_X1  g606(.A1(new_n806), .A2(new_n807), .A3(new_n679), .ZN(new_n808));
  OAI21_X1  g607(.A(KEYINPUT57), .B1(new_n776), .B2(new_n629), .ZN(new_n809));
  NOR3_X1   g608(.A1(new_n624), .A2(new_n436), .A3(new_n455), .ZN(new_n810));
  NAND3_X1  g609(.A1(new_n808), .A2(new_n809), .A3(new_n810), .ZN(new_n811));
  OAI21_X1  g610(.A(new_n372), .B1(new_n811), .B2(new_n259), .ZN(new_n812));
  NOR2_X1   g611(.A1(new_n624), .A2(new_n403), .ZN(new_n813));
  AND2_X1   g612(.A1(new_n778), .A2(new_n813), .ZN(new_n814));
  NOR2_X1   g613(.A1(new_n259), .A2(G141gat), .ZN(new_n815));
  XNOR2_X1  g614(.A(new_n815), .B(KEYINPUT118), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n814), .A2(new_n816), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n812), .A2(new_n817), .ZN(new_n818));
  INV_X1    g617(.A(KEYINPUT58), .ZN(new_n819));
  INV_X1    g618(.A(KEYINPUT117), .ZN(new_n820));
  AOI21_X1  g619(.A(new_n819), .B1(new_n817), .B2(new_n820), .ZN(new_n821));
  XNOR2_X1  g620(.A(new_n818), .B(new_n821), .ZN(G1344gat));
  NAND3_X1  g621(.A1(new_n814), .A2(new_n370), .A3(new_n610), .ZN(new_n823));
  INV_X1    g622(.A(KEYINPUT59), .ZN(new_n824));
  NAND3_X1  g623(.A1(new_n806), .A2(new_n807), .A3(new_n479), .ZN(new_n825));
  OAI21_X1  g624(.A(KEYINPUT57), .B1(new_n776), .B2(new_n403), .ZN(new_n826));
  NAND4_X1  g625(.A1(new_n825), .A2(new_n826), .A3(new_n610), .A4(new_n810), .ZN(new_n827));
  INV_X1    g626(.A(new_n827), .ZN(new_n828));
  AOI21_X1  g627(.A(new_n370), .B1(new_n828), .B2(KEYINPUT119), .ZN(new_n829));
  INV_X1    g628(.A(KEYINPUT119), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n827), .A2(new_n830), .ZN(new_n831));
  AOI21_X1  g630(.A(new_n824), .B1(new_n829), .B2(new_n831), .ZN(new_n832));
  AND3_X1   g631(.A1(new_n808), .A2(new_n809), .A3(new_n810), .ZN(new_n833));
  AOI211_X1 g632(.A(KEYINPUT59), .B(new_n370), .C1(new_n833), .C2(new_n610), .ZN(new_n834));
  OAI21_X1  g633(.A(new_n823), .B1(new_n832), .B2(new_n834), .ZN(G1345gat));
  NAND3_X1  g634(.A1(new_n833), .A2(G155gat), .A3(new_n559), .ZN(new_n836));
  NAND3_X1  g635(.A1(new_n778), .A2(new_n559), .A3(new_n813), .ZN(new_n837));
  AND2_X1   g636(.A1(new_n837), .A2(KEYINPUT120), .ZN(new_n838));
  OAI21_X1  g637(.A(new_n357), .B1(new_n837), .B2(KEYINPUT120), .ZN(new_n839));
  OAI21_X1  g638(.A(new_n836), .B1(new_n838), .B2(new_n839), .ZN(new_n840));
  INV_X1    g639(.A(KEYINPUT121), .ZN(new_n841));
  NAND2_X1  g640(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  OAI211_X1 g641(.A(new_n836), .B(KEYINPUT121), .C1(new_n838), .C2(new_n839), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n842), .A2(new_n843), .ZN(G1346gat));
  NAND2_X1  g643(.A1(new_n833), .A2(new_n645), .ZN(new_n845));
  INV_X1    g644(.A(KEYINPUT122), .ZN(new_n846));
  AOI21_X1  g645(.A(new_n358), .B1(new_n845), .B2(new_n846), .ZN(new_n847));
  OAI21_X1  g646(.A(new_n847), .B1(new_n846), .B2(new_n845), .ZN(new_n848));
  NAND3_X1  g647(.A1(new_n798), .A2(new_n358), .A3(new_n813), .ZN(new_n849));
  NAND2_X1  g648(.A1(new_n848), .A2(new_n849), .ZN(G1347gat));
  NOR2_X1   g649(.A1(new_n692), .A2(new_n456), .ZN(new_n851));
  XNOR2_X1  g650(.A(new_n851), .B(KEYINPUT123), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n785), .A2(new_n852), .ZN(new_n853));
  NOR3_X1   g652(.A1(new_n853), .A2(new_n250), .A3(new_n259), .ZN(new_n854));
  NOR3_X1   g653(.A1(new_n776), .A2(new_n435), .A3(new_n456), .ZN(new_n855));
  AND2_X1   g654(.A1(new_n855), .A2(new_n779), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n856), .A2(new_n258), .ZN(new_n857));
  AOI21_X1  g656(.A(new_n854), .B1(new_n857), .B2(new_n250), .ZN(G1348gat));
  NAND3_X1  g657(.A1(new_n856), .A2(new_n272), .A3(new_n610), .ZN(new_n859));
  OAI21_X1  g658(.A(G176gat), .B1(new_n853), .B2(new_n611), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n859), .A2(new_n860), .ZN(G1349gat));
  NAND3_X1  g660(.A1(new_n856), .A2(new_n293), .A3(new_n559), .ZN(new_n862));
  OAI21_X1  g661(.A(G183gat), .B1(new_n853), .B2(new_n633), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  XNOR2_X1  g663(.A(new_n864), .B(KEYINPUT60), .ZN(G1350gat));
  NAND3_X1  g664(.A1(new_n856), .A2(new_n294), .A3(new_n645), .ZN(new_n866));
  NAND3_X1  g665(.A1(new_n785), .A2(new_n645), .A3(new_n852), .ZN(new_n867));
  INV_X1    g666(.A(KEYINPUT61), .ZN(new_n868));
  AND3_X1   g667(.A1(new_n867), .A2(new_n868), .A3(G190gat), .ZN(new_n869));
  AOI21_X1  g668(.A(new_n868), .B1(new_n867), .B2(G190gat), .ZN(new_n870));
  OAI21_X1  g669(.A(new_n866), .B1(new_n869), .B2(new_n870), .ZN(G1351gat));
  AND2_X1   g670(.A1(new_n825), .A2(new_n826), .ZN(new_n872));
  INV_X1    g671(.A(KEYINPUT125), .ZN(new_n873));
  AND3_X1   g672(.A1(new_n852), .A2(new_n873), .A3(new_n625), .ZN(new_n874));
  AOI21_X1  g673(.A(new_n873), .B1(new_n852), .B2(new_n625), .ZN(new_n875));
  OR2_X1    g674(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  NAND2_X1  g675(.A1(new_n872), .A2(new_n876), .ZN(new_n877));
  NOR2_X1   g676(.A1(new_n877), .A2(new_n259), .ZN(new_n878));
  XOR2_X1   g677(.A(KEYINPUT124), .B(G197gat), .Z(new_n879));
  NAND2_X1  g678(.A1(new_n855), .A2(new_n813), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n258), .A2(new_n879), .ZN(new_n881));
  OAI22_X1  g680(.A1(new_n878), .A2(new_n879), .B1(new_n880), .B2(new_n881), .ZN(G1352gat));
  XOR2_X1   g681(.A(KEYINPUT126), .B(G204gat), .Z(new_n883));
  AND3_X1   g682(.A1(new_n610), .A2(new_n455), .A3(new_n883), .ZN(new_n884));
  NAND4_X1  g683(.A1(new_n806), .A2(new_n436), .A3(new_n813), .A4(new_n884), .ZN(new_n885));
  XOR2_X1   g684(.A(new_n885), .B(KEYINPUT62), .Z(new_n886));
  AND3_X1   g685(.A1(new_n872), .A2(new_n876), .A3(new_n610), .ZN(new_n887));
  OAI21_X1  g686(.A(new_n886), .B1(new_n887), .B2(new_n883), .ZN(G1353gat));
  OR3_X1    g687(.A1(new_n880), .A2(G211gat), .A3(new_n633), .ZN(new_n889));
  NAND3_X1  g688(.A1(new_n872), .A2(new_n876), .A3(new_n559), .ZN(new_n890));
  AND3_X1   g689(.A1(new_n890), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n891));
  AOI21_X1  g690(.A(KEYINPUT63), .B1(new_n890), .B2(G211gat), .ZN(new_n892));
  OAI21_X1  g691(.A(new_n889), .B1(new_n891), .B2(new_n892), .ZN(G1354gat));
  OAI21_X1  g692(.A(G218gat), .B1(new_n877), .B2(new_n593), .ZN(new_n894));
  OR2_X1    g693(.A1(new_n593), .A2(G218gat), .ZN(new_n895));
  OAI21_X1  g694(.A(new_n894), .B1(new_n880), .B2(new_n895), .ZN(G1355gat));
endmodule


