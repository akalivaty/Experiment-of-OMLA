//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 1 1 1 0 1 0 1 1 0 1 0 1 0 1 0 0 1 1 1 1 1 1 1 0 0 1 0 1 1 1 0 1 1 0 0 1 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 0 1 1 1 1 1 1 0 1 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:23:56 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n613, new_n614, new_n615,
    new_n616, new_n618, new_n619, new_n620, new_n621, new_n622, new_n623,
    new_n624, new_n625, new_n626, new_n627, new_n628, new_n629, new_n630,
    new_n632, new_n633, new_n634, new_n635, new_n636, new_n637, new_n638,
    new_n639, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n673, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n684, new_n685,
    new_n686, new_n687, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n697, new_n698, new_n699, new_n700, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n723, new_n724,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n869,
    new_n870, new_n871, new_n872, new_n874, new_n875, new_n876, new_n877,
    new_n878, new_n879, new_n880, new_n881, new_n883, new_n884, new_n885,
    new_n886, new_n887, new_n888, new_n889, new_n890, new_n891, new_n892,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n906, new_n907, new_n908,
    new_n909, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n946, new_n947, new_n948, new_n949, new_n950, new_n951, new_n952,
    new_n953, new_n954, new_n955, new_n956, new_n957;
  XOR2_X1   g000(.A(KEYINPUT9), .B(G234), .Z(new_n187));
  INV_X1    g001(.A(new_n187), .ZN(new_n188));
  OAI21_X1  g002(.A(G221), .B1(new_n188), .B2(G902), .ZN(new_n189));
  XNOR2_X1  g003(.A(new_n189), .B(KEYINPUT80), .ZN(new_n190));
  XOR2_X1   g004(.A(G110), .B(G140), .Z(new_n191));
  INV_X1    g005(.A(G953), .ZN(new_n192));
  AND2_X1   g006(.A1(new_n192), .A2(G227), .ZN(new_n193));
  XNOR2_X1  g007(.A(new_n191), .B(new_n193), .ZN(new_n194));
  INV_X1    g008(.A(new_n194), .ZN(new_n195));
  NOR2_X1   g009(.A1(KEYINPUT81), .A2(KEYINPUT3), .ZN(new_n196));
  INV_X1    g010(.A(G107), .ZN(new_n197));
  NAND3_X1  g011(.A1(new_n196), .A2(G104), .A3(new_n197), .ZN(new_n198));
  INV_X1    g012(.A(G104), .ZN(new_n199));
  AOI22_X1  g013(.A1(new_n199), .A2(G107), .B1(KEYINPUT81), .B2(KEYINPUT3), .ZN(new_n200));
  OAI22_X1  g014(.A1(new_n199), .A2(G107), .B1(KEYINPUT81), .B2(KEYINPUT3), .ZN(new_n201));
  NAND3_X1  g015(.A1(new_n198), .A2(new_n200), .A3(new_n201), .ZN(new_n202));
  INV_X1    g016(.A(KEYINPUT4), .ZN(new_n203));
  NAND3_X1  g017(.A1(new_n202), .A2(new_n203), .A3(G101), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n202), .A2(G101), .ZN(new_n205));
  INV_X1    g019(.A(G101), .ZN(new_n206));
  NAND4_X1  g020(.A1(new_n198), .A2(new_n200), .A3(new_n201), .A4(new_n206), .ZN(new_n207));
  NAND3_X1  g021(.A1(new_n205), .A2(KEYINPUT4), .A3(new_n207), .ZN(new_n208));
  INV_X1    g022(.A(G143), .ZN(new_n209));
  OAI21_X1  g023(.A(KEYINPUT64), .B1(new_n209), .B2(G146), .ZN(new_n210));
  INV_X1    g024(.A(KEYINPUT64), .ZN(new_n211));
  INV_X1    g025(.A(G146), .ZN(new_n212));
  NAND3_X1  g026(.A1(new_n211), .A2(new_n212), .A3(G143), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n209), .A2(G146), .ZN(new_n214));
  NAND3_X1  g028(.A1(new_n210), .A2(new_n213), .A3(new_n214), .ZN(new_n215));
  AND2_X1   g029(.A1(KEYINPUT0), .A2(G128), .ZN(new_n216));
  NOR2_X1   g030(.A1(KEYINPUT0), .A2(G128), .ZN(new_n217));
  NOR2_X1   g031(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n215), .A2(new_n218), .ZN(new_n219));
  INV_X1    g033(.A(KEYINPUT65), .ZN(new_n220));
  AOI21_X1  g034(.A(new_n220), .B1(G143), .B2(new_n212), .ZN(new_n221));
  NOR3_X1   g035(.A1(new_n209), .A2(KEYINPUT65), .A3(G146), .ZN(new_n222));
  OAI211_X1 g036(.A(new_n216), .B(new_n214), .C1(new_n221), .C2(new_n222), .ZN(new_n223));
  INV_X1    g037(.A(KEYINPUT69), .ZN(new_n224));
  AND3_X1   g038(.A1(new_n219), .A2(new_n223), .A3(new_n224), .ZN(new_n225));
  AOI21_X1  g039(.A(new_n224), .B1(new_n219), .B2(new_n223), .ZN(new_n226));
  OAI211_X1 g040(.A(new_n204), .B(new_n208), .C1(new_n225), .C2(new_n226), .ZN(new_n227));
  OAI21_X1  g041(.A(KEYINPUT65), .B1(new_n209), .B2(G146), .ZN(new_n228));
  NAND3_X1  g042(.A1(new_n220), .A2(new_n212), .A3(G143), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  INV_X1    g044(.A(KEYINPUT1), .ZN(new_n231));
  NAND4_X1  g045(.A1(new_n230), .A2(new_n231), .A3(G128), .A4(new_n214), .ZN(new_n232));
  NOR2_X1   g046(.A1(new_n209), .A2(G146), .ZN(new_n233));
  OAI21_X1  g047(.A(G128), .B1(new_n233), .B2(new_n231), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n215), .A2(new_n234), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n232), .A2(new_n235), .ZN(new_n236));
  NOR2_X1   g050(.A1(new_n197), .A2(G104), .ZN(new_n237));
  NOR2_X1   g051(.A1(new_n199), .A2(G107), .ZN(new_n238));
  OAI21_X1  g052(.A(G101), .B1(new_n237), .B2(new_n238), .ZN(new_n239));
  AND2_X1   g053(.A1(new_n207), .A2(new_n239), .ZN(new_n240));
  NAND3_X1  g054(.A1(new_n236), .A2(new_n240), .A3(KEYINPUT10), .ZN(new_n241));
  INV_X1    g055(.A(KEYINPUT83), .ZN(new_n242));
  OAI211_X1 g056(.A(G128), .B(new_n214), .C1(new_n221), .C2(new_n222), .ZN(new_n243));
  AOI22_X1  g057(.A1(new_n228), .A2(new_n229), .B1(new_n209), .B2(G146), .ZN(new_n244));
  INV_X1    g058(.A(G128), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n212), .A2(G143), .ZN(new_n246));
  AOI21_X1  g060(.A(new_n245), .B1(new_n246), .B2(KEYINPUT1), .ZN(new_n247));
  OAI22_X1  g061(.A1(new_n243), .A2(KEYINPUT1), .B1(new_n244), .B2(new_n247), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n248), .A2(new_n240), .ZN(new_n249));
  XNOR2_X1  g063(.A(KEYINPUT82), .B(KEYINPUT10), .ZN(new_n250));
  INV_X1    g064(.A(new_n250), .ZN(new_n251));
  AOI21_X1  g065(.A(new_n242), .B1(new_n249), .B2(new_n251), .ZN(new_n252));
  AOI211_X1 g066(.A(KEYINPUT83), .B(new_n250), .C1(new_n248), .C2(new_n240), .ZN(new_n253));
  OAI211_X1 g067(.A(new_n227), .B(new_n241), .C1(new_n252), .C2(new_n253), .ZN(new_n254));
  INV_X1    g068(.A(KEYINPUT11), .ZN(new_n255));
  INV_X1    g069(.A(G134), .ZN(new_n256));
  OAI21_X1  g070(.A(new_n255), .B1(new_n256), .B2(G137), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n256), .A2(G137), .ZN(new_n258));
  INV_X1    g072(.A(G137), .ZN(new_n259));
  NAND3_X1  g073(.A1(new_n259), .A2(KEYINPUT11), .A3(G134), .ZN(new_n260));
  NAND3_X1  g074(.A1(new_n257), .A2(new_n258), .A3(new_n260), .ZN(new_n261));
  OR2_X1    g075(.A1(new_n261), .A2(G131), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n261), .A2(G131), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n262), .A2(new_n263), .ZN(new_n264));
  XOR2_X1   g078(.A(new_n264), .B(KEYINPUT84), .Z(new_n265));
  INV_X1    g079(.A(new_n265), .ZN(new_n266));
  NOR2_X1   g080(.A1(new_n254), .A2(new_n266), .ZN(new_n267));
  INV_X1    g081(.A(new_n264), .ZN(new_n268));
  INV_X1    g082(.A(new_n241), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n207), .A2(new_n239), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n230), .A2(new_n214), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n271), .A2(new_n234), .ZN(new_n272));
  AOI21_X1  g086(.A(new_n270), .B1(new_n272), .B2(new_n232), .ZN(new_n273));
  OAI21_X1  g087(.A(KEYINPUT83), .B1(new_n273), .B2(new_n250), .ZN(new_n274));
  NAND3_X1  g088(.A1(new_n249), .A2(new_n242), .A3(new_n251), .ZN(new_n275));
  AOI21_X1  g089(.A(new_n269), .B1(new_n274), .B2(new_n275), .ZN(new_n276));
  AOI21_X1  g090(.A(new_n268), .B1(new_n276), .B2(new_n227), .ZN(new_n277));
  OAI21_X1  g091(.A(new_n195), .B1(new_n267), .B2(new_n277), .ZN(new_n278));
  INV_X1    g092(.A(KEYINPUT85), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  OAI211_X1 g094(.A(KEYINPUT85), .B(new_n195), .C1(new_n267), .C2(new_n277), .ZN(new_n281));
  NOR2_X1   g095(.A1(new_n267), .A2(new_n195), .ZN(new_n282));
  NOR2_X1   g096(.A1(new_n236), .A2(new_n240), .ZN(new_n283));
  OAI21_X1  g097(.A(new_n264), .B1(new_n283), .B2(new_n273), .ZN(new_n284));
  XOR2_X1   g098(.A(new_n284), .B(KEYINPUT12), .Z(new_n285));
  NAND2_X1  g099(.A1(new_n282), .A2(new_n285), .ZN(new_n286));
  NAND3_X1  g100(.A1(new_n280), .A2(new_n281), .A3(new_n286), .ZN(new_n287));
  INV_X1    g101(.A(G469), .ZN(new_n288));
  INV_X1    g102(.A(G902), .ZN(new_n289));
  NAND3_X1  g103(.A1(new_n287), .A2(new_n288), .A3(new_n289), .ZN(new_n290));
  INV_X1    g104(.A(new_n277), .ZN(new_n291));
  NAND3_X1  g105(.A1(new_n276), .A2(new_n227), .A3(new_n265), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n285), .A2(new_n292), .ZN(new_n293));
  AOI22_X1  g107(.A1(new_n291), .A2(new_n282), .B1(new_n293), .B2(new_n195), .ZN(new_n294));
  OAI21_X1  g108(.A(G469), .B1(new_n294), .B2(G902), .ZN(new_n295));
  AOI21_X1  g109(.A(new_n190), .B1(new_n290), .B2(new_n295), .ZN(new_n296));
  OAI21_X1  g110(.A(G214), .B1(G237), .B2(G902), .ZN(new_n297));
  INV_X1    g111(.A(new_n297), .ZN(new_n298));
  AND2_X1   g112(.A1(new_n192), .A2(G952), .ZN(new_n299));
  INV_X1    g113(.A(G234), .ZN(new_n300));
  INV_X1    g114(.A(G237), .ZN(new_n301));
  OAI21_X1  g115(.A(new_n299), .B1(new_n300), .B2(new_n301), .ZN(new_n302));
  XOR2_X1   g116(.A(new_n302), .B(KEYINPUT99), .Z(new_n303));
  INV_X1    g117(.A(new_n303), .ZN(new_n304));
  OAI211_X1 g118(.A(G902), .B(G953), .C1(new_n300), .C2(new_n301), .ZN(new_n305));
  XNOR2_X1  g119(.A(new_n305), .B(KEYINPUT100), .ZN(new_n306));
  XNOR2_X1  g120(.A(KEYINPUT21), .B(G898), .ZN(new_n307));
  AOI21_X1  g121(.A(new_n304), .B1(new_n306), .B2(new_n307), .ZN(new_n308));
  XOR2_X1   g122(.A(new_n308), .B(KEYINPUT101), .Z(new_n309));
  INV_X1    g123(.A(new_n309), .ZN(new_n310));
  INV_X1    g124(.A(KEYINPUT5), .ZN(new_n311));
  INV_X1    g125(.A(G119), .ZN(new_n312));
  NAND3_X1  g126(.A1(new_n311), .A2(new_n312), .A3(G116), .ZN(new_n313));
  INV_X1    g127(.A(KEYINPUT68), .ZN(new_n314));
  OAI21_X1  g128(.A(new_n314), .B1(new_n312), .B2(G116), .ZN(new_n315));
  INV_X1    g129(.A(KEYINPUT67), .ZN(new_n316));
  INV_X1    g130(.A(G116), .ZN(new_n317));
  OAI21_X1  g131(.A(new_n316), .B1(new_n317), .B2(G119), .ZN(new_n318));
  NAND3_X1  g132(.A1(new_n317), .A2(KEYINPUT68), .A3(G119), .ZN(new_n319));
  NAND3_X1  g133(.A1(new_n312), .A2(KEYINPUT67), .A3(G116), .ZN(new_n320));
  NAND4_X1  g134(.A1(new_n315), .A2(new_n318), .A3(new_n319), .A4(new_n320), .ZN(new_n321));
  OAI211_X1 g135(.A(G113), .B(new_n313), .C1(new_n321), .C2(new_n311), .ZN(new_n322));
  XNOR2_X1  g136(.A(KEYINPUT2), .B(G113), .ZN(new_n323));
  OR2_X1    g137(.A1(new_n321), .A2(new_n323), .ZN(new_n324));
  AND2_X1   g138(.A1(new_n322), .A2(new_n324), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n325), .A2(new_n240), .ZN(new_n326));
  XOR2_X1   g140(.A(new_n321), .B(new_n323), .Z(new_n327));
  NAND2_X1  g141(.A1(new_n208), .A2(new_n204), .ZN(new_n328));
  OAI21_X1  g142(.A(new_n326), .B1(new_n327), .B2(new_n328), .ZN(new_n329));
  XOR2_X1   g143(.A(G110), .B(G122), .Z(new_n330));
  NAND2_X1  g144(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  INV_X1    g145(.A(new_n330), .ZN(new_n332));
  OAI211_X1 g146(.A(new_n326), .B(new_n332), .C1(new_n327), .C2(new_n328), .ZN(new_n333));
  NAND3_X1  g147(.A1(new_n331), .A2(KEYINPUT6), .A3(new_n333), .ZN(new_n334));
  INV_X1    g148(.A(KEYINPUT6), .ZN(new_n335));
  NAND3_X1  g149(.A1(new_n329), .A2(new_n335), .A3(new_n330), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n219), .A2(new_n223), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n337), .A2(G125), .ZN(new_n338));
  OAI21_X1  g152(.A(new_n338), .B1(G125), .B2(new_n236), .ZN(new_n339));
  INV_X1    g153(.A(G224), .ZN(new_n340));
  NOR2_X1   g154(.A1(new_n340), .A2(G953), .ZN(new_n341));
  XNOR2_X1  g155(.A(new_n339), .B(new_n341), .ZN(new_n342));
  NAND3_X1  g156(.A1(new_n334), .A2(new_n336), .A3(new_n342), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n240), .A2(KEYINPUT86), .ZN(new_n344));
  XOR2_X1   g158(.A(new_n325), .B(new_n344), .Z(new_n345));
  XOR2_X1   g159(.A(new_n330), .B(KEYINPUT8), .Z(new_n346));
  NAND2_X1  g160(.A1(new_n345), .A2(new_n346), .ZN(new_n347));
  INV_X1    g161(.A(KEYINPUT87), .ZN(new_n348));
  INV_X1    g162(.A(new_n341), .ZN(new_n349));
  AOI22_X1  g163(.A1(new_n338), .A2(new_n348), .B1(KEYINPUT7), .B2(new_n349), .ZN(new_n350));
  OR2_X1    g164(.A1(new_n350), .A2(new_n339), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n350), .A2(new_n339), .ZN(new_n352));
  NAND4_X1  g166(.A1(new_n347), .A2(new_n351), .A3(new_n333), .A4(new_n352), .ZN(new_n353));
  NAND3_X1  g167(.A1(new_n343), .A2(new_n353), .A3(new_n289), .ZN(new_n354));
  OAI21_X1  g168(.A(G210), .B1(G237), .B2(G902), .ZN(new_n355));
  XNOR2_X1  g169(.A(new_n355), .B(KEYINPUT89), .ZN(new_n356));
  NAND3_X1  g170(.A1(new_n354), .A2(KEYINPUT88), .A3(new_n356), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n356), .A2(KEYINPUT88), .ZN(new_n358));
  NAND4_X1  g172(.A1(new_n343), .A2(new_n353), .A3(new_n289), .A4(new_n358), .ZN(new_n359));
  AOI211_X1 g173(.A(new_n298), .B(new_n310), .C1(new_n357), .C2(new_n359), .ZN(new_n360));
  INV_X1    g174(.A(KEYINPUT97), .ZN(new_n361));
  INV_X1    g175(.A(KEYINPUT96), .ZN(new_n362));
  INV_X1    g176(.A(G122), .ZN(new_n363));
  OAI21_X1  g177(.A(KEYINPUT94), .B1(new_n363), .B2(G116), .ZN(new_n364));
  INV_X1    g178(.A(KEYINPUT94), .ZN(new_n365));
  NAND3_X1  g179(.A1(new_n365), .A2(new_n317), .A3(G122), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n364), .A2(new_n366), .ZN(new_n367));
  AOI21_X1  g181(.A(new_n362), .B1(new_n367), .B2(KEYINPUT14), .ZN(new_n368));
  INV_X1    g182(.A(KEYINPUT14), .ZN(new_n369));
  AOI211_X1 g183(.A(KEYINPUT96), .B(new_n369), .C1(new_n364), .C2(new_n366), .ZN(new_n370));
  NAND3_X1  g184(.A1(new_n364), .A2(new_n366), .A3(new_n369), .ZN(new_n371));
  OAI21_X1  g185(.A(KEYINPUT93), .B1(new_n317), .B2(G122), .ZN(new_n372));
  INV_X1    g186(.A(KEYINPUT93), .ZN(new_n373));
  NAND3_X1  g187(.A1(new_n373), .A2(new_n363), .A3(G116), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n372), .A2(new_n374), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n371), .A2(new_n375), .ZN(new_n376));
  NOR3_X1   g190(.A1(new_n368), .A2(new_n370), .A3(new_n376), .ZN(new_n377));
  OAI21_X1  g191(.A(new_n361), .B1(new_n377), .B2(new_n197), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n367), .A2(KEYINPUT14), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n379), .A2(KEYINPUT96), .ZN(new_n380));
  NAND3_X1  g194(.A1(new_n367), .A2(new_n362), .A3(KEYINPUT14), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n380), .A2(new_n381), .ZN(new_n382));
  OAI211_X1 g196(.A(KEYINPUT97), .B(G107), .C1(new_n382), .C2(new_n376), .ZN(new_n383));
  NAND3_X1  g197(.A1(new_n375), .A2(new_n367), .A3(new_n197), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n209), .A2(G128), .ZN(new_n385));
  XNOR2_X1  g199(.A(new_n385), .B(KEYINPUT95), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n245), .A2(G143), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  XNOR2_X1  g202(.A(new_n388), .B(G134), .ZN(new_n389));
  NAND4_X1  g203(.A1(new_n378), .A2(new_n383), .A3(new_n384), .A4(new_n389), .ZN(new_n390));
  INV_X1    g204(.A(KEYINPUT13), .ZN(new_n391));
  AOI21_X1  g205(.A(new_n256), .B1(new_n387), .B2(new_n391), .ZN(new_n392));
  XOR2_X1   g206(.A(new_n388), .B(new_n392), .Z(new_n393));
  NAND2_X1  g207(.A1(new_n375), .A2(new_n367), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n394), .A2(G107), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n395), .A2(new_n384), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n393), .A2(new_n396), .ZN(new_n397));
  NAND3_X1  g211(.A1(new_n187), .A2(G217), .A3(new_n192), .ZN(new_n398));
  INV_X1    g212(.A(new_n398), .ZN(new_n399));
  AND3_X1   g213(.A1(new_n390), .A2(new_n397), .A3(new_n399), .ZN(new_n400));
  AOI21_X1  g214(.A(new_n399), .B1(new_n390), .B2(new_n397), .ZN(new_n401));
  OAI211_X1 g215(.A(KEYINPUT98), .B(new_n289), .C1(new_n400), .C2(new_n401), .ZN(new_n402));
  INV_X1    g216(.A(new_n402), .ZN(new_n403));
  INV_X1    g217(.A(G478), .ZN(new_n404));
  NOR2_X1   g218(.A1(new_n404), .A2(KEYINPUT15), .ZN(new_n405));
  INV_X1    g219(.A(new_n405), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n403), .A2(new_n406), .ZN(new_n407));
  OAI21_X1  g221(.A(new_n289), .B1(new_n400), .B2(new_n401), .ZN(new_n408));
  INV_X1    g222(.A(KEYINPUT98), .ZN(new_n409));
  AOI21_X1  g223(.A(new_n405), .B1(new_n408), .B2(new_n409), .ZN(new_n410));
  OAI21_X1  g224(.A(new_n407), .B1(new_n410), .B2(new_n403), .ZN(new_n411));
  NOR2_X1   g225(.A1(G475), .A2(G902), .ZN(new_n412));
  XNOR2_X1  g226(.A(new_n412), .B(KEYINPUT92), .ZN(new_n413));
  INV_X1    g227(.A(G125), .ZN(new_n414));
  INV_X1    g228(.A(G140), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n414), .A2(new_n415), .ZN(new_n416));
  NAND2_X1  g230(.A1(G125), .A2(G140), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n418), .A2(KEYINPUT16), .ZN(new_n419));
  NOR3_X1   g233(.A1(new_n414), .A2(KEYINPUT16), .A3(G140), .ZN(new_n420));
  INV_X1    g234(.A(new_n420), .ZN(new_n421));
  NAND3_X1  g235(.A1(new_n419), .A2(G146), .A3(new_n421), .ZN(new_n422));
  INV_X1    g236(.A(KEYINPUT16), .ZN(new_n423));
  AOI21_X1  g237(.A(new_n423), .B1(new_n416), .B2(new_n417), .ZN(new_n424));
  OAI21_X1  g238(.A(new_n212), .B1(new_n424), .B2(new_n420), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n422), .A2(new_n425), .ZN(new_n426));
  INV_X1    g240(.A(KEYINPUT90), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n426), .A2(new_n427), .ZN(new_n428));
  NAND3_X1  g242(.A1(new_n301), .A2(new_n192), .A3(G214), .ZN(new_n429));
  XNOR2_X1  g243(.A(new_n429), .B(G143), .ZN(new_n430));
  INV_X1    g244(.A(new_n430), .ZN(new_n431));
  NAND3_X1  g245(.A1(new_n431), .A2(KEYINPUT17), .A3(G131), .ZN(new_n432));
  NAND3_X1  g246(.A1(new_n422), .A2(new_n425), .A3(KEYINPUT90), .ZN(new_n433));
  NAND3_X1  g247(.A1(new_n428), .A2(new_n432), .A3(new_n433), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n434), .A2(KEYINPUT91), .ZN(new_n435));
  XNOR2_X1  g249(.A(new_n430), .B(G131), .ZN(new_n436));
  INV_X1    g250(.A(KEYINPUT17), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n436), .A2(new_n437), .ZN(new_n438));
  INV_X1    g252(.A(KEYINPUT91), .ZN(new_n439));
  NAND4_X1  g253(.A1(new_n428), .A2(new_n439), .A3(new_n432), .A4(new_n433), .ZN(new_n440));
  NAND3_X1  g254(.A1(new_n435), .A2(new_n438), .A3(new_n440), .ZN(new_n441));
  XNOR2_X1  g255(.A(G113), .B(G122), .ZN(new_n442));
  XNOR2_X1  g256(.A(new_n442), .B(new_n199), .ZN(new_n443));
  NAND3_X1  g257(.A1(new_n431), .A2(KEYINPUT18), .A3(G131), .ZN(new_n444));
  INV_X1    g258(.A(KEYINPUT18), .ZN(new_n445));
  INV_X1    g259(.A(G131), .ZN(new_n446));
  OAI21_X1  g260(.A(new_n430), .B1(new_n445), .B2(new_n446), .ZN(new_n447));
  XNOR2_X1  g261(.A(new_n418), .B(new_n212), .ZN(new_n448));
  NAND3_X1  g262(.A1(new_n444), .A2(new_n447), .A3(new_n448), .ZN(new_n449));
  NAND3_X1  g263(.A1(new_n441), .A2(new_n443), .A3(new_n449), .ZN(new_n450));
  XOR2_X1   g264(.A(new_n418), .B(KEYINPUT19), .Z(new_n451));
  OAI21_X1  g265(.A(new_n422), .B1(new_n451), .B2(G146), .ZN(new_n452));
  OAI21_X1  g266(.A(new_n449), .B1(new_n452), .B2(new_n436), .ZN(new_n453));
  INV_X1    g267(.A(new_n443), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  AOI21_X1  g269(.A(new_n413), .B1(new_n450), .B2(new_n455), .ZN(new_n456));
  OR2_X1    g270(.A1(new_n456), .A2(KEYINPUT20), .ZN(new_n457));
  AND3_X1   g271(.A1(new_n441), .A2(new_n443), .A3(new_n449), .ZN(new_n458));
  AOI21_X1  g272(.A(new_n443), .B1(new_n441), .B2(new_n449), .ZN(new_n459));
  OAI21_X1  g273(.A(new_n289), .B1(new_n458), .B2(new_n459), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n460), .A2(G475), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n456), .A2(KEYINPUT20), .ZN(new_n462));
  NAND3_X1  g276(.A1(new_n457), .A2(new_n461), .A3(new_n462), .ZN(new_n463));
  NOR2_X1   g277(.A1(new_n411), .A2(new_n463), .ZN(new_n464));
  AND3_X1   g278(.A1(new_n296), .A2(new_n360), .A3(new_n464), .ZN(new_n465));
  XOR2_X1   g279(.A(KEYINPUT26), .B(G101), .Z(new_n466));
  NAND3_X1  g280(.A1(new_n301), .A2(new_n192), .A3(G210), .ZN(new_n467));
  XNOR2_X1  g281(.A(new_n466), .B(new_n467), .ZN(new_n468));
  XNOR2_X1  g282(.A(KEYINPUT71), .B(KEYINPUT27), .ZN(new_n469));
  XNOR2_X1  g283(.A(new_n468), .B(new_n469), .ZN(new_n470));
  XOR2_X1   g284(.A(new_n470), .B(KEYINPUT73), .Z(new_n471));
  INV_X1    g285(.A(new_n471), .ZN(new_n472));
  INV_X1    g286(.A(KEYINPUT28), .ZN(new_n473));
  INV_X1    g287(.A(new_n258), .ZN(new_n474));
  NOR2_X1   g288(.A1(new_n256), .A2(G137), .ZN(new_n475));
  OAI21_X1  g289(.A(G131), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  NAND3_X1  g290(.A1(new_n236), .A2(new_n262), .A3(new_n476), .ZN(new_n477));
  INV_X1    g291(.A(new_n477), .ZN(new_n478));
  OAI21_X1  g292(.A(new_n264), .B1(new_n225), .B2(new_n226), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n479), .A2(KEYINPUT70), .ZN(new_n480));
  INV_X1    g294(.A(KEYINPUT70), .ZN(new_n481));
  OAI211_X1 g295(.A(new_n481), .B(new_n264), .C1(new_n225), .C2(new_n226), .ZN(new_n482));
  AOI21_X1  g296(.A(new_n478), .B1(new_n480), .B2(new_n482), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n483), .A2(new_n327), .ZN(new_n484));
  INV_X1    g298(.A(KEYINPUT66), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n477), .A2(new_n485), .ZN(new_n486));
  NAND3_X1  g300(.A1(new_n264), .A2(new_n223), .A3(new_n219), .ZN(new_n487));
  NAND4_X1  g301(.A1(new_n236), .A2(KEYINPUT66), .A3(new_n262), .A4(new_n476), .ZN(new_n488));
  NAND3_X1  g302(.A1(new_n486), .A2(new_n487), .A3(new_n488), .ZN(new_n489));
  INV_X1    g303(.A(new_n327), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  AOI21_X1  g305(.A(new_n473), .B1(new_n484), .B2(new_n491), .ZN(new_n492));
  INV_X1    g306(.A(new_n492), .ZN(new_n493));
  NAND3_X1  g307(.A1(new_n479), .A2(new_n327), .A3(new_n477), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n494), .A2(new_n473), .ZN(new_n495));
  XOR2_X1   g309(.A(new_n495), .B(KEYINPUT74), .Z(new_n496));
  AOI21_X1  g310(.A(new_n472), .B1(new_n493), .B2(new_n496), .ZN(new_n497));
  INV_X1    g311(.A(new_n497), .ZN(new_n498));
  INV_X1    g312(.A(new_n470), .ZN(new_n499));
  AOI211_X1 g313(.A(new_n490), .B(new_n478), .C1(new_n480), .C2(new_n482), .ZN(new_n500));
  INV_X1    g314(.A(KEYINPUT30), .ZN(new_n501));
  NAND4_X1  g315(.A1(new_n486), .A2(new_n501), .A3(new_n487), .A4(new_n488), .ZN(new_n502));
  OAI21_X1  g316(.A(new_n502), .B1(new_n483), .B2(new_n501), .ZN(new_n503));
  AOI211_X1 g317(.A(new_n499), .B(new_n500), .C1(new_n503), .C2(new_n490), .ZN(new_n504));
  AOI21_X1  g318(.A(KEYINPUT31), .B1(new_n504), .B2(KEYINPUT72), .ZN(new_n505));
  INV_X1    g319(.A(new_n502), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n337), .A2(KEYINPUT69), .ZN(new_n507));
  NAND3_X1  g321(.A1(new_n219), .A2(new_n223), .A3(new_n224), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  AOI21_X1  g323(.A(new_n481), .B1(new_n509), .B2(new_n264), .ZN(new_n510));
  INV_X1    g324(.A(new_n482), .ZN(new_n511));
  OAI21_X1  g325(.A(new_n477), .B1(new_n510), .B2(new_n511), .ZN(new_n512));
  AOI21_X1  g326(.A(new_n506), .B1(new_n512), .B2(KEYINPUT30), .ZN(new_n513));
  OAI211_X1 g327(.A(new_n484), .B(new_n470), .C1(new_n513), .C2(new_n327), .ZN(new_n514));
  INV_X1    g328(.A(KEYINPUT72), .ZN(new_n515));
  INV_X1    g329(.A(KEYINPUT31), .ZN(new_n516));
  NOR3_X1   g330(.A1(new_n514), .A2(new_n515), .A3(new_n516), .ZN(new_n517));
  OAI21_X1  g331(.A(new_n498), .B1(new_n505), .B2(new_n517), .ZN(new_n518));
  NOR2_X1   g332(.A1(G472), .A2(G902), .ZN(new_n519));
  NAND3_X1  g333(.A1(new_n518), .A2(KEYINPUT32), .A3(new_n519), .ZN(new_n520));
  XNOR2_X1  g334(.A(KEYINPUT75), .B(KEYINPUT32), .ZN(new_n521));
  INV_X1    g335(.A(new_n521), .ZN(new_n522));
  OAI21_X1  g336(.A(new_n516), .B1(new_n514), .B2(new_n515), .ZN(new_n523));
  AOI21_X1  g337(.A(new_n500), .B1(new_n503), .B2(new_n490), .ZN(new_n524));
  NAND4_X1  g338(.A1(new_n524), .A2(KEYINPUT72), .A3(KEYINPUT31), .A4(new_n470), .ZN(new_n525));
  AOI21_X1  g339(.A(new_n497), .B1(new_n523), .B2(new_n525), .ZN(new_n526));
  INV_X1    g340(.A(new_n519), .ZN(new_n527));
  OAI21_X1  g341(.A(new_n522), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  XNOR2_X1  g342(.A(new_n495), .B(KEYINPUT74), .ZN(new_n529));
  NOR3_X1   g343(.A1(new_n492), .A2(new_n529), .A3(new_n471), .ZN(new_n530));
  NOR2_X1   g344(.A1(new_n524), .A2(new_n470), .ZN(new_n531));
  NOR3_X1   g345(.A1(new_n530), .A2(new_n531), .A3(KEYINPUT29), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n512), .A2(new_n490), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n533), .A2(new_n484), .ZN(new_n534));
  AOI21_X1  g348(.A(new_n529), .B1(new_n534), .B2(KEYINPUT28), .ZN(new_n535));
  AND2_X1   g349(.A1(new_n470), .A2(KEYINPUT29), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n537), .A2(new_n289), .ZN(new_n538));
  OAI21_X1  g352(.A(G472), .B1(new_n532), .B2(new_n538), .ZN(new_n539));
  NAND3_X1  g353(.A1(new_n520), .A2(new_n528), .A3(new_n539), .ZN(new_n540));
  NOR2_X1   g354(.A1(new_n312), .A2(G128), .ZN(new_n541));
  AND2_X1   g355(.A1(KEYINPUT77), .A2(KEYINPUT23), .ZN(new_n542));
  NOR2_X1   g356(.A1(KEYINPUT77), .A2(KEYINPUT23), .ZN(new_n543));
  OAI21_X1  g357(.A(new_n541), .B1(new_n542), .B2(new_n543), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n312), .A2(G128), .ZN(new_n545));
  OAI211_X1 g359(.A(new_n544), .B(new_n545), .C1(new_n541), .C2(new_n542), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n546), .A2(G110), .ZN(new_n547));
  INV_X1    g361(.A(KEYINPUT78), .ZN(new_n548));
  XNOR2_X1  g362(.A(new_n547), .B(new_n548), .ZN(new_n549));
  XNOR2_X1  g363(.A(new_n541), .B(KEYINPUT76), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n550), .A2(new_n545), .ZN(new_n551));
  XNOR2_X1  g365(.A(KEYINPUT24), .B(G110), .ZN(new_n552));
  OAI211_X1 g366(.A(new_n549), .B(new_n426), .C1(new_n551), .C2(new_n552), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n551), .A2(new_n552), .ZN(new_n554));
  OAI21_X1  g368(.A(new_n554), .B1(G110), .B2(new_n546), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n418), .A2(new_n212), .ZN(new_n556));
  NAND3_X1  g370(.A1(new_n555), .A2(new_n422), .A3(new_n556), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n553), .A2(new_n557), .ZN(new_n558));
  NAND3_X1  g372(.A1(new_n192), .A2(G221), .A3(G234), .ZN(new_n559));
  XNOR2_X1  g373(.A(new_n559), .B(KEYINPUT22), .ZN(new_n560));
  XNOR2_X1  g374(.A(new_n560), .B(G137), .ZN(new_n561));
  INV_X1    g375(.A(new_n561), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n558), .A2(new_n562), .ZN(new_n563));
  NAND3_X1  g377(.A1(new_n553), .A2(new_n557), .A3(new_n561), .ZN(new_n564));
  NAND3_X1  g378(.A1(new_n563), .A2(new_n289), .A3(new_n564), .ZN(new_n565));
  INV_X1    g379(.A(KEYINPUT79), .ZN(new_n566));
  INV_X1    g380(.A(KEYINPUT25), .ZN(new_n567));
  NAND3_X1  g381(.A1(new_n565), .A2(new_n566), .A3(new_n567), .ZN(new_n568));
  INV_X1    g382(.A(G217), .ZN(new_n569));
  AOI21_X1  g383(.A(new_n569), .B1(G234), .B2(new_n289), .ZN(new_n570));
  AND2_X1   g384(.A1(new_n568), .A2(new_n570), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n565), .A2(new_n567), .ZN(new_n572));
  NAND4_X1  g386(.A1(new_n563), .A2(KEYINPUT25), .A3(new_n289), .A4(new_n564), .ZN(new_n573));
  NAND3_X1  g387(.A1(new_n572), .A2(KEYINPUT79), .A3(new_n573), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n571), .A2(new_n574), .ZN(new_n575));
  OR2_X1    g389(.A1(new_n565), .A2(new_n570), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  INV_X1    g391(.A(new_n577), .ZN(new_n578));
  AND3_X1   g392(.A1(new_n465), .A2(new_n540), .A3(new_n578), .ZN(new_n579));
  XNOR2_X1  g393(.A(new_n579), .B(new_n206), .ZN(G3));
  NOR2_X1   g394(.A1(new_n526), .A2(new_n527), .ZN(new_n581));
  OAI21_X1  g395(.A(G472), .B1(new_n526), .B2(G902), .ZN(new_n582));
  AOI21_X1  g396(.A(new_n581), .B1(new_n582), .B2(KEYINPUT102), .ZN(new_n583));
  NOR2_X1   g397(.A1(new_n577), .A2(new_n190), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n518), .A2(new_n289), .ZN(new_n585));
  INV_X1    g399(.A(KEYINPUT102), .ZN(new_n586));
  NAND3_X1  g400(.A1(new_n585), .A2(new_n586), .A3(G472), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n290), .A2(new_n295), .ZN(new_n588));
  NAND4_X1  g402(.A1(new_n583), .A2(new_n584), .A3(new_n587), .A4(new_n588), .ZN(new_n589));
  INV_X1    g403(.A(new_n589), .ZN(new_n590));
  INV_X1    g404(.A(new_n463), .ZN(new_n591));
  INV_X1    g405(.A(new_n356), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n354), .A2(new_n592), .ZN(new_n593));
  NAND4_X1  g407(.A1(new_n343), .A2(new_n353), .A3(new_n289), .A4(new_n356), .ZN(new_n594));
  NAND3_X1  g408(.A1(new_n593), .A2(new_n297), .A3(new_n594), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n390), .A2(new_n397), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n596), .A2(new_n398), .ZN(new_n597));
  NAND3_X1  g411(.A1(new_n390), .A2(new_n397), .A3(new_n399), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n597), .A2(KEYINPUT103), .ZN(new_n600));
  NAND3_X1  g414(.A1(new_n599), .A2(new_n600), .A3(KEYINPUT33), .ZN(new_n601));
  INV_X1    g415(.A(KEYINPUT33), .ZN(new_n602));
  OAI211_X1 g416(.A(new_n597), .B(new_n598), .C1(KEYINPUT103), .C2(new_n602), .ZN(new_n603));
  NAND3_X1  g417(.A1(new_n601), .A2(G478), .A3(new_n603), .ZN(new_n604));
  NAND3_X1  g418(.A1(new_n599), .A2(new_n404), .A3(new_n289), .ZN(new_n605));
  NAND2_X1  g419(.A1(G478), .A2(G902), .ZN(new_n606));
  NAND3_X1  g420(.A1(new_n604), .A2(new_n605), .A3(new_n606), .ZN(new_n607));
  NOR4_X1   g421(.A1(new_n591), .A2(new_n595), .A3(new_n607), .A4(new_n310), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n590), .A2(new_n608), .ZN(new_n609));
  XNOR2_X1  g423(.A(KEYINPUT34), .B(G104), .ZN(new_n610));
  XOR2_X1   g424(.A(new_n610), .B(KEYINPUT104), .Z(new_n611));
  XNOR2_X1  g425(.A(new_n609), .B(new_n611), .ZN(G6));
  INV_X1    g426(.A(new_n411), .ZN(new_n613));
  NOR4_X1   g427(.A1(new_n613), .A2(new_n595), .A3(new_n463), .A4(new_n310), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n590), .A2(new_n614), .ZN(new_n615));
  XOR2_X1   g429(.A(KEYINPUT35), .B(G107), .Z(new_n616));
  XNOR2_X1  g430(.A(new_n615), .B(new_n616), .ZN(G9));
  NAND2_X1  g431(.A1(new_n558), .A2(KEYINPUT105), .ZN(new_n618));
  INV_X1    g432(.A(new_n618), .ZN(new_n619));
  NOR2_X1   g433(.A1(new_n558), .A2(KEYINPUT105), .ZN(new_n620));
  OAI22_X1  g434(.A1(new_n619), .A2(new_n620), .B1(KEYINPUT36), .B2(new_n562), .ZN(new_n621));
  INV_X1    g435(.A(new_n620), .ZN(new_n622));
  NOR2_X1   g436(.A1(new_n562), .A2(KEYINPUT36), .ZN(new_n623));
  NAND3_X1  g437(.A1(new_n622), .A2(new_n623), .A3(new_n618), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n621), .A2(new_n624), .ZN(new_n625));
  NOR2_X1   g439(.A1(new_n570), .A2(G902), .ZN(new_n626));
  INV_X1    g440(.A(new_n626), .ZN(new_n627));
  OAI21_X1  g441(.A(new_n575), .B1(new_n625), .B2(new_n627), .ZN(new_n628));
  NAND4_X1  g442(.A1(new_n465), .A2(new_n583), .A3(new_n587), .A4(new_n628), .ZN(new_n629));
  XOR2_X1   g443(.A(new_n629), .B(KEYINPUT37), .Z(new_n630));
  XNOR2_X1  g444(.A(new_n630), .B(G110), .ZN(G12));
  INV_X1    g445(.A(G900), .ZN(new_n632));
  NAND2_X1  g446(.A1(new_n306), .A2(new_n632), .ZN(new_n633));
  AND2_X1   g447(.A1(new_n633), .A2(KEYINPUT106), .ZN(new_n634));
  NOR2_X1   g448(.A1(new_n633), .A2(KEYINPUT106), .ZN(new_n635));
  OAI21_X1  g449(.A(new_n303), .B1(new_n634), .B2(new_n635), .ZN(new_n636));
  INV_X1    g450(.A(new_n636), .ZN(new_n637));
  NOR4_X1   g451(.A1(new_n613), .A2(new_n595), .A3(new_n463), .A4(new_n637), .ZN(new_n638));
  NAND4_X1  g452(.A1(new_n540), .A2(new_n296), .A3(new_n628), .A4(new_n638), .ZN(new_n639));
  XNOR2_X1  g453(.A(new_n639), .B(G128), .ZN(G30));
  AND2_X1   g454(.A1(new_n520), .A2(new_n528), .ZN(new_n641));
  AOI21_X1  g455(.A(new_n504), .B1(new_n471), .B2(new_n534), .ZN(new_n642));
  OAI21_X1  g456(.A(G472), .B1(new_n642), .B2(G902), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n641), .A2(new_n643), .ZN(new_n644));
  INV_X1    g458(.A(new_n644), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n411), .A2(new_n463), .ZN(new_n646));
  NOR2_X1   g460(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n357), .A2(new_n359), .ZN(new_n648));
  XNOR2_X1  g462(.A(new_n648), .B(KEYINPUT38), .ZN(new_n649));
  XOR2_X1   g463(.A(new_n636), .B(KEYINPUT39), .Z(new_n650));
  INV_X1    g464(.A(new_n650), .ZN(new_n651));
  NAND2_X1  g465(.A1(new_n296), .A2(new_n651), .ZN(new_n652));
  NOR2_X1   g466(.A1(new_n652), .A2(KEYINPUT40), .ZN(new_n653));
  NOR2_X1   g467(.A1(new_n653), .A2(new_n628), .ZN(new_n654));
  AOI21_X1  g468(.A(new_n298), .B1(new_n652), .B2(KEYINPUT40), .ZN(new_n655));
  NAND4_X1  g469(.A1(new_n647), .A2(new_n649), .A3(new_n654), .A4(new_n655), .ZN(new_n656));
  XNOR2_X1  g470(.A(new_n656), .B(G143), .ZN(G45));
  AND2_X1   g471(.A1(new_n540), .A2(new_n296), .ZN(new_n658));
  INV_X1    g472(.A(new_n607), .ZN(new_n659));
  AND3_X1   g473(.A1(new_n593), .A2(new_n297), .A3(new_n594), .ZN(new_n660));
  NAND4_X1  g474(.A1(new_n659), .A2(new_n660), .A3(new_n463), .A4(new_n636), .ZN(new_n661));
  NOR2_X1   g475(.A1(new_n661), .A2(KEYINPUT107), .ZN(new_n662));
  INV_X1    g476(.A(new_n662), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n661), .A2(KEYINPUT107), .ZN(new_n664));
  NAND4_X1  g478(.A1(new_n658), .A2(new_n628), .A3(new_n663), .A4(new_n664), .ZN(new_n665));
  XNOR2_X1  g479(.A(new_n665), .B(G146), .ZN(G48));
  INV_X1    g480(.A(new_n290), .ZN(new_n667));
  AOI21_X1  g481(.A(new_n288), .B1(new_n287), .B2(new_n289), .ZN(new_n668));
  NOR3_X1   g482(.A1(new_n667), .A2(new_n668), .A3(new_n190), .ZN(new_n669));
  NAND4_X1  g483(.A1(new_n540), .A2(new_n608), .A3(new_n578), .A4(new_n669), .ZN(new_n670));
  XNOR2_X1  g484(.A(KEYINPUT41), .B(G113), .ZN(new_n671));
  XNOR2_X1  g485(.A(new_n670), .B(new_n671), .ZN(G15));
  AND4_X1   g486(.A1(new_n540), .A2(new_n578), .A3(new_n614), .A4(new_n669), .ZN(new_n673));
  XNOR2_X1  g487(.A(new_n673), .B(new_n317), .ZN(G18));
  NAND2_X1  g488(.A1(new_n540), .A2(new_n464), .ZN(new_n675));
  NAND4_X1  g489(.A1(new_n669), .A2(new_n628), .A3(new_n309), .A4(new_n660), .ZN(new_n676));
  OAI21_X1  g490(.A(KEYINPUT108), .B1(new_n675), .B2(new_n676), .ZN(new_n677));
  NAND2_X1  g491(.A1(new_n287), .A2(new_n289), .ZN(new_n678));
  NAND2_X1  g492(.A1(new_n678), .A2(G469), .ZN(new_n679));
  INV_X1    g493(.A(new_n190), .ZN(new_n680));
  NAND4_X1  g494(.A1(new_n679), .A2(new_n660), .A3(new_n680), .A4(new_n290), .ZN(new_n681));
  INV_X1    g495(.A(new_n625), .ZN(new_n682));
  AOI22_X1  g496(.A1(new_n682), .A2(new_n626), .B1(new_n571), .B2(new_n574), .ZN(new_n683));
  NOR3_X1   g497(.A1(new_n681), .A2(new_n683), .A3(new_n310), .ZN(new_n684));
  INV_X1    g498(.A(KEYINPUT108), .ZN(new_n685));
  NAND4_X1  g499(.A1(new_n684), .A2(new_n685), .A3(new_n540), .A4(new_n464), .ZN(new_n686));
  NAND2_X1  g500(.A1(new_n677), .A2(new_n686), .ZN(new_n687));
  XNOR2_X1  g501(.A(new_n687), .B(G119), .ZN(G21));
  NOR4_X1   g502(.A1(new_n646), .A2(new_n667), .A3(new_n668), .A4(new_n190), .ZN(new_n689));
  NAND2_X1  g503(.A1(new_n523), .A2(new_n525), .ZN(new_n690));
  OR2_X1    g504(.A1(new_n535), .A2(new_n472), .ZN(new_n691));
  AOI21_X1  g505(.A(new_n527), .B1(new_n690), .B2(new_n691), .ZN(new_n692));
  AOI21_X1  g506(.A(new_n692), .B1(new_n585), .B2(G472), .ZN(new_n693));
  NOR2_X1   g507(.A1(new_n595), .A2(new_n310), .ZN(new_n694));
  NAND4_X1  g508(.A1(new_n689), .A2(new_n693), .A3(new_n578), .A4(new_n694), .ZN(new_n695));
  XNOR2_X1  g509(.A(new_n695), .B(G122), .ZN(G24));
  NOR2_X1   g510(.A1(new_n681), .A2(new_n683), .ZN(new_n697));
  NAND2_X1  g511(.A1(new_n659), .A2(new_n463), .ZN(new_n698));
  NOR2_X1   g512(.A1(new_n698), .A2(new_n637), .ZN(new_n699));
  NAND3_X1  g513(.A1(new_n697), .A2(new_n699), .A3(new_n693), .ZN(new_n700));
  XNOR2_X1  g514(.A(new_n700), .B(G125), .ZN(G27));
  INV_X1    g515(.A(KEYINPUT32), .ZN(new_n702));
  OAI21_X1  g516(.A(new_n702), .B1(new_n526), .B2(new_n527), .ZN(new_n703));
  NAND3_X1  g517(.A1(new_n520), .A2(new_n703), .A3(new_n539), .ZN(new_n704));
  NAND3_X1  g518(.A1(new_n704), .A2(new_n699), .A3(new_n578), .ZN(new_n705));
  AND3_X1   g519(.A1(new_n357), .A2(new_n359), .A3(new_n297), .ZN(new_n706));
  NAND3_X1  g520(.A1(new_n588), .A2(new_n706), .A3(new_n680), .ZN(new_n707));
  NAND2_X1  g521(.A1(new_n707), .A2(KEYINPUT109), .ZN(new_n708));
  INV_X1    g522(.A(KEYINPUT109), .ZN(new_n709));
  NAND3_X1  g523(.A1(new_n296), .A2(new_n709), .A3(new_n706), .ZN(new_n710));
  NAND2_X1  g524(.A1(new_n708), .A2(new_n710), .ZN(new_n711));
  OAI21_X1  g525(.A(KEYINPUT42), .B1(new_n705), .B2(new_n711), .ZN(new_n712));
  AND2_X1   g526(.A1(new_n540), .A2(new_n578), .ZN(new_n713));
  AND4_X1   g527(.A1(new_n709), .A2(new_n588), .A3(new_n680), .A4(new_n706), .ZN(new_n714));
  AOI21_X1  g528(.A(new_n709), .B1(new_n296), .B2(new_n706), .ZN(new_n715));
  NOR2_X1   g529(.A1(new_n714), .A2(new_n715), .ZN(new_n716));
  NOR2_X1   g530(.A1(new_n591), .A2(new_n607), .ZN(new_n717));
  NAND2_X1  g531(.A1(new_n717), .A2(new_n636), .ZN(new_n718));
  NOR2_X1   g532(.A1(new_n718), .A2(KEYINPUT42), .ZN(new_n719));
  NAND3_X1  g533(.A1(new_n713), .A2(new_n716), .A3(new_n719), .ZN(new_n720));
  NAND2_X1  g534(.A1(new_n712), .A2(new_n720), .ZN(new_n721));
  XNOR2_X1  g535(.A(new_n721), .B(new_n446), .ZN(G33));
  NOR3_X1   g536(.A1(new_n613), .A2(new_n463), .A3(new_n637), .ZN(new_n723));
  NAND3_X1  g537(.A1(new_n713), .A2(new_n723), .A3(new_n716), .ZN(new_n724));
  XNOR2_X1  g538(.A(new_n724), .B(G134), .ZN(G36));
  AOI21_X1  g539(.A(new_n683), .B1(new_n583), .B2(new_n587), .ZN(new_n726));
  XOR2_X1   g540(.A(new_n726), .B(KEYINPUT112), .Z(new_n727));
  NOR3_X1   g541(.A1(new_n607), .A2(new_n463), .A3(KEYINPUT43), .ZN(new_n728));
  XNOR2_X1  g542(.A(new_n463), .B(KEYINPUT111), .ZN(new_n729));
  NAND2_X1  g543(.A1(new_n729), .A2(new_n659), .ZN(new_n730));
  AOI21_X1  g544(.A(new_n728), .B1(new_n730), .B2(KEYINPUT43), .ZN(new_n731));
  NAND2_X1  g545(.A1(new_n727), .A2(new_n731), .ZN(new_n732));
  INV_X1    g546(.A(KEYINPUT44), .ZN(new_n733));
  NAND2_X1  g547(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  OR2_X1    g548(.A1(new_n294), .A2(KEYINPUT45), .ZN(new_n735));
  NAND2_X1  g549(.A1(new_n294), .A2(KEYINPUT45), .ZN(new_n736));
  NAND3_X1  g550(.A1(new_n735), .A2(G469), .A3(new_n736), .ZN(new_n737));
  NAND2_X1  g551(.A1(G469), .A2(G902), .ZN(new_n738));
  NAND2_X1  g552(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  INV_X1    g553(.A(KEYINPUT46), .ZN(new_n740));
  AOI21_X1  g554(.A(new_n667), .B1(new_n739), .B2(new_n740), .ZN(new_n741));
  OAI21_X1  g555(.A(new_n741), .B1(new_n740), .B2(new_n739), .ZN(new_n742));
  NAND2_X1  g556(.A1(new_n742), .A2(new_n680), .ZN(new_n743));
  INV_X1    g557(.A(new_n743), .ZN(new_n744));
  NAND3_X1  g558(.A1(new_n744), .A2(KEYINPUT110), .A3(new_n651), .ZN(new_n745));
  INV_X1    g559(.A(KEYINPUT110), .ZN(new_n746));
  OAI21_X1  g560(.A(new_n746), .B1(new_n743), .B2(new_n650), .ZN(new_n747));
  AND2_X1   g561(.A1(new_n745), .A2(new_n747), .ZN(new_n748));
  NAND3_X1  g562(.A1(new_n727), .A2(KEYINPUT44), .A3(new_n731), .ZN(new_n749));
  NAND4_X1  g563(.A1(new_n734), .A2(new_n748), .A3(new_n706), .A4(new_n749), .ZN(new_n750));
  XNOR2_X1  g564(.A(new_n750), .B(KEYINPUT113), .ZN(new_n751));
  XNOR2_X1  g565(.A(new_n751), .B(G137), .ZN(G39));
  NAND2_X1  g566(.A1(new_n744), .A2(KEYINPUT47), .ZN(new_n753));
  INV_X1    g567(.A(KEYINPUT47), .ZN(new_n754));
  NAND2_X1  g568(.A1(new_n743), .A2(new_n754), .ZN(new_n755));
  AOI21_X1  g569(.A(new_n540), .B1(new_n753), .B2(new_n755), .ZN(new_n756));
  NAND4_X1  g570(.A1(new_n756), .A2(new_n577), .A3(new_n699), .A4(new_n706), .ZN(new_n757));
  XNOR2_X1  g571(.A(new_n757), .B(G140), .ZN(G42));
  AND2_X1   g572(.A1(new_n731), .A2(new_n304), .ZN(new_n759));
  NAND2_X1  g573(.A1(new_n669), .A2(new_n706), .ZN(new_n760));
  INV_X1    g574(.A(new_n760), .ZN(new_n761));
  AND4_X1   g575(.A1(new_n628), .A2(new_n759), .A3(new_n693), .A4(new_n761), .ZN(new_n762));
  NAND4_X1  g576(.A1(new_n645), .A2(new_n578), .A3(new_n304), .A4(new_n761), .ZN(new_n763));
  NOR3_X1   g577(.A1(new_n763), .A2(new_n463), .A3(new_n659), .ZN(new_n764));
  NOR2_X1   g578(.A1(new_n762), .A2(new_n764), .ZN(new_n765));
  INV_X1    g579(.A(new_n669), .ZN(new_n766));
  NOR3_X1   g580(.A1(new_n766), .A2(new_n649), .A3(new_n297), .ZN(new_n767));
  XOR2_X1   g581(.A(new_n767), .B(KEYINPUT117), .Z(new_n768));
  AND2_X1   g582(.A1(new_n693), .A2(new_n578), .ZN(new_n769));
  NAND3_X1  g583(.A1(new_n768), .A2(new_n769), .A3(new_n759), .ZN(new_n770));
  NAND2_X1  g584(.A1(new_n770), .A2(KEYINPUT50), .ZN(new_n771));
  NOR2_X1   g585(.A1(new_n667), .A2(new_n668), .ZN(new_n772));
  NAND2_X1  g586(.A1(new_n772), .A2(new_n190), .ZN(new_n773));
  NAND3_X1  g587(.A1(new_n753), .A2(new_n755), .A3(new_n773), .ZN(new_n774));
  INV_X1    g588(.A(KEYINPUT50), .ZN(new_n775));
  AOI22_X1  g589(.A1(new_n774), .A2(new_n706), .B1(new_n775), .B2(new_n768), .ZN(new_n776));
  NAND2_X1  g590(.A1(new_n759), .A2(new_n769), .ZN(new_n777));
  OAI211_X1 g591(.A(new_n765), .B(new_n771), .C1(new_n776), .C2(new_n777), .ZN(new_n778));
  XNOR2_X1  g592(.A(new_n778), .B(KEYINPUT51), .ZN(new_n779));
  AND2_X1   g593(.A1(new_n704), .A2(new_n578), .ZN(new_n780));
  NAND3_X1  g594(.A1(new_n759), .A2(new_n780), .A3(new_n761), .ZN(new_n781));
  XNOR2_X1  g595(.A(new_n781), .B(KEYINPUT48), .ZN(new_n782));
  OR2_X1    g596(.A1(new_n763), .A2(new_n698), .ZN(new_n783));
  OR2_X1    g597(.A1(new_n777), .A2(new_n681), .ZN(new_n784));
  NAND4_X1  g598(.A1(new_n782), .A2(new_n299), .A3(new_n783), .A4(new_n784), .ZN(new_n785));
  XOR2_X1   g599(.A(new_n785), .B(KEYINPUT118), .Z(new_n786));
  NAND2_X1  g600(.A1(new_n779), .A2(new_n786), .ZN(new_n787));
  INV_X1    g601(.A(KEYINPUT116), .ZN(new_n788));
  INV_X1    g602(.A(KEYINPUT53), .ZN(new_n789));
  NAND3_X1  g603(.A1(new_n712), .A2(new_n720), .A3(new_n724), .ZN(new_n790));
  NAND4_X1  g604(.A1(new_n708), .A2(new_n693), .A3(new_n699), .A4(new_n710), .ZN(new_n791));
  NAND2_X1  g605(.A1(new_n411), .A2(KEYINPUT114), .ZN(new_n792));
  INV_X1    g606(.A(KEYINPUT114), .ZN(new_n793));
  OAI211_X1 g607(.A(new_n407), .B(new_n793), .C1(new_n403), .C2(new_n410), .ZN(new_n794));
  AND4_X1   g608(.A1(new_n591), .A2(new_n792), .A3(new_n636), .A4(new_n794), .ZN(new_n795));
  NAND4_X1  g609(.A1(new_n540), .A2(new_n795), .A3(new_n296), .A4(new_n706), .ZN(new_n796));
  AOI21_X1  g610(.A(new_n683), .B1(new_n791), .B2(new_n796), .ZN(new_n797));
  NOR2_X1   g611(.A1(new_n790), .A2(new_n797), .ZN(new_n798));
  INV_X1    g612(.A(new_n673), .ZN(new_n799));
  AND2_X1   g613(.A1(new_n695), .A2(new_n670), .ZN(new_n800));
  AND3_X1   g614(.A1(new_n687), .A2(new_n799), .A3(new_n800), .ZN(new_n801));
  INV_X1    g615(.A(new_n579), .ZN(new_n802));
  AOI21_X1  g616(.A(new_n463), .B1(new_n792), .B2(new_n794), .ZN(new_n803));
  INV_X1    g617(.A(KEYINPUT115), .ZN(new_n804));
  NAND2_X1  g618(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  INV_X1    g619(.A(new_n805), .ZN(new_n806));
  OAI21_X1  g620(.A(new_n698), .B1(new_n803), .B2(new_n804), .ZN(new_n807));
  OAI21_X1  g621(.A(new_n360), .B1(new_n806), .B2(new_n807), .ZN(new_n808));
  OAI211_X1 g622(.A(new_n802), .B(new_n629), .C1(new_n808), .C2(new_n589), .ZN(new_n809));
  INV_X1    g623(.A(new_n809), .ZN(new_n810));
  NAND3_X1  g624(.A1(new_n798), .A2(new_n801), .A3(new_n810), .ZN(new_n811));
  NAND4_X1  g625(.A1(new_n664), .A2(new_n540), .A3(new_n296), .A4(new_n628), .ZN(new_n812));
  OAI211_X1 g626(.A(new_n639), .B(new_n700), .C1(new_n812), .C2(new_n662), .ZN(new_n813));
  NAND3_X1  g627(.A1(new_n660), .A2(new_n463), .A3(new_n411), .ZN(new_n814));
  NOR2_X1   g628(.A1(new_n628), .A2(new_n814), .ZN(new_n815));
  AND2_X1   g629(.A1(new_n296), .A2(new_n636), .ZN(new_n816));
  NAND3_X1  g630(.A1(new_n644), .A2(new_n815), .A3(new_n816), .ZN(new_n817));
  INV_X1    g631(.A(new_n817), .ZN(new_n818));
  OAI21_X1  g632(.A(KEYINPUT52), .B1(new_n813), .B2(new_n818), .ZN(new_n819));
  AND2_X1   g633(.A1(new_n700), .A2(new_n639), .ZN(new_n820));
  INV_X1    g634(.A(KEYINPUT52), .ZN(new_n821));
  NAND4_X1  g635(.A1(new_n820), .A2(new_n665), .A3(new_n821), .A4(new_n817), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n819), .A2(new_n822), .ZN(new_n823));
  OAI21_X1  g637(.A(new_n789), .B1(new_n811), .B2(new_n823), .ZN(new_n824));
  AOI21_X1  g638(.A(new_n673), .B1(new_n677), .B2(new_n686), .ZN(new_n825));
  INV_X1    g639(.A(new_n360), .ZN(new_n826));
  OR2_X1    g640(.A1(new_n410), .A2(new_n403), .ZN(new_n827));
  AOI21_X1  g641(.A(new_n793), .B1(new_n827), .B2(new_n407), .ZN(new_n828));
  INV_X1    g642(.A(new_n794), .ZN(new_n829));
  OAI21_X1  g643(.A(new_n591), .B1(new_n828), .B2(new_n829), .ZN(new_n830));
  AOI21_X1  g644(.A(new_n717), .B1(new_n830), .B2(KEYINPUT115), .ZN(new_n831));
  AOI21_X1  g645(.A(new_n826), .B1(new_n831), .B2(new_n805), .ZN(new_n832));
  AOI21_X1  g646(.A(new_n579), .B1(new_n832), .B2(new_n590), .ZN(new_n833));
  NAND4_X1  g647(.A1(new_n825), .A2(new_n833), .A3(new_n629), .A4(new_n800), .ZN(new_n834));
  NAND2_X1  g648(.A1(new_n791), .A2(new_n796), .ZN(new_n835));
  NAND2_X1  g649(.A1(new_n835), .A2(new_n628), .ZN(new_n836));
  NAND4_X1  g650(.A1(new_n836), .A2(new_n712), .A3(new_n720), .A4(new_n724), .ZN(new_n837));
  NOR2_X1   g651(.A1(new_n834), .A2(new_n837), .ZN(new_n838));
  AND2_X1   g652(.A1(new_n819), .A2(new_n822), .ZN(new_n839));
  NAND3_X1  g653(.A1(new_n838), .A2(KEYINPUT53), .A3(new_n839), .ZN(new_n840));
  AND3_X1   g654(.A1(new_n824), .A2(KEYINPUT54), .A3(new_n840), .ZN(new_n841));
  AOI21_X1  g655(.A(KEYINPUT54), .B1(new_n824), .B2(new_n840), .ZN(new_n842));
  OAI21_X1  g656(.A(new_n788), .B1(new_n841), .B2(new_n842), .ZN(new_n843));
  INV_X1    g657(.A(KEYINPUT54), .ZN(new_n844));
  AOI21_X1  g658(.A(KEYINPUT53), .B1(new_n838), .B2(new_n839), .ZN(new_n845));
  NOR4_X1   g659(.A1(new_n823), .A2(new_n834), .A3(new_n789), .A4(new_n837), .ZN(new_n846));
  OAI21_X1  g660(.A(new_n844), .B1(new_n845), .B2(new_n846), .ZN(new_n847));
  NAND3_X1  g661(.A1(new_n824), .A2(new_n840), .A3(KEYINPUT54), .ZN(new_n848));
  NAND3_X1  g662(.A1(new_n847), .A2(KEYINPUT116), .A3(new_n848), .ZN(new_n849));
  NAND2_X1  g663(.A1(new_n843), .A2(new_n849), .ZN(new_n850));
  OAI22_X1  g664(.A1(new_n787), .A2(new_n850), .B1(G952), .B2(G953), .ZN(new_n851));
  INV_X1    g665(.A(new_n584), .ZN(new_n852));
  NOR4_X1   g666(.A1(new_n852), .A2(new_n730), .A3(new_n649), .A4(new_n298), .ZN(new_n853));
  XNOR2_X1  g667(.A(new_n772), .B(KEYINPUT49), .ZN(new_n854));
  NAND3_X1  g668(.A1(new_n853), .A2(new_n645), .A3(new_n854), .ZN(new_n855));
  NAND2_X1  g669(.A1(new_n851), .A2(new_n855), .ZN(G75));
  AOI21_X1  g670(.A(new_n289), .B1(new_n824), .B2(new_n840), .ZN(new_n857));
  NAND2_X1  g671(.A1(new_n857), .A2(new_n356), .ZN(new_n858));
  INV_X1    g672(.A(KEYINPUT56), .ZN(new_n859));
  NAND3_X1  g673(.A1(new_n858), .A2(KEYINPUT120), .A3(new_n859), .ZN(new_n860));
  NAND2_X1  g674(.A1(new_n334), .A2(new_n336), .ZN(new_n861));
  XOR2_X1   g675(.A(new_n861), .B(new_n342), .Z(new_n862));
  XNOR2_X1  g676(.A(KEYINPUT119), .B(KEYINPUT55), .ZN(new_n863));
  XNOR2_X1  g677(.A(new_n862), .B(new_n863), .ZN(new_n864));
  AND2_X1   g678(.A1(new_n860), .A2(new_n864), .ZN(new_n865));
  NOR2_X1   g679(.A1(new_n860), .A2(new_n864), .ZN(new_n866));
  NOR2_X1   g680(.A1(new_n192), .A2(G952), .ZN(new_n867));
  NOR3_X1   g681(.A1(new_n865), .A2(new_n866), .A3(new_n867), .ZN(G51));
  XOR2_X1   g682(.A(new_n738), .B(KEYINPUT57), .Z(new_n869));
  NAND3_X1  g683(.A1(new_n847), .A2(new_n848), .A3(new_n869), .ZN(new_n870));
  NAND2_X1  g684(.A1(new_n870), .A2(new_n287), .ZN(new_n871));
  NAND4_X1  g685(.A1(new_n857), .A2(G469), .A3(new_n735), .A4(new_n736), .ZN(new_n872));
  AOI21_X1  g686(.A(new_n867), .B1(new_n871), .B2(new_n872), .ZN(G54));
  INV_X1    g687(.A(new_n867), .ZN(new_n874));
  NAND3_X1  g688(.A1(new_n857), .A2(KEYINPUT58), .A3(G475), .ZN(new_n875));
  NAND2_X1  g689(.A1(new_n450), .A2(new_n455), .ZN(new_n876));
  INV_X1    g690(.A(new_n876), .ZN(new_n877));
  OAI21_X1  g691(.A(new_n874), .B1(new_n875), .B2(new_n877), .ZN(new_n878));
  NAND2_X1  g692(.A1(new_n875), .A2(new_n877), .ZN(new_n879));
  OR2_X1    g693(.A1(new_n879), .A2(KEYINPUT121), .ZN(new_n880));
  NAND2_X1  g694(.A1(new_n879), .A2(KEYINPUT121), .ZN(new_n881));
  AOI21_X1  g695(.A(new_n878), .B1(new_n880), .B2(new_n881), .ZN(G60));
  NAND2_X1  g696(.A1(new_n601), .A2(new_n603), .ZN(new_n883));
  XNOR2_X1  g697(.A(new_n606), .B(KEYINPUT59), .ZN(new_n884));
  AND2_X1   g698(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  NAND3_X1  g699(.A1(new_n847), .A2(new_n848), .A3(new_n885), .ZN(new_n886));
  NAND2_X1  g700(.A1(new_n886), .A2(KEYINPUT122), .ZN(new_n887));
  INV_X1    g701(.A(KEYINPUT122), .ZN(new_n888));
  NAND4_X1  g702(.A1(new_n847), .A2(new_n888), .A3(new_n848), .A4(new_n885), .ZN(new_n889));
  NAND2_X1  g703(.A1(new_n887), .A2(new_n889), .ZN(new_n890));
  NAND2_X1  g704(.A1(new_n890), .A2(new_n874), .ZN(new_n891));
  AOI21_X1  g705(.A(new_n883), .B1(new_n850), .B2(new_n884), .ZN(new_n892));
  NOR2_X1   g706(.A1(new_n891), .A2(new_n892), .ZN(G63));
  XNOR2_X1  g707(.A(KEYINPUT123), .B(KEYINPUT60), .ZN(new_n894));
  NOR2_X1   g708(.A1(new_n569), .A2(new_n289), .ZN(new_n895));
  XNOR2_X1  g709(.A(new_n894), .B(new_n895), .ZN(new_n896));
  OAI21_X1  g710(.A(new_n896), .B1(new_n845), .B2(new_n846), .ZN(new_n897));
  OR2_X1    g711(.A1(new_n897), .A2(new_n625), .ZN(new_n898));
  NAND2_X1  g712(.A1(new_n563), .A2(new_n564), .ZN(new_n899));
  NAND2_X1  g713(.A1(new_n897), .A2(new_n899), .ZN(new_n900));
  NAND3_X1  g714(.A1(new_n898), .A2(new_n874), .A3(new_n900), .ZN(new_n901));
  INV_X1    g715(.A(KEYINPUT61), .ZN(new_n902));
  NAND2_X1  g716(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  NAND4_X1  g717(.A1(new_n898), .A2(KEYINPUT61), .A3(new_n874), .A4(new_n900), .ZN(new_n904));
  NAND2_X1  g718(.A1(new_n903), .A2(new_n904), .ZN(G66));
  NAND2_X1  g719(.A1(new_n834), .A2(new_n192), .ZN(new_n906));
  OAI21_X1  g720(.A(G953), .B1(new_n307), .B2(new_n340), .ZN(new_n907));
  NAND2_X1  g721(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  OAI21_X1  g722(.A(new_n861), .B1(G898), .B2(new_n192), .ZN(new_n909));
  XNOR2_X1  g723(.A(new_n908), .B(new_n909), .ZN(G69));
  AOI21_X1  g724(.A(new_n192), .B1(G227), .B2(G900), .ZN(new_n911));
  XNOR2_X1  g725(.A(new_n513), .B(new_n451), .ZN(new_n912));
  XNOR2_X1  g726(.A(new_n912), .B(KEYINPUT124), .ZN(new_n913));
  INV_X1    g727(.A(new_n913), .ZN(new_n914));
  AND2_X1   g728(.A1(new_n750), .A2(new_n757), .ZN(new_n915));
  INV_X1    g729(.A(KEYINPUT126), .ZN(new_n916));
  INV_X1    g730(.A(KEYINPUT62), .ZN(new_n917));
  NOR2_X1   g731(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  INV_X1    g732(.A(KEYINPUT125), .ZN(new_n919));
  XNOR2_X1  g733(.A(new_n813), .B(new_n919), .ZN(new_n920));
  NAND2_X1  g734(.A1(new_n920), .A2(new_n656), .ZN(new_n921));
  NAND2_X1  g735(.A1(new_n916), .A2(new_n917), .ZN(new_n922));
  AOI21_X1  g736(.A(new_n918), .B1(new_n921), .B2(new_n922), .ZN(new_n923));
  INV_X1    g737(.A(new_n923), .ZN(new_n924));
  NAND2_X1  g738(.A1(new_n921), .A2(new_n918), .ZN(new_n925));
  NAND2_X1  g739(.A1(new_n831), .A2(new_n805), .ZN(new_n926));
  INV_X1    g740(.A(new_n707), .ZN(new_n927));
  NAND4_X1  g741(.A1(new_n926), .A2(new_n713), .A3(new_n651), .A4(new_n927), .ZN(new_n928));
  NAND4_X1  g742(.A1(new_n915), .A2(new_n924), .A3(new_n925), .A4(new_n928), .ZN(new_n929));
  AOI21_X1  g743(.A(new_n914), .B1(new_n929), .B2(new_n192), .ZN(new_n930));
  NAND2_X1  g744(.A1(G900), .A2(G953), .ZN(new_n931));
  INV_X1    g745(.A(new_n814), .ZN(new_n932));
  NAND4_X1  g746(.A1(new_n745), .A2(new_n780), .A3(new_n747), .A4(new_n932), .ZN(new_n933));
  AND4_X1   g747(.A1(new_n712), .A2(new_n933), .A3(new_n720), .A4(new_n724), .ZN(new_n934));
  NAND4_X1  g748(.A1(new_n934), .A2(new_n750), .A3(new_n757), .A4(new_n920), .ZN(new_n935));
  OAI211_X1 g749(.A(new_n912), .B(new_n931), .C1(new_n935), .C2(G953), .ZN(new_n936));
  INV_X1    g750(.A(new_n936), .ZN(new_n937));
  OAI21_X1  g751(.A(new_n911), .B1(new_n930), .B2(new_n937), .ZN(new_n938));
  NAND3_X1  g752(.A1(new_n750), .A2(new_n925), .A3(new_n757), .ZN(new_n939));
  INV_X1    g753(.A(new_n928), .ZN(new_n940));
  NOR3_X1   g754(.A1(new_n939), .A2(new_n923), .A3(new_n940), .ZN(new_n941));
  OAI21_X1  g755(.A(new_n913), .B1(new_n941), .B2(G953), .ZN(new_n942));
  INV_X1    g756(.A(new_n911), .ZN(new_n943));
  NAND3_X1  g757(.A1(new_n942), .A2(new_n943), .A3(new_n936), .ZN(new_n944));
  NAND2_X1  g758(.A1(new_n938), .A2(new_n944), .ZN(G72));
  XNOR2_X1  g759(.A(new_n524), .B(KEYINPUT127), .ZN(new_n946));
  INV_X1    g760(.A(new_n946), .ZN(new_n947));
  NOR4_X1   g761(.A1(new_n939), .A2(new_n834), .A3(new_n923), .A4(new_n940), .ZN(new_n948));
  NAND2_X1  g762(.A1(G472), .A2(G902), .ZN(new_n949));
  XOR2_X1   g763(.A(new_n949), .B(KEYINPUT63), .Z(new_n950));
  INV_X1    g764(.A(new_n950), .ZN(new_n951));
  OAI211_X1 g765(.A(new_n470), .B(new_n947), .C1(new_n948), .C2(new_n951), .ZN(new_n952));
  NOR2_X1   g766(.A1(new_n531), .A2(new_n504), .ZN(new_n953));
  AOI21_X1  g767(.A(new_n953), .B1(new_n824), .B2(new_n840), .ZN(new_n954));
  AOI21_X1  g768(.A(new_n867), .B1(new_n954), .B2(new_n950), .ZN(new_n955));
  OAI21_X1  g769(.A(new_n950), .B1(new_n935), .B2(new_n834), .ZN(new_n956));
  NAND3_X1  g770(.A1(new_n956), .A2(new_n499), .A3(new_n946), .ZN(new_n957));
  AND3_X1   g771(.A1(new_n952), .A2(new_n955), .A3(new_n957), .ZN(G57));
endmodule


