//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 1 1 1 0 0 1 1 0 1 0 1 1 1 1 0 1 1 0 1 1 0 0 0 0 0 1 1 1 1 0 0 1 1 0 1 1 0 0 1 0 0 1 1 0 0 0 0 1 0 1 0 0 1 0 1 0 0 0 0 1 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:24:38 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n703,
    new_n704, new_n705, new_n706, new_n707, new_n708, new_n709, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n737, new_n738, new_n739, new_n740, new_n741, new_n742,
    new_n743, new_n744, new_n745, new_n746, new_n747, new_n749, new_n750,
    new_n751, new_n752, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n769, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n801, new_n802, new_n803,
    new_n804, new_n805, new_n806, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n917, new_n918, new_n919,
    new_n921, new_n922, new_n923, new_n924, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n952, new_n953, new_n954, new_n955, new_n956, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n980,
    new_n981, new_n982, new_n983, new_n984, new_n985, new_n986, new_n987,
    new_n988, new_n989, new_n990, new_n991, new_n992, new_n993, new_n994,
    new_n995, new_n996, new_n997;
  INV_X1    g000(.A(G902), .ZN(new_n187));
  XNOR2_X1  g001(.A(G110), .B(G140), .ZN(new_n188));
  INV_X1    g002(.A(G227), .ZN(new_n189));
  NOR2_X1   g003(.A1(new_n189), .A2(G953), .ZN(new_n190));
  XNOR2_X1  g004(.A(new_n188), .B(new_n190), .ZN(new_n191));
  INV_X1    g005(.A(new_n191), .ZN(new_n192));
  NAND2_X1  g006(.A1(KEYINPUT76), .A2(KEYINPUT3), .ZN(new_n193));
  INV_X1    g007(.A(G104), .ZN(new_n194));
  NOR2_X1   g008(.A1(new_n194), .A2(G107), .ZN(new_n195));
  NOR2_X1   g009(.A1(KEYINPUT76), .A2(KEYINPUT3), .ZN(new_n196));
  OAI21_X1  g010(.A(new_n193), .B1(new_n195), .B2(new_n196), .ZN(new_n197));
  INV_X1    g011(.A(G107), .ZN(new_n198));
  OAI21_X1  g012(.A(KEYINPUT77), .B1(new_n198), .B2(G104), .ZN(new_n199));
  INV_X1    g013(.A(KEYINPUT77), .ZN(new_n200));
  NAND3_X1  g014(.A1(new_n200), .A2(new_n194), .A3(G107), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n199), .A2(new_n201), .ZN(new_n202));
  INV_X1    g016(.A(G101), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n198), .A2(G104), .ZN(new_n204));
  NAND3_X1  g018(.A1(new_n204), .A2(KEYINPUT76), .A3(KEYINPUT3), .ZN(new_n205));
  NAND4_X1  g019(.A1(new_n197), .A2(new_n202), .A3(new_n203), .A4(new_n205), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n194), .A2(G107), .ZN(new_n207));
  NAND3_X1  g021(.A1(new_n204), .A2(new_n207), .A3(KEYINPUT78), .ZN(new_n208));
  OAI211_X1 g022(.A(new_n208), .B(G101), .C1(KEYINPUT78), .C2(new_n207), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n206), .A2(new_n209), .ZN(new_n210));
  INV_X1    g024(.A(G143), .ZN(new_n211));
  AND3_X1   g025(.A1(new_n211), .A2(KEYINPUT1), .A3(G146), .ZN(new_n212));
  INV_X1    g026(.A(G146), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n213), .A2(G143), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n211), .A2(G146), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n214), .A2(new_n215), .ZN(new_n216));
  INV_X1    g030(.A(G128), .ZN(new_n217));
  AOI21_X1  g031(.A(new_n212), .B1(new_n216), .B2(new_n217), .ZN(new_n218));
  NOR2_X1   g032(.A1(new_n217), .A2(KEYINPUT1), .ZN(new_n219));
  NAND3_X1  g033(.A1(new_n219), .A2(new_n214), .A3(new_n215), .ZN(new_n220));
  AND2_X1   g034(.A1(new_n218), .A2(new_n220), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n210), .A2(new_n221), .ZN(new_n222));
  INV_X1    g036(.A(KEYINPUT79), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n220), .A2(new_n223), .ZN(new_n224));
  NAND4_X1  g038(.A1(new_n219), .A2(new_n214), .A3(new_n215), .A4(KEYINPUT79), .ZN(new_n225));
  NAND3_X1  g039(.A1(new_n218), .A2(new_n224), .A3(new_n225), .ZN(new_n226));
  NAND3_X1  g040(.A1(new_n226), .A2(new_n206), .A3(new_n209), .ZN(new_n227));
  NAND3_X1  g041(.A1(new_n222), .A2(new_n227), .A3(KEYINPUT81), .ZN(new_n228));
  INV_X1    g042(.A(KEYINPUT81), .ZN(new_n229));
  NAND3_X1  g043(.A1(new_n210), .A2(new_n221), .A3(new_n229), .ZN(new_n230));
  INV_X1    g044(.A(G134), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n231), .A2(G137), .ZN(new_n232));
  INV_X1    g046(.A(G137), .ZN(new_n233));
  AOI21_X1  g047(.A(KEYINPUT65), .B1(new_n233), .B2(G134), .ZN(new_n234));
  INV_X1    g048(.A(KEYINPUT11), .ZN(new_n235));
  OAI21_X1  g049(.A(new_n232), .B1(new_n234), .B2(new_n235), .ZN(new_n236));
  INV_X1    g050(.A(KEYINPUT65), .ZN(new_n237));
  OAI211_X1 g051(.A(new_n237), .B(new_n235), .C1(new_n231), .C2(G137), .ZN(new_n238));
  INV_X1    g052(.A(new_n238), .ZN(new_n239));
  NOR3_X1   g053(.A1(new_n236), .A2(new_n239), .A3(G131), .ZN(new_n240));
  INV_X1    g054(.A(G131), .ZN(new_n241));
  NOR2_X1   g055(.A1(new_n233), .A2(G134), .ZN(new_n242));
  OAI21_X1  g056(.A(new_n237), .B1(new_n231), .B2(G137), .ZN(new_n243));
  AOI21_X1  g057(.A(new_n242), .B1(new_n243), .B2(KEYINPUT11), .ZN(new_n244));
  AOI21_X1  g058(.A(new_n241), .B1(new_n244), .B2(new_n238), .ZN(new_n245));
  NOR2_X1   g059(.A1(new_n240), .A2(new_n245), .ZN(new_n246));
  XNOR2_X1  g060(.A(KEYINPUT80), .B(KEYINPUT12), .ZN(new_n247));
  NOR2_X1   g061(.A1(new_n246), .A2(new_n247), .ZN(new_n248));
  NAND3_X1  g062(.A1(new_n228), .A2(new_n230), .A3(new_n248), .ZN(new_n249));
  INV_X1    g063(.A(KEYINPUT69), .ZN(new_n250));
  OAI21_X1  g064(.A(new_n250), .B1(new_n240), .B2(new_n245), .ZN(new_n251));
  OAI21_X1  g065(.A(G131), .B1(new_n236), .B2(new_n239), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n243), .A2(KEYINPUT11), .ZN(new_n253));
  NAND4_X1  g067(.A1(new_n253), .A2(new_n241), .A3(new_n238), .A4(new_n232), .ZN(new_n254));
  NAND3_X1  g068(.A1(new_n252), .A2(KEYINPUT69), .A3(new_n254), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n251), .A2(new_n255), .ZN(new_n256));
  NAND3_X1  g070(.A1(new_n228), .A2(new_n256), .A3(new_n230), .ZN(new_n257));
  INV_X1    g071(.A(KEYINPUT82), .ZN(new_n258));
  INV_X1    g072(.A(KEYINPUT12), .ZN(new_n259));
  AND3_X1   g073(.A1(new_n257), .A2(new_n258), .A3(new_n259), .ZN(new_n260));
  AOI21_X1  g074(.A(new_n258), .B1(new_n257), .B2(new_n259), .ZN(new_n261));
  OAI21_X1  g075(.A(new_n249), .B1(new_n260), .B2(new_n261), .ZN(new_n262));
  INV_X1    g076(.A(KEYINPUT10), .ZN(new_n263));
  INV_X1    g077(.A(new_n210), .ZN(new_n264));
  AOI21_X1  g078(.A(new_n263), .B1(new_n218), .B2(new_n220), .ZN(new_n265));
  AOI22_X1  g079(.A1(new_n227), .A2(new_n263), .B1(new_n264), .B2(new_n265), .ZN(new_n266));
  AND3_X1   g080(.A1(new_n252), .A2(KEYINPUT69), .A3(new_n254), .ZN(new_n267));
  AOI21_X1  g081(.A(KEYINPUT69), .B1(new_n252), .B2(new_n254), .ZN(new_n268));
  NOR2_X1   g082(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  NAND3_X1  g083(.A1(new_n197), .A2(new_n202), .A3(new_n205), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n270), .A2(G101), .ZN(new_n271));
  NAND3_X1  g085(.A1(new_n271), .A2(KEYINPUT4), .A3(new_n206), .ZN(new_n272));
  AND2_X1   g086(.A1(KEYINPUT0), .A2(G128), .ZN(new_n273));
  NOR2_X1   g087(.A1(KEYINPUT0), .A2(G128), .ZN(new_n274));
  NOR2_X1   g088(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  AOI21_X1  g089(.A(new_n275), .B1(new_n214), .B2(new_n215), .ZN(new_n276));
  NOR2_X1   g090(.A1(new_n216), .A2(new_n273), .ZN(new_n277));
  NOR2_X1   g091(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  INV_X1    g092(.A(new_n278), .ZN(new_n279));
  INV_X1    g093(.A(KEYINPUT4), .ZN(new_n280));
  NAND3_X1  g094(.A1(new_n270), .A2(new_n280), .A3(G101), .ZN(new_n281));
  NAND3_X1  g095(.A1(new_n272), .A2(new_n279), .A3(new_n281), .ZN(new_n282));
  NAND3_X1  g096(.A1(new_n266), .A2(new_n269), .A3(new_n282), .ZN(new_n283));
  AOI21_X1  g097(.A(new_n192), .B1(new_n262), .B2(new_n283), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n266), .A2(new_n282), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n285), .A2(new_n256), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n283), .A2(new_n192), .ZN(new_n287));
  INV_X1    g101(.A(KEYINPUT83), .ZN(new_n288));
  OAI21_X1  g102(.A(new_n286), .B1(new_n287), .B2(new_n288), .ZN(new_n289));
  AOI21_X1  g103(.A(new_n289), .B1(new_n288), .B2(new_n287), .ZN(new_n290));
  OAI21_X1  g104(.A(new_n187), .B1(new_n284), .B2(new_n290), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n291), .A2(G469), .ZN(new_n292));
  INV_X1    g106(.A(KEYINPUT84), .ZN(new_n293));
  INV_X1    g107(.A(new_n287), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n262), .A2(new_n294), .ZN(new_n295));
  AOI21_X1  g109(.A(new_n192), .B1(new_n286), .B2(new_n283), .ZN(new_n296));
  INV_X1    g110(.A(new_n296), .ZN(new_n297));
  AOI21_X1  g111(.A(G902), .B1(new_n295), .B2(new_n297), .ZN(new_n298));
  INV_X1    g112(.A(G469), .ZN(new_n299));
  AOI21_X1  g113(.A(new_n293), .B1(new_n298), .B2(new_n299), .ZN(new_n300));
  AOI21_X1  g114(.A(new_n296), .B1(new_n262), .B2(new_n294), .ZN(new_n301));
  NOR4_X1   g115(.A1(new_n301), .A2(KEYINPUT84), .A3(G469), .A4(G902), .ZN(new_n302));
  OAI21_X1  g116(.A(new_n292), .B1(new_n300), .B2(new_n302), .ZN(new_n303));
  INV_X1    g117(.A(G478), .ZN(new_n304));
  NOR2_X1   g118(.A1(new_n304), .A2(KEYINPUT15), .ZN(new_n305));
  OR2_X1    g119(.A1(KEYINPUT67), .A2(G116), .ZN(new_n306));
  NAND2_X1  g120(.A1(KEYINPUT67), .A2(G116), .ZN(new_n307));
  NAND3_X1  g121(.A1(new_n306), .A2(G122), .A3(new_n307), .ZN(new_n308));
  INV_X1    g122(.A(G116), .ZN(new_n309));
  OR2_X1    g123(.A1(new_n309), .A2(G122), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n308), .A2(new_n310), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n311), .A2(G107), .ZN(new_n312));
  NAND3_X1  g126(.A1(new_n308), .A2(new_n198), .A3(new_n310), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  INV_X1    g128(.A(KEYINPUT92), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  NAND3_X1  g130(.A1(new_n312), .A2(KEYINPUT92), .A3(new_n313), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n211), .A2(G128), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n217), .A2(G143), .ZN(new_n319));
  AND3_X1   g133(.A1(new_n318), .A2(new_n319), .A3(new_n231), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n319), .A2(KEYINPUT13), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n321), .A2(new_n318), .ZN(new_n322));
  INV_X1    g136(.A(KEYINPUT93), .ZN(new_n323));
  NOR2_X1   g137(.A1(new_n217), .A2(G143), .ZN(new_n324));
  AOI21_X1  g138(.A(new_n323), .B1(new_n324), .B2(KEYINPUT13), .ZN(new_n325));
  AOI21_X1  g139(.A(new_n231), .B1(new_n322), .B2(new_n325), .ZN(new_n326));
  NAND3_X1  g140(.A1(new_n321), .A2(new_n323), .A3(new_n318), .ZN(new_n327));
  AOI21_X1  g141(.A(new_n320), .B1(new_n326), .B2(new_n327), .ZN(new_n328));
  NAND3_X1  g142(.A1(new_n316), .A2(new_n317), .A3(new_n328), .ZN(new_n329));
  AOI21_X1  g143(.A(new_n231), .B1(new_n318), .B2(new_n319), .ZN(new_n330));
  INV_X1    g144(.A(KEYINPUT94), .ZN(new_n331));
  OR3_X1    g145(.A1(new_n320), .A2(new_n330), .A3(new_n331), .ZN(new_n332));
  NAND4_X1  g146(.A1(new_n306), .A2(KEYINPUT14), .A3(G122), .A4(new_n307), .ZN(new_n333));
  OAI211_X1 g147(.A(G107), .B(new_n333), .C1(new_n311), .C2(KEYINPUT14), .ZN(new_n334));
  OAI21_X1  g148(.A(new_n331), .B1(new_n320), .B2(new_n330), .ZN(new_n335));
  NAND4_X1  g149(.A1(new_n332), .A2(new_n334), .A3(new_n313), .A4(new_n335), .ZN(new_n336));
  XNOR2_X1  g150(.A(KEYINPUT9), .B(G234), .ZN(new_n337));
  INV_X1    g151(.A(new_n337), .ZN(new_n338));
  INV_X1    g152(.A(G953), .ZN(new_n339));
  NAND3_X1  g153(.A1(new_n338), .A2(G217), .A3(new_n339), .ZN(new_n340));
  INV_X1    g154(.A(new_n340), .ZN(new_n341));
  AND3_X1   g155(.A1(new_n329), .A2(new_n336), .A3(new_n341), .ZN(new_n342));
  AOI21_X1  g156(.A(new_n341), .B1(new_n329), .B2(new_n336), .ZN(new_n343));
  OAI21_X1  g157(.A(new_n187), .B1(new_n342), .B2(new_n343), .ZN(new_n344));
  INV_X1    g158(.A(KEYINPUT95), .ZN(new_n345));
  AOI21_X1  g159(.A(new_n305), .B1(new_n344), .B2(new_n345), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n329), .A2(new_n336), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n347), .A2(new_n340), .ZN(new_n348));
  NAND3_X1  g162(.A1(new_n329), .A2(new_n336), .A3(new_n341), .ZN(new_n349));
  AOI21_X1  g163(.A(G902), .B1(new_n348), .B2(new_n349), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n350), .A2(KEYINPUT95), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n344), .A2(new_n345), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n351), .A2(new_n352), .ZN(new_n353));
  AOI21_X1  g167(.A(new_n346), .B1(new_n353), .B2(new_n305), .ZN(new_n354));
  INV_X1    g168(.A(KEYINPUT89), .ZN(new_n355));
  INV_X1    g169(.A(G237), .ZN(new_n356));
  NAND3_X1  g170(.A1(new_n356), .A2(new_n339), .A3(G214), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n357), .A2(new_n211), .ZN(new_n358));
  NOR2_X1   g172(.A1(G237), .A2(G953), .ZN(new_n359));
  NAND3_X1  g173(.A1(new_n359), .A2(G143), .A3(G214), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n358), .A2(new_n360), .ZN(new_n361));
  AND2_X1   g175(.A1(KEYINPUT18), .A2(G131), .ZN(new_n362));
  OR2_X1    g176(.A1(new_n361), .A2(new_n362), .ZN(new_n363));
  INV_X1    g177(.A(G140), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n364), .A2(G125), .ZN(new_n365));
  INV_X1    g179(.A(G125), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n366), .A2(G140), .ZN(new_n367));
  AND2_X1   g181(.A1(new_n365), .A2(new_n367), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n368), .A2(new_n213), .ZN(new_n369));
  INV_X1    g183(.A(KEYINPUT75), .ZN(new_n370));
  NAND3_X1  g184(.A1(new_n365), .A2(new_n367), .A3(new_n370), .ZN(new_n371));
  NAND3_X1  g185(.A1(new_n366), .A2(KEYINPUT75), .A3(G140), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  OAI21_X1  g187(.A(new_n369), .B1(new_n373), .B2(new_n213), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n361), .A2(new_n362), .ZN(new_n375));
  AND3_X1   g189(.A1(new_n363), .A2(new_n374), .A3(new_n375), .ZN(new_n376));
  NAND3_X1  g190(.A1(new_n371), .A2(KEYINPUT16), .A3(new_n372), .ZN(new_n377));
  INV_X1    g191(.A(KEYINPUT16), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n365), .A2(new_n378), .ZN(new_n379));
  AOI21_X1  g193(.A(new_n213), .B1(new_n377), .B2(new_n379), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n373), .A2(KEYINPUT19), .ZN(new_n381));
  OAI21_X1  g195(.A(new_n381), .B1(KEYINPUT19), .B2(new_n368), .ZN(new_n382));
  AOI21_X1  g196(.A(new_n380), .B1(new_n382), .B2(new_n213), .ZN(new_n383));
  OAI21_X1  g197(.A(KEYINPUT88), .B1(new_n361), .B2(G131), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n361), .A2(G131), .ZN(new_n385));
  INV_X1    g199(.A(KEYINPUT88), .ZN(new_n386));
  NAND4_X1  g200(.A1(new_n358), .A2(new_n386), .A3(new_n241), .A4(new_n360), .ZN(new_n387));
  NAND3_X1  g201(.A1(new_n384), .A2(new_n385), .A3(new_n387), .ZN(new_n388));
  AOI21_X1  g202(.A(new_n376), .B1(new_n383), .B2(new_n388), .ZN(new_n389));
  XNOR2_X1  g203(.A(G113), .B(G122), .ZN(new_n390));
  XNOR2_X1  g204(.A(new_n390), .B(new_n194), .ZN(new_n391));
  OAI21_X1  g205(.A(new_n355), .B1(new_n389), .B2(new_n391), .ZN(new_n392));
  INV_X1    g206(.A(new_n380), .ZN(new_n393));
  NOR2_X1   g207(.A1(new_n368), .A2(KEYINPUT19), .ZN(new_n394));
  AOI21_X1  g208(.A(new_n394), .B1(new_n373), .B2(KEYINPUT19), .ZN(new_n395));
  OAI211_X1 g209(.A(new_n388), .B(new_n393), .C1(G146), .C2(new_n395), .ZN(new_n396));
  INV_X1    g210(.A(new_n376), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n396), .A2(new_n397), .ZN(new_n398));
  INV_X1    g212(.A(new_n391), .ZN(new_n399));
  NAND3_X1  g213(.A1(new_n398), .A2(KEYINPUT89), .A3(new_n399), .ZN(new_n400));
  NAND3_X1  g214(.A1(new_n377), .A2(new_n213), .A3(new_n379), .ZN(new_n401));
  NAND3_X1  g215(.A1(new_n361), .A2(KEYINPUT17), .A3(G131), .ZN(new_n402));
  AND3_X1   g216(.A1(new_n393), .A2(new_n401), .A3(new_n402), .ZN(new_n403));
  INV_X1    g217(.A(KEYINPUT17), .ZN(new_n404));
  NAND4_X1  g218(.A1(new_n384), .A2(new_n404), .A3(new_n385), .A4(new_n387), .ZN(new_n405));
  AOI21_X1  g219(.A(new_n376), .B1(new_n403), .B2(new_n405), .ZN(new_n406));
  XOR2_X1   g220(.A(new_n391), .B(KEYINPUT90), .Z(new_n407));
  AOI22_X1  g221(.A1(new_n392), .A2(new_n400), .B1(new_n406), .B2(new_n407), .ZN(new_n408));
  NOR2_X1   g222(.A1(G475), .A2(G902), .ZN(new_n409));
  INV_X1    g223(.A(new_n409), .ZN(new_n410));
  OAI21_X1  g224(.A(KEYINPUT20), .B1(new_n408), .B2(new_n410), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n406), .A2(new_n407), .ZN(new_n412));
  AOI21_X1  g226(.A(KEYINPUT89), .B1(new_n398), .B2(new_n399), .ZN(new_n413));
  AOI211_X1 g227(.A(new_n355), .B(new_n391), .C1(new_n396), .C2(new_n397), .ZN(new_n414));
  OAI21_X1  g228(.A(new_n412), .B1(new_n413), .B2(new_n414), .ZN(new_n415));
  INV_X1    g229(.A(KEYINPUT20), .ZN(new_n416));
  NAND3_X1  g230(.A1(new_n415), .A2(new_n416), .A3(new_n409), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n411), .A2(new_n417), .ZN(new_n418));
  OAI21_X1  g232(.A(new_n412), .B1(new_n406), .B2(new_n391), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n419), .A2(new_n187), .ZN(new_n420));
  XOR2_X1   g234(.A(KEYINPUT91), .B(G475), .Z(new_n421));
  INV_X1    g235(.A(new_n421), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n420), .A2(new_n422), .ZN(new_n423));
  NAND2_X1  g237(.A1(G234), .A2(G237), .ZN(new_n424));
  NAND3_X1  g238(.A1(new_n424), .A2(G952), .A3(new_n339), .ZN(new_n425));
  XNOR2_X1  g239(.A(KEYINPUT21), .B(G898), .ZN(new_n426));
  INV_X1    g240(.A(new_n426), .ZN(new_n427));
  NAND3_X1  g241(.A1(new_n424), .A2(G902), .A3(G953), .ZN(new_n428));
  OAI21_X1  g242(.A(new_n425), .B1(new_n427), .B2(new_n428), .ZN(new_n429));
  NAND4_X1  g243(.A1(new_n354), .A2(new_n418), .A3(new_n423), .A4(new_n429), .ZN(new_n430));
  OAI21_X1  g244(.A(G214), .B1(G237), .B2(G902), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n339), .A2(G224), .ZN(new_n432));
  OR2_X1    g246(.A1(new_n432), .A2(KEYINPUT86), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n432), .A2(KEYINPUT86), .ZN(new_n434));
  NAND3_X1  g248(.A1(new_n433), .A2(KEYINPUT7), .A3(new_n434), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n218), .A2(new_n220), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n436), .A2(new_n366), .ZN(new_n437));
  OAI21_X1  g251(.A(G125), .B1(new_n276), .B2(new_n277), .ZN(new_n438));
  AOI21_X1  g252(.A(new_n435), .B1(new_n437), .B2(new_n438), .ZN(new_n439));
  NOR2_X1   g253(.A1(new_n439), .A2(KEYINPUT87), .ZN(new_n440));
  INV_X1    g254(.A(KEYINPUT87), .ZN(new_n441));
  AOI211_X1 g255(.A(new_n441), .B(new_n435), .C1(new_n437), .C2(new_n438), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n437), .A2(new_n438), .ZN(new_n443));
  AND2_X1   g257(.A1(new_n432), .A2(KEYINPUT7), .ZN(new_n444));
  OAI22_X1  g258(.A1(new_n440), .A2(new_n442), .B1(new_n443), .B2(new_n444), .ZN(new_n445));
  XNOR2_X1  g259(.A(G110), .B(G122), .ZN(new_n446));
  XOR2_X1   g260(.A(new_n446), .B(KEYINPUT8), .Z(new_n447));
  INV_X1    g261(.A(KEYINPUT68), .ZN(new_n448));
  NAND4_X1  g262(.A1(new_n306), .A2(new_n448), .A3(G119), .A4(new_n307), .ZN(new_n449));
  AND3_X1   g263(.A1(new_n306), .A2(G119), .A3(new_n307), .ZN(new_n450));
  OAI21_X1  g264(.A(KEYINPUT68), .B1(new_n309), .B2(G119), .ZN(new_n451));
  OAI21_X1  g265(.A(new_n449), .B1(new_n450), .B2(new_n451), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n452), .A2(KEYINPUT5), .ZN(new_n453));
  INV_X1    g267(.A(G113), .ZN(new_n454));
  NOR2_X1   g268(.A1(new_n309), .A2(G119), .ZN(new_n455));
  INV_X1    g269(.A(KEYINPUT5), .ZN(new_n456));
  AOI21_X1  g270(.A(new_n454), .B1(new_n455), .B2(new_n456), .ZN(new_n457));
  XNOR2_X1  g271(.A(new_n457), .B(KEYINPUT85), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n453), .A2(new_n458), .ZN(new_n459));
  XNOR2_X1  g273(.A(KEYINPUT2), .B(G113), .ZN(new_n460));
  INV_X1    g274(.A(new_n460), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n452), .A2(new_n461), .ZN(new_n462));
  NAND3_X1  g276(.A1(new_n459), .A2(new_n264), .A3(new_n462), .ZN(new_n463));
  INV_X1    g277(.A(new_n462), .ZN(new_n464));
  INV_X1    g278(.A(new_n457), .ZN(new_n465));
  AOI21_X1  g279(.A(new_n465), .B1(new_n452), .B2(KEYINPUT5), .ZN(new_n466));
  OAI21_X1  g280(.A(new_n210), .B1(new_n464), .B2(new_n466), .ZN(new_n467));
  AOI21_X1  g281(.A(new_n447), .B1(new_n463), .B2(new_n467), .ZN(new_n468));
  NOR2_X1   g282(.A1(new_n445), .A2(new_n468), .ZN(new_n469));
  OAI211_X1 g283(.A(KEYINPUT66), .B(new_n449), .C1(new_n450), .C2(new_n451), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n470), .A2(new_n461), .ZN(new_n471));
  NAND3_X1  g285(.A1(new_n306), .A2(G119), .A3(new_n307), .ZN(new_n472));
  OAI211_X1 g286(.A(new_n472), .B(KEYINPUT68), .C1(new_n309), .C2(G119), .ZN(new_n473));
  NAND4_X1  g287(.A1(new_n473), .A2(KEYINPUT66), .A3(new_n449), .A4(new_n460), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n471), .A2(new_n474), .ZN(new_n475));
  NAND3_X1  g289(.A1(new_n475), .A2(new_n281), .A3(new_n272), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n453), .A2(new_n457), .ZN(new_n477));
  NAND3_X1  g291(.A1(new_n477), .A2(new_n264), .A3(new_n462), .ZN(new_n478));
  NAND3_X1  g292(.A1(new_n476), .A2(new_n446), .A3(new_n478), .ZN(new_n479));
  AOI21_X1  g293(.A(G902), .B1(new_n469), .B2(new_n479), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n476), .A2(new_n478), .ZN(new_n481));
  INV_X1    g295(.A(new_n446), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  NAND3_X1  g297(.A1(new_n483), .A2(KEYINPUT6), .A3(new_n479), .ZN(new_n484));
  XNOR2_X1  g298(.A(new_n443), .B(new_n432), .ZN(new_n485));
  INV_X1    g299(.A(KEYINPUT6), .ZN(new_n486));
  NAND3_X1  g300(.A1(new_n481), .A2(new_n486), .A3(new_n482), .ZN(new_n487));
  NAND3_X1  g301(.A1(new_n484), .A2(new_n485), .A3(new_n487), .ZN(new_n488));
  OAI21_X1  g302(.A(G210), .B1(G237), .B2(G902), .ZN(new_n489));
  AND3_X1   g303(.A1(new_n480), .A2(new_n488), .A3(new_n489), .ZN(new_n490));
  AOI21_X1  g304(.A(new_n489), .B1(new_n480), .B2(new_n488), .ZN(new_n491));
  OAI21_X1  g305(.A(new_n431), .B1(new_n490), .B2(new_n491), .ZN(new_n492));
  NOR2_X1   g306(.A1(new_n430), .A2(new_n492), .ZN(new_n493));
  INV_X1    g307(.A(G221), .ZN(new_n494));
  AOI21_X1  g308(.A(new_n494), .B1(new_n338), .B2(new_n187), .ZN(new_n495));
  INV_X1    g309(.A(new_n495), .ZN(new_n496));
  NAND3_X1  g310(.A1(new_n303), .A2(new_n493), .A3(new_n496), .ZN(new_n497));
  INV_X1    g311(.A(KEYINPUT96), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  OAI21_X1  g313(.A(new_n279), .B1(new_n267), .B2(new_n268), .ZN(new_n500));
  NOR2_X1   g314(.A1(new_n231), .A2(G137), .ZN(new_n501));
  OAI21_X1  g315(.A(G131), .B1(new_n501), .B2(new_n242), .ZN(new_n502));
  AOI21_X1  g316(.A(KEYINPUT70), .B1(new_n254), .B2(new_n502), .ZN(new_n503));
  INV_X1    g317(.A(new_n503), .ZN(new_n504));
  NAND3_X1  g318(.A1(new_n254), .A2(KEYINPUT70), .A3(new_n502), .ZN(new_n505));
  NAND3_X1  g319(.A1(new_n504), .A2(new_n505), .A3(new_n436), .ZN(new_n506));
  INV_X1    g320(.A(new_n475), .ZN(new_n507));
  NAND3_X1  g321(.A1(new_n500), .A2(new_n506), .A3(new_n507), .ZN(new_n508));
  INV_X1    g322(.A(KEYINPUT28), .ZN(new_n509));
  AOI21_X1  g323(.A(KEYINPUT71), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  AND3_X1   g324(.A1(new_n508), .A2(KEYINPUT71), .A3(new_n509), .ZN(new_n511));
  AOI21_X1  g325(.A(new_n278), .B1(new_n251), .B2(new_n255), .ZN(new_n512));
  AND3_X1   g326(.A1(new_n254), .A2(KEYINPUT70), .A3(new_n502), .ZN(new_n513));
  NOR3_X1   g327(.A1(new_n513), .A2(new_n503), .A3(new_n221), .ZN(new_n514));
  NOR2_X1   g328(.A1(new_n512), .A2(new_n514), .ZN(new_n515));
  XNOR2_X1  g329(.A(new_n515), .B(new_n507), .ZN(new_n516));
  AOI211_X1 g330(.A(new_n510), .B(new_n511), .C1(new_n516), .C2(KEYINPUT28), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n359), .A2(G210), .ZN(new_n518));
  XNOR2_X1  g332(.A(new_n518), .B(KEYINPUT27), .ZN(new_n519));
  XNOR2_X1  g333(.A(KEYINPUT26), .B(G101), .ZN(new_n520));
  XNOR2_X1  g334(.A(new_n519), .B(new_n520), .ZN(new_n521));
  INV_X1    g335(.A(new_n521), .ZN(new_n522));
  INV_X1    g336(.A(KEYINPUT29), .ZN(new_n523));
  NOR2_X1   g337(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n517), .A2(new_n524), .ZN(new_n525));
  NAND3_X1  g339(.A1(new_n500), .A2(KEYINPUT30), .A3(new_n506), .ZN(new_n526));
  NAND3_X1  g340(.A1(new_n436), .A2(new_n254), .A3(new_n502), .ZN(new_n527));
  OAI21_X1  g341(.A(new_n527), .B1(new_n278), .B2(new_n246), .ZN(new_n528));
  XNOR2_X1  g342(.A(KEYINPUT64), .B(KEYINPUT30), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  NAND3_X1  g344(.A1(new_n526), .A2(new_n475), .A3(new_n530), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n531), .A2(new_n508), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n532), .A2(new_n522), .ZN(new_n533));
  INV_X1    g347(.A(KEYINPUT71), .ZN(new_n534));
  NOR3_X1   g348(.A1(new_n512), .A2(new_n514), .A3(new_n475), .ZN(new_n535));
  OAI21_X1  g349(.A(new_n534), .B1(new_n535), .B2(KEYINPUT28), .ZN(new_n536));
  AND2_X1   g350(.A1(new_n528), .A2(new_n475), .ZN(new_n537));
  OAI21_X1  g351(.A(KEYINPUT28), .B1(new_n535), .B2(new_n537), .ZN(new_n538));
  NAND3_X1  g352(.A1(new_n508), .A2(KEYINPUT71), .A3(new_n509), .ZN(new_n539));
  NAND3_X1  g353(.A1(new_n536), .A2(new_n538), .A3(new_n539), .ZN(new_n540));
  OAI211_X1 g354(.A(new_n523), .B(new_n533), .C1(new_n540), .C2(new_n522), .ZN(new_n541));
  NAND3_X1  g355(.A1(new_n525), .A2(new_n187), .A3(new_n541), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n542), .A2(G472), .ZN(new_n543));
  INV_X1    g357(.A(KEYINPUT32), .ZN(new_n544));
  NOR2_X1   g358(.A1(new_n511), .A2(new_n510), .ZN(new_n545));
  AOI21_X1  g359(.A(new_n521), .B1(new_n545), .B2(new_n538), .ZN(new_n546));
  AOI21_X1  g360(.A(new_n522), .B1(new_n515), .B2(new_n507), .ZN(new_n547));
  AND3_X1   g361(.A1(new_n547), .A2(new_n531), .A3(KEYINPUT31), .ZN(new_n548));
  AOI21_X1  g362(.A(KEYINPUT31), .B1(new_n547), .B2(new_n531), .ZN(new_n549));
  NOR2_X1   g363(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  OAI21_X1  g364(.A(KEYINPUT72), .B1(new_n546), .B2(new_n550), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n540), .A2(new_n522), .ZN(new_n552));
  INV_X1    g366(.A(KEYINPUT31), .ZN(new_n553));
  AND3_X1   g367(.A1(new_n526), .A2(new_n475), .A3(new_n530), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n508), .A2(new_n521), .ZN(new_n555));
  OAI21_X1  g369(.A(new_n553), .B1(new_n554), .B2(new_n555), .ZN(new_n556));
  NAND3_X1  g370(.A1(new_n547), .A2(new_n531), .A3(KEYINPUT31), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  INV_X1    g372(.A(KEYINPUT72), .ZN(new_n559));
  NAND3_X1  g373(.A1(new_n552), .A2(new_n558), .A3(new_n559), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n551), .A2(new_n560), .ZN(new_n561));
  NOR2_X1   g375(.A1(G472), .A2(G902), .ZN(new_n562));
  AOI21_X1  g376(.A(new_n544), .B1(new_n561), .B2(new_n562), .ZN(new_n563));
  INV_X1    g377(.A(new_n562), .ZN(new_n564));
  AOI211_X1 g378(.A(KEYINPUT32), .B(new_n564), .C1(new_n551), .C2(new_n560), .ZN(new_n565));
  OAI21_X1  g379(.A(new_n543), .B1(new_n563), .B2(new_n565), .ZN(new_n566));
  INV_X1    g380(.A(G234), .ZN(new_n567));
  OAI21_X1  g381(.A(G217), .B1(new_n567), .B2(G902), .ZN(new_n568));
  XNOR2_X1  g382(.A(new_n568), .B(KEYINPUT73), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n393), .A2(new_n401), .ZN(new_n570));
  XOR2_X1   g384(.A(G119), .B(G128), .Z(new_n571));
  XNOR2_X1  g385(.A(KEYINPUT24), .B(G110), .ZN(new_n572));
  NOR2_X1   g386(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  INV_X1    g387(.A(KEYINPUT74), .ZN(new_n574));
  AOI21_X1  g388(.A(new_n574), .B1(G119), .B2(new_n217), .ZN(new_n575));
  OAI21_X1  g389(.A(KEYINPUT23), .B1(new_n217), .B2(G119), .ZN(new_n576));
  XNOR2_X1  g390(.A(new_n575), .B(new_n576), .ZN(new_n577));
  AOI21_X1  g391(.A(new_n573), .B1(new_n577), .B2(G110), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n570), .A2(new_n578), .ZN(new_n579));
  NOR2_X1   g393(.A1(new_n577), .A2(G110), .ZN(new_n580));
  AND2_X1   g394(.A1(new_n571), .A2(new_n572), .ZN(new_n581));
  OAI211_X1 g395(.A(new_n393), .B(new_n369), .C1(new_n580), .C2(new_n581), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n579), .A2(new_n582), .ZN(new_n583));
  XNOR2_X1  g397(.A(KEYINPUT22), .B(G137), .ZN(new_n584));
  NOR3_X1   g398(.A1(new_n494), .A2(new_n567), .A3(G953), .ZN(new_n585));
  XOR2_X1   g399(.A(new_n584), .B(new_n585), .Z(new_n586));
  INV_X1    g400(.A(new_n586), .ZN(new_n587));
  NOR2_X1   g401(.A1(new_n583), .A2(new_n587), .ZN(new_n588));
  AOI21_X1  g402(.A(new_n586), .B1(new_n579), .B2(new_n582), .ZN(new_n589));
  NOR2_X1   g403(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  AOI21_X1  g404(.A(KEYINPUT25), .B1(new_n590), .B2(new_n187), .ZN(new_n591));
  INV_X1    g405(.A(KEYINPUT25), .ZN(new_n592));
  NOR4_X1   g406(.A1(new_n588), .A2(new_n589), .A3(new_n592), .A4(G902), .ZN(new_n593));
  OAI21_X1  g407(.A(new_n569), .B1(new_n591), .B2(new_n593), .ZN(new_n594));
  NOR2_X1   g408(.A1(new_n569), .A2(G902), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n590), .A2(new_n595), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n594), .A2(new_n596), .ZN(new_n597));
  INV_X1    g411(.A(new_n597), .ZN(new_n598));
  NAND4_X1  g412(.A1(new_n303), .A2(new_n493), .A3(KEYINPUT96), .A4(new_n496), .ZN(new_n599));
  NAND4_X1  g413(.A1(new_n499), .A2(new_n566), .A3(new_n598), .A4(new_n599), .ZN(new_n600));
  XNOR2_X1  g414(.A(new_n600), .B(G101), .ZN(G3));
  NAND2_X1  g415(.A1(new_n303), .A2(new_n496), .ZN(new_n602));
  AND3_X1   g416(.A1(new_n552), .A2(new_n558), .A3(new_n559), .ZN(new_n603));
  AOI21_X1  g417(.A(new_n559), .B1(new_n552), .B2(new_n558), .ZN(new_n604));
  OAI21_X1  g418(.A(new_n562), .B1(new_n603), .B2(new_n604), .ZN(new_n605));
  AOI21_X1  g419(.A(G902), .B1(new_n551), .B2(new_n560), .ZN(new_n606));
  INV_X1    g420(.A(G472), .ZN(new_n607));
  OAI21_X1  g421(.A(new_n605), .B1(new_n606), .B2(new_n607), .ZN(new_n608));
  NOR3_X1   g422(.A1(new_n602), .A2(new_n608), .A3(new_n597), .ZN(new_n609));
  INV_X1    g423(.A(new_n431), .ZN(new_n610));
  INV_X1    g424(.A(new_n491), .ZN(new_n611));
  NAND3_X1  g425(.A1(new_n480), .A2(new_n488), .A3(new_n489), .ZN(new_n612));
  AOI21_X1  g426(.A(new_n610), .B1(new_n611), .B2(new_n612), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n613), .A2(new_n429), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n418), .A2(new_n423), .ZN(new_n615));
  INV_X1    g429(.A(KEYINPUT33), .ZN(new_n616));
  OAI21_X1  g430(.A(new_n616), .B1(new_n342), .B2(new_n343), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n617), .A2(KEYINPUT97), .ZN(new_n618));
  INV_X1    g432(.A(KEYINPUT97), .ZN(new_n619));
  OAI211_X1 g433(.A(new_n619), .B(new_n616), .C1(new_n342), .C2(new_n343), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n618), .A2(new_n620), .ZN(new_n621));
  NAND3_X1  g435(.A1(new_n348), .A2(KEYINPUT33), .A3(new_n349), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n622), .A2(KEYINPUT98), .ZN(new_n623));
  INV_X1    g437(.A(KEYINPUT98), .ZN(new_n624));
  NAND4_X1  g438(.A1(new_n348), .A2(new_n624), .A3(KEYINPUT33), .A4(new_n349), .ZN(new_n625));
  NAND2_X1  g439(.A1(new_n623), .A2(new_n625), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n621), .A2(new_n626), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n627), .A2(G478), .ZN(new_n628));
  NOR2_X1   g442(.A1(new_n304), .A2(new_n187), .ZN(new_n629));
  AOI21_X1  g443(.A(new_n629), .B1(new_n350), .B2(new_n304), .ZN(new_n630));
  NAND3_X1  g444(.A1(new_n615), .A2(new_n628), .A3(new_n630), .ZN(new_n631));
  NOR2_X1   g445(.A1(new_n614), .A2(new_n631), .ZN(new_n632));
  NAND2_X1  g446(.A1(new_n609), .A2(new_n632), .ZN(new_n633));
  XOR2_X1   g447(.A(KEYINPUT34), .B(G104), .Z(new_n634));
  XNOR2_X1  g448(.A(new_n633), .B(new_n634), .ZN(G6));
  INV_X1    g449(.A(KEYINPUT99), .ZN(new_n636));
  OR2_X1    g450(.A1(new_n411), .A2(new_n636), .ZN(new_n637));
  NAND3_X1  g451(.A1(new_n411), .A2(new_n417), .A3(new_n636), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  INV_X1    g453(.A(new_n639), .ZN(new_n640));
  INV_X1    g454(.A(new_n354), .ZN(new_n641));
  NAND3_X1  g455(.A1(new_n640), .A2(new_n641), .A3(new_n423), .ZN(new_n642));
  NOR2_X1   g456(.A1(new_n642), .A2(new_n614), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n609), .A2(new_n643), .ZN(new_n644));
  XOR2_X1   g458(.A(KEYINPUT35), .B(G107), .Z(new_n645));
  XNOR2_X1  g459(.A(new_n644), .B(new_n645), .ZN(G9));
  NOR2_X1   g460(.A1(new_n587), .A2(KEYINPUT36), .ZN(new_n647));
  XNOR2_X1  g461(.A(new_n583), .B(new_n647), .ZN(new_n648));
  NAND2_X1  g462(.A1(new_n648), .A2(new_n595), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n594), .A2(new_n649), .ZN(new_n650));
  OAI211_X1 g464(.A(new_n605), .B(new_n650), .C1(new_n606), .C2(new_n607), .ZN(new_n651));
  INV_X1    g465(.A(new_n651), .ZN(new_n652));
  NAND3_X1  g466(.A1(new_n499), .A2(new_n599), .A3(new_n652), .ZN(new_n653));
  XNOR2_X1  g467(.A(KEYINPUT37), .B(G110), .ZN(new_n654));
  XNOR2_X1  g468(.A(new_n653), .B(new_n654), .ZN(new_n655));
  XOR2_X1   g469(.A(KEYINPUT100), .B(KEYINPUT101), .Z(new_n656));
  XNOR2_X1  g470(.A(new_n655), .B(new_n656), .ZN(G12));
  NAND2_X1  g471(.A1(new_n257), .A2(new_n259), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n658), .A2(KEYINPUT82), .ZN(new_n659));
  NAND3_X1  g473(.A1(new_n257), .A2(new_n258), .A3(new_n259), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  AOI21_X1  g475(.A(new_n287), .B1(new_n661), .B2(new_n249), .ZN(new_n662));
  OAI211_X1 g476(.A(new_n299), .B(new_n187), .C1(new_n662), .C2(new_n296), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n663), .A2(KEYINPUT84), .ZN(new_n664));
  NAND3_X1  g478(.A1(new_n298), .A2(new_n293), .A3(new_n299), .ZN(new_n665));
  AOI22_X1  g479(.A1(new_n664), .A2(new_n665), .B1(G469), .B2(new_n291), .ZN(new_n666));
  OAI211_X1 g480(.A(new_n650), .B(new_n431), .C1(new_n491), .C2(new_n490), .ZN(new_n667));
  NOR3_X1   g481(.A1(new_n666), .A2(new_n495), .A3(new_n667), .ZN(new_n668));
  OR2_X1    g482(.A1(new_n428), .A2(G900), .ZN(new_n669));
  NAND2_X1  g483(.A1(new_n669), .A2(new_n425), .ZN(new_n670));
  NAND2_X1  g484(.A1(new_n423), .A2(new_n670), .ZN(new_n671));
  NOR3_X1   g485(.A1(new_n639), .A2(new_n354), .A3(new_n671), .ZN(new_n672));
  NAND3_X1  g486(.A1(new_n668), .A2(new_n566), .A3(new_n672), .ZN(new_n673));
  INV_X1    g487(.A(KEYINPUT102), .ZN(new_n674));
  NAND2_X1  g488(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  INV_X1    g489(.A(new_n672), .ZN(new_n676));
  NAND2_X1  g490(.A1(new_n605), .A2(KEYINPUT32), .ZN(new_n677));
  NAND3_X1  g491(.A1(new_n561), .A2(new_n544), .A3(new_n562), .ZN(new_n678));
  NAND2_X1  g492(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  AOI21_X1  g493(.A(new_n676), .B1(new_n679), .B2(new_n543), .ZN(new_n680));
  NAND3_X1  g494(.A1(new_n680), .A2(KEYINPUT102), .A3(new_n668), .ZN(new_n681));
  NAND2_X1  g495(.A1(new_n675), .A2(new_n681), .ZN(new_n682));
  XNOR2_X1  g496(.A(new_n682), .B(G128), .ZN(G30));
  NAND2_X1  g497(.A1(new_n516), .A2(new_n522), .ZN(new_n684));
  NAND2_X1  g498(.A1(new_n547), .A2(new_n531), .ZN(new_n685));
  NAND2_X1  g499(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  AOI21_X1  g500(.A(new_n607), .B1(new_n686), .B2(new_n187), .ZN(new_n687));
  AOI21_X1  g501(.A(new_n687), .B1(new_n677), .B2(new_n678), .ZN(new_n688));
  NOR2_X1   g502(.A1(new_n688), .A2(new_n650), .ZN(new_n689));
  NOR2_X1   g503(.A1(new_n490), .A2(new_n491), .ZN(new_n690));
  XNOR2_X1  g504(.A(new_n690), .B(KEYINPUT38), .ZN(new_n691));
  NAND2_X1  g505(.A1(new_n615), .A2(new_n641), .ZN(new_n692));
  NOR3_X1   g506(.A1(new_n691), .A2(new_n610), .A3(new_n692), .ZN(new_n693));
  NAND2_X1  g507(.A1(new_n689), .A2(new_n693), .ZN(new_n694));
  XOR2_X1   g508(.A(new_n694), .B(KEYINPUT103), .Z(new_n695));
  INV_X1    g509(.A(new_n602), .ZN(new_n696));
  XNOR2_X1  g510(.A(KEYINPUT104), .B(KEYINPUT39), .ZN(new_n697));
  XNOR2_X1  g511(.A(new_n670), .B(new_n697), .ZN(new_n698));
  NAND2_X1  g512(.A1(new_n696), .A2(new_n698), .ZN(new_n699));
  XNOR2_X1  g513(.A(new_n699), .B(KEYINPUT40), .ZN(new_n700));
  NOR2_X1   g514(.A1(new_n695), .A2(new_n700), .ZN(new_n701));
  XNOR2_X1  g515(.A(new_n701), .B(new_n211), .ZN(G45));
  AOI22_X1  g516(.A1(new_n620), .A2(new_n618), .B1(new_n623), .B2(new_n625), .ZN(new_n703));
  OAI21_X1  g517(.A(new_n630), .B1(new_n703), .B2(new_n304), .ZN(new_n704));
  AOI22_X1  g518(.A1(new_n411), .A2(new_n417), .B1(new_n420), .B2(new_n422), .ZN(new_n705));
  INV_X1    g519(.A(new_n670), .ZN(new_n706));
  NOR3_X1   g520(.A1(new_n704), .A2(new_n705), .A3(new_n706), .ZN(new_n707));
  NAND3_X1  g521(.A1(new_n668), .A2(new_n566), .A3(new_n707), .ZN(new_n708));
  XOR2_X1   g522(.A(KEYINPUT105), .B(G146), .Z(new_n709));
  XNOR2_X1  g523(.A(new_n708), .B(new_n709), .ZN(G48));
  AOI22_X1  g524(.A1(new_n677), .A2(new_n678), .B1(G472), .B2(new_n542), .ZN(new_n711));
  NOR2_X1   g525(.A1(new_n711), .A2(new_n597), .ZN(new_n712));
  OAI21_X1  g526(.A(G469), .B1(new_n301), .B2(G902), .ZN(new_n713));
  OAI211_X1 g527(.A(new_n496), .B(new_n713), .C1(new_n300), .C2(new_n302), .ZN(new_n714));
  INV_X1    g528(.A(KEYINPUT106), .ZN(new_n715));
  NAND2_X1  g529(.A1(new_n714), .A2(new_n715), .ZN(new_n716));
  NAND2_X1  g530(.A1(new_n664), .A2(new_n665), .ZN(new_n717));
  NAND4_X1  g531(.A1(new_n717), .A2(KEYINPUT106), .A3(new_n496), .A4(new_n713), .ZN(new_n718));
  AND2_X1   g532(.A1(new_n716), .A2(new_n718), .ZN(new_n719));
  NAND3_X1  g533(.A1(new_n712), .A2(new_n719), .A3(new_n632), .ZN(new_n720));
  XNOR2_X1  g534(.A(KEYINPUT41), .B(G113), .ZN(new_n721));
  XNOR2_X1  g535(.A(new_n720), .B(new_n721), .ZN(G15));
  NAND4_X1  g536(.A1(new_n566), .A2(new_n598), .A3(new_n716), .A4(new_n718), .ZN(new_n723));
  INV_X1    g537(.A(new_n643), .ZN(new_n724));
  OAI21_X1  g538(.A(KEYINPUT107), .B1(new_n723), .B2(new_n724), .ZN(new_n725));
  INV_X1    g539(.A(KEYINPUT107), .ZN(new_n726));
  NAND4_X1  g540(.A1(new_n712), .A2(new_n719), .A3(new_n726), .A4(new_n643), .ZN(new_n727));
  NAND2_X1  g541(.A1(new_n725), .A2(new_n727), .ZN(new_n728));
  XNOR2_X1  g542(.A(new_n728), .B(G116), .ZN(G18));
  NAND2_X1  g543(.A1(new_n650), .A2(new_n354), .ZN(new_n730));
  INV_X1    g544(.A(new_n429), .ZN(new_n731));
  NOR3_X1   g545(.A1(new_n730), .A2(new_n615), .A3(new_n731), .ZN(new_n732));
  NAND2_X1  g546(.A1(new_n566), .A2(new_n732), .ZN(new_n733));
  NAND3_X1  g547(.A1(new_n716), .A2(new_n613), .A3(new_n718), .ZN(new_n734));
  NOR2_X1   g548(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  XOR2_X1   g549(.A(new_n735), .B(G119), .Z(G21));
  OR2_X1    g550(.A1(new_n517), .A2(new_n521), .ZN(new_n737));
  AOI21_X1  g551(.A(new_n564), .B1(new_n737), .B2(new_n558), .ZN(new_n738));
  OAI21_X1  g552(.A(KEYINPUT108), .B1(new_n606), .B2(new_n607), .ZN(new_n739));
  OAI21_X1  g553(.A(new_n187), .B1(new_n603), .B2(new_n604), .ZN(new_n740));
  INV_X1    g554(.A(KEYINPUT108), .ZN(new_n741));
  NAND3_X1  g555(.A1(new_n740), .A2(new_n741), .A3(G472), .ZN(new_n742));
  AOI21_X1  g556(.A(new_n738), .B1(new_n739), .B2(new_n742), .ZN(new_n743));
  NAND2_X1  g557(.A1(new_n743), .A2(new_n598), .ZN(new_n744));
  NOR2_X1   g558(.A1(new_n614), .A2(new_n692), .ZN(new_n745));
  NAND3_X1  g559(.A1(new_n716), .A2(new_n718), .A3(new_n745), .ZN(new_n746));
  NOR2_X1   g560(.A1(new_n744), .A2(new_n746), .ZN(new_n747));
  XOR2_X1   g561(.A(new_n747), .B(G122), .Z(G24));
  AND3_X1   g562(.A1(new_n743), .A2(new_n650), .A3(new_n707), .ZN(new_n749));
  INV_X1    g563(.A(new_n734), .ZN(new_n750));
  NAND2_X1  g564(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  XOR2_X1   g565(.A(KEYINPUT109), .B(G125), .Z(new_n752));
  XNOR2_X1  g566(.A(new_n751), .B(new_n752), .ZN(G27));
  NAND2_X1  g567(.A1(new_n690), .A2(new_n431), .ZN(new_n754));
  NOR3_X1   g568(.A1(new_n666), .A2(new_n495), .A3(new_n754), .ZN(new_n755));
  NAND4_X1  g569(.A1(new_n755), .A2(new_n566), .A3(new_n598), .A4(new_n707), .ZN(new_n756));
  INV_X1    g570(.A(KEYINPUT42), .ZN(new_n757));
  NAND2_X1  g571(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  OAI21_X1  g572(.A(KEYINPUT110), .B1(new_n563), .B2(new_n565), .ZN(new_n759));
  INV_X1    g573(.A(KEYINPUT110), .ZN(new_n760));
  NAND3_X1  g574(.A1(new_n677), .A2(new_n678), .A3(new_n760), .ZN(new_n761));
  NAND3_X1  g575(.A1(new_n759), .A2(new_n761), .A3(new_n543), .ZN(new_n762));
  INV_X1    g576(.A(new_n754), .ZN(new_n763));
  NAND4_X1  g577(.A1(new_n303), .A2(new_n763), .A3(new_n496), .A4(new_n707), .ZN(new_n764));
  NOR2_X1   g578(.A1(new_n764), .A2(new_n757), .ZN(new_n765));
  NAND3_X1  g579(.A1(new_n762), .A2(new_n765), .A3(new_n598), .ZN(new_n766));
  NAND2_X1  g580(.A1(new_n758), .A2(new_n766), .ZN(new_n767));
  XNOR2_X1  g581(.A(new_n767), .B(G131), .ZN(G33));
  NAND4_X1  g582(.A1(new_n755), .A2(new_n566), .A3(new_n598), .A4(new_n672), .ZN(new_n769));
  XNOR2_X1  g583(.A(new_n769), .B(G134), .ZN(G36));
  INV_X1    g584(.A(new_n608), .ZN(new_n771));
  INV_X1    g585(.A(new_n650), .ZN(new_n772));
  NOR2_X1   g586(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  NOR2_X1   g587(.A1(new_n704), .A2(new_n615), .ZN(new_n774));
  XOR2_X1   g588(.A(KEYINPUT111), .B(KEYINPUT43), .Z(new_n775));
  NAND2_X1  g589(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  INV_X1    g590(.A(KEYINPUT43), .ZN(new_n777));
  OAI22_X1  g591(.A1(new_n704), .A2(new_n615), .B1(KEYINPUT111), .B2(new_n777), .ZN(new_n778));
  NAND2_X1  g592(.A1(new_n776), .A2(new_n778), .ZN(new_n779));
  INV_X1    g593(.A(new_n779), .ZN(new_n780));
  NOR2_X1   g594(.A1(new_n780), .A2(KEYINPUT112), .ZN(new_n781));
  AND3_X1   g595(.A1(new_n776), .A2(KEYINPUT112), .A3(new_n778), .ZN(new_n782));
  OAI21_X1  g596(.A(new_n773), .B1(new_n781), .B2(new_n782), .ZN(new_n783));
  INV_X1    g597(.A(KEYINPUT44), .ZN(new_n784));
  NOR2_X1   g598(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  INV_X1    g599(.A(KEYINPUT113), .ZN(new_n786));
  XNOR2_X1  g600(.A(new_n785), .B(new_n786), .ZN(new_n787));
  NOR2_X1   g601(.A1(new_n284), .A2(new_n290), .ZN(new_n788));
  OR2_X1    g602(.A1(new_n788), .A2(KEYINPUT45), .ZN(new_n789));
  NAND2_X1  g603(.A1(new_n788), .A2(KEYINPUT45), .ZN(new_n790));
  NAND3_X1  g604(.A1(new_n789), .A2(G469), .A3(new_n790), .ZN(new_n791));
  NAND2_X1  g605(.A1(G469), .A2(G902), .ZN(new_n792));
  NAND2_X1  g606(.A1(new_n791), .A2(new_n792), .ZN(new_n793));
  INV_X1    g607(.A(KEYINPUT46), .ZN(new_n794));
  AOI22_X1  g608(.A1(new_n793), .A2(new_n794), .B1(new_n665), .B2(new_n664), .ZN(new_n795));
  OAI21_X1  g609(.A(new_n795), .B1(new_n794), .B2(new_n793), .ZN(new_n796));
  AND3_X1   g610(.A1(new_n796), .A2(new_n496), .A3(new_n698), .ZN(new_n797));
  AOI21_X1  g611(.A(new_n754), .B1(new_n783), .B2(new_n784), .ZN(new_n798));
  NAND3_X1  g612(.A1(new_n787), .A2(new_n797), .A3(new_n798), .ZN(new_n799));
  XNOR2_X1  g613(.A(new_n799), .B(G137), .ZN(G39));
  AND3_X1   g614(.A1(new_n763), .A2(new_n597), .A3(new_n707), .ZN(new_n801));
  AND3_X1   g615(.A1(new_n796), .A2(KEYINPUT47), .A3(new_n496), .ZN(new_n802));
  AOI21_X1  g616(.A(KEYINPUT47), .B1(new_n796), .B2(new_n496), .ZN(new_n803));
  OAI211_X1 g617(.A(new_n711), .B(new_n801), .C1(new_n802), .C2(new_n803), .ZN(new_n804));
  XNOR2_X1  g618(.A(new_n804), .B(KEYINPUT114), .ZN(new_n805));
  XOR2_X1   g619(.A(KEYINPUT115), .B(G140), .Z(new_n806));
  XNOR2_X1  g620(.A(new_n805), .B(new_n806), .ZN(G42));
  AND2_X1   g621(.A1(new_n717), .A2(new_n713), .ZN(new_n808));
  XNOR2_X1  g622(.A(new_n808), .B(KEYINPUT49), .ZN(new_n809));
  AND4_X1   g623(.A1(new_n598), .A2(new_n774), .A3(new_n496), .A4(new_n431), .ZN(new_n810));
  NAND4_X1  g624(.A1(new_n809), .A2(new_n688), .A3(new_n691), .A4(new_n810), .ZN(new_n811));
  INV_X1    g625(.A(new_n632), .ZN(new_n812));
  OAI22_X1  g626(.A1(new_n723), .A2(new_n812), .B1(new_n733), .B2(new_n734), .ZN(new_n813));
  NOR2_X1   g627(.A1(new_n813), .A2(new_n747), .ZN(new_n814));
  AND2_X1   g628(.A1(new_n814), .A2(new_n728), .ZN(new_n815));
  OAI21_X1  g629(.A(KEYINPUT116), .B1(new_n615), .B2(new_n354), .ZN(new_n816));
  INV_X1    g630(.A(KEYINPUT116), .ZN(new_n817));
  NAND3_X1  g631(.A1(new_n641), .A2(new_n705), .A3(new_n817), .ZN(new_n818));
  NAND3_X1  g632(.A1(new_n816), .A2(new_n631), .A3(new_n818), .ZN(new_n819));
  INV_X1    g633(.A(new_n614), .ZN(new_n820));
  AND2_X1   g634(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  NAND4_X1  g635(.A1(new_n821), .A2(new_n598), .A3(new_n696), .A4(new_n771), .ZN(new_n822));
  AND3_X1   g636(.A1(new_n600), .A2(new_n822), .A3(new_n653), .ZN(new_n823));
  INV_X1    g637(.A(new_n764), .ZN(new_n824));
  NAND3_X1  g638(.A1(new_n824), .A2(new_n743), .A3(new_n650), .ZN(new_n825));
  NOR3_X1   g639(.A1(new_n730), .A2(new_n639), .A3(new_n671), .ZN(new_n826));
  NAND3_X1  g640(.A1(new_n755), .A2(new_n566), .A3(new_n826), .ZN(new_n827));
  AND3_X1   g641(.A1(new_n825), .A2(new_n769), .A3(new_n827), .ZN(new_n828));
  AND3_X1   g642(.A1(new_n823), .A2(new_n767), .A3(new_n828), .ZN(new_n829));
  AOI21_X1  g643(.A(KEYINPUT102), .B1(new_n680), .B2(new_n668), .ZN(new_n830));
  AND4_X1   g644(.A1(KEYINPUT102), .A2(new_n668), .A3(new_n566), .A4(new_n672), .ZN(new_n831));
  OAI21_X1  g645(.A(new_n708), .B1(new_n830), .B2(new_n831), .ZN(new_n832));
  NAND3_X1  g646(.A1(new_n613), .A2(new_n641), .A3(new_n615), .ZN(new_n833));
  NOR3_X1   g647(.A1(new_n602), .A2(new_n706), .A3(new_n833), .ZN(new_n834));
  NAND2_X1  g648(.A1(new_n689), .A2(new_n834), .ZN(new_n835));
  NAND3_X1  g649(.A1(new_n743), .A2(new_n650), .A3(new_n707), .ZN(new_n836));
  OAI21_X1  g650(.A(new_n835), .B1(new_n836), .B2(new_n734), .ZN(new_n837));
  INV_X1    g651(.A(KEYINPUT52), .ZN(new_n838));
  NOR3_X1   g652(.A1(new_n832), .A2(new_n837), .A3(new_n838), .ZN(new_n839));
  INV_X1    g653(.A(new_n708), .ZN(new_n840));
  AOI21_X1  g654(.A(new_n840), .B1(new_n675), .B2(new_n681), .ZN(new_n841));
  AOI22_X1  g655(.A1(new_n749), .A2(new_n750), .B1(new_n689), .B2(new_n834), .ZN(new_n842));
  AOI21_X1  g656(.A(KEYINPUT52), .B1(new_n841), .B2(new_n842), .ZN(new_n843));
  OAI211_X1 g657(.A(new_n815), .B(new_n829), .C1(new_n839), .C2(new_n843), .ZN(new_n844));
  INV_X1    g658(.A(KEYINPUT53), .ZN(new_n845));
  XNOR2_X1  g659(.A(new_n844), .B(new_n845), .ZN(new_n846));
  INV_X1    g660(.A(KEYINPUT117), .ZN(new_n847));
  NAND3_X1  g661(.A1(new_n846), .A2(new_n847), .A3(KEYINPUT54), .ZN(new_n848));
  NAND2_X1  g662(.A1(new_n844), .A2(new_n845), .ZN(new_n849));
  INV_X1    g663(.A(KEYINPUT118), .ZN(new_n850));
  AND3_X1   g664(.A1(new_n814), .A2(new_n850), .A3(new_n728), .ZN(new_n851));
  AOI21_X1  g665(.A(new_n850), .B1(new_n814), .B2(new_n728), .ZN(new_n852));
  NOR2_X1   g666(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  NAND4_X1  g667(.A1(new_n823), .A2(new_n767), .A3(new_n828), .A4(KEYINPUT53), .ZN(new_n854));
  OAI21_X1  g668(.A(new_n838), .B1(new_n832), .B2(new_n837), .ZN(new_n855));
  NAND3_X1  g669(.A1(new_n841), .A2(new_n842), .A3(KEYINPUT52), .ZN(new_n856));
  AOI21_X1  g670(.A(new_n854), .B1(new_n855), .B2(new_n856), .ZN(new_n857));
  NAND2_X1  g671(.A1(new_n853), .A2(new_n857), .ZN(new_n858));
  NAND2_X1  g672(.A1(new_n849), .A2(new_n858), .ZN(new_n859));
  OAI21_X1  g673(.A(new_n848), .B1(KEYINPUT54), .B2(new_n859), .ZN(new_n860));
  NAND3_X1  g674(.A1(new_n719), .A2(new_n610), .A3(new_n691), .ZN(new_n861));
  INV_X1    g675(.A(KEYINPUT119), .ZN(new_n862));
  OR2_X1    g676(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  NAND2_X1  g677(.A1(new_n861), .A2(new_n862), .ZN(new_n864));
  NOR3_X1   g678(.A1(new_n744), .A2(new_n425), .A3(new_n780), .ZN(new_n865));
  NAND3_X1  g679(.A1(new_n863), .A2(new_n864), .A3(new_n865), .ZN(new_n866));
  XOR2_X1   g680(.A(new_n866), .B(KEYINPUT50), .Z(new_n867));
  AND2_X1   g681(.A1(new_n719), .A2(new_n763), .ZN(new_n868));
  NOR2_X1   g682(.A1(new_n597), .A2(new_n425), .ZN(new_n869));
  AND3_X1   g683(.A1(new_n868), .A2(new_n688), .A3(new_n869), .ZN(new_n870));
  NAND3_X1  g684(.A1(new_n870), .A2(new_n705), .A3(new_n704), .ZN(new_n871));
  XNOR2_X1  g685(.A(new_n871), .B(KEYINPUT120), .ZN(new_n872));
  OR2_X1    g686(.A1(new_n802), .A2(new_n803), .ZN(new_n873));
  AND2_X1   g687(.A1(new_n808), .A2(new_n495), .ZN(new_n874));
  OAI211_X1 g688(.A(new_n763), .B(new_n865), .C1(new_n873), .C2(new_n874), .ZN(new_n875));
  NOR2_X1   g689(.A1(new_n780), .A2(new_n425), .ZN(new_n876));
  NAND4_X1  g690(.A1(new_n868), .A2(new_n650), .A3(new_n743), .A4(new_n876), .ZN(new_n877));
  NAND4_X1  g691(.A1(new_n867), .A2(new_n872), .A3(new_n875), .A4(new_n877), .ZN(new_n878));
  INV_X1    g692(.A(KEYINPUT51), .ZN(new_n879));
  NAND2_X1  g693(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  NAND2_X1  g694(.A1(new_n865), .A2(new_n750), .ZN(new_n881));
  NAND3_X1  g695(.A1(new_n881), .A2(G952), .A3(new_n339), .ZN(new_n882));
  NAND4_X1  g696(.A1(new_n868), .A2(new_n598), .A3(new_n762), .A4(new_n876), .ZN(new_n883));
  XOR2_X1   g697(.A(new_n883), .B(KEYINPUT48), .Z(new_n884));
  INV_X1    g698(.A(new_n631), .ZN(new_n885));
  AOI211_X1 g699(.A(new_n882), .B(new_n884), .C1(new_n885), .C2(new_n870), .ZN(new_n886));
  NAND2_X1  g700(.A1(new_n880), .A2(new_n886), .ZN(new_n887));
  AOI21_X1  g701(.A(new_n847), .B1(new_n846), .B2(KEYINPUT54), .ZN(new_n888));
  NOR2_X1   g702(.A1(new_n878), .A2(new_n879), .ZN(new_n889));
  NOR4_X1   g703(.A1(new_n860), .A2(new_n887), .A3(new_n888), .A4(new_n889), .ZN(new_n890));
  NOR2_X1   g704(.A1(G952), .A2(G953), .ZN(new_n891));
  OAI21_X1  g705(.A(new_n811), .B1(new_n890), .B2(new_n891), .ZN(G75));
  NOR2_X1   g706(.A1(new_n339), .A2(G952), .ZN(new_n893));
  INV_X1    g707(.A(new_n893), .ZN(new_n894));
  AOI22_X1  g708(.A1(new_n845), .A2(new_n844), .B1(new_n853), .B2(new_n857), .ZN(new_n895));
  NOR2_X1   g709(.A1(new_n895), .A2(new_n187), .ZN(new_n896));
  AOI21_X1  g710(.A(KEYINPUT56), .B1(new_n896), .B2(G210), .ZN(new_n897));
  AND2_X1   g711(.A1(new_n484), .A2(new_n487), .ZN(new_n898));
  XNOR2_X1  g712(.A(new_n898), .B(new_n485), .ZN(new_n899));
  XOR2_X1   g713(.A(new_n899), .B(KEYINPUT55), .Z(new_n900));
  OAI21_X1  g714(.A(new_n894), .B1(new_n897), .B2(new_n900), .ZN(new_n901));
  NAND2_X1  g715(.A1(new_n896), .A2(KEYINPUT121), .ZN(new_n902));
  INV_X1    g716(.A(new_n489), .ZN(new_n903));
  INV_X1    g717(.A(KEYINPUT121), .ZN(new_n904));
  OAI21_X1  g718(.A(new_n904), .B1(new_n895), .B2(new_n187), .ZN(new_n905));
  NAND3_X1  g719(.A1(new_n902), .A2(new_n903), .A3(new_n905), .ZN(new_n906));
  INV_X1    g720(.A(KEYINPUT56), .ZN(new_n907));
  AND2_X1   g721(.A1(new_n900), .A2(new_n907), .ZN(new_n908));
  AOI21_X1  g722(.A(new_n901), .B1(new_n906), .B2(new_n908), .ZN(G51));
  XNOR2_X1  g723(.A(new_n859), .B(KEYINPUT54), .ZN(new_n910));
  XOR2_X1   g724(.A(new_n792), .B(KEYINPUT57), .Z(new_n911));
  NAND2_X1  g725(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  OAI21_X1  g726(.A(new_n912), .B1(new_n662), .B2(new_n296), .ZN(new_n913));
  INV_X1    g727(.A(new_n791), .ZN(new_n914));
  NAND3_X1  g728(.A1(new_n902), .A2(new_n914), .A3(new_n905), .ZN(new_n915));
  AOI21_X1  g729(.A(new_n893), .B1(new_n913), .B2(new_n915), .ZN(G54));
  NAND4_X1  g730(.A1(new_n902), .A2(KEYINPUT58), .A3(G475), .A4(new_n905), .ZN(new_n917));
  AND2_X1   g731(.A1(new_n917), .A2(new_n408), .ZN(new_n918));
  NOR2_X1   g732(.A1(new_n917), .A2(new_n408), .ZN(new_n919));
  NOR3_X1   g733(.A1(new_n918), .A2(new_n919), .A3(new_n893), .ZN(G60));
  XNOR2_X1  g734(.A(new_n629), .B(KEYINPUT59), .ZN(new_n921));
  INV_X1    g735(.A(new_n921), .ZN(new_n922));
  AND3_X1   g736(.A1(new_n910), .A2(new_n703), .A3(new_n922), .ZN(new_n923));
  OAI21_X1  g737(.A(new_n922), .B1(new_n860), .B2(new_n888), .ZN(new_n924));
  AOI211_X1 g738(.A(new_n893), .B(new_n923), .C1(new_n627), .C2(new_n924), .ZN(G63));
  XNOR2_X1  g739(.A(KEYINPUT122), .B(KEYINPUT61), .ZN(new_n926));
  NAND2_X1  g740(.A1(G217), .A2(G902), .ZN(new_n927));
  XNOR2_X1  g741(.A(new_n927), .B(KEYINPUT60), .ZN(new_n928));
  OAI21_X1  g742(.A(KEYINPUT123), .B1(new_n895), .B2(new_n928), .ZN(new_n929));
  INV_X1    g743(.A(new_n590), .ZN(new_n930));
  INV_X1    g744(.A(KEYINPUT123), .ZN(new_n931));
  INV_X1    g745(.A(new_n928), .ZN(new_n932));
  NAND2_X1  g746(.A1(new_n855), .A2(new_n856), .ZN(new_n933));
  INV_X1    g747(.A(new_n852), .ZN(new_n934));
  INV_X1    g748(.A(new_n854), .ZN(new_n935));
  NAND3_X1  g749(.A1(new_n814), .A2(new_n850), .A3(new_n728), .ZN(new_n936));
  AND4_X1   g750(.A1(new_n933), .A2(new_n934), .A3(new_n935), .A4(new_n936), .ZN(new_n937));
  NAND2_X1  g751(.A1(new_n814), .A2(new_n728), .ZN(new_n938));
  NAND3_X1  g752(.A1(new_n823), .A2(new_n767), .A3(new_n828), .ZN(new_n939));
  NOR2_X1   g753(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  AOI21_X1  g754(.A(KEYINPUT53), .B1(new_n940), .B2(new_n933), .ZN(new_n941));
  OAI211_X1 g755(.A(new_n931), .B(new_n932), .C1(new_n937), .C2(new_n941), .ZN(new_n942));
  NAND3_X1  g756(.A1(new_n929), .A2(new_n930), .A3(new_n942), .ZN(new_n943));
  NAND3_X1  g757(.A1(new_n943), .A2(KEYINPUT124), .A3(new_n894), .ZN(new_n944));
  NAND2_X1  g758(.A1(new_n929), .A2(new_n942), .ZN(new_n945));
  NAND2_X1  g759(.A1(new_n945), .A2(new_n648), .ZN(new_n946));
  NAND2_X1  g760(.A1(new_n944), .A2(new_n946), .ZN(new_n947));
  AOI21_X1  g761(.A(KEYINPUT124), .B1(new_n943), .B2(new_n894), .ZN(new_n948));
  OAI21_X1  g762(.A(new_n926), .B1(new_n947), .B2(new_n948), .ZN(new_n949));
  NAND4_X1  g763(.A1(new_n946), .A2(KEYINPUT61), .A3(new_n894), .A4(new_n943), .ZN(new_n950));
  NAND2_X1  g764(.A1(new_n949), .A2(new_n950), .ZN(G66));
  AOI21_X1  g765(.A(new_n339), .B1(new_n427), .B2(G224), .ZN(new_n952));
  NAND2_X1  g766(.A1(new_n815), .A2(new_n823), .ZN(new_n953));
  AOI21_X1  g767(.A(new_n952), .B1(new_n953), .B2(new_n339), .ZN(new_n954));
  INV_X1    g768(.A(G898), .ZN(new_n955));
  AOI21_X1  g769(.A(new_n898), .B1(new_n955), .B2(G953), .ZN(new_n956));
  XNOR2_X1  g770(.A(new_n954), .B(new_n956), .ZN(G69));
  NAND2_X1  g771(.A1(new_n526), .A2(new_n530), .ZN(new_n958));
  XNOR2_X1  g772(.A(new_n958), .B(new_n395), .ZN(new_n959));
  INV_X1    g773(.A(new_n699), .ZN(new_n960));
  NAND4_X1  g774(.A1(new_n960), .A2(new_n712), .A3(new_n763), .A4(new_n819), .ZN(new_n961));
  NAND2_X1  g775(.A1(new_n799), .A2(new_n961), .ZN(new_n962));
  NOR2_X1   g776(.A1(new_n962), .A2(new_n805), .ZN(new_n963));
  NAND2_X1  g777(.A1(new_n841), .A2(new_n751), .ZN(new_n964));
  XNOR2_X1  g778(.A(new_n964), .B(KEYINPUT125), .ZN(new_n965));
  OAI21_X1  g779(.A(KEYINPUT62), .B1(new_n965), .B2(new_n701), .ZN(new_n966));
  OR3_X1    g780(.A1(new_n965), .A2(KEYINPUT62), .A3(new_n701), .ZN(new_n967));
  NAND3_X1  g781(.A1(new_n963), .A2(new_n966), .A3(new_n967), .ZN(new_n968));
  AOI21_X1  g782(.A(new_n959), .B1(new_n968), .B2(new_n339), .ZN(new_n969));
  INV_X1    g783(.A(G900), .ZN(new_n970));
  OAI21_X1  g784(.A(new_n959), .B1(new_n970), .B2(new_n339), .ZN(new_n971));
  INV_X1    g785(.A(new_n833), .ZN(new_n972));
  NAND4_X1  g786(.A1(new_n797), .A2(new_n598), .A3(new_n762), .A4(new_n972), .ZN(new_n973));
  NAND4_X1  g787(.A1(new_n799), .A2(new_n767), .A3(new_n769), .A4(new_n973), .ZN(new_n974));
  NOR3_X1   g788(.A1(new_n974), .A2(new_n805), .A3(new_n965), .ZN(new_n975));
  AOI21_X1  g789(.A(new_n971), .B1(new_n975), .B2(new_n339), .ZN(new_n976));
  NOR2_X1   g790(.A1(new_n969), .A2(new_n976), .ZN(new_n977));
  OAI21_X1  g791(.A(G953), .B1(new_n189), .B2(new_n970), .ZN(new_n978));
  XNOR2_X1  g792(.A(new_n977), .B(new_n978), .ZN(G72));
  XNOR2_X1  g793(.A(new_n532), .B(KEYINPUT126), .ZN(new_n980));
  NOR2_X1   g794(.A1(new_n980), .A2(new_n521), .ZN(new_n981));
  NOR4_X1   g795(.A1(new_n974), .A2(new_n805), .A3(new_n953), .A4(new_n965), .ZN(new_n982));
  NAND2_X1  g796(.A1(G472), .A2(G902), .ZN(new_n983));
  XOR2_X1   g797(.A(new_n983), .B(KEYINPUT63), .Z(new_n984));
  INV_X1    g798(.A(new_n984), .ZN(new_n985));
  OAI21_X1  g799(.A(new_n981), .B1(new_n982), .B2(new_n985), .ZN(new_n986));
  AOI21_X1  g800(.A(new_n985), .B1(new_n533), .B2(new_n685), .ZN(new_n987));
  AOI21_X1  g801(.A(new_n893), .B1(new_n846), .B2(new_n987), .ZN(new_n988));
  NAND2_X1  g802(.A1(new_n986), .A2(new_n988), .ZN(new_n989));
  NAND2_X1  g803(.A1(new_n980), .A2(new_n521), .ZN(new_n990));
  INV_X1    g804(.A(new_n953), .ZN(new_n991));
  NAND4_X1  g805(.A1(new_n963), .A2(new_n966), .A3(new_n991), .A4(new_n967), .ZN(new_n992));
  AOI21_X1  g806(.A(new_n990), .B1(new_n992), .B2(new_n984), .ZN(new_n993));
  OAI21_X1  g807(.A(KEYINPUT127), .B1(new_n989), .B2(new_n993), .ZN(new_n994));
  INV_X1    g808(.A(new_n993), .ZN(new_n995));
  INV_X1    g809(.A(KEYINPUT127), .ZN(new_n996));
  NAND4_X1  g810(.A1(new_n995), .A2(new_n996), .A3(new_n986), .A4(new_n988), .ZN(new_n997));
  NAND2_X1  g811(.A1(new_n994), .A2(new_n997), .ZN(G57));
endmodule


