

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361,
         n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372,
         n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383,
         n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394,
         n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405,
         n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416,
         n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427,
         n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438,
         n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449,
         n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460,
         n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471,
         n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482,
         n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493,
         n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504,
         n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515,
         n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526,
         n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537,
         n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
         n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559,
         n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570,
         n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581,
         n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592,
         n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603,
         n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614,
         n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625,
         n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636,
         n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647,
         n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658,
         n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669,
         n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680,
         n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691,
         n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702,
         n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713,
         n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724,
         n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735,
         n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746,
         n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757,
         n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768,
         n769, n770, n771, n772, n773, n774, n775, n776;

  OR2_X1 U373 ( .A1(n723), .A2(n383), .ZN(n389) );
  AND2_X1 U374 ( .A1(n550), .A2(n687), .ZN(n354) );
  AND2_X1 U375 ( .A1(n611), .A2(n610), .ZN(n612) );
  XNOR2_X1 U376 ( .A(n697), .B(KEYINPUT6), .ZN(n610) );
  XNOR2_X1 U377 ( .A(n455), .B(n454), .ZN(n513) );
  INV_X1 U378 ( .A(KEYINPUT3), .ZN(n453) );
  NAND2_X2 U379 ( .A1(n579), .A2(n580), .ZN(n582) );
  XNOR2_X1 U380 ( .A(n622), .B(KEYINPUT39), .ZN(n627) );
  XOR2_X1 U381 ( .A(n514), .B(n513), .Z(n351) );
  BUF_X2 U382 ( .A(n596), .Z(n697) );
  AND2_X1 U383 ( .A1(n614), .A2(n550), .ZN(n749) );
  XNOR2_X2 U384 ( .A(n600), .B(KEYINPUT110), .ZN(n617) );
  AND2_X2 U385 ( .A1(n409), .A2(n547), .ZN(n651) );
  OR2_X2 U386 ( .A1(n613), .A2(n356), .ZN(n628) );
  XNOR2_X2 U387 ( .A(n560), .B(KEYINPUT101), .ZN(n590) );
  XNOR2_X2 U388 ( .A(n554), .B(KEYINPUT35), .ZN(n774) );
  XNOR2_X2 U389 ( .A(n459), .B(n759), .ZN(n638) );
  NOR2_X2 U390 ( .A1(n387), .A2(n385), .ZN(n554) );
  AND2_X2 U391 ( .A1(n578), .A2(n360), .ZN(n579) );
  XNOR2_X2 U392 ( .A(n457), .B(n458), .ZN(n759) );
  OR2_X2 U393 ( .A1(n774), .A2(n555), .ZN(n557) );
  XNOR2_X2 U394 ( .A(n552), .B(n551), .ZN(n723) );
  AND2_X2 U395 ( .A1(n610), .A2(n354), .ZN(n552) );
  INV_X1 U396 ( .A(G953), .ZN(n767) );
  INV_X2 U397 ( .A(n668), .ZN(n675) );
  OR2_X1 U398 ( .A1(n621), .A2(n620), .ZN(n622) );
  NAND2_X1 U399 ( .A1(n420), .A2(n418), .ZN(n417) );
  AND2_X1 U400 ( .A1(n424), .A2(n422), .ZN(n421) );
  NAND2_X1 U401 ( .A1(n401), .A2(n633), .ZN(n390) );
  XNOR2_X1 U402 ( .A(n402), .B(n626), .ZN(n401) );
  NAND2_X1 U403 ( .A1(n404), .A2(n403), .ZN(n402) );
  NOR2_X1 U404 ( .A1(n776), .A2(n650), .ZN(n625) );
  AND2_X1 U405 ( .A1(n593), .A2(n592), .ZN(n605) );
  NAND2_X1 U406 ( .A1(n440), .A2(n594), .ZN(n621) );
  XNOR2_X1 U407 ( .A(n499), .B(G478), .ZN(n569) );
  XNOR2_X1 U408 ( .A(n489), .B(n488), .ZN(n570) );
  XOR2_X1 U409 ( .A(G146), .B(G125), .Z(n477) );
  XNOR2_X2 U410 ( .A(n352), .B(n353), .ZN(n598) );
  NOR2_X1 U411 ( .A1(n678), .A2(G902), .ZN(n352) );
  XOR2_X1 U412 ( .A(n523), .B(G469), .Z(n353) );
  INV_X1 U413 ( .A(n390), .ZN(n420) );
  XNOR2_X1 U414 ( .A(n453), .B(G113), .ZN(n455) );
  INV_X1 U415 ( .A(G128), .ZN(n447) );
  XNOR2_X1 U416 ( .A(n376), .B(n462), .ZN(n587) );
  NOR2_X1 U417 ( .A1(n570), .A2(n567), .ZN(n589) );
  BUF_X1 U418 ( .A(n587), .Z(n426) );
  INV_X1 U419 ( .A(KEYINPUT87), .ZN(n398) );
  INV_X1 U420 ( .A(KEYINPUT47), .ZN(n406) );
  NAND2_X1 U421 ( .A1(n408), .A2(n366), .ZN(n407) );
  INV_X1 U422 ( .A(n602), .ZN(n408) );
  OR2_X2 U423 ( .A1(n735), .A2(n741), .ZN(n371) );
  XNOR2_X1 U424 ( .A(n431), .B(n363), .ZN(n601) );
  NOR2_X1 U425 ( .A1(n587), .A2(n432), .ZN(n431) );
  XNOR2_X1 U426 ( .A(n493), .B(n492), .ZN(n494) );
  INV_X1 U427 ( .A(KEYINPUT7), .ZN(n373) );
  INV_X1 U428 ( .A(G134), .ZN(n495) );
  XNOR2_X1 U429 ( .A(n428), .B(n427), .ZN(n704) );
  INV_X1 U430 ( .A(KEYINPUT41), .ZN(n427) );
  NOR2_X1 U431 ( .A1(n711), .A2(n710), .ZN(n428) );
  XNOR2_X1 U432 ( .A(n544), .B(n382), .ZN(n381) );
  INV_X1 U433 ( .A(KEYINPUT106), .ZN(n382) );
  NAND2_X1 U434 ( .A1(n590), .A2(n358), .ZN(n591) );
  INV_X1 U435 ( .A(n426), .ZN(n588) );
  XNOR2_X1 U436 ( .A(n487), .B(n667), .ZN(n488) );
  INV_X1 U437 ( .A(n610), .ZN(n437) );
  INV_X1 U438 ( .A(n591), .ZN(n400) );
  XNOR2_X1 U439 ( .A(n442), .B(n441), .ZN(n440) );
  INV_X1 U440 ( .A(KEYINPUT30), .ZN(n441) );
  NAND2_X1 U441 ( .A1(n369), .A2(n708), .ZN(n442) );
  NOR2_X1 U442 ( .A1(n621), .A2(n398), .ZN(n394) );
  AND2_X1 U443 ( .A1(n397), .A2(n396), .ZN(n395) );
  AND2_X1 U444 ( .A1(n407), .A2(n405), .ZN(n374) );
  NAND2_X1 U445 ( .A1(n603), .A2(n406), .ZN(n405) );
  NAND2_X1 U446 ( .A1(n378), .A2(n362), .ZN(n377) );
  NOR2_X1 U447 ( .A1(KEYINPUT47), .A2(n607), .ZN(n608) );
  XNOR2_X1 U448 ( .A(n371), .B(n370), .ZN(n607) );
  INV_X1 U449 ( .A(KEYINPUT86), .ZN(n370) );
  INV_X1 U450 ( .A(n371), .ZN(n712) );
  NAND2_X1 U451 ( .A1(G234), .A2(G237), .ZN(n464) );
  NOR2_X1 U452 ( .A1(n596), .A2(n609), .ZN(n597) );
  XNOR2_X1 U453 ( .A(n368), .B(KEYINPUT8), .ZN(n491) );
  INV_X1 U454 ( .A(KEYINPUT88), .ZN(n368) );
  NOR2_X1 U455 ( .A1(G953), .A2(G237), .ZN(n508) );
  XNOR2_X1 U456 ( .A(KEYINPUT66), .B(G101), .ZN(n506) );
  XNOR2_X1 U457 ( .A(n477), .B(n503), .ZN(n445) );
  XNOR2_X1 U458 ( .A(KEYINPUT18), .B(KEYINPUT17), .ZN(n443) );
  XOR2_X1 U459 ( .A(KEYINPUT93), .B(KEYINPUT78), .Z(n444) );
  AND2_X1 U460 ( .A1(n419), .A2(KEYINPUT2), .ZN(n418) );
  INV_X1 U461 ( .A(KEYINPUT89), .ZN(n419) );
  NAND2_X1 U462 ( .A1(n423), .A2(KEYINPUT89), .ZN(n422) );
  INV_X1 U463 ( .A(KEYINPUT2), .ZN(n423) );
  XNOR2_X1 U464 ( .A(n426), .B(KEYINPUT38), .ZN(n707) );
  AND2_X1 U465 ( .A1(n693), .A2(n692), .ZN(n687) );
  INV_X1 U466 ( .A(G237), .ZN(n460) );
  INV_X1 U467 ( .A(G902), .ZN(n535) );
  NOR2_X1 U468 ( .A1(n601), .A2(n468), .ZN(n469) );
  XNOR2_X1 U469 ( .A(n522), .B(n351), .ZN(n515) );
  XNOR2_X1 U470 ( .A(KEYINPUT98), .B(KEYINPUT23), .ZN(n529) );
  XNOR2_X1 U471 ( .A(KEYINPUT68), .B(KEYINPUT10), .ZN(n476) );
  XNOR2_X1 U472 ( .A(G902), .B(KEYINPUT15), .ZN(n635) );
  INV_X1 U473 ( .A(n704), .ZN(n722) );
  BUF_X1 U474 ( .A(n549), .Z(n565) );
  INV_X1 U475 ( .A(n769), .ZN(n391) );
  XNOR2_X1 U476 ( .A(n498), .B(n372), .ZN(n663) );
  XNOR2_X1 U477 ( .A(n494), .B(n373), .ZN(n372) );
  XOR2_X1 U478 ( .A(G116), .B(G107), .Z(n497) );
  XNOR2_X1 U479 ( .A(n638), .B(n639), .ZN(n640) );
  XNOR2_X1 U480 ( .A(n643), .B(KEYINPUT92), .ZN(n681) );
  AND2_X1 U481 ( .A1(n631), .A2(n426), .ZN(n752) );
  NAND2_X1 U482 ( .A1(n704), .A2(n378), .ZN(n619) );
  XNOR2_X1 U483 ( .A(n624), .B(n623), .ZN(n650) );
  XNOR2_X1 U484 ( .A(n430), .B(KEYINPUT36), .ZN(n614) );
  NOR2_X2 U485 ( .A1(n628), .A2(n426), .ZN(n430) );
  NAND2_X1 U486 ( .A1(n386), .A2(n357), .ZN(n385) );
  XNOR2_X1 U487 ( .A(n411), .B(n367), .ZN(n775) );
  NAND2_X1 U488 ( .A1(n381), .A2(n437), .ZN(n380) );
  XNOR2_X1 U489 ( .A(n568), .B(KEYINPUT105), .ZN(n735) );
  OR2_X1 U490 ( .A1(n570), .A2(n569), .ZN(n744) );
  NAND2_X1 U491 ( .A1(n438), .A2(n437), .ZN(n574) );
  INV_X1 U492 ( .A(n621), .ZN(n392) );
  AND2_X1 U493 ( .A1(n378), .A2(n602), .ZN(n355) );
  OR2_X1 U494 ( .A1(n744), .A2(n432), .ZN(n356) );
  XOR2_X1 U495 ( .A(KEYINPUT79), .B(n589), .Z(n357) );
  AND2_X1 U496 ( .A1(n589), .A2(n588), .ZN(n358) );
  OR2_X1 U497 ( .A1(G953), .A2(n720), .ZN(n359) );
  AND2_X1 U498 ( .A1(n577), .A2(n576), .ZN(n360) );
  OR2_X1 U499 ( .A1(n584), .A2(G900), .ZN(n361) );
  AND2_X1 U500 ( .A1(n602), .A2(n603), .ZN(n362) );
  XOR2_X1 U501 ( .A(KEYINPUT65), .B(KEYINPUT19), .Z(n363) );
  INV_X1 U502 ( .A(n708), .ZN(n432) );
  XOR2_X1 U503 ( .A(KEYINPUT109), .B(KEYINPUT28), .Z(n364) );
  XOR2_X1 U504 ( .A(n553), .B(KEYINPUT80), .Z(n365) );
  AND2_X1 U505 ( .A1(KEYINPUT85), .A2(KEYINPUT47), .ZN(n366) );
  XOR2_X1 U506 ( .A(KEYINPUT81), .B(KEYINPUT32), .Z(n367) );
  INV_X1 U507 ( .A(n596), .ZN(n369) );
  XNOR2_X2 U508 ( .A(n516), .B(n652), .ZN(n596) );
  NOR2_X1 U509 ( .A1(n756), .A2(n390), .ZN(n634) );
  INV_X1 U510 ( .A(n569), .ZN(n567) );
  NAND2_X1 U511 ( .A1(n569), .A2(n570), .ZN(n568) );
  NAND2_X1 U512 ( .A1(n389), .A2(n388), .ZN(n387) );
  NAND2_X1 U513 ( .A1(n515), .A2(n535), .ZN(n516) );
  INV_X1 U514 ( .A(n515), .ZN(n654) );
  XNOR2_X2 U515 ( .A(n765), .B(n507), .ZN(n522) );
  XNOR2_X2 U516 ( .A(n505), .B(n504), .ZN(n765) );
  AND2_X1 U517 ( .A1(n375), .A2(n374), .ZN(n379) );
  NAND2_X1 U518 ( .A1(n617), .A2(n366), .ZN(n375) );
  NAND2_X1 U519 ( .A1(n638), .A2(n635), .ZN(n376) );
  NAND2_X1 U520 ( .A1(n379), .A2(n377), .ZN(n604) );
  INV_X1 U521 ( .A(n617), .ZN(n378) );
  NOR2_X1 U522 ( .A1(n546), .A2(n380), .ZN(n411) );
  INV_X1 U523 ( .A(n565), .ZN(n559) );
  NAND2_X1 U524 ( .A1(n565), .A2(n384), .ZN(n383) );
  INV_X1 U525 ( .A(n365), .ZN(n384) );
  NAND2_X1 U526 ( .A1(n559), .A2(n365), .ZN(n386) );
  NAND2_X1 U527 ( .A1(n723), .A2(n365), .ZN(n388) );
  NAND2_X1 U528 ( .A1(n390), .A2(KEYINPUT89), .ZN(n424) );
  XNOR2_X1 U529 ( .A(n420), .B(n391), .ZN(n768) );
  NAND2_X1 U530 ( .A1(n621), .A2(n398), .ZN(n396) );
  NAND2_X1 U531 ( .A1(n400), .A2(n392), .ZN(n399) );
  NAND2_X1 U532 ( .A1(n395), .A2(n393), .ZN(n593) );
  NAND2_X1 U533 ( .A1(n394), .A2(n400), .ZN(n393) );
  NAND2_X1 U534 ( .A1(n591), .A2(n398), .ZN(n397) );
  XNOR2_X1 U535 ( .A(n399), .B(G143), .ZN(G45) );
  NOR2_X1 U536 ( .A1(n546), .A2(n545), .ZN(n410) );
  XNOR2_X1 U537 ( .A(n625), .B(KEYINPUT46), .ZN(n403) );
  XNOR2_X1 U538 ( .A(n429), .B(n439), .ZN(n404) );
  INV_X1 U539 ( .A(n546), .ZN(n438) );
  NOR2_X2 U540 ( .A1(n775), .A2(n651), .ZN(n556) );
  XNOR2_X1 U541 ( .A(n410), .B(KEYINPUT64), .ZN(n409) );
  XNOR2_X1 U542 ( .A(n412), .B(KEYINPUT73), .ZN(n616) );
  NAND2_X1 U543 ( .A1(n415), .A2(n413), .ZN(n412) );
  NAND2_X1 U544 ( .A1(n414), .A2(n355), .ZN(n413) );
  XNOR2_X1 U545 ( .A(n608), .B(KEYINPUT74), .ZN(n414) );
  XNOR2_X1 U546 ( .A(n416), .B(n606), .ZN(n415) );
  NAND2_X1 U547 ( .A1(n604), .A2(n605), .ZN(n416) );
  NAND2_X1 U548 ( .A1(n421), .A2(n417), .ZN(n425) );
  NAND2_X1 U549 ( .A1(n425), .A2(n636), .ZN(n685) );
  XNOR2_X1 U550 ( .A(n469), .B(KEYINPUT0), .ZN(n549) );
  NAND2_X1 U551 ( .A1(n616), .A2(n615), .ZN(n429) );
  NAND2_X1 U552 ( .A1(n433), .A2(n774), .ZN(n580) );
  NAND2_X1 U553 ( .A1(n434), .A2(KEYINPUT90), .ZN(n433) );
  NAND2_X1 U554 ( .A1(n435), .A2(n548), .ZN(n434) );
  XNOR2_X1 U555 ( .A(n556), .B(n436), .ZN(n435) );
  INV_X1 U556 ( .A(KEYINPUT91), .ZN(n436) );
  XNOR2_X2 U557 ( .A(n502), .B(KEYINPUT22), .ZN(n546) );
  INV_X1 U558 ( .A(KEYINPUT70), .ZN(n439) );
  INV_X1 U559 ( .A(KEYINPUT84), .ZN(n606) );
  INV_X1 U560 ( .A(KEYINPUT11), .ZN(n480) );
  XNOR2_X1 U561 ( .A(n481), .B(n480), .ZN(n482) );
  XNOR2_X1 U562 ( .A(n483), .B(n482), .ZN(n485) );
  INV_X1 U563 ( .A(KEYINPUT34), .ZN(n553) );
  INV_X1 U564 ( .A(KEYINPUT56), .ZN(n645) );
  XNOR2_X1 U565 ( .A(n444), .B(n443), .ZN(n446) );
  XNOR2_X1 U566 ( .A(KEYINPUT67), .B(KEYINPUT4), .ZN(n503) );
  XNOR2_X1 U567 ( .A(n446), .B(n445), .ZN(n452) );
  XNOR2_X2 U568 ( .A(G143), .B(KEYINPUT82), .ZN(n448) );
  XNOR2_X2 U569 ( .A(n448), .B(n447), .ZN(n496) );
  NAND2_X1 U570 ( .A1(G224), .A2(n767), .ZN(n449) );
  XNOR2_X1 U571 ( .A(n506), .B(n449), .ZN(n450) );
  XNOR2_X1 U572 ( .A(n496), .B(n450), .ZN(n451) );
  XNOR2_X1 U573 ( .A(n452), .B(n451), .ZN(n459) );
  XOR2_X1 U574 ( .A(G122), .B(KEYINPUT16), .Z(n458) );
  XNOR2_X1 U575 ( .A(G119), .B(G116), .ZN(n454) );
  XNOR2_X1 U576 ( .A(G110), .B(G107), .ZN(n456) );
  XNOR2_X1 U577 ( .A(n456), .B(G104), .ZN(n520) );
  XNOR2_X1 U578 ( .A(n513), .B(n520), .ZN(n457) );
  NAND2_X1 U579 ( .A1(n535), .A2(n460), .ZN(n463) );
  NAND2_X1 U580 ( .A1(n463), .A2(G210), .ZN(n461) );
  XNOR2_X1 U581 ( .A(n461), .B(KEYINPUT94), .ZN(n462) );
  NAND2_X1 U582 ( .A1(n463), .A2(G214), .ZN(n708) );
  XNOR2_X1 U583 ( .A(n464), .B(KEYINPUT14), .ZN(n465) );
  NAND2_X1 U584 ( .A1(n465), .A2(G952), .ZN(n720) );
  XNOR2_X1 U585 ( .A(KEYINPUT95), .B(n359), .ZN(n585) );
  NAND2_X1 U586 ( .A1(G902), .A2(n465), .ZN(n466) );
  XOR2_X1 U587 ( .A(n466), .B(KEYINPUT97), .Z(n583) );
  XOR2_X1 U588 ( .A(G898), .B(KEYINPUT96), .Z(n755) );
  NAND2_X1 U589 ( .A1(G953), .A2(n755), .ZN(n761) );
  NOR2_X1 U590 ( .A1(n583), .A2(n761), .ZN(n467) );
  NOR2_X1 U591 ( .A1(n585), .A2(n467), .ZN(n468) );
  NAND2_X1 U592 ( .A1(n635), .A2(G234), .ZN(n471) );
  INV_X1 U593 ( .A(KEYINPUT20), .ZN(n470) );
  XNOR2_X1 U594 ( .A(n471), .B(n470), .ZN(n536) );
  INV_X1 U595 ( .A(G221), .ZN(n472) );
  OR2_X1 U596 ( .A1(n536), .A2(n472), .ZN(n475) );
  INV_X1 U597 ( .A(KEYINPUT100), .ZN(n473) );
  XNOR2_X1 U598 ( .A(n473), .B(KEYINPUT21), .ZN(n474) );
  XNOR2_X1 U599 ( .A(n475), .B(n474), .ZN(n692) );
  XNOR2_X1 U600 ( .A(G140), .B(G131), .ZN(n518) );
  XNOR2_X1 U601 ( .A(n477), .B(n476), .ZN(n525) );
  XOR2_X1 U602 ( .A(n518), .B(n525), .Z(n766) );
  XOR2_X1 U603 ( .A(KEYINPUT12), .B(KEYINPUT103), .Z(n479) );
  XNOR2_X1 U604 ( .A(G104), .B(G122), .ZN(n478) );
  XNOR2_X1 U605 ( .A(n479), .B(n478), .ZN(n483) );
  XNOR2_X1 U606 ( .A(G113), .B(G143), .ZN(n481) );
  NAND2_X1 U607 ( .A1(n508), .A2(G214), .ZN(n484) );
  XNOR2_X1 U608 ( .A(n485), .B(n484), .ZN(n486) );
  XNOR2_X1 U609 ( .A(n766), .B(n486), .ZN(n669) );
  NOR2_X1 U610 ( .A1(G902), .A2(n669), .ZN(n489) );
  XNOR2_X1 U611 ( .A(KEYINPUT13), .B(KEYINPUT104), .ZN(n487) );
  INV_X1 U612 ( .A(G475), .ZN(n667) );
  XOR2_X1 U613 ( .A(G122), .B(KEYINPUT9), .Z(n493) );
  NAND2_X1 U614 ( .A1(G234), .A2(n767), .ZN(n490) );
  XNOR2_X1 U615 ( .A(n491), .B(n490), .ZN(n524) );
  NAND2_X1 U616 ( .A1(G217), .A2(n524), .ZN(n492) );
  XNOR2_X2 U617 ( .A(n496), .B(n495), .ZN(n505) );
  XNOR2_X1 U618 ( .A(n505), .B(n497), .ZN(n498) );
  NAND2_X1 U619 ( .A1(n663), .A2(n535), .ZN(n499) );
  INV_X1 U620 ( .A(G478), .ZN(n662) );
  NAND2_X1 U621 ( .A1(n570), .A2(n567), .ZN(n710) );
  INV_X1 U622 ( .A(n710), .ZN(n500) );
  AND2_X1 U623 ( .A1(n692), .A2(n500), .ZN(n501) );
  NAND2_X1 U624 ( .A1(n549), .A2(n501), .ZN(n502) );
  XNOR2_X1 U625 ( .A(n503), .B(G137), .ZN(n504) );
  XNOR2_X1 U626 ( .A(n506), .B(G146), .ZN(n507) );
  NAND2_X1 U627 ( .A1(n508), .A2(G210), .ZN(n509) );
  XNOR2_X1 U628 ( .A(n509), .B(KEYINPUT5), .ZN(n512) );
  INV_X1 U629 ( .A(KEYINPUT75), .ZN(n510) );
  XNOR2_X1 U630 ( .A(n510), .B(G131), .ZN(n511) );
  XNOR2_X1 U631 ( .A(n512), .B(n511), .ZN(n514) );
  INV_X1 U632 ( .A(G472), .ZN(n652) );
  NAND2_X1 U633 ( .A1(n767), .A2(G227), .ZN(n517) );
  XNOR2_X1 U634 ( .A(n518), .B(n517), .ZN(n519) );
  XNOR2_X1 U635 ( .A(n520), .B(n519), .ZN(n521) );
  XNOR2_X1 U636 ( .A(n522), .B(n521), .ZN(n678) );
  INV_X1 U637 ( .A(KEYINPUT71), .ZN(n523) );
  XNOR2_X2 U638 ( .A(n598), .B(KEYINPUT1), .ZN(n550) );
  NAND2_X1 U639 ( .A1(n524), .A2(G221), .ZN(n526) );
  XNOR2_X1 U640 ( .A(n526), .B(n525), .ZN(n534) );
  XNOR2_X1 U641 ( .A(G128), .B(G137), .ZN(n528) );
  XNOR2_X1 U642 ( .A(G110), .B(G140), .ZN(n527) );
  XNOR2_X1 U643 ( .A(n528), .B(n527), .ZN(n532) );
  XNOR2_X1 U644 ( .A(G119), .B(KEYINPUT24), .ZN(n530) );
  XNOR2_X1 U645 ( .A(n530), .B(n529), .ZN(n531) );
  XNOR2_X1 U646 ( .A(n532), .B(n531), .ZN(n533) );
  XNOR2_X1 U647 ( .A(n534), .B(n533), .ZN(n660) );
  NAND2_X1 U648 ( .A1(n660), .A2(n535), .ZN(n543) );
  INV_X1 U649 ( .A(n536), .ZN(n537) );
  AND2_X1 U650 ( .A1(n537), .A2(G217), .ZN(n541) );
  XNOR2_X1 U651 ( .A(KEYINPUT77), .B(KEYINPUT99), .ZN(n539) );
  XNOR2_X1 U652 ( .A(KEYINPUT25), .B(KEYINPUT76), .ZN(n538) );
  XNOR2_X1 U653 ( .A(n539), .B(n538), .ZN(n540) );
  XNOR2_X1 U654 ( .A(n541), .B(n540), .ZN(n542) );
  XNOR2_X1 U655 ( .A(n543), .B(n542), .ZN(n693) );
  INV_X1 U656 ( .A(n693), .ZN(n547) );
  NAND2_X1 U657 ( .A1(n550), .A2(n547), .ZN(n544) );
  INV_X1 U658 ( .A(n697), .ZN(n562) );
  OR2_X1 U659 ( .A1(n550), .A2(n562), .ZN(n545) );
  INV_X1 U660 ( .A(KEYINPUT44), .ZN(n548) );
  XNOR2_X1 U661 ( .A(KEYINPUT33), .B(KEYINPUT72), .ZN(n551) );
  INV_X1 U662 ( .A(KEYINPUT90), .ZN(n555) );
  NAND2_X1 U663 ( .A1(n557), .A2(n556), .ZN(n558) );
  NAND2_X1 U664 ( .A1(n558), .A2(KEYINPUT44), .ZN(n578) );
  NOR2_X1 U665 ( .A1(n559), .A2(n562), .ZN(n561) );
  NAND2_X1 U666 ( .A1(n598), .A2(n687), .ZN(n560) );
  NAND2_X1 U667 ( .A1(n561), .A2(n590), .ZN(n736) );
  INV_X1 U668 ( .A(n550), .ZN(n689) );
  NAND2_X1 U669 ( .A1(n562), .A2(n687), .ZN(n563) );
  NOR2_X1 U670 ( .A1(n689), .A2(n563), .ZN(n564) );
  XNOR2_X1 U671 ( .A(n564), .B(KEYINPUT102), .ZN(n701) );
  AND2_X1 U672 ( .A1(n565), .A2(n701), .ZN(n566) );
  XNOR2_X1 U673 ( .A(n566), .B(KEYINPUT31), .ZN(n746) );
  NAND2_X1 U674 ( .A1(n736), .A2(n746), .ZN(n572) );
  INV_X1 U675 ( .A(n744), .ZN(n741) );
  INV_X1 U676 ( .A(n607), .ZN(n571) );
  NAND2_X1 U677 ( .A1(n572), .A2(n571), .ZN(n577) );
  NAND2_X1 U678 ( .A1(n689), .A2(n693), .ZN(n573) );
  NOR2_X1 U679 ( .A1(n574), .A2(n573), .ZN(n733) );
  NOR2_X1 U680 ( .A1(KEYINPUT44), .A2(KEYINPUT90), .ZN(n575) );
  NOR2_X1 U681 ( .A1(n733), .A2(n575), .ZN(n576) );
  INV_X1 U682 ( .A(KEYINPUT45), .ZN(n581) );
  XNOR2_X2 U683 ( .A(n582), .B(n581), .ZN(n756) );
  OR2_X1 U684 ( .A1(n767), .A2(n583), .ZN(n584) );
  INV_X1 U685 ( .A(n585), .ZN(n586) );
  NAND2_X1 U686 ( .A1(n361), .A2(n586), .ZN(n594) );
  NAND2_X1 U687 ( .A1(n712), .A2(KEYINPUT47), .ZN(n592) );
  NAND2_X1 U688 ( .A1(n594), .A2(n692), .ZN(n595) );
  OR2_X1 U689 ( .A1(n693), .A2(n595), .ZN(n609) );
  XNOR2_X1 U690 ( .A(n597), .B(n364), .ZN(n599) );
  NAND2_X1 U691 ( .A1(n599), .A2(n598), .ZN(n600) );
  INV_X1 U692 ( .A(n601), .ZN(n602) );
  INV_X1 U693 ( .A(KEYINPUT85), .ZN(n603) );
  INV_X1 U694 ( .A(n609), .ZN(n611) );
  XNOR2_X1 U695 ( .A(KEYINPUT107), .B(n612), .ZN(n613) );
  INV_X1 U696 ( .A(n749), .ZN(n615) );
  NAND2_X1 U697 ( .A1(n708), .A2(n707), .ZN(n711) );
  XNOR2_X1 U698 ( .A(KEYINPUT111), .B(KEYINPUT42), .ZN(n618) );
  XNOR2_X1 U699 ( .A(n619), .B(n618), .ZN(n776) );
  NAND2_X1 U700 ( .A1(n707), .A2(n590), .ZN(n620) );
  NAND2_X1 U701 ( .A1(n627), .A2(n741), .ZN(n624) );
  INV_X1 U702 ( .A(KEYINPUT40), .ZN(n623) );
  XNOR2_X1 U703 ( .A(KEYINPUT69), .B(KEYINPUT48), .ZN(n626) );
  NAND2_X1 U704 ( .A1(n627), .A2(n735), .ZN(n649) );
  OR2_X1 U705 ( .A1(n550), .A2(n628), .ZN(n630) );
  XNOR2_X1 U706 ( .A(KEYINPUT108), .B(KEYINPUT43), .ZN(n629) );
  XNOR2_X1 U707 ( .A(n630), .B(n629), .ZN(n631) );
  INV_X1 U708 ( .A(n752), .ZN(n632) );
  AND2_X1 U709 ( .A1(n649), .A2(n632), .ZN(n633) );
  NOR2_X1 U710 ( .A1(n634), .A2(KEYINPUT2), .ZN(n684) );
  NOR2_X1 U711 ( .A1(n684), .A2(n635), .ZN(n637) );
  INV_X1 U712 ( .A(n756), .ZN(n636) );
  NAND2_X2 U713 ( .A1(n637), .A2(n685), .ZN(n668) );
  NAND2_X1 U714 ( .A1(n675), .A2(G210), .ZN(n641) );
  XOR2_X1 U715 ( .A(KEYINPUT54), .B(KEYINPUT55), .Z(n639) );
  XNOR2_X1 U716 ( .A(n641), .B(n640), .ZN(n644) );
  INV_X1 U717 ( .A(G952), .ZN(n642) );
  NAND2_X1 U718 ( .A1(n642), .A2(G953), .ZN(n643) );
  NAND2_X1 U719 ( .A1(n644), .A2(n681), .ZN(n646) );
  XNOR2_X1 U720 ( .A(n646), .B(n645), .ZN(G51) );
  NAND2_X1 U721 ( .A1(n355), .A2(n735), .ZN(n648) );
  XOR2_X1 U722 ( .A(G128), .B(KEYINPUT29), .Z(n647) );
  XNOR2_X1 U723 ( .A(n648), .B(n647), .ZN(G30) );
  XNOR2_X1 U724 ( .A(n649), .B(G134), .ZN(G36) );
  XOR2_X1 U725 ( .A(G131), .B(n650), .Z(G33) );
  XOR2_X1 U726 ( .A(n651), .B(G110), .Z(G12) );
  NOR2_X1 U727 ( .A1(n668), .A2(n652), .ZN(n656) );
  XNOR2_X1 U728 ( .A(KEYINPUT112), .B(KEYINPUT62), .ZN(n653) );
  XNOR2_X1 U729 ( .A(n654), .B(n653), .ZN(n655) );
  XNOR2_X1 U730 ( .A(n656), .B(n655), .ZN(n657) );
  NAND2_X1 U731 ( .A1(n657), .A2(n681), .ZN(n658) );
  XNOR2_X1 U732 ( .A(n658), .B(KEYINPUT63), .ZN(G57) );
  NAND2_X1 U733 ( .A1(n675), .A2(G217), .ZN(n659) );
  XOR2_X1 U734 ( .A(n660), .B(n659), .Z(n661) );
  INV_X1 U735 ( .A(n681), .ZN(n665) );
  NOR2_X1 U736 ( .A1(n661), .A2(n665), .ZN(G66) );
  NOR2_X1 U737 ( .A1(n668), .A2(n662), .ZN(n664) );
  XNOR2_X1 U738 ( .A(n663), .B(n664), .ZN(n666) );
  NOR2_X1 U739 ( .A1(n666), .A2(n665), .ZN(G63) );
  NOR2_X1 U740 ( .A1(n668), .A2(n667), .ZN(n671) );
  XOR2_X1 U741 ( .A(KEYINPUT59), .B(n669), .Z(n670) );
  XNOR2_X1 U742 ( .A(n671), .B(n670), .ZN(n672) );
  NAND2_X1 U743 ( .A1(n672), .A2(n681), .ZN(n674) );
  XOR2_X1 U744 ( .A(KEYINPUT126), .B(KEYINPUT60), .Z(n673) );
  XNOR2_X1 U745 ( .A(n674), .B(n673), .ZN(G60) );
  NAND2_X1 U746 ( .A1(n675), .A2(G469), .ZN(n680) );
  XNOR2_X1 U747 ( .A(KEYINPUT124), .B(KEYINPUT57), .ZN(n676) );
  XNOR2_X1 U748 ( .A(n676), .B(KEYINPUT58), .ZN(n677) );
  XNOR2_X1 U749 ( .A(n678), .B(n677), .ZN(n679) );
  XNOR2_X1 U750 ( .A(n680), .B(n679), .ZN(n682) );
  NAND2_X1 U751 ( .A1(n682), .A2(n681), .ZN(n683) );
  XNOR2_X1 U752 ( .A(n683), .B(KEYINPUT125), .ZN(G54) );
  XNOR2_X1 U753 ( .A(n684), .B(KEYINPUT83), .ZN(n686) );
  NAND2_X1 U754 ( .A1(n686), .A2(n685), .ZN(n728) );
  XOR2_X1 U755 ( .A(KEYINPUT118), .B(KEYINPUT50), .Z(n691) );
  INV_X1 U756 ( .A(n687), .ZN(n688) );
  NAND2_X1 U757 ( .A1(n689), .A2(n688), .ZN(n690) );
  XNOR2_X1 U758 ( .A(n691), .B(n690), .ZN(n700) );
  NOR2_X1 U759 ( .A1(n693), .A2(n692), .ZN(n695) );
  XNOR2_X1 U760 ( .A(KEYINPUT116), .B(KEYINPUT49), .ZN(n694) );
  XNOR2_X1 U761 ( .A(n695), .B(n694), .ZN(n696) );
  NAND2_X1 U762 ( .A1(n697), .A2(n696), .ZN(n698) );
  XOR2_X1 U763 ( .A(KEYINPUT117), .B(n698), .Z(n699) );
  NOR2_X1 U764 ( .A1(n700), .A2(n699), .ZN(n702) );
  NOR2_X1 U765 ( .A1(n702), .A2(n701), .ZN(n703) );
  XNOR2_X1 U766 ( .A(KEYINPUT51), .B(n703), .ZN(n705) );
  NAND2_X1 U767 ( .A1(n705), .A2(n704), .ZN(n706) );
  XNOR2_X1 U768 ( .A(n706), .B(KEYINPUT119), .ZN(n718) );
  NOR2_X1 U769 ( .A1(n708), .A2(n707), .ZN(n709) );
  NOR2_X1 U770 ( .A1(n710), .A2(n709), .ZN(n715) );
  NOR2_X1 U771 ( .A1(n712), .A2(n711), .ZN(n713) );
  XNOR2_X1 U772 ( .A(n713), .B(KEYINPUT120), .ZN(n714) );
  NOR2_X1 U773 ( .A1(n715), .A2(n714), .ZN(n716) );
  NOR2_X1 U774 ( .A1(n723), .A2(n716), .ZN(n717) );
  NOR2_X1 U775 ( .A1(n718), .A2(n717), .ZN(n719) );
  XNOR2_X1 U776 ( .A(n719), .B(KEYINPUT52), .ZN(n721) );
  NOR2_X1 U777 ( .A1(n721), .A2(n720), .ZN(n726) );
  NOR2_X1 U778 ( .A1(n723), .A2(n722), .ZN(n724) );
  XOR2_X1 U779 ( .A(n724), .B(KEYINPUT121), .Z(n725) );
  NOR2_X1 U780 ( .A1(n726), .A2(n725), .ZN(n727) );
  NAND2_X1 U781 ( .A1(n728), .A2(n727), .ZN(n729) );
  XNOR2_X1 U782 ( .A(n729), .B(KEYINPUT122), .ZN(n730) );
  NOR2_X1 U783 ( .A1(n730), .A2(G953), .ZN(n732) );
  XOR2_X1 U784 ( .A(KEYINPUT123), .B(KEYINPUT53), .Z(n731) );
  XNOR2_X1 U785 ( .A(n732), .B(n731), .ZN(G75) );
  XOR2_X1 U786 ( .A(G101), .B(n733), .Z(G3) );
  NOR2_X1 U787 ( .A1(n744), .A2(n736), .ZN(n734) );
  XOR2_X1 U788 ( .A(G104), .B(n734), .Z(G6) );
  INV_X1 U789 ( .A(n735), .ZN(n747) );
  NOR2_X1 U790 ( .A1(n736), .A2(n747), .ZN(n740) );
  XOR2_X1 U791 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n738) );
  XNOR2_X1 U792 ( .A(G107), .B(KEYINPUT113), .ZN(n737) );
  XNOR2_X1 U793 ( .A(n738), .B(n737), .ZN(n739) );
  XNOR2_X1 U794 ( .A(n740), .B(n739), .ZN(G9) );
  NAND2_X1 U795 ( .A1(n355), .A2(n741), .ZN(n742) );
  XNOR2_X1 U796 ( .A(n742), .B(KEYINPUT114), .ZN(n743) );
  XNOR2_X1 U797 ( .A(G146), .B(n743), .ZN(G48) );
  NOR2_X1 U798 ( .A1(n744), .A2(n746), .ZN(n745) );
  XOR2_X1 U799 ( .A(G113), .B(n745), .Z(G15) );
  NOR2_X1 U800 ( .A1(n747), .A2(n746), .ZN(n748) );
  XOR2_X1 U801 ( .A(G116), .B(n748), .Z(G18) );
  XOR2_X1 U802 ( .A(KEYINPUT115), .B(KEYINPUT37), .Z(n751) );
  XNOR2_X1 U803 ( .A(n749), .B(G125), .ZN(n750) );
  XNOR2_X1 U804 ( .A(n751), .B(n750), .ZN(G27) );
  XOR2_X1 U805 ( .A(G140), .B(n752), .Z(G42) );
  NAND2_X1 U806 ( .A1(G953), .A2(G224), .ZN(n753) );
  XOR2_X1 U807 ( .A(KEYINPUT61), .B(n753), .Z(n754) );
  NOR2_X1 U808 ( .A1(n755), .A2(n754), .ZN(n758) );
  NOR2_X1 U809 ( .A1(G953), .A2(n756), .ZN(n757) );
  NOR2_X1 U810 ( .A1(n758), .A2(n757), .ZN(n764) );
  XNOR2_X1 U811 ( .A(n759), .B(G101), .ZN(n760) );
  XNOR2_X1 U812 ( .A(n760), .B(KEYINPUT127), .ZN(n762) );
  NAND2_X1 U813 ( .A1(n762), .A2(n761), .ZN(n763) );
  XNOR2_X1 U814 ( .A(n764), .B(n763), .ZN(G69) );
  XNOR2_X1 U815 ( .A(n765), .B(n766), .ZN(n769) );
  NAND2_X1 U816 ( .A1(n768), .A2(n767), .ZN(n773) );
  XNOR2_X1 U817 ( .A(n769), .B(G227), .ZN(n770) );
  NAND2_X1 U818 ( .A1(n770), .A2(G900), .ZN(n771) );
  NAND2_X1 U819 ( .A1(n771), .A2(G953), .ZN(n772) );
  NAND2_X1 U820 ( .A1(n773), .A2(n772), .ZN(G72) );
  XNOR2_X1 U821 ( .A(G122), .B(n774), .ZN(G24) );
  XOR2_X1 U822 ( .A(n775), .B(G119), .Z(G21) );
  XOR2_X1 U823 ( .A(G137), .B(n776), .Z(G39) );
endmodule

