//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 0 1 0 1 1 1 1 1 1 1 1 1 0 1 1 1 1 0 0 0 1 1 0 0 1 1 1 0 0 0 0 1 0 1 0 0 0 1 0 1 1 0 1 1 0 0 0 1 1 0 1 1 1 0 0 1 0 0 0 1 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:22:20 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n659, new_n660, new_n661, new_n662, new_n663, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n711, new_n712, new_n713, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n728, new_n730, new_n731, new_n732, new_n734, new_n735,
    new_n736, new_n737, new_n738, new_n739, new_n740, new_n741, new_n742,
    new_n743, new_n745, new_n746, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n761, new_n762, new_n763, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n790, new_n791, new_n792, new_n793, new_n794, new_n795, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n931, new_n932, new_n933, new_n934,
    new_n935, new_n936, new_n937, new_n938, new_n939, new_n940, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n952, new_n953, new_n954, new_n955, new_n956, new_n957,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n991, new_n992, new_n993, new_n994,
    new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001;
  OAI21_X1  g000(.A(G214), .B1(G237), .B2(G902), .ZN(new_n187));
  INV_X1    g001(.A(G952), .ZN(new_n188));
  AOI211_X1 g002(.A(G953), .B(new_n188), .C1(G234), .C2(G237), .ZN(new_n189));
  INV_X1    g003(.A(G953), .ZN(new_n190));
  XOR2_X1   g004(.A(KEYINPUT72), .B(G902), .Z(new_n191));
  AOI211_X1 g005(.A(new_n190), .B(new_n191), .C1(G234), .C2(G237), .ZN(new_n192));
  XNOR2_X1  g006(.A(KEYINPUT21), .B(G898), .ZN(new_n193));
  AOI21_X1  g007(.A(new_n189), .B1(new_n192), .B2(new_n193), .ZN(new_n194));
  INV_X1    g008(.A(new_n194), .ZN(new_n195));
  XNOR2_X1  g009(.A(G128), .B(G143), .ZN(new_n196));
  OR2_X1    g010(.A1(new_n196), .A2(G134), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n196), .A2(G134), .ZN(new_n198));
  INV_X1    g012(.A(G128), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n199), .A2(G143), .ZN(new_n200));
  INV_X1    g014(.A(KEYINPUT13), .ZN(new_n201));
  NAND3_X1  g015(.A1(new_n200), .A2(new_n201), .A3(G134), .ZN(new_n202));
  NAND3_X1  g016(.A1(new_n197), .A2(new_n198), .A3(new_n202), .ZN(new_n203));
  NAND4_X1  g017(.A1(new_n196), .A2(new_n201), .A3(G134), .A4(new_n200), .ZN(new_n204));
  INV_X1    g018(.A(KEYINPUT96), .ZN(new_n205));
  INV_X1    g019(.A(G116), .ZN(new_n206));
  OAI21_X1  g020(.A(new_n205), .B1(new_n206), .B2(G122), .ZN(new_n207));
  INV_X1    g021(.A(G122), .ZN(new_n208));
  NAND3_X1  g022(.A1(new_n208), .A2(KEYINPUT96), .A3(G116), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n207), .A2(new_n209), .ZN(new_n210));
  INV_X1    g024(.A(G107), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n211), .A2(KEYINPUT78), .ZN(new_n212));
  INV_X1    g026(.A(KEYINPUT78), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n213), .A2(G107), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n212), .A2(new_n214), .ZN(new_n215));
  INV_X1    g029(.A(new_n215), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n206), .A2(G122), .ZN(new_n217));
  AND3_X1   g031(.A1(new_n210), .A2(new_n216), .A3(new_n217), .ZN(new_n218));
  AOI21_X1  g032(.A(new_n216), .B1(new_n210), .B2(new_n217), .ZN(new_n219));
  OAI211_X1 g033(.A(new_n203), .B(new_n204), .C1(new_n218), .C2(new_n219), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n217), .A2(KEYINPUT14), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n210), .A2(new_n221), .ZN(new_n222));
  INV_X1    g036(.A(KEYINPUT98), .ZN(new_n223));
  OAI22_X1  g037(.A1(new_n222), .A2(new_n223), .B1(KEYINPUT14), .B2(new_n217), .ZN(new_n224));
  INV_X1    g038(.A(new_n224), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n222), .A2(new_n223), .ZN(new_n226));
  AOI21_X1  g040(.A(new_n211), .B1(new_n225), .B2(new_n226), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n218), .A2(KEYINPUT97), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n197), .A2(new_n198), .ZN(new_n229));
  INV_X1    g043(.A(new_n229), .ZN(new_n230));
  NAND3_X1  g044(.A1(new_n216), .A2(new_n210), .A3(new_n217), .ZN(new_n231));
  INV_X1    g045(.A(KEYINPUT97), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n231), .A2(new_n232), .ZN(new_n233));
  NAND3_X1  g047(.A1(new_n228), .A2(new_n230), .A3(new_n233), .ZN(new_n234));
  OAI21_X1  g048(.A(new_n220), .B1(new_n227), .B2(new_n234), .ZN(new_n235));
  XNOR2_X1  g049(.A(KEYINPUT9), .B(G234), .ZN(new_n236));
  INV_X1    g050(.A(G217), .ZN(new_n237));
  NOR3_X1   g051(.A1(new_n236), .A2(new_n237), .A3(G953), .ZN(new_n238));
  INV_X1    g052(.A(new_n238), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n235), .A2(new_n239), .ZN(new_n240));
  OAI211_X1 g054(.A(new_n238), .B(new_n220), .C1(new_n227), .C2(new_n234), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n240), .A2(new_n241), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n242), .A2(new_n191), .ZN(new_n243));
  INV_X1    g057(.A(G478), .ZN(new_n244));
  NOR2_X1   g058(.A1(new_n244), .A2(KEYINPUT15), .ZN(new_n245));
  NOR2_X1   g059(.A1(new_n243), .A2(new_n245), .ZN(new_n246));
  AOI21_X1  g060(.A(KEYINPUT99), .B1(new_n242), .B2(new_n191), .ZN(new_n247));
  INV_X1    g061(.A(KEYINPUT99), .ZN(new_n248));
  INV_X1    g062(.A(new_n191), .ZN(new_n249));
  AOI211_X1 g063(.A(new_n248), .B(new_n249), .C1(new_n240), .C2(new_n241), .ZN(new_n250));
  NOR2_X1   g064(.A1(new_n247), .A2(new_n250), .ZN(new_n251));
  AOI21_X1  g065(.A(new_n246), .B1(new_n251), .B2(new_n245), .ZN(new_n252));
  NOR2_X1   g066(.A1(G475), .A2(G902), .ZN(new_n253));
  XNOR2_X1  g067(.A(G113), .B(G122), .ZN(new_n254));
  INV_X1    g068(.A(G104), .ZN(new_n255));
  XNOR2_X1  g069(.A(new_n254), .B(new_n255), .ZN(new_n256));
  INV_X1    g070(.A(KEYINPUT16), .ZN(new_n257));
  INV_X1    g071(.A(G140), .ZN(new_n258));
  NAND3_X1  g072(.A1(new_n257), .A2(new_n258), .A3(G125), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n258), .A2(G125), .ZN(new_n260));
  INV_X1    g074(.A(G125), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n261), .A2(G140), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n260), .A2(new_n262), .ZN(new_n263));
  OAI211_X1 g077(.A(G146), .B(new_n259), .C1(new_n263), .C2(new_n257), .ZN(new_n264));
  INV_X1    g078(.A(G237), .ZN(new_n265));
  NAND3_X1  g079(.A1(new_n265), .A2(new_n190), .A3(G214), .ZN(new_n266));
  INV_X1    g080(.A(G143), .ZN(new_n267));
  OR2_X1    g081(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n266), .A2(new_n267), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n270), .A2(G131), .ZN(new_n271));
  INV_X1    g085(.A(G131), .ZN(new_n272));
  NAND3_X1  g086(.A1(new_n268), .A2(new_n272), .A3(new_n269), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n271), .A2(new_n273), .ZN(new_n274));
  AND2_X1   g088(.A1(new_n260), .A2(new_n262), .ZN(new_n275));
  XOR2_X1   g089(.A(KEYINPUT91), .B(KEYINPUT19), .Z(new_n276));
  NAND2_X1  g090(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n263), .A2(KEYINPUT19), .ZN(new_n278));
  NAND3_X1  g092(.A1(new_n277), .A2(KEYINPUT92), .A3(new_n278), .ZN(new_n279));
  OAI21_X1  g093(.A(new_n279), .B1(KEYINPUT92), .B2(new_n277), .ZN(new_n280));
  INV_X1    g094(.A(G146), .ZN(new_n281));
  AND3_X1   g095(.A1(new_n280), .A2(KEYINPUT93), .A3(new_n281), .ZN(new_n282));
  AOI21_X1  g096(.A(KEYINPUT93), .B1(new_n280), .B2(new_n281), .ZN(new_n283));
  OAI211_X1 g097(.A(new_n264), .B(new_n274), .C1(new_n282), .C2(new_n283), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n275), .A2(new_n281), .ZN(new_n285));
  XNOR2_X1  g099(.A(new_n285), .B(KEYINPUT77), .ZN(new_n286));
  OAI21_X1  g100(.A(new_n286), .B1(new_n281), .B2(new_n275), .ZN(new_n287));
  NAND2_X1  g101(.A1(KEYINPUT18), .A2(G131), .ZN(new_n288));
  NAND3_X1  g102(.A1(new_n268), .A2(new_n269), .A3(new_n288), .ZN(new_n289));
  NAND3_X1  g103(.A1(new_n270), .A2(KEYINPUT18), .A3(G131), .ZN(new_n290));
  NAND3_X1  g104(.A1(new_n287), .A2(new_n289), .A3(new_n290), .ZN(new_n291));
  AOI21_X1  g105(.A(new_n256), .B1(new_n284), .B2(new_n291), .ZN(new_n292));
  OAI21_X1  g106(.A(KEYINPUT94), .B1(new_n274), .B2(KEYINPUT17), .ZN(new_n293));
  OAI21_X1  g107(.A(new_n259), .B1(new_n263), .B2(new_n257), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n294), .A2(new_n281), .ZN(new_n295));
  NAND3_X1  g109(.A1(new_n295), .A2(KEYINPUT74), .A3(new_n264), .ZN(new_n296));
  INV_X1    g110(.A(KEYINPUT74), .ZN(new_n297));
  NAND3_X1  g111(.A1(new_n294), .A2(new_n297), .A3(new_n281), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n296), .A2(new_n298), .ZN(new_n299));
  NAND3_X1  g113(.A1(new_n270), .A2(KEYINPUT17), .A3(G131), .ZN(new_n300));
  INV_X1    g114(.A(KEYINPUT94), .ZN(new_n301));
  INV_X1    g115(.A(KEYINPUT17), .ZN(new_n302));
  NAND4_X1  g116(.A1(new_n271), .A2(new_n301), .A3(new_n302), .A4(new_n273), .ZN(new_n303));
  NAND4_X1  g117(.A1(new_n293), .A2(new_n299), .A3(new_n300), .A4(new_n303), .ZN(new_n304));
  NAND3_X1  g118(.A1(new_n304), .A2(new_n256), .A3(new_n291), .ZN(new_n305));
  INV_X1    g119(.A(new_n305), .ZN(new_n306));
  OAI21_X1  g120(.A(new_n253), .B1(new_n292), .B2(new_n306), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n307), .A2(KEYINPUT20), .ZN(new_n308));
  INV_X1    g122(.A(KEYINPUT20), .ZN(new_n309));
  OAI211_X1 g123(.A(new_n309), .B(new_n253), .C1(new_n292), .C2(new_n306), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n308), .A2(new_n310), .ZN(new_n311));
  INV_X1    g125(.A(G902), .ZN(new_n312));
  AOI21_X1  g126(.A(new_n256), .B1(new_n304), .B2(new_n291), .ZN(new_n313));
  OAI21_X1  g127(.A(new_n312), .B1(new_n306), .B2(new_n313), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n314), .A2(KEYINPUT95), .ZN(new_n315));
  INV_X1    g129(.A(KEYINPUT95), .ZN(new_n316));
  OAI211_X1 g130(.A(new_n316), .B(new_n312), .C1(new_n306), .C2(new_n313), .ZN(new_n317));
  NAND3_X1  g131(.A1(new_n315), .A2(G475), .A3(new_n317), .ZN(new_n318));
  AND4_X1   g132(.A1(new_n195), .A2(new_n252), .A3(new_n311), .A4(new_n318), .ZN(new_n319));
  XNOR2_X1  g133(.A(G116), .B(G119), .ZN(new_n320));
  INV_X1    g134(.A(new_n320), .ZN(new_n321));
  XNOR2_X1  g135(.A(KEYINPUT2), .B(G113), .ZN(new_n322));
  NOR2_X1   g136(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  INV_X1    g137(.A(new_n323), .ZN(new_n324));
  XNOR2_X1  g138(.A(new_n320), .B(KEYINPUT68), .ZN(new_n325));
  INV_X1    g139(.A(KEYINPUT5), .ZN(new_n326));
  NOR2_X1   g140(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  INV_X1    g141(.A(G119), .ZN(new_n328));
  NAND3_X1  g142(.A1(new_n326), .A2(new_n328), .A3(G116), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n329), .A2(G113), .ZN(new_n330));
  OAI21_X1  g144(.A(new_n324), .B1(new_n327), .B2(new_n330), .ZN(new_n331));
  NOR2_X1   g145(.A1(new_n255), .A2(KEYINPUT3), .ZN(new_n332));
  INV_X1    g146(.A(KEYINPUT79), .ZN(new_n333));
  NAND4_X1  g147(.A1(new_n332), .A2(new_n212), .A3(new_n214), .A4(new_n333), .ZN(new_n334));
  AND3_X1   g148(.A1(new_n332), .A2(new_n212), .A3(new_n214), .ZN(new_n335));
  NOR2_X1   g149(.A1(new_n255), .A2(G107), .ZN(new_n336));
  INV_X1    g150(.A(KEYINPUT3), .ZN(new_n337));
  OAI21_X1  g151(.A(KEYINPUT79), .B1(new_n336), .B2(new_n337), .ZN(new_n338));
  OAI21_X1  g152(.A(new_n334), .B1(new_n335), .B2(new_n338), .ZN(new_n339));
  XOR2_X1   g153(.A(KEYINPUT81), .B(G101), .Z(new_n340));
  NOR2_X1   g154(.A1(new_n211), .A2(G104), .ZN(new_n341));
  INV_X1    g155(.A(new_n341), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n340), .A2(new_n342), .ZN(new_n343));
  INV_X1    g157(.A(new_n343), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n339), .A2(new_n344), .ZN(new_n345));
  INV_X1    g159(.A(G101), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n215), .A2(new_n255), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n211), .A2(G104), .ZN(new_n348));
  AOI21_X1  g162(.A(new_n346), .B1(new_n347), .B2(new_n348), .ZN(new_n349));
  INV_X1    g163(.A(new_n349), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n345), .A2(new_n350), .ZN(new_n351));
  OR2_X1    g165(.A1(new_n331), .A2(new_n351), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n345), .A2(KEYINPUT4), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n339), .A2(new_n342), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n354), .A2(KEYINPUT80), .ZN(new_n355));
  INV_X1    g169(.A(KEYINPUT80), .ZN(new_n356));
  NAND3_X1  g170(.A1(new_n339), .A2(new_n356), .A3(new_n342), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n355), .A2(new_n357), .ZN(new_n358));
  AOI21_X1  g172(.A(new_n353), .B1(new_n358), .B2(G101), .ZN(new_n359));
  NOR2_X1   g173(.A1(new_n346), .A2(KEYINPUT4), .ZN(new_n360));
  AOI21_X1  g174(.A(new_n356), .B1(new_n339), .B2(new_n342), .ZN(new_n361));
  NAND3_X1  g175(.A1(new_n332), .A2(new_n212), .A3(new_n214), .ZN(new_n362));
  AOI21_X1  g176(.A(new_n333), .B1(new_n348), .B2(KEYINPUT3), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n362), .A2(new_n363), .ZN(new_n364));
  AOI211_X1 g178(.A(KEYINPUT80), .B(new_n341), .C1(new_n364), .C2(new_n334), .ZN(new_n365));
  OAI21_X1  g179(.A(new_n360), .B1(new_n361), .B2(new_n365), .ZN(new_n366));
  AOI21_X1  g180(.A(new_n323), .B1(new_n325), .B2(new_n322), .ZN(new_n367));
  INV_X1    g181(.A(new_n367), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n366), .A2(new_n368), .ZN(new_n369));
  OAI21_X1  g183(.A(new_n352), .B1(new_n359), .B2(new_n369), .ZN(new_n370));
  XNOR2_X1  g184(.A(G110), .B(G122), .ZN(new_n371));
  INV_X1    g185(.A(new_n371), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n370), .A2(new_n372), .ZN(new_n373));
  OAI211_X1 g187(.A(new_n352), .B(new_n371), .C1(new_n359), .C2(new_n369), .ZN(new_n374));
  NAND3_X1  g188(.A1(new_n373), .A2(KEYINPUT6), .A3(new_n374), .ZN(new_n375));
  INV_X1    g189(.A(KEYINPUT6), .ZN(new_n376));
  NAND3_X1  g190(.A1(new_n370), .A2(new_n376), .A3(new_n372), .ZN(new_n377));
  INV_X1    g191(.A(KEYINPUT87), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n281), .A2(G143), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n267), .A2(G146), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n379), .A2(new_n380), .ZN(new_n381));
  NAND2_X1  g195(.A1(KEYINPUT0), .A2(G128), .ZN(new_n382));
  OR2_X1    g196(.A1(KEYINPUT0), .A2(G128), .ZN(new_n383));
  NAND3_X1  g197(.A1(new_n381), .A2(new_n382), .A3(new_n383), .ZN(new_n384));
  OAI21_X1  g198(.A(KEYINPUT64), .B1(new_n267), .B2(G146), .ZN(new_n385));
  INV_X1    g199(.A(KEYINPUT64), .ZN(new_n386));
  NAND3_X1  g200(.A1(new_n386), .A2(new_n281), .A3(G143), .ZN(new_n387));
  INV_X1    g201(.A(new_n382), .ZN(new_n388));
  NAND4_X1  g202(.A1(new_n385), .A2(new_n387), .A3(new_n388), .A4(new_n380), .ZN(new_n389));
  AND2_X1   g203(.A1(new_n384), .A2(new_n389), .ZN(new_n390));
  OAI21_X1  g204(.A(new_n378), .B1(new_n390), .B2(new_n261), .ZN(new_n391));
  OR2_X1    g205(.A1(KEYINPUT67), .A2(KEYINPUT1), .ZN(new_n392));
  NAND2_X1  g206(.A1(KEYINPUT67), .A2(KEYINPUT1), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n392), .A2(new_n393), .ZN(new_n394));
  AOI21_X1  g208(.A(new_n199), .B1(new_n394), .B2(new_n379), .ZN(new_n395));
  XNOR2_X1  g209(.A(G143), .B(G146), .ZN(new_n396));
  NAND3_X1  g210(.A1(new_n385), .A2(new_n387), .A3(new_n380), .ZN(new_n397));
  NAND3_X1  g211(.A1(new_n392), .A2(G128), .A3(new_n393), .ZN(new_n398));
  OAI22_X1  g212(.A1(new_n395), .A2(new_n396), .B1(new_n397), .B2(new_n398), .ZN(new_n399));
  MUX2_X1   g213(.A(new_n390), .B(new_n399), .S(new_n261), .Z(new_n400));
  OAI21_X1  g214(.A(new_n391), .B1(new_n400), .B2(new_n378), .ZN(new_n401));
  XNOR2_X1  g215(.A(KEYINPUT88), .B(G224), .ZN(new_n402));
  INV_X1    g216(.A(new_n402), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n403), .A2(new_n190), .ZN(new_n404));
  XNOR2_X1  g218(.A(new_n404), .B(KEYINPUT89), .ZN(new_n405));
  XNOR2_X1  g219(.A(new_n401), .B(new_n405), .ZN(new_n406));
  NAND3_X1  g220(.A1(new_n375), .A2(new_n377), .A3(new_n406), .ZN(new_n407));
  INV_X1    g221(.A(KEYINPUT7), .ZN(new_n408));
  NOR2_X1   g222(.A1(new_n405), .A2(new_n408), .ZN(new_n409));
  OR2_X1    g223(.A1(new_n400), .A2(new_n409), .ZN(new_n410));
  OAI211_X1 g224(.A(new_n391), .B(new_n409), .C1(new_n400), .C2(new_n378), .ZN(new_n411));
  AOI21_X1  g225(.A(new_n343), .B1(new_n364), .B2(new_n334), .ZN(new_n412));
  NOR2_X1   g226(.A1(new_n412), .A2(new_n349), .ZN(new_n413));
  NOR2_X1   g227(.A1(new_n321), .A2(new_n326), .ZN(new_n414));
  OAI21_X1  g228(.A(new_n324), .B1(new_n414), .B2(new_n330), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n413), .A2(new_n415), .ZN(new_n416));
  XNOR2_X1  g230(.A(new_n371), .B(KEYINPUT8), .ZN(new_n417));
  OAI211_X1 g231(.A(new_n416), .B(new_n417), .C1(new_n331), .C2(new_n413), .ZN(new_n418));
  AND3_X1   g232(.A1(new_n410), .A2(new_n411), .A3(new_n418), .ZN(new_n419));
  AOI21_X1  g233(.A(G902), .B1(new_n419), .B2(new_n374), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n407), .A2(new_n420), .ZN(new_n421));
  OAI21_X1  g235(.A(G210), .B1(G237), .B2(G902), .ZN(new_n422));
  INV_X1    g236(.A(new_n422), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n421), .A2(new_n423), .ZN(new_n424));
  NAND3_X1  g238(.A1(new_n407), .A2(new_n420), .A3(new_n422), .ZN(new_n425));
  NAND3_X1  g239(.A1(new_n424), .A2(KEYINPUT90), .A3(new_n425), .ZN(new_n426));
  AOI21_X1  g240(.A(new_n422), .B1(new_n407), .B2(new_n420), .ZN(new_n427));
  INV_X1    g241(.A(KEYINPUT90), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n427), .A2(new_n428), .ZN(new_n429));
  AND4_X1   g243(.A1(new_n187), .A2(new_n319), .A3(new_n426), .A4(new_n429), .ZN(new_n430));
  XNOR2_X1  g244(.A(G110), .B(G140), .ZN(new_n431));
  AND2_X1   g245(.A1(new_n190), .A2(G227), .ZN(new_n432));
  XNOR2_X1  g246(.A(new_n431), .B(new_n432), .ZN(new_n433));
  INV_X1    g247(.A(KEYINPUT82), .ZN(new_n434));
  OAI21_X1  g248(.A(new_n434), .B1(new_n397), .B2(new_n398), .ZN(new_n435));
  INV_X1    g249(.A(KEYINPUT83), .ZN(new_n436));
  OAI211_X1 g250(.A(new_n436), .B(KEYINPUT1), .C1(new_n267), .C2(G146), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n437), .A2(G128), .ZN(new_n438));
  AOI21_X1  g252(.A(new_n436), .B1(new_n379), .B2(KEYINPUT1), .ZN(new_n439));
  OAI21_X1  g253(.A(new_n397), .B1(new_n438), .B2(new_n439), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n435), .A2(new_n440), .ZN(new_n441));
  NOR3_X1   g255(.A1(new_n397), .A2(new_n398), .A3(new_n434), .ZN(new_n442));
  OAI211_X1 g256(.A(new_n345), .B(new_n350), .C1(new_n441), .C2(new_n442), .ZN(new_n443));
  NOR2_X1   g257(.A1(new_n397), .A2(new_n398), .ZN(new_n444));
  AND2_X1   g258(.A1(KEYINPUT67), .A2(KEYINPUT1), .ZN(new_n445));
  NOR2_X1   g259(.A1(KEYINPUT67), .A2(KEYINPUT1), .ZN(new_n446));
  OAI21_X1  g260(.A(new_n379), .B1(new_n445), .B2(new_n446), .ZN(new_n447));
  AOI21_X1  g261(.A(new_n396), .B1(new_n447), .B2(G128), .ZN(new_n448));
  NOR2_X1   g262(.A1(new_n444), .A2(new_n448), .ZN(new_n449));
  OAI21_X1  g263(.A(new_n449), .B1(new_n412), .B2(new_n349), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n443), .A2(new_n450), .ZN(new_n451));
  INV_X1    g265(.A(G134), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n452), .A2(G137), .ZN(new_n453));
  NOR2_X1   g267(.A1(new_n452), .A2(G137), .ZN(new_n454));
  INV_X1    g268(.A(KEYINPUT11), .ZN(new_n455));
  NOR2_X1   g269(.A1(new_n455), .A2(KEYINPUT65), .ZN(new_n456));
  OAI21_X1  g270(.A(new_n453), .B1(new_n454), .B2(new_n456), .ZN(new_n457));
  INV_X1    g271(.A(G137), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n458), .A2(G134), .ZN(new_n459));
  INV_X1    g273(.A(KEYINPUT65), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n460), .A2(KEYINPUT11), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n455), .A2(KEYINPUT65), .ZN(new_n462));
  AOI21_X1  g276(.A(new_n459), .B1(new_n461), .B2(new_n462), .ZN(new_n463));
  NOR3_X1   g277(.A1(new_n457), .A2(new_n463), .A3(G131), .ZN(new_n464));
  NOR2_X1   g278(.A1(new_n458), .A2(G134), .ZN(new_n465));
  AOI21_X1  g279(.A(new_n465), .B1(new_n459), .B2(new_n461), .ZN(new_n466));
  NOR2_X1   g280(.A1(new_n460), .A2(KEYINPUT11), .ZN(new_n467));
  OAI21_X1  g281(.A(new_n454), .B1(new_n456), .B2(new_n467), .ZN(new_n468));
  AOI21_X1  g282(.A(new_n272), .B1(new_n466), .B2(new_n468), .ZN(new_n469));
  NOR2_X1   g283(.A1(new_n464), .A2(new_n469), .ZN(new_n470));
  INV_X1    g284(.A(new_n470), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n451), .A2(new_n471), .ZN(new_n472));
  XNOR2_X1  g286(.A(new_n472), .B(KEYINPUT12), .ZN(new_n473));
  AOI21_X1  g287(.A(new_n346), .B1(new_n355), .B2(new_n357), .ZN(new_n474));
  OAI211_X1 g288(.A(new_n390), .B(new_n366), .C1(new_n474), .C2(new_n353), .ZN(new_n475));
  INV_X1    g289(.A(KEYINPUT84), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n399), .A2(KEYINPUT10), .ZN(new_n477));
  OAI21_X1  g291(.A(new_n476), .B1(new_n351), .B2(new_n477), .ZN(new_n478));
  INV_X1    g292(.A(KEYINPUT10), .ZN(new_n479));
  NOR2_X1   g293(.A1(new_n449), .A2(new_n479), .ZN(new_n480));
  NAND3_X1  g294(.A1(new_n480), .A2(new_n413), .A3(KEYINPUT84), .ZN(new_n481));
  AOI22_X1  g295(.A1(new_n478), .A2(new_n481), .B1(new_n479), .B2(new_n443), .ZN(new_n482));
  AND3_X1   g296(.A1(new_n475), .A2(new_n482), .A3(new_n470), .ZN(new_n483));
  OAI21_X1  g297(.A(new_n433), .B1(new_n473), .B2(new_n483), .ZN(new_n484));
  AOI21_X1  g298(.A(new_n470), .B1(new_n475), .B2(new_n482), .ZN(new_n485));
  NAND3_X1  g299(.A1(new_n475), .A2(new_n482), .A3(new_n470), .ZN(new_n486));
  INV_X1    g300(.A(new_n433), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n486), .A2(new_n487), .ZN(new_n488));
  OAI211_X1 g302(.A(new_n484), .B(G469), .C1(new_n485), .C2(new_n488), .ZN(new_n489));
  NAND2_X1  g303(.A1(G469), .A2(G902), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  OAI21_X1  g305(.A(new_n433), .B1(new_n483), .B2(new_n485), .ZN(new_n492));
  INV_X1    g306(.A(new_n488), .ZN(new_n493));
  INV_X1    g307(.A(KEYINPUT12), .ZN(new_n494));
  XNOR2_X1  g308(.A(new_n472), .B(new_n494), .ZN(new_n495));
  AOI22_X1  g309(.A1(new_n492), .A2(KEYINPUT85), .B1(new_n493), .B2(new_n495), .ZN(new_n496));
  INV_X1    g310(.A(KEYINPUT85), .ZN(new_n497));
  OAI211_X1 g311(.A(new_n497), .B(new_n433), .C1(new_n483), .C2(new_n485), .ZN(new_n498));
  AOI21_X1  g312(.A(new_n249), .B1(new_n496), .B2(new_n498), .ZN(new_n499));
  INV_X1    g313(.A(G469), .ZN(new_n500));
  AOI21_X1  g314(.A(new_n491), .B1(new_n499), .B2(new_n500), .ZN(new_n501));
  INV_X1    g315(.A(G221), .ZN(new_n502));
  INV_X1    g316(.A(new_n236), .ZN(new_n503));
  AOI21_X1  g317(.A(new_n502), .B1(new_n503), .B2(new_n312), .ZN(new_n504));
  OAI21_X1  g318(.A(KEYINPUT86), .B1(new_n501), .B2(new_n504), .ZN(new_n505));
  OAI21_X1  g319(.A(new_n390), .B1(new_n464), .B2(new_n469), .ZN(new_n506));
  NAND3_X1  g320(.A1(new_n466), .A2(new_n468), .A3(new_n272), .ZN(new_n507));
  INV_X1    g321(.A(KEYINPUT66), .ZN(new_n508));
  NAND3_X1  g322(.A1(new_n459), .A2(new_n453), .A3(new_n508), .ZN(new_n509));
  OAI211_X1 g323(.A(new_n509), .B(G131), .C1(new_n508), .C2(new_n459), .ZN(new_n510));
  OAI211_X1 g324(.A(new_n507), .B(new_n510), .C1(new_n444), .C2(new_n448), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n506), .A2(new_n511), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n512), .A2(KEYINPUT30), .ZN(new_n513));
  INV_X1    g327(.A(KEYINPUT30), .ZN(new_n514));
  NAND3_X1  g328(.A1(new_n506), .A2(new_n514), .A3(new_n511), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n513), .A2(new_n515), .ZN(new_n516));
  NAND3_X1  g330(.A1(new_n506), .A2(new_n367), .A3(new_n511), .ZN(new_n517));
  NAND3_X1  g331(.A1(new_n265), .A2(new_n190), .A3(G210), .ZN(new_n518));
  XNOR2_X1  g332(.A(new_n518), .B(KEYINPUT27), .ZN(new_n519));
  XNOR2_X1  g333(.A(KEYINPUT26), .B(G101), .ZN(new_n520));
  XNOR2_X1  g334(.A(new_n519), .B(new_n520), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n517), .A2(new_n521), .ZN(new_n522));
  AOI22_X1  g336(.A1(new_n516), .A2(new_n368), .B1(KEYINPUT69), .B2(new_n522), .ZN(new_n523));
  INV_X1    g337(.A(KEYINPUT31), .ZN(new_n524));
  INV_X1    g338(.A(KEYINPUT69), .ZN(new_n525));
  NAND3_X1  g339(.A1(new_n517), .A2(new_n525), .A3(new_n521), .ZN(new_n526));
  NAND4_X1  g340(.A1(new_n523), .A2(KEYINPUT70), .A3(new_n524), .A4(new_n526), .ZN(new_n527));
  AND3_X1   g341(.A1(new_n506), .A2(new_n514), .A3(new_n511), .ZN(new_n528));
  AOI21_X1  g342(.A(new_n514), .B1(new_n506), .B2(new_n511), .ZN(new_n529));
  OAI21_X1  g343(.A(new_n368), .B1(new_n528), .B2(new_n529), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n522), .A2(KEYINPUT69), .ZN(new_n531));
  NAND4_X1  g345(.A1(new_n530), .A2(new_n531), .A3(new_n524), .A4(new_n526), .ZN(new_n532));
  INV_X1    g346(.A(KEYINPUT70), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  NAND3_X1  g348(.A1(new_n530), .A2(new_n531), .A3(new_n526), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n535), .A2(KEYINPUT31), .ZN(new_n536));
  INV_X1    g350(.A(new_n521), .ZN(new_n537));
  INV_X1    g351(.A(KEYINPUT28), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n512), .A2(new_n368), .ZN(new_n539));
  AOI21_X1  g353(.A(new_n538), .B1(new_n539), .B2(new_n517), .ZN(new_n540));
  AND2_X1   g354(.A1(new_n517), .A2(new_n538), .ZN(new_n541));
  OAI21_X1  g355(.A(new_n537), .B1(new_n540), .B2(new_n541), .ZN(new_n542));
  NAND4_X1  g356(.A1(new_n527), .A2(new_n534), .A3(new_n536), .A4(new_n542), .ZN(new_n543));
  NOR2_X1   g357(.A1(G472), .A2(G902), .ZN(new_n544));
  AOI21_X1  g358(.A(KEYINPUT32), .B1(new_n543), .B2(new_n544), .ZN(new_n545));
  INV_X1    g359(.A(new_n545), .ZN(new_n546));
  NAND3_X1  g360(.A1(new_n543), .A2(KEYINPUT32), .A3(new_n544), .ZN(new_n547));
  NOR2_X1   g361(.A1(new_n540), .A2(new_n541), .ZN(new_n548));
  INV_X1    g362(.A(KEYINPUT71), .ZN(new_n549));
  NOR2_X1   g363(.A1(new_n549), .A2(KEYINPUT29), .ZN(new_n550));
  OAI21_X1  g364(.A(new_n521), .B1(new_n548), .B2(new_n550), .ZN(new_n551));
  AOI21_X1  g365(.A(new_n551), .B1(new_n548), .B2(new_n550), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n530), .A2(new_n517), .ZN(new_n553));
  INV_X1    g367(.A(new_n553), .ZN(new_n554));
  NAND3_X1  g368(.A1(new_n554), .A2(new_n537), .A3(new_n550), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n555), .A2(new_n191), .ZN(new_n556));
  OAI21_X1  g370(.A(G472), .B1(new_n552), .B2(new_n556), .ZN(new_n557));
  NAND3_X1  g371(.A1(new_n546), .A2(new_n547), .A3(new_n557), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n199), .A2(G119), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n328), .A2(G128), .ZN(new_n560));
  NAND4_X1  g374(.A1(new_n559), .A2(new_n560), .A3(KEYINPUT73), .A4(KEYINPUT23), .ZN(new_n561));
  OR2_X1    g375(.A1(KEYINPUT73), .A2(KEYINPUT23), .ZN(new_n562));
  NAND2_X1  g376(.A1(KEYINPUT73), .A2(KEYINPUT23), .ZN(new_n563));
  NAND4_X1  g377(.A1(new_n562), .A2(G119), .A3(new_n199), .A4(new_n563), .ZN(new_n564));
  NAND3_X1  g378(.A1(new_n561), .A2(new_n564), .A3(G110), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n559), .A2(new_n560), .ZN(new_n566));
  XNOR2_X1  g380(.A(KEYINPUT24), .B(G110), .ZN(new_n567));
  OR2_X1    g381(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  AND2_X1   g382(.A1(new_n565), .A2(new_n568), .ZN(new_n569));
  NAND3_X1  g383(.A1(new_n296), .A2(new_n298), .A3(new_n569), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n570), .A2(KEYINPUT75), .ZN(new_n571));
  INV_X1    g385(.A(KEYINPUT75), .ZN(new_n572));
  NAND4_X1  g386(.A1(new_n296), .A2(new_n569), .A3(new_n572), .A4(new_n298), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n571), .A2(new_n573), .ZN(new_n574));
  AOI21_X1  g388(.A(G110), .B1(new_n561), .B2(new_n564), .ZN(new_n575));
  OR2_X1    g389(.A1(new_n575), .A2(KEYINPUT76), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n575), .A2(KEYINPUT76), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n566), .A2(new_n567), .ZN(new_n578));
  NAND3_X1  g392(.A1(new_n576), .A2(new_n577), .A3(new_n578), .ZN(new_n579));
  NAND3_X1  g393(.A1(new_n579), .A2(new_n264), .A3(new_n286), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n574), .A2(new_n580), .ZN(new_n581));
  XNOR2_X1  g395(.A(KEYINPUT22), .B(G137), .ZN(new_n582));
  AND3_X1   g396(.A1(new_n190), .A2(G221), .A3(G234), .ZN(new_n583));
  XOR2_X1   g397(.A(new_n582), .B(new_n583), .Z(new_n584));
  INV_X1    g398(.A(new_n584), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n581), .A2(new_n585), .ZN(new_n586));
  AOI21_X1  g400(.A(new_n237), .B1(new_n191), .B2(G234), .ZN(new_n587));
  NOR2_X1   g401(.A1(new_n587), .A2(G902), .ZN(new_n588));
  NAND3_X1  g402(.A1(new_n574), .A2(new_n580), .A3(new_n584), .ZN(new_n589));
  AND3_X1   g403(.A1(new_n586), .A2(new_n588), .A3(new_n589), .ZN(new_n590));
  NAND3_X1  g404(.A1(new_n586), .A2(new_n191), .A3(new_n589), .ZN(new_n591));
  INV_X1    g405(.A(KEYINPUT25), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  NAND4_X1  g407(.A1(new_n586), .A2(KEYINPUT25), .A3(new_n191), .A4(new_n589), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  AOI21_X1  g409(.A(new_n590), .B1(new_n595), .B2(new_n587), .ZN(new_n596));
  AND2_X1   g410(.A1(new_n558), .A2(new_n596), .ZN(new_n597));
  NAND3_X1  g411(.A1(new_n495), .A2(new_n487), .A3(new_n486), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n366), .A2(new_n390), .ZN(new_n599));
  NOR2_X1   g413(.A1(new_n359), .A2(new_n599), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n443), .A2(new_n479), .ZN(new_n601));
  NOR3_X1   g415(.A1(new_n351), .A2(new_n477), .A3(new_n476), .ZN(new_n602));
  AOI21_X1  g416(.A(KEYINPUT84), .B1(new_n480), .B2(new_n413), .ZN(new_n603));
  OAI21_X1  g417(.A(new_n601), .B1(new_n602), .B2(new_n603), .ZN(new_n604));
  OAI21_X1  g418(.A(new_n471), .B1(new_n600), .B2(new_n604), .ZN(new_n605));
  AOI21_X1  g419(.A(new_n487), .B1(new_n605), .B2(new_n486), .ZN(new_n606));
  OAI21_X1  g420(.A(new_n598), .B1(new_n606), .B2(new_n497), .ZN(new_n607));
  INV_X1    g421(.A(new_n498), .ZN(new_n608));
  OAI211_X1 g422(.A(new_n500), .B(new_n191), .C1(new_n607), .C2(new_n608), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n495), .A2(new_n486), .ZN(new_n610));
  AOI22_X1  g424(.A1(new_n605), .A2(new_n493), .B1(new_n610), .B2(new_n433), .ZN(new_n611));
  OAI21_X1  g425(.A(G469), .B1(new_n611), .B2(G902), .ZN(new_n612));
  AOI21_X1  g426(.A(new_n504), .B1(new_n609), .B2(new_n612), .ZN(new_n613));
  INV_X1    g427(.A(KEYINPUT86), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  NAND4_X1  g429(.A1(new_n430), .A2(new_n505), .A3(new_n597), .A4(new_n615), .ZN(new_n616));
  XOR2_X1   g430(.A(new_n616), .B(new_n340), .Z(G3));
  NAND2_X1  g431(.A1(new_n609), .A2(new_n612), .ZN(new_n618));
  INV_X1    g432(.A(new_n504), .ZN(new_n619));
  AOI21_X1  g433(.A(new_n614), .B1(new_n618), .B2(new_n619), .ZN(new_n620));
  AOI211_X1 g434(.A(KEYINPUT86), .B(new_n504), .C1(new_n609), .C2(new_n612), .ZN(new_n621));
  NOR2_X1   g435(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n543), .A2(new_n191), .ZN(new_n623));
  AOI22_X1  g437(.A1(new_n623), .A2(G472), .B1(new_n543), .B2(new_n544), .ZN(new_n624));
  AND2_X1   g438(.A1(new_n624), .A2(new_n596), .ZN(new_n625));
  NAND2_X1  g439(.A1(new_n622), .A2(new_n625), .ZN(new_n626));
  AND3_X1   g440(.A1(new_n407), .A2(new_n420), .A3(new_n422), .ZN(new_n627));
  OAI21_X1  g441(.A(new_n187), .B1(new_n627), .B2(new_n427), .ZN(new_n628));
  INV_X1    g442(.A(KEYINPUT100), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  OAI211_X1 g444(.A(KEYINPUT100), .B(new_n187), .C1(new_n627), .C2(new_n427), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  INV_X1    g446(.A(new_n632), .ZN(new_n633));
  AND2_X1   g447(.A1(new_n231), .A2(new_n232), .ZN(new_n634));
  NOR2_X1   g448(.A1(new_n231), .A2(new_n232), .ZN(new_n635));
  NOR3_X1   g449(.A1(new_n634), .A2(new_n635), .A3(new_n229), .ZN(new_n636));
  INV_X1    g450(.A(new_n226), .ZN(new_n637));
  OAI21_X1  g451(.A(G107), .B1(new_n637), .B2(new_n224), .ZN(new_n638));
  AND2_X1   g452(.A1(new_n203), .A2(new_n204), .ZN(new_n639));
  OR2_X1    g453(.A1(new_n218), .A2(new_n219), .ZN(new_n640));
  AOI22_X1  g454(.A1(new_n636), .A2(new_n638), .B1(new_n639), .B2(new_n640), .ZN(new_n641));
  OAI21_X1  g455(.A(KEYINPUT101), .B1(new_n641), .B2(new_n238), .ZN(new_n642));
  NAND3_X1  g456(.A1(new_n242), .A2(KEYINPUT33), .A3(new_n642), .ZN(new_n643));
  INV_X1    g457(.A(KEYINPUT33), .ZN(new_n644));
  OAI211_X1 g458(.A(new_n240), .B(new_n241), .C1(KEYINPUT101), .C2(new_n644), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n643), .A2(new_n645), .ZN(new_n646));
  NOR2_X1   g460(.A1(new_n249), .A2(new_n244), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  AOI22_X1  g462(.A1(new_n648), .A2(KEYINPUT102), .B1(new_n251), .B2(new_n244), .ZN(new_n649));
  INV_X1    g463(.A(KEYINPUT102), .ZN(new_n650));
  NAND3_X1  g464(.A1(new_n646), .A2(new_n650), .A3(new_n647), .ZN(new_n651));
  AOI22_X1  g465(.A1(new_n649), .A2(new_n651), .B1(new_n318), .B2(new_n311), .ZN(new_n652));
  INV_X1    g466(.A(new_n652), .ZN(new_n653));
  NOR2_X1   g467(.A1(new_n653), .A2(new_n194), .ZN(new_n654));
  NAND2_X1  g468(.A1(new_n633), .A2(new_n654), .ZN(new_n655));
  NOR2_X1   g469(.A1(new_n626), .A2(new_n655), .ZN(new_n656));
  XNOR2_X1  g470(.A(KEYINPUT34), .B(G104), .ZN(new_n657));
  XNOR2_X1  g471(.A(new_n656), .B(new_n657), .ZN(G6));
  NAND2_X1  g472(.A1(new_n318), .A2(new_n311), .ZN(new_n659));
  NOR3_X1   g473(.A1(new_n659), .A2(new_n194), .A3(new_n252), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n633), .A2(new_n660), .ZN(new_n661));
  NOR2_X1   g475(.A1(new_n626), .A2(new_n661), .ZN(new_n662));
  XNOR2_X1  g476(.A(KEYINPUT35), .B(G107), .ZN(new_n663));
  XNOR2_X1  g477(.A(new_n662), .B(new_n663), .ZN(G9));
  INV_X1    g478(.A(new_n587), .ZN(new_n665));
  AOI21_X1  g479(.A(new_n665), .B1(new_n593), .B2(new_n594), .ZN(new_n666));
  NOR2_X1   g480(.A1(new_n585), .A2(KEYINPUT36), .ZN(new_n667));
  XNOR2_X1  g481(.A(new_n581), .B(new_n667), .ZN(new_n668));
  NAND2_X1  g482(.A1(new_n668), .A2(new_n588), .ZN(new_n669));
  INV_X1    g483(.A(new_n669), .ZN(new_n670));
  NOR2_X1   g484(.A1(new_n666), .A2(new_n670), .ZN(new_n671));
  INV_X1    g485(.A(new_n671), .ZN(new_n672));
  NAND2_X1  g486(.A1(new_n672), .A2(new_n624), .ZN(new_n673));
  INV_X1    g487(.A(new_n673), .ZN(new_n674));
  NAND3_X1  g488(.A1(new_n622), .A2(new_n430), .A3(new_n674), .ZN(new_n675));
  XOR2_X1   g489(.A(KEYINPUT37), .B(G110), .Z(new_n676));
  XNOR2_X1  g490(.A(new_n676), .B(KEYINPUT103), .ZN(new_n677));
  XNOR2_X1  g491(.A(new_n675), .B(new_n677), .ZN(G12));
  AND3_X1   g492(.A1(new_n630), .A2(new_n558), .A3(new_n631), .ZN(new_n679));
  INV_X1    g493(.A(G900), .ZN(new_n680));
  NAND2_X1  g494(.A1(new_n192), .A2(new_n680), .ZN(new_n681));
  OR2_X1    g495(.A1(new_n681), .A2(KEYINPUT104), .ZN(new_n682));
  INV_X1    g496(.A(new_n189), .ZN(new_n683));
  NAND2_X1  g497(.A1(new_n681), .A2(KEYINPUT104), .ZN(new_n684));
  NAND3_X1  g498(.A1(new_n682), .A2(new_n683), .A3(new_n684), .ZN(new_n685));
  INV_X1    g499(.A(new_n685), .ZN(new_n686));
  NOR4_X1   g500(.A1(new_n671), .A2(new_n659), .A3(new_n252), .A4(new_n686), .ZN(new_n687));
  NAND3_X1  g501(.A1(new_n622), .A2(new_n679), .A3(new_n687), .ZN(new_n688));
  XNOR2_X1  g502(.A(new_n688), .B(G128), .ZN(G30));
  INV_X1    g503(.A(new_n659), .ZN(new_n690));
  INV_X1    g504(.A(new_n187), .ZN(new_n691));
  NOR4_X1   g505(.A1(new_n672), .A2(new_n690), .A3(new_n691), .A4(new_n252), .ZN(new_n692));
  INV_X1    g506(.A(KEYINPUT105), .ZN(new_n693));
  NAND2_X1  g507(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  AOI21_X1  g508(.A(new_n521), .B1(new_n539), .B2(new_n517), .ZN(new_n695));
  AOI21_X1  g509(.A(new_n695), .B1(new_n523), .B2(new_n526), .ZN(new_n696));
  OAI21_X1  g510(.A(G472), .B1(new_n696), .B2(G902), .ZN(new_n697));
  NAND3_X1  g511(.A1(new_n546), .A2(new_n547), .A3(new_n697), .ZN(new_n698));
  NAND2_X1  g512(.A1(new_n694), .A2(new_n698), .ZN(new_n699));
  NAND2_X1  g513(.A1(new_n426), .A2(new_n429), .ZN(new_n700));
  XNOR2_X1  g514(.A(new_n700), .B(KEYINPUT38), .ZN(new_n701));
  NOR2_X1   g515(.A1(new_n692), .A2(new_n693), .ZN(new_n702));
  NOR3_X1   g516(.A1(new_n699), .A2(new_n701), .A3(new_n702), .ZN(new_n703));
  XNOR2_X1  g517(.A(new_n685), .B(KEYINPUT39), .ZN(new_n704));
  NAND2_X1  g518(.A1(new_n622), .A2(new_n704), .ZN(new_n705));
  OR2_X1    g519(.A1(new_n705), .A2(KEYINPUT40), .ZN(new_n706));
  NAND2_X1  g520(.A1(new_n705), .A2(KEYINPUT40), .ZN(new_n707));
  AND3_X1   g521(.A1(new_n703), .A2(new_n706), .A3(new_n707), .ZN(new_n708));
  XOR2_X1   g522(.A(KEYINPUT106), .B(G143), .Z(new_n709));
  XNOR2_X1  g523(.A(new_n708), .B(new_n709), .ZN(G45));
  NAND2_X1  g524(.A1(new_n652), .A2(new_n685), .ZN(new_n711));
  NOR2_X1   g525(.A1(new_n711), .A2(new_n671), .ZN(new_n712));
  NAND3_X1  g526(.A1(new_n622), .A2(new_n679), .A3(new_n712), .ZN(new_n713));
  XNOR2_X1  g527(.A(new_n713), .B(G146), .ZN(G48));
  OAI21_X1  g528(.A(new_n191), .B1(new_n607), .B2(new_n608), .ZN(new_n715));
  NOR2_X1   g529(.A1(new_n500), .A2(KEYINPUT107), .ZN(new_n716));
  NAND2_X1  g530(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  INV_X1    g531(.A(new_n716), .ZN(new_n718));
  OAI211_X1 g532(.A(new_n191), .B(new_n718), .C1(new_n607), .C2(new_n608), .ZN(new_n719));
  NAND3_X1  g533(.A1(new_n717), .A2(new_n619), .A3(new_n719), .ZN(new_n720));
  INV_X1    g534(.A(new_n558), .ZN(new_n721));
  INV_X1    g535(.A(new_n596), .ZN(new_n722));
  NOR3_X1   g536(.A1(new_n720), .A2(new_n721), .A3(new_n722), .ZN(new_n723));
  INV_X1    g537(.A(new_n723), .ZN(new_n724));
  NOR2_X1   g538(.A1(new_n655), .A2(new_n724), .ZN(new_n725));
  XOR2_X1   g539(.A(KEYINPUT41), .B(G113), .Z(new_n726));
  XNOR2_X1  g540(.A(new_n725), .B(new_n726), .ZN(G15));
  NOR2_X1   g541(.A1(new_n661), .A2(new_n724), .ZN(new_n728));
  XNOR2_X1  g542(.A(new_n728), .B(new_n206), .ZN(G18));
  NOR2_X1   g543(.A1(new_n632), .A2(new_n720), .ZN(new_n730));
  AND3_X1   g544(.A1(new_n558), .A2(new_n319), .A3(new_n672), .ZN(new_n731));
  NAND2_X1  g545(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  XNOR2_X1  g546(.A(new_n732), .B(G119), .ZN(G21));
  NAND4_X1  g547(.A1(new_n717), .A2(new_n619), .A3(new_n195), .A4(new_n719), .ZN(new_n734));
  INV_X1    g548(.A(KEYINPUT108), .ZN(new_n735));
  AOI21_X1  g549(.A(new_n735), .B1(new_n624), .B2(new_n596), .ZN(new_n736));
  NAND2_X1  g550(.A1(new_n623), .A2(G472), .ZN(new_n737));
  NAND2_X1  g551(.A1(new_n543), .A2(new_n544), .ZN(new_n738));
  AND4_X1   g552(.A1(new_n735), .A2(new_n737), .A3(new_n596), .A4(new_n738), .ZN(new_n739));
  NOR3_X1   g553(.A1(new_n734), .A2(new_n736), .A3(new_n739), .ZN(new_n740));
  NOR2_X1   g554(.A1(new_n690), .A2(new_n252), .ZN(new_n741));
  AND3_X1   g555(.A1(new_n630), .A2(new_n631), .A3(new_n741), .ZN(new_n742));
  NAND2_X1  g556(.A1(new_n740), .A2(new_n742), .ZN(new_n743));
  XNOR2_X1  g557(.A(new_n743), .B(G122), .ZN(G24));
  NAND4_X1  g558(.A1(new_n652), .A2(new_n624), .A3(new_n672), .A4(new_n685), .ZN(new_n745));
  NOR3_X1   g559(.A1(new_n632), .A2(new_n720), .A3(new_n745), .ZN(new_n746));
  XNOR2_X1  g560(.A(new_n746), .B(new_n261), .ZN(G27));
  AOI21_X1  g561(.A(new_n691), .B1(new_n426), .B2(new_n429), .ZN(new_n748));
  AND2_X1   g562(.A1(new_n748), .A2(new_n613), .ZN(new_n749));
  INV_X1    g563(.A(new_n711), .ZN(new_n750));
  OAI211_X1 g564(.A(new_n557), .B(new_n547), .C1(KEYINPUT109), .C2(new_n545), .ZN(new_n751));
  AND2_X1   g565(.A1(new_n545), .A2(KEYINPUT109), .ZN(new_n752));
  OAI21_X1  g566(.A(new_n596), .B1(new_n751), .B2(new_n752), .ZN(new_n753));
  INV_X1    g567(.A(new_n753), .ZN(new_n754));
  NAND3_X1  g568(.A1(new_n749), .A2(new_n750), .A3(new_n754), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n755), .A2(KEYINPUT42), .ZN(new_n756));
  NOR2_X1   g570(.A1(new_n711), .A2(KEYINPUT42), .ZN(new_n757));
  NAND3_X1  g571(.A1(new_n749), .A2(new_n597), .A3(new_n757), .ZN(new_n758));
  AND2_X1   g572(.A1(new_n756), .A2(new_n758), .ZN(new_n759));
  XNOR2_X1  g573(.A(new_n759), .B(G131), .ZN(G33));
  INV_X1    g574(.A(new_n252), .ZN(new_n761));
  NOR2_X1   g575(.A1(new_n659), .A2(new_n686), .ZN(new_n762));
  NAND4_X1  g576(.A1(new_n749), .A2(new_n597), .A3(new_n761), .A4(new_n762), .ZN(new_n763));
  XNOR2_X1  g577(.A(new_n763), .B(G134), .ZN(G36));
  AND2_X1   g578(.A1(new_n649), .A2(new_n651), .ZN(new_n765));
  NOR2_X1   g579(.A1(new_n765), .A2(new_n659), .ZN(new_n766));
  INV_X1    g580(.A(KEYINPUT43), .ZN(new_n767));
  INV_X1    g581(.A(KEYINPUT111), .ZN(new_n768));
  OAI21_X1  g582(.A(new_n767), .B1(new_n659), .B2(new_n768), .ZN(new_n769));
  XNOR2_X1  g583(.A(new_n766), .B(new_n769), .ZN(new_n770));
  NOR2_X1   g584(.A1(new_n624), .A2(new_n671), .ZN(new_n771));
  NAND2_X1  g585(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  INV_X1    g586(.A(KEYINPUT44), .ZN(new_n773));
  NAND2_X1  g587(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  NAND3_X1  g588(.A1(new_n770), .A2(KEYINPUT44), .A3(new_n771), .ZN(new_n775));
  NAND3_X1  g589(.A1(new_n774), .A2(new_n748), .A3(new_n775), .ZN(new_n776));
  OAI21_X1  g590(.A(new_n484), .B1(new_n485), .B2(new_n488), .ZN(new_n777));
  INV_X1    g591(.A(KEYINPUT45), .ZN(new_n778));
  AOI21_X1  g592(.A(new_n500), .B1(new_n777), .B2(new_n778), .ZN(new_n779));
  OAI21_X1  g593(.A(new_n779), .B1(new_n778), .B2(new_n777), .ZN(new_n780));
  AND2_X1   g594(.A1(new_n780), .A2(new_n490), .ZN(new_n781));
  OAI21_X1  g595(.A(KEYINPUT110), .B1(new_n781), .B2(KEYINPUT46), .ZN(new_n782));
  NAND2_X1  g596(.A1(new_n781), .A2(KEYINPUT46), .ZN(new_n783));
  NAND3_X1  g597(.A1(new_n782), .A2(new_n609), .A3(new_n783), .ZN(new_n784));
  NOR3_X1   g598(.A1(new_n781), .A2(KEYINPUT110), .A3(KEYINPUT46), .ZN(new_n785));
  OAI211_X1 g599(.A(new_n619), .B(new_n704), .C1(new_n784), .C2(new_n785), .ZN(new_n786));
  NOR2_X1   g600(.A1(new_n776), .A2(new_n786), .ZN(new_n787));
  XNOR2_X1  g601(.A(KEYINPUT112), .B(G137), .ZN(new_n788));
  XNOR2_X1  g602(.A(new_n787), .B(new_n788), .ZN(G39));
  NAND4_X1  g603(.A1(new_n750), .A2(new_n722), .A3(new_n748), .A4(new_n721), .ZN(new_n790));
  OAI21_X1  g604(.A(new_n619), .B1(new_n784), .B2(new_n785), .ZN(new_n791));
  INV_X1    g605(.A(KEYINPUT47), .ZN(new_n792));
  NAND2_X1  g606(.A1(new_n791), .A2(new_n792), .ZN(new_n793));
  OAI211_X1 g607(.A(KEYINPUT47), .B(new_n619), .C1(new_n784), .C2(new_n785), .ZN(new_n794));
  AOI21_X1  g608(.A(new_n790), .B1(new_n793), .B2(new_n794), .ZN(new_n795));
  XNOR2_X1  g609(.A(new_n795), .B(new_n258), .ZN(G42));
  NAND4_X1  g610(.A1(new_n766), .A2(new_n596), .A3(new_n619), .A4(new_n187), .ZN(new_n797));
  NAND2_X1  g611(.A1(new_n717), .A2(new_n719), .ZN(new_n798));
  AOI211_X1 g612(.A(new_n698), .B(new_n797), .C1(KEYINPUT49), .C2(new_n798), .ZN(new_n799));
  NOR2_X1   g613(.A1(new_n798), .A2(KEYINPUT49), .ZN(new_n800));
  XOR2_X1   g614(.A(new_n800), .B(KEYINPUT113), .Z(new_n801));
  NAND3_X1  g615(.A1(new_n799), .A2(new_n701), .A3(new_n801), .ZN(new_n802));
  INV_X1    g616(.A(KEYINPUT54), .ZN(new_n803));
  NOR3_X1   g617(.A1(new_n666), .A2(new_n670), .A3(new_n686), .ZN(new_n804));
  AOI21_X1  g618(.A(KEYINPUT117), .B1(new_n613), .B2(new_n804), .ZN(new_n805));
  AND3_X1   g619(.A1(new_n613), .A2(KEYINPUT117), .A3(new_n804), .ZN(new_n806));
  OAI211_X1 g620(.A(new_n742), .B(new_n698), .C1(new_n805), .C2(new_n806), .ZN(new_n807));
  INV_X1    g621(.A(new_n745), .ZN(new_n808));
  NAND2_X1  g622(.A1(new_n730), .A2(new_n808), .ZN(new_n809));
  NAND4_X1  g623(.A1(new_n807), .A2(new_n688), .A3(new_n713), .A4(new_n809), .ZN(new_n810));
  INV_X1    g624(.A(KEYINPUT52), .ZN(new_n811));
  NAND2_X1  g625(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  NAND3_X1  g626(.A1(new_n630), .A2(new_n558), .A3(new_n631), .ZN(new_n813));
  NOR3_X1   g627(.A1(new_n813), .A2(new_n620), .A3(new_n621), .ZN(new_n814));
  AOI21_X1  g628(.A(new_n746), .B1(new_n814), .B2(new_n687), .ZN(new_n815));
  NAND4_X1  g629(.A1(new_n815), .A2(KEYINPUT52), .A3(new_n713), .A4(new_n807), .ZN(new_n816));
  AOI21_X1  g630(.A(KEYINPUT116), .B1(new_n812), .B2(new_n816), .ZN(new_n817));
  NOR2_X1   g631(.A1(new_n817), .A2(KEYINPUT53), .ZN(new_n818));
  AOI22_X1  g632(.A1(new_n730), .A2(new_n731), .B1(new_n740), .B2(new_n742), .ZN(new_n819));
  AND3_X1   g633(.A1(new_n426), .A2(new_n187), .A3(new_n429), .ZN(new_n820));
  INV_X1    g634(.A(KEYINPUT115), .ZN(new_n821));
  NOR2_X1   g635(.A1(new_n761), .A2(new_n821), .ZN(new_n822));
  NOR2_X1   g636(.A1(new_n252), .A2(KEYINPUT115), .ZN(new_n823));
  OAI211_X1 g637(.A(new_n195), .B(new_n690), .C1(new_n822), .C2(new_n823), .ZN(new_n824));
  INV_X1    g638(.A(new_n824), .ZN(new_n825));
  NAND4_X1  g639(.A1(new_n622), .A2(new_n820), .A3(new_n625), .A4(new_n825), .ZN(new_n826));
  OAI211_X1 g640(.A(new_n723), .B(new_n633), .C1(new_n654), .C2(new_n660), .ZN(new_n827));
  NAND4_X1  g641(.A1(new_n819), .A2(new_n675), .A3(new_n826), .A4(new_n827), .ZN(new_n828));
  INV_X1    g642(.A(KEYINPUT114), .ZN(new_n829));
  NAND4_X1  g643(.A1(new_n505), .A2(new_n820), .A3(new_n615), .A4(new_n625), .ZN(new_n830));
  INV_X1    g644(.A(new_n654), .ZN(new_n831));
  OAI211_X1 g645(.A(new_n616), .B(new_n829), .C1(new_n830), .C2(new_n831), .ZN(new_n832));
  INV_X1    g646(.A(new_n832), .ZN(new_n833));
  NAND4_X1  g647(.A1(new_n622), .A2(new_n820), .A3(new_n625), .A4(new_n654), .ZN(new_n834));
  AOI21_X1  g648(.A(new_n829), .B1(new_n834), .B2(new_n616), .ZN(new_n835));
  NOR3_X1   g649(.A1(new_n828), .A2(new_n833), .A3(new_n835), .ZN(new_n836));
  NAND2_X1  g650(.A1(new_n812), .A2(new_n816), .ZN(new_n837));
  NAND2_X1  g651(.A1(new_n700), .A2(new_n187), .ZN(new_n838));
  XNOR2_X1  g652(.A(new_n252), .B(new_n821), .ZN(new_n839));
  NAND3_X1  g653(.A1(new_n839), .A2(new_n672), .A3(new_n762), .ZN(new_n840));
  NOR3_X1   g654(.A1(new_n838), .A2(new_n840), .A3(new_n721), .ZN(new_n841));
  AOI22_X1  g655(.A1(new_n841), .A2(new_n622), .B1(new_n749), .B2(new_n808), .ZN(new_n842));
  NAND4_X1  g656(.A1(new_n842), .A2(new_n756), .A3(new_n758), .A4(new_n763), .ZN(new_n843));
  INV_X1    g657(.A(new_n843), .ZN(new_n844));
  NAND3_X1  g658(.A1(new_n836), .A2(new_n837), .A3(new_n844), .ZN(new_n845));
  NAND2_X1  g659(.A1(new_n818), .A2(new_n845), .ZN(new_n846));
  AOI21_X1  g660(.A(new_n843), .B1(new_n812), .B2(new_n816), .ZN(new_n847));
  OAI211_X1 g661(.A(new_n847), .B(new_n836), .C1(new_n817), .C2(KEYINPUT53), .ZN(new_n848));
  AOI21_X1  g662(.A(new_n803), .B1(new_n846), .B2(new_n848), .ZN(new_n849));
  NAND2_X1  g663(.A1(new_n845), .A2(KEYINPUT53), .ZN(new_n850));
  INV_X1    g664(.A(KEYINPUT53), .ZN(new_n851));
  NAND3_X1  g665(.A1(new_n847), .A2(new_n851), .A3(new_n836), .ZN(new_n852));
  AOI21_X1  g666(.A(KEYINPUT54), .B1(new_n850), .B2(new_n852), .ZN(new_n853));
  NOR2_X1   g667(.A1(new_n849), .A2(new_n853), .ZN(new_n854));
  AND2_X1   g668(.A1(new_n770), .A2(new_n189), .ZN(new_n855));
  NOR2_X1   g669(.A1(new_n838), .A2(new_n720), .ZN(new_n856));
  AND2_X1   g670(.A1(new_n855), .A2(new_n856), .ZN(new_n857));
  NAND2_X1  g671(.A1(new_n857), .A2(new_n754), .ZN(new_n858));
  XNOR2_X1  g672(.A(new_n858), .B(KEYINPUT48), .ZN(new_n859));
  NOR3_X1   g673(.A1(new_n698), .A2(new_n722), .A3(new_n683), .ZN(new_n860));
  AND2_X1   g674(.A1(new_n856), .A2(new_n860), .ZN(new_n861));
  NAND2_X1  g675(.A1(new_n861), .A2(new_n652), .ZN(new_n862));
  NOR2_X1   g676(.A1(new_n739), .A2(new_n736), .ZN(new_n863));
  NAND2_X1  g677(.A1(new_n855), .A2(new_n863), .ZN(new_n864));
  INV_X1    g678(.A(new_n864), .ZN(new_n865));
  AOI211_X1 g679(.A(new_n188), .B(G953), .C1(new_n865), .C2(new_n730), .ZN(new_n866));
  NAND3_X1  g680(.A1(new_n859), .A2(new_n862), .A3(new_n866), .ZN(new_n867));
  NAND2_X1  g681(.A1(new_n857), .A2(new_n674), .ZN(new_n868));
  NAND3_X1  g682(.A1(new_n861), .A2(new_n690), .A3(new_n765), .ZN(new_n869));
  NAND2_X1  g683(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  OAI211_X1 g684(.A(new_n793), .B(new_n794), .C1(new_n619), .C2(new_n798), .ZN(new_n871));
  NOR2_X1   g685(.A1(new_n864), .A2(new_n838), .ZN(new_n872));
  AOI21_X1  g686(.A(new_n870), .B1(new_n871), .B2(new_n872), .ZN(new_n873));
  INV_X1    g687(.A(KEYINPUT51), .ZN(new_n874));
  NOR2_X1   g688(.A1(new_n720), .A2(new_n187), .ZN(new_n875));
  AND2_X1   g689(.A1(new_n701), .A2(new_n875), .ZN(new_n876));
  NAND2_X1  g690(.A1(new_n865), .A2(new_n876), .ZN(new_n877));
  INV_X1    g691(.A(KEYINPUT50), .ZN(new_n878));
  NAND2_X1  g692(.A1(new_n877), .A2(new_n878), .ZN(new_n879));
  NAND3_X1  g693(.A1(new_n865), .A2(KEYINPUT50), .A3(new_n876), .ZN(new_n880));
  AOI21_X1  g694(.A(new_n874), .B1(new_n879), .B2(new_n880), .ZN(new_n881));
  AOI21_X1  g695(.A(new_n867), .B1(new_n873), .B2(new_n881), .ZN(new_n882));
  NAND2_X1  g696(.A1(new_n879), .A2(new_n880), .ZN(new_n883));
  INV_X1    g697(.A(KEYINPUT118), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  NAND3_X1  g699(.A1(new_n879), .A2(KEYINPUT118), .A3(new_n880), .ZN(new_n886));
  NAND3_X1  g700(.A1(new_n885), .A2(new_n873), .A3(new_n886), .ZN(new_n887));
  NAND2_X1  g701(.A1(new_n887), .A2(new_n874), .ZN(new_n888));
  AND3_X1   g702(.A1(new_n854), .A2(new_n882), .A3(new_n888), .ZN(new_n889));
  NAND2_X1  g703(.A1(new_n188), .A2(new_n190), .ZN(new_n890));
  XNOR2_X1  g704(.A(new_n890), .B(KEYINPUT119), .ZN(new_n891));
  OAI21_X1  g705(.A(new_n802), .B1(new_n889), .B2(new_n891), .ZN(G75));
  NOR2_X1   g706(.A1(new_n190), .A2(G952), .ZN(new_n893));
  AND2_X1   g707(.A1(new_n375), .A2(new_n377), .ZN(new_n894));
  XNOR2_X1  g708(.A(new_n894), .B(new_n406), .ZN(new_n895));
  XOR2_X1   g709(.A(new_n895), .B(KEYINPUT55), .Z(new_n896));
  NAND4_X1  g710(.A1(new_n850), .A2(new_n249), .A3(new_n423), .A4(new_n852), .ZN(new_n897));
  INV_X1    g711(.A(KEYINPUT56), .ZN(new_n898));
  AOI21_X1  g712(.A(new_n896), .B1(new_n897), .B2(new_n898), .ZN(new_n899));
  XOR2_X1   g713(.A(new_n896), .B(KEYINPUT120), .Z(new_n900));
  NAND3_X1  g714(.A1(new_n897), .A2(new_n898), .A3(new_n900), .ZN(new_n901));
  OR2_X1    g715(.A1(new_n901), .A2(KEYINPUT121), .ZN(new_n902));
  NAND2_X1  g716(.A1(new_n901), .A2(KEYINPUT121), .ZN(new_n903));
  AOI211_X1 g717(.A(new_n893), .B(new_n899), .C1(new_n902), .C2(new_n903), .ZN(G51));
  AND3_X1   g718(.A1(new_n847), .A2(new_n851), .A3(new_n836), .ZN(new_n905));
  AOI21_X1  g719(.A(new_n851), .B1(new_n847), .B2(new_n836), .ZN(new_n906));
  NOR4_X1   g720(.A1(new_n905), .A2(new_n906), .A3(new_n191), .A4(new_n780), .ZN(new_n907));
  XOR2_X1   g721(.A(new_n490), .B(KEYINPUT57), .Z(new_n908));
  NOR3_X1   g722(.A1(new_n905), .A2(new_n906), .A3(new_n803), .ZN(new_n909));
  OAI21_X1  g723(.A(new_n908), .B1(new_n909), .B2(new_n853), .ZN(new_n910));
  NOR2_X1   g724(.A1(new_n607), .A2(new_n608), .ZN(new_n911));
  INV_X1    g725(.A(new_n911), .ZN(new_n912));
  AOI21_X1  g726(.A(new_n907), .B1(new_n910), .B2(new_n912), .ZN(new_n913));
  OAI21_X1  g727(.A(KEYINPUT122), .B1(new_n913), .B2(new_n893), .ZN(new_n914));
  INV_X1    g728(.A(KEYINPUT122), .ZN(new_n915));
  INV_X1    g729(.A(new_n893), .ZN(new_n916));
  OAI21_X1  g730(.A(new_n803), .B1(new_n905), .B2(new_n906), .ZN(new_n917));
  NAND3_X1  g731(.A1(new_n850), .A2(KEYINPUT54), .A3(new_n852), .ZN(new_n918));
  NAND2_X1  g732(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  AOI21_X1  g733(.A(new_n911), .B1(new_n919), .B2(new_n908), .ZN(new_n920));
  OAI211_X1 g734(.A(new_n915), .B(new_n916), .C1(new_n920), .C2(new_n907), .ZN(new_n921));
  NAND2_X1  g735(.A1(new_n914), .A2(new_n921), .ZN(G54));
  NOR3_X1   g736(.A1(new_n905), .A2(new_n906), .A3(new_n191), .ZN(new_n923));
  NAND3_X1  g737(.A1(new_n923), .A2(KEYINPUT58), .A3(G475), .ZN(new_n924));
  NOR2_X1   g738(.A1(new_n292), .A2(new_n306), .ZN(new_n925));
  OAI21_X1  g739(.A(KEYINPUT123), .B1(new_n924), .B2(new_n925), .ZN(new_n926));
  AOI21_X1  g740(.A(new_n893), .B1(new_n924), .B2(new_n925), .ZN(new_n927));
  NAND2_X1  g741(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  NOR3_X1   g742(.A1(new_n924), .A2(KEYINPUT123), .A3(new_n925), .ZN(new_n929));
  NOR2_X1   g743(.A1(new_n928), .A2(new_n929), .ZN(G60));
  NAND2_X1  g744(.A1(G478), .A2(G902), .ZN(new_n931));
  XOR2_X1   g745(.A(new_n931), .B(KEYINPUT59), .Z(new_n932));
  INV_X1    g746(.A(new_n932), .ZN(new_n933));
  NAND3_X1  g747(.A1(new_n919), .A2(new_n646), .A3(new_n933), .ZN(new_n934));
  NAND2_X1  g748(.A1(new_n934), .A2(new_n916), .ZN(new_n935));
  INV_X1    g749(.A(new_n646), .ZN(new_n936));
  OAI21_X1  g750(.A(new_n936), .B1(new_n854), .B2(new_n932), .ZN(new_n937));
  INV_X1    g751(.A(KEYINPUT124), .ZN(new_n938));
  NAND2_X1  g752(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  OAI211_X1 g753(.A(KEYINPUT124), .B(new_n936), .C1(new_n854), .C2(new_n932), .ZN(new_n940));
  AOI21_X1  g754(.A(new_n935), .B1(new_n939), .B2(new_n940), .ZN(G63));
  NAND2_X1  g755(.A1(G217), .A2(G902), .ZN(new_n942));
  XNOR2_X1  g756(.A(new_n942), .B(KEYINPUT60), .ZN(new_n943));
  NOR3_X1   g757(.A1(new_n905), .A2(new_n906), .A3(new_n943), .ZN(new_n944));
  NAND2_X1  g758(.A1(new_n944), .A2(new_n668), .ZN(new_n945));
  INV_X1    g759(.A(new_n586), .ZN(new_n946));
  INV_X1    g760(.A(new_n589), .ZN(new_n947));
  NOR2_X1   g761(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  OAI211_X1 g762(.A(new_n945), .B(new_n916), .C1(new_n948), .C2(new_n944), .ZN(new_n949));
  INV_X1    g763(.A(KEYINPUT61), .ZN(new_n950));
  XNOR2_X1  g764(.A(new_n949), .B(new_n950), .ZN(G66));
  INV_X1    g765(.A(new_n193), .ZN(new_n952));
  AOI21_X1  g766(.A(new_n190), .B1(new_n403), .B2(new_n952), .ZN(new_n953));
  INV_X1    g767(.A(new_n836), .ZN(new_n954));
  AOI21_X1  g768(.A(new_n953), .B1(new_n954), .B2(new_n190), .ZN(new_n955));
  INV_X1    g769(.A(G898), .ZN(new_n956));
  AOI21_X1  g770(.A(new_n894), .B1(new_n956), .B2(G953), .ZN(new_n957));
  XNOR2_X1  g771(.A(new_n955), .B(new_n957), .ZN(G69));
  INV_X1    g772(.A(KEYINPUT126), .ZN(new_n959));
  INV_X1    g773(.A(new_n786), .ZN(new_n960));
  INV_X1    g774(.A(new_n776), .ZN(new_n961));
  AND2_X1   g775(.A1(new_n742), .A2(new_n754), .ZN(new_n962));
  OAI21_X1  g776(.A(new_n960), .B1(new_n961), .B2(new_n962), .ZN(new_n963));
  INV_X1    g777(.A(new_n795), .ZN(new_n964));
  NAND2_X1  g778(.A1(new_n759), .A2(new_n763), .ZN(new_n965));
  NAND2_X1  g779(.A1(new_n815), .A2(new_n713), .ZN(new_n966));
  NOR2_X1   g780(.A1(new_n965), .A2(new_n966), .ZN(new_n967));
  NAND3_X1  g781(.A1(new_n963), .A2(new_n964), .A3(new_n967), .ZN(new_n968));
  OR2_X1    g782(.A1(new_n968), .A2(G953), .ZN(new_n969));
  XNOR2_X1  g783(.A(new_n516), .B(new_n280), .ZN(new_n970));
  INV_X1    g784(.A(new_n970), .ZN(new_n971));
  AOI21_X1  g785(.A(new_n971), .B1(G900), .B2(G953), .ZN(new_n972));
  AOI21_X1  g786(.A(new_n959), .B1(new_n969), .B2(new_n972), .ZN(new_n973));
  INV_X1    g787(.A(KEYINPUT125), .ZN(new_n974));
  OR3_X1    g788(.A1(new_n708), .A2(KEYINPUT62), .A3(new_n966), .ZN(new_n975));
  OAI21_X1  g789(.A(KEYINPUT62), .B1(new_n708), .B2(new_n966), .ZN(new_n976));
  OAI21_X1  g790(.A(new_n653), .B1(new_n659), .B2(new_n839), .ZN(new_n977));
  NAND3_X1  g791(.A1(new_n977), .A2(new_n597), .A3(new_n748), .ZN(new_n978));
  NOR2_X1   g792(.A1(new_n705), .A2(new_n978), .ZN(new_n979));
  NOR2_X1   g793(.A1(new_n787), .A2(new_n979), .ZN(new_n980));
  NAND4_X1  g794(.A1(new_n975), .A2(new_n964), .A3(new_n976), .A4(new_n980), .ZN(new_n981));
  NAND2_X1  g795(.A1(new_n981), .A2(new_n190), .ZN(new_n982));
  AOI21_X1  g796(.A(new_n974), .B1(new_n982), .B2(new_n971), .ZN(new_n983));
  AOI211_X1 g797(.A(KEYINPUT125), .B(new_n970), .C1(new_n981), .C2(new_n190), .ZN(new_n984));
  OAI21_X1  g798(.A(new_n973), .B1(new_n983), .B2(new_n984), .ZN(new_n985));
  AOI21_X1  g799(.A(new_n190), .B1(G227), .B2(G900), .ZN(new_n986));
  NAND2_X1  g800(.A1(new_n985), .A2(new_n986), .ZN(new_n987));
  INV_X1    g801(.A(new_n986), .ZN(new_n988));
  OAI211_X1 g802(.A(new_n988), .B(new_n973), .C1(new_n983), .C2(new_n984), .ZN(new_n989));
  NAND2_X1  g803(.A1(new_n987), .A2(new_n989), .ZN(G72));
  NAND2_X1  g804(.A1(G472), .A2(G902), .ZN(new_n991));
  XOR2_X1   g805(.A(new_n991), .B(KEYINPUT63), .Z(new_n992));
  OAI21_X1  g806(.A(new_n992), .B1(new_n981), .B2(new_n954), .ZN(new_n993));
  NAND3_X1  g807(.A1(new_n993), .A2(new_n521), .A3(new_n553), .ZN(new_n994));
  NAND2_X1  g808(.A1(new_n846), .A2(new_n848), .ZN(new_n995));
  OAI21_X1  g809(.A(new_n535), .B1(new_n554), .B2(new_n521), .ZN(new_n996));
  NAND3_X1  g810(.A1(new_n995), .A2(new_n992), .A3(new_n996), .ZN(new_n997));
  OAI21_X1  g811(.A(new_n992), .B1(new_n968), .B2(new_n954), .ZN(new_n998));
  NAND2_X1  g812(.A1(new_n554), .A2(new_n537), .ZN(new_n999));
  XNOR2_X1  g813(.A(new_n999), .B(KEYINPUT127), .ZN(new_n1000));
  AOI21_X1  g814(.A(new_n893), .B1(new_n998), .B2(new_n1000), .ZN(new_n1001));
  AND3_X1   g815(.A1(new_n994), .A2(new_n997), .A3(new_n1001), .ZN(G57));
endmodule


