//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 1 1 0 0 0 1 0 1 0 1 1 1 0 0 1 1 1 0 1 1 0 1 1 1 1 0 1 1 0 0 1 0 1 1 0 0 0 1 0 1 1 0 0 0 0 0 0 1 1 0 1 0 1 0 1 1 0 1 0 0 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:37:21 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n203, new_n204, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n245, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n600, new_n601, new_n602, new_n603, new_n604, new_n605,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n805, new_n806,
    new_n807, new_n808, new_n809, new_n810, new_n811, new_n812, new_n813,
    new_n814, new_n815, new_n816, new_n817, new_n818, new_n819, new_n820,
    new_n821, new_n822, new_n823, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n984, new_n985, new_n986, new_n987, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1018, new_n1019, new_n1020, new_n1021, new_n1022,
    new_n1023, new_n1024, new_n1025, new_n1026, new_n1027, new_n1028,
    new_n1029, new_n1030, new_n1031, new_n1032, new_n1033, new_n1034,
    new_n1035, new_n1036, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1046, new_n1047,
    new_n1048, new_n1049, new_n1050, new_n1051, new_n1052, new_n1053,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1115, new_n1116, new_n1117, new_n1118, new_n1119, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1179, new_n1180, new_n1181,
    new_n1182, new_n1183, new_n1184, new_n1185, new_n1186, new_n1187,
    new_n1188, new_n1189, new_n1190, new_n1191, new_n1192, new_n1193,
    new_n1194, new_n1195, new_n1196, new_n1197, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1205, new_n1206, new_n1207,
    new_n1208, new_n1210, new_n1211, new_n1212, new_n1213, new_n1214,
    new_n1215, new_n1216, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1267, new_n1268, new_n1269,
    new_n1270, new_n1271, new_n1272, new_n1273;
  NOR4_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .A4(G77), .ZN(G353));
  OAI21_X1  g0001(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0002(.A1(G1), .A2(G20), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G13), .ZN(new_n204));
  OAI211_X1 g0004(.A(new_n204), .B(G250), .C1(G257), .C2(G264), .ZN(new_n205));
  XOR2_X1   g0005(.A(new_n205), .B(KEYINPUT0), .Z(new_n206));
  AOI22_X1  g0006(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n207));
  INV_X1    g0007(.A(G68), .ZN(new_n208));
  INV_X1    g0008(.A(G238), .ZN(new_n209));
  INV_X1    g0009(.A(G107), .ZN(new_n210));
  INV_X1    g0010(.A(G264), .ZN(new_n211));
  OAI221_X1 g0011(.A(new_n207), .B1(new_n208), .B2(new_n209), .C1(new_n210), .C2(new_n211), .ZN(new_n212));
  AOI21_X1  g0012(.A(new_n212), .B1(G116), .B2(G270), .ZN(new_n213));
  INV_X1    g0013(.A(G50), .ZN(new_n214));
  INV_X1    g0014(.A(G226), .ZN(new_n215));
  INV_X1    g0015(.A(G77), .ZN(new_n216));
  INV_X1    g0016(.A(G244), .ZN(new_n217));
  OAI221_X1 g0017(.A(new_n213), .B1(new_n214), .B2(new_n215), .C1(new_n216), .C2(new_n217), .ZN(new_n218));
  INV_X1    g0018(.A(G58), .ZN(new_n219));
  INV_X1    g0019(.A(G232), .ZN(new_n220));
  NOR2_X1   g0020(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  OAI21_X1  g0021(.A(new_n203), .B1(new_n218), .B2(new_n221), .ZN(new_n222));
  XNOR2_X1  g0022(.A(new_n222), .B(KEYINPUT1), .ZN(new_n223));
  NAND2_X1  g0023(.A1(G1), .A2(G13), .ZN(new_n224));
  INV_X1    g0024(.A(G20), .ZN(new_n225));
  NOR2_X1   g0025(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  OAI21_X1  g0026(.A(G50), .B1(G58), .B2(G68), .ZN(new_n227));
  INV_X1    g0027(.A(new_n227), .ZN(new_n228));
  AOI211_X1 g0028(.A(new_n206), .B(new_n223), .C1(new_n226), .C2(new_n228), .ZN(G361));
  XNOR2_X1  g0029(.A(G238), .B(G244), .ZN(new_n230));
  XNOR2_X1  g0030(.A(G226), .B(G232), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n230), .B(new_n231), .ZN(new_n232));
  XNOR2_X1  g0032(.A(KEYINPUT64), .B(KEYINPUT2), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n232), .B(new_n233), .ZN(new_n234));
  XNOR2_X1  g0034(.A(G250), .B(G257), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n235), .B(new_n211), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n236), .B(G270), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n234), .B(new_n237), .ZN(G358));
  XNOR2_X1  g0038(.A(G50), .B(G58), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n239), .B(KEYINPUT65), .ZN(new_n240));
  XNOR2_X1  g0040(.A(G68), .B(G77), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XOR2_X1   g0042(.A(G97), .B(G107), .Z(new_n243));
  XNOR2_X1  g0043(.A(G87), .B(G116), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n242), .B(new_n245), .ZN(G351));
  NAND3_X1  g0046(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n247));
  NAND2_X1  g0047(.A1(new_n247), .A2(new_n224), .ZN(new_n248));
  XNOR2_X1  g0048(.A(KEYINPUT8), .B(G58), .ZN(new_n249));
  NAND2_X1  g0049(.A1(new_n225), .A2(G33), .ZN(new_n250));
  NOR2_X1   g0050(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  NOR3_X1   g0051(.A1(G50), .A2(G58), .A3(G68), .ZN(new_n252));
  INV_X1    g0052(.A(G33), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n225), .A2(new_n253), .ZN(new_n254));
  INV_X1    g0054(.A(G150), .ZN(new_n255));
  OAI22_X1  g0055(.A1(new_n252), .A2(new_n225), .B1(new_n254), .B2(new_n255), .ZN(new_n256));
  OAI21_X1  g0056(.A(new_n248), .B1(new_n251), .B2(new_n256), .ZN(new_n257));
  XNOR2_X1  g0057(.A(new_n257), .B(KEYINPUT67), .ZN(new_n258));
  INV_X1    g0058(.A(G1), .ZN(new_n259));
  NAND3_X1  g0059(.A1(new_n259), .A2(G13), .A3(G20), .ZN(new_n260));
  INV_X1    g0060(.A(new_n260), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n261), .A2(new_n214), .ZN(new_n262));
  AOI21_X1  g0062(.A(new_n248), .B1(new_n259), .B2(G20), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n263), .A2(G50), .ZN(new_n264));
  NAND3_X1  g0064(.A1(new_n258), .A2(new_n262), .A3(new_n264), .ZN(new_n265));
  INV_X1    g0065(.A(new_n265), .ZN(new_n266));
  INV_X1    g0066(.A(KEYINPUT3), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n267), .A2(new_n253), .ZN(new_n268));
  NAND2_X1  g0068(.A1(KEYINPUT3), .A2(G33), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  INV_X1    g0070(.A(G1698), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n271), .A2(G222), .ZN(new_n272));
  NAND2_X1  g0072(.A1(G223), .A2(G1698), .ZN(new_n273));
  NAND3_X1  g0073(.A1(new_n270), .A2(new_n272), .A3(new_n273), .ZN(new_n274));
  AOI21_X1  g0074(.A(new_n224), .B1(G33), .B2(G41), .ZN(new_n275));
  OAI211_X1 g0075(.A(new_n274), .B(new_n275), .C1(G77), .C2(new_n270), .ZN(new_n276));
  OAI21_X1  g0076(.A(new_n259), .B1(G41), .B2(G45), .ZN(new_n277));
  INV_X1    g0077(.A(G274), .ZN(new_n278));
  NOR2_X1   g0078(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  INV_X1    g0079(.A(new_n279), .ZN(new_n280));
  INV_X1    g0080(.A(G41), .ZN(new_n281));
  OAI211_X1 g0081(.A(G1), .B(G13), .C1(new_n253), .C2(new_n281), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n282), .A2(new_n277), .ZN(new_n283));
  OAI211_X1 g0083(.A(new_n276), .B(new_n280), .C1(new_n215), .C2(new_n283), .ZN(new_n284));
  INV_X1    g0084(.A(KEYINPUT66), .ZN(new_n285));
  XNOR2_X1  g0085(.A(new_n284), .B(new_n285), .ZN(new_n286));
  AOI22_X1  g0086(.A1(KEYINPUT9), .A2(new_n266), .B1(new_n286), .B2(G190), .ZN(new_n287));
  INV_X1    g0087(.A(new_n286), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n288), .A2(G200), .ZN(new_n289));
  OAI211_X1 g0089(.A(new_n287), .B(new_n289), .C1(KEYINPUT9), .C2(new_n266), .ZN(new_n290));
  XNOR2_X1  g0090(.A(new_n290), .B(KEYINPUT10), .ZN(new_n291));
  INV_X1    g0091(.A(G169), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n288), .A2(new_n292), .ZN(new_n293));
  INV_X1    g0093(.A(G179), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n286), .A2(new_n294), .ZN(new_n295));
  NAND3_X1  g0095(.A1(new_n293), .A2(new_n265), .A3(new_n295), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n291), .A2(new_n296), .ZN(new_n297));
  INV_X1    g0097(.A(new_n297), .ZN(new_n298));
  NAND2_X1  g0098(.A1(G238), .A2(G1698), .ZN(new_n299));
  OAI211_X1 g0099(.A(new_n270), .B(new_n299), .C1(new_n220), .C2(G1698), .ZN(new_n300));
  OAI211_X1 g0100(.A(new_n300), .B(new_n275), .C1(G107), .C2(new_n270), .ZN(new_n301));
  OAI211_X1 g0101(.A(new_n301), .B(new_n280), .C1(new_n217), .C2(new_n283), .ZN(new_n302));
  XNOR2_X1  g0102(.A(new_n302), .B(KEYINPUT68), .ZN(new_n303));
  INV_X1    g0103(.A(new_n303), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n304), .A2(G200), .ZN(new_n305));
  INV_X1    g0105(.A(new_n249), .ZN(new_n306));
  INV_X1    g0106(.A(new_n254), .ZN(new_n307));
  AOI22_X1  g0107(.A1(new_n306), .A2(new_n307), .B1(G20), .B2(G77), .ZN(new_n308));
  XOR2_X1   g0108(.A(KEYINPUT15), .B(G87), .Z(new_n309));
  INV_X1    g0109(.A(new_n309), .ZN(new_n310));
  OAI21_X1  g0110(.A(new_n308), .B1(new_n250), .B2(new_n310), .ZN(new_n311));
  AOI22_X1  g0111(.A1(new_n311), .A2(new_n248), .B1(G77), .B2(new_n263), .ZN(new_n312));
  OAI21_X1  g0112(.A(new_n312), .B1(G77), .B2(new_n260), .ZN(new_n313));
  INV_X1    g0113(.A(new_n313), .ZN(new_n314));
  AND3_X1   g0114(.A1(new_n303), .A2(KEYINPUT69), .A3(G190), .ZN(new_n315));
  AOI21_X1  g0115(.A(KEYINPUT69), .B1(new_n303), .B2(G190), .ZN(new_n316));
  OAI211_X1 g0116(.A(new_n305), .B(new_n314), .C1(new_n315), .C2(new_n316), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n303), .A2(new_n294), .ZN(new_n318));
  OAI211_X1 g0118(.A(new_n318), .B(new_n313), .C1(G169), .C2(new_n303), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n317), .A2(new_n319), .ZN(new_n320));
  XNOR2_X1  g0120(.A(new_n320), .B(KEYINPUT70), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n215), .A2(G1698), .ZN(new_n322));
  AND2_X1   g0122(.A1(KEYINPUT3), .A2(G33), .ZN(new_n323));
  NOR2_X1   g0123(.A1(KEYINPUT3), .A2(G33), .ZN(new_n324));
  OAI221_X1 g0124(.A(new_n322), .B1(G223), .B2(G1698), .C1(new_n323), .C2(new_n324), .ZN(new_n325));
  NAND2_X1  g0125(.A1(G33), .A2(G87), .ZN(new_n326));
  AOI21_X1  g0126(.A(new_n282), .B1(new_n325), .B2(new_n326), .ZN(new_n327));
  NOR2_X1   g0127(.A1(new_n283), .A2(new_n220), .ZN(new_n328));
  NOR3_X1   g0128(.A1(new_n327), .A2(new_n328), .A3(new_n279), .ZN(new_n329));
  INV_X1    g0129(.A(G200), .ZN(new_n330));
  OR2_X1    g0130(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  INV_X1    g0131(.A(KEYINPUT16), .ZN(new_n332));
  INV_X1    g0132(.A(G159), .ZN(new_n333));
  NOR2_X1   g0133(.A1(new_n254), .A2(new_n333), .ZN(new_n334));
  INV_X1    g0134(.A(new_n334), .ZN(new_n335));
  INV_X1    g0135(.A(KEYINPUT73), .ZN(new_n336));
  XNOR2_X1  g0136(.A(G58), .B(G68), .ZN(new_n337));
  AOI21_X1  g0137(.A(new_n336), .B1(new_n337), .B2(G20), .ZN(new_n338));
  AND2_X1   g0138(.A1(G58), .A2(G68), .ZN(new_n339));
  NOR2_X1   g0139(.A1(G58), .A2(G68), .ZN(new_n340));
  OAI211_X1 g0140(.A(new_n336), .B(G20), .C1(new_n339), .C2(new_n340), .ZN(new_n341));
  INV_X1    g0141(.A(new_n341), .ZN(new_n342));
  OAI21_X1  g0142(.A(new_n335), .B1(new_n338), .B2(new_n342), .ZN(new_n343));
  NAND3_X1  g0143(.A1(new_n268), .A2(new_n225), .A3(new_n269), .ZN(new_n344));
  INV_X1    g0144(.A(KEYINPUT7), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n344), .A2(new_n345), .ZN(new_n346));
  NAND4_X1  g0146(.A1(new_n268), .A2(KEYINPUT7), .A3(new_n225), .A4(new_n269), .ZN(new_n347));
  AOI21_X1  g0147(.A(new_n208), .B1(new_n346), .B2(new_n347), .ZN(new_n348));
  OAI21_X1  g0148(.A(new_n332), .B1(new_n343), .B2(new_n348), .ZN(new_n349));
  NOR2_X1   g0149(.A1(new_n323), .A2(new_n324), .ZN(new_n350));
  AOI21_X1  g0150(.A(KEYINPUT7), .B1(new_n350), .B2(new_n225), .ZN(new_n351));
  INV_X1    g0151(.A(new_n347), .ZN(new_n352));
  OAI21_X1  g0152(.A(G68), .B1(new_n351), .B2(new_n352), .ZN(new_n353));
  OAI21_X1  g0153(.A(G20), .B1(new_n339), .B2(new_n340), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n354), .A2(KEYINPUT73), .ZN(new_n355));
  AOI21_X1  g0155(.A(new_n334), .B1(new_n355), .B2(new_n341), .ZN(new_n356));
  NAND3_X1  g0156(.A1(new_n353), .A2(new_n356), .A3(KEYINPUT16), .ZN(new_n357));
  NAND3_X1  g0157(.A1(new_n349), .A2(new_n357), .A3(new_n248), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n329), .A2(G190), .ZN(new_n359));
  NOR2_X1   g0159(.A1(new_n306), .A2(new_n260), .ZN(new_n360));
  AOI21_X1  g0160(.A(new_n360), .B1(new_n306), .B2(new_n263), .ZN(new_n361));
  NAND4_X1  g0161(.A1(new_n331), .A2(new_n358), .A3(new_n359), .A4(new_n361), .ZN(new_n362));
  XNOR2_X1  g0162(.A(new_n362), .B(KEYINPUT17), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n358), .A2(new_n361), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n325), .A2(new_n326), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n365), .A2(new_n275), .ZN(new_n366));
  INV_X1    g0166(.A(new_n328), .ZN(new_n367));
  NAND4_X1  g0167(.A1(new_n366), .A2(new_n367), .A3(G179), .A4(new_n280), .ZN(new_n368));
  OAI21_X1  g0168(.A(new_n368), .B1(new_n329), .B2(new_n292), .ZN(new_n369));
  AOI21_X1  g0169(.A(KEYINPUT18), .B1(new_n364), .B2(new_n369), .ZN(new_n370));
  AND3_X1   g0170(.A1(new_n364), .A2(KEYINPUT18), .A3(new_n369), .ZN(new_n371));
  OAI21_X1  g0171(.A(new_n363), .B1(new_n370), .B2(new_n371), .ZN(new_n372));
  INV_X1    g0172(.A(new_n372), .ZN(new_n373));
  NAND2_X1  g0173(.A1(G33), .A2(G97), .ZN(new_n374));
  OAI21_X1  g0174(.A(new_n270), .B1(G232), .B2(new_n271), .ZN(new_n375));
  NOR2_X1   g0175(.A1(G226), .A2(G1698), .ZN(new_n376));
  OAI21_X1  g0176(.A(new_n374), .B1(new_n375), .B2(new_n376), .ZN(new_n377));
  AOI21_X1  g0177(.A(new_n279), .B1(new_n377), .B2(new_n275), .ZN(new_n378));
  NAND3_X1  g0178(.A1(new_n282), .A2(G238), .A3(new_n277), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n378), .A2(new_n379), .ZN(new_n380));
  NOR2_X1   g0180(.A1(new_n380), .A2(KEYINPUT13), .ZN(new_n381));
  INV_X1    g0181(.A(KEYINPUT13), .ZN(new_n382));
  AOI21_X1  g0182(.A(new_n382), .B1(new_n378), .B2(new_n379), .ZN(new_n383));
  OR2_X1    g0183(.A1(new_n381), .A2(new_n383), .ZN(new_n384));
  INV_X1    g0184(.A(KEYINPUT14), .ZN(new_n385));
  NAND3_X1  g0185(.A1(new_n384), .A2(new_n385), .A3(G169), .ZN(new_n386));
  NOR2_X1   g0186(.A1(new_n381), .A2(new_n383), .ZN(new_n387));
  OAI21_X1  g0187(.A(KEYINPUT14), .B1(new_n387), .B2(new_n292), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n387), .A2(G179), .ZN(new_n389));
  NAND3_X1  g0189(.A1(new_n386), .A2(new_n388), .A3(new_n389), .ZN(new_n390));
  OAI22_X1  g0190(.A1(new_n254), .A2(new_n214), .B1(new_n225), .B2(G68), .ZN(new_n391));
  NOR2_X1   g0191(.A1(new_n250), .A2(new_n216), .ZN(new_n392));
  OAI21_X1  g0192(.A(new_n248), .B1(new_n391), .B2(new_n392), .ZN(new_n393));
  XNOR2_X1  g0193(.A(new_n393), .B(KEYINPUT11), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n263), .A2(G68), .ZN(new_n395));
  OAI21_X1  g0195(.A(KEYINPUT71), .B1(new_n260), .B2(G68), .ZN(new_n396));
  XOR2_X1   g0196(.A(new_n396), .B(KEYINPUT12), .Z(new_n397));
  AND3_X1   g0197(.A1(new_n394), .A2(new_n395), .A3(new_n397), .ZN(new_n398));
  XNOR2_X1  g0198(.A(new_n398), .B(KEYINPUT72), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n390), .A2(new_n399), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n384), .A2(G200), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n387), .A2(G190), .ZN(new_n402));
  NAND3_X1  g0202(.A1(new_n401), .A2(new_n402), .A3(new_n398), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n400), .A2(new_n403), .ZN(new_n404));
  INV_X1    g0204(.A(new_n404), .ZN(new_n405));
  NAND4_X1  g0205(.A1(new_n298), .A2(new_n321), .A3(new_n373), .A4(new_n405), .ZN(new_n406));
  INV_X1    g0206(.A(new_n406), .ZN(new_n407));
  NOR2_X1   g0207(.A1(KEYINPUT83), .A2(KEYINPUT20), .ZN(new_n408));
  INV_X1    g0208(.A(G97), .ZN(new_n409));
  OAI21_X1  g0209(.A(new_n225), .B1(new_n409), .B2(G33), .ZN(new_n410));
  NAND2_X1  g0210(.A1(G33), .A2(G283), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n411), .A2(KEYINPUT75), .ZN(new_n412));
  INV_X1    g0212(.A(KEYINPUT75), .ZN(new_n413));
  NAND3_X1  g0213(.A1(new_n413), .A2(G33), .A3(G283), .ZN(new_n414));
  AOI21_X1  g0214(.A(new_n410), .B1(new_n412), .B2(new_n414), .ZN(new_n415));
  INV_X1    g0215(.A(G116), .ZN(new_n416));
  AOI22_X1  g0216(.A1(new_n247), .A2(new_n224), .B1(G20), .B2(new_n416), .ZN(new_n417));
  INV_X1    g0217(.A(new_n417), .ZN(new_n418));
  OAI21_X1  g0218(.A(new_n408), .B1(new_n415), .B2(new_n418), .ZN(new_n419));
  INV_X1    g0219(.A(new_n408), .ZN(new_n420));
  AND2_X1   g0220(.A1(new_n412), .A2(new_n414), .ZN(new_n421));
  OAI211_X1 g0221(.A(new_n417), .B(new_n420), .C1(new_n421), .C2(new_n410), .ZN(new_n422));
  NAND2_X1  g0222(.A1(KEYINPUT83), .A2(KEYINPUT20), .ZN(new_n423));
  NAND3_X1  g0223(.A1(new_n419), .A2(new_n422), .A3(new_n423), .ZN(new_n424));
  AND2_X1   g0224(.A1(new_n247), .A2(new_n224), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n259), .A2(G33), .ZN(new_n426));
  NAND3_X1  g0226(.A1(new_n425), .A2(new_n260), .A3(new_n426), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n427), .A2(G116), .ZN(new_n428));
  OAI21_X1  g0228(.A(new_n428), .B1(G116), .B2(new_n261), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n424), .A2(new_n429), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n271), .A2(G257), .ZN(new_n431));
  NAND2_X1  g0231(.A1(G264), .A2(G1698), .ZN(new_n432));
  OAI211_X1 g0232(.A(new_n431), .B(new_n432), .C1(new_n323), .C2(new_n324), .ZN(new_n433));
  INV_X1    g0233(.A(G303), .ZN(new_n434));
  NAND3_X1  g0234(.A1(new_n268), .A2(new_n434), .A3(new_n269), .ZN(new_n435));
  NAND3_X1  g0235(.A1(new_n433), .A2(new_n275), .A3(new_n435), .ZN(new_n436));
  INV_X1    g0236(.A(G45), .ZN(new_n437));
  NOR2_X1   g0237(.A1(new_n437), .A2(G1), .ZN(new_n438));
  AND2_X1   g0238(.A1(KEYINPUT5), .A2(G41), .ZN(new_n439));
  NOR2_X1   g0239(.A1(KEYINPUT5), .A2(G41), .ZN(new_n440));
  OAI21_X1  g0240(.A(new_n438), .B1(new_n439), .B2(new_n440), .ZN(new_n441));
  NAND3_X1  g0241(.A1(new_n441), .A2(G270), .A3(new_n282), .ZN(new_n442));
  OAI211_X1 g0242(.A(new_n438), .B(G274), .C1(new_n440), .C2(new_n439), .ZN(new_n443));
  NAND3_X1  g0243(.A1(new_n436), .A2(new_n442), .A3(new_n443), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n444), .A2(G169), .ZN(new_n445));
  INV_X1    g0245(.A(KEYINPUT21), .ZN(new_n446));
  NOR2_X1   g0246(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  NOR2_X1   g0247(.A1(new_n444), .A2(new_n294), .ZN(new_n448));
  OAI21_X1  g0248(.A(new_n430), .B1(new_n447), .B2(new_n448), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n444), .A2(G200), .ZN(new_n450));
  INV_X1    g0250(.A(G190), .ZN(new_n451));
  OAI21_X1  g0251(.A(new_n450), .B1(new_n451), .B2(new_n444), .ZN(new_n452));
  OR2_X1    g0252(.A1(new_n452), .A2(new_n430), .ZN(new_n453));
  AOI21_X1  g0253(.A(new_n445), .B1(new_n429), .B2(new_n424), .ZN(new_n454));
  NOR3_X1   g0254(.A1(new_n454), .A2(KEYINPUT84), .A3(KEYINPUT21), .ZN(new_n455));
  INV_X1    g0255(.A(KEYINPUT84), .ZN(new_n456));
  INV_X1    g0256(.A(new_n445), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n430), .A2(new_n457), .ZN(new_n458));
  AOI21_X1  g0258(.A(new_n456), .B1(new_n458), .B2(new_n446), .ZN(new_n459));
  OAI211_X1 g0259(.A(new_n449), .B(new_n453), .C1(new_n455), .C2(new_n459), .ZN(new_n460));
  INV_X1    g0260(.A(KEYINPUT85), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  OAI21_X1  g0262(.A(KEYINPUT84), .B1(new_n454), .B2(KEYINPUT21), .ZN(new_n463));
  NAND3_X1  g0263(.A1(new_n458), .A2(new_n456), .A3(new_n446), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  NAND4_X1  g0265(.A1(new_n465), .A2(KEYINPUT85), .A3(new_n449), .A4(new_n453), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n462), .A2(new_n466), .ZN(new_n467));
  OR2_X1    g0267(.A1(G250), .A2(G1698), .ZN(new_n468));
  OAI211_X1 g0268(.A(new_n270), .B(new_n468), .C1(G257), .C2(new_n271), .ZN(new_n469));
  NAND2_X1  g0269(.A1(G33), .A2(G294), .ZN(new_n470));
  AOI21_X1  g0270(.A(new_n282), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  AND3_X1   g0271(.A1(new_n441), .A2(G264), .A3(new_n282), .ZN(new_n472));
  NOR2_X1   g0272(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n473), .A2(new_n443), .ZN(new_n474));
  NAND3_X1  g0274(.A1(new_n474), .A2(KEYINPUT89), .A3(G169), .ZN(new_n475));
  INV_X1    g0275(.A(KEYINPUT89), .ZN(new_n476));
  INV_X1    g0276(.A(new_n443), .ZN(new_n477));
  NOR3_X1   g0277(.A1(new_n471), .A2(new_n472), .A3(new_n477), .ZN(new_n478));
  OAI21_X1  g0278(.A(new_n476), .B1(new_n478), .B2(new_n292), .ZN(new_n479));
  OAI211_X1 g0279(.A(new_n475), .B(new_n479), .C1(new_n294), .C2(new_n474), .ZN(new_n480));
  NOR2_X1   g0280(.A1(new_n225), .A2(G107), .ZN(new_n481));
  XNOR2_X1  g0281(.A(new_n481), .B(KEYINPUT23), .ZN(new_n482));
  NOR2_X1   g0282(.A1(new_n253), .A2(new_n416), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n483), .A2(new_n225), .ZN(new_n484));
  NAND3_X1  g0284(.A1(new_n270), .A2(new_n225), .A3(G87), .ZN(new_n485));
  AND2_X1   g0285(.A1(new_n485), .A2(KEYINPUT22), .ZN(new_n486));
  NOR2_X1   g0286(.A1(new_n485), .A2(KEYINPUT22), .ZN(new_n487));
  OAI211_X1 g0287(.A(new_n482), .B(new_n484), .C1(new_n486), .C2(new_n487), .ZN(new_n488));
  XNOR2_X1  g0288(.A(KEYINPUT86), .B(KEYINPUT24), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  XNOR2_X1  g0290(.A(new_n485), .B(KEYINPUT22), .ZN(new_n491));
  INV_X1    g0291(.A(new_n489), .ZN(new_n492));
  NAND4_X1  g0292(.A1(new_n491), .A2(new_n492), .A3(new_n482), .A4(new_n484), .ZN(new_n493));
  NAND3_X1  g0293(.A1(new_n490), .A2(new_n493), .A3(new_n248), .ZN(new_n494));
  INV_X1    g0294(.A(KEYINPUT74), .ZN(new_n495));
  OR2_X1    g0295(.A1(new_n427), .A2(new_n495), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n427), .A2(new_n495), .ZN(new_n497));
  AND2_X1   g0297(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n498), .A2(G107), .ZN(new_n499));
  AOI21_X1  g0299(.A(KEYINPUT25), .B1(new_n261), .B2(new_n210), .ZN(new_n500));
  XOR2_X1   g0300(.A(new_n500), .B(KEYINPUT88), .Z(new_n501));
  NAND3_X1  g0301(.A1(new_n261), .A2(KEYINPUT25), .A3(new_n210), .ZN(new_n502));
  XNOR2_X1  g0302(.A(new_n502), .B(KEYINPUT87), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n501), .A2(new_n503), .ZN(new_n504));
  NAND3_X1  g0304(.A1(new_n494), .A2(new_n499), .A3(new_n504), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n480), .A2(new_n505), .ZN(new_n506));
  INV_X1    g0306(.A(new_n506), .ZN(new_n507));
  NOR2_X1   g0307(.A1(new_n478), .A2(new_n330), .ZN(new_n508));
  NOR2_X1   g0308(.A1(new_n474), .A2(new_n451), .ZN(new_n509));
  NOR3_X1   g0309(.A1(new_n505), .A2(new_n508), .A3(new_n509), .ZN(new_n510));
  NOR2_X1   g0310(.A1(new_n507), .A2(new_n510), .ZN(new_n511));
  INV_X1    g0311(.A(KEYINPUT19), .ZN(new_n512));
  OAI21_X1  g0312(.A(new_n225), .B1(new_n374), .B2(new_n512), .ZN(new_n513));
  XNOR2_X1  g0313(.A(KEYINPUT79), .B(G87), .ZN(new_n514));
  INV_X1    g0314(.A(KEYINPUT80), .ZN(new_n515));
  NOR2_X1   g0315(.A1(G97), .A2(G107), .ZN(new_n516));
  NAND3_X1  g0316(.A1(new_n514), .A2(new_n515), .A3(new_n516), .ZN(new_n517));
  INV_X1    g0317(.A(new_n517), .ZN(new_n518));
  AOI21_X1  g0318(.A(new_n515), .B1(new_n514), .B2(new_n516), .ZN(new_n519));
  OAI21_X1  g0319(.A(new_n513), .B1(new_n518), .B2(new_n519), .ZN(new_n520));
  INV_X1    g0320(.A(KEYINPUT81), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  OAI21_X1  g0322(.A(new_n512), .B1(new_n250), .B2(new_n409), .ZN(new_n523));
  INV_X1    g0323(.A(KEYINPUT82), .ZN(new_n524));
  OR2_X1    g0324(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  OAI211_X1 g0325(.A(KEYINPUT81), .B(new_n513), .C1(new_n518), .C2(new_n519), .ZN(new_n526));
  NOR2_X1   g0326(.A1(new_n350), .A2(G20), .ZN(new_n527));
  AOI22_X1  g0327(.A1(new_n527), .A2(G68), .B1(new_n524), .B2(new_n523), .ZN(new_n528));
  NAND4_X1  g0328(.A1(new_n522), .A2(new_n525), .A3(new_n526), .A4(new_n528), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n529), .A2(new_n248), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n310), .A2(new_n261), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n498), .A2(new_n309), .ZN(new_n532));
  NAND3_X1  g0332(.A1(new_n530), .A2(new_n531), .A3(new_n532), .ZN(new_n533));
  NAND3_X1  g0333(.A1(new_n270), .A2(G238), .A3(new_n271), .ZN(new_n534));
  INV_X1    g0334(.A(new_n483), .ZN(new_n535));
  AND2_X1   g0335(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  OAI211_X1 g0336(.A(G244), .B(G1698), .C1(new_n323), .C2(new_n324), .ZN(new_n537));
  INV_X1    g0337(.A(KEYINPUT77), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  NAND4_X1  g0339(.A1(new_n270), .A2(KEYINPUT77), .A3(G244), .A4(G1698), .ZN(new_n540));
  NAND4_X1  g0340(.A1(new_n536), .A2(KEYINPUT78), .A3(new_n539), .A4(new_n540), .ZN(new_n541));
  NAND4_X1  g0341(.A1(new_n539), .A2(new_n540), .A3(new_n535), .A4(new_n534), .ZN(new_n542));
  INV_X1    g0342(.A(KEYINPUT78), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  AOI21_X1  g0344(.A(new_n282), .B1(new_n541), .B2(new_n544), .ZN(new_n545));
  OAI21_X1  g0345(.A(new_n282), .B1(G250), .B2(new_n438), .ZN(new_n546));
  AOI21_X1  g0346(.A(new_n546), .B1(new_n278), .B2(new_n438), .ZN(new_n547));
  NOR2_X1   g0347(.A1(new_n545), .A2(new_n547), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n548), .A2(new_n294), .ZN(new_n549));
  OAI21_X1  g0349(.A(new_n292), .B1(new_n545), .B2(new_n547), .ZN(new_n550));
  NAND3_X1  g0350(.A1(new_n533), .A2(new_n549), .A3(new_n550), .ZN(new_n551));
  OAI211_X1 g0351(.A(G244), .B(new_n271), .C1(new_n323), .C2(new_n324), .ZN(new_n552));
  INV_X1    g0352(.A(KEYINPUT4), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  NAND4_X1  g0354(.A1(new_n270), .A2(KEYINPUT4), .A3(G244), .A4(new_n271), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n412), .A2(new_n414), .ZN(new_n556));
  NAND3_X1  g0356(.A1(new_n270), .A2(G250), .A3(G1698), .ZN(new_n557));
  NAND4_X1  g0357(.A1(new_n554), .A2(new_n555), .A3(new_n556), .A4(new_n557), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n558), .A2(new_n275), .ZN(new_n559));
  AND2_X1   g0359(.A1(new_n441), .A2(new_n282), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n560), .A2(G257), .ZN(new_n561));
  NAND3_X1  g0361(.A1(new_n559), .A2(new_n443), .A3(new_n561), .ZN(new_n562));
  INV_X1    g0362(.A(KEYINPUT76), .ZN(new_n563));
  NOR2_X1   g0363(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  AOI22_X1  g0364(.A1(new_n558), .A2(new_n275), .B1(G257), .B2(new_n560), .ZN(new_n565));
  AOI21_X1  g0365(.A(KEYINPUT76), .B1(new_n565), .B2(new_n443), .ZN(new_n566));
  OAI21_X1  g0366(.A(G190), .B1(new_n564), .B2(new_n566), .ZN(new_n567));
  NOR2_X1   g0367(.A1(new_n260), .A2(G97), .ZN(new_n568));
  AND3_X1   g0368(.A1(new_n496), .A2(G97), .A3(new_n497), .ZN(new_n569));
  AOI21_X1  g0369(.A(new_n210), .B1(new_n346), .B2(new_n347), .ZN(new_n570));
  NAND3_X1  g0370(.A1(new_n210), .A2(KEYINPUT6), .A3(G97), .ZN(new_n571));
  NOR2_X1   g0371(.A1(new_n409), .A2(new_n210), .ZN(new_n572));
  NOR2_X1   g0372(.A1(new_n572), .A2(new_n516), .ZN(new_n573));
  OAI21_X1  g0373(.A(new_n571), .B1(new_n573), .B2(KEYINPUT6), .ZN(new_n574));
  AOI21_X1  g0374(.A(new_n570), .B1(G20), .B2(new_n574), .ZN(new_n575));
  NOR2_X1   g0375(.A1(new_n254), .A2(new_n216), .ZN(new_n576));
  INV_X1    g0376(.A(new_n576), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n575), .A2(new_n577), .ZN(new_n578));
  AOI211_X1 g0378(.A(new_n568), .B(new_n569), .C1(new_n578), .C2(new_n248), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n562), .A2(G200), .ZN(new_n580));
  NAND3_X1  g0380(.A1(new_n567), .A2(new_n579), .A3(new_n580), .ZN(new_n581));
  INV_X1    g0381(.A(new_n545), .ZN(new_n582));
  INV_X1    g0382(.A(new_n547), .ZN(new_n583));
  NAND3_X1  g0383(.A1(new_n582), .A2(G190), .A3(new_n583), .ZN(new_n584));
  AOI22_X1  g0384(.A1(new_n529), .A2(new_n248), .B1(new_n261), .B2(new_n310), .ZN(new_n585));
  OAI21_X1  g0385(.A(G200), .B1(new_n545), .B2(new_n547), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n498), .A2(G87), .ZN(new_n587));
  NAND4_X1  g0387(.A1(new_n584), .A2(new_n585), .A3(new_n586), .A4(new_n587), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n562), .A2(new_n563), .ZN(new_n589));
  NAND3_X1  g0389(.A1(new_n565), .A2(KEYINPUT76), .A3(new_n443), .ZN(new_n590));
  NAND3_X1  g0390(.A1(new_n589), .A2(new_n292), .A3(new_n590), .ZN(new_n591));
  NAND3_X1  g0391(.A1(new_n565), .A2(new_n294), .A3(new_n443), .ZN(new_n592));
  INV_X1    g0392(.A(new_n568), .ZN(new_n593));
  INV_X1    g0393(.A(new_n569), .ZN(new_n594));
  AOI211_X1 g0394(.A(new_n576), .B(new_n570), .C1(G20), .C2(new_n574), .ZN(new_n595));
  OAI211_X1 g0395(.A(new_n593), .B(new_n594), .C1(new_n595), .C2(new_n425), .ZN(new_n596));
  NAND3_X1  g0396(.A1(new_n591), .A2(new_n592), .A3(new_n596), .ZN(new_n597));
  AND4_X1   g0397(.A1(new_n551), .A2(new_n581), .A3(new_n588), .A4(new_n597), .ZN(new_n598));
  AND4_X1   g0398(.A1(new_n407), .A2(new_n467), .A3(new_n511), .A4(new_n598), .ZN(G372));
  AND3_X1   g0399(.A1(new_n584), .A2(new_n585), .A3(new_n587), .ZN(new_n600));
  INV_X1    g0400(.A(KEYINPUT90), .ZN(new_n601));
  NOR2_X1   g0401(.A1(new_n545), .A2(new_n601), .ZN(new_n602));
  AOI211_X1 g0402(.A(KEYINPUT90), .B(new_n282), .C1(new_n541), .C2(new_n544), .ZN(new_n603));
  OAI21_X1  g0403(.A(new_n583), .B1(new_n602), .B2(new_n603), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n604), .A2(G200), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n604), .A2(new_n292), .ZN(new_n606));
  AOI22_X1  g0406(.A1(new_n585), .A2(new_n532), .B1(new_n548), .B2(new_n294), .ZN(new_n607));
  AOI22_X1  g0407(.A1(new_n600), .A2(new_n605), .B1(new_n606), .B2(new_n607), .ZN(new_n608));
  INV_X1    g0408(.A(KEYINPUT26), .ZN(new_n609));
  INV_X1    g0409(.A(new_n597), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n610), .A2(KEYINPUT91), .ZN(new_n611));
  INV_X1    g0411(.A(KEYINPUT91), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n597), .A2(new_n612), .ZN(new_n613));
  NAND4_X1  g0413(.A1(new_n608), .A2(new_n609), .A3(new_n611), .A4(new_n613), .ZN(new_n614));
  AOI21_X1  g0414(.A(new_n510), .B1(new_n600), .B2(new_n605), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n581), .A2(new_n597), .ZN(new_n616));
  INV_X1    g0416(.A(new_n616), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n465), .A2(new_n449), .ZN(new_n618));
  INV_X1    g0418(.A(new_n618), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n619), .A2(new_n506), .ZN(new_n620));
  NAND3_X1  g0420(.A1(new_n615), .A2(new_n617), .A3(new_n620), .ZN(new_n621));
  NAND3_X1  g0421(.A1(new_n610), .A2(new_n551), .A3(new_n588), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n622), .A2(KEYINPUT26), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n606), .A2(new_n607), .ZN(new_n624));
  NAND4_X1  g0424(.A1(new_n614), .A2(new_n621), .A3(new_n623), .A4(new_n624), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n407), .A2(new_n625), .ZN(new_n626));
  NOR2_X1   g0426(.A1(new_n371), .A2(new_n370), .ZN(new_n627));
  INV_X1    g0427(.A(new_n403), .ZN(new_n628));
  OAI21_X1  g0428(.A(new_n400), .B1(new_n319), .B2(new_n628), .ZN(new_n629));
  AOI21_X1  g0429(.A(new_n627), .B1(new_n629), .B2(new_n363), .ZN(new_n630));
  INV_X1    g0430(.A(new_n291), .ZN(new_n631));
  OAI21_X1  g0431(.A(new_n296), .B1(new_n630), .B2(new_n631), .ZN(new_n632));
  INV_X1    g0432(.A(new_n632), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n626), .A2(new_n633), .ZN(G369));
  INV_X1    g0434(.A(G13), .ZN(new_n635));
  NOR2_X1   g0435(.A1(new_n635), .A2(G20), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n636), .A2(new_n259), .ZN(new_n637));
  OR2_X1    g0437(.A1(new_n637), .A2(KEYINPUT27), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n637), .A2(KEYINPUT27), .ZN(new_n639));
  AND3_X1   g0439(.A1(new_n638), .A2(G213), .A3(new_n639), .ZN(new_n640));
  INV_X1    g0440(.A(new_n640), .ZN(new_n641));
  INV_X1    g0441(.A(G343), .ZN(new_n642));
  NOR2_X1   g0442(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n643), .A2(new_n430), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n467), .A2(new_n644), .ZN(new_n645));
  OAI21_X1  g0445(.A(new_n645), .B1(new_n619), .B2(new_n644), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n646), .A2(G330), .ZN(new_n647));
  INV_X1    g0447(.A(new_n647), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n505), .A2(new_n643), .ZN(new_n649));
  AOI22_X1  g0449(.A1(new_n511), .A2(new_n649), .B1(new_n507), .B2(new_n643), .ZN(new_n650));
  INV_X1    g0450(.A(new_n650), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n648), .A2(new_n651), .ZN(new_n652));
  INV_X1    g0452(.A(new_n643), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n618), .A2(new_n653), .ZN(new_n654));
  NOR3_X1   g0454(.A1(new_n654), .A2(new_n507), .A3(new_n510), .ZN(new_n655));
  AOI21_X1  g0455(.A(new_n655), .B1(new_n507), .B2(new_n653), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n652), .A2(new_n656), .ZN(G399));
  NOR2_X1   g0457(.A1(new_n518), .A2(new_n519), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n658), .A2(new_n416), .ZN(new_n659));
  INV_X1    g0459(.A(new_n659), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n204), .A2(new_n281), .ZN(new_n661));
  NAND3_X1  g0461(.A1(new_n660), .A2(G1), .A3(new_n661), .ZN(new_n662));
  OAI21_X1  g0462(.A(new_n662), .B1(new_n227), .B2(new_n661), .ZN(new_n663));
  XNOR2_X1  g0463(.A(new_n663), .B(KEYINPUT28), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n625), .A2(new_n653), .ZN(new_n665));
  INV_X1    g0465(.A(KEYINPUT29), .ZN(new_n666));
  AOI21_X1  g0466(.A(KEYINPUT94), .B1(new_n665), .B2(new_n666), .ZN(new_n667));
  NOR2_X1   g0467(.A1(new_n622), .A2(KEYINPUT26), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n600), .A2(new_n605), .ZN(new_n669));
  NAND4_X1  g0469(.A1(new_n611), .A2(new_n669), .A3(new_n624), .A4(new_n613), .ZN(new_n670));
  AOI21_X1  g0470(.A(new_n668), .B1(new_n670), .B2(KEYINPUT26), .ZN(new_n671));
  AOI21_X1  g0471(.A(new_n616), .B1(new_n619), .B2(new_n506), .ZN(new_n672));
  AOI22_X1  g0472(.A1(new_n672), .A2(new_n615), .B1(new_n607), .B2(new_n606), .ZN(new_n673));
  AOI21_X1  g0473(.A(new_n643), .B1(new_n671), .B2(new_n673), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n674), .A2(KEYINPUT29), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n667), .A2(new_n675), .ZN(new_n676));
  NAND3_X1  g0476(.A1(new_n674), .A2(KEYINPUT94), .A3(KEYINPUT29), .ZN(new_n677));
  AND2_X1   g0477(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  NAND4_X1  g0478(.A1(new_n598), .A2(new_n467), .A3(new_n511), .A4(new_n653), .ZN(new_n679));
  NAND3_X1  g0479(.A1(new_n562), .A2(new_n474), .A3(KEYINPUT93), .ZN(new_n680));
  INV_X1    g0480(.A(KEYINPUT93), .ZN(new_n681));
  OAI211_X1 g0481(.A(new_n681), .B(new_n443), .C1(new_n565), .C2(new_n473), .ZN(new_n682));
  AOI21_X1  g0482(.A(G179), .B1(new_n680), .B2(new_n682), .ZN(new_n683));
  NAND3_X1  g0483(.A1(new_n604), .A2(new_n444), .A3(new_n683), .ZN(new_n684));
  INV_X1    g0484(.A(KEYINPUT30), .ZN(new_n685));
  OAI21_X1  g0485(.A(new_n448), .B1(new_n564), .B2(new_n566), .ZN(new_n686));
  NAND3_X1  g0486(.A1(new_n582), .A2(new_n473), .A3(new_n583), .ZN(new_n687));
  OAI21_X1  g0487(.A(new_n685), .B1(new_n686), .B2(new_n687), .ZN(new_n688));
  NOR4_X1   g0488(.A1(new_n545), .A2(new_n472), .A3(new_n471), .A4(new_n547), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n589), .A2(new_n590), .ZN(new_n690));
  NAND4_X1  g0490(.A1(new_n689), .A2(new_n690), .A3(KEYINPUT30), .A4(new_n448), .ZN(new_n691));
  NAND3_X1  g0491(.A1(new_n684), .A2(new_n688), .A3(new_n691), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n692), .A2(new_n643), .ZN(new_n693));
  INV_X1    g0493(.A(KEYINPUT31), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  XNOR2_X1  g0495(.A(KEYINPUT92), .B(KEYINPUT31), .ZN(new_n696));
  INV_X1    g0496(.A(new_n696), .ZN(new_n697));
  OAI211_X1 g0497(.A(new_n679), .B(new_n695), .C1(new_n693), .C2(new_n697), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n698), .A2(G330), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n678), .A2(new_n699), .ZN(new_n700));
  INV_X1    g0500(.A(new_n700), .ZN(new_n701));
  OAI21_X1  g0501(.A(new_n664), .B1(new_n701), .B2(G1), .ZN(G364));
  NAND2_X1  g0502(.A1(new_n636), .A2(G45), .ZN(new_n703));
  NAND3_X1  g0503(.A1(new_n661), .A2(G1), .A3(new_n703), .ZN(new_n704));
  INV_X1    g0504(.A(new_n704), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n350), .A2(new_n204), .ZN(new_n706));
  XOR2_X1   g0506(.A(new_n706), .B(KEYINPUT96), .Z(new_n707));
  OAI21_X1  g0507(.A(new_n707), .B1(G45), .B2(new_n227), .ZN(new_n708));
  XNOR2_X1  g0508(.A(new_n708), .B(KEYINPUT97), .ZN(new_n709));
  OAI21_X1  g0509(.A(new_n709), .B1(new_n437), .B2(new_n242), .ZN(new_n710));
  NAND3_X1  g0510(.A1(new_n270), .A2(G355), .A3(new_n204), .ZN(new_n711));
  OAI21_X1  g0511(.A(new_n711), .B1(G116), .B2(new_n204), .ZN(new_n712));
  XNOR2_X1  g0512(.A(new_n712), .B(KEYINPUT95), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n710), .A2(new_n713), .ZN(new_n714));
  NOR3_X1   g0514(.A1(G13), .A2(G20), .A3(G33), .ZN(new_n715));
  XOR2_X1   g0515(.A(new_n715), .B(KEYINPUT98), .Z(new_n716));
  INV_X1    g0516(.A(new_n716), .ZN(new_n717));
  AOI21_X1  g0517(.A(new_n224), .B1(G20), .B2(new_n292), .ZN(new_n718));
  NOR2_X1   g0518(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  NOR2_X1   g0519(.A1(new_n225), .A2(new_n451), .ZN(new_n720));
  NOR2_X1   g0520(.A1(new_n330), .A2(G179), .ZN(new_n721));
  NAND2_X1  g0521(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  NOR2_X1   g0522(.A1(new_n225), .A2(G190), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n723), .A2(new_n721), .ZN(new_n724));
  OAI22_X1  g0524(.A1(new_n722), .A2(new_n514), .B1(new_n724), .B2(new_n210), .ZN(new_n725));
  NOR2_X1   g0525(.A1(new_n294), .A2(G200), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n720), .A2(new_n726), .ZN(new_n727));
  INV_X1    g0527(.A(new_n727), .ZN(new_n728));
  AOI211_X1 g0528(.A(new_n350), .B(new_n725), .C1(G58), .C2(new_n728), .ZN(new_n729));
  NOR2_X1   g0529(.A1(G179), .A2(G200), .ZN(new_n730));
  AOI21_X1  g0530(.A(new_n225), .B1(new_n730), .B2(G190), .ZN(new_n731));
  INV_X1    g0531(.A(new_n731), .ZN(new_n732));
  NAND2_X1  g0532(.A1(new_n732), .A2(G97), .ZN(new_n733));
  NAND2_X1  g0533(.A1(new_n723), .A2(new_n730), .ZN(new_n734));
  NOR2_X1   g0534(.A1(new_n734), .A2(new_n333), .ZN(new_n735));
  XNOR2_X1  g0535(.A(new_n735), .B(KEYINPUT32), .ZN(new_n736));
  NOR2_X1   g0536(.A1(new_n294), .A2(new_n330), .ZN(new_n737));
  NAND2_X1  g0537(.A1(new_n737), .A2(new_n723), .ZN(new_n738));
  NAND2_X1  g0538(.A1(new_n723), .A2(new_n726), .ZN(new_n739));
  OAI22_X1  g0539(.A1(new_n738), .A2(new_n208), .B1(new_n739), .B2(new_n216), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n720), .A2(new_n737), .ZN(new_n741));
  INV_X1    g0541(.A(new_n741), .ZN(new_n742));
  AOI21_X1  g0542(.A(new_n740), .B1(G50), .B2(new_n742), .ZN(new_n743));
  NAND4_X1  g0543(.A1(new_n729), .A2(new_n733), .A3(new_n736), .A4(new_n743), .ZN(new_n744));
  INV_X1    g0544(.A(new_n738), .ZN(new_n745));
  INV_X1    g0545(.A(G317), .ZN(new_n746));
  NAND2_X1  g0546(.A1(new_n746), .A2(KEYINPUT33), .ZN(new_n747));
  OR2_X1    g0547(.A1(new_n746), .A2(KEYINPUT33), .ZN(new_n748));
  NAND3_X1  g0548(.A1(new_n745), .A2(new_n747), .A3(new_n748), .ZN(new_n749));
  NAND2_X1  g0549(.A1(new_n742), .A2(G326), .ZN(new_n750));
  INV_X1    g0550(.A(new_n734), .ZN(new_n751));
  NAND2_X1  g0551(.A1(new_n751), .A2(G329), .ZN(new_n752));
  INV_X1    g0552(.A(new_n724), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n753), .A2(G283), .ZN(new_n754));
  NAND4_X1  g0554(.A1(new_n749), .A2(new_n750), .A3(new_n752), .A4(new_n754), .ZN(new_n755));
  AOI21_X1  g0555(.A(new_n755), .B1(G294), .B2(new_n732), .ZN(new_n756));
  AOI21_X1  g0556(.A(new_n270), .B1(new_n728), .B2(G322), .ZN(new_n757));
  OAI211_X1 g0557(.A(new_n756), .B(new_n757), .C1(new_n434), .C2(new_n722), .ZN(new_n758));
  INV_X1    g0558(.A(G311), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n739), .A2(new_n759), .ZN(new_n760));
  OAI21_X1  g0560(.A(new_n744), .B1(new_n758), .B2(new_n760), .ZN(new_n761));
  AOI22_X1  g0561(.A1(new_n714), .A2(new_n719), .B1(new_n718), .B2(new_n761), .ZN(new_n762));
  OAI211_X1 g0562(.A(new_n705), .B(new_n762), .C1(new_n646), .C2(new_n716), .ZN(new_n763));
  NAND2_X1  g0563(.A1(new_n647), .A2(new_n704), .ZN(new_n764));
  NOR2_X1   g0564(.A1(new_n646), .A2(G330), .ZN(new_n765));
  OAI21_X1  g0565(.A(new_n763), .B1(new_n764), .B2(new_n765), .ZN(G396));
  OAI21_X1  g0566(.A(new_n317), .B1(new_n314), .B2(new_n653), .ZN(new_n767));
  NAND2_X1  g0567(.A1(new_n767), .A2(new_n319), .ZN(new_n768));
  NOR2_X1   g0568(.A1(new_n319), .A2(new_n643), .ZN(new_n769));
  INV_X1    g0569(.A(new_n769), .ZN(new_n770));
  NAND2_X1  g0570(.A1(new_n768), .A2(new_n770), .ZN(new_n771));
  NAND2_X1  g0571(.A1(new_n665), .A2(new_n771), .ZN(new_n772));
  AOI21_X1  g0572(.A(new_n769), .B1(new_n767), .B2(new_n319), .ZN(new_n773));
  NAND3_X1  g0573(.A1(new_n625), .A2(new_n653), .A3(new_n773), .ZN(new_n774));
  NAND2_X1  g0574(.A1(new_n772), .A2(new_n774), .ZN(new_n775));
  INV_X1    g0575(.A(new_n699), .ZN(new_n776));
  XNOR2_X1  g0576(.A(new_n775), .B(new_n776), .ZN(new_n777));
  NAND2_X1  g0577(.A1(new_n777), .A2(new_n704), .ZN(new_n778));
  INV_X1    g0578(.A(new_n739), .ZN(new_n779));
  AOI22_X1  g0579(.A1(G143), .A2(new_n728), .B1(new_n779), .B2(G159), .ZN(new_n780));
  INV_X1    g0580(.A(G137), .ZN(new_n781));
  OAI221_X1 g0581(.A(new_n780), .B1(new_n781), .B2(new_n741), .C1(new_n255), .C2(new_n738), .ZN(new_n782));
  XOR2_X1   g0582(.A(new_n782), .B(KEYINPUT34), .Z(new_n783));
  INV_X1    g0583(.A(new_n722), .ZN(new_n784));
  AOI21_X1  g0584(.A(new_n783), .B1(G50), .B2(new_n784), .ZN(new_n785));
  NAND2_X1  g0585(.A1(new_n732), .A2(G58), .ZN(new_n786));
  NAND2_X1  g0586(.A1(new_n753), .A2(G68), .ZN(new_n787));
  NAND3_X1  g0587(.A1(new_n785), .A2(new_n786), .A3(new_n787), .ZN(new_n788));
  AOI211_X1 g0588(.A(new_n350), .B(new_n788), .C1(G132), .C2(new_n751), .ZN(new_n789));
  INV_X1    g0589(.A(G87), .ZN(new_n790));
  OAI22_X1  g0590(.A1(new_n790), .A2(new_n724), .B1(new_n739), .B2(new_n416), .ZN(new_n791));
  AOI211_X1 g0591(.A(new_n270), .B(new_n791), .C1(G294), .C2(new_n728), .ZN(new_n792));
  OAI221_X1 g0592(.A(new_n733), .B1(new_n210), .B2(new_n722), .C1(new_n759), .C2(new_n734), .ZN(new_n793));
  INV_X1    g0593(.A(new_n793), .ZN(new_n794));
  INV_X1    g0594(.A(G283), .ZN(new_n795));
  OAI211_X1 g0595(.A(new_n792), .B(new_n794), .C1(new_n795), .C2(new_n738), .ZN(new_n796));
  AOI21_X1  g0596(.A(new_n796), .B1(G303), .B2(new_n742), .ZN(new_n797));
  OAI21_X1  g0597(.A(new_n718), .B1(new_n789), .B2(new_n797), .ZN(new_n798));
  NOR2_X1   g0598(.A1(G13), .A2(G33), .ZN(new_n799));
  NOR2_X1   g0599(.A1(new_n718), .A2(new_n799), .ZN(new_n800));
  NAND2_X1  g0600(.A1(new_n800), .A2(new_n216), .ZN(new_n801));
  NAND2_X1  g0601(.A1(new_n771), .A2(new_n799), .ZN(new_n802));
  NAND4_X1  g0602(.A1(new_n798), .A2(new_n705), .A3(new_n801), .A4(new_n802), .ZN(new_n803));
  NAND2_X1  g0603(.A1(new_n778), .A2(new_n803), .ZN(G384));
  NOR2_X1   g0604(.A1(new_n678), .A2(new_n406), .ZN(new_n805));
  NOR2_X1   g0605(.A1(new_n805), .A2(new_n632), .ZN(new_n806));
  INV_X1    g0606(.A(KEYINPUT38), .ZN(new_n807));
  AND3_X1   g0607(.A1(new_n349), .A2(new_n357), .A3(new_n248), .ZN(new_n808));
  INV_X1    g0608(.A(new_n361), .ZN(new_n809));
  OAI22_X1  g0609(.A1(new_n808), .A2(new_n809), .B1(new_n369), .B2(new_n640), .ZN(new_n810));
  INV_X1    g0610(.A(KEYINPUT37), .ZN(new_n811));
  NAND3_X1  g0611(.A1(new_n810), .A2(new_n811), .A3(new_n362), .ZN(new_n812));
  INV_X1    g0612(.A(KEYINPUT101), .ZN(new_n813));
  NAND2_X1  g0613(.A1(new_n812), .A2(new_n813), .ZN(new_n814));
  NAND4_X1  g0614(.A1(new_n810), .A2(KEYINPUT101), .A3(new_n811), .A4(new_n362), .ZN(new_n815));
  AND2_X1   g0615(.A1(new_n814), .A2(new_n815), .ZN(new_n816));
  AOI21_X1  g0616(.A(KEYINPUT16), .B1(new_n353), .B2(new_n356), .ZN(new_n817));
  OAI21_X1  g0617(.A(KEYINPUT99), .B1(new_n817), .B2(new_n425), .ZN(new_n818));
  INV_X1    g0618(.A(KEYINPUT99), .ZN(new_n819));
  NAND3_X1  g0619(.A1(new_n349), .A2(new_n819), .A3(new_n248), .ZN(new_n820));
  NAND3_X1  g0620(.A1(new_n818), .A2(new_n820), .A3(new_n357), .ZN(new_n821));
  NAND2_X1  g0621(.A1(new_n821), .A2(new_n361), .ZN(new_n822));
  NAND2_X1  g0622(.A1(new_n822), .A2(KEYINPUT100), .ZN(new_n823));
  INV_X1    g0623(.A(KEYINPUT100), .ZN(new_n824));
  NAND3_X1  g0624(.A1(new_n821), .A2(new_n824), .A3(new_n361), .ZN(new_n825));
  NAND3_X1  g0625(.A1(new_n823), .A2(new_n369), .A3(new_n825), .ZN(new_n826));
  NAND3_X1  g0626(.A1(new_n823), .A2(new_n640), .A3(new_n825), .ZN(new_n827));
  NAND3_X1  g0627(.A1(new_n826), .A2(new_n827), .A3(new_n362), .ZN(new_n828));
  AOI21_X1  g0628(.A(new_n816), .B1(KEYINPUT37), .B2(new_n828), .ZN(new_n829));
  AND3_X1   g0629(.A1(new_n821), .A2(new_n824), .A3(new_n361), .ZN(new_n830));
  AOI21_X1  g0630(.A(new_n824), .B1(new_n821), .B2(new_n361), .ZN(new_n831));
  NOR2_X1   g0631(.A1(new_n830), .A2(new_n831), .ZN(new_n832));
  NAND3_X1  g0632(.A1(new_n372), .A2(new_n640), .A3(new_n832), .ZN(new_n833));
  INV_X1    g0633(.A(new_n833), .ZN(new_n834));
  OAI21_X1  g0634(.A(new_n807), .B1(new_n829), .B2(new_n834), .ZN(new_n835));
  INV_X1    g0635(.A(new_n362), .ZN(new_n836));
  AOI21_X1  g0636(.A(new_n836), .B1(new_n832), .B2(new_n640), .ZN(new_n837));
  AOI21_X1  g0637(.A(new_n811), .B1(new_n837), .B2(new_n826), .ZN(new_n838));
  OAI211_X1 g0638(.A(KEYINPUT38), .B(new_n833), .C1(new_n838), .C2(new_n816), .ZN(new_n839));
  NAND2_X1  g0639(.A1(new_n835), .A2(new_n839), .ZN(new_n840));
  INV_X1    g0640(.A(KEYINPUT104), .ZN(new_n841));
  NAND2_X1  g0641(.A1(new_n814), .A2(new_n815), .ZN(new_n842));
  INV_X1    g0642(.A(new_n810), .ZN(new_n843));
  OAI21_X1  g0643(.A(KEYINPUT37), .B1(new_n843), .B2(new_n836), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n842), .A2(new_n844), .ZN(new_n845));
  INV_X1    g0645(.A(KEYINPUT103), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  NAND3_X1  g0647(.A1(new_n372), .A2(new_n364), .A3(new_n640), .ZN(new_n848));
  NAND3_X1  g0648(.A1(new_n842), .A2(KEYINPUT103), .A3(new_n844), .ZN(new_n849));
  NAND3_X1  g0649(.A1(new_n847), .A2(new_n848), .A3(new_n849), .ZN(new_n850));
  XNOR2_X1  g0650(.A(KEYINPUT102), .B(KEYINPUT38), .ZN(new_n851));
  AOI21_X1  g0651(.A(new_n841), .B1(new_n850), .B2(new_n851), .ZN(new_n852));
  OAI21_X1  g0652(.A(KEYINPUT39), .B1(new_n840), .B2(new_n852), .ZN(new_n853));
  NAND2_X1  g0653(.A1(new_n850), .A2(new_n851), .ZN(new_n854));
  INV_X1    g0654(.A(KEYINPUT39), .ZN(new_n855));
  NAND4_X1  g0655(.A1(new_n854), .A2(new_n841), .A3(new_n855), .A4(new_n839), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n853), .A2(new_n856), .ZN(new_n857));
  NOR2_X1   g0657(.A1(new_n400), .A2(new_n643), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n399), .A2(new_n643), .ZN(new_n860));
  NAND3_X1  g0660(.A1(new_n400), .A2(new_n403), .A3(new_n860), .ZN(new_n861));
  OAI211_X1 g0661(.A(new_n399), .B(new_n643), .C1(new_n628), .C2(new_n390), .ZN(new_n862));
  AND2_X1   g0662(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  AOI21_X1  g0663(.A(new_n863), .B1(new_n774), .B2(new_n770), .ZN(new_n864));
  AOI22_X1  g0664(.A1(new_n864), .A2(new_n840), .B1(new_n627), .B2(new_n641), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n859), .A2(new_n865), .ZN(new_n866));
  XNOR2_X1  g0666(.A(new_n806), .B(new_n866), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n854), .A2(new_n839), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n868), .A2(KEYINPUT40), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n861), .A2(new_n862), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n870), .A2(new_n773), .ZN(new_n871));
  INV_X1    g0671(.A(new_n871), .ZN(new_n872));
  INV_X1    g0672(.A(KEYINPUT105), .ZN(new_n873));
  AOI21_X1  g0673(.A(new_n696), .B1(new_n692), .B2(new_n643), .ZN(new_n874));
  AND2_X1   g0674(.A1(new_n692), .A2(new_n643), .ZN(new_n875));
  AOI21_X1  g0675(.A(new_n874), .B1(KEYINPUT31), .B2(new_n875), .ZN(new_n876));
  AOI21_X1  g0676(.A(new_n873), .B1(new_n876), .B2(new_n679), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n693), .A2(new_n697), .ZN(new_n878));
  NAND3_X1  g0678(.A1(new_n692), .A2(KEYINPUT31), .A3(new_n643), .ZN(new_n879));
  NAND4_X1  g0679(.A1(new_n679), .A2(new_n878), .A3(new_n873), .A4(new_n879), .ZN(new_n880));
  INV_X1    g0680(.A(new_n880), .ZN(new_n881));
  OAI21_X1  g0681(.A(new_n872), .B1(new_n877), .B2(new_n881), .ZN(new_n882));
  OAI21_X1  g0682(.A(KEYINPUT106), .B1(new_n869), .B2(new_n882), .ZN(new_n883));
  INV_X1    g0683(.A(KEYINPUT40), .ZN(new_n884));
  AOI21_X1  g0684(.A(new_n884), .B1(new_n854), .B2(new_n839), .ZN(new_n885));
  NAND3_X1  g0685(.A1(new_n679), .A2(new_n878), .A3(new_n879), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n886), .A2(KEYINPUT105), .ZN(new_n887));
  AOI21_X1  g0687(.A(new_n871), .B1(new_n887), .B2(new_n880), .ZN(new_n888));
  INV_X1    g0688(.A(KEYINPUT106), .ZN(new_n889));
  NAND3_X1  g0689(.A1(new_n885), .A2(new_n888), .A3(new_n889), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n883), .A2(new_n890), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n887), .A2(new_n880), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n888), .A2(new_n840), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n893), .A2(new_n884), .ZN(new_n894));
  NAND4_X1  g0694(.A1(new_n891), .A2(new_n407), .A3(new_n892), .A4(new_n894), .ZN(new_n895));
  AND3_X1   g0695(.A1(new_n885), .A2(new_n888), .A3(new_n889), .ZN(new_n896));
  AOI21_X1  g0696(.A(new_n889), .B1(new_n885), .B2(new_n888), .ZN(new_n897));
  OAI211_X1 g0697(.A(new_n894), .B(G330), .C1(new_n896), .C2(new_n897), .ZN(new_n898));
  INV_X1    g0698(.A(new_n898), .ZN(new_n899));
  INV_X1    g0699(.A(G330), .ZN(new_n900));
  AOI21_X1  g0700(.A(new_n900), .B1(new_n887), .B2(new_n880), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n407), .A2(new_n901), .ZN(new_n902));
  INV_X1    g0702(.A(new_n902), .ZN(new_n903));
  OAI21_X1  g0703(.A(new_n895), .B1(new_n899), .B2(new_n903), .ZN(new_n904));
  XNOR2_X1  g0704(.A(new_n867), .B(new_n904), .ZN(new_n905));
  OAI21_X1  g0705(.A(new_n905), .B1(new_n259), .B2(new_n636), .ZN(new_n906));
  AOI21_X1  g0706(.A(new_n416), .B1(new_n574), .B2(KEYINPUT35), .ZN(new_n907));
  OAI211_X1 g0707(.A(new_n907), .B(new_n226), .C1(KEYINPUT35), .C2(new_n574), .ZN(new_n908));
  XNOR2_X1  g0708(.A(new_n908), .B(KEYINPUT36), .ZN(new_n909));
  OAI21_X1  g0709(.A(G77), .B1(new_n219), .B2(new_n208), .ZN(new_n910));
  OAI22_X1  g0710(.A1(new_n910), .A2(new_n227), .B1(G50), .B2(new_n208), .ZN(new_n911));
  NAND3_X1  g0711(.A1(new_n911), .A2(G1), .A3(new_n635), .ZN(new_n912));
  NAND3_X1  g0712(.A1(new_n906), .A2(new_n909), .A3(new_n912), .ZN(G367));
  NAND2_X1  g0713(.A1(new_n672), .A2(new_n655), .ZN(new_n914));
  XOR2_X1   g0714(.A(new_n914), .B(KEYINPUT42), .Z(new_n915));
  AOI21_X1  g0715(.A(new_n610), .B1(new_n507), .B2(new_n581), .ZN(new_n916));
  OR2_X1    g0716(.A1(new_n916), .A2(new_n643), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n585), .A2(new_n587), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n918), .A2(new_n643), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n608), .A2(new_n919), .ZN(new_n920));
  OR2_X1    g0720(.A1(new_n624), .A2(new_n919), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  AOI22_X1  g0722(.A1(new_n915), .A2(new_n917), .B1(KEYINPUT43), .B2(new_n922), .ZN(new_n923));
  NOR2_X1   g0723(.A1(new_n922), .A2(KEYINPUT43), .ZN(new_n924));
  XNOR2_X1  g0724(.A(new_n923), .B(new_n924), .ZN(new_n925));
  INV_X1    g0725(.A(new_n652), .ZN(new_n926));
  OAI21_X1  g0726(.A(new_n617), .B1(new_n579), .B2(new_n653), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n610), .A2(new_n643), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n926), .A2(new_n929), .ZN(new_n930));
  XNOR2_X1  g0730(.A(new_n925), .B(new_n930), .ZN(new_n931));
  XOR2_X1   g0731(.A(new_n661), .B(KEYINPUT41), .Z(new_n932));
  INV_X1    g0732(.A(new_n932), .ZN(new_n933));
  AOI21_X1  g0733(.A(new_n655), .B1(new_n650), .B2(new_n654), .ZN(new_n934));
  XOR2_X1   g0734(.A(new_n647), .B(new_n934), .Z(new_n935));
  INV_X1    g0735(.A(new_n935), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n701), .A2(new_n936), .ZN(new_n937));
  INV_X1    g0737(.A(KEYINPUT108), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n656), .A2(new_n929), .ZN(new_n940));
  XNOR2_X1  g0740(.A(new_n940), .B(KEYINPUT107), .ZN(new_n941));
  XNOR2_X1  g0741(.A(new_n941), .B(KEYINPUT45), .ZN(new_n942));
  NOR2_X1   g0742(.A1(new_n656), .A2(new_n929), .ZN(new_n943));
  XNOR2_X1  g0743(.A(new_n943), .B(KEYINPUT44), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n942), .A2(new_n944), .ZN(new_n945));
  INV_X1    g0745(.A(KEYINPUT109), .ZN(new_n946));
  NAND3_X1  g0746(.A1(new_n945), .A2(new_n946), .A3(new_n652), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n652), .A2(new_n946), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n926), .A2(KEYINPUT109), .ZN(new_n949));
  NAND4_X1  g0749(.A1(new_n942), .A2(new_n948), .A3(new_n949), .A4(new_n944), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n947), .A2(new_n950), .ZN(new_n951));
  NOR2_X1   g0751(.A1(new_n700), .A2(new_n935), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n952), .A2(KEYINPUT108), .ZN(new_n953));
  NAND3_X1  g0753(.A1(new_n939), .A2(new_n951), .A3(new_n953), .ZN(new_n954));
  AOI21_X1  g0754(.A(new_n933), .B1(new_n954), .B2(new_n701), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n703), .A2(G1), .ZN(new_n956));
  OAI21_X1  g0756(.A(new_n931), .B1(new_n955), .B2(new_n956), .ZN(new_n957));
  NAND3_X1  g0757(.A1(new_n920), .A2(new_n717), .A3(new_n921), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n753), .A2(G97), .ZN(new_n959));
  OAI221_X1 g0759(.A(new_n959), .B1(new_n434), .B2(new_n727), .C1(new_n746), .C2(new_n734), .ZN(new_n960));
  AOI211_X1 g0760(.A(new_n270), .B(new_n960), .C1(G107), .C2(new_n732), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n742), .A2(G311), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n784), .A2(G116), .ZN(new_n963));
  XNOR2_X1  g0763(.A(new_n963), .B(KEYINPUT46), .ZN(new_n964));
  AOI22_X1  g0764(.A1(G294), .A2(new_n745), .B1(new_n779), .B2(G283), .ZN(new_n965));
  NAND4_X1  g0765(.A1(new_n961), .A2(new_n962), .A3(new_n964), .A4(new_n965), .ZN(new_n966));
  NOR2_X1   g0766(.A1(new_n738), .A2(new_n333), .ZN(new_n967));
  NOR2_X1   g0767(.A1(new_n722), .A2(new_n219), .ZN(new_n968));
  OAI22_X1  g0768(.A1(new_n739), .A2(new_n214), .B1(new_n734), .B2(new_n781), .ZN(new_n969));
  AOI211_X1 g0769(.A(new_n968), .B(new_n969), .C1(G143), .C2(new_n742), .ZN(new_n970));
  NOR2_X1   g0770(.A1(new_n731), .A2(new_n208), .ZN(new_n971));
  INV_X1    g0771(.A(new_n971), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n728), .A2(G150), .ZN(new_n973));
  OAI21_X1  g0773(.A(new_n270), .B1(new_n724), .B2(new_n216), .ZN(new_n974));
  XNOR2_X1  g0774(.A(new_n974), .B(KEYINPUT110), .ZN(new_n975));
  NAND4_X1  g0775(.A1(new_n970), .A2(new_n972), .A3(new_n973), .A4(new_n975), .ZN(new_n976));
  OAI21_X1  g0776(.A(new_n966), .B1(new_n967), .B2(new_n976), .ZN(new_n977));
  XNOR2_X1  g0777(.A(new_n977), .B(KEYINPUT47), .ZN(new_n978));
  NAND2_X1  g0778(.A1(new_n978), .A2(new_n718), .ZN(new_n979));
  INV_X1    g0779(.A(new_n707), .ZN(new_n980));
  OAI221_X1 g0780(.A(new_n719), .B1(new_n204), .B2(new_n310), .C1(new_n237), .C2(new_n980), .ZN(new_n981));
  NAND4_X1  g0781(.A1(new_n958), .A2(new_n979), .A3(new_n705), .A4(new_n981), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n957), .A2(new_n982), .ZN(G387));
  OAI221_X1 g0783(.A(new_n959), .B1(new_n208), .B2(new_n739), .C1(new_n249), .C2(new_n738), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n732), .A2(new_n309), .ZN(new_n985));
  OAI21_X1  g0785(.A(new_n985), .B1(new_n214), .B2(new_n727), .ZN(new_n986));
  NOR2_X1   g0786(.A1(new_n722), .A2(new_n216), .ZN(new_n987));
  OAI21_X1  g0787(.A(new_n270), .B1(new_n741), .B2(new_n333), .ZN(new_n988));
  OR3_X1    g0788(.A1(new_n986), .A2(new_n987), .A3(new_n988), .ZN(new_n989));
  AOI211_X1 g0789(.A(new_n984), .B(new_n989), .C1(G150), .C2(new_n751), .ZN(new_n990));
  XNOR2_X1  g0790(.A(new_n990), .B(KEYINPUT112), .ZN(new_n991));
  AOI22_X1  g0791(.A1(G322), .A2(new_n742), .B1(new_n745), .B2(G311), .ZN(new_n992));
  OAI221_X1 g0792(.A(new_n992), .B1(new_n434), .B2(new_n739), .C1(new_n746), .C2(new_n727), .ZN(new_n993));
  XNOR2_X1  g0793(.A(new_n993), .B(KEYINPUT48), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n784), .A2(G294), .ZN(new_n995));
  OAI211_X1 g0795(.A(new_n994), .B(new_n995), .C1(new_n795), .C2(new_n731), .ZN(new_n996));
  XOR2_X1   g0796(.A(new_n996), .B(KEYINPUT49), .Z(new_n997));
  AOI21_X1  g0797(.A(new_n270), .B1(new_n751), .B2(G326), .ZN(new_n998));
  OAI21_X1  g0798(.A(new_n998), .B1(new_n416), .B2(new_n724), .ZN(new_n999));
  OAI21_X1  g0799(.A(new_n991), .B1(new_n997), .B2(new_n999), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n1000), .A2(new_n718), .ZN(new_n1001));
  OAI21_X1  g0801(.A(new_n1001), .B1(new_n651), .B2(new_n716), .ZN(new_n1002));
  NAND3_X1  g0802(.A1(new_n659), .A2(new_n204), .A3(new_n270), .ZN(new_n1003));
  OAI21_X1  g0803(.A(new_n1003), .B1(G107), .B2(new_n204), .ZN(new_n1004));
  XNOR2_X1  g0804(.A(new_n1004), .B(KEYINPUT111), .ZN(new_n1005));
  OAI21_X1  g0805(.A(new_n707), .B1(new_n234), .B2(new_n437), .ZN(new_n1006));
  NAND2_X1  g0806(.A1(new_n306), .A2(new_n214), .ZN(new_n1007));
  OAI21_X1  g0807(.A(new_n660), .B1(KEYINPUT50), .B2(new_n1007), .ZN(new_n1008));
  NOR2_X1   g0808(.A1(new_n208), .A2(new_n216), .ZN(new_n1009));
  AND2_X1   g0809(.A1(new_n1007), .A2(KEYINPUT50), .ZN(new_n1010));
  NOR4_X1   g0810(.A1(new_n1008), .A2(G45), .A3(new_n1009), .A4(new_n1010), .ZN(new_n1011));
  OAI21_X1  g0811(.A(new_n1005), .B1(new_n1006), .B2(new_n1011), .ZN(new_n1012));
  AOI21_X1  g0812(.A(new_n1002), .B1(new_n719), .B2(new_n1012), .ZN(new_n1013));
  AOI22_X1  g0813(.A1(new_n936), .A2(new_n956), .B1(new_n1013), .B2(new_n705), .ZN(new_n1014));
  INV_X1    g0814(.A(new_n661), .ZN(new_n1015));
  OAI21_X1  g0815(.A(new_n1015), .B1(new_n701), .B2(new_n936), .ZN(new_n1016));
  OAI21_X1  g0816(.A(new_n1014), .B1(new_n1016), .B2(new_n952), .ZN(G393));
  NAND2_X1  g0817(.A1(new_n951), .A2(new_n956), .ZN(new_n1018));
  NAND3_X1  g0818(.A1(new_n927), .A2(new_n717), .A3(new_n928), .ZN(new_n1019));
  OAI221_X1 g0819(.A(new_n719), .B1(new_n409), .B2(new_n204), .C1(new_n980), .C2(new_n245), .ZN(new_n1020));
  OAI22_X1  g0820(.A1(new_n741), .A2(new_n255), .B1(new_n727), .B2(new_n333), .ZN(new_n1021));
  XNOR2_X1  g0821(.A(new_n1021), .B(KEYINPUT51), .ZN(new_n1022));
  AOI22_X1  g0822(.A1(G87), .A2(new_n753), .B1(new_n732), .B2(G77), .ZN(new_n1023));
  NAND2_X1  g0823(.A1(new_n751), .A2(G143), .ZN(new_n1024));
  NAND3_X1  g0824(.A1(new_n1022), .A2(new_n1023), .A3(new_n1024), .ZN(new_n1025));
  OAI22_X1  g0825(.A1(new_n738), .A2(new_n214), .B1(new_n739), .B2(new_n249), .ZN(new_n1026));
  XNOR2_X1  g0826(.A(new_n1026), .B(KEYINPUT113), .ZN(new_n1027));
  OAI21_X1  g0827(.A(new_n270), .B1(new_n722), .B2(new_n208), .ZN(new_n1028));
  NOR3_X1   g0828(.A1(new_n1025), .A2(new_n1027), .A3(new_n1028), .ZN(new_n1029));
  XNOR2_X1  g0829(.A(new_n1029), .B(KEYINPUT114), .ZN(new_n1030));
  AOI22_X1  g0830(.A1(G107), .A2(new_n753), .B1(new_n779), .B2(G294), .ZN(new_n1031));
  NAND2_X1  g0831(.A1(new_n751), .A2(G322), .ZN(new_n1032));
  OAI211_X1 g0832(.A(new_n1031), .B(new_n1032), .C1(new_n434), .C2(new_n738), .ZN(new_n1033));
  AOI211_X1 g0833(.A(new_n270), .B(new_n1033), .C1(G283), .C2(new_n784), .ZN(new_n1034));
  OAI21_X1  g0834(.A(new_n1034), .B1(new_n416), .B2(new_n731), .ZN(new_n1035));
  OAI22_X1  g0835(.A1(new_n741), .A2(new_n746), .B1(new_n727), .B2(new_n759), .ZN(new_n1036));
  XOR2_X1   g0836(.A(new_n1036), .B(KEYINPUT52), .Z(new_n1037));
  NOR2_X1   g0837(.A1(new_n1035), .A2(new_n1037), .ZN(new_n1038));
  OAI21_X1  g0838(.A(new_n718), .B1(new_n1030), .B2(new_n1038), .ZN(new_n1039));
  NAND4_X1  g0839(.A1(new_n1019), .A2(new_n705), .A3(new_n1020), .A4(new_n1039), .ZN(new_n1040));
  NAND2_X1  g0840(.A1(new_n1018), .A2(new_n1040), .ZN(new_n1041));
  NAND3_X1  g0841(.A1(new_n937), .A2(new_n947), .A3(new_n950), .ZN(new_n1042));
  AND2_X1   g0842(.A1(new_n954), .A2(new_n1042), .ZN(new_n1043));
  AOI21_X1  g0843(.A(new_n1041), .B1(new_n1043), .B2(new_n1015), .ZN(new_n1044));
  INV_X1    g0844(.A(new_n1044), .ZN(G390));
  INV_X1    g0845(.A(new_n858), .ZN(new_n1046));
  AOI21_X1  g0846(.A(new_n769), .B1(new_n674), .B2(new_n768), .ZN(new_n1047));
  OAI211_X1 g0847(.A(new_n868), .B(new_n1046), .C1(new_n1047), .C2(new_n863), .ZN(new_n1048));
  NAND2_X1  g0848(.A1(new_n774), .A2(new_n770), .ZN(new_n1049));
  AOI21_X1  g0849(.A(new_n858), .B1(new_n1049), .B2(new_n870), .ZN(new_n1050));
  OAI21_X1  g0850(.A(new_n1048), .B1(new_n857), .B2(new_n1050), .ZN(new_n1051));
  INV_X1    g0851(.A(KEYINPUT116), .ZN(new_n1052));
  NOR3_X1   g0852(.A1(new_n699), .A2(new_n863), .A3(new_n771), .ZN(new_n1053));
  NOR3_X1   g0853(.A1(new_n1051), .A2(new_n1052), .A3(new_n1053), .ZN(new_n1054));
  NAND3_X1  g0854(.A1(new_n892), .A2(G330), .A3(new_n872), .ZN(new_n1055));
  NAND2_X1  g0855(.A1(new_n1055), .A2(KEYINPUT115), .ZN(new_n1056));
  INV_X1    g0856(.A(KEYINPUT115), .ZN(new_n1057));
  NAND3_X1  g0857(.A1(new_n901), .A2(new_n1057), .A3(new_n872), .ZN(new_n1058));
  NAND2_X1  g0858(.A1(new_n1056), .A2(new_n1058), .ZN(new_n1059));
  NAND2_X1  g0859(.A1(new_n1051), .A2(new_n1059), .ZN(new_n1060));
  NAND2_X1  g0860(.A1(new_n1060), .A2(KEYINPUT116), .ZN(new_n1061));
  OR2_X1    g0861(.A1(new_n857), .A2(new_n1050), .ZN(new_n1062));
  INV_X1    g0862(.A(new_n1053), .ZN(new_n1063));
  NAND3_X1  g0863(.A1(new_n1062), .A2(new_n1048), .A3(new_n1063), .ZN(new_n1064));
  AOI21_X1  g0864(.A(new_n1054), .B1(new_n1061), .B2(new_n1064), .ZN(new_n1065));
  NAND2_X1  g0865(.A1(new_n1065), .A2(new_n956), .ZN(new_n1066));
  NAND3_X1  g0866(.A1(new_n853), .A2(new_n799), .A3(new_n856), .ZN(new_n1067));
  NAND2_X1  g0867(.A1(new_n800), .A2(new_n249), .ZN(new_n1068));
  XOR2_X1   g0868(.A(KEYINPUT54), .B(G143), .Z(new_n1069));
  XNOR2_X1  g0869(.A(new_n1069), .B(KEYINPUT118), .ZN(new_n1070));
  AOI22_X1  g0870(.A1(new_n1070), .A2(new_n779), .B1(G50), .B2(new_n753), .ZN(new_n1071));
  AOI22_X1  g0871(.A1(G132), .A2(new_n728), .B1(new_n745), .B2(G137), .ZN(new_n1072));
  INV_X1    g0872(.A(G125), .ZN(new_n1073));
  OAI211_X1 g0873(.A(new_n1071), .B(new_n1072), .C1(new_n1073), .C2(new_n734), .ZN(new_n1074));
  NOR3_X1   g0874(.A1(new_n722), .A2(KEYINPUT53), .A3(new_n255), .ZN(new_n1075));
  NOR2_X1   g0875(.A1(new_n731), .A2(new_n333), .ZN(new_n1076));
  OAI21_X1  g0876(.A(KEYINPUT53), .B1(new_n722), .B2(new_n255), .ZN(new_n1077));
  INV_X1    g0877(.A(G128), .ZN(new_n1078));
  OAI211_X1 g0878(.A(new_n1077), .B(new_n270), .C1(new_n1078), .C2(new_n741), .ZN(new_n1079));
  NOR4_X1   g0879(.A1(new_n1074), .A2(new_n1075), .A3(new_n1076), .A4(new_n1079), .ZN(new_n1080));
  NOR2_X1   g0880(.A1(new_n722), .A2(new_n790), .ZN(new_n1081));
  AOI22_X1  g0881(.A1(G283), .A2(new_n742), .B1(new_n753), .B2(G68), .ZN(new_n1082));
  AOI22_X1  g0882(.A1(G294), .A2(new_n751), .B1(new_n732), .B2(G77), .ZN(new_n1083));
  NAND2_X1  g0883(.A1(new_n779), .A2(G97), .ZN(new_n1084));
  AOI21_X1  g0884(.A(new_n270), .B1(new_n728), .B2(G116), .ZN(new_n1085));
  NAND4_X1  g0885(.A1(new_n1082), .A2(new_n1083), .A3(new_n1084), .A4(new_n1085), .ZN(new_n1086));
  AOI211_X1 g0886(.A(new_n1081), .B(new_n1086), .C1(G107), .C2(new_n745), .ZN(new_n1087));
  OAI21_X1  g0887(.A(new_n718), .B1(new_n1080), .B2(new_n1087), .ZN(new_n1088));
  NAND4_X1  g0888(.A1(new_n1067), .A2(new_n705), .A3(new_n1068), .A4(new_n1088), .ZN(new_n1089));
  NAND2_X1  g0889(.A1(new_n1066), .A2(new_n1089), .ZN(new_n1090));
  OAI211_X1 g0890(.A(new_n902), .B(new_n633), .C1(new_n678), .C2(new_n406), .ZN(new_n1091));
  AOI21_X1  g0891(.A(new_n870), .B1(new_n901), .B2(new_n773), .ZN(new_n1092));
  NAND2_X1  g0892(.A1(new_n671), .A2(new_n673), .ZN(new_n1093));
  NAND3_X1  g0893(.A1(new_n1093), .A2(new_n653), .A3(new_n768), .ZN(new_n1094));
  NAND2_X1  g0894(.A1(new_n1094), .A2(new_n770), .ZN(new_n1095));
  NOR4_X1   g0895(.A1(new_n1092), .A2(KEYINPUT117), .A3(new_n1053), .A4(new_n1095), .ZN(new_n1096));
  INV_X1    g0896(.A(KEYINPUT117), .ZN(new_n1097));
  OAI211_X1 g0897(.A(G330), .B(new_n773), .C1(new_n877), .C2(new_n881), .ZN(new_n1098));
  AOI21_X1  g0898(.A(new_n1095), .B1(new_n1098), .B2(new_n863), .ZN(new_n1099));
  AOI21_X1  g0899(.A(new_n1097), .B1(new_n1099), .B2(new_n1063), .ZN(new_n1100));
  NOR2_X1   g0900(.A1(new_n1096), .A2(new_n1100), .ZN(new_n1101));
  OAI21_X1  g0901(.A(new_n863), .B1(new_n699), .B2(new_n771), .ZN(new_n1102));
  NAND3_X1  g0902(.A1(new_n1056), .A2(new_n1058), .A3(new_n1102), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n1103), .A2(new_n1049), .ZN(new_n1104));
  AOI21_X1  g0904(.A(new_n1091), .B1(new_n1101), .B2(new_n1104), .ZN(new_n1105));
  AOI21_X1  g0905(.A(new_n661), .B1(new_n1065), .B2(new_n1105), .ZN(new_n1106));
  INV_X1    g0906(.A(new_n1105), .ZN(new_n1107));
  NAND4_X1  g0907(.A1(new_n1062), .A2(KEYINPUT116), .A3(new_n1048), .A4(new_n1063), .ZN(new_n1108));
  AOI21_X1  g0908(.A(new_n1052), .B1(new_n1051), .B2(new_n1059), .ZN(new_n1109));
  NOR2_X1   g0909(.A1(new_n1051), .A2(new_n1053), .ZN(new_n1110));
  OAI21_X1  g0910(.A(new_n1108), .B1(new_n1109), .B2(new_n1110), .ZN(new_n1111));
  NAND2_X1  g0911(.A1(new_n1107), .A2(new_n1111), .ZN(new_n1112));
  AOI21_X1  g0912(.A(new_n1090), .B1(new_n1106), .B2(new_n1112), .ZN(new_n1113));
  INV_X1    g0913(.A(new_n1113), .ZN(G378));
  AOI21_X1  g0914(.A(new_n1091), .B1(new_n1065), .B2(new_n1105), .ZN(new_n1115));
  AOI21_X1  g0915(.A(KEYINPUT124), .B1(new_n859), .B2(new_n865), .ZN(new_n1116));
  XOR2_X1   g0916(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1117));
  XNOR2_X1  g0917(.A(new_n297), .B(new_n1117), .ZN(new_n1118));
  NAND2_X1  g0918(.A1(new_n265), .A2(new_n640), .ZN(new_n1119));
  XNOR2_X1  g0919(.A(new_n1118), .B(new_n1119), .ZN(new_n1120));
  INV_X1    g0920(.A(new_n1120), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n898), .A2(new_n1121), .ZN(new_n1122));
  NAND4_X1  g0922(.A1(new_n891), .A2(G330), .A3(new_n894), .A4(new_n1120), .ZN(new_n1123));
  AOI21_X1  g0923(.A(new_n1116), .B1(new_n1122), .B2(new_n1123), .ZN(new_n1124));
  NAND2_X1  g0924(.A1(new_n1122), .A2(new_n1123), .ZN(new_n1125));
  INV_X1    g0925(.A(new_n1125), .ZN(new_n1126));
  INV_X1    g0926(.A(new_n1116), .ZN(new_n1127));
  NAND3_X1  g0927(.A1(new_n859), .A2(KEYINPUT124), .A3(new_n865), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n1127), .A2(new_n1128), .ZN(new_n1129));
  AOI21_X1  g0929(.A(new_n1124), .B1(new_n1126), .B2(new_n1129), .ZN(new_n1130));
  OAI21_X1  g0930(.A(KEYINPUT57), .B1(new_n1115), .B2(new_n1130), .ZN(new_n1131));
  INV_X1    g0931(.A(new_n1091), .ZN(new_n1132));
  NAND2_X1  g0932(.A1(new_n1099), .A2(new_n1063), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n1133), .A2(KEYINPUT117), .ZN(new_n1134));
  NAND3_X1  g0934(.A1(new_n1099), .A2(new_n1097), .A3(new_n1063), .ZN(new_n1135));
  NAND3_X1  g0935(.A1(new_n1134), .A2(new_n1104), .A3(new_n1135), .ZN(new_n1136));
  INV_X1    g0936(.A(new_n1136), .ZN(new_n1137));
  OAI21_X1  g0937(.A(new_n1132), .B1(new_n1111), .B2(new_n1137), .ZN(new_n1138));
  AOI21_X1  g0938(.A(KEYINPUT122), .B1(new_n1122), .B2(new_n1123), .ZN(new_n1139));
  INV_X1    g0939(.A(KEYINPUT123), .ZN(new_n1140));
  OAI21_X1  g0940(.A(new_n866), .B1(new_n1139), .B2(new_n1140), .ZN(new_n1141));
  INV_X1    g0941(.A(KEYINPUT57), .ZN(new_n1142));
  NOR2_X1   g0942(.A1(new_n866), .A2(new_n1140), .ZN(new_n1143));
  OAI211_X1 g0943(.A(new_n1123), .B(new_n1122), .C1(new_n1143), .C2(KEYINPUT122), .ZN(new_n1144));
  NAND4_X1  g0944(.A1(new_n1138), .A2(new_n1141), .A3(new_n1142), .A4(new_n1144), .ZN(new_n1145));
  AOI21_X1  g0945(.A(new_n661), .B1(new_n1131), .B2(new_n1145), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n1141), .A2(new_n1144), .ZN(new_n1147));
  INV_X1    g0947(.A(new_n956), .ZN(new_n1148));
  NOR2_X1   g0948(.A1(new_n1147), .A2(new_n1148), .ZN(new_n1149));
  NOR2_X1   g0949(.A1(new_n1146), .A2(new_n1149), .ZN(new_n1150));
  AOI22_X1  g0950(.A1(new_n1120), .A2(new_n799), .B1(new_n214), .B2(new_n800), .ZN(new_n1151));
  OAI22_X1  g0951(.A1(new_n741), .A2(new_n416), .B1(new_n734), .B2(new_n795), .ZN(new_n1152));
  AOI22_X1  g0952(.A1(new_n745), .A2(G97), .B1(new_n779), .B2(new_n309), .ZN(new_n1153));
  OR2_X1    g0953(.A1(new_n1153), .A2(KEYINPUT120), .ZN(new_n1154));
  NAND2_X1  g0954(.A1(new_n1153), .A2(KEYINPUT120), .ZN(new_n1155));
  AOI211_X1 g0955(.A(G41), .B(new_n1152), .C1(new_n1154), .C2(new_n1155), .ZN(new_n1156));
  NOR2_X1   g0956(.A1(new_n724), .A2(new_n219), .ZN(new_n1157));
  XNOR2_X1  g0957(.A(new_n1157), .B(KEYINPUT119), .ZN(new_n1158));
  NAND2_X1  g0958(.A1(new_n1158), .A2(new_n972), .ZN(new_n1159));
  NOR3_X1   g0959(.A1(new_n1159), .A2(new_n270), .A3(new_n987), .ZN(new_n1160));
  OAI211_X1 g0960(.A(new_n1156), .B(new_n1160), .C1(new_n210), .C2(new_n727), .ZN(new_n1161));
  XOR2_X1   g0961(.A(new_n1161), .B(KEYINPUT58), .Z(new_n1162));
  OAI21_X1  g0962(.A(new_n214), .B1(new_n323), .B2(G41), .ZN(new_n1163));
  NOR2_X1   g0963(.A1(new_n727), .A2(new_n1078), .ZN(new_n1164));
  OAI22_X1  g0964(.A1(new_n741), .A2(new_n1073), .B1(new_n731), .B2(new_n255), .ZN(new_n1165));
  AOI211_X1 g0965(.A(new_n1164), .B(new_n1165), .C1(new_n1070), .C2(new_n784), .ZN(new_n1166));
  NAND2_X1  g0966(.A1(new_n745), .A2(G132), .ZN(new_n1167));
  OAI211_X1 g0967(.A(new_n1166), .B(new_n1167), .C1(new_n781), .C2(new_n739), .ZN(new_n1168));
  OR2_X1    g0968(.A1(new_n1168), .A2(KEYINPUT59), .ZN(new_n1169));
  NAND2_X1  g0969(.A1(new_n753), .A2(G159), .ZN(new_n1170));
  AOI21_X1  g0970(.A(G41), .B1(new_n751), .B2(G124), .ZN(new_n1171));
  NAND4_X1  g0971(.A1(new_n1169), .A2(new_n253), .A3(new_n1170), .A4(new_n1171), .ZN(new_n1172));
  AND2_X1   g0972(.A1(new_n1168), .A2(KEYINPUT59), .ZN(new_n1173));
  OAI21_X1  g0973(.A(new_n1163), .B1(new_n1172), .B2(new_n1173), .ZN(new_n1174));
  OAI21_X1  g0974(.A(new_n718), .B1(new_n1162), .B2(new_n1174), .ZN(new_n1175));
  NAND3_X1  g0975(.A1(new_n1151), .A2(new_n705), .A3(new_n1175), .ZN(new_n1176));
  XNOR2_X1  g0976(.A(new_n1176), .B(KEYINPUT121), .ZN(new_n1177));
  NAND2_X1  g0977(.A1(new_n1150), .A2(new_n1177), .ZN(G375));
  OAI21_X1  g0978(.A(new_n1158), .B1(new_n1078), .B2(new_n734), .ZN(new_n1179));
  AOI22_X1  g0979(.A1(G137), .A2(new_n728), .B1(new_n779), .B2(G150), .ZN(new_n1180));
  AOI21_X1  g0980(.A(new_n350), .B1(new_n742), .B2(G132), .ZN(new_n1181));
  OAI211_X1 g0981(.A(new_n1180), .B(new_n1181), .C1(new_n214), .C2(new_n731), .ZN(new_n1182));
  AND2_X1   g0982(.A1(new_n1070), .A2(new_n745), .ZN(new_n1183));
  NOR2_X1   g0983(.A1(new_n722), .A2(new_n333), .ZN(new_n1184));
  NOR4_X1   g0984(.A1(new_n1179), .A2(new_n1182), .A3(new_n1183), .A4(new_n1184), .ZN(new_n1185));
  AOI22_X1  g0985(.A1(G294), .A2(new_n742), .B1(new_n753), .B2(G77), .ZN(new_n1186));
  OAI211_X1 g0986(.A(new_n1186), .B(new_n985), .C1(new_n434), .C2(new_n734), .ZN(new_n1187));
  OAI221_X1 g0987(.A(new_n350), .B1(new_n739), .B2(new_n210), .C1(new_n409), .C2(new_n722), .ZN(new_n1188));
  NOR2_X1   g0988(.A1(new_n727), .A2(new_n795), .ZN(new_n1189));
  NOR2_X1   g0989(.A1(new_n738), .A2(new_n416), .ZN(new_n1190));
  NOR4_X1   g0990(.A1(new_n1187), .A2(new_n1188), .A3(new_n1189), .A4(new_n1190), .ZN(new_n1191));
  OAI21_X1  g0991(.A(new_n718), .B1(new_n1185), .B2(new_n1191), .ZN(new_n1192));
  INV_X1    g0992(.A(new_n799), .ZN(new_n1193));
  OAI211_X1 g0993(.A(new_n705), .B(new_n1192), .C1(new_n870), .C2(new_n1193), .ZN(new_n1194));
  AOI21_X1  g0994(.A(new_n1194), .B1(new_n208), .B2(new_n800), .ZN(new_n1195));
  AOI21_X1  g0995(.A(new_n1195), .B1(new_n1136), .B2(new_n956), .ZN(new_n1196));
  OAI21_X1  g0996(.A(new_n932), .B1(new_n1136), .B2(new_n1132), .ZN(new_n1197));
  OAI21_X1  g0997(.A(new_n1196), .B1(new_n1197), .B2(new_n1105), .ZN(G381));
  NOR2_X1   g0998(.A1(G375), .A2(G378), .ZN(new_n1199));
  INV_X1    g0999(.A(G384), .ZN(new_n1200));
  INV_X1    g1000(.A(G381), .ZN(new_n1201));
  NAND3_X1  g1001(.A1(new_n1044), .A2(new_n957), .A3(new_n982), .ZN(new_n1202));
  NOR3_X1   g1002(.A1(new_n1202), .A2(G396), .A3(G393), .ZN(new_n1203));
  NAND4_X1  g1003(.A1(new_n1199), .A2(new_n1200), .A3(new_n1201), .A4(new_n1203), .ZN(G407));
  NAND2_X1  g1004(.A1(new_n642), .A2(G213), .ZN(new_n1205));
  XOR2_X1   g1005(.A(new_n1205), .B(KEYINPUT125), .Z(new_n1206));
  INV_X1    g1006(.A(new_n1206), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n1199), .A2(new_n1207), .ZN(new_n1208));
  NAND3_X1  g1008(.A1(G407), .A2(G213), .A3(new_n1208), .ZN(G409));
  XNOR2_X1  g1009(.A(G393), .B(G396), .ZN(new_n1210));
  XNOR2_X1  g1010(.A(new_n1210), .B(KEYINPUT126), .ZN(new_n1211));
  INV_X1    g1011(.A(new_n1202), .ZN(new_n1212));
  AOI21_X1  g1012(.A(new_n1044), .B1(new_n957), .B2(new_n982), .ZN(new_n1213));
  OAI21_X1  g1013(.A(new_n1211), .B1(new_n1212), .B2(new_n1213), .ZN(new_n1214));
  NAND2_X1  g1014(.A1(G387), .A2(G390), .ZN(new_n1215));
  INV_X1    g1015(.A(KEYINPUT126), .ZN(new_n1216));
  XNOR2_X1  g1016(.A(new_n1210), .B(new_n1216), .ZN(new_n1217));
  NAND3_X1  g1017(.A1(new_n1215), .A2(new_n1217), .A3(new_n1202), .ZN(new_n1218));
  AND2_X1   g1018(.A1(new_n1214), .A2(new_n1218), .ZN(new_n1219));
  NAND3_X1  g1019(.A1(new_n1137), .A2(KEYINPUT60), .A3(new_n1091), .ZN(new_n1220));
  INV_X1    g1020(.A(KEYINPUT60), .ZN(new_n1221));
  OAI21_X1  g1021(.A(new_n1221), .B1(new_n1136), .B2(new_n1132), .ZN(new_n1222));
  NAND4_X1  g1022(.A1(new_n1220), .A2(new_n1107), .A3(new_n1015), .A4(new_n1222), .ZN(new_n1223));
  NAND3_X1  g1023(.A1(new_n1223), .A2(G384), .A3(new_n1196), .ZN(new_n1224));
  INV_X1    g1024(.A(new_n1224), .ZN(new_n1225));
  AOI21_X1  g1025(.A(G384), .B1(new_n1223), .B2(new_n1196), .ZN(new_n1226));
  NOR2_X1   g1026(.A1(new_n1225), .A2(new_n1226), .ZN(new_n1227));
  INV_X1    g1027(.A(new_n1177), .ZN(new_n1228));
  NOR4_X1   g1028(.A1(new_n1146), .A2(new_n1113), .A3(new_n1149), .A4(new_n1228), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n1138), .A2(new_n932), .ZN(new_n1230));
  OAI221_X1 g1030(.A(new_n1176), .B1(new_n1148), .B2(new_n1130), .C1(new_n1230), .C2(new_n1147), .ZN(new_n1231));
  NAND2_X1  g1031(.A1(new_n1231), .A2(new_n1113), .ZN(new_n1232));
  INV_X1    g1032(.A(new_n1232), .ZN(new_n1233));
  OAI211_X1 g1033(.A(new_n1205), .B(new_n1227), .C1(new_n1229), .C2(new_n1233), .ZN(new_n1234));
  INV_X1    g1034(.A(KEYINPUT62), .ZN(new_n1235));
  INV_X1    g1035(.A(new_n1145), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n1126), .A2(new_n1129), .ZN(new_n1237));
  INV_X1    g1037(.A(new_n1124), .ZN(new_n1238));
  NAND2_X1  g1038(.A1(new_n1237), .A2(new_n1238), .ZN(new_n1239));
  AOI21_X1  g1039(.A(new_n1142), .B1(new_n1239), .B2(new_n1138), .ZN(new_n1240));
  OAI21_X1  g1040(.A(new_n1015), .B1(new_n1236), .B2(new_n1240), .ZN(new_n1241));
  INV_X1    g1041(.A(new_n1149), .ZN(new_n1242));
  NAND4_X1  g1042(.A1(new_n1241), .A2(G378), .A3(new_n1242), .A4(new_n1177), .ZN(new_n1243));
  AOI21_X1  g1043(.A(new_n1207), .B1(new_n1243), .B2(new_n1232), .ZN(new_n1244));
  INV_X1    g1044(.A(new_n1227), .ZN(new_n1245));
  NOR2_X1   g1045(.A1(new_n1245), .A2(new_n1235), .ZN(new_n1246));
  AOI22_X1  g1046(.A1(new_n1234), .A2(new_n1235), .B1(new_n1244), .B2(new_n1246), .ZN(new_n1247));
  INV_X1    g1047(.A(KEYINPUT61), .ZN(new_n1248));
  INV_X1    g1048(.A(new_n1226), .ZN(new_n1249));
  AOI21_X1  g1049(.A(new_n1206), .B1(new_n1249), .B2(new_n1224), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(new_n1250), .A2(G2897), .ZN(new_n1251));
  NAND3_X1  g1051(.A1(new_n642), .A2(G213), .A3(G2897), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(new_n1227), .A2(new_n1252), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(new_n1251), .A2(new_n1253), .ZN(new_n1254));
  OAI21_X1  g1054(.A(new_n1248), .B1(new_n1254), .B2(new_n1244), .ZN(new_n1255));
  OAI21_X1  g1055(.A(new_n1219), .B1(new_n1247), .B2(new_n1255), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(new_n1214), .A2(new_n1218), .ZN(new_n1257));
  INV_X1    g1057(.A(KEYINPUT63), .ZN(new_n1258));
  NOR2_X1   g1058(.A1(new_n1245), .A2(new_n1258), .ZN(new_n1259));
  AOI21_X1  g1059(.A(KEYINPUT61), .B1(new_n1244), .B2(new_n1259), .ZN(new_n1260));
  OAI21_X1  g1060(.A(new_n1205), .B1(new_n1229), .B2(new_n1233), .ZN(new_n1261));
  AOI22_X1  g1061(.A1(new_n1250), .A2(G2897), .B1(new_n1227), .B2(new_n1252), .ZN(new_n1262));
  AOI21_X1  g1062(.A(new_n1258), .B1(new_n1261), .B2(new_n1262), .ZN(new_n1263));
  INV_X1    g1063(.A(new_n1234), .ZN(new_n1264));
  OAI211_X1 g1064(.A(new_n1257), .B(new_n1260), .C1(new_n1263), .C2(new_n1264), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(new_n1256), .A2(new_n1265), .ZN(G405));
  AOI21_X1  g1066(.A(G378), .B1(new_n1150), .B2(new_n1177), .ZN(new_n1267));
  INV_X1    g1067(.A(new_n1267), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1227), .A2(KEYINPUT127), .ZN(new_n1269));
  NAND3_X1  g1069(.A1(new_n1268), .A2(new_n1243), .A3(new_n1269), .ZN(new_n1270));
  OAI211_X1 g1070(.A(KEYINPUT127), .B(new_n1227), .C1(new_n1267), .C2(new_n1229), .ZN(new_n1271));
  AND3_X1   g1071(.A1(new_n1270), .A2(new_n1219), .A3(new_n1271), .ZN(new_n1272));
  AOI21_X1  g1072(.A(new_n1219), .B1(new_n1271), .B2(new_n1270), .ZN(new_n1273));
  NOR2_X1   g1073(.A1(new_n1272), .A2(new_n1273), .ZN(G402));
endmodule


