

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
         n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706,
         n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717,
         n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
         n729, n730, n731, n732, n733, n734;

  XNOR2_X2 U377 ( .A(n372), .B(n357), .ZN(n567) );
  NOR2_X2 U378 ( .A1(n543), .A2(n374), .ZN(n373) );
  XNOR2_X2 U379 ( .A(n427), .B(n426), .ZN(n543) );
  NOR2_X1 U380 ( .A1(n648), .A2(n647), .ZN(n580) );
  XNOR2_X2 U381 ( .A(n510), .B(n509), .ZN(n560) );
  XNOR2_X1 U382 ( .A(n537), .B(n536), .ZN(n596) );
  AND2_X1 U383 ( .A1(n583), .A2(n409), .ZN(n557) );
  NAND2_X1 U384 ( .A1(n394), .A2(n393), .ZN(n583) );
  XNOR2_X1 U385 ( .A(n466), .B(n407), .ZN(n651) );
  XNOR2_X1 U386 ( .A(n384), .B(G131), .ZN(n485) );
  XNOR2_X1 U387 ( .A(n382), .B(G107), .ZN(n432) );
  INV_X2 U388 ( .A(G953), .ZN(n721) );
  XNOR2_X1 U389 ( .A(KEYINPUT4), .B(G146), .ZN(n487) );
  XNOR2_X1 U390 ( .A(n401), .B(n413), .ZN(n437) );
  INV_X1 U391 ( .A(G143), .ZN(n413) );
  XNOR2_X1 U392 ( .A(G128), .B(KEYINPUT65), .ZN(n401) );
  XNOR2_X1 U393 ( .A(n452), .B(n451), .ZN(n525) );
  OR2_X1 U394 ( .A1(n687), .A2(G902), .ZN(n391) );
  XOR2_X1 U395 ( .A(G134), .B(n437), .Z(n488) );
  XNOR2_X1 U396 ( .A(G116), .B(G119), .ZN(n478) );
  XOR2_X1 U397 ( .A(KEYINPUT5), .B(KEYINPUT96), .Z(n479) );
  XNOR2_X1 U398 ( .A(n574), .B(n573), .ZN(n376) );
  NOR2_X1 U399 ( .A1(n592), .A2(n572), .ZN(n574) );
  XNOR2_X1 U400 ( .A(n400), .B(n399), .ZN(n398) );
  XNOR2_X1 U401 ( .A(n414), .B(KEYINPUT88), .ZN(n400) );
  NAND2_X1 U402 ( .A1(n721), .A2(G224), .ZN(n399) );
  XNOR2_X1 U403 ( .A(n487), .B(n364), .ZN(n418) );
  INV_X1 U404 ( .A(KEYINPUT17), .ZN(n364) );
  XNOR2_X1 U405 ( .A(KEYINPUT78), .B(KEYINPUT86), .ZN(n415) );
  XOR2_X1 U406 ( .A(G125), .B(KEYINPUT89), .Z(n416) );
  INV_X1 U407 ( .A(n560), .ZN(n576) );
  NAND2_X1 U408 ( .A1(n651), .A2(n477), .ZN(n511) );
  OR2_X1 U409 ( .A1(n602), .A2(G902), .ZN(n372) );
  XNOR2_X1 U410 ( .A(n424), .B(n423), .ZN(n481) );
  XOR2_X1 U411 ( .A(KEYINPUT73), .B(KEYINPUT3), .Z(n423) );
  INV_X1 U412 ( .A(KEYINPUT74), .ZN(n421) );
  INV_X1 U413 ( .A(G116), .ZN(n382) );
  INV_X1 U414 ( .A(KEYINPUT102), .ZN(n433) );
  XNOR2_X1 U415 ( .A(n449), .B(n448), .ZN(n691) );
  XNOR2_X1 U416 ( .A(n447), .B(n408), .ZN(n448) );
  XNOR2_X1 U417 ( .A(G113), .B(G143), .ZN(n408) );
  XNOR2_X1 U418 ( .A(n489), .B(n488), .ZN(n717) );
  XNOR2_X1 U419 ( .A(n355), .B(n487), .ZN(n489) );
  XOR2_X1 U420 ( .A(KEYINPUT71), .B(G137), .Z(n486) );
  XNOR2_X1 U421 ( .A(G101), .B(G104), .ZN(n492) );
  XOR2_X1 U422 ( .A(G110), .B(G107), .Z(n493) );
  AND2_X1 U423 ( .A1(n596), .A2(n367), .ZN(n599) );
  AND2_X1 U424 ( .A1(n598), .A2(n635), .ZN(n367) );
  NAND2_X1 U425 ( .A1(n390), .A2(n389), .ZN(n388) );
  INV_X1 U426 ( .A(KEYINPUT34), .ZN(n578) );
  NOR2_X1 U427 ( .A1(n648), .A2(n561), .ZN(n562) );
  XNOR2_X1 U428 ( .A(n373), .B(KEYINPUT19), .ZN(n552) );
  INV_X1 U429 ( .A(n638), .ZN(n374) );
  XNOR2_X1 U430 ( .A(n441), .B(n440), .ZN(n526) );
  XNOR2_X1 U431 ( .A(KEYINPUT85), .B(n571), .ZN(n592) );
  XNOR2_X1 U432 ( .A(G113), .B(G101), .ZN(n422) );
  XNOR2_X1 U433 ( .A(n406), .B(n405), .ZN(n719) );
  INV_X1 U434 ( .A(G125), .ZN(n405) );
  XNOR2_X1 U435 ( .A(KEYINPUT10), .B(G140), .ZN(n406) );
  INV_X1 U436 ( .A(KEYINPUT70), .ZN(n384) );
  XNOR2_X1 U437 ( .A(KEYINPUT48), .B(KEYINPUT83), .ZN(n536) );
  NOR2_X1 U438 ( .A1(n526), .A2(n525), .ZN(n554) );
  INV_X1 U439 ( .A(n501), .ZN(n369) );
  XNOR2_X1 U440 ( .A(n490), .B(n717), .ZN(n602) );
  XNOR2_X1 U441 ( .A(n380), .B(G122), .ZN(n442) );
  INV_X1 U442 ( .A(G104), .ZN(n380) );
  INV_X1 U443 ( .A(KEYINPUT16), .ZN(n379) );
  NAND2_X1 U444 ( .A1(n377), .A2(n376), .ZN(n375) );
  NOR2_X1 U445 ( .A1(n365), .A2(n356), .ZN(n377) );
  XNOR2_X1 U446 ( .A(n719), .B(G146), .ZN(n457) );
  XNOR2_X1 U447 ( .A(G128), .B(G137), .ZN(n454) );
  XNOR2_X1 U448 ( .A(n383), .B(G110), .ZN(n458) );
  INV_X1 U449 ( .A(G119), .ZN(n383) );
  NAND2_X1 U450 ( .A1(n359), .A2(n362), .ZN(n361) );
  INV_X1 U451 ( .A(n595), .ZN(n362) );
  XNOR2_X1 U452 ( .A(n437), .B(n398), .ZN(n420) );
  NOR2_X1 U453 ( .A1(n527), .A2(n503), .ZN(n505) );
  INV_X1 U454 ( .A(KEYINPUT1), .ZN(n366) );
  NAND2_X1 U455 ( .A1(n370), .A2(n368), .ZN(n527) );
  XNOR2_X1 U456 ( .A(n500), .B(n371), .ZN(n370) );
  AND2_X1 U457 ( .A1(n584), .A2(n369), .ZN(n368) );
  INV_X1 U458 ( .A(KEYINPUT30), .ZN(n371) );
  OR2_X1 U459 ( .A1(n552), .A2(n358), .ZN(n393) );
  AND2_X1 U460 ( .A1(n396), .A2(n395), .ZN(n394) );
  BUF_X1 U461 ( .A(n567), .Z(n657) );
  XNOR2_X1 U462 ( .A(n465), .B(n467), .ZN(n407) );
  NOR2_X1 U463 ( .A1(G902), .A2(n704), .ZN(n466) );
  INV_X1 U464 ( .A(KEYINPUT6), .ZN(n508) );
  XNOR2_X1 U465 ( .A(n481), .B(n425), .ZN(n712) );
  XNOR2_X1 U466 ( .A(n381), .B(n378), .ZN(n425) );
  XNOR2_X1 U467 ( .A(n442), .B(n379), .ZN(n378) );
  XNOR2_X1 U468 ( .A(n432), .B(n458), .ZN(n381) );
  XNOR2_X1 U469 ( .A(n436), .B(n435), .ZN(n439) );
  XNOR2_X1 U470 ( .A(n434), .B(n433), .ZN(n435) );
  XNOR2_X1 U471 ( .A(n692), .B(KEYINPUT122), .ZN(n693) );
  XNOR2_X1 U472 ( .A(n717), .B(n497), .ZN(n687) );
  XOR2_X1 U473 ( .A(KEYINPUT87), .B(n607), .Z(n706) );
  XNOR2_X1 U474 ( .A(n403), .B(n402), .ZN(n734) );
  XNOR2_X1 U475 ( .A(KEYINPUT42), .B(KEYINPUT107), .ZN(n402) );
  NOR2_X1 U476 ( .A1(n669), .A2(n518), .ZN(n403) );
  INV_X1 U477 ( .A(n579), .ZN(n386) );
  XOR2_X1 U478 ( .A(KEYINPUT31), .B(n582), .Z(n628) );
  NOR2_X1 U479 ( .A1(n581), .A2(n659), .ZN(n582) );
  AND2_X1 U480 ( .A1(n526), .A2(n519), .ZN(n627) );
  AND2_X1 U481 ( .A1(n677), .A2(n721), .ZN(n678) );
  NOR2_X1 U482 ( .A1(n675), .A2(n674), .ZN(n676) );
  XOR2_X1 U483 ( .A(n486), .B(n485), .Z(n355) );
  NAND2_X1 U484 ( .A1(n590), .A2(n575), .ZN(n356) );
  XOR2_X1 U485 ( .A(G472), .B(KEYINPUT97), .Z(n357) );
  OR2_X1 U486 ( .A1(n553), .A2(n397), .ZN(n358) );
  AND2_X1 U487 ( .A1(n392), .A2(n720), .ZN(n359) );
  XNOR2_X1 U488 ( .A(n404), .B(KEYINPUT40), .ZN(n732) );
  XNOR2_X1 U489 ( .A(KEYINPUT68), .B(n412), .ZN(n360) );
  NAND2_X1 U490 ( .A1(n589), .A2(n593), .ZN(n365) );
  NAND2_X1 U491 ( .A1(n361), .A2(n360), .ZN(n410) );
  XNOR2_X1 U492 ( .A(n712), .B(n363), .ZN(n680) );
  XNOR2_X1 U493 ( .A(n419), .B(n420), .ZN(n363) );
  XNOR2_X2 U494 ( .A(n507), .B(n366), .ZN(n648) );
  XNOR2_X2 U495 ( .A(n391), .B(n498), .ZN(n507) );
  INV_X1 U496 ( .A(n567), .ZN(n510) );
  XNOR2_X2 U497 ( .A(n375), .B(n594), .ZN(n392) );
  XNOR2_X2 U498 ( .A(n385), .B(KEYINPUT35), .ZN(n728) );
  NAND2_X1 U499 ( .A1(n387), .A2(n386), .ZN(n385) );
  XNOR2_X1 U500 ( .A(n388), .B(n578), .ZN(n387) );
  INV_X1 U501 ( .A(n581), .ZN(n389) );
  INV_X1 U502 ( .A(n668), .ZN(n390) );
  NAND2_X1 U503 ( .A1(n392), .A2(n599), .ZN(n600) );
  NAND2_X1 U504 ( .A1(n392), .A2(n721), .ZN(n710) );
  NAND2_X1 U505 ( .A1(n553), .A2(n397), .ZN(n395) );
  NAND2_X1 U506 ( .A1(n552), .A2(n397), .ZN(n396) );
  INV_X1 U507 ( .A(KEYINPUT0), .ZN(n397) );
  NAND2_X1 U508 ( .A1(n732), .A2(n734), .ZN(n506) );
  NAND2_X1 U509 ( .A1(n538), .A2(n623), .ZN(n404) );
  XNOR2_X1 U510 ( .A(n505), .B(n504), .ZN(n538) );
  NOR2_X1 U511 ( .A1(n510), .A2(n511), .ZN(n491) );
  XNOR2_X1 U512 ( .A(n457), .B(n443), .ZN(n444) );
  AND2_X1 U513 ( .A1(n555), .A2(n554), .ZN(n409) );
  XNOR2_X1 U514 ( .A(n442), .B(KEYINPUT99), .ZN(n443) );
  XNOR2_X1 U515 ( .A(n422), .B(n421), .ZN(n424) );
  XNOR2_X1 U516 ( .A(KEYINPUT75), .B(KEYINPUT39), .ZN(n504) );
  XNOR2_X1 U517 ( .A(n450), .B(G475), .ZN(n451) );
  XNOR2_X1 U518 ( .A(n508), .B(KEYINPUT104), .ZN(n509) );
  XNOR2_X1 U519 ( .A(n604), .B(n603), .ZN(n605) );
  XNOR2_X1 U520 ( .A(n687), .B(n686), .ZN(n688) );
  XNOR2_X1 U521 ( .A(n689), .B(n688), .ZN(n690) );
  XNOR2_X1 U522 ( .A(G902), .B(KEYINPUT15), .ZN(n595) );
  XOR2_X1 U523 ( .A(n595), .B(KEYINPUT82), .Z(n411) );
  NAND2_X1 U524 ( .A1(n411), .A2(KEYINPUT2), .ZN(n412) );
  INV_X1 U525 ( .A(KEYINPUT18), .ZN(n414) );
  XNOR2_X1 U526 ( .A(n416), .B(n415), .ZN(n417) );
  XNOR2_X1 U527 ( .A(n418), .B(n417), .ZN(n419) );
  NAND2_X1 U528 ( .A1(n680), .A2(n595), .ZN(n427) );
  OR2_X1 U529 ( .A1(G237), .A2(G902), .ZN(n428) );
  NAND2_X1 U530 ( .A1(G210), .A2(n428), .ZN(n426) );
  INV_X1 U531 ( .A(n543), .ZN(n528) );
  XOR2_X1 U532 ( .A(KEYINPUT38), .B(n528), .Z(n639) );
  NAND2_X1 U533 ( .A1(G214), .A2(n428), .ZN(n638) );
  NAND2_X1 U534 ( .A1(n639), .A2(n638), .ZN(n642) );
  XOR2_X1 U535 ( .A(KEYINPUT7), .B(KEYINPUT9), .Z(n431) );
  NAND2_X1 U536 ( .A1(G234), .A2(n721), .ZN(n429) );
  XOR2_X1 U537 ( .A(KEYINPUT8), .B(n429), .Z(n459) );
  NAND2_X1 U538 ( .A1(G217), .A2(n459), .ZN(n430) );
  XNOR2_X1 U539 ( .A(n431), .B(n430), .ZN(n436) );
  XNOR2_X1 U540 ( .A(n432), .B(G122), .ZN(n434) );
  INV_X1 U541 ( .A(n488), .ZN(n438) );
  XOR2_X1 U542 ( .A(n439), .B(n438), .Z(n700) );
  NOR2_X1 U543 ( .A1(G902), .A2(n700), .ZN(n441) );
  XNOR2_X1 U544 ( .A(KEYINPUT103), .B(G478), .ZN(n440) );
  XNOR2_X1 U545 ( .A(n444), .B(n485), .ZN(n449) );
  XOR2_X1 U546 ( .A(KEYINPUT12), .B(KEYINPUT11), .Z(n446) );
  NOR2_X1 U547 ( .A1(G953), .A2(G237), .ZN(n482) );
  NAND2_X1 U548 ( .A1(G214), .A2(n482), .ZN(n445) );
  XNOR2_X1 U549 ( .A(n446), .B(n445), .ZN(n447) );
  NOR2_X1 U550 ( .A1(G902), .A2(n691), .ZN(n452) );
  XNOR2_X1 U551 ( .A(KEYINPUT100), .B(KEYINPUT13), .ZN(n450) );
  INV_X1 U552 ( .A(n554), .ZN(n641) );
  NOR2_X1 U553 ( .A1(n642), .A2(n641), .ZN(n453) );
  XNOR2_X1 U554 ( .A(KEYINPUT41), .B(n453), .ZN(n669) );
  XNOR2_X1 U555 ( .A(KEYINPUT93), .B(KEYINPUT25), .ZN(n467) );
  XOR2_X1 U556 ( .A(KEYINPUT24), .B(KEYINPUT92), .Z(n455) );
  XNOR2_X1 U557 ( .A(n455), .B(n454), .ZN(n456) );
  XNOR2_X1 U558 ( .A(n457), .B(n456), .ZN(n463) );
  XOR2_X1 U559 ( .A(n458), .B(KEYINPUT23), .Z(n461) );
  NAND2_X1 U560 ( .A1(G221), .A2(n459), .ZN(n460) );
  XNOR2_X1 U561 ( .A(n461), .B(n460), .ZN(n462) );
  XNOR2_X1 U562 ( .A(n463), .B(n462), .ZN(n704) );
  NAND2_X1 U563 ( .A1(G234), .A2(n595), .ZN(n464) );
  XNOR2_X1 U564 ( .A(KEYINPUT20), .B(n464), .ZN(n473) );
  NAND2_X1 U565 ( .A1(G217), .A2(n473), .ZN(n465) );
  NAND2_X1 U566 ( .A1(G234), .A2(G237), .ZN(n468) );
  XNOR2_X1 U567 ( .A(n468), .B(KEYINPUT90), .ZN(n469) );
  XNOR2_X1 U568 ( .A(KEYINPUT14), .B(n469), .ZN(n470) );
  NAND2_X1 U569 ( .A1(G952), .A2(n470), .ZN(n667) );
  NOR2_X1 U570 ( .A1(G953), .A2(n667), .ZN(n551) );
  NAND2_X1 U571 ( .A1(n470), .A2(G902), .ZN(n549) );
  OR2_X1 U572 ( .A1(n721), .A2(n549), .ZN(n471) );
  NOR2_X1 U573 ( .A1(G900), .A2(n471), .ZN(n472) );
  NOR2_X1 U574 ( .A1(n551), .A2(n472), .ZN(n501) );
  NAND2_X1 U575 ( .A1(n473), .A2(G221), .ZN(n476) );
  XNOR2_X1 U576 ( .A(KEYINPUT95), .B(KEYINPUT21), .ZN(n474) );
  XNOR2_X1 U577 ( .A(n474), .B(KEYINPUT94), .ZN(n475) );
  XOR2_X1 U578 ( .A(n476), .B(n475), .Z(n650) );
  NOR2_X1 U579 ( .A1(n501), .A2(n650), .ZN(n477) );
  XNOR2_X1 U580 ( .A(n479), .B(n478), .ZN(n480) );
  XOR2_X1 U581 ( .A(n481), .B(n480), .Z(n484) );
  NAND2_X1 U582 ( .A1(n482), .A2(G210), .ZN(n483) );
  XNOR2_X1 U583 ( .A(n484), .B(n483), .ZN(n490) );
  XNOR2_X1 U584 ( .A(n491), .B(KEYINPUT28), .ZN(n499) );
  XNOR2_X1 U585 ( .A(n493), .B(n492), .ZN(n494) );
  XOR2_X1 U586 ( .A(G140), .B(n494), .Z(n496) );
  NAND2_X1 U587 ( .A1(G227), .A2(n721), .ZN(n495) );
  XNOR2_X1 U588 ( .A(n496), .B(n495), .ZN(n497) );
  XNOR2_X1 U589 ( .A(KEYINPUT72), .B(G469), .ZN(n498) );
  NAND2_X1 U590 ( .A1(n499), .A2(n507), .ZN(n518) );
  NAND2_X1 U591 ( .A1(n567), .A2(n638), .ZN(n500) );
  INV_X1 U592 ( .A(n507), .ZN(n502) );
  INV_X1 U593 ( .A(n650), .ZN(n555) );
  INV_X1 U594 ( .A(n651), .ZN(n568) );
  NAND2_X1 U595 ( .A1(n555), .A2(n568), .ZN(n647) );
  NOR2_X1 U596 ( .A1(n502), .A2(n647), .ZN(n584) );
  INV_X1 U597 ( .A(n639), .ZN(n503) );
  XNOR2_X1 U598 ( .A(n525), .B(KEYINPUT101), .ZN(n519) );
  NOR2_X1 U599 ( .A1(n526), .A2(n519), .ZN(n520) );
  BUF_X1 U600 ( .A(n520), .Z(n623) );
  XNOR2_X1 U601 ( .A(n506), .B(KEYINPUT46), .ZN(n517) );
  NAND2_X1 U602 ( .A1(n520), .A2(n576), .ZN(n512) );
  NOR2_X1 U603 ( .A1(n512), .A2(n511), .ZN(n539) );
  AND2_X1 U604 ( .A1(n528), .A2(n638), .ZN(n513) );
  AND2_X1 U605 ( .A1(n539), .A2(n513), .ZN(n514) );
  XOR2_X1 U606 ( .A(KEYINPUT36), .B(n514), .Z(n515) );
  NOR2_X1 U607 ( .A1(n648), .A2(n515), .ZN(n630) );
  XNOR2_X1 U608 ( .A(KEYINPUT84), .B(n630), .ZN(n516) );
  NOR2_X1 U609 ( .A1(n517), .A2(n516), .ZN(n535) );
  NOR2_X1 U610 ( .A1(n518), .A2(n552), .ZN(n621) );
  INV_X1 U611 ( .A(n621), .ZN(n523) );
  NOR2_X1 U612 ( .A1(n520), .A2(n627), .ZN(n643) );
  XOR2_X1 U613 ( .A(n643), .B(KEYINPUT81), .Z(n588) );
  NOR2_X1 U614 ( .A1(KEYINPUT47), .A2(n588), .ZN(n521) );
  XOR2_X1 U615 ( .A(KEYINPUT76), .B(n521), .Z(n522) );
  NOR2_X1 U616 ( .A1(n523), .A2(n522), .ZN(n533) );
  OR2_X1 U617 ( .A1(n643), .A2(n523), .ZN(n524) );
  NAND2_X1 U618 ( .A1(n524), .A2(KEYINPUT47), .ZN(n531) );
  NAND2_X1 U619 ( .A1(n526), .A2(n525), .ZN(n579) );
  NOR2_X1 U620 ( .A1(n527), .A2(n579), .ZN(n529) );
  NAND2_X1 U621 ( .A1(n529), .A2(n528), .ZN(n530) );
  XNOR2_X1 U622 ( .A(n530), .B(KEYINPUT106), .ZN(n733) );
  NAND2_X1 U623 ( .A1(n531), .A2(n733), .ZN(n532) );
  NOR2_X1 U624 ( .A1(n533), .A2(n532), .ZN(n534) );
  NAND2_X1 U625 ( .A1(n535), .A2(n534), .ZN(n537) );
  NAND2_X1 U626 ( .A1(n627), .A2(n538), .ZN(n633) );
  INV_X1 U627 ( .A(n633), .ZN(n546) );
  NAND2_X1 U628 ( .A1(n539), .A2(n638), .ZN(n540) );
  XNOR2_X1 U629 ( .A(KEYINPUT105), .B(n540), .ZN(n541) );
  NAND2_X1 U630 ( .A1(n541), .A2(n648), .ZN(n542) );
  XNOR2_X1 U631 ( .A(n542), .B(KEYINPUT43), .ZN(n544) );
  NAND2_X1 U632 ( .A1(n544), .A2(n543), .ZN(n635) );
  INV_X1 U633 ( .A(n635), .ZN(n545) );
  NOR2_X1 U634 ( .A1(n546), .A2(n545), .ZN(n547) );
  AND2_X1 U635 ( .A1(n596), .A2(n547), .ZN(n720) );
  INV_X1 U636 ( .A(n648), .ZN(n558) );
  NOR2_X1 U637 ( .A1(G898), .A2(n721), .ZN(n548) );
  XNOR2_X1 U638 ( .A(KEYINPUT91), .B(n548), .ZN(n714) );
  NOR2_X1 U639 ( .A1(n549), .A2(n714), .ZN(n550) );
  NOR2_X1 U640 ( .A1(n551), .A2(n550), .ZN(n553) );
  XNOR2_X1 U641 ( .A(KEYINPUT67), .B(KEYINPUT22), .ZN(n556) );
  XNOR2_X1 U642 ( .A(n557), .B(n556), .ZN(n564) );
  NOR2_X1 U643 ( .A1(n558), .A2(n564), .ZN(n570) );
  NAND2_X1 U644 ( .A1(n560), .A2(n570), .ZN(n559) );
  NOR2_X1 U645 ( .A1(n651), .A2(n559), .ZN(n610) );
  INV_X1 U646 ( .A(n610), .ZN(n575) );
  NAND2_X1 U647 ( .A1(n651), .A2(n560), .ZN(n561) );
  XNOR2_X1 U648 ( .A(n562), .B(KEYINPUT79), .ZN(n563) );
  NOR2_X1 U649 ( .A1(n564), .A2(n563), .ZN(n566) );
  INV_X1 U650 ( .A(KEYINPUT32), .ZN(n565) );
  XNOR2_X1 U651 ( .A(n566), .B(n565), .ZN(n729) );
  NOR2_X1 U652 ( .A1(n657), .A2(n568), .ZN(n569) );
  NAND2_X1 U653 ( .A1(n570), .A2(n569), .ZN(n618) );
  NAND2_X1 U654 ( .A1(n729), .A2(n618), .ZN(n571) );
  INV_X1 U655 ( .A(KEYINPUT44), .ZN(n572) );
  INV_X1 U656 ( .A(KEYINPUT66), .ZN(n573) );
  AND2_X1 U657 ( .A1(n576), .A2(n580), .ZN(n577) );
  XNOR2_X2 U658 ( .A(n577), .B(KEYINPUT33), .ZN(n668) );
  INV_X1 U659 ( .A(n583), .ZN(n581) );
  NAND2_X1 U660 ( .A1(n728), .A2(KEYINPUT44), .ZN(n590) );
  NAND2_X1 U661 ( .A1(n657), .A2(n580), .ZN(n659) );
  NAND2_X1 U662 ( .A1(n584), .A2(n583), .ZN(n585) );
  NOR2_X1 U663 ( .A1(n657), .A2(n585), .ZN(n615) );
  NOR2_X1 U664 ( .A1(n628), .A2(n615), .ZN(n586) );
  XNOR2_X1 U665 ( .A(n586), .B(KEYINPUT98), .ZN(n587) );
  OR2_X1 U666 ( .A1(n588), .A2(n587), .ZN(n589) );
  NOR2_X1 U667 ( .A1(n728), .A2(KEYINPUT44), .ZN(n591) );
  NAND2_X1 U668 ( .A1(n592), .A2(n591), .ZN(n593) );
  XNOR2_X1 U669 ( .A(KEYINPUT45), .B(KEYINPUT64), .ZN(n594) );
  NAND2_X1 U670 ( .A1(KEYINPUT2), .A2(n633), .ZN(n597) );
  XOR2_X1 U671 ( .A(KEYINPUT80), .B(n597), .Z(n598) );
  XNOR2_X1 U672 ( .A(n600), .B(KEYINPUT77), .ZN(n637) );
  INV_X1 U673 ( .A(n637), .ZN(n601) );
  AND2_X2 U674 ( .A1(n410), .A2(n601), .ZN(n702) );
  NAND2_X1 U675 ( .A1(n702), .A2(G472), .ZN(n606) );
  XNOR2_X1 U676 ( .A(n602), .B(KEYINPUT108), .ZN(n604) );
  XNOR2_X1 U677 ( .A(KEYINPUT109), .B(KEYINPUT62), .ZN(n603) );
  XNOR2_X1 U678 ( .A(n606), .B(n605), .ZN(n608) );
  NOR2_X1 U679 ( .A1(G952), .A2(n721), .ZN(n607) );
  INV_X1 U680 ( .A(n706), .ZN(n695) );
  NAND2_X1 U681 ( .A1(n608), .A2(n695), .ZN(n609) );
  XNOR2_X1 U682 ( .A(n609), .B(KEYINPUT63), .ZN(G57) );
  XOR2_X1 U683 ( .A(G101), .B(n610), .Z(G3) );
  NAND2_X1 U684 ( .A1(n615), .A2(n623), .ZN(n611) );
  XNOR2_X1 U685 ( .A(n611), .B(G104), .ZN(G6) );
  XOR2_X1 U686 ( .A(KEYINPUT27), .B(KEYINPUT111), .Z(n613) );
  XNOR2_X1 U687 ( .A(G107), .B(KEYINPUT110), .ZN(n612) );
  XNOR2_X1 U688 ( .A(n613), .B(n612), .ZN(n614) );
  XOR2_X1 U689 ( .A(KEYINPUT26), .B(n614), .Z(n617) );
  NAND2_X1 U690 ( .A1(n615), .A2(n627), .ZN(n616) );
  XNOR2_X1 U691 ( .A(n617), .B(n616), .ZN(G9) );
  XNOR2_X1 U692 ( .A(G110), .B(n618), .ZN(G12) );
  XOR2_X1 U693 ( .A(G128), .B(KEYINPUT29), .Z(n620) );
  NAND2_X1 U694 ( .A1(n627), .A2(n621), .ZN(n619) );
  XNOR2_X1 U695 ( .A(n620), .B(n619), .ZN(G30) );
  NAND2_X1 U696 ( .A1(n621), .A2(n623), .ZN(n622) );
  XNOR2_X1 U697 ( .A(n622), .B(G146), .ZN(G48) );
  XOR2_X1 U698 ( .A(KEYINPUT112), .B(KEYINPUT113), .Z(n625) );
  NAND2_X1 U699 ( .A1(n628), .A2(n623), .ZN(n624) );
  XNOR2_X1 U700 ( .A(n625), .B(n624), .ZN(n626) );
  XNOR2_X1 U701 ( .A(G113), .B(n626), .ZN(G15) );
  NAND2_X1 U702 ( .A1(n628), .A2(n627), .ZN(n629) );
  XNOR2_X1 U703 ( .A(n629), .B(G116), .ZN(G18) );
  XNOR2_X1 U704 ( .A(n630), .B(KEYINPUT37), .ZN(n631) );
  XNOR2_X1 U705 ( .A(n631), .B(KEYINPUT114), .ZN(n632) );
  XNOR2_X1 U706 ( .A(G125), .B(n632), .ZN(G27) );
  XOR2_X1 U707 ( .A(G134), .B(n633), .Z(n634) );
  XNOR2_X1 U708 ( .A(n634), .B(KEYINPUT115), .ZN(G36) );
  XNOR2_X1 U709 ( .A(G140), .B(n635), .ZN(G42) );
  NOR2_X1 U710 ( .A1(KEYINPUT2), .A2(n359), .ZN(n636) );
  NOR2_X1 U711 ( .A1(n637), .A2(n636), .ZN(n675) );
  NOR2_X1 U712 ( .A1(n639), .A2(n638), .ZN(n640) );
  NOR2_X1 U713 ( .A1(n641), .A2(n640), .ZN(n645) );
  NOR2_X1 U714 ( .A1(n643), .A2(n642), .ZN(n644) );
  NOR2_X1 U715 ( .A1(n645), .A2(n644), .ZN(n646) );
  NOR2_X1 U716 ( .A1(n646), .A2(n668), .ZN(n664) );
  NAND2_X1 U717 ( .A1(n648), .A2(n647), .ZN(n649) );
  XNOR2_X1 U718 ( .A(KEYINPUT50), .B(n649), .ZN(n655) );
  XOR2_X1 U719 ( .A(KEYINPUT116), .B(KEYINPUT49), .Z(n653) );
  NAND2_X1 U720 ( .A1(n651), .A2(n650), .ZN(n652) );
  XNOR2_X1 U721 ( .A(n653), .B(n652), .ZN(n654) );
  NAND2_X1 U722 ( .A1(n655), .A2(n654), .ZN(n656) );
  NOR2_X1 U723 ( .A1(n657), .A2(n656), .ZN(n658) );
  XNOR2_X1 U724 ( .A(n658), .B(KEYINPUT117), .ZN(n660) );
  NAND2_X1 U725 ( .A1(n660), .A2(n659), .ZN(n661) );
  XNOR2_X1 U726 ( .A(KEYINPUT51), .B(n661), .ZN(n662) );
  NOR2_X1 U727 ( .A1(n669), .A2(n662), .ZN(n663) );
  NOR2_X1 U728 ( .A1(n664), .A2(n663), .ZN(n665) );
  XNOR2_X1 U729 ( .A(n665), .B(KEYINPUT52), .ZN(n666) );
  NOR2_X1 U730 ( .A1(n667), .A2(n666), .ZN(n672) );
  NOR2_X1 U731 ( .A1(n669), .A2(n668), .ZN(n670) );
  XNOR2_X1 U732 ( .A(n670), .B(KEYINPUT118), .ZN(n671) );
  NOR2_X1 U733 ( .A1(n672), .A2(n671), .ZN(n673) );
  XNOR2_X1 U734 ( .A(n673), .B(KEYINPUT119), .ZN(n674) );
  XNOR2_X1 U735 ( .A(n676), .B(KEYINPUT120), .ZN(n677) );
  XNOR2_X1 U736 ( .A(KEYINPUT53), .B(n678), .ZN(G75) );
  NAND2_X1 U737 ( .A1(n702), .A2(G210), .ZN(n682) );
  XOR2_X1 U738 ( .A(KEYINPUT54), .B(KEYINPUT55), .Z(n679) );
  XNOR2_X1 U739 ( .A(n680), .B(n679), .ZN(n681) );
  XNOR2_X1 U740 ( .A(n682), .B(n681), .ZN(n683) );
  NAND2_X1 U741 ( .A1(n683), .A2(n695), .ZN(n685) );
  XNOR2_X1 U742 ( .A(KEYINPUT56), .B(KEYINPUT121), .ZN(n684) );
  XNOR2_X1 U743 ( .A(n685), .B(n684), .ZN(G51) );
  NAND2_X1 U744 ( .A1(n702), .A2(G469), .ZN(n689) );
  XOR2_X1 U745 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n686) );
  NOR2_X1 U746 ( .A1(n706), .A2(n690), .ZN(G54) );
  NAND2_X1 U747 ( .A1(n702), .A2(G475), .ZN(n694) );
  XNOR2_X1 U748 ( .A(KEYINPUT59), .B(n691), .ZN(n692) );
  XNOR2_X1 U749 ( .A(n694), .B(n693), .ZN(n696) );
  NAND2_X1 U750 ( .A1(n696), .A2(n695), .ZN(n698) );
  XNOR2_X1 U751 ( .A(KEYINPUT60), .B(KEYINPUT69), .ZN(n697) );
  XNOR2_X1 U752 ( .A(n698), .B(n697), .ZN(G60) );
  NAND2_X1 U753 ( .A1(G478), .A2(n702), .ZN(n699) );
  XNOR2_X1 U754 ( .A(n700), .B(n699), .ZN(n701) );
  NOR2_X1 U755 ( .A1(n706), .A2(n701), .ZN(G63) );
  NAND2_X1 U756 ( .A1(G217), .A2(n702), .ZN(n703) );
  XNOR2_X1 U757 ( .A(n704), .B(n703), .ZN(n705) );
  NOR2_X1 U758 ( .A1(n706), .A2(n705), .ZN(G66) );
  XOR2_X1 U759 ( .A(KEYINPUT123), .B(KEYINPUT61), .Z(n708) );
  NAND2_X1 U760 ( .A1(G224), .A2(G953), .ZN(n707) );
  XNOR2_X1 U761 ( .A(n708), .B(n707), .ZN(n709) );
  NAND2_X1 U762 ( .A1(n709), .A2(G898), .ZN(n711) );
  NAND2_X1 U763 ( .A1(n711), .A2(n710), .ZN(n716) );
  XNOR2_X1 U764 ( .A(n712), .B(KEYINPUT124), .ZN(n713) );
  NAND2_X1 U765 ( .A1(n714), .A2(n713), .ZN(n715) );
  XOR2_X1 U766 ( .A(n716), .B(n715), .Z(G69) );
  XOR2_X1 U767 ( .A(n717), .B(KEYINPUT125), .Z(n718) );
  XOR2_X1 U768 ( .A(n719), .B(n718), .Z(n723) );
  XOR2_X1 U769 ( .A(n723), .B(n720), .Z(n722) );
  NAND2_X1 U770 ( .A1(n722), .A2(n721), .ZN(n727) );
  XNOR2_X1 U771 ( .A(G227), .B(n723), .ZN(n724) );
  NAND2_X1 U772 ( .A1(n724), .A2(G900), .ZN(n725) );
  NAND2_X1 U773 ( .A1(G953), .A2(n725), .ZN(n726) );
  NAND2_X1 U774 ( .A1(n727), .A2(n726), .ZN(G72) );
  XOR2_X1 U775 ( .A(n728), .B(G122), .Z(G24) );
  BUF_X1 U776 ( .A(n729), .Z(n730) );
  XNOR2_X1 U777 ( .A(G119), .B(n730), .ZN(n731) );
  XNOR2_X1 U778 ( .A(n731), .B(KEYINPUT126), .ZN(G21) );
  XNOR2_X1 U779 ( .A(G131), .B(n732), .ZN(G33) );
  XNOR2_X1 U780 ( .A(G143), .B(n733), .ZN(G45) );
  XNOR2_X1 U781 ( .A(G137), .B(n734), .ZN(G39) );
endmodule

