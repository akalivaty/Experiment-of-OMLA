//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 1 1 0 0 1 1 0 1 0 0 0 1 0 1 1 0 1 1 0 1 0 0 0 1 0 1 1 1 1 1 1 0 0 1 0 1 0 1 0 0 0 1 0 0 1 0 0 0 1 1 1 0 1 0 1 0 1 0 0 0 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:28:32 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n444, new_n448, new_n449, new_n451, new_n454, new_n455,
    new_n456, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n522, new_n523, new_n524, new_n525,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n531, new_n532,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n541, new_n542,
    new_n543, new_n544, new_n545, new_n546, new_n547, new_n548, new_n549,
    new_n550, new_n553, new_n554, new_n556, new_n557, new_n558, new_n559,
    new_n560, new_n561, new_n562, new_n563, new_n564, new_n565, new_n566,
    new_n567, new_n568, new_n569, new_n570, new_n571, new_n572, new_n573,
    new_n574, new_n575, new_n576, new_n577, new_n578, new_n579, new_n582,
    new_n583, new_n584, new_n586, new_n587, new_n588, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n620, new_n621, new_n624, new_n626,
    new_n627, new_n628, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1191, new_n1192, new_n1193, new_n1194, new_n1195, new_n1196,
    new_n1197, new_n1198, new_n1199, new_n1200, new_n1201;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  XNOR2_X1  g012(.A(KEYINPUT64), .B(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  XOR2_X1   g014(.A(KEYINPUT65), .B(G57), .Z(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  AND2_X1   g016(.A1(G2072), .A2(G2078), .ZN(new_n442));
  NAND3_X1  g017(.A1(new_n442), .A2(G2084), .A3(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(new_n444));
  XNOR2_X1  g019(.A(new_n444), .B(KEYINPUT66), .ZN(G259));
  BUF_X1    g020(.A(G452), .Z(G391));
  AND2_X1   g021(.A1(G94), .A2(G452), .ZN(G173));
  XNOR2_X1  g022(.A(KEYINPUT67), .B(KEYINPUT1), .ZN(new_n448));
  AND2_X1   g023(.A1(G7), .A2(G661), .ZN(new_n449));
  XNOR2_X1  g024(.A(new_n448), .B(new_n449), .ZN(G223));
  NAND2_X1  g025(.A1(new_n449), .A2(G567), .ZN(new_n451));
  XOR2_X1   g026(.A(new_n451), .B(KEYINPUT68), .Z(G234));
  NAND2_X1  g027(.A1(new_n449), .A2(G2106), .ZN(G217));
  NOR4_X1   g028(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n454));
  XOR2_X1   g029(.A(new_n454), .B(KEYINPUT2), .Z(new_n455));
  OR4_X1    g030(.A1(G238), .A2(G237), .A3(G236), .A4(G235), .ZN(new_n456));
  NOR2_X1   g031(.A1(new_n455), .A2(new_n456), .ZN(G325));
  INV_X1    g032(.A(G325), .ZN(G261));
  AOI22_X1  g033(.A1(new_n455), .A2(G2106), .B1(G567), .B2(new_n456), .ZN(G319));
  INV_X1    g034(.A(G2105), .ZN(new_n460));
  AND2_X1   g035(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n461));
  NOR2_X1   g036(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n462));
  OAI21_X1  g037(.A(KEYINPUT69), .B1(new_n461), .B2(new_n462), .ZN(new_n463));
  INV_X1    g038(.A(KEYINPUT3), .ZN(new_n464));
  INV_X1    g039(.A(G2104), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  INV_X1    g041(.A(KEYINPUT69), .ZN(new_n467));
  NAND2_X1  g042(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n468));
  NAND3_X1  g043(.A1(new_n466), .A2(new_n467), .A3(new_n468), .ZN(new_n469));
  NAND3_X1  g044(.A1(new_n463), .A2(new_n469), .A3(G125), .ZN(new_n470));
  NAND2_X1  g045(.A1(G113), .A2(G2104), .ZN(new_n471));
  XNOR2_X1  g046(.A(new_n471), .B(KEYINPUT70), .ZN(new_n472));
  AOI21_X1  g047(.A(new_n460), .B1(new_n470), .B2(new_n472), .ZN(new_n473));
  AOI21_X1  g048(.A(G2105), .B1(new_n466), .B2(new_n468), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n474), .A2(G137), .ZN(new_n475));
  NAND3_X1  g050(.A1(new_n460), .A2(G101), .A3(G2104), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  NOR2_X1   g052(.A1(new_n473), .A2(new_n477), .ZN(G160));
  OAI21_X1  g053(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n479));
  INV_X1    g054(.A(G112), .ZN(new_n480));
  AOI21_X1  g055(.A(new_n479), .B1(new_n480), .B2(G2105), .ZN(new_n481));
  AOI21_X1  g056(.A(new_n460), .B1(new_n466), .B2(new_n468), .ZN(new_n482));
  XNOR2_X1  g057(.A(new_n482), .B(KEYINPUT71), .ZN(new_n483));
  AND2_X1   g058(.A1(new_n483), .A2(G124), .ZN(new_n484));
  AOI211_X1 g059(.A(new_n481), .B(new_n484), .C1(G136), .C2(new_n474), .ZN(G162));
  INV_X1    g060(.A(G138), .ZN(new_n486));
  NOR3_X1   g061(.A1(new_n486), .A2(KEYINPUT4), .A3(G2105), .ZN(new_n487));
  NAND3_X1  g062(.A1(new_n463), .A2(new_n469), .A3(new_n487), .ZN(new_n488));
  OAI211_X1 g063(.A(G138), .B(new_n460), .C1(new_n461), .C2(new_n462), .ZN(new_n489));
  NAND2_X1  g064(.A1(new_n489), .A2(KEYINPUT4), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n488), .A2(new_n490), .ZN(new_n491));
  INV_X1    g066(.A(KEYINPUT72), .ZN(new_n492));
  NOR2_X1   g067(.A1(new_n460), .A2(G114), .ZN(new_n493));
  OAI21_X1  g068(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n494));
  OAI21_X1  g069(.A(new_n492), .B1(new_n493), .B2(new_n494), .ZN(new_n495));
  OR2_X1    g070(.A1(G102), .A2(G2105), .ZN(new_n496));
  INV_X1    g071(.A(G114), .ZN(new_n497));
  NAND2_X1  g072(.A1(new_n497), .A2(G2105), .ZN(new_n498));
  NAND4_X1  g073(.A1(new_n496), .A2(new_n498), .A3(KEYINPUT72), .A4(G2104), .ZN(new_n499));
  AOI22_X1  g074(.A1(new_n495), .A2(new_n499), .B1(new_n482), .B2(G126), .ZN(new_n500));
  NAND2_X1  g075(.A1(new_n491), .A2(new_n500), .ZN(new_n501));
  INV_X1    g076(.A(new_n501), .ZN(G164));
  NAND2_X1  g077(.A1(KEYINPUT73), .A2(KEYINPUT5), .ZN(new_n503));
  INV_X1    g078(.A(G543), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  NAND3_X1  g080(.A1(KEYINPUT73), .A2(KEYINPUT5), .A3(G543), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  AOI22_X1  g082(.A1(new_n507), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n508));
  INV_X1    g083(.A(G651), .ZN(new_n509));
  OR2_X1    g084(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  AND2_X1   g085(.A1(KEYINPUT6), .A2(G651), .ZN(new_n511));
  NOR2_X1   g086(.A1(KEYINPUT6), .A2(G651), .ZN(new_n512));
  OR2_X1    g087(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  NAND3_X1  g088(.A1(new_n513), .A2(G88), .A3(new_n507), .ZN(new_n514));
  INV_X1    g089(.A(KEYINPUT74), .ZN(new_n515));
  OAI211_X1 g090(.A(G50), .B(G543), .C1(new_n511), .C2(new_n512), .ZN(new_n516));
  NAND3_X1  g091(.A1(new_n514), .A2(new_n515), .A3(new_n516), .ZN(new_n517));
  INV_X1    g092(.A(new_n517), .ZN(new_n518));
  AOI21_X1  g093(.A(new_n515), .B1(new_n514), .B2(new_n516), .ZN(new_n519));
  OAI21_X1  g094(.A(new_n510), .B1(new_n518), .B2(new_n519), .ZN(new_n520));
  INV_X1    g095(.A(new_n520), .ZN(G166));
  INV_X1    g096(.A(new_n506), .ZN(new_n522));
  AOI21_X1  g097(.A(G543), .B1(KEYINPUT73), .B2(KEYINPUT5), .ZN(new_n523));
  OAI22_X1  g098(.A1(new_n522), .A2(new_n523), .B1(new_n511), .B2(new_n512), .ZN(new_n524));
  INV_X1    g099(.A(new_n524), .ZN(new_n525));
  AND2_X1   g100(.A1(new_n525), .A2(G89), .ZN(new_n526));
  NAND3_X1  g101(.A1(new_n507), .A2(G63), .A3(G651), .ZN(new_n527));
  NAND3_X1  g102(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n528));
  XNOR2_X1  g103(.A(new_n528), .B(KEYINPUT7), .ZN(new_n529));
  NAND2_X1  g104(.A1(new_n513), .A2(G543), .ZN(new_n530));
  INV_X1    g105(.A(G51), .ZN(new_n531));
  OAI211_X1 g106(.A(new_n527), .B(new_n529), .C1(new_n530), .C2(new_n531), .ZN(new_n532));
  OR2_X1    g107(.A1(new_n526), .A2(new_n532), .ZN(G286));
  INV_X1    g108(.A(G286), .ZN(G168));
  INV_X1    g109(.A(G52), .ZN(new_n535));
  INV_X1    g110(.A(G90), .ZN(new_n536));
  OAI22_X1  g111(.A1(new_n530), .A2(new_n535), .B1(new_n524), .B2(new_n536), .ZN(new_n537));
  AOI22_X1  g112(.A1(new_n507), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n538));
  NOR2_X1   g113(.A1(new_n538), .A2(new_n509), .ZN(new_n539));
  NOR2_X1   g114(.A1(new_n537), .A2(new_n539), .ZN(G171));
  NAND2_X1  g115(.A1(G68), .A2(G543), .ZN(new_n541));
  INV_X1    g116(.A(new_n507), .ZN(new_n542));
  INV_X1    g117(.A(G56), .ZN(new_n543));
  OAI21_X1  g118(.A(new_n541), .B1(new_n542), .B2(new_n543), .ZN(new_n544));
  AOI21_X1  g119(.A(new_n509), .B1(new_n544), .B2(KEYINPUT75), .ZN(new_n545));
  OAI21_X1  g120(.A(new_n545), .B1(KEYINPUT75), .B2(new_n544), .ZN(new_n546));
  INV_X1    g121(.A(new_n530), .ZN(new_n547));
  AOI22_X1  g122(.A1(new_n547), .A2(G43), .B1(new_n525), .B2(G81), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n546), .A2(new_n548), .ZN(new_n549));
  INV_X1    g124(.A(new_n549), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n550), .A2(G860), .ZN(G153));
  NAND4_X1  g126(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g127(.A1(G1), .A2(G3), .ZN(new_n553));
  XNOR2_X1  g128(.A(new_n553), .B(KEYINPUT8), .ZN(new_n554));
  NAND4_X1  g129(.A1(G319), .A2(G483), .A3(G661), .A4(new_n554), .ZN(G188));
  INV_X1    g130(.A(KEYINPUT76), .ZN(new_n556));
  NAND3_X1  g131(.A1(new_n513), .A2(G53), .A3(G543), .ZN(new_n557));
  INV_X1    g132(.A(KEYINPUT77), .ZN(new_n558));
  OAI21_X1  g133(.A(new_n556), .B1(new_n557), .B2(new_n558), .ZN(new_n559));
  OR2_X1    g134(.A1(new_n559), .A2(KEYINPUT9), .ZN(new_n560));
  OAI211_X1 g135(.A(new_n559), .B(KEYINPUT9), .C1(new_n556), .C2(new_n557), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n525), .A2(G91), .ZN(new_n562));
  NAND3_X1  g137(.A1(new_n560), .A2(new_n561), .A3(new_n562), .ZN(new_n563));
  INV_X1    g138(.A(new_n563), .ZN(new_n564));
  INV_X1    g139(.A(KEYINPUT80), .ZN(new_n565));
  NAND2_X1  g140(.A1(G78), .A2(G543), .ZN(new_n566));
  XNOR2_X1  g141(.A(new_n507), .B(KEYINPUT78), .ZN(new_n567));
  INV_X1    g142(.A(G65), .ZN(new_n568));
  OAI211_X1 g143(.A(KEYINPUT79), .B(new_n566), .C1(new_n567), .C2(new_n568), .ZN(new_n569));
  AND2_X1   g144(.A1(new_n569), .A2(G651), .ZN(new_n570));
  INV_X1    g145(.A(KEYINPUT79), .ZN(new_n571));
  NAND2_X1  g146(.A1(new_n542), .A2(KEYINPUT78), .ZN(new_n572));
  INV_X1    g147(.A(KEYINPUT78), .ZN(new_n573));
  NAND2_X1  g148(.A1(new_n507), .A2(new_n573), .ZN(new_n574));
  AOI21_X1  g149(.A(new_n568), .B1(new_n572), .B2(new_n574), .ZN(new_n575));
  INV_X1    g150(.A(new_n566), .ZN(new_n576));
  OAI21_X1  g151(.A(new_n571), .B1(new_n575), .B2(new_n576), .ZN(new_n577));
  AOI21_X1  g152(.A(new_n565), .B1(new_n570), .B2(new_n577), .ZN(new_n578));
  AND4_X1   g153(.A1(new_n565), .A2(new_n577), .A3(new_n569), .A4(G651), .ZN(new_n579));
  OAI21_X1  g154(.A(new_n564), .B1(new_n578), .B2(new_n579), .ZN(G299));
  INV_X1    g155(.A(G171), .ZN(G301));
  NAND2_X1  g156(.A1(new_n520), .A2(KEYINPUT81), .ZN(new_n582));
  INV_X1    g157(.A(KEYINPUT81), .ZN(new_n583));
  OAI211_X1 g158(.A(new_n583), .B(new_n510), .C1(new_n518), .C2(new_n519), .ZN(new_n584));
  AND2_X1   g159(.A1(new_n582), .A2(new_n584), .ZN(G303));
  NAND2_X1  g160(.A1(new_n547), .A2(G49), .ZN(new_n586));
  OAI21_X1  g161(.A(G651), .B1(new_n507), .B2(G74), .ZN(new_n587));
  NAND2_X1  g162(.A1(new_n525), .A2(G87), .ZN(new_n588));
  NAND3_X1  g163(.A1(new_n586), .A2(new_n587), .A3(new_n588), .ZN(G288));
  NAND2_X1  g164(.A1(new_n525), .A2(G86), .ZN(new_n590));
  INV_X1    g165(.A(G61), .ZN(new_n591));
  AOI21_X1  g166(.A(new_n591), .B1(new_n505), .B2(new_n506), .ZN(new_n592));
  NAND2_X1  g167(.A1(G73), .A2(G543), .ZN(new_n593));
  INV_X1    g168(.A(new_n593), .ZN(new_n594));
  OAI21_X1  g169(.A(G651), .B1(new_n592), .B2(new_n594), .ZN(new_n595));
  NAND3_X1  g170(.A1(new_n513), .A2(G48), .A3(G543), .ZN(new_n596));
  NAND3_X1  g171(.A1(new_n590), .A2(new_n595), .A3(new_n596), .ZN(G305));
  AND2_X1   g172(.A1(new_n525), .A2(G85), .ZN(new_n598));
  NAND2_X1  g173(.A1(G72), .A2(G543), .ZN(new_n599));
  INV_X1    g174(.A(G60), .ZN(new_n600));
  OAI21_X1  g175(.A(new_n599), .B1(new_n542), .B2(new_n600), .ZN(new_n601));
  AOI21_X1  g176(.A(KEYINPUT82), .B1(new_n601), .B2(G651), .ZN(new_n602));
  AOI211_X1 g177(.A(new_n598), .B(new_n602), .C1(G47), .C2(new_n547), .ZN(new_n603));
  NAND3_X1  g178(.A1(new_n601), .A2(KEYINPUT82), .A3(G651), .ZN(new_n604));
  NAND2_X1  g179(.A1(new_n603), .A2(new_n604), .ZN(G290));
  NAND2_X1  g180(.A1(G301), .A2(G868), .ZN(new_n606));
  INV_X1    g181(.A(G66), .ZN(new_n607));
  NOR2_X1   g182(.A1(new_n567), .A2(new_n607), .ZN(new_n608));
  AND2_X1   g183(.A1(G79), .A2(G543), .ZN(new_n609));
  OAI21_X1  g184(.A(G651), .B1(new_n608), .B2(new_n609), .ZN(new_n610));
  NAND3_X1  g185(.A1(new_n525), .A2(KEYINPUT10), .A3(G92), .ZN(new_n611));
  INV_X1    g186(.A(KEYINPUT10), .ZN(new_n612));
  INV_X1    g187(.A(G92), .ZN(new_n613));
  OAI21_X1  g188(.A(new_n612), .B1(new_n524), .B2(new_n613), .ZN(new_n614));
  AOI22_X1  g189(.A1(new_n611), .A2(new_n614), .B1(G54), .B2(new_n547), .ZN(new_n615));
  NAND2_X1  g190(.A1(new_n610), .A2(new_n615), .ZN(new_n616));
  INV_X1    g191(.A(new_n616), .ZN(new_n617));
  OAI21_X1  g192(.A(new_n606), .B1(new_n617), .B2(G868), .ZN(G284));
  OAI21_X1  g193(.A(new_n606), .B1(new_n617), .B2(G868), .ZN(G321));
  NAND2_X1  g194(.A1(G286), .A2(G868), .ZN(new_n620));
  INV_X1    g195(.A(G299), .ZN(new_n621));
  OAI21_X1  g196(.A(new_n620), .B1(new_n621), .B2(G868), .ZN(G297));
  OAI21_X1  g197(.A(new_n620), .B1(new_n621), .B2(G868), .ZN(G280));
  INV_X1    g198(.A(G559), .ZN(new_n624));
  OAI21_X1  g199(.A(new_n617), .B1(new_n624), .B2(G860), .ZN(G148));
  INV_X1    g200(.A(G868), .ZN(new_n626));
  NAND2_X1  g201(.A1(new_n549), .A2(new_n626), .ZN(new_n627));
  NOR2_X1   g202(.A1(new_n616), .A2(G559), .ZN(new_n628));
  OAI21_X1  g203(.A(new_n627), .B1(new_n628), .B2(new_n626), .ZN(G323));
  XNOR2_X1  g204(.A(G323), .B(KEYINPUT11), .ZN(G282));
  AND2_X1   g205(.A1(new_n463), .A2(new_n469), .ZN(new_n631));
  NAND3_X1  g206(.A1(new_n631), .A2(G2104), .A3(new_n460), .ZN(new_n632));
  XNOR2_X1  g207(.A(new_n632), .B(KEYINPUT12), .ZN(new_n633));
  XNOR2_X1  g208(.A(new_n633), .B(KEYINPUT13), .ZN(new_n634));
  INV_X1    g209(.A(G2100), .ZN(new_n635));
  OR2_X1    g210(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  NAND2_X1  g211(.A1(new_n634), .A2(new_n635), .ZN(new_n637));
  NAND2_X1  g212(.A1(new_n474), .A2(G135), .ZN(new_n638));
  NOR2_X1   g213(.A1(new_n460), .A2(G111), .ZN(new_n639));
  OAI21_X1  g214(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n640));
  INV_X1    g215(.A(KEYINPUT71), .ZN(new_n641));
  XNOR2_X1  g216(.A(new_n482), .B(new_n641), .ZN(new_n642));
  INV_X1    g217(.A(G123), .ZN(new_n643));
  OAI221_X1 g218(.A(new_n638), .B1(new_n639), .B2(new_n640), .C1(new_n642), .C2(new_n643), .ZN(new_n644));
  XOR2_X1   g219(.A(new_n644), .B(G2096), .Z(new_n645));
  NAND3_X1  g220(.A1(new_n636), .A2(new_n637), .A3(new_n645), .ZN(G156));
  XOR2_X1   g221(.A(G2451), .B(G2454), .Z(new_n647));
  XNOR2_X1  g222(.A(new_n647), .B(KEYINPUT16), .ZN(new_n648));
  XNOR2_X1  g223(.A(G1341), .B(G1348), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n648), .B(new_n649), .ZN(new_n650));
  INV_X1    g225(.A(KEYINPUT14), .ZN(new_n651));
  XNOR2_X1  g226(.A(G2427), .B(G2438), .ZN(new_n652));
  XNOR2_X1  g227(.A(new_n652), .B(G2430), .ZN(new_n653));
  XNOR2_X1  g228(.A(KEYINPUT15), .B(G2435), .ZN(new_n654));
  AOI21_X1  g229(.A(new_n651), .B1(new_n653), .B2(new_n654), .ZN(new_n655));
  OAI21_X1  g230(.A(new_n655), .B1(new_n654), .B2(new_n653), .ZN(new_n656));
  XOR2_X1   g231(.A(new_n650), .B(new_n656), .Z(new_n657));
  XNOR2_X1  g232(.A(G2443), .B(G2446), .ZN(new_n658));
  OR2_X1    g233(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  NAND2_X1  g234(.A1(new_n657), .A2(new_n658), .ZN(new_n660));
  AND3_X1   g235(.A1(new_n659), .A2(G14), .A3(new_n660), .ZN(G401));
  INV_X1    g236(.A(KEYINPUT18), .ZN(new_n662));
  XOR2_X1   g237(.A(G2084), .B(G2090), .Z(new_n663));
  XNOR2_X1  g238(.A(new_n663), .B(KEYINPUT83), .ZN(new_n664));
  XNOR2_X1  g239(.A(G2067), .B(G2678), .ZN(new_n665));
  NAND2_X1  g240(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  NAND2_X1  g241(.A1(new_n666), .A2(KEYINPUT17), .ZN(new_n667));
  NOR2_X1   g242(.A1(new_n664), .A2(new_n665), .ZN(new_n668));
  OAI21_X1  g243(.A(new_n662), .B1(new_n667), .B2(new_n668), .ZN(new_n669));
  XOR2_X1   g244(.A(KEYINPUT84), .B(G2100), .Z(new_n670));
  XOR2_X1   g245(.A(new_n669), .B(new_n670), .Z(new_n671));
  NOR2_X1   g246(.A1(G2072), .A2(G2078), .ZN(new_n672));
  NOR2_X1   g247(.A1(new_n442), .A2(new_n672), .ZN(new_n673));
  AOI21_X1  g248(.A(new_n673), .B1(new_n666), .B2(KEYINPUT18), .ZN(new_n674));
  XOR2_X1   g249(.A(new_n674), .B(G2096), .Z(new_n675));
  XNOR2_X1  g250(.A(new_n671), .B(new_n675), .ZN(G227));
  XNOR2_X1  g251(.A(G1956), .B(G2474), .ZN(new_n677));
  INV_X1    g252(.A(KEYINPUT85), .ZN(new_n678));
  XNOR2_X1  g253(.A(new_n677), .B(new_n678), .ZN(new_n679));
  XOR2_X1   g254(.A(G1961), .B(G1966), .Z(new_n680));
  OR2_X1    g255(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  XNOR2_X1  g256(.A(G1971), .B(G1976), .ZN(new_n682));
  XNOR2_X1  g257(.A(new_n682), .B(KEYINPUT19), .ZN(new_n683));
  NAND2_X1  g258(.A1(new_n679), .A2(new_n680), .ZN(new_n684));
  NAND3_X1  g259(.A1(new_n681), .A2(new_n683), .A3(new_n684), .ZN(new_n685));
  NOR2_X1   g260(.A1(new_n684), .A2(new_n683), .ZN(new_n686));
  INV_X1    g261(.A(KEYINPUT20), .ZN(new_n687));
  NOR2_X1   g262(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  NOR3_X1   g263(.A1(new_n684), .A2(KEYINPUT20), .A3(new_n683), .ZN(new_n689));
  OAI221_X1 g264(.A(new_n685), .B1(new_n683), .B2(new_n681), .C1(new_n688), .C2(new_n689), .ZN(new_n690));
  XNOR2_X1  g265(.A(new_n690), .B(KEYINPUT86), .ZN(new_n691));
  XNOR2_X1  g266(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n692));
  XNOR2_X1  g267(.A(new_n691), .B(new_n692), .ZN(new_n693));
  XNOR2_X1  g268(.A(G1991), .B(G1996), .ZN(new_n694));
  XNOR2_X1  g269(.A(new_n693), .B(new_n694), .ZN(new_n695));
  XNOR2_X1  g270(.A(G1981), .B(G1986), .ZN(new_n696));
  XNOR2_X1  g271(.A(new_n695), .B(new_n696), .ZN(new_n697));
  INV_X1    g272(.A(new_n697), .ZN(G229));
  NAND2_X1  g273(.A1(new_n483), .A2(G129), .ZN(new_n699));
  NAND2_X1  g274(.A1(new_n474), .A2(G141), .ZN(new_n700));
  NAND3_X1  g275(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n701));
  XOR2_X1   g276(.A(new_n701), .B(KEYINPUT26), .Z(new_n702));
  NAND3_X1  g277(.A1(new_n460), .A2(G105), .A3(G2104), .ZN(new_n703));
  NAND4_X1  g278(.A1(new_n699), .A2(new_n700), .A3(new_n702), .A4(new_n703), .ZN(new_n704));
  MUX2_X1   g279(.A(G32), .B(new_n704), .S(G29), .Z(new_n705));
  XOR2_X1   g280(.A(KEYINPUT27), .B(G1996), .Z(new_n706));
  INV_X1    g281(.A(G16), .ZN(new_n707));
  NAND2_X1  g282(.A1(new_n707), .A2(G5), .ZN(new_n708));
  OAI21_X1  g283(.A(new_n708), .B1(G171), .B2(new_n707), .ZN(new_n709));
  AOI22_X1  g284(.A1(new_n705), .A2(new_n706), .B1(G1961), .B2(new_n709), .ZN(new_n710));
  INV_X1    g285(.A(G2067), .ZN(new_n711));
  INV_X1    g286(.A(G29), .ZN(new_n712));
  AND3_X1   g287(.A1(new_n712), .A2(KEYINPUT28), .A3(G26), .ZN(new_n713));
  AOI21_X1  g288(.A(KEYINPUT28), .B1(new_n712), .B2(G26), .ZN(new_n714));
  NAND2_X1  g289(.A1(new_n474), .A2(G140), .ZN(new_n715));
  NOR2_X1   g290(.A1(new_n460), .A2(G116), .ZN(new_n716));
  OAI21_X1  g291(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n717));
  INV_X1    g292(.A(G128), .ZN(new_n718));
  OAI221_X1 g293(.A(new_n715), .B1(new_n716), .B2(new_n717), .C1(new_n642), .C2(new_n718), .ZN(new_n719));
  AOI211_X1 g294(.A(new_n713), .B(new_n714), .C1(new_n719), .C2(G29), .ZN(new_n720));
  INV_X1    g295(.A(G2078), .ZN(new_n721));
  NAND2_X1  g296(.A1(G164), .A2(G29), .ZN(new_n722));
  OAI21_X1  g297(.A(new_n722), .B1(G27), .B2(G29), .ZN(new_n723));
  OAI221_X1 g298(.A(new_n710), .B1(new_n711), .B2(new_n720), .C1(new_n721), .C2(new_n723), .ZN(new_n724));
  NAND2_X1  g299(.A1(new_n707), .A2(G21), .ZN(new_n725));
  OAI21_X1  g300(.A(new_n725), .B1(G168), .B2(new_n707), .ZN(new_n726));
  XNOR2_X1  g301(.A(new_n726), .B(G1966), .ZN(new_n727));
  XOR2_X1   g302(.A(KEYINPUT31), .B(G11), .Z(new_n728));
  XNOR2_X1  g303(.A(new_n728), .B(KEYINPUT93), .ZN(new_n729));
  INV_X1    g304(.A(G28), .ZN(new_n730));
  OR2_X1    g305(.A1(new_n730), .A2(KEYINPUT30), .ZN(new_n731));
  AOI21_X1  g306(.A(G29), .B1(new_n730), .B2(KEYINPUT30), .ZN(new_n732));
  AOI21_X1  g307(.A(new_n729), .B1(new_n731), .B2(new_n732), .ZN(new_n733));
  OAI221_X1 g308(.A(new_n733), .B1(new_n644), .B2(new_n712), .C1(new_n709), .C2(G1961), .ZN(new_n734));
  OR3_X1    g309(.A1(new_n724), .A2(new_n727), .A3(new_n734), .ZN(new_n735));
  NAND2_X1  g310(.A1(new_n712), .A2(G33), .ZN(new_n736));
  NAND3_X1  g311(.A1(new_n460), .A2(G103), .A3(G2104), .ZN(new_n737));
  XNOR2_X1  g312(.A(new_n737), .B(KEYINPUT25), .ZN(new_n738));
  AOI22_X1  g313(.A1(new_n631), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n739));
  NOR2_X1   g314(.A1(new_n739), .A2(new_n460), .ZN(new_n740));
  AOI211_X1 g315(.A(new_n738), .B(new_n740), .C1(G139), .C2(new_n474), .ZN(new_n741));
  OAI21_X1  g316(.A(new_n736), .B1(new_n741), .B2(new_n712), .ZN(new_n742));
  OR2_X1    g317(.A1(new_n742), .A2(G2072), .ZN(new_n743));
  INV_X1    g318(.A(KEYINPUT24), .ZN(new_n744));
  OAI21_X1  g319(.A(new_n712), .B1(new_n744), .B2(G34), .ZN(new_n745));
  AOI21_X1  g320(.A(new_n745), .B1(new_n744), .B2(G34), .ZN(new_n746));
  AOI21_X1  g321(.A(new_n746), .B1(G160), .B2(G29), .ZN(new_n747));
  AOI22_X1  g322(.A1(new_n742), .A2(G2072), .B1(G2084), .B2(new_n747), .ZN(new_n748));
  OR2_X1    g323(.A1(new_n747), .A2(G2084), .ZN(new_n749));
  NAND3_X1  g324(.A1(new_n743), .A2(new_n748), .A3(new_n749), .ZN(new_n750));
  NAND2_X1  g325(.A1(new_n707), .A2(G19), .ZN(new_n751));
  XNOR2_X1  g326(.A(new_n751), .B(KEYINPUT92), .ZN(new_n752));
  OAI21_X1  g327(.A(new_n752), .B1(new_n550), .B2(new_n707), .ZN(new_n753));
  XNOR2_X1  g328(.A(new_n753), .B(G1341), .ZN(new_n754));
  NAND2_X1  g329(.A1(new_n707), .A2(G4), .ZN(new_n755));
  OAI21_X1  g330(.A(new_n755), .B1(new_n617), .B2(new_n707), .ZN(new_n756));
  XOR2_X1   g331(.A(KEYINPUT91), .B(G1348), .Z(new_n757));
  XOR2_X1   g332(.A(new_n756), .B(new_n757), .Z(new_n758));
  NOR4_X1   g333(.A1(new_n735), .A2(new_n750), .A3(new_n754), .A4(new_n758), .ZN(new_n759));
  NAND2_X1  g334(.A1(new_n707), .A2(G20), .ZN(new_n760));
  XNOR2_X1  g335(.A(new_n760), .B(KEYINPUT94), .ZN(new_n761));
  XNOR2_X1  g336(.A(new_n761), .B(KEYINPUT23), .ZN(new_n762));
  OAI21_X1  g337(.A(new_n762), .B1(new_n621), .B2(new_n707), .ZN(new_n763));
  XOR2_X1   g338(.A(KEYINPUT95), .B(G1956), .Z(new_n764));
  XNOR2_X1  g339(.A(new_n763), .B(new_n764), .ZN(new_n765));
  NAND2_X1  g340(.A1(new_n712), .A2(G35), .ZN(new_n766));
  OAI21_X1  g341(.A(new_n766), .B1(G162), .B2(new_n712), .ZN(new_n767));
  XOR2_X1   g342(.A(new_n767), .B(KEYINPUT29), .Z(new_n768));
  INV_X1    g343(.A(G2090), .ZN(new_n769));
  NAND2_X1  g344(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  NOR2_X1   g345(.A1(new_n768), .A2(new_n769), .ZN(new_n771));
  AOI22_X1  g346(.A1(new_n720), .A2(new_n711), .B1(new_n721), .B2(new_n723), .ZN(new_n772));
  OAI21_X1  g347(.A(new_n772), .B1(new_n705), .B2(new_n706), .ZN(new_n773));
  NOR2_X1   g348(.A1(new_n771), .A2(new_n773), .ZN(new_n774));
  NAND4_X1  g349(.A1(new_n759), .A2(new_n765), .A3(new_n770), .A4(new_n774), .ZN(new_n775));
  XNOR2_X1  g350(.A(new_n775), .B(KEYINPUT96), .ZN(new_n776));
  NAND2_X1  g351(.A1(new_n707), .A2(G23), .ZN(new_n777));
  INV_X1    g352(.A(G288), .ZN(new_n778));
  OAI21_X1  g353(.A(new_n777), .B1(new_n778), .B2(new_n707), .ZN(new_n779));
  XNOR2_X1  g354(.A(new_n779), .B(KEYINPUT33), .ZN(new_n780));
  INV_X1    g355(.A(G1976), .ZN(new_n781));
  XNOR2_X1  g356(.A(new_n780), .B(new_n781), .ZN(new_n782));
  MUX2_X1   g357(.A(G6), .B(G305), .S(G16), .Z(new_n783));
  XOR2_X1   g358(.A(KEYINPUT32), .B(G1981), .Z(new_n784));
  XNOR2_X1  g359(.A(new_n784), .B(KEYINPUT89), .ZN(new_n785));
  XNOR2_X1  g360(.A(new_n783), .B(new_n785), .ZN(new_n786));
  XNOR2_X1  g361(.A(new_n786), .B(KEYINPUT90), .ZN(new_n787));
  NOR2_X1   g362(.A1(G16), .A2(G22), .ZN(new_n788));
  AOI21_X1  g363(.A(new_n788), .B1(G166), .B2(G16), .ZN(new_n789));
  XNOR2_X1  g364(.A(new_n789), .B(G1971), .ZN(new_n790));
  NOR3_X1   g365(.A1(new_n782), .A2(new_n787), .A3(new_n790), .ZN(new_n791));
  INV_X1    g366(.A(KEYINPUT34), .ZN(new_n792));
  OR2_X1    g367(.A1(new_n791), .A2(new_n792), .ZN(new_n793));
  NAND2_X1  g368(.A1(new_n791), .A2(new_n792), .ZN(new_n794));
  INV_X1    g369(.A(G25), .ZN(new_n795));
  OR3_X1    g370(.A1(new_n795), .A2(KEYINPUT87), .A3(G29), .ZN(new_n796));
  OAI21_X1  g371(.A(KEYINPUT87), .B1(new_n795), .B2(G29), .ZN(new_n797));
  NAND2_X1  g372(.A1(new_n483), .A2(G119), .ZN(new_n798));
  OAI21_X1  g373(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n799));
  INV_X1    g374(.A(G107), .ZN(new_n800));
  AOI21_X1  g375(.A(new_n799), .B1(new_n800), .B2(G2105), .ZN(new_n801));
  AOI21_X1  g376(.A(new_n801), .B1(new_n474), .B2(G131), .ZN(new_n802));
  NAND2_X1  g377(.A1(new_n798), .A2(new_n802), .ZN(new_n803));
  INV_X1    g378(.A(new_n803), .ZN(new_n804));
  OAI211_X1 g379(.A(new_n796), .B(new_n797), .C1(new_n804), .C2(new_n712), .ZN(new_n805));
  XOR2_X1   g380(.A(KEYINPUT35), .B(G1991), .Z(new_n806));
  XNOR2_X1  g381(.A(new_n805), .B(new_n806), .ZN(new_n807));
  NAND2_X1  g382(.A1(new_n707), .A2(G24), .ZN(new_n808));
  XNOR2_X1  g383(.A(new_n808), .B(KEYINPUT88), .ZN(new_n809));
  AOI21_X1  g384(.A(new_n809), .B1(G290), .B2(G16), .ZN(new_n810));
  XNOR2_X1  g385(.A(new_n810), .B(G1986), .ZN(new_n811));
  NAND4_X1  g386(.A1(new_n793), .A2(new_n794), .A3(new_n807), .A4(new_n811), .ZN(new_n812));
  XOR2_X1   g387(.A(new_n812), .B(KEYINPUT36), .Z(new_n813));
  NOR2_X1   g388(.A1(new_n776), .A2(new_n813), .ZN(G311));
  INV_X1    g389(.A(G311), .ZN(G150));
  INV_X1    g390(.A(G55), .ZN(new_n816));
  INV_X1    g391(.A(G93), .ZN(new_n817));
  OAI22_X1  g392(.A1(new_n530), .A2(new_n816), .B1(new_n524), .B2(new_n817), .ZN(new_n818));
  XNOR2_X1  g393(.A(new_n818), .B(KEYINPUT97), .ZN(new_n819));
  AOI22_X1  g394(.A1(new_n507), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n820));
  OR2_X1    g395(.A1(new_n820), .A2(new_n509), .ZN(new_n821));
  NAND2_X1  g396(.A1(new_n819), .A2(new_n821), .ZN(new_n822));
  NAND2_X1  g397(.A1(new_n822), .A2(G860), .ZN(new_n823));
  XOR2_X1   g398(.A(KEYINPUT99), .B(KEYINPUT37), .Z(new_n824));
  XNOR2_X1  g399(.A(new_n823), .B(new_n824), .ZN(new_n825));
  NAND2_X1  g400(.A1(new_n617), .A2(G559), .ZN(new_n826));
  XOR2_X1   g401(.A(new_n826), .B(KEYINPUT38), .Z(new_n827));
  INV_X1    g402(.A(KEYINPUT98), .ZN(new_n828));
  NAND3_X1  g403(.A1(new_n819), .A2(new_n828), .A3(new_n821), .ZN(new_n829));
  INV_X1    g404(.A(new_n829), .ZN(new_n830));
  AOI21_X1  g405(.A(new_n828), .B1(new_n819), .B2(new_n821), .ZN(new_n831));
  NOR2_X1   g406(.A1(new_n830), .A2(new_n831), .ZN(new_n832));
  NAND2_X1  g407(.A1(new_n832), .A2(new_n550), .ZN(new_n833));
  OAI21_X1  g408(.A(new_n549), .B1(new_n830), .B2(new_n831), .ZN(new_n834));
  NAND2_X1  g409(.A1(new_n833), .A2(new_n834), .ZN(new_n835));
  XNOR2_X1  g410(.A(new_n827), .B(new_n835), .ZN(new_n836));
  INV_X1    g411(.A(new_n836), .ZN(new_n837));
  AND2_X1   g412(.A1(new_n837), .A2(KEYINPUT39), .ZN(new_n838));
  INV_X1    g413(.A(G860), .ZN(new_n839));
  OAI21_X1  g414(.A(new_n839), .B1(new_n837), .B2(KEYINPUT39), .ZN(new_n840));
  OAI21_X1  g415(.A(new_n825), .B1(new_n838), .B2(new_n840), .ZN(G145));
  NAND2_X1  g416(.A1(new_n474), .A2(G142), .ZN(new_n842));
  NOR2_X1   g417(.A1(new_n460), .A2(G118), .ZN(new_n843));
  OAI21_X1  g418(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n844));
  OAI21_X1  g419(.A(new_n842), .B1(new_n843), .B2(new_n844), .ZN(new_n845));
  AOI21_X1  g420(.A(new_n845), .B1(new_n483), .B2(G130), .ZN(new_n846));
  XNOR2_X1  g421(.A(new_n633), .B(new_n846), .ZN(new_n847));
  XNOR2_X1  g422(.A(new_n847), .B(new_n804), .ZN(new_n848));
  OR2_X1    g423(.A1(new_n848), .A2(KEYINPUT100), .ZN(new_n849));
  NAND2_X1  g424(.A1(new_n848), .A2(KEYINPUT100), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n849), .A2(new_n850), .ZN(new_n851));
  XNOR2_X1  g426(.A(new_n704), .B(new_n501), .ZN(new_n852));
  XNOR2_X1  g427(.A(new_n852), .B(new_n719), .ZN(new_n853));
  XNOR2_X1  g428(.A(new_n853), .B(new_n741), .ZN(new_n854));
  XNOR2_X1  g429(.A(new_n851), .B(new_n854), .ZN(new_n855));
  XNOR2_X1  g430(.A(new_n644), .B(G160), .ZN(new_n856));
  XNOR2_X1  g431(.A(new_n856), .B(G162), .ZN(new_n857));
  NAND2_X1  g432(.A1(new_n855), .A2(new_n857), .ZN(new_n858));
  INV_X1    g433(.A(G37), .ZN(new_n859));
  INV_X1    g434(.A(new_n854), .ZN(new_n860));
  AOI21_X1  g435(.A(new_n857), .B1(new_n860), .B2(new_n848), .ZN(new_n861));
  INV_X1    g436(.A(new_n851), .ZN(new_n862));
  OAI21_X1  g437(.A(new_n861), .B1(new_n862), .B2(new_n860), .ZN(new_n863));
  NAND3_X1  g438(.A1(new_n858), .A2(new_n859), .A3(new_n863), .ZN(new_n864));
  XNOR2_X1  g439(.A(new_n864), .B(KEYINPUT40), .ZN(G395));
  XNOR2_X1  g440(.A(G290), .B(G166), .ZN(new_n866));
  XNOR2_X1  g441(.A(G288), .B(G305), .ZN(new_n867));
  XNOR2_X1  g442(.A(new_n866), .B(new_n867), .ZN(new_n868));
  INV_X1    g443(.A(KEYINPUT42), .ZN(new_n869));
  XOR2_X1   g444(.A(new_n835), .B(new_n628), .Z(new_n870));
  INV_X1    g445(.A(new_n870), .ZN(new_n871));
  NOR2_X1   g446(.A1(G299), .A2(new_n616), .ZN(new_n872));
  INV_X1    g447(.A(new_n872), .ZN(new_n873));
  NAND2_X1  g448(.A1(G299), .A2(new_n616), .ZN(new_n874));
  NAND2_X1  g449(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n871), .A2(new_n875), .ZN(new_n876));
  NAND3_X1  g451(.A1(new_n873), .A2(KEYINPUT41), .A3(new_n874), .ZN(new_n877));
  INV_X1    g452(.A(new_n877), .ZN(new_n878));
  INV_X1    g453(.A(KEYINPUT41), .ZN(new_n879));
  INV_X1    g454(.A(new_n874), .ZN(new_n880));
  OAI21_X1  g455(.A(new_n879), .B1(new_n880), .B2(new_n872), .ZN(new_n881));
  INV_X1    g456(.A(new_n881), .ZN(new_n882));
  OAI21_X1  g457(.A(new_n870), .B1(new_n878), .B2(new_n882), .ZN(new_n883));
  AOI21_X1  g458(.A(new_n869), .B1(new_n876), .B2(new_n883), .ZN(new_n884));
  INV_X1    g459(.A(new_n884), .ZN(new_n885));
  NAND3_X1  g460(.A1(new_n876), .A2(new_n869), .A3(new_n883), .ZN(new_n886));
  AOI21_X1  g461(.A(new_n868), .B1(new_n885), .B2(new_n886), .ZN(new_n887));
  INV_X1    g462(.A(new_n886), .ZN(new_n888));
  INV_X1    g463(.A(new_n868), .ZN(new_n889));
  NOR3_X1   g464(.A1(new_n888), .A2(new_n889), .A3(new_n884), .ZN(new_n890));
  OAI21_X1  g465(.A(G868), .B1(new_n887), .B2(new_n890), .ZN(new_n891));
  INV_X1    g466(.A(KEYINPUT101), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n822), .A2(new_n626), .ZN(new_n893));
  NAND3_X1  g468(.A1(new_n891), .A2(new_n892), .A3(new_n893), .ZN(new_n894));
  OAI21_X1  g469(.A(new_n889), .B1(new_n888), .B2(new_n884), .ZN(new_n895));
  NAND3_X1  g470(.A1(new_n885), .A2(new_n886), .A3(new_n868), .ZN(new_n896));
  AOI21_X1  g471(.A(new_n626), .B1(new_n895), .B2(new_n896), .ZN(new_n897));
  INV_X1    g472(.A(new_n893), .ZN(new_n898));
  OAI21_X1  g473(.A(KEYINPUT101), .B1(new_n897), .B2(new_n898), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n894), .A2(new_n899), .ZN(G295));
  NAND2_X1  g475(.A1(new_n891), .A2(new_n893), .ZN(G331));
  INV_X1    g476(.A(KEYINPUT44), .ZN(new_n902));
  XNOR2_X1  g477(.A(G301), .B(G286), .ZN(new_n903));
  INV_X1    g478(.A(new_n903), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n835), .A2(new_n904), .ZN(new_n905));
  NAND3_X1  g480(.A1(new_n833), .A2(new_n834), .A3(new_n903), .ZN(new_n906));
  NAND2_X1  g481(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  NAND3_X1  g482(.A1(new_n907), .A2(new_n881), .A3(new_n877), .ZN(new_n908));
  NAND4_X1  g483(.A1(new_n905), .A2(new_n874), .A3(new_n873), .A4(new_n906), .ZN(new_n909));
  AOI21_X1  g484(.A(new_n889), .B1(new_n908), .B2(new_n909), .ZN(new_n910));
  INV_X1    g485(.A(new_n910), .ZN(new_n911));
  NAND3_X1  g486(.A1(new_n911), .A2(KEYINPUT102), .A3(new_n859), .ZN(new_n912));
  NAND3_X1  g487(.A1(new_n908), .A2(new_n889), .A3(new_n909), .ZN(new_n913));
  INV_X1    g488(.A(KEYINPUT43), .ZN(new_n914));
  AND2_X1   g489(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  INV_X1    g490(.A(KEYINPUT102), .ZN(new_n916));
  OAI21_X1  g491(.A(new_n916), .B1(new_n910), .B2(G37), .ZN(new_n917));
  NAND3_X1  g492(.A1(new_n912), .A2(new_n915), .A3(new_n917), .ZN(new_n918));
  NOR2_X1   g493(.A1(new_n910), .A2(G37), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n919), .A2(new_n913), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n920), .A2(KEYINPUT43), .ZN(new_n921));
  AOI21_X1  g496(.A(new_n902), .B1(new_n918), .B2(new_n921), .ZN(new_n922));
  NAND3_X1  g497(.A1(new_n912), .A2(new_n913), .A3(new_n917), .ZN(new_n923));
  AOI22_X1  g498(.A1(new_n923), .A2(KEYINPUT43), .B1(new_n919), .B2(new_n915), .ZN(new_n924));
  AOI21_X1  g499(.A(new_n922), .B1(new_n902), .B2(new_n924), .ZN(G397));
  INV_X1    g500(.A(G1384), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n501), .A2(new_n926), .ZN(new_n927));
  INV_X1    g502(.A(KEYINPUT45), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  NAND2_X1  g504(.A1(G160), .A2(G40), .ZN(new_n930));
  NOR2_X1   g505(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  NAND3_X1  g506(.A1(new_n931), .A2(G1996), .A3(new_n704), .ZN(new_n932));
  XNOR2_X1  g507(.A(new_n932), .B(KEYINPUT103), .ZN(new_n933));
  XNOR2_X1  g508(.A(new_n719), .B(new_n711), .ZN(new_n934));
  INV_X1    g509(.A(new_n934), .ZN(new_n935));
  NOR2_X1   g510(.A1(new_n704), .A2(G1996), .ZN(new_n936));
  OAI21_X1  g511(.A(new_n931), .B1(new_n935), .B2(new_n936), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n933), .A2(new_n937), .ZN(new_n938));
  XOR2_X1   g513(.A(new_n803), .B(new_n806), .Z(new_n939));
  AOI21_X1  g514(.A(new_n938), .B1(new_n931), .B2(new_n939), .ZN(new_n940));
  AND2_X1   g515(.A1(G290), .A2(G1986), .ZN(new_n941));
  NOR2_X1   g516(.A1(G290), .A2(G1986), .ZN(new_n942));
  OAI21_X1  g517(.A(new_n931), .B1(new_n941), .B2(new_n942), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n940), .A2(new_n943), .ZN(new_n944));
  NAND4_X1  g519(.A1(G303), .A2(KEYINPUT107), .A3(KEYINPUT55), .A4(G8), .ZN(new_n945));
  INV_X1    g520(.A(KEYINPUT107), .ZN(new_n946));
  NAND3_X1  g521(.A1(new_n582), .A2(G8), .A3(new_n584), .ZN(new_n947));
  INV_X1    g522(.A(KEYINPUT55), .ZN(new_n948));
  OAI21_X1  g523(.A(new_n946), .B1(new_n947), .B2(new_n948), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n947), .A2(new_n948), .ZN(new_n950));
  NAND3_X1  g525(.A1(new_n945), .A2(new_n949), .A3(new_n950), .ZN(new_n951));
  INV_X1    g526(.A(G40), .ZN(new_n952));
  NOR3_X1   g527(.A1(new_n473), .A2(new_n952), .A3(new_n477), .ZN(new_n953));
  NAND3_X1  g528(.A1(new_n501), .A2(KEYINPUT45), .A3(new_n926), .ZN(new_n954));
  NAND3_X1  g529(.A1(new_n929), .A2(new_n953), .A3(new_n954), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n955), .A2(KEYINPUT104), .ZN(new_n956));
  INV_X1    g531(.A(KEYINPUT104), .ZN(new_n957));
  NAND4_X1  g532(.A1(new_n929), .A2(new_n957), .A3(new_n953), .A4(new_n954), .ZN(new_n958));
  XNOR2_X1  g533(.A(KEYINPUT105), .B(G1971), .ZN(new_n959));
  NAND3_X1  g534(.A1(new_n956), .A2(new_n958), .A3(new_n959), .ZN(new_n960));
  AOI21_X1  g535(.A(new_n930), .B1(KEYINPUT50), .B2(new_n927), .ZN(new_n961));
  INV_X1    g536(.A(KEYINPUT106), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n927), .A2(new_n962), .ZN(new_n963));
  INV_X1    g538(.A(KEYINPUT50), .ZN(new_n964));
  NAND3_X1  g539(.A1(new_n501), .A2(KEYINPUT106), .A3(new_n926), .ZN(new_n965));
  NAND3_X1  g540(.A1(new_n963), .A2(new_n964), .A3(new_n965), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n961), .A2(new_n966), .ZN(new_n967));
  OAI21_X1  g542(.A(new_n960), .B1(G2090), .B2(new_n967), .ZN(new_n968));
  AND3_X1   g543(.A1(new_n951), .A2(new_n968), .A3(G8), .ZN(new_n969));
  NAND3_X1  g544(.A1(new_n963), .A2(new_n953), .A3(new_n965), .ZN(new_n970));
  XNOR2_X1  g545(.A(KEYINPUT108), .B(G8), .ZN(new_n971));
  INV_X1    g546(.A(new_n971), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n778), .A2(G1976), .ZN(new_n973));
  NAND3_X1  g548(.A1(new_n970), .A2(new_n972), .A3(new_n973), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n974), .A2(KEYINPUT109), .ZN(new_n975));
  INV_X1    g550(.A(KEYINPUT109), .ZN(new_n976));
  NAND4_X1  g551(.A1(new_n970), .A2(new_n976), .A3(new_n972), .A4(new_n973), .ZN(new_n977));
  NAND3_X1  g552(.A1(new_n975), .A2(KEYINPUT52), .A3(new_n977), .ZN(new_n978));
  INV_X1    g553(.A(G86), .ZN(new_n979));
  OAI21_X1  g554(.A(new_n596), .B1(new_n524), .B2(new_n979), .ZN(new_n980));
  INV_X1    g555(.A(new_n595), .ZN(new_n981));
  OAI21_X1  g556(.A(G1981), .B1(new_n980), .B2(new_n981), .ZN(new_n982));
  INV_X1    g557(.A(G1981), .ZN(new_n983));
  NAND4_X1  g558(.A1(new_n590), .A2(new_n983), .A3(new_n595), .A4(new_n596), .ZN(new_n984));
  AND3_X1   g559(.A1(new_n982), .A2(new_n984), .A3(KEYINPUT49), .ZN(new_n985));
  AOI21_X1  g560(.A(KEYINPUT49), .B1(new_n982), .B2(new_n984), .ZN(new_n986));
  NOR2_X1   g561(.A1(new_n985), .A2(new_n986), .ZN(new_n987));
  NAND3_X1  g562(.A1(new_n987), .A2(new_n972), .A3(new_n970), .ZN(new_n988));
  AOI21_X1  g563(.A(KEYINPUT52), .B1(G288), .B2(new_n781), .ZN(new_n989));
  NAND4_X1  g564(.A1(new_n970), .A2(new_n972), .A3(new_n973), .A4(new_n989), .ZN(new_n990));
  AND2_X1   g565(.A1(new_n988), .A2(new_n990), .ZN(new_n991));
  NAND3_X1  g566(.A1(new_n969), .A2(new_n978), .A3(new_n991), .ZN(new_n992));
  NAND2_X1  g567(.A1(new_n970), .A2(new_n972), .ZN(new_n993));
  NAND2_X1  g568(.A1(new_n993), .A2(KEYINPUT110), .ZN(new_n994));
  OR2_X1    g569(.A1(new_n993), .A2(KEYINPUT110), .ZN(new_n995));
  AND3_X1   g570(.A1(new_n988), .A2(new_n781), .A3(new_n778), .ZN(new_n996));
  INV_X1    g571(.A(new_n984), .ZN(new_n997));
  OAI211_X1 g572(.A(new_n994), .B(new_n995), .C1(new_n996), .C2(new_n997), .ZN(new_n998));
  INV_X1    g573(.A(KEYINPUT62), .ZN(new_n999));
  INV_X1    g574(.A(G2084), .ZN(new_n1000));
  AND3_X1   g575(.A1(new_n961), .A2(new_n1000), .A3(new_n966), .ZN(new_n1001));
  AOI21_X1  g576(.A(KEYINPUT106), .B1(new_n501), .B2(new_n926), .ZN(new_n1002));
  AOI211_X1 g577(.A(new_n962), .B(G1384), .C1(new_n491), .C2(new_n500), .ZN(new_n1003));
  OAI21_X1  g578(.A(new_n928), .B1(new_n1002), .B2(new_n1003), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n954), .A2(new_n953), .ZN(new_n1005));
  INV_X1    g580(.A(new_n1005), .ZN(new_n1006));
  AOI21_X1  g581(.A(G1966), .B1(new_n1004), .B2(new_n1006), .ZN(new_n1007));
  OAI211_X1 g582(.A(G286), .B(new_n972), .C1(new_n1001), .C2(new_n1007), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n1008), .A2(KEYINPUT51), .ZN(new_n1009));
  NOR2_X1   g584(.A1(G168), .A2(new_n971), .ZN(new_n1010));
  INV_X1    g585(.A(G8), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n1004), .A2(new_n1006), .ZN(new_n1012));
  INV_X1    g587(.A(G1966), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n1012), .A2(new_n1013), .ZN(new_n1014));
  NAND3_X1  g589(.A1(new_n961), .A2(new_n966), .A3(new_n1000), .ZN(new_n1015));
  AOI21_X1  g590(.A(new_n1011), .B1(new_n1014), .B2(new_n1015), .ZN(new_n1016));
  AOI21_X1  g591(.A(new_n1010), .B1(new_n1016), .B2(KEYINPUT122), .ZN(new_n1017));
  OAI21_X1  g592(.A(G8), .B1(new_n1001), .B2(new_n1007), .ZN(new_n1018));
  INV_X1    g593(.A(KEYINPUT122), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n1018), .A2(new_n1019), .ZN(new_n1020));
  AOI21_X1  g595(.A(new_n1009), .B1(new_n1017), .B2(new_n1020), .ZN(new_n1021));
  AOI21_X1  g596(.A(new_n971), .B1(new_n1014), .B2(new_n1015), .ZN(new_n1022));
  NOR3_X1   g597(.A1(new_n1022), .A2(KEYINPUT51), .A3(new_n1010), .ZN(new_n1023));
  OAI21_X1  g598(.A(new_n999), .B1(new_n1021), .B2(new_n1023), .ZN(new_n1024));
  INV_X1    g599(.A(G1961), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n967), .A2(new_n1025), .ZN(new_n1026));
  AND2_X1   g601(.A1(new_n721), .A2(KEYINPUT53), .ZN(new_n1027));
  NAND3_X1  g602(.A1(new_n1004), .A2(new_n1006), .A3(new_n1027), .ZN(new_n1028));
  AOI21_X1  g603(.A(G2078), .B1(new_n956), .B2(new_n958), .ZN(new_n1029));
  OAI211_X1 g604(.A(new_n1026), .B(new_n1028), .C1(new_n1029), .C2(KEYINPUT53), .ZN(new_n1030));
  INV_X1    g605(.A(new_n1030), .ZN(new_n1031));
  NOR2_X1   g606(.A1(new_n1031), .A2(G301), .ZN(new_n1032));
  INV_X1    g607(.A(KEYINPUT51), .ZN(new_n1033));
  AOI21_X1  g608(.A(new_n1033), .B1(new_n1022), .B2(G286), .ZN(new_n1034));
  INV_X1    g609(.A(new_n1010), .ZN(new_n1035));
  OAI21_X1  g610(.A(new_n1035), .B1(new_n1018), .B2(new_n1019), .ZN(new_n1036));
  NOR2_X1   g611(.A1(new_n1016), .A2(KEYINPUT122), .ZN(new_n1037));
  OAI21_X1  g612(.A(new_n1034), .B1(new_n1036), .B2(new_n1037), .ZN(new_n1038));
  INV_X1    g613(.A(new_n1023), .ZN(new_n1039));
  NAND3_X1  g614(.A1(new_n1038), .A2(KEYINPUT62), .A3(new_n1039), .ZN(new_n1040));
  NAND3_X1  g615(.A1(new_n1024), .A2(new_n1032), .A3(new_n1040), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n991), .A2(new_n978), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n1042), .A2(KEYINPUT113), .ZN(new_n1043));
  INV_X1    g618(.A(KEYINPUT113), .ZN(new_n1044));
  NAND3_X1  g619(.A1(new_n991), .A2(new_n978), .A3(new_n1044), .ZN(new_n1045));
  AOI21_X1  g620(.A(new_n969), .B1(new_n1043), .B2(new_n1045), .ZN(new_n1046));
  NOR2_X1   g621(.A1(new_n1002), .A2(new_n1003), .ZN(new_n1047));
  OAI21_X1  g622(.A(new_n953), .B1(new_n1047), .B2(new_n964), .ZN(new_n1048));
  INV_X1    g623(.A(KEYINPUT111), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n1048), .A2(new_n1049), .ZN(new_n1050));
  NAND3_X1  g625(.A1(new_n501), .A2(new_n964), .A3(new_n926), .ZN(new_n1051));
  OAI211_X1 g626(.A(KEYINPUT111), .B(new_n953), .C1(new_n1047), .C2(new_n964), .ZN(new_n1052));
  NAND4_X1  g627(.A1(new_n1050), .A2(new_n769), .A3(new_n1051), .A4(new_n1052), .ZN(new_n1053));
  INV_X1    g628(.A(KEYINPUT112), .ZN(new_n1054));
  NAND3_X1  g629(.A1(new_n1053), .A2(new_n1054), .A3(new_n960), .ZN(new_n1055));
  INV_X1    g630(.A(new_n1055), .ZN(new_n1056));
  AOI21_X1  g631(.A(new_n1054), .B1(new_n1053), .B2(new_n960), .ZN(new_n1057));
  NOR3_X1   g632(.A1(new_n1056), .A2(new_n1057), .A3(new_n971), .ZN(new_n1058));
  OAI21_X1  g633(.A(new_n1046), .B1(new_n1058), .B2(new_n951), .ZN(new_n1059));
  OAI211_X1 g634(.A(new_n992), .B(new_n998), .C1(new_n1041), .C2(new_n1059), .ZN(new_n1060));
  INV_X1    g635(.A(G1956), .ZN(new_n1061));
  AND2_X1   g636(.A1(new_n1048), .A2(new_n1049), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n1052), .A2(new_n1051), .ZN(new_n1063));
  OAI21_X1  g638(.A(new_n1061), .B1(new_n1062), .B2(new_n1063), .ZN(new_n1064));
  XOR2_X1   g639(.A(KEYINPUT56), .B(G2072), .Z(new_n1065));
  OR2_X1    g640(.A1(new_n955), .A2(new_n1065), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n1064), .A2(new_n1066), .ZN(new_n1067));
  XNOR2_X1  g642(.A(KEYINPUT115), .B(KEYINPUT57), .ZN(new_n1068));
  OAI211_X1 g643(.A(new_n564), .B(new_n1068), .C1(new_n578), .C2(new_n579), .ZN(new_n1069));
  INV_X1    g644(.A(new_n1068), .ZN(new_n1070));
  NAND2_X1  g645(.A1(G299), .A2(new_n1070), .ZN(new_n1071));
  NAND3_X1  g646(.A1(new_n1067), .A2(new_n1069), .A3(new_n1071), .ZN(new_n1072));
  INV_X1    g647(.A(KEYINPUT118), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n967), .A2(new_n757), .ZN(new_n1074));
  INV_X1    g649(.A(KEYINPUT116), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n970), .A2(new_n1075), .ZN(new_n1076));
  NAND4_X1  g651(.A1(new_n963), .A2(KEYINPUT116), .A3(new_n953), .A4(new_n965), .ZN(new_n1077));
  AOI21_X1  g652(.A(G2067), .B1(new_n1076), .B2(new_n1077), .ZN(new_n1078));
  INV_X1    g653(.A(KEYINPUT117), .ZN(new_n1079));
  OAI21_X1  g654(.A(new_n1074), .B1(new_n1078), .B2(new_n1079), .ZN(new_n1080));
  AOI21_X1  g655(.A(KEYINPUT116), .B1(new_n1047), .B2(new_n953), .ZN(new_n1081));
  INV_X1    g656(.A(new_n1077), .ZN(new_n1082));
  OAI211_X1 g657(.A(new_n1079), .B(new_n711), .C1(new_n1081), .C2(new_n1082), .ZN(new_n1083));
  INV_X1    g658(.A(new_n1083), .ZN(new_n1084));
  OAI21_X1  g659(.A(new_n1073), .B1(new_n1080), .B2(new_n1084), .ZN(new_n1085));
  OAI21_X1  g660(.A(new_n711), .B1(new_n1081), .B2(new_n1082), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n1086), .A2(KEYINPUT117), .ZN(new_n1087));
  NAND4_X1  g662(.A1(new_n1087), .A2(KEYINPUT118), .A3(new_n1083), .A4(new_n1074), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n1085), .A2(new_n1088), .ZN(new_n1089));
  OAI21_X1  g664(.A(new_n1072), .B1(new_n1089), .B2(new_n616), .ZN(new_n1090));
  NAND2_X1  g665(.A1(new_n1071), .A2(new_n1069), .ZN(new_n1091));
  NAND3_X1  g666(.A1(new_n1091), .A2(new_n1064), .A3(new_n1066), .ZN(new_n1092));
  NAND2_X1  g667(.A1(new_n1090), .A2(new_n1092), .ZN(new_n1093));
  NOR2_X1   g668(.A1(new_n617), .A2(KEYINPUT121), .ZN(new_n1094));
  INV_X1    g669(.A(new_n1094), .ZN(new_n1095));
  INV_X1    g670(.A(KEYINPUT121), .ZN(new_n1096));
  OAI21_X1  g671(.A(KEYINPUT60), .B1(new_n616), .B2(new_n1096), .ZN(new_n1097));
  INV_X1    g672(.A(new_n1097), .ZN(new_n1098));
  AOI21_X1  g673(.A(new_n1095), .B1(new_n1089), .B2(new_n1098), .ZN(new_n1099));
  AOI211_X1 g674(.A(new_n1097), .B(new_n1094), .C1(new_n1085), .C2(new_n1088), .ZN(new_n1100));
  INV_X1    g675(.A(KEYINPUT60), .ZN(new_n1101));
  NAND3_X1  g676(.A1(new_n1085), .A2(new_n1101), .A3(new_n1088), .ZN(new_n1102));
  INV_X1    g677(.A(new_n1102), .ZN(new_n1103));
  NOR3_X1   g678(.A1(new_n1099), .A2(new_n1100), .A3(new_n1103), .ZN(new_n1104));
  NAND3_X1  g679(.A1(new_n1072), .A2(KEYINPUT61), .A3(new_n1092), .ZN(new_n1105));
  INV_X1    g680(.A(KEYINPUT61), .ZN(new_n1106));
  AND3_X1   g681(.A1(new_n1091), .A2(new_n1064), .A3(new_n1066), .ZN(new_n1107));
  AOI21_X1  g682(.A(new_n1091), .B1(new_n1064), .B2(new_n1066), .ZN(new_n1108));
  OAI21_X1  g683(.A(new_n1106), .B1(new_n1107), .B2(new_n1108), .ZN(new_n1109));
  XNOR2_X1  g684(.A(KEYINPUT119), .B(KEYINPUT58), .ZN(new_n1110));
  XNOR2_X1  g685(.A(new_n1110), .B(G1341), .ZN(new_n1111));
  NAND3_X1  g686(.A1(new_n1076), .A2(new_n1077), .A3(new_n1111), .ZN(new_n1112));
  INV_X1    g687(.A(KEYINPUT120), .ZN(new_n1113));
  OAI22_X1  g688(.A1(new_n1112), .A2(new_n1113), .B1(new_n955), .B2(G1996), .ZN(new_n1114));
  AND2_X1   g689(.A1(new_n1112), .A2(new_n1113), .ZN(new_n1115));
  OAI21_X1  g690(.A(new_n550), .B1(new_n1114), .B2(new_n1115), .ZN(new_n1116));
  INV_X1    g691(.A(KEYINPUT59), .ZN(new_n1117));
  OR2_X1    g692(.A1(new_n1116), .A2(new_n1117), .ZN(new_n1118));
  NAND2_X1  g693(.A1(new_n1116), .A2(new_n1117), .ZN(new_n1119));
  NAND4_X1  g694(.A1(new_n1105), .A2(new_n1109), .A3(new_n1118), .A4(new_n1119), .ZN(new_n1120));
  OAI21_X1  g695(.A(new_n1093), .B1(new_n1104), .B2(new_n1120), .ZN(new_n1121));
  INV_X1    g696(.A(KEYINPUT54), .ZN(new_n1122));
  INV_X1    g697(.A(KEYINPUT123), .ZN(new_n1123));
  AND3_X1   g698(.A1(new_n929), .A2(new_n1123), .A3(new_n953), .ZN(new_n1124));
  AOI21_X1  g699(.A(new_n1123), .B1(new_n929), .B2(new_n953), .ZN(new_n1125));
  OAI211_X1 g700(.A(new_n954), .B(new_n1027), .C1(new_n1124), .C2(new_n1125), .ZN(new_n1126));
  OAI211_X1 g701(.A(new_n1126), .B(new_n1026), .C1(new_n1029), .C2(KEYINPUT53), .ZN(new_n1127));
  NOR2_X1   g702(.A1(new_n1127), .A2(G171), .ZN(new_n1128));
  OAI21_X1  g703(.A(new_n1122), .B1(new_n1032), .B2(new_n1128), .ZN(new_n1129));
  NOR2_X1   g704(.A1(new_n1021), .A2(new_n1023), .ZN(new_n1130));
  NAND2_X1  g705(.A1(new_n1031), .A2(G301), .ZN(new_n1131));
  AOI21_X1  g706(.A(new_n1122), .B1(new_n1127), .B2(G171), .ZN(new_n1132));
  AND3_X1   g707(.A1(new_n1131), .A2(new_n1132), .A3(KEYINPUT124), .ZN(new_n1133));
  AOI21_X1  g708(.A(KEYINPUT124), .B1(new_n1131), .B2(new_n1132), .ZN(new_n1134));
  OAI211_X1 g709(.A(new_n1129), .B(new_n1130), .C1(new_n1133), .C2(new_n1134), .ZN(new_n1135));
  NOR2_X1   g710(.A1(new_n1135), .A2(new_n1059), .ZN(new_n1136));
  AOI21_X1  g711(.A(new_n1060), .B1(new_n1121), .B2(new_n1136), .ZN(new_n1137));
  INV_X1    g712(.A(new_n1022), .ZN(new_n1138));
  NOR2_X1   g713(.A1(new_n1138), .A2(G286), .ZN(new_n1139));
  OAI211_X1 g714(.A(new_n1046), .B(new_n1139), .C1(new_n1058), .C2(new_n951), .ZN(new_n1140));
  INV_X1    g715(.A(KEYINPUT63), .ZN(new_n1141));
  NAND2_X1  g716(.A1(new_n1140), .A2(new_n1141), .ZN(new_n1142));
  INV_X1    g717(.A(KEYINPUT114), .ZN(new_n1143));
  NAND2_X1  g718(.A1(new_n1142), .A2(new_n1143), .ZN(new_n1144));
  NAND3_X1  g719(.A1(new_n1140), .A2(KEYINPUT114), .A3(new_n1141), .ZN(new_n1145));
  INV_X1    g720(.A(new_n969), .ZN(new_n1146));
  NAND3_X1  g721(.A1(new_n1146), .A2(KEYINPUT63), .A3(new_n1139), .ZN(new_n1147));
  AND2_X1   g722(.A1(new_n968), .A2(G8), .ZN(new_n1148));
  OAI211_X1 g723(.A(new_n978), .B(new_n991), .C1(new_n1148), .C2(new_n951), .ZN(new_n1149));
  OAI211_X1 g724(.A(new_n1144), .B(new_n1145), .C1(new_n1147), .C2(new_n1149), .ZN(new_n1150));
  AOI21_X1  g725(.A(new_n944), .B1(new_n1137), .B2(new_n1150), .ZN(new_n1151));
  NAND2_X1  g726(.A1(new_n942), .A2(new_n931), .ZN(new_n1152));
  XNOR2_X1  g727(.A(new_n1152), .B(KEYINPUT48), .ZN(new_n1153));
  NAND2_X1  g728(.A1(new_n940), .A2(new_n1153), .ZN(new_n1154));
  AND4_X1   g729(.A1(new_n806), .A2(new_n933), .A3(new_n804), .A4(new_n937), .ZN(new_n1155));
  NOR2_X1   g730(.A1(new_n719), .A2(G2067), .ZN(new_n1156));
  OAI21_X1  g731(.A(new_n931), .B1(new_n1155), .B2(new_n1156), .ZN(new_n1157));
  NOR3_X1   g732(.A1(new_n929), .A2(new_n930), .A3(G1996), .ZN(new_n1158));
  XOR2_X1   g733(.A(new_n1158), .B(KEYINPUT46), .Z(new_n1159));
  OAI21_X1  g734(.A(new_n931), .B1(new_n935), .B2(new_n704), .ZN(new_n1160));
  NAND2_X1  g735(.A1(new_n1159), .A2(new_n1160), .ZN(new_n1161));
  XOR2_X1   g736(.A(KEYINPUT125), .B(KEYINPUT47), .Z(new_n1162));
  XNOR2_X1  g737(.A(new_n1161), .B(new_n1162), .ZN(new_n1163));
  NAND3_X1  g738(.A1(new_n1154), .A2(new_n1157), .A3(new_n1163), .ZN(new_n1164));
  OAI21_X1  g739(.A(KEYINPUT126), .B1(new_n1151), .B2(new_n1164), .ZN(new_n1165));
  INV_X1    g740(.A(new_n944), .ZN(new_n1166));
  NAND2_X1  g741(.A1(new_n992), .A2(new_n998), .ZN(new_n1167));
  INV_X1    g742(.A(new_n1041), .ZN(new_n1168));
  INV_X1    g743(.A(new_n1059), .ZN(new_n1169));
  AOI21_X1  g744(.A(new_n1167), .B1(new_n1168), .B2(new_n1169), .ZN(new_n1170));
  AND2_X1   g745(.A1(new_n1090), .A2(new_n1092), .ZN(new_n1171));
  AND4_X1   g746(.A1(new_n1105), .A2(new_n1109), .A3(new_n1118), .A4(new_n1119), .ZN(new_n1172));
  NAND2_X1  g747(.A1(new_n1089), .A2(new_n1098), .ZN(new_n1173));
  NAND2_X1  g748(.A1(new_n1173), .A2(new_n1094), .ZN(new_n1174));
  NAND3_X1  g749(.A1(new_n1089), .A2(new_n1098), .A3(new_n1095), .ZN(new_n1175));
  NAND3_X1  g750(.A1(new_n1174), .A2(new_n1102), .A3(new_n1175), .ZN(new_n1176));
  AOI21_X1  g751(.A(new_n1171), .B1(new_n1172), .B2(new_n1176), .ZN(new_n1177));
  AND2_X1   g752(.A1(new_n1130), .A2(new_n1129), .ZN(new_n1178));
  OAI211_X1 g753(.A(new_n1169), .B(new_n1178), .C1(new_n1134), .C2(new_n1133), .ZN(new_n1179));
  OAI21_X1  g754(.A(new_n1170), .B1(new_n1177), .B2(new_n1179), .ZN(new_n1180));
  INV_X1    g755(.A(new_n1145), .ZN(new_n1181));
  AOI21_X1  g756(.A(KEYINPUT114), .B1(new_n1140), .B2(new_n1141), .ZN(new_n1182));
  NOR2_X1   g757(.A1(new_n1147), .A2(new_n1149), .ZN(new_n1183));
  NOR3_X1   g758(.A1(new_n1181), .A2(new_n1182), .A3(new_n1183), .ZN(new_n1184));
  OAI21_X1  g759(.A(new_n1166), .B1(new_n1180), .B2(new_n1184), .ZN(new_n1185));
  INV_X1    g760(.A(KEYINPUT126), .ZN(new_n1186));
  INV_X1    g761(.A(new_n1164), .ZN(new_n1187));
  NAND3_X1  g762(.A1(new_n1185), .A2(new_n1186), .A3(new_n1187), .ZN(new_n1188));
  NAND2_X1  g763(.A1(new_n1165), .A2(new_n1188), .ZN(G329));
  assign    G231 = 1'b0;
  NAND2_X1  g764(.A1(new_n923), .A2(KEYINPUT43), .ZN(new_n1191));
  NAND2_X1  g765(.A1(new_n915), .A2(new_n919), .ZN(new_n1192));
  NAND2_X1  g766(.A1(new_n1191), .A2(new_n1192), .ZN(new_n1193));
  INV_X1    g767(.A(KEYINPUT127), .ZN(new_n1194));
  INV_X1    g768(.A(G401), .ZN(new_n1195));
  NAND2_X1  g769(.A1(new_n1195), .A2(G319), .ZN(new_n1196));
  NOR2_X1   g770(.A1(new_n1196), .A2(G227), .ZN(new_n1197));
  NAND3_X1  g771(.A1(new_n697), .A2(new_n864), .A3(new_n1197), .ZN(new_n1198));
  INV_X1    g772(.A(new_n1198), .ZN(new_n1199));
  NAND3_X1  g773(.A1(new_n1193), .A2(new_n1194), .A3(new_n1199), .ZN(new_n1200));
  OAI21_X1  g774(.A(KEYINPUT127), .B1(new_n924), .B2(new_n1198), .ZN(new_n1201));
  AND2_X1   g775(.A1(new_n1200), .A2(new_n1201), .ZN(G308));
  NAND2_X1  g776(.A1(new_n1200), .A2(new_n1201), .ZN(G225));
endmodule


