//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 1 1 1 1 0 0 1 1 1 1 0 0 0 1 1 0 1 1 1 1 0 0 0 0 0 0 1 1 0 1 0 1 1 1 1 0 1 1 0 0 1 1 1 0 0 0 1 1 0 0 1 1 0 0 0 1 1 0 1 0 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:23:07 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n709, new_n710,
    new_n711, new_n712, new_n713, new_n714, new_n715, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n728, new_n729, new_n731, new_n732, new_n733, new_n734,
    new_n736, new_n737, new_n738, new_n739, new_n740, new_n741, new_n742,
    new_n743, new_n744, new_n745, new_n746, new_n748, new_n749, new_n750,
    new_n751, new_n752, new_n753, new_n754, new_n755, new_n756, new_n757,
    new_n758, new_n759, new_n760, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n791, new_n792, new_n793, new_n794,
    new_n795, new_n796, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n821, new_n822, new_n823, new_n824,
    new_n825, new_n826, new_n827, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n964, new_n965, new_n966,
    new_n967, new_n968, new_n969, new_n970, new_n971, new_n972, new_n973,
    new_n974, new_n975, new_n976, new_n977, new_n978, new_n979, new_n980,
    new_n981, new_n982, new_n983, new_n984, new_n985, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1013, new_n1014, new_n1015, new_n1016,
    new_n1017, new_n1018, new_n1019, new_n1020, new_n1021, new_n1022,
    new_n1023, new_n1024, new_n1025, new_n1027, new_n1028, new_n1029,
    new_n1031, new_n1032, new_n1033, new_n1034, new_n1035, new_n1036,
    new_n1037, new_n1038, new_n1039, new_n1040, new_n1041, new_n1042,
    new_n1043, new_n1044, new_n1045, new_n1046, new_n1047, new_n1048,
    new_n1049, new_n1050, new_n1051, new_n1052, new_n1053, new_n1054,
    new_n1055, new_n1057, new_n1058, new_n1059, new_n1060, new_n1061,
    new_n1062, new_n1063, new_n1064, new_n1065, new_n1066, new_n1067,
    new_n1068, new_n1069, new_n1070, new_n1071, new_n1072, new_n1073;
  INV_X1    g000(.A(G472), .ZN(new_n187));
  INV_X1    g001(.A(KEYINPUT11), .ZN(new_n188));
  INV_X1    g002(.A(G134), .ZN(new_n189));
  OAI21_X1  g003(.A(new_n188), .B1(new_n189), .B2(G137), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n189), .A2(G137), .ZN(new_n191));
  INV_X1    g005(.A(G137), .ZN(new_n192));
  NAND3_X1  g006(.A1(new_n192), .A2(KEYINPUT11), .A3(G134), .ZN(new_n193));
  NAND3_X1  g007(.A1(new_n190), .A2(new_n191), .A3(new_n193), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n194), .A2(G131), .ZN(new_n195));
  INV_X1    g009(.A(G131), .ZN(new_n196));
  NAND4_X1  g010(.A1(new_n190), .A2(new_n193), .A3(new_n196), .A4(new_n191), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n195), .A2(new_n197), .ZN(new_n198));
  INV_X1    g012(.A(G146), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n199), .A2(G143), .ZN(new_n200));
  INV_X1    g014(.A(G143), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n201), .A2(G146), .ZN(new_n202));
  NAND4_X1  g016(.A1(new_n200), .A2(new_n202), .A3(KEYINPUT0), .A4(G128), .ZN(new_n203));
  INV_X1    g017(.A(KEYINPUT64), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  XNOR2_X1  g019(.A(G143), .B(G146), .ZN(new_n206));
  NAND4_X1  g020(.A1(new_n206), .A2(KEYINPUT64), .A3(KEYINPUT0), .A4(G128), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n205), .A2(new_n207), .ZN(new_n208));
  XNOR2_X1  g022(.A(KEYINPUT0), .B(G128), .ZN(new_n209));
  NOR2_X1   g023(.A1(new_n206), .A2(new_n209), .ZN(new_n210));
  INV_X1    g024(.A(new_n210), .ZN(new_n211));
  NAND3_X1  g025(.A1(new_n198), .A2(new_n208), .A3(new_n211), .ZN(new_n212));
  AND3_X1   g026(.A1(new_n200), .A2(new_n202), .A3(G128), .ZN(new_n213));
  INV_X1    g027(.A(KEYINPUT1), .ZN(new_n214));
  OAI21_X1  g028(.A(KEYINPUT1), .B1(new_n201), .B2(G146), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n215), .A2(G128), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n200), .A2(new_n202), .ZN(new_n217));
  AOI22_X1  g031(.A1(new_n213), .A2(new_n214), .B1(new_n216), .B2(new_n217), .ZN(new_n218));
  INV_X1    g032(.A(new_n191), .ZN(new_n219));
  NOR2_X1   g033(.A1(new_n189), .A2(G137), .ZN(new_n220));
  OAI21_X1  g034(.A(G131), .B1(new_n219), .B2(new_n220), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n221), .A2(new_n197), .ZN(new_n222));
  OAI21_X1  g036(.A(KEYINPUT65), .B1(new_n218), .B2(new_n222), .ZN(new_n223));
  NAND4_X1  g037(.A1(new_n200), .A2(new_n202), .A3(new_n214), .A4(G128), .ZN(new_n224));
  INV_X1    g038(.A(G128), .ZN(new_n225));
  AOI21_X1  g039(.A(new_n225), .B1(new_n200), .B2(KEYINPUT1), .ZN(new_n226));
  OAI21_X1  g040(.A(new_n224), .B1(new_n226), .B2(new_n206), .ZN(new_n227));
  INV_X1    g041(.A(KEYINPUT65), .ZN(new_n228));
  NAND4_X1  g042(.A1(new_n227), .A2(new_n228), .A3(new_n221), .A4(new_n197), .ZN(new_n229));
  NAND3_X1  g043(.A1(new_n212), .A2(new_n223), .A3(new_n229), .ZN(new_n230));
  INV_X1    g044(.A(KEYINPUT30), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n230), .A2(new_n231), .ZN(new_n232));
  INV_X1    g046(.A(KEYINPUT66), .ZN(new_n233));
  INV_X1    g047(.A(G116), .ZN(new_n234));
  OAI21_X1  g048(.A(new_n233), .B1(new_n234), .B2(G119), .ZN(new_n235));
  INV_X1    g049(.A(G119), .ZN(new_n236));
  NAND3_X1  g050(.A1(new_n236), .A2(KEYINPUT66), .A3(G116), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n234), .A2(G119), .ZN(new_n238));
  NAND3_X1  g052(.A1(new_n235), .A2(new_n237), .A3(new_n238), .ZN(new_n239));
  XNOR2_X1  g053(.A(KEYINPUT2), .B(G113), .ZN(new_n240));
  XNOR2_X1  g054(.A(new_n239), .B(new_n240), .ZN(new_n241));
  NAND3_X1  g055(.A1(new_n227), .A2(new_n221), .A3(new_n197), .ZN(new_n242));
  NAND3_X1  g056(.A1(new_n212), .A2(KEYINPUT30), .A3(new_n242), .ZN(new_n243));
  NAND3_X1  g057(.A1(new_n232), .A2(new_n241), .A3(new_n243), .ZN(new_n244));
  XOR2_X1   g058(.A(new_n239), .B(new_n240), .Z(new_n245));
  NAND3_X1  g059(.A1(new_n212), .A2(new_n245), .A3(new_n242), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n244), .A2(new_n246), .ZN(new_n247));
  OR2_X1    g061(.A1(KEYINPUT67), .A2(G953), .ZN(new_n248));
  INV_X1    g062(.A(G237), .ZN(new_n249));
  NAND2_X1  g063(.A1(KEYINPUT67), .A2(G953), .ZN(new_n250));
  NAND4_X1  g064(.A1(new_n248), .A2(G210), .A3(new_n249), .A4(new_n250), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n251), .A2(KEYINPUT69), .ZN(new_n252));
  AND2_X1   g066(.A1(KEYINPUT67), .A2(G953), .ZN(new_n253));
  NOR2_X1   g067(.A1(KEYINPUT67), .A2(G953), .ZN(new_n254));
  NOR2_X1   g068(.A1(new_n253), .A2(new_n254), .ZN(new_n255));
  INV_X1    g069(.A(KEYINPUT69), .ZN(new_n256));
  NAND4_X1  g070(.A1(new_n255), .A2(new_n256), .A3(G210), .A4(new_n249), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n252), .A2(new_n257), .ZN(new_n258));
  XNOR2_X1  g072(.A(KEYINPUT26), .B(G101), .ZN(new_n259));
  XNOR2_X1  g073(.A(KEYINPUT68), .B(KEYINPUT27), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  INV_X1    g075(.A(new_n261), .ZN(new_n262));
  NOR2_X1   g076(.A1(new_n259), .A2(new_n260), .ZN(new_n263));
  OAI21_X1  g077(.A(new_n258), .B1(new_n262), .B2(new_n263), .ZN(new_n264));
  OR2_X1    g078(.A1(new_n259), .A2(new_n260), .ZN(new_n265));
  NAND4_X1  g079(.A1(new_n265), .A2(new_n252), .A3(new_n257), .A4(new_n261), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n264), .A2(new_n266), .ZN(new_n267));
  INV_X1    g081(.A(new_n267), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n247), .A2(new_n268), .ZN(new_n269));
  INV_X1    g083(.A(KEYINPUT29), .ZN(new_n270));
  XNOR2_X1  g084(.A(new_n246), .B(KEYINPUT28), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n230), .A2(new_n241), .ZN(new_n272));
  NAND3_X1  g086(.A1(new_n271), .A2(new_n272), .A3(new_n267), .ZN(new_n273));
  NAND3_X1  g087(.A1(new_n269), .A2(new_n270), .A3(new_n273), .ZN(new_n274));
  INV_X1    g088(.A(KEYINPUT28), .ZN(new_n275));
  XNOR2_X1  g089(.A(new_n246), .B(new_n275), .ZN(new_n276));
  AOI21_X1  g090(.A(new_n245), .B1(new_n212), .B2(new_n242), .ZN(new_n277));
  NOR2_X1   g091(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  NOR2_X1   g092(.A1(new_n268), .A2(new_n270), .ZN(new_n279));
  AOI21_X1  g093(.A(G902), .B1(new_n278), .B2(new_n279), .ZN(new_n280));
  AOI21_X1  g094(.A(new_n187), .B1(new_n274), .B2(new_n280), .ZN(new_n281));
  INV_X1    g095(.A(new_n281), .ZN(new_n282));
  AOI21_X1  g096(.A(new_n267), .B1(new_n271), .B2(new_n272), .ZN(new_n283));
  INV_X1    g097(.A(KEYINPUT31), .ZN(new_n284));
  INV_X1    g098(.A(KEYINPUT70), .ZN(new_n285));
  NAND3_X1  g099(.A1(new_n246), .A2(new_n267), .A3(new_n285), .ZN(new_n286));
  INV_X1    g100(.A(new_n286), .ZN(new_n287));
  AOI21_X1  g101(.A(new_n285), .B1(new_n246), .B2(new_n267), .ZN(new_n288));
  NOR2_X1   g102(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  AND3_X1   g103(.A1(new_n232), .A2(new_n241), .A3(new_n243), .ZN(new_n290));
  OAI21_X1  g104(.A(new_n284), .B1(new_n289), .B2(new_n290), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n246), .A2(new_n267), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n292), .A2(KEYINPUT70), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n293), .A2(new_n286), .ZN(new_n294));
  NAND3_X1  g108(.A1(new_n294), .A2(KEYINPUT31), .A3(new_n244), .ZN(new_n295));
  AOI21_X1  g109(.A(new_n283), .B1(new_n291), .B2(new_n295), .ZN(new_n296));
  NOR2_X1   g110(.A1(G472), .A2(G902), .ZN(new_n297));
  INV_X1    g111(.A(new_n297), .ZN(new_n298));
  NOR3_X1   g112(.A1(new_n296), .A2(KEYINPUT32), .A3(new_n298), .ZN(new_n299));
  INV_X1    g113(.A(KEYINPUT32), .ZN(new_n300));
  INV_X1    g114(.A(new_n283), .ZN(new_n301));
  AND3_X1   g115(.A1(new_n294), .A2(KEYINPUT31), .A3(new_n244), .ZN(new_n302));
  AOI21_X1  g116(.A(KEYINPUT31), .B1(new_n294), .B2(new_n244), .ZN(new_n303));
  OAI21_X1  g117(.A(new_n301), .B1(new_n302), .B2(new_n303), .ZN(new_n304));
  AOI21_X1  g118(.A(new_n300), .B1(new_n304), .B2(new_n297), .ZN(new_n305));
  OAI21_X1  g119(.A(new_n282), .B1(new_n299), .B2(new_n305), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n306), .A2(KEYINPUT71), .ZN(new_n307));
  OAI21_X1  g121(.A(KEYINPUT32), .B1(new_n296), .B2(new_n298), .ZN(new_n308));
  NAND3_X1  g122(.A1(new_n304), .A2(new_n300), .A3(new_n297), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n308), .A2(new_n309), .ZN(new_n310));
  INV_X1    g124(.A(KEYINPUT71), .ZN(new_n311));
  NAND3_X1  g125(.A1(new_n310), .A2(new_n311), .A3(new_n282), .ZN(new_n312));
  INV_X1    g126(.A(G234), .ZN(new_n313));
  OAI21_X1  g127(.A(G217), .B1(new_n313), .B2(G902), .ZN(new_n314));
  INV_X1    g128(.A(KEYINPUT72), .ZN(new_n315));
  INV_X1    g129(.A(G125), .ZN(new_n316));
  NAND3_X1  g130(.A1(new_n315), .A2(new_n316), .A3(G140), .ZN(new_n317));
  INV_X1    g131(.A(G140), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n318), .A2(G125), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n316), .A2(G140), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  OAI211_X1 g135(.A(KEYINPUT16), .B(new_n317), .C1(new_n321), .C2(new_n315), .ZN(new_n322));
  INV_X1    g136(.A(KEYINPUT16), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n319), .A2(new_n323), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n322), .A2(new_n324), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n325), .A2(G146), .ZN(new_n326));
  NAND3_X1  g140(.A1(new_n322), .A2(new_n199), .A3(new_n324), .ZN(new_n327));
  NAND3_X1  g141(.A1(new_n326), .A2(KEYINPUT73), .A3(new_n327), .ZN(new_n328));
  INV_X1    g142(.A(KEYINPUT73), .ZN(new_n329));
  NAND3_X1  g143(.A1(new_n325), .A2(new_n329), .A3(G146), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n236), .A2(G128), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n225), .A2(G119), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n331), .A2(new_n332), .ZN(new_n333));
  XNOR2_X1  g147(.A(KEYINPUT24), .B(G110), .ZN(new_n334));
  OR2_X1    g148(.A1(new_n333), .A2(new_n334), .ZN(new_n335));
  INV_X1    g149(.A(KEYINPUT23), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n332), .A2(new_n336), .ZN(new_n337));
  NAND3_X1  g151(.A1(new_n225), .A2(KEYINPUT23), .A3(G119), .ZN(new_n338));
  AND3_X1   g152(.A1(new_n337), .A2(new_n331), .A3(new_n338), .ZN(new_n339));
  INV_X1    g153(.A(G110), .ZN(new_n340));
  OR2_X1    g154(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  NAND4_X1  g155(.A1(new_n328), .A2(new_n330), .A3(new_n335), .A4(new_n341), .ZN(new_n342));
  NAND3_X1  g156(.A1(new_n319), .A2(new_n320), .A3(new_n199), .ZN(new_n343));
  AND2_X1   g157(.A1(new_n339), .A2(new_n340), .ZN(new_n344));
  AND2_X1   g158(.A1(new_n333), .A2(new_n334), .ZN(new_n345));
  OAI211_X1 g159(.A(new_n326), .B(new_n343), .C1(new_n344), .C2(new_n345), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n342), .A2(new_n346), .ZN(new_n347));
  NAND3_X1  g161(.A1(new_n255), .A2(G221), .A3(G234), .ZN(new_n348));
  XNOR2_X1  g162(.A(KEYINPUT22), .B(G137), .ZN(new_n349));
  XNOR2_X1  g163(.A(new_n348), .B(new_n349), .ZN(new_n350));
  INV_X1    g164(.A(new_n350), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n347), .A2(new_n351), .ZN(new_n352));
  NAND3_X1  g166(.A1(new_n342), .A2(new_n346), .A3(new_n350), .ZN(new_n353));
  INV_X1    g167(.A(KEYINPUT74), .ZN(new_n354));
  INV_X1    g168(.A(KEYINPUT25), .ZN(new_n355));
  AOI21_X1  g169(.A(G902), .B1(new_n354), .B2(new_n355), .ZN(new_n356));
  NAND3_X1  g170(.A1(new_n352), .A2(new_n353), .A3(new_n356), .ZN(new_n357));
  NOR2_X1   g171(.A1(new_n354), .A2(new_n355), .ZN(new_n358));
  AOI21_X1  g172(.A(new_n314), .B1(new_n357), .B2(new_n358), .ZN(new_n359));
  OAI21_X1  g173(.A(new_n359), .B1(new_n358), .B2(new_n357), .ZN(new_n360));
  AND2_X1   g174(.A1(new_n352), .A2(new_n353), .ZN(new_n361));
  AOI21_X1  g175(.A(G902), .B1(new_n313), .B2(G217), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n361), .A2(new_n362), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n360), .A2(new_n363), .ZN(new_n364));
  INV_X1    g178(.A(new_n364), .ZN(new_n365));
  NAND3_X1  g179(.A1(new_n307), .A2(new_n312), .A3(new_n365), .ZN(new_n366));
  INV_X1    g180(.A(KEYINPUT10), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n215), .A2(KEYINPUT77), .ZN(new_n368));
  INV_X1    g182(.A(KEYINPUT77), .ZN(new_n369));
  OAI211_X1 g183(.A(new_n369), .B(KEYINPUT1), .C1(new_n201), .C2(G146), .ZN(new_n370));
  NAND3_X1  g184(.A1(new_n368), .A2(G128), .A3(new_n370), .ZN(new_n371));
  AOI22_X1  g185(.A1(new_n371), .A2(new_n217), .B1(new_n214), .B2(new_n213), .ZN(new_n372));
  INV_X1    g186(.A(KEYINPUT3), .ZN(new_n373));
  INV_X1    g187(.A(G104), .ZN(new_n374));
  OAI21_X1  g188(.A(new_n373), .B1(new_n374), .B2(G107), .ZN(new_n375));
  INV_X1    g189(.A(G107), .ZN(new_n376));
  NAND3_X1  g190(.A1(new_n376), .A2(KEYINPUT3), .A3(G104), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n375), .A2(new_n377), .ZN(new_n378));
  INV_X1    g192(.A(G101), .ZN(new_n379));
  OAI21_X1  g193(.A(KEYINPUT76), .B1(new_n376), .B2(G104), .ZN(new_n380));
  INV_X1    g194(.A(KEYINPUT76), .ZN(new_n381));
  NAND3_X1  g195(.A1(new_n381), .A2(new_n374), .A3(G107), .ZN(new_n382));
  NAND4_X1  g196(.A1(new_n378), .A2(new_n379), .A3(new_n380), .A4(new_n382), .ZN(new_n383));
  NOR2_X1   g197(.A1(new_n374), .A2(G107), .ZN(new_n384));
  NOR2_X1   g198(.A1(new_n376), .A2(G104), .ZN(new_n385));
  OAI21_X1  g199(.A(G101), .B1(new_n384), .B2(new_n385), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n383), .A2(new_n386), .ZN(new_n387));
  OAI21_X1  g201(.A(new_n367), .B1(new_n372), .B2(new_n387), .ZN(new_n388));
  INV_X1    g202(.A(KEYINPUT78), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n388), .A2(new_n389), .ZN(new_n390));
  AND2_X1   g204(.A1(new_n383), .A2(new_n386), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n370), .A2(G128), .ZN(new_n392));
  AOI21_X1  g206(.A(new_n369), .B1(new_n200), .B2(KEYINPUT1), .ZN(new_n393));
  OAI21_X1  g207(.A(new_n217), .B1(new_n392), .B2(new_n393), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n394), .A2(new_n224), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n391), .A2(new_n395), .ZN(new_n396));
  NAND3_X1  g210(.A1(new_n396), .A2(KEYINPUT78), .A3(new_n367), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n390), .A2(new_n397), .ZN(new_n398));
  AND3_X1   g212(.A1(new_n376), .A2(KEYINPUT3), .A3(G104), .ZN(new_n399));
  AOI21_X1  g213(.A(KEYINPUT3), .B1(new_n376), .B2(G104), .ZN(new_n400));
  OAI211_X1 g214(.A(new_n380), .B(new_n382), .C1(new_n399), .C2(new_n400), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n401), .A2(G101), .ZN(new_n402));
  NAND3_X1  g216(.A1(new_n402), .A2(KEYINPUT4), .A3(new_n383), .ZN(new_n403));
  AOI21_X1  g217(.A(new_n210), .B1(new_n205), .B2(new_n207), .ZN(new_n404));
  INV_X1    g218(.A(KEYINPUT4), .ZN(new_n405));
  NAND3_X1  g219(.A1(new_n401), .A2(new_n405), .A3(G101), .ZN(new_n406));
  NAND3_X1  g220(.A1(new_n403), .A2(new_n404), .A3(new_n406), .ZN(new_n407));
  NAND3_X1  g221(.A1(new_n391), .A2(KEYINPUT10), .A3(new_n227), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n407), .A2(new_n408), .ZN(new_n409));
  INV_X1    g223(.A(new_n409), .ZN(new_n410));
  INV_X1    g224(.A(new_n198), .ZN(new_n411));
  NAND3_X1  g225(.A1(new_n398), .A2(new_n410), .A3(new_n411), .ZN(new_n412));
  INV_X1    g226(.A(KEYINPUT80), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n387), .A2(new_n218), .ZN(new_n414));
  INV_X1    g228(.A(KEYINPUT79), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n414), .A2(new_n415), .ZN(new_n416));
  AOI21_X1  g230(.A(new_n227), .B1(new_n383), .B2(new_n386), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n417), .A2(KEYINPUT79), .ZN(new_n418));
  NAND3_X1  g232(.A1(new_n416), .A2(new_n418), .A3(new_n396), .ZN(new_n419));
  AOI211_X1 g233(.A(new_n413), .B(KEYINPUT12), .C1(new_n419), .C2(new_n198), .ZN(new_n420));
  NOR2_X1   g234(.A1(new_n413), .A2(KEYINPUT12), .ZN(new_n421));
  OAI22_X1  g235(.A1(new_n417), .A2(KEYINPUT79), .B1(new_n372), .B2(new_n387), .ZN(new_n422));
  NOR2_X1   g236(.A1(new_n414), .A2(new_n415), .ZN(new_n423));
  OAI21_X1  g237(.A(new_n198), .B1(new_n422), .B2(new_n423), .ZN(new_n424));
  INV_X1    g238(.A(KEYINPUT12), .ZN(new_n425));
  NOR2_X1   g239(.A1(new_n425), .A2(KEYINPUT80), .ZN(new_n426));
  INV_X1    g240(.A(new_n426), .ZN(new_n427));
  AOI21_X1  g241(.A(new_n421), .B1(new_n424), .B2(new_n427), .ZN(new_n428));
  OAI21_X1  g242(.A(new_n412), .B1(new_n420), .B2(new_n428), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n255), .A2(G227), .ZN(new_n430));
  XOR2_X1   g244(.A(G110), .B(G140), .Z(new_n431));
  XNOR2_X1  g245(.A(new_n430), .B(new_n431), .ZN(new_n432));
  INV_X1    g246(.A(new_n432), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n429), .A2(new_n433), .ZN(new_n434));
  INV_X1    g248(.A(G469), .ZN(new_n435));
  INV_X1    g249(.A(G902), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n398), .A2(new_n410), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n437), .A2(new_n198), .ZN(new_n438));
  NAND3_X1  g252(.A1(new_n438), .A2(new_n432), .A3(new_n412), .ZN(new_n439));
  NAND4_X1  g253(.A1(new_n434), .A2(new_n435), .A3(new_n436), .A4(new_n439), .ZN(new_n440));
  NOR2_X1   g254(.A1(new_n435), .A2(new_n436), .ZN(new_n441));
  INV_X1    g255(.A(new_n441), .ZN(new_n442));
  NAND3_X1  g256(.A1(new_n438), .A2(new_n433), .A3(new_n412), .ZN(new_n443));
  INV_X1    g257(.A(new_n421), .ZN(new_n444));
  AOI22_X1  g258(.A1(new_n414), .A2(new_n415), .B1(new_n391), .B2(new_n395), .ZN(new_n445));
  AOI21_X1  g259(.A(new_n411), .B1(new_n445), .B2(new_n418), .ZN(new_n446));
  OAI21_X1  g260(.A(new_n444), .B1(new_n446), .B2(new_n426), .ZN(new_n447));
  NAND3_X1  g261(.A1(new_n424), .A2(KEYINPUT80), .A3(new_n425), .ZN(new_n448));
  AOI21_X1  g262(.A(new_n409), .B1(new_n390), .B2(new_n397), .ZN(new_n449));
  AOI22_X1  g263(.A1(new_n447), .A2(new_n448), .B1(new_n411), .B2(new_n449), .ZN(new_n450));
  OAI211_X1 g264(.A(G469), .B(new_n443), .C1(new_n450), .C2(new_n433), .ZN(new_n451));
  NAND3_X1  g265(.A1(new_n440), .A2(new_n442), .A3(new_n451), .ZN(new_n452));
  INV_X1    g266(.A(G221), .ZN(new_n453));
  XNOR2_X1  g267(.A(KEYINPUT9), .B(G234), .ZN(new_n454));
  INV_X1    g268(.A(KEYINPUT75), .ZN(new_n455));
  XNOR2_X1  g269(.A(new_n454), .B(new_n455), .ZN(new_n456));
  AOI21_X1  g270(.A(new_n453), .B1(new_n456), .B2(new_n436), .ZN(new_n457));
  INV_X1    g271(.A(new_n457), .ZN(new_n458));
  AND2_X1   g272(.A1(new_n452), .A2(new_n458), .ZN(new_n459));
  INV_X1    g273(.A(G217), .ZN(new_n460));
  NOR2_X1   g274(.A1(new_n460), .A2(G953), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n456), .A2(new_n461), .ZN(new_n462));
  INV_X1    g276(.A(KEYINPUT92), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  NAND3_X1  g278(.A1(new_n456), .A2(KEYINPUT92), .A3(new_n461), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  INV_X1    g280(.A(KEYINPUT90), .ZN(new_n467));
  INV_X1    g281(.A(G122), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n468), .A2(G116), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n234), .A2(G122), .ZN(new_n470));
  NAND3_X1  g284(.A1(new_n469), .A2(new_n470), .A3(new_n376), .ZN(new_n471));
  INV_X1    g285(.A(new_n471), .ZN(new_n472));
  AOI21_X1  g286(.A(new_n376), .B1(new_n469), .B2(new_n470), .ZN(new_n473));
  OAI21_X1  g287(.A(new_n467), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  INV_X1    g288(.A(new_n473), .ZN(new_n475));
  NAND3_X1  g289(.A1(new_n475), .A2(KEYINPUT90), .A3(new_n471), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n201), .A2(G128), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n225), .A2(G143), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  INV_X1    g293(.A(new_n479), .ZN(new_n480));
  INV_X1    g294(.A(KEYINPUT13), .ZN(new_n481));
  AOI21_X1  g295(.A(new_n189), .B1(new_n478), .B2(new_n481), .ZN(new_n482));
  OR2_X1    g296(.A1(new_n480), .A2(new_n482), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n480), .A2(new_n482), .ZN(new_n484));
  AOI22_X1  g298(.A1(new_n474), .A2(new_n476), .B1(new_n483), .B2(new_n484), .ZN(new_n485));
  INV_X1    g299(.A(new_n485), .ZN(new_n486));
  NAND3_X1  g300(.A1(new_n470), .A2(KEYINPUT91), .A3(KEYINPUT14), .ZN(new_n487));
  INV_X1    g301(.A(new_n487), .ZN(new_n488));
  AOI21_X1  g302(.A(KEYINPUT91), .B1(new_n470), .B2(KEYINPUT14), .ZN(new_n489));
  OAI221_X1 g303(.A(new_n469), .B1(KEYINPUT14), .B2(new_n470), .C1(new_n488), .C2(new_n489), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n490), .A2(G107), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n480), .A2(G134), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n479), .A2(new_n189), .ZN(new_n493));
  NAND3_X1  g307(.A1(new_n492), .A2(new_n471), .A3(new_n493), .ZN(new_n494));
  INV_X1    g308(.A(new_n494), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n491), .A2(new_n495), .ZN(new_n496));
  NAND3_X1  g310(.A1(new_n466), .A2(new_n486), .A3(new_n496), .ZN(new_n497));
  AOI21_X1  g311(.A(new_n494), .B1(new_n490), .B2(G107), .ZN(new_n498));
  OAI211_X1 g312(.A(new_n464), .B(new_n465), .C1(new_n498), .C2(new_n485), .ZN(new_n499));
  AOI21_X1  g313(.A(G902), .B1(new_n497), .B2(new_n499), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n500), .A2(KEYINPUT93), .ZN(new_n501));
  INV_X1    g315(.A(G478), .ZN(new_n502));
  NOR2_X1   g316(.A1(new_n502), .A2(KEYINPUT15), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n501), .A2(new_n503), .ZN(new_n504));
  INV_X1    g318(.A(new_n503), .ZN(new_n505));
  NAND3_X1  g319(.A1(new_n500), .A2(KEYINPUT93), .A3(new_n505), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n504), .A2(new_n506), .ZN(new_n507));
  INV_X1    g321(.A(new_n507), .ZN(new_n508));
  INV_X1    g322(.A(G475), .ZN(new_n509));
  OAI21_X1  g323(.A(new_n317), .B1(new_n321), .B2(new_n315), .ZN(new_n510));
  OAI21_X1  g324(.A(new_n343), .B1(new_n510), .B2(new_n199), .ZN(new_n511));
  NAND4_X1  g325(.A1(new_n248), .A2(G214), .A3(new_n249), .A4(new_n250), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n512), .A2(new_n201), .ZN(new_n513));
  NAND4_X1  g327(.A1(new_n255), .A2(G143), .A3(G214), .A4(new_n249), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  AND2_X1   g329(.A1(KEYINPUT18), .A2(G131), .ZN(new_n516));
  OAI21_X1  g330(.A(new_n511), .B1(new_n515), .B2(new_n516), .ZN(new_n517));
  AND2_X1   g331(.A1(new_n515), .A2(new_n516), .ZN(new_n518));
  NOR2_X1   g332(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n515), .A2(G131), .ZN(new_n520));
  INV_X1    g334(.A(KEYINPUT85), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  NAND3_X1  g336(.A1(new_n515), .A2(KEYINPUT85), .A3(G131), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  AOI22_X1  g338(.A1(new_n524), .A2(KEYINPUT17), .B1(new_n330), .B2(new_n328), .ZN(new_n525));
  AOI21_X1  g339(.A(KEYINPUT85), .B1(new_n515), .B2(G131), .ZN(new_n526));
  AOI211_X1 g340(.A(new_n521), .B(new_n196), .C1(new_n513), .C2(new_n514), .ZN(new_n527));
  NOR2_X1   g341(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  INV_X1    g342(.A(KEYINPUT17), .ZN(new_n529));
  INV_X1    g343(.A(KEYINPUT84), .ZN(new_n530));
  OAI21_X1  g344(.A(new_n530), .B1(new_n515), .B2(G131), .ZN(new_n531));
  NAND4_X1  g345(.A1(new_n513), .A2(new_n514), .A3(KEYINPUT84), .A4(new_n196), .ZN(new_n532));
  NAND4_X1  g346(.A1(new_n528), .A2(new_n529), .A3(new_n531), .A4(new_n532), .ZN(new_n533));
  AOI21_X1  g347(.A(new_n519), .B1(new_n525), .B2(new_n533), .ZN(new_n534));
  XNOR2_X1  g348(.A(G113), .B(G122), .ZN(new_n535));
  XNOR2_X1  g349(.A(new_n535), .B(G104), .ZN(new_n536));
  INV_X1    g350(.A(new_n536), .ZN(new_n537));
  NOR2_X1   g351(.A1(new_n537), .A2(KEYINPUT89), .ZN(new_n538));
  NOR2_X1   g352(.A1(new_n534), .A2(new_n538), .ZN(new_n539));
  INV_X1    g353(.A(new_n539), .ZN(new_n540));
  AOI21_X1  g354(.A(G902), .B1(new_n534), .B2(new_n538), .ZN(new_n541));
  AOI21_X1  g355(.A(new_n509), .B1(new_n540), .B2(new_n541), .ZN(new_n542));
  INV_X1    g356(.A(KEYINPUT87), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n328), .A2(new_n330), .ZN(new_n544));
  OAI21_X1  g358(.A(KEYINPUT17), .B1(new_n526), .B2(new_n527), .ZN(new_n545));
  NAND4_X1  g359(.A1(new_n522), .A2(new_n523), .A3(new_n531), .A4(new_n532), .ZN(new_n546));
  OAI211_X1 g360(.A(new_n544), .B(new_n545), .C1(new_n546), .C2(KEYINPUT17), .ZN(new_n547));
  INV_X1    g361(.A(new_n519), .ZN(new_n548));
  AOI21_X1  g362(.A(new_n536), .B1(new_n547), .B2(new_n548), .ZN(new_n549));
  OAI21_X1  g363(.A(new_n536), .B1(new_n517), .B2(new_n518), .ZN(new_n550));
  INV_X1    g364(.A(new_n326), .ZN(new_n551));
  NOR3_X1   g365(.A1(new_n321), .A2(KEYINPUT86), .A3(KEYINPUT19), .ZN(new_n552));
  INV_X1    g366(.A(KEYINPUT86), .ZN(new_n553));
  OAI21_X1  g367(.A(new_n510), .B1(new_n553), .B2(new_n321), .ZN(new_n554));
  AOI21_X1  g368(.A(new_n552), .B1(new_n554), .B2(KEYINPUT19), .ZN(new_n555));
  AOI21_X1  g369(.A(new_n551), .B1(new_n555), .B2(new_n199), .ZN(new_n556));
  AOI21_X1  g370(.A(new_n550), .B1(new_n556), .B2(new_n546), .ZN(new_n557));
  OAI21_X1  g371(.A(new_n543), .B1(new_n549), .B2(new_n557), .ZN(new_n558));
  NOR2_X1   g372(.A1(G475), .A2(G902), .ZN(new_n559));
  INV_X1    g373(.A(new_n557), .ZN(new_n560));
  OAI211_X1 g374(.A(KEYINPUT87), .B(new_n560), .C1(new_n534), .C2(new_n536), .ZN(new_n561));
  NAND3_X1  g375(.A1(new_n558), .A2(new_n559), .A3(new_n561), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n562), .A2(KEYINPUT20), .ZN(new_n563));
  INV_X1    g377(.A(KEYINPUT88), .ZN(new_n564));
  NOR2_X1   g378(.A1(new_n546), .A2(KEYINPUT17), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n544), .A2(new_n545), .ZN(new_n566));
  OAI21_X1  g380(.A(new_n548), .B1(new_n565), .B2(new_n566), .ZN(new_n567));
  AOI21_X1  g381(.A(new_n557), .B1(new_n567), .B2(new_n537), .ZN(new_n568));
  NOR3_X1   g382(.A1(KEYINPUT20), .A2(G475), .A3(G902), .ZN(new_n569));
  AOI21_X1  g383(.A(new_n564), .B1(new_n568), .B2(new_n569), .ZN(new_n570));
  INV_X1    g384(.A(new_n569), .ZN(new_n571));
  NOR4_X1   g385(.A1(new_n549), .A2(KEYINPUT88), .A3(new_n557), .A4(new_n571), .ZN(new_n572));
  NOR2_X1   g386(.A1(new_n570), .A2(new_n572), .ZN(new_n573));
  AOI21_X1  g387(.A(new_n542), .B1(new_n563), .B2(new_n573), .ZN(new_n574));
  NAND3_X1  g388(.A1(new_n403), .A2(new_n241), .A3(new_n406), .ZN(new_n575));
  OR2_X1    g389(.A1(new_n239), .A2(new_n240), .ZN(new_n576));
  INV_X1    g390(.A(KEYINPUT5), .ZN(new_n577));
  NAND3_X1  g391(.A1(new_n577), .A2(new_n236), .A3(G116), .ZN(new_n578));
  OAI211_X1 g392(.A(G113), .B(new_n578), .C1(new_n239), .C2(new_n577), .ZN(new_n579));
  NAND3_X1  g393(.A1(new_n391), .A2(new_n576), .A3(new_n579), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n575), .A2(new_n580), .ZN(new_n581));
  XNOR2_X1  g395(.A(G110), .B(G122), .ZN(new_n582));
  INV_X1    g396(.A(new_n582), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n581), .A2(new_n583), .ZN(new_n584));
  NAND3_X1  g398(.A1(new_n575), .A2(new_n582), .A3(new_n580), .ZN(new_n585));
  NAND3_X1  g399(.A1(new_n584), .A2(KEYINPUT6), .A3(new_n585), .ZN(new_n586));
  INV_X1    g400(.A(KEYINPUT6), .ZN(new_n587));
  NAND3_X1  g401(.A1(new_n581), .A2(new_n587), .A3(new_n583), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n218), .A2(new_n316), .ZN(new_n589));
  OAI21_X1  g403(.A(new_n589), .B1(new_n404), .B2(new_n316), .ZN(new_n590));
  INV_X1    g404(.A(G224), .ZN(new_n591));
  NOR2_X1   g405(.A1(new_n591), .A2(G953), .ZN(new_n592));
  XNOR2_X1  g406(.A(new_n590), .B(new_n592), .ZN(new_n593));
  NAND3_X1  g407(.A1(new_n586), .A2(new_n588), .A3(new_n593), .ZN(new_n594));
  XNOR2_X1  g408(.A(new_n582), .B(KEYINPUT8), .ZN(new_n595));
  AND4_X1   g409(.A1(new_n576), .A2(new_n579), .A3(new_n383), .A4(new_n386), .ZN(new_n596));
  AOI22_X1  g410(.A1(new_n579), .A2(new_n576), .B1(new_n383), .B2(new_n386), .ZN(new_n597));
  OAI21_X1  g411(.A(new_n595), .B1(new_n596), .B2(new_n597), .ZN(new_n598));
  AND2_X1   g412(.A1(new_n585), .A2(new_n598), .ZN(new_n599));
  NAND2_X1  g413(.A1(KEYINPUT81), .A2(KEYINPUT7), .ZN(new_n600));
  OAI211_X1 g414(.A(new_n589), .B(new_n600), .C1(new_n404), .C2(new_n316), .ZN(new_n601));
  INV_X1    g415(.A(KEYINPUT7), .ZN(new_n602));
  NOR2_X1   g416(.A1(new_n592), .A2(new_n602), .ZN(new_n603));
  XNOR2_X1  g417(.A(new_n601), .B(new_n603), .ZN(new_n604));
  AOI21_X1  g418(.A(G902), .B1(new_n599), .B2(new_n604), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n594), .A2(new_n605), .ZN(new_n606));
  OAI21_X1  g420(.A(G210), .B1(G237), .B2(G902), .ZN(new_n607));
  XOR2_X1   g421(.A(new_n607), .B(KEYINPUT83), .Z(new_n608));
  NAND2_X1  g422(.A1(new_n608), .A2(KEYINPUT82), .ZN(new_n609));
  XNOR2_X1  g423(.A(new_n606), .B(new_n609), .ZN(new_n610));
  OAI21_X1  g424(.A(G214), .B1(G237), .B2(G902), .ZN(new_n611));
  INV_X1    g425(.A(new_n611), .ZN(new_n612));
  INV_X1    g426(.A(G952), .ZN(new_n613));
  NOR2_X1   g427(.A1(new_n613), .A2(G953), .ZN(new_n614));
  NAND2_X1  g428(.A1(G234), .A2(G237), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  INV_X1    g430(.A(new_n616), .ZN(new_n617));
  INV_X1    g431(.A(new_n255), .ZN(new_n618));
  NAND3_X1  g432(.A1(new_n618), .A2(G902), .A3(new_n615), .ZN(new_n619));
  INV_X1    g433(.A(new_n619), .ZN(new_n620));
  XNOR2_X1  g434(.A(KEYINPUT21), .B(G898), .ZN(new_n621));
  AOI21_X1  g435(.A(new_n617), .B1(new_n620), .B2(new_n621), .ZN(new_n622));
  NOR3_X1   g436(.A1(new_n610), .A2(new_n612), .A3(new_n622), .ZN(new_n623));
  NAND4_X1  g437(.A1(new_n459), .A2(new_n508), .A3(new_n574), .A4(new_n623), .ZN(new_n624));
  OR2_X1    g438(.A1(new_n366), .A2(new_n624), .ZN(new_n625));
  XOR2_X1   g439(.A(KEYINPUT94), .B(G101), .Z(new_n626));
  XNOR2_X1  g440(.A(new_n626), .B(KEYINPUT95), .ZN(new_n627));
  XNOR2_X1  g441(.A(new_n625), .B(new_n627), .ZN(G3));
  NAND2_X1  g442(.A1(new_n304), .A2(new_n436), .ZN(new_n629));
  AOI22_X1  g443(.A1(new_n629), .A2(G472), .B1(new_n297), .B2(new_n304), .ZN(new_n630));
  NAND3_X1  g444(.A1(new_n459), .A2(new_n630), .A3(new_n365), .ZN(new_n631));
  INV_X1    g445(.A(new_n631), .ZN(new_n632));
  INV_X1    g446(.A(KEYINPUT33), .ZN(new_n633));
  AOI21_X1  g447(.A(new_n633), .B1(new_n497), .B2(KEYINPUT96), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n497), .A2(new_n499), .ZN(new_n635));
  XNOR2_X1  g449(.A(new_n634), .B(new_n635), .ZN(new_n636));
  NAND3_X1  g450(.A1(new_n636), .A2(G478), .A3(new_n436), .ZN(new_n637));
  XNOR2_X1  g451(.A(KEYINPUT97), .B(G478), .ZN(new_n638));
  OR2_X1    g452(.A1(new_n500), .A2(new_n638), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n637), .A2(new_n639), .ZN(new_n640));
  INV_X1    g454(.A(new_n640), .ZN(new_n641));
  NAND3_X1  g455(.A1(new_n594), .A2(new_n605), .A3(new_n608), .ZN(new_n642));
  INV_X1    g456(.A(new_n642), .ZN(new_n643));
  AOI21_X1  g457(.A(new_n608), .B1(new_n594), .B2(new_n605), .ZN(new_n644));
  NOR3_X1   g458(.A1(new_n643), .A2(new_n644), .A3(new_n612), .ZN(new_n645));
  INV_X1    g459(.A(new_n622), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  NOR3_X1   g461(.A1(new_n574), .A2(new_n641), .A3(new_n647), .ZN(new_n648));
  NAND2_X1  g462(.A1(new_n632), .A2(new_n648), .ZN(new_n649));
  XOR2_X1   g463(.A(KEYINPUT34), .B(G104), .Z(new_n650));
  XNOR2_X1  g464(.A(new_n649), .B(new_n650), .ZN(G6));
  INV_X1    g465(.A(new_n538), .ZN(new_n652));
  OAI21_X1  g466(.A(new_n436), .B1(new_n567), .B2(new_n652), .ZN(new_n653));
  OAI21_X1  g467(.A(G475), .B1(new_n653), .B2(new_n539), .ZN(new_n654));
  NAND2_X1  g468(.A1(new_n654), .A2(new_n507), .ZN(new_n655));
  NAND3_X1  g469(.A1(new_n558), .A2(new_n561), .A3(new_n569), .ZN(new_n656));
  AOI21_X1  g470(.A(new_n655), .B1(new_n563), .B2(new_n656), .ZN(new_n657));
  NOR4_X1   g471(.A1(new_n643), .A2(new_n644), .A3(new_n612), .A4(new_n622), .ZN(new_n658));
  AOI21_X1  g472(.A(KEYINPUT98), .B1(new_n657), .B2(new_n658), .ZN(new_n659));
  INV_X1    g473(.A(new_n659), .ZN(new_n660));
  NAND3_X1  g474(.A1(new_n657), .A2(KEYINPUT98), .A3(new_n658), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  NAND2_X1  g476(.A1(new_n662), .A2(new_n632), .ZN(new_n663));
  XOR2_X1   g477(.A(KEYINPUT35), .B(G107), .Z(new_n664));
  XNOR2_X1  g478(.A(new_n663), .B(new_n664), .ZN(G9));
  NAND2_X1  g479(.A1(new_n459), .A2(new_n630), .ZN(new_n666));
  NOR2_X1   g480(.A1(new_n351), .A2(KEYINPUT36), .ZN(new_n667));
  XNOR2_X1  g481(.A(new_n347), .B(new_n667), .ZN(new_n668));
  NAND2_X1  g482(.A1(new_n668), .A2(new_n362), .ZN(new_n669));
  NAND2_X1  g483(.A1(new_n360), .A2(new_n669), .ZN(new_n670));
  NAND4_X1  g484(.A1(new_n623), .A2(new_n574), .A3(new_n508), .A4(new_n670), .ZN(new_n671));
  OR2_X1    g485(.A1(new_n666), .A2(new_n671), .ZN(new_n672));
  XOR2_X1   g486(.A(KEYINPUT37), .B(G110), .Z(new_n673));
  XNOR2_X1  g487(.A(new_n672), .B(new_n673), .ZN(G12));
  AND4_X1   g488(.A1(new_n307), .A2(new_n312), .A3(new_n459), .A4(new_n670), .ZN(new_n675));
  NAND2_X1  g489(.A1(new_n563), .A2(new_n656), .ZN(new_n676));
  INV_X1    g490(.A(new_n655), .ZN(new_n677));
  XNOR2_X1  g491(.A(new_n616), .B(KEYINPUT99), .ZN(new_n678));
  INV_X1    g492(.A(new_n678), .ZN(new_n679));
  INV_X1    g493(.A(G900), .ZN(new_n680));
  AOI21_X1  g494(.A(new_n679), .B1(new_n620), .B2(new_n680), .ZN(new_n681));
  INV_X1    g495(.A(new_n681), .ZN(new_n682));
  NAND4_X1  g496(.A1(new_n676), .A2(new_n645), .A3(new_n677), .A4(new_n682), .ZN(new_n683));
  INV_X1    g497(.A(KEYINPUT100), .ZN(new_n684));
  NAND2_X1  g498(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  NAND4_X1  g499(.A1(new_n657), .A2(KEYINPUT100), .A3(new_n645), .A4(new_n682), .ZN(new_n686));
  NAND2_X1  g500(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  NAND2_X1  g501(.A1(new_n675), .A2(new_n687), .ZN(new_n688));
  XNOR2_X1  g502(.A(new_n688), .B(G128), .ZN(G30));
  NAND2_X1  g503(.A1(new_n563), .A2(new_n573), .ZN(new_n690));
  NAND2_X1  g504(.A1(new_n690), .A2(new_n654), .ZN(new_n691));
  XOR2_X1   g505(.A(new_n610), .B(KEYINPUT38), .Z(new_n692));
  NOR2_X1   g506(.A1(new_n670), .A2(new_n508), .ZN(new_n693));
  AND4_X1   g507(.A1(new_n691), .A2(new_n692), .A3(new_n611), .A4(new_n693), .ZN(new_n694));
  NAND2_X1  g508(.A1(new_n294), .A2(new_n244), .ZN(new_n695));
  INV_X1    g509(.A(new_n246), .ZN(new_n696));
  OAI21_X1  g510(.A(new_n268), .B1(new_n696), .B2(new_n277), .ZN(new_n697));
  AND2_X1   g511(.A1(new_n695), .A2(new_n697), .ZN(new_n698));
  OAI21_X1  g512(.A(G472), .B1(new_n698), .B2(G902), .ZN(new_n699));
  NAND2_X1  g513(.A1(new_n310), .A2(new_n699), .ZN(new_n700));
  XNOR2_X1  g514(.A(new_n700), .B(KEYINPUT101), .ZN(new_n701));
  INV_X1    g515(.A(new_n701), .ZN(new_n702));
  XOR2_X1   g516(.A(new_n681), .B(KEYINPUT39), .Z(new_n703));
  NAND2_X1  g517(.A1(new_n459), .A2(new_n703), .ZN(new_n704));
  OR2_X1    g518(.A1(new_n704), .A2(KEYINPUT40), .ZN(new_n705));
  NAND2_X1  g519(.A1(new_n704), .A2(KEYINPUT40), .ZN(new_n706));
  NAND4_X1  g520(.A1(new_n694), .A2(new_n702), .A3(new_n705), .A4(new_n706), .ZN(new_n707));
  XNOR2_X1  g521(.A(new_n707), .B(G143), .ZN(G45));
  AOI21_X1  g522(.A(new_n311), .B1(new_n310), .B2(new_n282), .ZN(new_n709));
  AOI211_X1 g523(.A(KEYINPUT71), .B(new_n281), .C1(new_n308), .C2(new_n309), .ZN(new_n710));
  INV_X1    g524(.A(new_n670), .ZN(new_n711));
  NOR3_X1   g525(.A1(new_n709), .A2(new_n710), .A3(new_n711), .ZN(new_n712));
  INV_X1    g526(.A(new_n645), .ZN(new_n713));
  NOR4_X1   g527(.A1(new_n574), .A2(new_n713), .A3(new_n641), .A4(new_n681), .ZN(new_n714));
  NAND3_X1  g528(.A1(new_n712), .A2(new_n459), .A3(new_n714), .ZN(new_n715));
  XNOR2_X1  g529(.A(new_n715), .B(G146), .ZN(G48));
  NOR2_X1   g530(.A1(new_n709), .A2(new_n710), .ZN(new_n717));
  OAI211_X1 g531(.A(new_n436), .B(new_n439), .C1(new_n450), .C2(new_n432), .ZN(new_n718));
  NAND2_X1  g532(.A1(new_n718), .A2(G469), .ZN(new_n719));
  NAND3_X1  g533(.A1(new_n719), .A2(new_n458), .A3(new_n440), .ZN(new_n720));
  NAND2_X1  g534(.A1(new_n720), .A2(KEYINPUT102), .ZN(new_n721));
  INV_X1    g535(.A(KEYINPUT102), .ZN(new_n722));
  NAND4_X1  g536(.A1(new_n719), .A2(new_n440), .A3(new_n722), .A4(new_n458), .ZN(new_n723));
  AND2_X1   g537(.A1(new_n721), .A2(new_n723), .ZN(new_n724));
  NAND4_X1  g538(.A1(new_n717), .A2(new_n724), .A3(new_n365), .A4(new_n648), .ZN(new_n725));
  XNOR2_X1  g539(.A(KEYINPUT41), .B(G113), .ZN(new_n726));
  XNOR2_X1  g540(.A(new_n725), .B(new_n726), .ZN(G15));
  NOR3_X1   g541(.A1(new_n709), .A2(new_n710), .A3(new_n364), .ZN(new_n728));
  NAND3_X1  g542(.A1(new_n662), .A2(new_n728), .A3(new_n724), .ZN(new_n729));
  XNOR2_X1  g543(.A(new_n729), .B(G116), .ZN(G18));
  NAND3_X1  g544(.A1(new_n690), .A2(new_n508), .A3(new_n654), .ZN(new_n731));
  NAND4_X1  g545(.A1(new_n658), .A2(new_n458), .A3(new_n440), .A4(new_n719), .ZN(new_n732));
  NOR2_X1   g546(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  NAND3_X1  g547(.A1(new_n717), .A2(new_n733), .A3(new_n670), .ZN(new_n734));
  XNOR2_X1  g548(.A(new_n734), .B(G119), .ZN(G21));
  AND3_X1   g549(.A1(new_n721), .A2(new_n646), .A3(new_n723), .ZN(new_n736));
  NOR3_X1   g550(.A1(new_n574), .A2(new_n508), .A3(new_n713), .ZN(new_n737));
  NAND2_X1  g551(.A1(new_n291), .A2(new_n295), .ZN(new_n738));
  OAI21_X1  g552(.A(new_n268), .B1(new_n276), .B2(new_n277), .ZN(new_n739));
  AOI21_X1  g553(.A(new_n298), .B1(new_n738), .B2(new_n739), .ZN(new_n740));
  OAI21_X1  g554(.A(G472), .B1(new_n296), .B2(G902), .ZN(new_n741));
  NAND2_X1  g555(.A1(new_n741), .A2(KEYINPUT103), .ZN(new_n742));
  INV_X1    g556(.A(KEYINPUT103), .ZN(new_n743));
  NAND3_X1  g557(.A1(new_n629), .A2(new_n743), .A3(G472), .ZN(new_n744));
  AOI211_X1 g558(.A(new_n740), .B(new_n364), .C1(new_n742), .C2(new_n744), .ZN(new_n745));
  NAND3_X1  g559(.A1(new_n736), .A2(new_n737), .A3(new_n745), .ZN(new_n746));
  XNOR2_X1  g560(.A(new_n746), .B(G122), .ZN(G24));
  NAND3_X1  g561(.A1(new_n568), .A2(new_n564), .A3(new_n569), .ZN(new_n748));
  OAI211_X1 g562(.A(new_n560), .B(new_n569), .C1(new_n534), .C2(new_n536), .ZN(new_n749));
  NAND2_X1  g563(.A1(new_n749), .A2(KEYINPUT88), .ZN(new_n750));
  NAND2_X1  g564(.A1(new_n748), .A2(new_n750), .ZN(new_n751));
  AOI21_X1  g565(.A(new_n751), .B1(KEYINPUT20), .B2(new_n562), .ZN(new_n752));
  OAI211_X1 g566(.A(new_n640), .B(new_n682), .C1(new_n752), .C2(new_n542), .ZN(new_n753));
  INV_X1    g567(.A(new_n740), .ZN(new_n754));
  AOI21_X1  g568(.A(new_n743), .B1(new_n629), .B2(G472), .ZN(new_n755));
  AOI211_X1 g569(.A(KEYINPUT103), .B(new_n187), .C1(new_n304), .C2(new_n436), .ZN(new_n756));
  OAI211_X1 g570(.A(new_n670), .B(new_n754), .C1(new_n755), .C2(new_n756), .ZN(new_n757));
  NOR2_X1   g571(.A1(new_n753), .A2(new_n757), .ZN(new_n758));
  NOR2_X1   g572(.A1(new_n720), .A2(new_n713), .ZN(new_n759));
  NAND2_X1  g573(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  XNOR2_X1  g574(.A(new_n760), .B(G125), .ZN(G27));
  NOR2_X1   g575(.A1(new_n753), .A2(KEYINPUT42), .ZN(new_n762));
  OAI21_X1  g576(.A(KEYINPUT104), .B1(new_n450), .B2(new_n433), .ZN(new_n763));
  INV_X1    g577(.A(KEYINPUT104), .ZN(new_n764));
  NAND3_X1  g578(.A1(new_n429), .A2(new_n764), .A3(new_n432), .ZN(new_n765));
  NAND4_X1  g579(.A1(new_n763), .A2(new_n765), .A3(G469), .A4(new_n443), .ZN(new_n766));
  NAND2_X1  g580(.A1(new_n766), .A2(KEYINPUT105), .ZN(new_n767));
  AND3_X1   g581(.A1(new_n438), .A2(new_n433), .A3(new_n412), .ZN(new_n768));
  NAND2_X1  g582(.A1(new_n447), .A2(new_n448), .ZN(new_n769));
  AOI21_X1  g583(.A(new_n433), .B1(new_n769), .B2(new_n412), .ZN(new_n770));
  AOI21_X1  g584(.A(new_n768), .B1(new_n770), .B2(new_n764), .ZN(new_n771));
  INV_X1    g585(.A(KEYINPUT105), .ZN(new_n772));
  NAND4_X1  g586(.A1(new_n771), .A2(new_n772), .A3(G469), .A4(new_n763), .ZN(new_n773));
  NAND4_X1  g587(.A1(new_n767), .A2(new_n773), .A3(new_n440), .A4(new_n442), .ZN(new_n774));
  AND3_X1   g588(.A1(new_n610), .A2(new_n458), .A3(new_n611), .ZN(new_n775));
  AND3_X1   g589(.A1(new_n774), .A2(KEYINPUT106), .A3(new_n775), .ZN(new_n776));
  AOI21_X1  g590(.A(KEYINPUT106), .B1(new_n774), .B2(new_n775), .ZN(new_n777));
  OAI211_X1 g591(.A(new_n728), .B(new_n762), .C1(new_n776), .C2(new_n777), .ZN(new_n778));
  AOI21_X1  g592(.A(new_n641), .B1(new_n690), .B2(new_n654), .ZN(new_n779));
  NAND4_X1  g593(.A1(new_n779), .A2(new_n306), .A3(new_n365), .A4(new_n682), .ZN(new_n780));
  OAI211_X1 g594(.A(new_n440), .B(new_n442), .C1(new_n766), .C2(KEYINPUT105), .ZN(new_n781));
  AND2_X1   g595(.A1(new_n766), .A2(KEYINPUT105), .ZN(new_n782));
  OAI21_X1  g596(.A(new_n775), .B1(new_n781), .B2(new_n782), .ZN(new_n783));
  INV_X1    g597(.A(KEYINPUT106), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  NAND3_X1  g599(.A1(new_n774), .A2(KEYINPUT106), .A3(new_n775), .ZN(new_n786));
  AOI21_X1  g600(.A(new_n780), .B1(new_n785), .B2(new_n786), .ZN(new_n787));
  INV_X1    g601(.A(KEYINPUT42), .ZN(new_n788));
  OAI21_X1  g602(.A(new_n778), .B1(new_n787), .B2(new_n788), .ZN(new_n789));
  XNOR2_X1  g603(.A(new_n789), .B(new_n196), .ZN(G33));
  INV_X1    g604(.A(KEYINPUT107), .ZN(new_n791));
  AND3_X1   g605(.A1(new_n657), .A2(new_n791), .A3(new_n682), .ZN(new_n792));
  AOI21_X1  g606(.A(new_n791), .B1(new_n657), .B2(new_n682), .ZN(new_n793));
  NOR2_X1   g607(.A1(new_n792), .A2(new_n793), .ZN(new_n794));
  OAI211_X1 g608(.A(new_n794), .B(new_n728), .C1(new_n776), .C2(new_n777), .ZN(new_n795));
  XNOR2_X1  g609(.A(KEYINPUT108), .B(G134), .ZN(new_n796));
  XNOR2_X1  g610(.A(new_n795), .B(new_n796), .ZN(G36));
  INV_X1    g611(.A(KEYINPUT109), .ZN(new_n798));
  OAI21_X1  g612(.A(new_n798), .B1(new_n691), .B2(new_n641), .ZN(new_n799));
  INV_X1    g613(.A(KEYINPUT43), .ZN(new_n800));
  NAND2_X1  g614(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  OAI211_X1 g615(.A(new_n798), .B(KEYINPUT43), .C1(new_n691), .C2(new_n641), .ZN(new_n802));
  AND2_X1   g616(.A1(new_n801), .A2(new_n802), .ZN(new_n803));
  NOR2_X1   g617(.A1(new_n711), .A2(new_n630), .ZN(new_n804));
  XOR2_X1   g618(.A(new_n804), .B(KEYINPUT110), .Z(new_n805));
  AOI21_X1  g619(.A(KEYINPUT44), .B1(new_n803), .B2(new_n805), .ZN(new_n806));
  XNOR2_X1  g620(.A(new_n806), .B(KEYINPUT111), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n610), .A2(new_n611), .ZN(new_n808));
  NAND3_X1  g622(.A1(new_n771), .A2(KEYINPUT45), .A3(new_n763), .ZN(new_n809));
  OAI21_X1  g623(.A(new_n443), .B1(new_n450), .B2(new_n433), .ZN(new_n810));
  INV_X1    g624(.A(KEYINPUT45), .ZN(new_n811));
  AOI21_X1  g625(.A(new_n435), .B1(new_n810), .B2(new_n811), .ZN(new_n812));
  AOI21_X1  g626(.A(new_n441), .B1(new_n809), .B2(new_n812), .ZN(new_n813));
  AND2_X1   g627(.A1(new_n813), .A2(KEYINPUT46), .ZN(new_n814));
  OAI21_X1  g628(.A(new_n440), .B1(new_n813), .B2(KEYINPUT46), .ZN(new_n815));
  OAI211_X1 g629(.A(new_n458), .B(new_n703), .C1(new_n814), .C2(new_n815), .ZN(new_n816));
  AND2_X1   g630(.A1(new_n803), .A2(new_n805), .ZN(new_n817));
  AOI211_X1 g631(.A(new_n808), .B(new_n816), .C1(new_n817), .C2(KEYINPUT44), .ZN(new_n818));
  NAND2_X1  g632(.A1(new_n807), .A2(new_n818), .ZN(new_n819));
  XNOR2_X1  g633(.A(new_n819), .B(G137), .ZN(G39));
  NOR3_X1   g634(.A1(new_n717), .A2(new_n365), .A3(new_n808), .ZN(new_n821));
  NAND3_X1  g635(.A1(new_n821), .A2(new_n779), .A3(new_n682), .ZN(new_n822));
  OAI21_X1  g636(.A(new_n458), .B1(new_n814), .B2(new_n815), .ZN(new_n823));
  INV_X1    g637(.A(KEYINPUT47), .ZN(new_n824));
  NAND2_X1  g638(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  OAI211_X1 g639(.A(KEYINPUT47), .B(new_n458), .C1(new_n814), .C2(new_n815), .ZN(new_n826));
  AOI21_X1  g640(.A(new_n822), .B1(new_n825), .B2(new_n826), .ZN(new_n827));
  XNOR2_X1  g641(.A(new_n827), .B(new_n318), .ZN(G42));
  INV_X1    g642(.A(KEYINPUT120), .ZN(new_n829));
  NOR2_X1   g643(.A1(new_n720), .A2(new_n808), .ZN(new_n830));
  NAND4_X1  g644(.A1(new_n701), .A2(new_n365), .A3(new_n617), .A4(new_n830), .ZN(new_n831));
  NOR3_X1   g645(.A1(new_n831), .A2(new_n691), .A3(new_n640), .ZN(new_n832));
  NAND3_X1  g646(.A1(new_n803), .A2(new_n679), .A3(new_n830), .ZN(new_n833));
  INV_X1    g647(.A(new_n833), .ZN(new_n834));
  INV_X1    g648(.A(new_n757), .ZN(new_n835));
  AOI21_X1  g649(.A(new_n832), .B1(new_n834), .B2(new_n835), .ZN(new_n836));
  NAND2_X1  g650(.A1(new_n719), .A2(new_n440), .ZN(new_n837));
  OAI211_X1 g651(.A(new_n825), .B(new_n826), .C1(new_n458), .C2(new_n837), .ZN(new_n838));
  INV_X1    g652(.A(new_n808), .ZN(new_n839));
  NAND4_X1  g653(.A1(new_n801), .A2(new_n679), .A3(new_n745), .A4(new_n802), .ZN(new_n840));
  INV_X1    g654(.A(new_n840), .ZN(new_n841));
  NAND3_X1  g655(.A1(new_n838), .A2(new_n839), .A3(new_n841), .ZN(new_n842));
  NAND2_X1  g656(.A1(new_n836), .A2(new_n842), .ZN(new_n843));
  INV_X1    g657(.A(KEYINPUT119), .ZN(new_n844));
  INV_X1    g658(.A(KEYINPUT50), .ZN(new_n845));
  INV_X1    g659(.A(KEYINPUT117), .ZN(new_n846));
  OR3_X1    g660(.A1(new_n692), .A2(new_n611), .A3(new_n720), .ZN(new_n847));
  NOR3_X1   g661(.A1(new_n840), .A2(new_n846), .A3(new_n847), .ZN(new_n848));
  OAI21_X1  g662(.A(new_n845), .B1(new_n848), .B2(KEYINPUT118), .ZN(new_n849));
  OAI21_X1  g663(.A(KEYINPUT117), .B1(new_n845), .B2(KEYINPUT118), .ZN(new_n850));
  OAI21_X1  g664(.A(new_n850), .B1(new_n840), .B2(new_n847), .ZN(new_n851));
  NAND2_X1  g665(.A1(new_n849), .A2(new_n851), .ZN(new_n852));
  AOI21_X1  g666(.A(new_n843), .B1(new_n844), .B2(new_n852), .ZN(new_n853));
  NAND3_X1  g667(.A1(new_n849), .A2(KEYINPUT119), .A3(new_n851), .ZN(new_n854));
  AOI21_X1  g668(.A(KEYINPUT51), .B1(new_n853), .B2(new_n854), .ZN(new_n855));
  NAND2_X1  g669(.A1(new_n306), .A2(new_n365), .ZN(new_n856));
  NOR2_X1   g670(.A1(new_n833), .A2(new_n856), .ZN(new_n857));
  INV_X1    g671(.A(KEYINPUT48), .ZN(new_n858));
  XNOR2_X1  g672(.A(new_n857), .B(new_n858), .ZN(new_n859));
  INV_X1    g673(.A(new_n779), .ZN(new_n860));
  OAI21_X1  g674(.A(new_n614), .B1(new_n831), .B2(new_n860), .ZN(new_n861));
  AOI21_X1  g675(.A(new_n861), .B1(new_n841), .B2(new_n759), .ZN(new_n862));
  AND2_X1   g676(.A1(new_n859), .A2(new_n862), .ZN(new_n863));
  AND2_X1   g677(.A1(new_n836), .A2(new_n842), .ZN(new_n864));
  INV_X1    g678(.A(new_n852), .ZN(new_n865));
  NAND3_X1  g679(.A1(new_n864), .A2(new_n865), .A3(KEYINPUT51), .ZN(new_n866));
  NAND2_X1  g680(.A1(new_n863), .A2(new_n866), .ZN(new_n867));
  OAI21_X1  g681(.A(new_n829), .B1(new_n855), .B2(new_n867), .ZN(new_n868));
  NAND2_X1  g682(.A1(new_n852), .A2(new_n844), .ZN(new_n869));
  NAND3_X1  g683(.A1(new_n869), .A2(new_n864), .A3(new_n854), .ZN(new_n870));
  INV_X1    g684(.A(KEYINPUT51), .ZN(new_n871));
  NAND2_X1  g685(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  NAND4_X1  g686(.A1(new_n872), .A2(KEYINPUT120), .A3(new_n866), .A4(new_n863), .ZN(new_n873));
  NAND2_X1  g687(.A1(new_n868), .A2(new_n873), .ZN(new_n874));
  NAND4_X1  g688(.A1(new_n307), .A2(new_n312), .A3(new_n459), .A4(new_n670), .ZN(new_n875));
  INV_X1    g689(.A(KEYINPUT112), .ZN(new_n876));
  AND3_X1   g690(.A1(new_n500), .A2(KEYINPUT93), .A3(new_n505), .ZN(new_n877));
  AOI21_X1  g691(.A(new_n505), .B1(new_n500), .B2(KEYINPUT93), .ZN(new_n878));
  OAI21_X1  g692(.A(new_n876), .B1(new_n877), .B2(new_n878), .ZN(new_n879));
  NAND3_X1  g693(.A1(new_n504), .A2(KEYINPUT112), .A3(new_n506), .ZN(new_n880));
  NAND2_X1  g694(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  INV_X1    g695(.A(new_n881), .ZN(new_n882));
  NOR3_X1   g696(.A1(new_n882), .A2(new_n542), .A3(new_n681), .ZN(new_n883));
  NAND3_X1  g697(.A1(new_n883), .A2(new_n676), .A3(new_n839), .ZN(new_n884));
  NOR2_X1   g698(.A1(new_n875), .A2(new_n884), .ZN(new_n885));
  AOI21_X1  g699(.A(new_n366), .B1(new_n785), .B2(new_n786), .ZN(new_n886));
  AOI21_X1  g700(.A(new_n885), .B1(new_n886), .B2(new_n794), .ZN(new_n887));
  INV_X1    g701(.A(KEYINPUT113), .ZN(new_n888));
  OAI211_X1 g702(.A(new_n888), .B(new_n758), .C1(new_n776), .C2(new_n777), .ZN(new_n889));
  INV_X1    g703(.A(new_n889), .ZN(new_n890));
  NAND2_X1  g704(.A1(new_n785), .A2(new_n786), .ZN(new_n891));
  AOI21_X1  g705(.A(new_n888), .B1(new_n891), .B2(new_n758), .ZN(new_n892));
  OAI21_X1  g706(.A(new_n887), .B1(new_n890), .B2(new_n892), .ZN(new_n893));
  OAI22_X1  g707(.A1(new_n366), .A2(new_n624), .B1(new_n666), .B2(new_n671), .ZN(new_n894));
  AOI211_X1 g708(.A(new_n542), .B(new_n881), .C1(new_n563), .C2(new_n573), .ZN(new_n895));
  OAI21_X1  g709(.A(new_n623), .B1(new_n779), .B2(new_n895), .ZN(new_n896));
  NOR2_X1   g710(.A1(new_n896), .A2(new_n631), .ZN(new_n897));
  NOR2_X1   g711(.A1(new_n894), .A2(new_n897), .ZN(new_n898));
  OAI211_X1 g712(.A(new_n507), .B(new_n645), .C1(new_n752), .C2(new_n542), .ZN(new_n899));
  OAI211_X1 g713(.A(new_n365), .B(new_n754), .C1(new_n755), .C2(new_n756), .ZN(new_n900));
  NOR2_X1   g714(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  AOI22_X1  g715(.A1(new_n736), .A2(new_n901), .B1(new_n712), .B2(new_n733), .ZN(new_n902));
  NAND4_X1  g716(.A1(new_n898), .A2(new_n725), .A3(new_n729), .A4(new_n902), .ZN(new_n903));
  NOR3_X1   g717(.A1(new_n893), .A2(new_n903), .A3(new_n789), .ZN(new_n904));
  NOR4_X1   g718(.A1(new_n670), .A2(new_n457), .A3(new_n508), .A4(new_n681), .ZN(new_n905));
  NOR2_X1   g719(.A1(new_n574), .A2(new_n713), .ZN(new_n906));
  NAND4_X1  g720(.A1(new_n905), .A2(new_n906), .A3(new_n700), .A4(new_n774), .ZN(new_n907));
  NAND4_X1  g721(.A1(new_n688), .A2(new_n715), .A3(new_n760), .A4(new_n907), .ZN(new_n908));
  NAND2_X1  g722(.A1(new_n908), .A2(KEYINPUT52), .ZN(new_n909));
  AOI22_X1  g723(.A1(new_n675), .A2(new_n687), .B1(new_n758), .B2(new_n759), .ZN(new_n910));
  INV_X1    g724(.A(KEYINPUT52), .ZN(new_n911));
  NAND4_X1  g725(.A1(new_n910), .A2(new_n911), .A3(new_n715), .A4(new_n907), .ZN(new_n912));
  NAND2_X1  g726(.A1(new_n909), .A2(new_n912), .ZN(new_n913));
  INV_X1    g727(.A(new_n913), .ZN(new_n914));
  AOI21_X1  g728(.A(KEYINPUT53), .B1(new_n904), .B2(new_n914), .ZN(new_n915));
  INV_X1    g729(.A(new_n885), .ZN(new_n916));
  NAND2_X1  g730(.A1(new_n795), .A2(new_n916), .ZN(new_n917));
  NAND2_X1  g731(.A1(new_n891), .A2(new_n758), .ZN(new_n918));
  NAND2_X1  g732(.A1(new_n918), .A2(KEYINPUT113), .ZN(new_n919));
  AOI21_X1  g733(.A(new_n917), .B1(new_n919), .B2(new_n889), .ZN(new_n920));
  NAND2_X1  g734(.A1(new_n574), .A2(new_n882), .ZN(new_n921));
  NAND2_X1  g735(.A1(new_n860), .A2(new_n921), .ZN(new_n922));
  NAND3_X1  g736(.A1(new_n922), .A2(new_n632), .A3(new_n623), .ZN(new_n923));
  NAND4_X1  g737(.A1(new_n923), .A2(new_n625), .A3(KEYINPUT53), .A4(new_n672), .ZN(new_n924));
  NOR2_X1   g738(.A1(new_n789), .A2(new_n924), .ZN(new_n925));
  INV_X1    g739(.A(KEYINPUT115), .ZN(new_n926));
  NAND3_X1  g740(.A1(new_n725), .A2(new_n746), .A3(new_n734), .ZN(new_n927));
  AND3_X1   g741(.A1(new_n657), .A2(KEYINPUT98), .A3(new_n658), .ZN(new_n928));
  NOR2_X1   g742(.A1(new_n928), .A2(new_n659), .ZN(new_n929));
  NAND2_X1  g743(.A1(new_n721), .A2(new_n723), .ZN(new_n930));
  NOR3_X1   g744(.A1(new_n929), .A2(new_n366), .A3(new_n930), .ZN(new_n931));
  OAI21_X1  g745(.A(new_n926), .B1(new_n927), .B2(new_n931), .ZN(new_n932));
  NAND4_X1  g746(.A1(new_n902), .A2(KEYINPUT115), .A3(new_n729), .A4(new_n725), .ZN(new_n933));
  NAND4_X1  g747(.A1(new_n920), .A2(new_n925), .A3(new_n932), .A4(new_n933), .ZN(new_n934));
  AND3_X1   g748(.A1(new_n909), .A2(KEYINPUT114), .A3(new_n912), .ZN(new_n935));
  AOI21_X1  g749(.A(KEYINPUT114), .B1(new_n909), .B2(new_n912), .ZN(new_n936));
  NOR3_X1   g750(.A1(new_n934), .A2(new_n935), .A3(new_n936), .ZN(new_n937));
  AOI21_X1  g751(.A(new_n915), .B1(new_n937), .B2(KEYINPUT116), .ZN(new_n938));
  INV_X1    g752(.A(KEYINPUT54), .ZN(new_n939));
  INV_X1    g753(.A(KEYINPUT116), .ZN(new_n940));
  INV_X1    g754(.A(KEYINPUT114), .ZN(new_n941));
  NAND2_X1  g755(.A1(new_n913), .A2(new_n941), .ZN(new_n942));
  NAND3_X1  g756(.A1(new_n909), .A2(KEYINPUT114), .A3(new_n912), .ZN(new_n943));
  NAND2_X1  g757(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  OAI21_X1  g758(.A(new_n940), .B1(new_n944), .B2(new_n934), .ZN(new_n945));
  NAND3_X1  g759(.A1(new_n938), .A2(new_n939), .A3(new_n945), .ZN(new_n946));
  NOR2_X1   g760(.A1(new_n935), .A2(new_n936), .ZN(new_n947));
  INV_X1    g761(.A(KEYINPUT53), .ZN(new_n948));
  NAND3_X1  g762(.A1(new_n947), .A2(new_n948), .A3(new_n904), .ZN(new_n949));
  NOR4_X1   g763(.A1(new_n927), .A2(new_n931), .A3(new_n897), .A4(new_n894), .ZN(new_n950));
  NOR2_X1   g764(.A1(new_n753), .A2(new_n856), .ZN(new_n951));
  OAI21_X1  g765(.A(new_n951), .B1(new_n776), .B2(new_n777), .ZN(new_n952));
  NAND2_X1  g766(.A1(new_n952), .A2(KEYINPUT42), .ZN(new_n953));
  NAND4_X1  g767(.A1(new_n920), .A2(new_n950), .A3(new_n953), .A4(new_n778), .ZN(new_n954));
  OAI21_X1  g768(.A(KEYINPUT53), .B1(new_n954), .B2(new_n913), .ZN(new_n955));
  NAND3_X1  g769(.A1(new_n949), .A2(KEYINPUT54), .A3(new_n955), .ZN(new_n956));
  NAND2_X1  g770(.A1(new_n946), .A2(new_n956), .ZN(new_n957));
  OAI22_X1  g771(.A1(new_n874), .A2(new_n957), .B1(G952), .B2(G953), .ZN(new_n958));
  NAND3_X1  g772(.A1(new_n640), .A2(new_n458), .A3(new_n611), .ZN(new_n959));
  NOR3_X1   g773(.A1(new_n692), .A2(new_n691), .A3(new_n959), .ZN(new_n960));
  XOR2_X1   g774(.A(new_n837), .B(KEYINPUT49), .Z(new_n961));
  NAND4_X1  g775(.A1(new_n960), .A2(new_n365), .A3(new_n701), .A4(new_n961), .ZN(new_n962));
  NAND2_X1  g776(.A1(new_n958), .A2(new_n962), .ZN(G75));
  NOR2_X1   g777(.A1(new_n255), .A2(G952), .ZN(new_n964));
  NAND2_X1  g778(.A1(new_n932), .A2(new_n933), .ZN(new_n965));
  NAND4_X1  g779(.A1(new_n898), .A2(new_n953), .A3(KEYINPUT53), .A4(new_n778), .ZN(new_n966));
  NOR3_X1   g780(.A1(new_n965), .A2(new_n893), .A3(new_n966), .ZN(new_n967));
  NAND4_X1  g781(.A1(new_n967), .A2(KEYINPUT116), .A3(new_n943), .A4(new_n942), .ZN(new_n968));
  OAI21_X1  g782(.A(new_n948), .B1(new_n954), .B2(new_n913), .ZN(new_n969));
  NAND2_X1  g783(.A1(new_n968), .A2(new_n969), .ZN(new_n970));
  AOI21_X1  g784(.A(KEYINPUT116), .B1(new_n947), .B2(new_n967), .ZN(new_n971));
  OAI211_X1 g785(.A(G902), .B(new_n608), .C1(new_n970), .C2(new_n971), .ZN(new_n972));
  INV_X1    g786(.A(KEYINPUT56), .ZN(new_n973));
  NAND2_X1  g787(.A1(new_n972), .A2(new_n973), .ZN(new_n974));
  NAND2_X1  g788(.A1(new_n586), .A2(new_n588), .ZN(new_n975));
  XOR2_X1   g789(.A(new_n975), .B(new_n593), .Z(new_n976));
  XNOR2_X1  g790(.A(new_n976), .B(KEYINPUT55), .ZN(new_n977));
  AOI21_X1  g791(.A(new_n964), .B1(new_n974), .B2(new_n977), .ZN(new_n978));
  INV_X1    g792(.A(KEYINPUT121), .ZN(new_n979));
  NAND2_X1  g793(.A1(new_n972), .A2(new_n979), .ZN(new_n980));
  NAND3_X1  g794(.A1(new_n945), .A2(new_n969), .A3(new_n968), .ZN(new_n981));
  NAND4_X1  g795(.A1(new_n981), .A2(KEYINPUT121), .A3(G902), .A4(new_n608), .ZN(new_n982));
  XNOR2_X1  g796(.A(KEYINPUT122), .B(KEYINPUT56), .ZN(new_n983));
  NOR2_X1   g797(.A1(new_n977), .A2(new_n983), .ZN(new_n984));
  NAND3_X1  g798(.A1(new_n980), .A2(new_n982), .A3(new_n984), .ZN(new_n985));
  AND2_X1   g799(.A1(new_n978), .A2(new_n985), .ZN(G51));
  XNOR2_X1  g800(.A(new_n441), .B(KEYINPUT57), .ZN(new_n987));
  AOI21_X1  g801(.A(new_n939), .B1(new_n938), .B2(new_n945), .ZN(new_n988));
  NOR3_X1   g802(.A1(new_n970), .A2(new_n971), .A3(KEYINPUT54), .ZN(new_n989));
  OAI21_X1  g803(.A(new_n987), .B1(new_n988), .B2(new_n989), .ZN(new_n990));
  AND2_X1   g804(.A1(new_n434), .A2(new_n439), .ZN(new_n991));
  NAND2_X1  g805(.A1(new_n990), .A2(new_n991), .ZN(new_n992));
  NAND2_X1  g806(.A1(new_n809), .A2(new_n812), .ZN(new_n993));
  INV_X1    g807(.A(new_n993), .ZN(new_n994));
  OAI211_X1 g808(.A(G902), .B(new_n994), .C1(new_n970), .C2(new_n971), .ZN(new_n995));
  NAND2_X1  g809(.A1(new_n995), .A2(KEYINPUT123), .ZN(new_n996));
  INV_X1    g810(.A(KEYINPUT123), .ZN(new_n997));
  NAND4_X1  g811(.A1(new_n981), .A2(new_n997), .A3(G902), .A4(new_n994), .ZN(new_n998));
  AND2_X1   g812(.A1(new_n996), .A2(new_n998), .ZN(new_n999));
  AOI21_X1  g813(.A(new_n964), .B1(new_n992), .B2(new_n999), .ZN(G54));
  NAND4_X1  g814(.A1(new_n981), .A2(KEYINPUT58), .A3(G475), .A4(G902), .ZN(new_n1001));
  NAND2_X1  g815(.A1(new_n558), .A2(new_n561), .ZN(new_n1002));
  AND2_X1   g816(.A1(new_n1001), .A2(new_n1002), .ZN(new_n1003));
  NOR2_X1   g817(.A1(new_n1001), .A2(new_n1002), .ZN(new_n1004));
  NOR3_X1   g818(.A1(new_n1003), .A2(new_n1004), .A3(new_n964), .ZN(G60));
  NAND2_X1  g819(.A1(G478), .A2(G902), .ZN(new_n1006));
  XNOR2_X1  g820(.A(new_n1006), .B(KEYINPUT59), .ZN(new_n1007));
  AOI21_X1  g821(.A(new_n636), .B1(new_n957), .B2(new_n1007), .ZN(new_n1008));
  NAND2_X1  g822(.A1(new_n636), .A2(new_n1007), .ZN(new_n1009));
  NAND2_X1  g823(.A1(new_n981), .A2(KEYINPUT54), .ZN(new_n1010));
  AOI21_X1  g824(.A(new_n1009), .B1(new_n1010), .B2(new_n946), .ZN(new_n1011));
  NOR3_X1   g825(.A1(new_n1008), .A2(new_n964), .A3(new_n1011), .ZN(G63));
  NAND2_X1  g826(.A1(G217), .A2(G902), .ZN(new_n1013));
  XNOR2_X1  g827(.A(new_n1013), .B(KEYINPUT60), .ZN(new_n1014));
  INV_X1    g828(.A(new_n1014), .ZN(new_n1015));
  NAND3_X1  g829(.A1(new_n981), .A2(new_n668), .A3(new_n1015), .ZN(new_n1016));
  INV_X1    g830(.A(new_n964), .ZN(new_n1017));
  AOI21_X1  g831(.A(new_n1014), .B1(new_n938), .B2(new_n945), .ZN(new_n1018));
  OAI211_X1 g832(.A(new_n1016), .B(new_n1017), .C1(new_n1018), .C2(new_n361), .ZN(new_n1019));
  INV_X1    g833(.A(KEYINPUT61), .ZN(new_n1020));
  NAND2_X1  g834(.A1(new_n1019), .A2(new_n1020), .ZN(new_n1021));
  NAND2_X1  g835(.A1(new_n981), .A2(new_n1015), .ZN(new_n1022));
  INV_X1    g836(.A(new_n361), .ZN(new_n1023));
  AOI21_X1  g837(.A(new_n964), .B1(new_n1022), .B2(new_n1023), .ZN(new_n1024));
  NAND3_X1  g838(.A1(new_n1024), .A2(KEYINPUT61), .A3(new_n1016), .ZN(new_n1025));
  NAND2_X1  g839(.A1(new_n1021), .A2(new_n1025), .ZN(G66));
  OAI21_X1  g840(.A(G953), .B1(new_n621), .B2(new_n591), .ZN(new_n1027));
  OAI21_X1  g841(.A(new_n1027), .B1(new_n950), .B2(new_n618), .ZN(new_n1028));
  OAI21_X1  g842(.A(new_n975), .B1(G898), .B2(new_n255), .ZN(new_n1029));
  XNOR2_X1  g843(.A(new_n1028), .B(new_n1029), .ZN(G69));
  AOI21_X1  g844(.A(new_n827), .B1(new_n807), .B2(new_n818), .ZN(new_n1031));
  NAND3_X1  g845(.A1(new_n910), .A2(new_n795), .A3(new_n715), .ZN(new_n1032));
  NOR3_X1   g846(.A1(new_n816), .A2(new_n899), .A3(new_n856), .ZN(new_n1033));
  NOR3_X1   g847(.A1(new_n1032), .A2(new_n789), .A3(new_n1033), .ZN(new_n1034));
  AND2_X1   g848(.A1(new_n1031), .A2(new_n1034), .ZN(new_n1035));
  NAND2_X1  g849(.A1(new_n1035), .A2(new_n255), .ZN(new_n1036));
  NAND2_X1  g850(.A1(new_n232), .A2(new_n243), .ZN(new_n1037));
  XOR2_X1   g851(.A(new_n1037), .B(KEYINPUT124), .Z(new_n1038));
  XNOR2_X1  g852(.A(new_n1038), .B(new_n555), .ZN(new_n1039));
  INV_X1    g853(.A(new_n1039), .ZN(new_n1040));
  AOI21_X1  g854(.A(new_n1040), .B1(G900), .B2(new_n618), .ZN(new_n1041));
  NAND2_X1  g855(.A1(new_n1036), .A2(new_n1041), .ZN(new_n1042));
  NAND3_X1  g856(.A1(new_n707), .A2(new_n715), .A3(new_n910), .ZN(new_n1043));
  XOR2_X1   g857(.A(new_n1043), .B(KEYINPUT62), .Z(new_n1044));
  NOR2_X1   g858(.A1(new_n704), .A2(new_n808), .ZN(new_n1045));
  NAND3_X1  g859(.A1(new_n1045), .A2(new_n922), .A3(new_n728), .ZN(new_n1046));
  AND3_X1   g860(.A1(new_n1031), .A2(new_n1044), .A3(new_n1046), .ZN(new_n1047));
  OAI21_X1  g861(.A(new_n1040), .B1(new_n1047), .B2(new_n618), .ZN(new_n1048));
  NAND2_X1  g862(.A1(new_n1042), .A2(new_n1048), .ZN(new_n1049));
  AOI21_X1  g863(.A(new_n255), .B1(G227), .B2(G900), .ZN(new_n1050));
  INV_X1    g864(.A(KEYINPUT125), .ZN(new_n1051));
  NAND2_X1  g865(.A1(new_n1050), .A2(new_n1051), .ZN(new_n1052));
  OR2_X1    g866(.A1(new_n1050), .A2(new_n1051), .ZN(new_n1053));
  NAND3_X1  g867(.A1(new_n1049), .A2(new_n1052), .A3(new_n1053), .ZN(new_n1054));
  NAND4_X1  g868(.A1(new_n1042), .A2(new_n1048), .A3(new_n1051), .A4(new_n1050), .ZN(new_n1055));
  AND2_X1   g869(.A1(new_n1054), .A2(new_n1055), .ZN(G72));
  NAND4_X1  g870(.A1(new_n1031), .A2(new_n950), .A3(new_n1044), .A4(new_n1046), .ZN(new_n1057));
  NAND2_X1  g871(.A1(G472), .A2(G902), .ZN(new_n1058));
  XOR2_X1   g872(.A(new_n1058), .B(KEYINPUT63), .Z(new_n1059));
  NAND2_X1  g873(.A1(new_n1057), .A2(new_n1059), .ZN(new_n1060));
  AOI21_X1  g874(.A(new_n268), .B1(new_n244), .B2(new_n246), .ZN(new_n1061));
  NAND2_X1  g875(.A1(new_n1060), .A2(new_n1061), .ZN(new_n1062));
  NAND2_X1  g876(.A1(new_n1062), .A2(KEYINPUT126), .ZN(new_n1063));
  INV_X1    g877(.A(KEYINPUT126), .ZN(new_n1064));
  NAND3_X1  g878(.A1(new_n1060), .A2(new_n1064), .A3(new_n1061), .ZN(new_n1065));
  NAND2_X1  g879(.A1(new_n1063), .A2(new_n1065), .ZN(new_n1066));
  NAND2_X1  g880(.A1(new_n269), .A2(new_n695), .ZN(new_n1067));
  NAND4_X1  g881(.A1(new_n949), .A2(new_n955), .A3(new_n1059), .A4(new_n1067), .ZN(new_n1068));
  XNOR2_X1  g882(.A(new_n1068), .B(KEYINPUT127), .ZN(new_n1069));
  NAND2_X1  g883(.A1(new_n1035), .A2(new_n950), .ZN(new_n1070));
  NAND2_X1  g884(.A1(new_n1070), .A2(new_n1059), .ZN(new_n1071));
  NOR2_X1   g885(.A1(new_n247), .A2(new_n267), .ZN(new_n1072));
  AOI21_X1  g886(.A(new_n964), .B1(new_n1071), .B2(new_n1072), .ZN(new_n1073));
  AND3_X1   g887(.A1(new_n1066), .A2(new_n1069), .A3(new_n1073), .ZN(G57));
endmodule


