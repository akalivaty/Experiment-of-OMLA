//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 0 0 0 0 0 1 1 0 1 0 0 0 0 1 0 1 0 1 1 1 0 0 0 1 0 1 1 0 1 1 0 1 0 0 1 1 1 1 1 0 0 0 0 1 0 1 1 1 1 1 0 0 1 0 1 1 0 0 0 1 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:36:55 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n228, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n236, new_n237, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1228, new_n1229, new_n1230,
    new_n1231, new_n1232, new_n1234, new_n1235, new_n1236, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1302, new_n1303, new_n1304, new_n1305,
    new_n1306;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0005(.A1(G1), .A2(G20), .ZN(new_n206));
  XNOR2_X1  g0006(.A(new_n206), .B(KEYINPUT64), .ZN(new_n207));
  AOI22_X1  g0007(.A1(G68), .A2(G238), .B1(G107), .B2(G264), .ZN(new_n208));
  INV_X1    g0008(.A(G226), .ZN(new_n209));
  INV_X1    g0009(.A(G87), .ZN(new_n210));
  INV_X1    g0010(.A(G250), .ZN(new_n211));
  OAI221_X1 g0011(.A(new_n208), .B1(new_n202), .B2(new_n209), .C1(new_n210), .C2(new_n211), .ZN(new_n212));
  AOI22_X1  g0012(.A1(G77), .A2(G244), .B1(G116), .B2(G270), .ZN(new_n213));
  AOI22_X1  g0013(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n214));
  NAND2_X1  g0014(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  OAI21_X1  g0015(.A(new_n207), .B1(new_n212), .B2(new_n215), .ZN(new_n216));
  XNOR2_X1  g0016(.A(new_n216), .B(KEYINPUT1), .ZN(new_n217));
  NOR2_X1   g0017(.A1(new_n207), .A2(G13), .ZN(new_n218));
  OAI211_X1 g0018(.A(new_n218), .B(G250), .C1(G257), .C2(G264), .ZN(new_n219));
  XOR2_X1   g0019(.A(new_n219), .B(KEYINPUT0), .Z(new_n220));
  NAND2_X1  g0020(.A1(G1), .A2(G13), .ZN(new_n221));
  INV_X1    g0021(.A(G20), .ZN(new_n222));
  NOR2_X1   g0022(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  INV_X1    g0023(.A(new_n201), .ZN(new_n224));
  NAND2_X1  g0024(.A1(new_n224), .A2(G50), .ZN(new_n225));
  INV_X1    g0025(.A(new_n225), .ZN(new_n226));
  AOI211_X1 g0026(.A(new_n217), .B(new_n220), .C1(new_n223), .C2(new_n226), .ZN(G361));
  XNOR2_X1  g0027(.A(G238), .B(G244), .ZN(new_n228));
  XNOR2_X1  g0028(.A(new_n228), .B(G232), .ZN(new_n229));
  XNOR2_X1  g0029(.A(KEYINPUT2), .B(G226), .ZN(new_n230));
  XNOR2_X1  g0030(.A(new_n229), .B(new_n230), .ZN(new_n231));
  XOR2_X1   g0031(.A(G264), .B(G270), .Z(new_n232));
  XNOR2_X1  g0032(.A(G250), .B(G257), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n232), .B(new_n233), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n231), .B(new_n234), .ZN(G358));
  XNOR2_X1  g0035(.A(G68), .B(G77), .ZN(new_n236));
  INV_X1    g0036(.A(G58), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XOR2_X1   g0038(.A(KEYINPUT65), .B(G50), .Z(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XOR2_X1   g0040(.A(G107), .B(G116), .Z(new_n241));
  XNOR2_X1  g0041(.A(G87), .B(G97), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n240), .B(new_n243), .ZN(G351));
  INV_X1    g0044(.A(KEYINPUT67), .ZN(new_n245));
  INV_X1    g0045(.A(KEYINPUT68), .ZN(new_n246));
  NAND3_X1  g0046(.A1(new_n245), .A2(new_n246), .A3(G58), .ZN(new_n247));
  OAI211_X1 g0047(.A(new_n247), .B(KEYINPUT8), .C1(new_n245), .C2(G58), .ZN(new_n248));
  OR3_X1    g0048(.A1(new_n237), .A2(KEYINPUT68), .A3(KEYINPUT8), .ZN(new_n249));
  NAND2_X1  g0049(.A1(new_n248), .A2(new_n249), .ZN(new_n250));
  INV_X1    g0050(.A(G33), .ZN(new_n251));
  NOR2_X1   g0051(.A1(new_n251), .A2(G20), .ZN(new_n252));
  NOR2_X1   g0052(.A1(G20), .A2(G33), .ZN(new_n253));
  AOI22_X1  g0053(.A1(new_n250), .A2(new_n252), .B1(G150), .B2(new_n253), .ZN(new_n254));
  AOI22_X1  g0054(.A1(new_n254), .A2(KEYINPUT69), .B1(G20), .B2(new_n203), .ZN(new_n255));
  OAI21_X1  g0055(.A(new_n255), .B1(KEYINPUT69), .B2(new_n254), .ZN(new_n256));
  OAI21_X1  g0056(.A(new_n221), .B1(new_n206), .B2(new_n251), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  INV_X1    g0058(.A(G1), .ZN(new_n259));
  NAND3_X1  g0059(.A1(new_n259), .A2(G13), .A3(G20), .ZN(new_n260));
  INV_X1    g0060(.A(KEYINPUT70), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  NAND4_X1  g0062(.A1(new_n259), .A2(KEYINPUT70), .A3(G13), .A4(G20), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n262), .A2(new_n263), .ZN(new_n264));
  INV_X1    g0064(.A(new_n257), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  NOR2_X1   g0066(.A1(new_n222), .A2(G1), .ZN(new_n267));
  NOR3_X1   g0067(.A1(new_n266), .A2(new_n202), .A3(new_n267), .ZN(new_n268));
  AND2_X1   g0068(.A1(new_n262), .A2(new_n263), .ZN(new_n269));
  AOI21_X1  g0069(.A(new_n268), .B1(new_n202), .B2(new_n269), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n258), .A2(new_n270), .ZN(new_n271));
  INV_X1    g0071(.A(new_n271), .ZN(new_n272));
  INV_X1    g0072(.A(G41), .ZN(new_n273));
  OAI211_X1 g0073(.A(G1), .B(G13), .C1(new_n251), .C2(new_n273), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n274), .A2(G274), .ZN(new_n275));
  INV_X1    g0075(.A(G45), .ZN(new_n276));
  AOI21_X1  g0076(.A(G1), .B1(new_n273), .B2(new_n276), .ZN(new_n277));
  INV_X1    g0077(.A(new_n277), .ZN(new_n278));
  NOR2_X1   g0078(.A1(new_n275), .A2(new_n278), .ZN(new_n279));
  AOI21_X1  g0079(.A(new_n221), .B1(G33), .B2(G41), .ZN(new_n280));
  NOR2_X1   g0080(.A1(new_n280), .A2(new_n277), .ZN(new_n281));
  XOR2_X1   g0081(.A(KEYINPUT66), .B(G226), .Z(new_n282));
  AND2_X1   g0082(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n251), .A2(KEYINPUT3), .ZN(new_n284));
  INV_X1    g0084(.A(KEYINPUT3), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n285), .A2(G33), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n284), .A2(new_n286), .ZN(new_n287));
  NOR2_X1   g0087(.A1(new_n287), .A2(G1698), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n288), .A2(G222), .ZN(new_n289));
  INV_X1    g0089(.A(G77), .ZN(new_n290));
  XNOR2_X1  g0090(.A(KEYINPUT3), .B(G33), .ZN(new_n291));
  INV_X1    g0091(.A(G223), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n291), .A2(G1698), .ZN(new_n293));
  OAI221_X1 g0093(.A(new_n289), .B1(new_n290), .B2(new_n291), .C1(new_n292), .C2(new_n293), .ZN(new_n294));
  AOI211_X1 g0094(.A(new_n279), .B(new_n283), .C1(new_n294), .C2(new_n280), .ZN(new_n295));
  INV_X1    g0095(.A(G179), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n295), .A2(new_n296), .ZN(new_n297));
  OAI21_X1  g0097(.A(new_n297), .B1(G169), .B2(new_n295), .ZN(new_n298));
  OR2_X1    g0098(.A1(new_n272), .A2(new_n298), .ZN(new_n299));
  INV_X1    g0099(.A(G1698), .ZN(new_n300));
  NAND3_X1  g0100(.A1(new_n291), .A2(G232), .A3(new_n300), .ZN(new_n301));
  INV_X1    g0101(.A(G107), .ZN(new_n302));
  INV_X1    g0102(.A(G238), .ZN(new_n303));
  OAI221_X1 g0103(.A(new_n301), .B1(new_n302), .B2(new_n291), .C1(new_n293), .C2(new_n303), .ZN(new_n304));
  INV_X1    g0104(.A(KEYINPUT71), .ZN(new_n305));
  AOI21_X1  g0105(.A(new_n274), .B1(new_n304), .B2(new_n305), .ZN(new_n306));
  OAI21_X1  g0106(.A(new_n306), .B1(new_n305), .B2(new_n304), .ZN(new_n307));
  AOI21_X1  g0107(.A(new_n279), .B1(G244), .B2(new_n281), .ZN(new_n308));
  AND2_X1   g0108(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  AND2_X1   g0109(.A1(new_n309), .A2(new_n296), .ZN(new_n310));
  INV_X1    g0110(.A(new_n266), .ZN(new_n311));
  INV_X1    g0111(.A(new_n267), .ZN(new_n312));
  NAND3_X1  g0112(.A1(new_n311), .A2(G77), .A3(new_n312), .ZN(new_n313));
  XOR2_X1   g0113(.A(KEYINPUT15), .B(G87), .Z(new_n314));
  INV_X1    g0114(.A(new_n314), .ZN(new_n315));
  INV_X1    g0115(.A(new_n252), .ZN(new_n316));
  NOR2_X1   g0116(.A1(new_n315), .A2(new_n316), .ZN(new_n317));
  XNOR2_X1  g0117(.A(KEYINPUT8), .B(G58), .ZN(new_n318));
  INV_X1    g0118(.A(new_n253), .ZN(new_n319));
  OAI22_X1  g0119(.A1(new_n318), .A2(new_n319), .B1(new_n222), .B2(new_n290), .ZN(new_n320));
  OAI21_X1  g0120(.A(new_n257), .B1(new_n317), .B2(new_n320), .ZN(new_n321));
  OAI211_X1 g0121(.A(new_n313), .B(new_n321), .C1(G77), .C2(new_n264), .ZN(new_n322));
  OAI21_X1  g0122(.A(new_n322), .B1(new_n309), .B2(G169), .ZN(new_n323));
  OR2_X1    g0123(.A1(new_n310), .A2(new_n323), .ZN(new_n324));
  AOI21_X1  g0124(.A(new_n322), .B1(new_n309), .B2(G190), .ZN(new_n325));
  INV_X1    g0125(.A(G200), .ZN(new_n326));
  OAI21_X1  g0126(.A(new_n325), .B1(new_n326), .B2(new_n309), .ZN(new_n327));
  AND2_X1   g0127(.A1(new_n324), .A2(new_n327), .ZN(new_n328));
  XNOR2_X1  g0128(.A(new_n271), .B(KEYINPUT9), .ZN(new_n329));
  INV_X1    g0129(.A(KEYINPUT10), .ZN(new_n330));
  NOR2_X1   g0130(.A1(new_n295), .A2(new_n326), .ZN(new_n331));
  AOI21_X1  g0131(.A(new_n331), .B1(G190), .B2(new_n295), .ZN(new_n332));
  NAND3_X1  g0132(.A1(new_n329), .A2(new_n330), .A3(new_n332), .ZN(new_n333));
  INV_X1    g0133(.A(new_n333), .ZN(new_n334));
  AOI21_X1  g0134(.A(new_n330), .B1(new_n329), .B2(new_n332), .ZN(new_n335));
  OAI211_X1 g0135(.A(new_n299), .B(new_n328), .C1(new_n334), .C2(new_n335), .ZN(new_n336));
  INV_X1    g0136(.A(KEYINPUT72), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n336), .A2(new_n337), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n329), .A2(new_n332), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n339), .A2(KEYINPUT10), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n340), .A2(new_n333), .ZN(new_n341));
  NAND4_X1  g0141(.A1(new_n341), .A2(KEYINPUT72), .A3(new_n299), .A4(new_n328), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n338), .A2(new_n342), .ZN(new_n343));
  INV_X1    g0143(.A(new_n250), .ZN(new_n344));
  NOR2_X1   g0144(.A1(new_n344), .A2(new_n267), .ZN(new_n345));
  AOI22_X1  g0145(.A1(new_n345), .A2(new_n311), .B1(new_n269), .B2(new_n344), .ZN(new_n346));
  INV_X1    g0146(.A(new_n346), .ZN(new_n347));
  INV_X1    g0147(.A(KEYINPUT16), .ZN(new_n348));
  XNOR2_X1  g0148(.A(KEYINPUT67), .B(G58), .ZN(new_n349));
  INV_X1    g0149(.A(G68), .ZN(new_n350));
  OAI21_X1  g0150(.A(new_n224), .B1(new_n349), .B2(new_n350), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n351), .A2(G20), .ZN(new_n352));
  INV_X1    g0152(.A(G159), .ZN(new_n353));
  NOR2_X1   g0153(.A1(new_n319), .A2(new_n353), .ZN(new_n354));
  INV_X1    g0154(.A(new_n354), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n352), .A2(new_n355), .ZN(new_n356));
  INV_X1    g0156(.A(KEYINPUT7), .ZN(new_n357));
  OAI21_X1  g0157(.A(new_n357), .B1(new_n291), .B2(G20), .ZN(new_n358));
  NOR2_X1   g0158(.A1(new_n285), .A2(G33), .ZN(new_n359));
  NOR2_X1   g0159(.A1(new_n251), .A2(KEYINPUT3), .ZN(new_n360));
  OAI211_X1 g0160(.A(KEYINPUT7), .B(new_n222), .C1(new_n359), .C2(new_n360), .ZN(new_n361));
  AOI21_X1  g0161(.A(new_n350), .B1(new_n358), .B2(new_n361), .ZN(new_n362));
  OAI21_X1  g0162(.A(new_n348), .B1(new_n356), .B2(new_n362), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n363), .A2(new_n257), .ZN(new_n364));
  INV_X1    g0164(.A(new_n364), .ZN(new_n365));
  INV_X1    g0165(.A(KEYINPUT75), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n358), .A2(new_n361), .ZN(new_n367));
  AOI21_X1  g0167(.A(new_n366), .B1(new_n367), .B2(G68), .ZN(new_n368));
  AOI211_X1 g0168(.A(KEYINPUT75), .B(new_n350), .C1(new_n358), .C2(new_n361), .ZN(new_n369));
  NOR2_X1   g0169(.A1(new_n368), .A2(new_n369), .ZN(new_n370));
  AOI211_X1 g0170(.A(new_n348), .B(new_n354), .C1(new_n351), .C2(G20), .ZN(new_n371));
  AOI21_X1  g0171(.A(KEYINPUT76), .B1(new_n370), .B2(new_n371), .ZN(new_n372));
  AOI21_X1  g0172(.A(KEYINPUT7), .B1(new_n287), .B2(new_n222), .ZN(new_n373));
  AOI211_X1 g0173(.A(new_n357), .B(G20), .C1(new_n284), .C2(new_n286), .ZN(new_n374));
  OAI21_X1  g0174(.A(G68), .B1(new_n373), .B2(new_n374), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n375), .A2(KEYINPUT75), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n362), .A2(new_n366), .ZN(new_n377));
  NAND4_X1  g0177(.A1(new_n376), .A2(new_n377), .A3(KEYINPUT76), .A4(new_n371), .ZN(new_n378));
  INV_X1    g0178(.A(new_n378), .ZN(new_n379));
  OAI21_X1  g0179(.A(new_n365), .B1(new_n372), .B2(new_n379), .ZN(new_n380));
  INV_X1    g0180(.A(KEYINPUT77), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n380), .A2(new_n381), .ZN(new_n382));
  NAND3_X1  g0182(.A1(new_n376), .A2(new_n377), .A3(new_n371), .ZN(new_n383));
  INV_X1    g0183(.A(KEYINPUT76), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n385), .A2(new_n378), .ZN(new_n386));
  NAND3_X1  g0186(.A1(new_n386), .A2(KEYINPUT77), .A3(new_n365), .ZN(new_n387));
  AOI21_X1  g0187(.A(new_n347), .B1(new_n382), .B2(new_n387), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n291), .A2(new_n300), .ZN(new_n389));
  OAI22_X1  g0189(.A1(new_n389), .A2(new_n292), .B1(new_n251), .B2(new_n210), .ZN(new_n390));
  NOR2_X1   g0190(.A1(new_n293), .A2(new_n209), .ZN(new_n391));
  OAI21_X1  g0191(.A(new_n280), .B1(new_n390), .B2(new_n391), .ZN(new_n392));
  AOI21_X1  g0192(.A(new_n279), .B1(G232), .B2(new_n281), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n392), .A2(new_n393), .ZN(new_n394));
  NOR2_X1   g0194(.A1(new_n394), .A2(new_n296), .ZN(new_n395));
  AOI21_X1  g0195(.A(new_n395), .B1(G169), .B2(new_n394), .ZN(new_n396));
  NOR3_X1   g0196(.A1(new_n388), .A2(new_n396), .A3(KEYINPUT18), .ZN(new_n397));
  INV_X1    g0197(.A(KEYINPUT18), .ZN(new_n398));
  AOI21_X1  g0198(.A(KEYINPUT77), .B1(new_n386), .B2(new_n365), .ZN(new_n399));
  AOI211_X1 g0199(.A(new_n381), .B(new_n364), .C1(new_n385), .C2(new_n378), .ZN(new_n400));
  OAI21_X1  g0200(.A(new_n346), .B1(new_n399), .B2(new_n400), .ZN(new_n401));
  INV_X1    g0201(.A(new_n396), .ZN(new_n402));
  AOI21_X1  g0202(.A(new_n398), .B1(new_n401), .B2(new_n402), .ZN(new_n403));
  NOR2_X1   g0203(.A1(new_n397), .A2(new_n403), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n394), .A2(new_n326), .ZN(new_n405));
  OAI21_X1  g0205(.A(new_n405), .B1(G190), .B2(new_n394), .ZN(new_n406));
  OAI211_X1 g0206(.A(new_n346), .B(new_n406), .C1(new_n399), .C2(new_n400), .ZN(new_n407));
  INV_X1    g0207(.A(KEYINPUT17), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n407), .A2(new_n408), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n382), .A2(new_n387), .ZN(new_n410));
  NAND4_X1  g0210(.A1(new_n410), .A2(KEYINPUT17), .A3(new_n346), .A4(new_n406), .ZN(new_n411));
  AND2_X1   g0211(.A1(new_n409), .A2(new_n411), .ZN(new_n412));
  NAND3_X1  g0212(.A1(new_n404), .A2(new_n412), .A3(KEYINPUT78), .ZN(new_n413));
  NAND3_X1  g0213(.A1(new_n291), .A2(G232), .A3(G1698), .ZN(new_n414));
  NAND2_X1  g0214(.A1(G33), .A2(G97), .ZN(new_n415));
  OAI211_X1 g0215(.A(new_n414), .B(new_n415), .C1(new_n389), .C2(new_n209), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n416), .A2(new_n280), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n281), .A2(G238), .ZN(new_n418));
  OAI211_X1 g0218(.A(new_n417), .B(new_n418), .C1(new_n278), .C2(new_n275), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n419), .A2(KEYINPUT13), .ZN(new_n420));
  AOI21_X1  g0220(.A(new_n279), .B1(G238), .B2(new_n281), .ZN(new_n421));
  INV_X1    g0221(.A(KEYINPUT13), .ZN(new_n422));
  NAND3_X1  g0222(.A1(new_n421), .A2(new_n417), .A3(new_n422), .ZN(new_n423));
  INV_X1    g0223(.A(KEYINPUT73), .ZN(new_n424));
  NAND3_X1  g0224(.A1(new_n420), .A2(new_n423), .A3(new_n424), .ZN(new_n425));
  NAND3_X1  g0225(.A1(new_n419), .A2(KEYINPUT73), .A3(KEYINPUT13), .ZN(new_n426));
  AND2_X1   g0226(.A1(new_n425), .A2(new_n426), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n427), .A2(G200), .ZN(new_n428));
  OAI22_X1  g0228(.A1(new_n316), .A2(new_n290), .B1(new_n222), .B2(G68), .ZN(new_n429));
  NOR2_X1   g0229(.A1(new_n319), .A2(new_n202), .ZN(new_n430));
  OAI21_X1  g0230(.A(new_n257), .B1(new_n429), .B2(new_n430), .ZN(new_n431));
  XNOR2_X1  g0231(.A(new_n431), .B(KEYINPUT11), .ZN(new_n432));
  NAND3_X1  g0232(.A1(new_n311), .A2(G68), .A3(new_n312), .ZN(new_n433));
  OAI22_X1  g0233(.A1(new_n264), .A2(G68), .B1(KEYINPUT74), .B2(KEYINPUT12), .ZN(new_n434));
  NAND2_X1  g0234(.A1(KEYINPUT74), .A2(KEYINPUT12), .ZN(new_n435));
  XNOR2_X1  g0235(.A(new_n434), .B(new_n435), .ZN(new_n436));
  NAND3_X1  g0236(.A1(new_n432), .A2(new_n433), .A3(new_n436), .ZN(new_n437));
  INV_X1    g0237(.A(new_n420), .ZN(new_n438));
  INV_X1    g0238(.A(G190), .ZN(new_n439));
  NOR2_X1   g0239(.A1(new_n438), .A2(new_n439), .ZN(new_n440));
  AOI21_X1  g0240(.A(new_n437), .B1(new_n440), .B2(new_n423), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n428), .A2(new_n441), .ZN(new_n442));
  INV_X1    g0242(.A(new_n423), .ZN(new_n443));
  NOR3_X1   g0243(.A1(new_n438), .A2(new_n296), .A3(new_n443), .ZN(new_n444));
  NAND3_X1  g0244(.A1(new_n427), .A2(KEYINPUT14), .A3(G169), .ZN(new_n445));
  NAND3_X1  g0245(.A1(new_n425), .A2(G169), .A3(new_n426), .ZN(new_n446));
  INV_X1    g0246(.A(KEYINPUT14), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n446), .A2(new_n447), .ZN(new_n448));
  AOI21_X1  g0248(.A(new_n444), .B1(new_n445), .B2(new_n448), .ZN(new_n449));
  INV_X1    g0249(.A(new_n437), .ZN(new_n450));
  OAI21_X1  g0250(.A(new_n442), .B1(new_n449), .B2(new_n450), .ZN(new_n451));
  INV_X1    g0251(.A(KEYINPUT78), .ZN(new_n452));
  OAI21_X1  g0252(.A(KEYINPUT18), .B1(new_n388), .B2(new_n396), .ZN(new_n453));
  NAND3_X1  g0253(.A1(new_n401), .A2(new_n398), .A3(new_n402), .ZN(new_n454));
  NAND4_X1  g0254(.A1(new_n453), .A2(new_n454), .A3(new_n409), .A4(new_n411), .ZN(new_n455));
  AOI21_X1  g0255(.A(new_n451), .B1(new_n452), .B2(new_n455), .ZN(new_n456));
  NAND3_X1  g0256(.A1(new_n343), .A2(new_n413), .A3(new_n456), .ZN(new_n457));
  INV_X1    g0257(.A(new_n457), .ZN(new_n458));
  NAND4_X1  g0258(.A1(new_n284), .A2(new_n286), .A3(G264), .A4(G1698), .ZN(new_n459));
  NAND4_X1  g0259(.A1(new_n284), .A2(new_n286), .A3(G257), .A4(new_n300), .ZN(new_n460));
  INV_X1    g0260(.A(G303), .ZN(new_n461));
  OAI211_X1 g0261(.A(new_n459), .B(new_n460), .C1(new_n461), .C2(new_n291), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n462), .A2(new_n280), .ZN(new_n463));
  OAI211_X1 g0263(.A(new_n259), .B(G45), .C1(new_n273), .C2(KEYINPUT5), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n464), .A2(KEYINPUT81), .ZN(new_n465));
  INV_X1    g0265(.A(new_n465), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n273), .A2(KEYINPUT5), .ZN(new_n467));
  OAI21_X1  g0267(.A(new_n467), .B1(new_n464), .B2(KEYINPUT81), .ZN(new_n468));
  OAI211_X1 g0268(.A(G270), .B(new_n274), .C1(new_n466), .C2(new_n468), .ZN(new_n469));
  AND2_X1   g0269(.A1(new_n274), .A2(G274), .ZN(new_n470));
  OR2_X1    g0270(.A1(new_n464), .A2(KEYINPUT81), .ZN(new_n471));
  NAND4_X1  g0271(.A1(new_n470), .A2(new_n471), .A3(new_n465), .A4(new_n467), .ZN(new_n472));
  NAND3_X1  g0272(.A1(new_n463), .A2(new_n469), .A3(new_n472), .ZN(new_n473));
  INV_X1    g0273(.A(KEYINPUT85), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  NAND4_X1  g0275(.A1(new_n463), .A2(new_n469), .A3(new_n472), .A4(KEYINPUT85), .ZN(new_n476));
  AND2_X1   g0276(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  NAND2_X1  g0277(.A1(G33), .A2(G283), .ZN(new_n478));
  INV_X1    g0278(.A(G97), .ZN(new_n479));
  OAI211_X1 g0279(.A(new_n478), .B(new_n222), .C1(G33), .C2(new_n479), .ZN(new_n480));
  OAI211_X1 g0280(.A(new_n480), .B(new_n257), .C1(new_n222), .C2(G116), .ZN(new_n481));
  INV_X1    g0281(.A(KEYINPUT20), .ZN(new_n482));
  OR3_X1    g0282(.A1(new_n481), .A2(KEYINPUT86), .A3(new_n482), .ZN(new_n483));
  OAI21_X1  g0283(.A(KEYINPUT86), .B1(new_n481), .B2(new_n482), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n481), .A2(new_n482), .ZN(new_n485));
  NAND3_X1  g0285(.A1(new_n483), .A2(new_n484), .A3(new_n485), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n259), .A2(G33), .ZN(new_n487));
  NAND3_X1  g0287(.A1(new_n311), .A2(G116), .A3(new_n487), .ZN(new_n488));
  INV_X1    g0288(.A(G116), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n269), .A2(new_n489), .ZN(new_n490));
  NAND3_X1  g0290(.A1(new_n486), .A2(new_n488), .A3(new_n490), .ZN(new_n491));
  NAND3_X1  g0291(.A1(new_n477), .A2(G169), .A3(new_n491), .ZN(new_n492));
  INV_X1    g0292(.A(KEYINPUT21), .ZN(new_n493));
  AOI21_X1  g0293(.A(KEYINPUT87), .B1(new_n492), .B2(new_n493), .ZN(new_n494));
  INV_X1    g0294(.A(new_n494), .ZN(new_n495));
  NAND3_X1  g0295(.A1(new_n492), .A2(KEYINPUT87), .A3(new_n493), .ZN(new_n496));
  NAND3_X1  g0296(.A1(new_n477), .A2(KEYINPUT21), .A3(G169), .ZN(new_n497));
  NOR2_X1   g0297(.A1(new_n473), .A2(new_n296), .ZN(new_n498));
  INV_X1    g0298(.A(new_n498), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n497), .A2(new_n499), .ZN(new_n500));
  AOI22_X1  g0300(.A1(new_n495), .A2(new_n496), .B1(new_n500), .B2(new_n491), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n475), .A2(new_n476), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n502), .A2(G190), .ZN(new_n503));
  INV_X1    g0303(.A(new_n491), .ZN(new_n504));
  OAI211_X1 g0304(.A(new_n503), .B(new_n504), .C1(new_n326), .C2(new_n502), .ZN(new_n505));
  INV_X1    g0305(.A(KEYINPUT88), .ZN(new_n506));
  XNOR2_X1  g0306(.A(new_n505), .B(new_n506), .ZN(new_n507));
  AND2_X1   g0307(.A1(new_n501), .A2(new_n507), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n253), .A2(G77), .ZN(new_n509));
  XNOR2_X1  g0309(.A(G97), .B(G107), .ZN(new_n510));
  INV_X1    g0310(.A(KEYINPUT79), .ZN(new_n511));
  OAI21_X1  g0311(.A(new_n510), .B1(new_n511), .B2(KEYINPUT6), .ZN(new_n512));
  MUX2_X1   g0312(.A(new_n511), .B(G97), .S(KEYINPUT6), .Z(new_n513));
  OAI21_X1  g0313(.A(new_n512), .B1(new_n510), .B2(new_n513), .ZN(new_n514));
  OAI21_X1  g0314(.A(new_n509), .B1(new_n514), .B2(new_n222), .ZN(new_n515));
  AOI21_X1  g0315(.A(new_n302), .B1(new_n358), .B2(new_n361), .ZN(new_n516));
  OAI21_X1  g0316(.A(new_n257), .B1(new_n515), .B2(new_n516), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n269), .A2(new_n479), .ZN(new_n518));
  AND2_X1   g0318(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n311), .A2(new_n487), .ZN(new_n520));
  INV_X1    g0320(.A(KEYINPUT80), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  NAND3_X1  g0322(.A1(new_n311), .A2(KEYINPUT80), .A3(new_n487), .ZN(new_n523));
  NAND3_X1  g0323(.A1(new_n522), .A2(G97), .A3(new_n523), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n519), .A2(new_n524), .ZN(new_n525));
  NAND3_X1  g0325(.A1(new_n288), .A2(KEYINPUT4), .A3(G244), .ZN(new_n526));
  OAI211_X1 g0326(.A(new_n526), .B(new_n478), .C1(new_n211), .C2(new_n293), .ZN(new_n527));
  AOI21_X1  g0327(.A(KEYINPUT4), .B1(new_n288), .B2(G244), .ZN(new_n528));
  OAI21_X1  g0328(.A(new_n280), .B1(new_n527), .B2(new_n528), .ZN(new_n529));
  OAI211_X1 g0329(.A(G257), .B(new_n274), .C1(new_n466), .C2(new_n468), .ZN(new_n530));
  AND2_X1   g0330(.A1(new_n530), .A2(new_n472), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n529), .A2(new_n531), .ZN(new_n532));
  NOR2_X1   g0332(.A1(new_n532), .A2(new_n296), .ZN(new_n533));
  INV_X1    g0333(.A(G169), .ZN(new_n534));
  AOI21_X1  g0334(.A(new_n534), .B1(new_n529), .B2(new_n531), .ZN(new_n535));
  OAI21_X1  g0335(.A(new_n525), .B1(new_n533), .B2(new_n535), .ZN(new_n536));
  NAND3_X1  g0336(.A1(new_n522), .A2(G107), .A3(new_n523), .ZN(new_n537));
  NOR2_X1   g0337(.A1(new_n264), .A2(G107), .ZN(new_n538));
  XNOR2_X1  g0338(.A(new_n538), .B(KEYINPUT25), .ZN(new_n539));
  AND2_X1   g0339(.A1(new_n537), .A2(new_n539), .ZN(new_n540));
  NAND4_X1  g0340(.A1(new_n291), .A2(KEYINPUT89), .A3(new_n222), .A4(G87), .ZN(new_n541));
  INV_X1    g0341(.A(KEYINPUT22), .ZN(new_n542));
  OR2_X1    g0342(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n541), .A2(new_n542), .ZN(new_n544));
  INV_X1    g0344(.A(KEYINPUT23), .ZN(new_n545));
  OAI21_X1  g0345(.A(new_n545), .B1(new_n222), .B2(G107), .ZN(new_n546));
  NAND3_X1  g0346(.A1(new_n302), .A2(KEYINPUT23), .A3(G20), .ZN(new_n547));
  NOR2_X1   g0347(.A1(new_n251), .A2(new_n489), .ZN(new_n548));
  AOI22_X1  g0348(.A1(new_n546), .A2(new_n547), .B1(new_n548), .B2(new_n222), .ZN(new_n549));
  NAND3_X1  g0349(.A1(new_n543), .A2(new_n544), .A3(new_n549), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n550), .A2(KEYINPUT24), .ZN(new_n551));
  INV_X1    g0351(.A(KEYINPUT24), .ZN(new_n552));
  NAND4_X1  g0352(.A1(new_n543), .A2(new_n552), .A3(new_n544), .A4(new_n549), .ZN(new_n553));
  AOI21_X1  g0353(.A(new_n265), .B1(new_n551), .B2(new_n553), .ZN(new_n554));
  INV_X1    g0354(.A(new_n554), .ZN(new_n555));
  NAND3_X1  g0355(.A1(new_n291), .A2(G257), .A3(G1698), .ZN(new_n556));
  INV_X1    g0356(.A(G294), .ZN(new_n557));
  OAI221_X1 g0357(.A(new_n556), .B1(new_n251), .B2(new_n557), .C1(new_n389), .C2(new_n211), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n558), .A2(new_n280), .ZN(new_n559));
  OAI211_X1 g0359(.A(G264), .B(new_n274), .C1(new_n466), .C2(new_n468), .ZN(new_n560));
  NAND3_X1  g0360(.A1(new_n559), .A2(new_n472), .A3(new_n560), .ZN(new_n561));
  INV_X1    g0361(.A(new_n561), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n562), .A2(G190), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n561), .A2(G200), .ZN(new_n564));
  NAND4_X1  g0364(.A1(new_n540), .A2(new_n555), .A3(new_n563), .A4(new_n564), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n532), .A2(G200), .ZN(new_n566));
  NAND3_X1  g0366(.A1(new_n529), .A2(G190), .A3(new_n531), .ZN(new_n567));
  NAND4_X1  g0367(.A1(new_n566), .A2(new_n519), .A3(new_n524), .A4(new_n567), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n562), .A2(new_n296), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n561), .A2(new_n534), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n537), .A2(new_n539), .ZN(new_n571));
  OAI211_X1 g0371(.A(new_n569), .B(new_n570), .C1(new_n571), .C2(new_n554), .ZN(new_n572));
  NAND4_X1  g0372(.A1(new_n536), .A2(new_n565), .A3(new_n568), .A4(new_n572), .ZN(new_n573));
  NOR2_X1   g0373(.A1(new_n276), .A2(G1), .ZN(new_n574));
  NOR3_X1   g0374(.A1(new_n280), .A2(new_n211), .A3(new_n574), .ZN(new_n575));
  INV_X1    g0375(.A(KEYINPUT82), .ZN(new_n576));
  INV_X1    g0376(.A(new_n574), .ZN(new_n577));
  OAI21_X1  g0377(.A(new_n576), .B1(new_n275), .B2(new_n577), .ZN(new_n578));
  NAND4_X1  g0378(.A1(new_n274), .A2(KEYINPUT82), .A3(G274), .A4(new_n574), .ZN(new_n579));
  AOI21_X1  g0379(.A(new_n575), .B1(new_n578), .B2(new_n579), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n303), .A2(new_n300), .ZN(new_n581));
  INV_X1    g0381(.A(G244), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n582), .A2(G1698), .ZN(new_n583));
  NAND3_X1  g0383(.A1(new_n291), .A2(new_n581), .A3(new_n583), .ZN(new_n584));
  INV_X1    g0384(.A(new_n548), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n586), .A2(new_n280), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n580), .A2(new_n587), .ZN(new_n588));
  NOR2_X1   g0388(.A1(new_n588), .A2(G179), .ZN(new_n589));
  AOI21_X1  g0389(.A(new_n589), .B1(new_n534), .B2(new_n588), .ZN(new_n590));
  NAND3_X1  g0390(.A1(new_n522), .A2(new_n314), .A3(new_n523), .ZN(new_n591));
  INV_X1    g0391(.A(KEYINPUT84), .ZN(new_n592));
  XOR2_X1   g0392(.A(KEYINPUT83), .B(G87), .Z(new_n593));
  NAND3_X1  g0393(.A1(new_n593), .A2(new_n479), .A3(new_n302), .ZN(new_n594));
  INV_X1    g0394(.A(KEYINPUT19), .ZN(new_n595));
  OAI21_X1  g0395(.A(new_n222), .B1(new_n415), .B2(new_n595), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n594), .A2(new_n596), .ZN(new_n597));
  NAND3_X1  g0397(.A1(new_n291), .A2(new_n222), .A3(G68), .ZN(new_n598));
  OAI21_X1  g0398(.A(new_n595), .B1(new_n316), .B2(new_n479), .ZN(new_n599));
  NAND3_X1  g0399(.A1(new_n597), .A2(new_n598), .A3(new_n599), .ZN(new_n600));
  AOI22_X1  g0400(.A1(new_n600), .A2(new_n257), .B1(new_n269), .B2(new_n315), .ZN(new_n601));
  AND3_X1   g0401(.A1(new_n591), .A2(new_n592), .A3(new_n601), .ZN(new_n602));
  AOI21_X1  g0402(.A(new_n592), .B1(new_n591), .B2(new_n601), .ZN(new_n603));
  OAI21_X1  g0403(.A(new_n590), .B1(new_n602), .B2(new_n603), .ZN(new_n604));
  INV_X1    g0404(.A(new_n588), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n605), .A2(G190), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n588), .A2(G200), .ZN(new_n607));
  NAND3_X1  g0407(.A1(new_n522), .A2(G87), .A3(new_n523), .ZN(new_n608));
  NAND4_X1  g0408(.A1(new_n606), .A2(new_n607), .A3(new_n608), .A4(new_n601), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n604), .A2(new_n609), .ZN(new_n610));
  NOR2_X1   g0410(.A1(new_n573), .A2(new_n610), .ZN(new_n611));
  AND3_X1   g0411(.A1(new_n458), .A2(new_n508), .A3(new_n611), .ZN(G372));
  NAND2_X1  g0412(.A1(new_n500), .A2(new_n491), .ZN(new_n613));
  INV_X1    g0413(.A(new_n496), .ZN(new_n614));
  OAI211_X1 g0414(.A(new_n613), .B(new_n572), .C1(new_n614), .C2(new_n494), .ZN(new_n615));
  NAND3_X1  g0415(.A1(new_n536), .A2(new_n565), .A3(new_n568), .ZN(new_n616));
  INV_X1    g0416(.A(new_n616), .ZN(new_n617));
  AOI21_X1  g0417(.A(KEYINPUT90), .B1(new_n586), .B2(new_n280), .ZN(new_n618));
  INV_X1    g0418(.A(KEYINPUT90), .ZN(new_n619));
  AOI211_X1 g0419(.A(new_n619), .B(new_n274), .C1(new_n584), .C2(new_n585), .ZN(new_n620));
  OAI21_X1  g0420(.A(new_n580), .B1(new_n618), .B2(new_n620), .ZN(new_n621));
  AOI21_X1  g0421(.A(new_n589), .B1(new_n534), .B2(new_n621), .ZN(new_n622));
  OAI21_X1  g0422(.A(new_n622), .B1(new_n602), .B2(new_n603), .ZN(new_n623));
  NAND3_X1  g0423(.A1(new_n606), .A2(new_n608), .A3(new_n601), .ZN(new_n624));
  INV_X1    g0424(.A(new_n621), .ZN(new_n625));
  NOR2_X1   g0425(.A1(new_n625), .A2(new_n326), .ZN(new_n626));
  OAI21_X1  g0426(.A(new_n623), .B1(new_n624), .B2(new_n626), .ZN(new_n627));
  INV_X1    g0427(.A(new_n627), .ZN(new_n628));
  NAND3_X1  g0428(.A1(new_n615), .A2(new_n617), .A3(new_n628), .ZN(new_n629));
  INV_X1    g0429(.A(KEYINPUT26), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n532), .A2(G169), .ZN(new_n631));
  OAI211_X1 g0431(.A(new_n631), .B(KEYINPUT91), .C1(new_n296), .C2(new_n532), .ZN(new_n632));
  INV_X1    g0432(.A(new_n525), .ZN(new_n633));
  AND2_X1   g0433(.A1(new_n529), .A2(new_n531), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n634), .A2(G179), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n635), .A2(new_n631), .ZN(new_n636));
  INV_X1    g0436(.A(KEYINPUT91), .ZN(new_n637));
  AOI21_X1  g0437(.A(new_n633), .B1(new_n636), .B2(new_n637), .ZN(new_n638));
  NAND4_X1  g0438(.A1(new_n628), .A2(new_n630), .A3(new_n632), .A4(new_n638), .ZN(new_n639));
  INV_X1    g0439(.A(new_n623), .ZN(new_n640));
  INV_X1    g0440(.A(new_n536), .ZN(new_n641));
  NAND3_X1  g0441(.A1(new_n641), .A2(new_n609), .A3(new_n604), .ZN(new_n642));
  AOI21_X1  g0442(.A(new_n640), .B1(new_n642), .B2(KEYINPUT26), .ZN(new_n643));
  NAND3_X1  g0443(.A1(new_n629), .A2(new_n639), .A3(new_n643), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n458), .A2(new_n644), .ZN(new_n645));
  INV_X1    g0445(.A(new_n299), .ZN(new_n646));
  AND3_X1   g0446(.A1(new_n453), .A2(KEYINPUT92), .A3(new_n454), .ZN(new_n647));
  AOI21_X1  g0447(.A(KEYINPUT92), .B1(new_n453), .B2(new_n454), .ZN(new_n648));
  NOR2_X1   g0448(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  INV_X1    g0449(.A(new_n649), .ZN(new_n650));
  INV_X1    g0450(.A(new_n442), .ZN(new_n651));
  OAI22_X1  g0451(.A1(new_n651), .A2(new_n324), .B1(new_n449), .B2(new_n450), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n652), .A2(new_n412), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n650), .A2(new_n653), .ZN(new_n654));
  AOI21_X1  g0454(.A(new_n646), .B1(new_n654), .B2(new_n341), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n645), .A2(new_n655), .ZN(G369));
  INV_X1    g0456(.A(new_n501), .ZN(new_n657));
  NAND3_X1  g0457(.A1(new_n259), .A2(new_n222), .A3(G13), .ZN(new_n658));
  OR2_X1    g0458(.A1(new_n658), .A2(KEYINPUT27), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n658), .A2(KEYINPUT27), .ZN(new_n660));
  NAND3_X1  g0460(.A1(new_n659), .A2(G213), .A3(new_n660), .ZN(new_n661));
  INV_X1    g0461(.A(G343), .ZN(new_n662));
  NOR2_X1   g0462(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  INV_X1    g0463(.A(new_n663), .ZN(new_n664));
  NOR2_X1   g0464(.A1(new_n504), .A2(new_n664), .ZN(new_n665));
  MUX2_X1   g0465(.A(new_n508), .B(new_n657), .S(new_n665), .Z(new_n666));
  NOR2_X1   g0466(.A1(new_n572), .A2(new_n663), .ZN(new_n667));
  OAI21_X1  g0467(.A(new_n663), .B1(new_n571), .B2(new_n554), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n565), .A2(new_n668), .ZN(new_n669));
  AOI21_X1  g0469(.A(new_n667), .B1(new_n669), .B2(new_n572), .ZN(new_n670));
  NAND3_X1  g0470(.A1(new_n666), .A2(G330), .A3(new_n670), .ZN(new_n671));
  NOR2_X1   g0471(.A1(new_n501), .A2(new_n663), .ZN(new_n672));
  AOI21_X1  g0472(.A(new_n667), .B1(new_n672), .B2(new_n670), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n671), .A2(new_n673), .ZN(G399));
  NOR3_X1   g0474(.A1(new_n594), .A2(new_n259), .A3(G116), .ZN(new_n675));
  INV_X1    g0475(.A(new_n218), .ZN(new_n676));
  NOR2_X1   g0476(.A1(new_n676), .A2(G41), .ZN(new_n677));
  MUX2_X1   g0477(.A(new_n675), .B(new_n226), .S(new_n677), .Z(new_n678));
  XNOR2_X1  g0478(.A(new_n678), .B(KEYINPUT28), .ZN(new_n679));
  INV_X1    g0479(.A(G330), .ZN(new_n680));
  AND4_X1   g0480(.A1(new_n501), .A2(new_n611), .A3(new_n507), .A4(new_n664), .ZN(new_n681));
  INV_X1    g0481(.A(KEYINPUT94), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n621), .A2(KEYINPUT93), .ZN(new_n683));
  INV_X1    g0483(.A(KEYINPUT93), .ZN(new_n684));
  OAI211_X1 g0484(.A(new_n580), .B(new_n684), .C1(new_n618), .C2(new_n620), .ZN(new_n685));
  NAND3_X1  g0485(.A1(new_n683), .A2(new_n296), .A3(new_n685), .ZN(new_n686));
  OAI21_X1  g0486(.A(new_n682), .B1(new_n686), .B2(new_n502), .ZN(new_n687));
  AND2_X1   g0487(.A1(new_n685), .A2(new_n296), .ZN(new_n688));
  NAND4_X1  g0488(.A1(new_n477), .A2(new_n688), .A3(KEYINPUT94), .A4(new_n683), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n687), .A2(new_n689), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n532), .A2(new_n561), .ZN(new_n691));
  INV_X1    g0491(.A(new_n691), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n690), .A2(new_n692), .ZN(new_n693));
  AND2_X1   g0493(.A1(new_n559), .A2(new_n560), .ZN(new_n694));
  AND2_X1   g0494(.A1(new_n694), .A2(new_n605), .ZN(new_n695));
  NAND4_X1  g0495(.A1(new_n695), .A2(KEYINPUT30), .A3(new_n634), .A4(new_n498), .ZN(new_n696));
  INV_X1    g0496(.A(KEYINPUT30), .ZN(new_n697));
  NAND4_X1  g0497(.A1(new_n694), .A2(new_n605), .A3(new_n529), .A4(new_n531), .ZN(new_n698));
  OAI21_X1  g0498(.A(new_n697), .B1(new_n698), .B2(new_n499), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n696), .A2(new_n699), .ZN(new_n700));
  INV_X1    g0500(.A(new_n700), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n693), .A2(new_n701), .ZN(new_n702));
  NAND4_X1  g0502(.A1(new_n702), .A2(KEYINPUT95), .A3(KEYINPUT31), .A4(new_n663), .ZN(new_n703));
  AOI21_X1  g0503(.A(new_n691), .B1(new_n687), .B2(new_n689), .ZN(new_n704));
  OAI211_X1 g0504(.A(KEYINPUT31), .B(new_n663), .C1(new_n704), .C2(new_n700), .ZN(new_n705));
  INV_X1    g0505(.A(KEYINPUT95), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  OAI21_X1  g0507(.A(new_n663), .B1(new_n704), .B2(new_n700), .ZN(new_n708));
  INV_X1    g0508(.A(KEYINPUT31), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  NAND3_X1  g0510(.A1(new_n703), .A2(new_n707), .A3(new_n710), .ZN(new_n711));
  INV_X1    g0511(.A(KEYINPUT96), .ZN(new_n712));
  AOI21_X1  g0512(.A(new_n681), .B1(new_n711), .B2(new_n712), .ZN(new_n713));
  NAND4_X1  g0513(.A1(new_n703), .A2(new_n707), .A3(KEYINPUT96), .A4(new_n710), .ZN(new_n714));
  AOI21_X1  g0514(.A(new_n680), .B1(new_n713), .B2(new_n714), .ZN(new_n715));
  INV_X1    g0515(.A(KEYINPUT29), .ZN(new_n716));
  NAND3_X1  g0516(.A1(new_n644), .A2(new_n716), .A3(new_n664), .ZN(new_n717));
  OAI21_X1  g0517(.A(new_n637), .B1(new_n533), .B2(new_n535), .ZN(new_n718));
  NAND3_X1  g0518(.A1(new_n718), .A2(new_n632), .A3(new_n525), .ZN(new_n719));
  OAI21_X1  g0519(.A(KEYINPUT26), .B1(new_n627), .B2(new_n719), .ZN(new_n720));
  NAND4_X1  g0520(.A1(new_n641), .A2(new_n604), .A3(new_n630), .A4(new_n609), .ZN(new_n721));
  AND3_X1   g0521(.A1(new_n720), .A2(new_n623), .A3(new_n721), .ZN(new_n722));
  AOI21_X1  g0522(.A(new_n663), .B1(new_n722), .B2(new_n629), .ZN(new_n723));
  OAI21_X1  g0523(.A(new_n717), .B1(new_n723), .B2(new_n716), .ZN(new_n724));
  OR2_X1    g0524(.A1(new_n715), .A2(new_n724), .ZN(new_n725));
  XNOR2_X1  g0525(.A(new_n725), .B(KEYINPUT97), .ZN(new_n726));
  INV_X1    g0526(.A(new_n726), .ZN(new_n727));
  OAI21_X1  g0527(.A(new_n679), .B1(new_n727), .B2(G1), .ZN(G364));
  INV_X1    g0528(.A(new_n677), .ZN(new_n729));
  INV_X1    g0529(.A(G13), .ZN(new_n730));
  NOR2_X1   g0530(.A1(new_n730), .A2(G20), .ZN(new_n731));
  AOI21_X1  g0531(.A(new_n259), .B1(new_n731), .B2(G45), .ZN(new_n732));
  NAND3_X1  g0532(.A1(new_n729), .A2(KEYINPUT98), .A3(new_n732), .ZN(new_n733));
  INV_X1    g0533(.A(KEYINPUT98), .ZN(new_n734));
  INV_X1    g0534(.A(new_n732), .ZN(new_n735));
  OAI21_X1  g0535(.A(new_n734), .B1(new_n677), .B2(new_n735), .ZN(new_n736));
  NAND2_X1  g0536(.A1(new_n733), .A2(new_n736), .ZN(new_n737));
  INV_X1    g0537(.A(new_n737), .ZN(new_n738));
  NAND3_X1  g0538(.A1(new_n218), .A2(G355), .A3(new_n291), .ZN(new_n739));
  OAI21_X1  g0539(.A(new_n739), .B1(G116), .B2(new_n218), .ZN(new_n740));
  OR2_X1    g0540(.A1(new_n240), .A2(new_n276), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n218), .A2(new_n287), .ZN(new_n742));
  AOI21_X1  g0542(.A(new_n742), .B1(new_n276), .B2(new_n226), .ZN(new_n743));
  AOI21_X1  g0543(.A(new_n740), .B1(new_n741), .B2(new_n743), .ZN(new_n744));
  NOR2_X1   g0544(.A1(G13), .A2(G33), .ZN(new_n745));
  INV_X1    g0545(.A(new_n745), .ZN(new_n746));
  NOR2_X1   g0546(.A1(new_n746), .A2(G20), .ZN(new_n747));
  AOI21_X1  g0547(.A(new_n221), .B1(G20), .B2(new_n534), .ZN(new_n748));
  NOR2_X1   g0548(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  INV_X1    g0549(.A(new_n749), .ZN(new_n750));
  OAI21_X1  g0550(.A(new_n738), .B1(new_n744), .B2(new_n750), .ZN(new_n751));
  INV_X1    g0551(.A(KEYINPUT99), .ZN(new_n752));
  AND2_X1   g0552(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  NOR2_X1   g0553(.A1(new_n222), .A2(new_n439), .ZN(new_n754));
  NOR2_X1   g0554(.A1(new_n296), .A2(G200), .ZN(new_n755));
  NAND2_X1  g0555(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  INV_X1    g0556(.A(KEYINPUT100), .ZN(new_n757));
  NAND2_X1  g0557(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  INV_X1    g0558(.A(new_n758), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n756), .A2(new_n757), .ZN(new_n760));
  NOR2_X1   g0560(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  NOR2_X1   g0561(.A1(new_n761), .A2(new_n349), .ZN(new_n762));
  NOR2_X1   g0562(.A1(new_n326), .A2(G179), .ZN(new_n763));
  NOR2_X1   g0563(.A1(new_n222), .A2(G190), .ZN(new_n764));
  NAND2_X1  g0564(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  NAND2_X1  g0565(.A1(new_n754), .A2(new_n763), .ZN(new_n766));
  OAI221_X1 g0566(.A(new_n291), .B1(new_n765), .B2(new_n302), .C1(new_n593), .C2(new_n766), .ZN(new_n767));
  NOR2_X1   g0567(.A1(new_n762), .A2(new_n767), .ZN(new_n768));
  NOR2_X1   g0568(.A1(G179), .A2(G200), .ZN(new_n769));
  NAND2_X1  g0569(.A1(new_n764), .A2(new_n769), .ZN(new_n770));
  NOR3_X1   g0570(.A1(new_n770), .A2(KEYINPUT32), .A3(new_n353), .ZN(new_n771));
  OAI21_X1  g0571(.A(KEYINPUT32), .B1(new_n770), .B2(new_n353), .ZN(new_n772));
  NAND2_X1  g0572(.A1(new_n769), .A2(G190), .ZN(new_n773));
  NAND2_X1  g0573(.A1(new_n773), .A2(G20), .ZN(new_n774));
  NAND2_X1  g0574(.A1(new_n774), .A2(G97), .ZN(new_n775));
  NAND2_X1  g0575(.A1(new_n772), .A2(new_n775), .ZN(new_n776));
  NAND3_X1  g0576(.A1(G20), .A2(G179), .A3(G200), .ZN(new_n777));
  XNOR2_X1  g0577(.A(new_n777), .B(KEYINPUT102), .ZN(new_n778));
  NOR2_X1   g0578(.A1(new_n778), .A2(G190), .ZN(new_n779));
  AOI211_X1 g0579(.A(new_n771), .B(new_n776), .C1(G68), .C2(new_n779), .ZN(new_n780));
  NAND2_X1  g0580(.A1(new_n755), .A2(new_n764), .ZN(new_n781));
  INV_X1    g0581(.A(KEYINPUT101), .ZN(new_n782));
  NAND2_X1  g0582(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  INV_X1    g0583(.A(new_n783), .ZN(new_n784));
  NOR2_X1   g0584(.A1(new_n781), .A2(new_n782), .ZN(new_n785));
  NOR2_X1   g0585(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  INV_X1    g0586(.A(new_n786), .ZN(new_n787));
  NAND2_X1  g0587(.A1(new_n787), .A2(G77), .ZN(new_n788));
  NOR2_X1   g0588(.A1(new_n778), .A2(new_n439), .ZN(new_n789));
  NAND2_X1  g0589(.A1(new_n789), .A2(G50), .ZN(new_n790));
  NAND4_X1  g0590(.A1(new_n768), .A2(new_n780), .A3(new_n788), .A4(new_n790), .ZN(new_n791));
  OR2_X1    g0591(.A1(new_n770), .A2(KEYINPUT104), .ZN(new_n792));
  NAND2_X1  g0592(.A1(new_n770), .A2(KEYINPUT104), .ZN(new_n793));
  NAND2_X1  g0593(.A1(new_n792), .A2(new_n793), .ZN(new_n794));
  INV_X1    g0594(.A(new_n794), .ZN(new_n795));
  AOI22_X1  g0595(.A1(new_n787), .A2(G311), .B1(new_n795), .B2(G329), .ZN(new_n796));
  INV_X1    g0596(.A(G283), .ZN(new_n797));
  OAI221_X1 g0597(.A(new_n287), .B1(new_n765), .B2(new_n797), .C1(new_n461), .C2(new_n766), .ZN(new_n798));
  INV_X1    g0598(.A(new_n761), .ZN(new_n799));
  AOI21_X1  g0599(.A(new_n798), .B1(new_n799), .B2(G322), .ZN(new_n800));
  AOI22_X1  g0600(.A1(new_n789), .A2(G326), .B1(G294), .B2(new_n774), .ZN(new_n801));
  INV_X1    g0601(.A(KEYINPUT103), .ZN(new_n802));
  NAND2_X1  g0602(.A1(new_n801), .A2(new_n802), .ZN(new_n803));
  XNOR2_X1  g0603(.A(KEYINPUT33), .B(G317), .ZN(new_n804));
  NAND2_X1  g0604(.A1(new_n779), .A2(new_n804), .ZN(new_n805));
  NAND4_X1  g0605(.A1(new_n796), .A2(new_n800), .A3(new_n803), .A4(new_n805), .ZN(new_n806));
  NOR2_X1   g0606(.A1(new_n801), .A2(new_n802), .ZN(new_n807));
  OAI21_X1  g0607(.A(new_n791), .B1(new_n806), .B2(new_n807), .ZN(new_n808));
  AOI21_X1  g0608(.A(new_n753), .B1(new_n748), .B2(new_n808), .ZN(new_n809));
  INV_X1    g0609(.A(new_n747), .ZN(new_n810));
  OAI221_X1 g0610(.A(new_n809), .B1(new_n752), .B2(new_n751), .C1(new_n666), .C2(new_n810), .ZN(new_n811));
  NAND2_X1  g0611(.A1(new_n666), .A2(G330), .ZN(new_n812));
  NAND2_X1  g0612(.A1(new_n812), .A2(new_n737), .ZN(new_n813));
  NOR2_X1   g0613(.A1(new_n666), .A2(G330), .ZN(new_n814));
  OAI21_X1  g0614(.A(new_n811), .B1(new_n813), .B2(new_n814), .ZN(new_n815));
  XNOR2_X1  g0615(.A(new_n815), .B(KEYINPUT105), .ZN(new_n816));
  INV_X1    g0616(.A(new_n816), .ZN(G396));
  NOR2_X1   g0617(.A1(new_n748), .A2(new_n745), .ZN(new_n818));
  AOI21_X1  g0618(.A(new_n737), .B1(new_n290), .B2(new_n818), .ZN(new_n819));
  INV_X1    g0619(.A(new_n748), .ZN(new_n820));
  OAI22_X1  g0620(.A1(new_n761), .A2(new_n557), .B1(new_n786), .B2(new_n489), .ZN(new_n821));
  INV_X1    g0621(.A(new_n765), .ZN(new_n822));
  AOI21_X1  g0622(.A(new_n291), .B1(new_n822), .B2(G87), .ZN(new_n823));
  OAI211_X1 g0623(.A(new_n823), .B(new_n775), .C1(new_n302), .C2(new_n766), .ZN(new_n824));
  AOI21_X1  g0624(.A(new_n824), .B1(G283), .B2(new_n779), .ZN(new_n825));
  INV_X1    g0625(.A(new_n789), .ZN(new_n826));
  OAI21_X1  g0626(.A(new_n825), .B1(new_n461), .B2(new_n826), .ZN(new_n827));
  AOI211_X1 g0627(.A(new_n821), .B(new_n827), .C1(G311), .C2(new_n795), .ZN(new_n828));
  INV_X1    g0628(.A(G132), .ZN(new_n829));
  NOR2_X1   g0629(.A1(new_n794), .A2(new_n829), .ZN(new_n830));
  AOI21_X1  g0630(.A(new_n287), .B1(new_n822), .B2(G68), .ZN(new_n831));
  INV_X1    g0631(.A(new_n774), .ZN(new_n832));
  OAI221_X1 g0632(.A(new_n831), .B1(new_n202), .B2(new_n766), .C1(new_n349), .C2(new_n832), .ZN(new_n833));
  AOI22_X1  g0633(.A1(G143), .A2(new_n799), .B1(new_n787), .B2(G159), .ZN(new_n834));
  AOI22_X1  g0634(.A1(G137), .A2(new_n789), .B1(new_n779), .B2(G150), .ZN(new_n835));
  INV_X1    g0635(.A(KEYINPUT106), .ZN(new_n836));
  AND2_X1   g0636(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  NOR2_X1   g0637(.A1(new_n835), .A2(new_n836), .ZN(new_n838));
  OAI21_X1  g0638(.A(new_n834), .B1(new_n837), .B2(new_n838), .ZN(new_n839));
  INV_X1    g0639(.A(KEYINPUT34), .ZN(new_n840));
  AOI211_X1 g0640(.A(new_n830), .B(new_n833), .C1(new_n839), .C2(new_n840), .ZN(new_n841));
  OR2_X1    g0641(.A1(new_n839), .A2(new_n840), .ZN(new_n842));
  AOI21_X1  g0642(.A(new_n828), .B1(new_n841), .B2(new_n842), .ZN(new_n843));
  NAND2_X1  g0643(.A1(new_n322), .A2(new_n663), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n327), .A2(new_n844), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n845), .A2(new_n324), .ZN(new_n846));
  OR3_X1    g0646(.A1(new_n310), .A2(new_n323), .A3(new_n663), .ZN(new_n847));
  NAND2_X1  g0647(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  INV_X1    g0648(.A(new_n848), .ZN(new_n849));
  OAI221_X1 g0649(.A(new_n819), .B1(new_n820), .B2(new_n843), .C1(new_n849), .C2(new_n746), .ZN(new_n850));
  INV_X1    g0650(.A(new_n715), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n644), .A2(new_n664), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n852), .A2(new_n848), .ZN(new_n853));
  NAND3_X1  g0653(.A1(new_n644), .A2(new_n664), .A3(new_n849), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  AOI21_X1  g0655(.A(new_n738), .B1(new_n851), .B2(new_n855), .ZN(new_n856));
  INV_X1    g0656(.A(new_n856), .ZN(new_n857));
  NOR2_X1   g0657(.A1(new_n851), .A2(new_n855), .ZN(new_n858));
  OAI21_X1  g0658(.A(new_n850), .B1(new_n857), .B2(new_n858), .ZN(G384));
  NOR2_X1   g0659(.A1(new_n731), .A2(new_n259), .ZN(new_n860));
  INV_X1    g0660(.A(KEYINPUT38), .ZN(new_n861));
  NAND4_X1  g0661(.A1(new_n376), .A2(new_n377), .A3(new_n352), .A4(new_n355), .ZN(new_n862));
  AOI21_X1  g0662(.A(new_n265), .B1(new_n862), .B2(new_n348), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n386), .A2(new_n863), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n864), .A2(new_n346), .ZN(new_n865));
  INV_X1    g0665(.A(new_n661), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  AOI21_X1  g0667(.A(new_n867), .B1(new_n404), .B2(new_n412), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n401), .A2(new_n402), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n401), .A2(new_n866), .ZN(new_n870));
  INV_X1    g0670(.A(KEYINPUT37), .ZN(new_n871));
  NAND4_X1  g0671(.A1(new_n869), .A2(new_n870), .A3(new_n871), .A4(new_n407), .ZN(new_n872));
  OAI21_X1  g0672(.A(new_n865), .B1(new_n402), .B2(new_n866), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n407), .A2(new_n873), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n874), .A2(KEYINPUT37), .ZN(new_n875));
  AND2_X1   g0675(.A1(new_n872), .A2(new_n875), .ZN(new_n876));
  OAI21_X1  g0676(.A(new_n861), .B1(new_n868), .B2(new_n876), .ZN(new_n877));
  AOI21_X1  g0677(.A(new_n861), .B1(new_n872), .B2(new_n875), .ZN(new_n878));
  INV_X1    g0678(.A(new_n867), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n455), .A2(new_n879), .ZN(new_n880));
  AND3_X1   g0680(.A1(new_n878), .A2(new_n880), .A3(KEYINPUT108), .ZN(new_n881));
  AOI21_X1  g0681(.A(KEYINPUT108), .B1(new_n878), .B2(new_n880), .ZN(new_n882));
  OAI21_X1  g0682(.A(new_n877), .B1(new_n881), .B2(new_n882), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n883), .A2(KEYINPUT109), .ZN(new_n884));
  INV_X1    g0684(.A(KEYINPUT109), .ZN(new_n885));
  OAI211_X1 g0685(.A(new_n885), .B(new_n877), .C1(new_n881), .C2(new_n882), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n884), .A2(new_n886), .ZN(new_n887));
  INV_X1    g0687(.A(new_n449), .ZN(new_n888));
  INV_X1    g0688(.A(KEYINPUT107), .ZN(new_n889));
  NAND3_X1  g0689(.A1(new_n888), .A2(new_n889), .A3(new_n437), .ZN(new_n890));
  OAI21_X1  g0690(.A(KEYINPUT107), .B1(new_n449), .B2(new_n450), .ZN(new_n891));
  NOR2_X1   g0691(.A1(new_n450), .A2(new_n664), .ZN(new_n892));
  NOR2_X1   g0692(.A1(new_n651), .A2(new_n892), .ZN(new_n893));
  NAND3_X1  g0693(.A1(new_n890), .A2(new_n891), .A3(new_n893), .ZN(new_n894));
  OAI21_X1  g0694(.A(new_n892), .B1(new_n888), .B2(new_n651), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  NAND4_X1  g0696(.A1(new_n501), .A2(new_n611), .A3(new_n507), .A4(new_n664), .ZN(new_n897));
  NAND3_X1  g0697(.A1(new_n897), .A2(new_n705), .A3(new_n710), .ZN(new_n898));
  NAND3_X1  g0698(.A1(new_n896), .A2(new_n849), .A3(new_n898), .ZN(new_n899));
  INV_X1    g0699(.A(new_n899), .ZN(new_n900));
  AOI21_X1  g0700(.A(KEYINPUT40), .B1(new_n887), .B2(new_n900), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n878), .A2(new_n880), .ZN(new_n902));
  OAI21_X1  g0702(.A(new_n412), .B1(new_n647), .B2(new_n648), .ZN(new_n903));
  INV_X1    g0703(.A(new_n870), .ZN(new_n904));
  NAND3_X1  g0704(.A1(new_n869), .A2(new_n870), .A3(new_n407), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n905), .A2(KEYINPUT37), .ZN(new_n906));
  AOI22_X1  g0706(.A1(new_n903), .A2(new_n904), .B1(new_n872), .B2(new_n906), .ZN(new_n907));
  OAI21_X1  g0707(.A(new_n902), .B1(new_n907), .B2(KEYINPUT38), .ZN(new_n908));
  INV_X1    g0708(.A(KEYINPUT40), .ZN(new_n909));
  NOR2_X1   g0709(.A1(new_n899), .A2(new_n909), .ZN(new_n910));
  AOI21_X1  g0710(.A(new_n901), .B1(new_n908), .B2(new_n910), .ZN(new_n911));
  AND2_X1   g0711(.A1(new_n458), .A2(new_n898), .ZN(new_n912));
  AOI21_X1  g0712(.A(new_n680), .B1(new_n911), .B2(new_n912), .ZN(new_n913));
  OAI21_X1  g0713(.A(new_n913), .B1(new_n911), .B2(new_n912), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n890), .A2(new_n891), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n915), .A2(new_n664), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n883), .A2(KEYINPUT39), .ZN(new_n917));
  INV_X1    g0717(.A(KEYINPUT39), .ZN(new_n918));
  OAI211_X1 g0718(.A(new_n918), .B(new_n902), .C1(new_n907), .C2(KEYINPUT38), .ZN(new_n919));
  AOI21_X1  g0719(.A(new_n916), .B1(new_n917), .B2(new_n919), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n854), .A2(new_n847), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n921), .A2(new_n896), .ZN(new_n922));
  AOI21_X1  g0722(.A(new_n922), .B1(new_n884), .B2(new_n886), .ZN(new_n923));
  NOR2_X1   g0723(.A1(new_n650), .A2(new_n866), .ZN(new_n924));
  NOR3_X1   g0724(.A1(new_n920), .A2(new_n923), .A3(new_n924), .ZN(new_n925));
  NAND4_X1  g0725(.A1(new_n724), .A2(new_n456), .A3(new_n413), .A4(new_n343), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n926), .A2(new_n655), .ZN(new_n927));
  XOR2_X1   g0727(.A(new_n925), .B(new_n927), .Z(new_n928));
  AOI21_X1  g0728(.A(new_n860), .B1(new_n914), .B2(new_n928), .ZN(new_n929));
  OAI21_X1  g0729(.A(new_n929), .B1(new_n928), .B2(new_n914), .ZN(new_n930));
  INV_X1    g0730(.A(KEYINPUT35), .ZN(new_n931));
  OAI211_X1 g0731(.A(G116), .B(new_n223), .C1(new_n514), .C2(new_n931), .ZN(new_n932));
  AOI21_X1  g0732(.A(new_n932), .B1(new_n931), .B2(new_n514), .ZN(new_n933));
  XOR2_X1   g0733(.A(new_n933), .B(KEYINPUT36), .Z(new_n934));
  OAI211_X1 g0734(.A(new_n226), .B(G77), .C1(new_n350), .C2(new_n349), .ZN(new_n935));
  OAI21_X1  g0735(.A(new_n935), .B1(G50), .B2(new_n350), .ZN(new_n936));
  NAND3_X1  g0736(.A1(new_n936), .A2(G1), .A3(new_n730), .ZN(new_n937));
  NAND3_X1  g0737(.A1(new_n930), .A2(new_n934), .A3(new_n937), .ZN(G367));
  OAI221_X1 g0738(.A(new_n749), .B1(new_n218), .B2(new_n315), .C1(new_n742), .C2(new_n234), .ZN(new_n939));
  AND2_X1   g0739(.A1(new_n738), .A2(new_n939), .ZN(new_n940));
  AOI21_X1  g0740(.A(new_n664), .B1(new_n608), .B2(new_n601), .ZN(new_n941));
  OR2_X1    g0741(.A1(new_n627), .A2(new_n941), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n640), .A2(new_n941), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  INV_X1    g0744(.A(new_n766), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n945), .A2(G116), .ZN(new_n946));
  XOR2_X1   g0746(.A(new_n946), .B(KEYINPUT46), .Z(new_n947));
  AOI21_X1  g0747(.A(new_n947), .B1(G107), .B2(new_n774), .ZN(new_n948));
  INV_X1    g0748(.A(new_n779), .ZN(new_n949));
  INV_X1    g0749(.A(G311), .ZN(new_n950));
  OAI221_X1 g0750(.A(new_n948), .B1(new_n557), .B2(new_n949), .C1(new_n950), .C2(new_n826), .ZN(new_n951));
  NOR2_X1   g0751(.A1(new_n765), .A2(new_n479), .ZN(new_n952));
  INV_X1    g0752(.A(new_n770), .ZN(new_n953));
  AOI211_X1 g0753(.A(new_n291), .B(new_n952), .C1(G317), .C2(new_n953), .ZN(new_n954));
  OAI221_X1 g0754(.A(new_n954), .B1(new_n797), .B2(new_n786), .C1(new_n461), .C2(new_n761), .ZN(new_n955));
  OAI21_X1  g0755(.A(new_n291), .B1(new_n766), .B2(new_n349), .ZN(new_n956));
  INV_X1    g0756(.A(G137), .ZN(new_n957));
  OAI22_X1  g0757(.A1(new_n765), .A2(new_n290), .B1(new_n770), .B2(new_n957), .ZN(new_n958));
  AOI211_X1 g0758(.A(new_n956), .B(new_n958), .C1(G68), .C2(new_n774), .ZN(new_n959));
  INV_X1    g0759(.A(G150), .ZN(new_n960));
  OAI221_X1 g0760(.A(new_n959), .B1(new_n202), .B2(new_n786), .C1(new_n960), .C2(new_n761), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n789), .A2(G143), .ZN(new_n962));
  OAI21_X1  g0762(.A(new_n962), .B1(new_n949), .B2(new_n353), .ZN(new_n963));
  OAI22_X1  g0763(.A1(new_n951), .A2(new_n955), .B1(new_n961), .B2(new_n963), .ZN(new_n964));
  XOR2_X1   g0764(.A(new_n964), .B(KEYINPUT47), .Z(new_n965));
  OAI221_X1 g0765(.A(new_n940), .B1(new_n944), .B2(new_n810), .C1(new_n965), .C2(new_n820), .ZN(new_n966));
  NAND3_X1  g0766(.A1(new_n638), .A2(new_n632), .A3(new_n663), .ZN(new_n967));
  OAI211_X1 g0767(.A(new_n536), .B(new_n568), .C1(new_n633), .C2(new_n664), .ZN(new_n968));
  AND2_X1   g0768(.A1(new_n967), .A2(new_n968), .ZN(new_n969));
  OR2_X1    g0769(.A1(new_n969), .A2(new_n572), .ZN(new_n970));
  AND2_X1   g0770(.A1(new_n970), .A2(new_n536), .ZN(new_n971));
  INV_X1    g0771(.A(KEYINPUT110), .ZN(new_n972));
  AOI21_X1  g0772(.A(new_n663), .B1(new_n971), .B2(new_n972), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n970), .A2(new_n536), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n974), .A2(KEYINPUT110), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n672), .A2(new_n670), .ZN(new_n976));
  OAI21_X1  g0776(.A(KEYINPUT111), .B1(new_n976), .B2(new_n969), .ZN(new_n977));
  INV_X1    g0777(.A(new_n969), .ZN(new_n978));
  INV_X1    g0778(.A(KEYINPUT111), .ZN(new_n979));
  NAND4_X1  g0779(.A1(new_n672), .A2(new_n978), .A3(new_n979), .A4(new_n670), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n977), .A2(new_n980), .ZN(new_n981));
  AOI22_X1  g0781(.A1(new_n973), .A2(new_n975), .B1(KEYINPUT42), .B2(new_n981), .ZN(new_n982));
  OR2_X1    g0782(.A1(new_n981), .A2(KEYINPUT42), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n982), .A2(new_n983), .ZN(new_n984));
  INV_X1    g0784(.A(new_n944), .ZN(new_n985));
  INV_X1    g0785(.A(KEYINPUT43), .ZN(new_n986));
  NAND2_X1  g0786(.A1(new_n985), .A2(new_n986), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n944), .A2(KEYINPUT43), .ZN(new_n988));
  NAND3_X1  g0788(.A1(new_n984), .A2(new_n987), .A3(new_n988), .ZN(new_n989));
  NAND4_X1  g0789(.A1(new_n982), .A2(new_n986), .A3(new_n985), .A4(new_n983), .ZN(new_n990));
  NAND2_X1  g0790(.A1(new_n989), .A2(new_n990), .ZN(new_n991));
  NOR2_X1   g0791(.A1(new_n671), .A2(new_n969), .ZN(new_n992));
  INV_X1    g0792(.A(new_n992), .ZN(new_n993));
  XNOR2_X1  g0793(.A(new_n991), .B(new_n993), .ZN(new_n994));
  INV_X1    g0794(.A(KEYINPUT45), .ZN(new_n995));
  INV_X1    g0795(.A(new_n667), .ZN(new_n996));
  NAND2_X1  g0796(.A1(new_n976), .A2(new_n996), .ZN(new_n997));
  OAI21_X1  g0797(.A(new_n995), .B1(new_n997), .B2(new_n969), .ZN(new_n998));
  NAND3_X1  g0798(.A1(new_n673), .A2(KEYINPUT45), .A3(new_n978), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n998), .A2(new_n999), .ZN(new_n1000));
  XOR2_X1   g0800(.A(KEYINPUT112), .B(KEYINPUT44), .Z(new_n1001));
  NAND3_X1  g0801(.A1(new_n997), .A2(new_n969), .A3(new_n1001), .ZN(new_n1002));
  INV_X1    g0802(.A(new_n1001), .ZN(new_n1003));
  OAI21_X1  g0803(.A(new_n1003), .B1(new_n673), .B2(new_n978), .ZN(new_n1004));
  NAND4_X1  g0804(.A1(new_n1000), .A2(new_n671), .A3(new_n1002), .A4(new_n1004), .ZN(new_n1005));
  NAND2_X1  g0805(.A1(new_n1005), .A2(KEYINPUT113), .ZN(new_n1006));
  NAND3_X1  g0806(.A1(new_n1000), .A2(new_n1002), .A3(new_n1004), .ZN(new_n1007));
  INV_X1    g0807(.A(new_n671), .ZN(new_n1008));
  NAND2_X1  g0808(.A1(new_n1007), .A2(new_n1008), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n1006), .A2(new_n1009), .ZN(new_n1010));
  NAND3_X1  g0810(.A1(new_n1007), .A2(KEYINPUT113), .A3(new_n1008), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n1010), .A2(new_n1011), .ZN(new_n1012));
  XOR2_X1   g0812(.A(new_n672), .B(new_n670), .Z(new_n1013));
  AOI21_X1  g0813(.A(KEYINPUT114), .B1(new_n666), .B2(G330), .ZN(new_n1014));
  NAND3_X1  g0814(.A1(new_n666), .A2(KEYINPUT114), .A3(G330), .ZN(new_n1015));
  INV_X1    g0815(.A(new_n1015), .ZN(new_n1016));
  OAI21_X1  g0816(.A(new_n1013), .B1(new_n1014), .B2(new_n1016), .ZN(new_n1017));
  OAI21_X1  g0817(.A(new_n1017), .B1(new_n1013), .B2(new_n1016), .ZN(new_n1018));
  OAI21_X1  g0818(.A(new_n727), .B1(new_n1012), .B2(new_n1018), .ZN(new_n1019));
  XOR2_X1   g0819(.A(new_n677), .B(KEYINPUT41), .Z(new_n1020));
  INV_X1    g0820(.A(new_n1020), .ZN(new_n1021));
  AOI21_X1  g0821(.A(new_n735), .B1(new_n1019), .B2(new_n1021), .ZN(new_n1022));
  OAI21_X1  g0822(.A(new_n966), .B1(new_n994), .B2(new_n1022), .ZN(G387));
  NOR2_X1   g0823(.A1(new_n726), .A2(new_n1018), .ZN(new_n1024));
  INV_X1    g0824(.A(new_n1024), .ZN(new_n1025));
  NAND2_X1  g0825(.A1(new_n726), .A2(new_n1018), .ZN(new_n1026));
  NAND3_X1  g0826(.A1(new_n1025), .A2(new_n1026), .A3(new_n677), .ZN(new_n1027));
  OR2_X1    g0827(.A1(new_n1018), .A2(new_n732), .ZN(new_n1028));
  AOI22_X1  g0828(.A1(G317), .A2(new_n799), .B1(new_n787), .B2(G303), .ZN(new_n1029));
  XOR2_X1   g0829(.A(KEYINPUT115), .B(G322), .Z(new_n1030));
  OAI221_X1 g0830(.A(new_n1029), .B1(new_n950), .B2(new_n949), .C1(new_n826), .C2(new_n1030), .ZN(new_n1031));
  INV_X1    g0831(.A(KEYINPUT48), .ZN(new_n1032));
  OR2_X1    g0832(.A1(new_n1031), .A2(new_n1032), .ZN(new_n1033));
  NAND2_X1  g0833(.A1(new_n1031), .A2(new_n1032), .ZN(new_n1034));
  AOI22_X1  g0834(.A1(new_n945), .A2(G294), .B1(new_n774), .B2(G283), .ZN(new_n1035));
  NAND3_X1  g0835(.A1(new_n1033), .A2(new_n1034), .A3(new_n1035), .ZN(new_n1036));
  XOR2_X1   g0836(.A(new_n1036), .B(KEYINPUT49), .Z(new_n1037));
  AOI21_X1  g0837(.A(new_n291), .B1(new_n953), .B2(G326), .ZN(new_n1038));
  OAI21_X1  g0838(.A(new_n1038), .B1(new_n489), .B2(new_n765), .ZN(new_n1039));
  NOR2_X1   g0839(.A1(new_n1037), .A2(new_n1039), .ZN(new_n1040));
  OAI22_X1  g0840(.A1(new_n761), .A2(new_n202), .B1(new_n786), .B2(new_n350), .ZN(new_n1041));
  OAI22_X1  g0841(.A1(new_n353), .A2(new_n826), .B1(new_n949), .B2(new_n344), .ZN(new_n1042));
  NOR2_X1   g0842(.A1(new_n766), .A2(new_n290), .ZN(new_n1043));
  AOI21_X1  g0843(.A(new_n1043), .B1(G150), .B2(new_n953), .ZN(new_n1044));
  NAND2_X1  g0844(.A1(new_n774), .A2(new_n314), .ZN(new_n1045));
  NOR2_X1   g0845(.A1(new_n952), .A2(new_n287), .ZN(new_n1046));
  NAND3_X1  g0846(.A1(new_n1044), .A2(new_n1045), .A3(new_n1046), .ZN(new_n1047));
  NOR3_X1   g0847(.A1(new_n1041), .A2(new_n1042), .A3(new_n1047), .ZN(new_n1048));
  OAI21_X1  g0848(.A(new_n748), .B1(new_n1040), .B2(new_n1048), .ZN(new_n1049));
  NOR3_X1   g0849(.A1(new_n231), .A2(new_n276), .A3(new_n291), .ZN(new_n1050));
  OR3_X1    g0850(.A1(new_n318), .A2(KEYINPUT50), .A3(G50), .ZN(new_n1051));
  OAI21_X1  g0851(.A(KEYINPUT50), .B1(new_n318), .B2(G50), .ZN(new_n1052));
  AOI21_X1  g0852(.A(G45), .B1(G68), .B2(G77), .ZN(new_n1053));
  NAND3_X1  g0853(.A1(new_n1051), .A2(new_n1052), .A3(new_n1053), .ZN(new_n1054));
  AOI211_X1 g0854(.A(G116), .B(new_n594), .C1(new_n1054), .C2(new_n287), .ZN(new_n1055));
  OAI21_X1  g0855(.A(new_n218), .B1(new_n1050), .B2(new_n1055), .ZN(new_n1056));
  AOI21_X1  g0856(.A(new_n750), .B1(new_n676), .B2(G107), .ZN(new_n1057));
  AOI21_X1  g0857(.A(new_n737), .B1(new_n1056), .B2(new_n1057), .ZN(new_n1058));
  OAI211_X1 g0858(.A(new_n1049), .B(new_n1058), .C1(new_n670), .C2(new_n810), .ZN(new_n1059));
  AND2_X1   g0859(.A1(new_n1028), .A2(new_n1059), .ZN(new_n1060));
  NAND2_X1  g0860(.A1(new_n1027), .A2(new_n1060), .ZN(G393));
  OAI221_X1 g0861(.A(new_n749), .B1(new_n479), .B2(new_n218), .C1(new_n742), .C2(new_n243), .ZN(new_n1062));
  NAND2_X1  g0862(.A1(new_n738), .A2(new_n1062), .ZN(new_n1063));
  NOR2_X1   g0863(.A1(new_n786), .A2(new_n557), .ZN(new_n1064));
  AOI21_X1  g0864(.A(new_n291), .B1(new_n822), .B2(G107), .ZN(new_n1065));
  OAI221_X1 g0865(.A(new_n1065), .B1(new_n797), .B2(new_n766), .C1(new_n770), .C2(new_n1030), .ZN(new_n1066));
  AOI211_X1 g0866(.A(new_n1064), .B(new_n1066), .C1(G116), .C2(new_n774), .ZN(new_n1067));
  OAI21_X1  g0867(.A(new_n1067), .B1(new_n461), .B2(new_n949), .ZN(new_n1068));
  AOI22_X1  g0868(.A1(new_n799), .A2(G311), .B1(G317), .B2(new_n789), .ZN(new_n1069));
  XNOR2_X1  g0869(.A(new_n1069), .B(KEYINPUT52), .ZN(new_n1070));
  AOI22_X1  g0870(.A1(G68), .A2(new_n945), .B1(new_n953), .B2(G143), .ZN(new_n1071));
  OAI211_X1 g0871(.A(new_n1071), .B(new_n291), .C1(new_n210), .C2(new_n765), .ZN(new_n1072));
  AOI21_X1  g0872(.A(new_n1072), .B1(G77), .B2(new_n774), .ZN(new_n1073));
  OAI221_X1 g0873(.A(new_n1073), .B1(new_n202), .B2(new_n949), .C1(new_n318), .C2(new_n786), .ZN(new_n1074));
  OAI22_X1  g0874(.A1(new_n761), .A2(new_n353), .B1(new_n826), .B2(new_n960), .ZN(new_n1075));
  XOR2_X1   g0875(.A(new_n1075), .B(KEYINPUT51), .Z(new_n1076));
  OAI22_X1  g0876(.A1(new_n1068), .A2(new_n1070), .B1(new_n1074), .B2(new_n1076), .ZN(new_n1077));
  AOI21_X1  g0877(.A(new_n1063), .B1(new_n1077), .B2(new_n748), .ZN(new_n1078));
  OAI21_X1  g0878(.A(new_n1078), .B1(new_n978), .B2(new_n810), .ZN(new_n1079));
  NAND2_X1  g0879(.A1(new_n1009), .A2(new_n1005), .ZN(new_n1080));
  OAI21_X1  g0880(.A(new_n1079), .B1(new_n1080), .B2(new_n732), .ZN(new_n1081));
  NAND2_X1  g0881(.A1(new_n1025), .A2(new_n1080), .ZN(new_n1082));
  INV_X1    g0882(.A(new_n1012), .ZN(new_n1083));
  AOI21_X1  g0883(.A(new_n729), .B1(new_n1024), .B2(new_n1083), .ZN(new_n1084));
  AOI21_X1  g0884(.A(new_n1081), .B1(new_n1082), .B2(new_n1084), .ZN(new_n1085));
  INV_X1    g0885(.A(new_n1085), .ZN(G390));
  NAND2_X1  g0886(.A1(new_n922), .A2(new_n916), .ZN(new_n1087));
  NAND3_X1  g0887(.A1(new_n917), .A2(new_n1087), .A3(new_n919), .ZN(new_n1088));
  NAND2_X1  g0888(.A1(new_n723), .A2(new_n846), .ZN(new_n1089));
  NAND2_X1  g0889(.A1(new_n1089), .A2(new_n847), .ZN(new_n1090));
  NAND2_X1  g0890(.A1(new_n1090), .A2(new_n896), .ZN(new_n1091));
  NAND3_X1  g0891(.A1(new_n1091), .A2(new_n908), .A3(new_n916), .ZN(new_n1092));
  NAND2_X1  g0892(.A1(new_n1088), .A2(new_n1092), .ZN(new_n1093));
  AND2_X1   g0893(.A1(new_n898), .A2(G330), .ZN(new_n1094));
  NAND3_X1  g0894(.A1(new_n1094), .A2(new_n896), .A3(new_n849), .ZN(new_n1095));
  INV_X1    g0895(.A(new_n1095), .ZN(new_n1096));
  NAND2_X1  g0896(.A1(new_n1093), .A2(new_n1096), .ZN(new_n1097));
  NAND3_X1  g0897(.A1(new_n715), .A2(new_n849), .A3(new_n896), .ZN(new_n1098));
  NAND3_X1  g0898(.A1(new_n1088), .A2(new_n1092), .A3(new_n1098), .ZN(new_n1099));
  NAND3_X1  g0899(.A1(new_n1097), .A2(new_n1099), .A3(new_n735), .ZN(new_n1100));
  NAND3_X1  g0900(.A1(new_n917), .A2(new_n745), .A3(new_n919), .ZN(new_n1101));
  INV_X1    g0901(.A(new_n818), .ZN(new_n1102));
  OAI21_X1  g0902(.A(new_n738), .B1(new_n250), .B2(new_n1102), .ZN(new_n1103));
  OAI22_X1  g0903(.A1(new_n794), .A2(new_n557), .B1(new_n350), .B2(new_n765), .ZN(new_n1104));
  XOR2_X1   g0904(.A(new_n1104), .B(KEYINPUT119), .Z(new_n1105));
  OAI221_X1 g0905(.A(new_n287), .B1(new_n766), .B2(new_n210), .C1(new_n832), .C2(new_n290), .ZN(new_n1106));
  AOI21_X1  g0906(.A(new_n1106), .B1(new_n799), .B2(G116), .ZN(new_n1107));
  AOI22_X1  g0907(.A1(new_n787), .A2(G97), .B1(new_n779), .B2(G107), .ZN(new_n1108));
  INV_X1    g0908(.A(KEYINPUT118), .ZN(new_n1109));
  OAI221_X1 g0909(.A(new_n1107), .B1(new_n797), .B2(new_n826), .C1(new_n1108), .C2(new_n1109), .ZN(new_n1110));
  AOI211_X1 g0910(.A(new_n1105), .B(new_n1110), .C1(new_n1109), .C2(new_n1108), .ZN(new_n1111));
  XNOR2_X1  g0911(.A(KEYINPUT54), .B(G143), .ZN(new_n1112));
  INV_X1    g0912(.A(G125), .ZN(new_n1113));
  OAI22_X1  g0913(.A1(new_n786), .A2(new_n1112), .B1(new_n794), .B2(new_n1113), .ZN(new_n1114));
  NOR2_X1   g0914(.A1(new_n766), .A2(new_n960), .ZN(new_n1115));
  XNOR2_X1  g0915(.A(KEYINPUT116), .B(KEYINPUT53), .ZN(new_n1116));
  OAI22_X1  g0916(.A1(new_n1115), .A2(new_n1116), .B1(new_n832), .B2(new_n353), .ZN(new_n1117));
  NAND2_X1  g0917(.A1(new_n1115), .A2(new_n1116), .ZN(new_n1118));
  OAI211_X1 g0918(.A(new_n1118), .B(new_n291), .C1(new_n202), .C2(new_n765), .ZN(new_n1119));
  AOI211_X1 g0919(.A(new_n1117), .B(new_n1119), .C1(G137), .C2(new_n779), .ZN(new_n1120));
  INV_X1    g0920(.A(G128), .ZN(new_n1121));
  OAI21_X1  g0921(.A(new_n1120), .B1(new_n1121), .B2(new_n826), .ZN(new_n1122));
  AOI211_X1 g0922(.A(new_n1114), .B(new_n1122), .C1(G132), .C2(new_n799), .ZN(new_n1123));
  INV_X1    g0923(.A(new_n1123), .ZN(new_n1124));
  AOI21_X1  g0924(.A(new_n1111), .B1(new_n1124), .B2(KEYINPUT117), .ZN(new_n1125));
  OAI21_X1  g0925(.A(new_n1125), .B1(KEYINPUT117), .B2(new_n1124), .ZN(new_n1126));
  AOI21_X1  g0926(.A(new_n1103), .B1(new_n1126), .B2(new_n748), .ZN(new_n1127));
  NAND2_X1  g0927(.A1(new_n1101), .A2(new_n1127), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n1100), .A2(new_n1128), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n1097), .A2(new_n1099), .ZN(new_n1130));
  NAND2_X1  g0930(.A1(new_n898), .A2(G330), .ZN(new_n1131));
  OAI211_X1 g0931(.A(new_n926), .B(new_n655), .C1(new_n457), .C2(new_n1131), .ZN(new_n1132));
  AOI21_X1  g0932(.A(new_n896), .B1(new_n715), .B2(new_n849), .ZN(new_n1133));
  OAI21_X1  g0933(.A(new_n921), .B1(new_n1133), .B2(new_n1096), .ZN(new_n1134));
  AOI21_X1  g0934(.A(new_n896), .B1(new_n1094), .B2(new_n849), .ZN(new_n1135));
  NOR2_X1   g0935(.A1(new_n1135), .A2(new_n1090), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n1136), .A2(new_n1098), .ZN(new_n1137));
  AOI21_X1  g0937(.A(new_n1132), .B1(new_n1134), .B2(new_n1137), .ZN(new_n1138));
  INV_X1    g0938(.A(new_n1138), .ZN(new_n1139));
  AOI21_X1  g0939(.A(new_n729), .B1(new_n1130), .B2(new_n1139), .ZN(new_n1140));
  NAND3_X1  g0940(.A1(new_n1097), .A2(new_n1138), .A3(new_n1099), .ZN(new_n1141));
  AOI21_X1  g0941(.A(new_n1129), .B1(new_n1140), .B2(new_n1141), .ZN(new_n1142));
  INV_X1    g0942(.A(new_n1142), .ZN(G378));
  INV_X1    g0943(.A(new_n925), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n341), .A2(new_n299), .ZN(new_n1145));
  NAND2_X1  g0945(.A1(new_n271), .A2(new_n866), .ZN(new_n1146));
  XNOR2_X1  g0946(.A(new_n1146), .B(KEYINPUT55), .ZN(new_n1147));
  XNOR2_X1  g0947(.A(new_n1145), .B(new_n1147), .ZN(new_n1148));
  XOR2_X1   g0948(.A(KEYINPUT121), .B(KEYINPUT56), .Z(new_n1149));
  XNOR2_X1  g0949(.A(new_n1148), .B(new_n1149), .ZN(new_n1150));
  INV_X1    g0950(.A(KEYINPUT108), .ZN(new_n1151));
  NAND2_X1  g0951(.A1(new_n902), .A2(new_n1151), .ZN(new_n1152));
  NAND3_X1  g0952(.A1(new_n878), .A2(new_n880), .A3(KEYINPUT108), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n1152), .A2(new_n1153), .ZN(new_n1154));
  AOI21_X1  g0954(.A(new_n885), .B1(new_n1154), .B2(new_n877), .ZN(new_n1155));
  INV_X1    g0955(.A(new_n886), .ZN(new_n1156));
  OAI21_X1  g0956(.A(new_n900), .B1(new_n1155), .B2(new_n1156), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n1157), .A2(new_n909), .ZN(new_n1158));
  AOI21_X1  g0958(.A(new_n680), .B1(new_n910), .B2(new_n908), .ZN(new_n1159));
  AOI21_X1  g0959(.A(new_n1150), .B1(new_n1158), .B2(new_n1159), .ZN(new_n1160));
  AOI21_X1  g0960(.A(new_n899), .B1(new_n884), .B2(new_n886), .ZN(new_n1161));
  OAI211_X1 g0961(.A(new_n1150), .B(new_n1159), .C1(new_n1161), .C2(KEYINPUT40), .ZN(new_n1162));
  INV_X1    g0962(.A(new_n1162), .ZN(new_n1163));
  OAI21_X1  g0963(.A(new_n1144), .B1(new_n1160), .B2(new_n1163), .ZN(new_n1164));
  INV_X1    g0964(.A(new_n1150), .ZN(new_n1165));
  INV_X1    g0965(.A(new_n1159), .ZN(new_n1166));
  OAI21_X1  g0966(.A(new_n1165), .B1(new_n901), .B2(new_n1166), .ZN(new_n1167));
  NAND3_X1  g0967(.A1(new_n1167), .A2(new_n925), .A3(new_n1162), .ZN(new_n1168));
  NAND3_X1  g0968(.A1(new_n1164), .A2(new_n735), .A3(new_n1168), .ZN(new_n1169));
  NAND2_X1  g0969(.A1(new_n287), .A2(new_n273), .ZN(new_n1170));
  OAI211_X1 g0970(.A(new_n1170), .B(new_n202), .C1(G33), .C2(G41), .ZN(new_n1171));
  NOR2_X1   g0971(.A1(new_n765), .A2(new_n349), .ZN(new_n1172));
  NOR3_X1   g0972(.A1(new_n1043), .A2(new_n1172), .A3(new_n1170), .ZN(new_n1173));
  OAI221_X1 g0973(.A(new_n1173), .B1(new_n350), .B2(new_n832), .C1(new_n949), .C2(new_n479), .ZN(new_n1174));
  AOI22_X1  g0974(.A1(new_n799), .A2(G107), .B1(new_n795), .B2(G283), .ZN(new_n1175));
  OAI21_X1  g0975(.A(new_n1175), .B1(new_n315), .B2(new_n786), .ZN(new_n1176));
  AOI211_X1 g0976(.A(new_n1174), .B(new_n1176), .C1(G116), .C2(new_n789), .ZN(new_n1177));
  OAI21_X1  g0977(.A(new_n1171), .B1(new_n1177), .B2(KEYINPUT58), .ZN(new_n1178));
  XOR2_X1   g0978(.A(new_n1178), .B(KEYINPUT120), .Z(new_n1179));
  OAI22_X1  g0979(.A1(new_n832), .A2(new_n960), .B1(new_n1112), .B2(new_n766), .ZN(new_n1180));
  AOI21_X1  g0980(.A(new_n1180), .B1(new_n799), .B2(G128), .ZN(new_n1181));
  AOI22_X1  g0981(.A1(G125), .A2(new_n789), .B1(new_n779), .B2(G132), .ZN(new_n1182));
  OAI211_X1 g0982(.A(new_n1181), .B(new_n1182), .C1(new_n957), .C2(new_n786), .ZN(new_n1183));
  OR2_X1    g0983(.A1(new_n1183), .A2(KEYINPUT59), .ZN(new_n1184));
  AOI211_X1 g0984(.A(G33), .B(G41), .C1(new_n953), .C2(G124), .ZN(new_n1185));
  OAI21_X1  g0985(.A(new_n1185), .B1(new_n353), .B2(new_n765), .ZN(new_n1186));
  AOI21_X1  g0986(.A(new_n1186), .B1(new_n1183), .B2(KEYINPUT59), .ZN(new_n1187));
  AOI22_X1  g0987(.A1(new_n1177), .A2(KEYINPUT58), .B1(new_n1184), .B2(new_n1187), .ZN(new_n1188));
  AND2_X1   g0988(.A1(new_n1179), .A2(new_n1188), .ZN(new_n1189));
  OAI221_X1 g0989(.A(new_n738), .B1(G50), .B2(new_n1102), .C1(new_n1189), .C2(new_n820), .ZN(new_n1190));
  AOI21_X1  g0990(.A(new_n1190), .B1(new_n1150), .B2(new_n745), .ZN(new_n1191));
  XOR2_X1   g0991(.A(new_n1191), .B(KEYINPUT122), .Z(new_n1192));
  INV_X1    g0992(.A(new_n1192), .ZN(new_n1193));
  NAND2_X1  g0993(.A1(new_n1169), .A2(new_n1193), .ZN(new_n1194));
  INV_X1    g0994(.A(new_n1132), .ZN(new_n1195));
  NAND2_X1  g0995(.A1(new_n1141), .A2(new_n1195), .ZN(new_n1196));
  NAND3_X1  g0996(.A1(new_n1164), .A2(new_n1196), .A3(new_n1168), .ZN(new_n1197));
  INV_X1    g0997(.A(KEYINPUT57), .ZN(new_n1198));
  AOI21_X1  g0998(.A(new_n729), .B1(new_n1197), .B2(new_n1198), .ZN(new_n1199));
  NAND4_X1  g0999(.A1(new_n1164), .A2(new_n1196), .A3(KEYINPUT57), .A4(new_n1168), .ZN(new_n1200));
  AOI21_X1  g1000(.A(new_n1194), .B1(new_n1199), .B2(new_n1200), .ZN(new_n1201));
  INV_X1    g1001(.A(new_n1201), .ZN(G375));
  NAND3_X1  g1002(.A1(new_n1134), .A2(new_n1132), .A3(new_n1137), .ZN(new_n1203));
  NAND3_X1  g1003(.A1(new_n1139), .A2(new_n1021), .A3(new_n1203), .ZN(new_n1204));
  NAND3_X1  g1004(.A1(new_n894), .A2(new_n745), .A3(new_n895), .ZN(new_n1205));
  OAI21_X1  g1005(.A(new_n738), .B1(G68), .B2(new_n1102), .ZN(new_n1206));
  OAI21_X1  g1006(.A(new_n1045), .B1(new_n761), .B2(new_n797), .ZN(new_n1207));
  XOR2_X1   g1007(.A(new_n1207), .B(KEYINPUT123), .Z(new_n1208));
  NOR2_X1   g1008(.A1(new_n786), .A2(new_n302), .ZN(new_n1209));
  OAI221_X1 g1009(.A(new_n287), .B1(new_n765), .B2(new_n290), .C1(new_n479), .C2(new_n766), .ZN(new_n1210));
  NOR2_X1   g1010(.A1(new_n1209), .A2(new_n1210), .ZN(new_n1211));
  AOI22_X1  g1011(.A1(G116), .A2(new_n779), .B1(new_n789), .B2(G294), .ZN(new_n1212));
  OAI211_X1 g1012(.A(new_n1211), .B(new_n1212), .C1(new_n461), .C2(new_n794), .ZN(new_n1213));
  AOI22_X1  g1013(.A1(G137), .A2(new_n799), .B1(new_n787), .B2(G150), .ZN(new_n1214));
  OAI21_X1  g1014(.A(new_n1214), .B1(new_n1121), .B2(new_n794), .ZN(new_n1215));
  OAI221_X1 g1015(.A(new_n291), .B1(new_n765), .B2(new_n349), .C1(new_n353), .C2(new_n766), .ZN(new_n1216));
  AOI21_X1  g1016(.A(new_n1216), .B1(G50), .B2(new_n774), .ZN(new_n1217));
  OAI221_X1 g1017(.A(new_n1217), .B1(new_n829), .B2(new_n826), .C1(new_n949), .C2(new_n1112), .ZN(new_n1218));
  OAI22_X1  g1018(.A1(new_n1208), .A2(new_n1213), .B1(new_n1215), .B2(new_n1218), .ZN(new_n1219));
  AOI21_X1  g1019(.A(new_n1206), .B1(new_n1219), .B2(new_n748), .ZN(new_n1220));
  NAND2_X1  g1020(.A1(new_n1205), .A2(new_n1220), .ZN(new_n1221));
  AOI211_X1 g1021(.A(new_n680), .B(new_n848), .C1(new_n713), .C2(new_n714), .ZN(new_n1222));
  OAI21_X1  g1022(.A(new_n1095), .B1(new_n1222), .B2(new_n896), .ZN(new_n1223));
  AOI22_X1  g1023(.A1(new_n1223), .A2(new_n921), .B1(new_n1098), .B2(new_n1136), .ZN(new_n1224));
  OAI21_X1  g1024(.A(new_n1221), .B1(new_n1224), .B2(new_n732), .ZN(new_n1225));
  INV_X1    g1025(.A(new_n1225), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n1204), .A2(new_n1226), .ZN(G381));
  NOR2_X1   g1027(.A1(G393), .A2(G396), .ZN(new_n1228));
  INV_X1    g1028(.A(G384), .ZN(new_n1229));
  NAND3_X1  g1029(.A1(new_n1228), .A2(new_n1229), .A3(new_n1085), .ZN(new_n1230));
  NOR2_X1   g1030(.A1(new_n1230), .A2(G381), .ZN(new_n1231));
  NOR2_X1   g1031(.A1(G387), .A2(G378), .ZN(new_n1232));
  NAND3_X1  g1032(.A1(new_n1231), .A2(new_n1201), .A3(new_n1232), .ZN(G407));
  NAND2_X1  g1033(.A1(new_n662), .A2(G213), .ZN(new_n1234));
  INV_X1    g1034(.A(new_n1234), .ZN(new_n1235));
  NAND3_X1  g1035(.A1(new_n1201), .A2(new_n1142), .A3(new_n1235), .ZN(new_n1236));
  NAND3_X1  g1036(.A1(G407), .A2(G213), .A3(new_n1236), .ZN(G409));
  AND2_X1   g1037(.A1(G387), .A2(new_n1085), .ZN(new_n1238));
  NOR2_X1   g1038(.A1(G387), .A2(new_n1085), .ZN(new_n1239));
  AOI21_X1  g1039(.A(new_n816), .B1(new_n1027), .B2(new_n1060), .ZN(new_n1240));
  OAI22_X1  g1040(.A1(new_n1238), .A2(new_n1239), .B1(new_n1228), .B2(new_n1240), .ZN(new_n1241));
  OR2_X1    g1041(.A1(G387), .A2(new_n1085), .ZN(new_n1242));
  NOR2_X1   g1042(.A1(new_n1228), .A2(new_n1240), .ZN(new_n1243));
  NAND2_X1  g1043(.A1(G387), .A2(new_n1085), .ZN(new_n1244));
  NAND3_X1  g1044(.A1(new_n1242), .A2(new_n1243), .A3(new_n1244), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n1241), .A2(new_n1245), .ZN(new_n1246));
  NAND4_X1  g1046(.A1(new_n1134), .A2(new_n1137), .A3(new_n1132), .A4(KEYINPUT60), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n1247), .A2(new_n677), .ZN(new_n1248));
  OAI21_X1  g1048(.A(KEYINPUT60), .B1(new_n1224), .B2(new_n1132), .ZN(new_n1249));
  AOI21_X1  g1049(.A(new_n1248), .B1(new_n1203), .B2(new_n1249), .ZN(new_n1250));
  OAI21_X1  g1050(.A(new_n1229), .B1(new_n1250), .B2(new_n1225), .ZN(new_n1251));
  INV_X1    g1051(.A(new_n1203), .ZN(new_n1252));
  AOI21_X1  g1052(.A(new_n1252), .B1(KEYINPUT60), .B2(new_n1139), .ZN(new_n1253));
  OAI211_X1 g1053(.A(G384), .B(new_n1226), .C1(new_n1253), .C2(new_n1248), .ZN(new_n1254));
  OR2_X1    g1054(.A1(new_n1234), .A2(KEYINPUT125), .ZN(new_n1255));
  NAND3_X1  g1055(.A1(new_n1251), .A2(new_n1254), .A3(new_n1255), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(new_n1235), .A2(G2897), .ZN(new_n1257));
  INV_X1    g1057(.A(new_n1257), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(new_n1256), .A2(new_n1258), .ZN(new_n1259));
  NAND4_X1  g1059(.A1(new_n1251), .A2(new_n1254), .A3(new_n1257), .A4(new_n1255), .ZN(new_n1260));
  AOI21_X1  g1060(.A(KEYINPUT62), .B1(new_n1259), .B2(new_n1260), .ZN(new_n1261));
  INV_X1    g1061(.A(KEYINPUT127), .ZN(new_n1262));
  AND3_X1   g1062(.A1(new_n1167), .A2(new_n925), .A3(new_n1162), .ZN(new_n1263));
  AOI21_X1  g1063(.A(new_n925), .B1(new_n1167), .B2(new_n1162), .ZN(new_n1264));
  NOR2_X1   g1064(.A1(new_n1263), .A2(new_n1264), .ZN(new_n1265));
  AOI21_X1  g1065(.A(new_n1192), .B1(new_n1265), .B2(new_n735), .ZN(new_n1266));
  NAND3_X1  g1066(.A1(new_n1265), .A2(new_n1021), .A3(new_n1196), .ZN(new_n1267));
  AOI21_X1  g1067(.A(G378), .B1(new_n1266), .B2(new_n1267), .ZN(new_n1268));
  AOI21_X1  g1068(.A(new_n1268), .B1(G378), .B2(new_n1201), .ZN(new_n1269));
  OAI21_X1  g1069(.A(new_n1262), .B1(new_n1269), .B2(new_n1235), .ZN(new_n1270));
  NAND2_X1  g1070(.A1(new_n1197), .A2(new_n1198), .ZN(new_n1271));
  NAND3_X1  g1071(.A1(new_n1271), .A2(new_n677), .A3(new_n1200), .ZN(new_n1272));
  NAND3_X1  g1072(.A1(new_n1272), .A2(G378), .A3(new_n1266), .ZN(new_n1273));
  NOR2_X1   g1073(.A1(new_n1197), .A2(new_n1020), .ZN(new_n1274));
  OAI21_X1  g1074(.A(new_n1142), .B1(new_n1274), .B2(new_n1194), .ZN(new_n1275));
  AOI21_X1  g1075(.A(new_n1235), .B1(new_n1273), .B2(new_n1275), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(new_n1276), .A2(KEYINPUT127), .ZN(new_n1277));
  AOI21_X1  g1077(.A(new_n1261), .B1(new_n1270), .B2(new_n1277), .ZN(new_n1278));
  AND2_X1   g1078(.A1(new_n1251), .A2(new_n1254), .ZN(new_n1279));
  INV_X1    g1079(.A(new_n1279), .ZN(new_n1280));
  AOI21_X1  g1080(.A(KEYINPUT61), .B1(new_n1280), .B2(KEYINPUT62), .ZN(new_n1281));
  AOI211_X1 g1081(.A(new_n1142), .B(new_n1194), .C1(new_n1199), .C2(new_n1200), .ZN(new_n1282));
  OAI211_X1 g1082(.A(new_n1234), .B(new_n1279), .C1(new_n1282), .C2(new_n1268), .ZN(new_n1283));
  OAI21_X1  g1083(.A(new_n1281), .B1(new_n1283), .B2(KEYINPUT62), .ZN(new_n1284));
  OAI21_X1  g1084(.A(new_n1246), .B1(new_n1278), .B2(new_n1284), .ZN(new_n1285));
  INV_X1    g1085(.A(KEYINPUT63), .ZN(new_n1286));
  NOR2_X1   g1086(.A1(new_n1280), .A2(new_n1286), .ZN(new_n1287));
  NAND3_X1  g1087(.A1(new_n1270), .A2(new_n1277), .A3(new_n1287), .ZN(new_n1288));
  INV_X1    g1088(.A(KEYINPUT61), .ZN(new_n1289));
  NAND3_X1  g1089(.A1(new_n1241), .A2(new_n1245), .A3(new_n1289), .ZN(new_n1290));
  INV_X1    g1090(.A(KEYINPUT126), .ZN(new_n1291));
  AOI21_X1  g1091(.A(new_n1291), .B1(new_n1259), .B2(new_n1260), .ZN(new_n1292));
  NAND2_X1  g1092(.A1(new_n1273), .A2(new_n1275), .ZN(new_n1293));
  AOI21_X1  g1093(.A(new_n1292), .B1(new_n1293), .B2(new_n1234), .ZN(new_n1294));
  NAND3_X1  g1094(.A1(new_n1259), .A2(new_n1291), .A3(new_n1260), .ZN(new_n1295));
  AOI21_X1  g1095(.A(new_n1290), .B1(new_n1294), .B2(new_n1295), .ZN(new_n1296));
  INV_X1    g1096(.A(KEYINPUT124), .ZN(new_n1297));
  AOI211_X1 g1097(.A(new_n1297), .B(KEYINPUT63), .C1(new_n1276), .C2(new_n1279), .ZN(new_n1298));
  AOI21_X1  g1098(.A(KEYINPUT124), .B1(new_n1283), .B2(new_n1286), .ZN(new_n1299));
  OAI211_X1 g1099(.A(new_n1288), .B(new_n1296), .C1(new_n1298), .C2(new_n1299), .ZN(new_n1300));
  NAND2_X1  g1100(.A1(new_n1285), .A2(new_n1300), .ZN(G405));
  NAND2_X1  g1101(.A1(G375), .A2(new_n1142), .ZN(new_n1302));
  NAND2_X1  g1102(.A1(new_n1302), .A2(new_n1273), .ZN(new_n1303));
  NAND2_X1  g1103(.A1(new_n1303), .A2(new_n1279), .ZN(new_n1304));
  NAND3_X1  g1104(.A1(new_n1302), .A2(new_n1273), .A3(new_n1280), .ZN(new_n1305));
  NAND2_X1  g1105(.A1(new_n1304), .A2(new_n1305), .ZN(new_n1306));
  XNOR2_X1  g1106(.A(new_n1306), .B(new_n1246), .ZN(G402));
endmodule


