

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582;

  XOR2_X1 U320 ( .A(n570), .B(KEYINPUT41), .Z(n553) );
  AND2_X1 U321 ( .A1(G232GAT), .A2(G233GAT), .ZN(n288) );
  XNOR2_X1 U322 ( .A(KEYINPUT65), .B(KEYINPUT45), .ZN(n498) );
  XNOR2_X1 U323 ( .A(n499), .B(n498), .ZN(n500) );
  XNOR2_X1 U324 ( .A(n423), .B(n288), .ZN(n424) );
  XNOR2_X1 U325 ( .A(n425), .B(n424), .ZN(n426) );
  INV_X1 U326 ( .A(KEYINPUT54), .ZN(n540) );
  XNOR2_X1 U327 ( .A(n431), .B(n430), .ZN(n432) );
  XNOR2_X1 U328 ( .A(n541), .B(n540), .ZN(n542) );
  XNOR2_X1 U329 ( .A(n433), .B(n432), .ZN(n437) );
  AND2_X1 U330 ( .A1(n547), .A2(n546), .ZN(n559) );
  XNOR2_X1 U331 ( .A(G148GAT), .B(KEYINPUT3), .ZN(n289) );
  XNOR2_X1 U332 ( .A(n289), .B(KEYINPUT87), .ZN(n290) );
  XOR2_X1 U333 ( .A(n290), .B(KEYINPUT2), .Z(n292) );
  XNOR2_X1 U334 ( .A(G141GAT), .B(G162GAT), .ZN(n291) );
  XNOR2_X1 U335 ( .A(n292), .B(n291), .ZN(n393) );
  XOR2_X1 U336 ( .A(KEYINPUT93), .B(KEYINPUT91), .Z(n294) );
  XNOR2_X1 U337 ( .A(KEYINPUT6), .B(KEYINPUT90), .ZN(n293) );
  XNOR2_X1 U338 ( .A(n294), .B(n293), .ZN(n298) );
  XOR2_X1 U339 ( .A(KEYINPUT5), .B(KEYINPUT92), .Z(n296) );
  NAND2_X1 U340 ( .A1(G225GAT), .A2(G233GAT), .ZN(n295) );
  XNOR2_X1 U341 ( .A(n296), .B(n295), .ZN(n297) );
  XOR2_X1 U342 ( .A(n298), .B(n297), .Z(n305) );
  XOR2_X1 U343 ( .A(KEYINPUT79), .B(KEYINPUT0), .Z(n300) );
  XNOR2_X1 U344 ( .A(KEYINPUT78), .B(G120GAT), .ZN(n299) );
  XNOR2_X1 U345 ( .A(n300), .B(n299), .ZN(n301) );
  XOR2_X1 U346 ( .A(G113GAT), .B(n301), .Z(n375) );
  XOR2_X1 U347 ( .A(G57GAT), .B(G155GAT), .Z(n303) );
  XNOR2_X1 U348 ( .A(G1GAT), .B(G127GAT), .ZN(n302) );
  XNOR2_X1 U349 ( .A(n303), .B(n302), .ZN(n414) );
  XNOR2_X1 U350 ( .A(n375), .B(n414), .ZN(n304) );
  XNOR2_X1 U351 ( .A(n305), .B(n304), .ZN(n306) );
  XOR2_X1 U352 ( .A(n306), .B(KEYINPUT1), .Z(n309) );
  XNOR2_X1 U353 ( .A(G29GAT), .B(G134GAT), .ZN(n307) );
  XNOR2_X1 U354 ( .A(n307), .B(G85GAT), .ZN(n434) );
  XNOR2_X1 U355 ( .A(n434), .B(KEYINPUT4), .ZN(n308) );
  XNOR2_X1 U356 ( .A(n309), .B(n308), .ZN(n310) );
  XNOR2_X1 U357 ( .A(n393), .B(n310), .ZN(n402) );
  XNOR2_X1 U358 ( .A(KEYINPUT94), .B(n402), .ZN(n543) );
  INV_X1 U359 ( .A(n543), .ZN(n479) );
  XOR2_X1 U360 ( .A(G141GAT), .B(G113GAT), .Z(n312) );
  XNOR2_X1 U361 ( .A(G169GAT), .B(G50GAT), .ZN(n311) );
  XNOR2_X1 U362 ( .A(n312), .B(n311), .ZN(n327) );
  XOR2_X1 U363 ( .A(G15GAT), .B(G22GAT), .Z(n409) );
  XOR2_X1 U364 ( .A(n409), .B(G29GAT), .Z(n316) );
  XOR2_X1 U365 ( .A(G43GAT), .B(KEYINPUT7), .Z(n314) );
  XNOR2_X1 U366 ( .A(KEYINPUT8), .B(KEYINPUT68), .ZN(n313) );
  XNOR2_X1 U367 ( .A(n314), .B(n313), .ZN(n435) );
  XNOR2_X1 U368 ( .A(G36GAT), .B(n435), .ZN(n315) );
  XNOR2_X1 U369 ( .A(n316), .B(n315), .ZN(n320) );
  XOR2_X1 U370 ( .A(G8GAT), .B(KEYINPUT69), .Z(n318) );
  NAND2_X1 U371 ( .A1(G229GAT), .A2(G233GAT), .ZN(n317) );
  XNOR2_X1 U372 ( .A(n318), .B(n317), .ZN(n319) );
  XOR2_X1 U373 ( .A(n320), .B(n319), .Z(n325) );
  XOR2_X1 U374 ( .A(KEYINPUT67), .B(KEYINPUT30), .Z(n322) );
  XNOR2_X1 U375 ( .A(G197GAT), .B(G1GAT), .ZN(n321) );
  XNOR2_X1 U376 ( .A(n322), .B(n321), .ZN(n323) );
  XNOR2_X1 U377 ( .A(n323), .B(KEYINPUT29), .ZN(n324) );
  XNOR2_X1 U378 ( .A(n325), .B(n324), .ZN(n326) );
  XOR2_X1 U379 ( .A(n327), .B(n326), .Z(n566) );
  INV_X1 U380 ( .A(n566), .ZN(n511) );
  XOR2_X1 U381 ( .A(KEYINPUT71), .B(KEYINPUT72), .Z(n329) );
  NAND2_X1 U382 ( .A1(G230GAT), .A2(G233GAT), .ZN(n328) );
  XNOR2_X1 U383 ( .A(n329), .B(n328), .ZN(n330) );
  XOR2_X1 U384 ( .A(n330), .B(KEYINPUT32), .Z(n338) );
  XOR2_X1 U385 ( .A(G85GAT), .B(G148GAT), .Z(n332) );
  XNOR2_X1 U386 ( .A(G120GAT), .B(G99GAT), .ZN(n331) );
  XNOR2_X1 U387 ( .A(n332), .B(n331), .ZN(n336) );
  XOR2_X1 U388 ( .A(KEYINPUT70), .B(KEYINPUT33), .Z(n334) );
  XNOR2_X1 U389 ( .A(G57GAT), .B(KEYINPUT31), .ZN(n333) );
  XNOR2_X1 U390 ( .A(n334), .B(n333), .ZN(n335) );
  XNOR2_X1 U391 ( .A(n336), .B(n335), .ZN(n337) );
  XNOR2_X1 U392 ( .A(n338), .B(n337), .ZN(n341) );
  XOR2_X1 U393 ( .A(G64GAT), .B(G92GAT), .Z(n340) );
  XNOR2_X1 U394 ( .A(G176GAT), .B(G204GAT), .ZN(n339) );
  XNOR2_X1 U395 ( .A(n340), .B(n339), .ZN(n347) );
  XOR2_X1 U396 ( .A(n341), .B(n347), .Z(n343) );
  XOR2_X1 U397 ( .A(G106GAT), .B(G78GAT), .Z(n377) );
  XOR2_X1 U398 ( .A(G71GAT), .B(KEYINPUT13), .Z(n418) );
  XNOR2_X1 U399 ( .A(n377), .B(n418), .ZN(n342) );
  XNOR2_X1 U400 ( .A(n343), .B(n342), .ZN(n570) );
  NAND2_X1 U401 ( .A1(n511), .A2(n570), .ZN(n344) );
  XNOR2_X1 U402 ( .A(n344), .B(KEYINPUT73), .ZN(n455) );
  XNOR2_X1 U403 ( .A(G36GAT), .B(G190GAT), .ZN(n345) );
  XNOR2_X1 U404 ( .A(n345), .B(G218GAT), .ZN(n427) );
  XNOR2_X1 U405 ( .A(G8GAT), .B(G183GAT), .ZN(n346) );
  XNOR2_X1 U406 ( .A(n346), .B(KEYINPUT76), .ZN(n413) );
  XOR2_X1 U407 ( .A(n413), .B(n347), .Z(n355) );
  XNOR2_X1 U408 ( .A(KEYINPUT83), .B(KEYINPUT17), .ZN(n348) );
  XNOR2_X1 U409 ( .A(n348), .B(KEYINPUT19), .ZN(n349) );
  XOR2_X1 U410 ( .A(n349), .B(KEYINPUT18), .Z(n351) );
  XNOR2_X1 U411 ( .A(G169GAT), .B(KEYINPUT82), .ZN(n350) );
  XNOR2_X1 U412 ( .A(n351), .B(n350), .ZN(n371) );
  XOR2_X1 U413 ( .A(G211GAT), .B(KEYINPUT21), .Z(n353) );
  XNOR2_X1 U414 ( .A(G197GAT), .B(KEYINPUT86), .ZN(n352) );
  XNOR2_X1 U415 ( .A(n353), .B(n352), .ZN(n385) );
  XNOR2_X1 U416 ( .A(n371), .B(n385), .ZN(n354) );
  XNOR2_X1 U417 ( .A(n355), .B(n354), .ZN(n356) );
  XOR2_X1 U418 ( .A(n427), .B(n356), .Z(n358) );
  NAND2_X1 U419 ( .A1(G226GAT), .A2(G233GAT), .ZN(n357) );
  XNOR2_X1 U420 ( .A(n358), .B(n357), .ZN(n537) );
  XOR2_X1 U421 ( .A(G183GAT), .B(KEYINPUT84), .Z(n360) );
  XNOR2_X1 U422 ( .A(KEYINPUT20), .B(KEYINPUT80), .ZN(n359) );
  XNOR2_X1 U423 ( .A(n360), .B(n359), .ZN(n364) );
  XOR2_X1 U424 ( .A(G71GAT), .B(G127GAT), .Z(n362) );
  XNOR2_X1 U425 ( .A(G176GAT), .B(KEYINPUT81), .ZN(n361) );
  XNOR2_X1 U426 ( .A(n362), .B(n361), .ZN(n363) );
  XOR2_X1 U427 ( .A(n364), .B(n363), .Z(n373) );
  XOR2_X1 U428 ( .A(G134GAT), .B(G190GAT), .Z(n366) );
  XNOR2_X1 U429 ( .A(G43GAT), .B(G99GAT), .ZN(n365) );
  XNOR2_X1 U430 ( .A(n366), .B(n365), .ZN(n367) );
  XOR2_X1 U431 ( .A(G15GAT), .B(n367), .Z(n369) );
  NAND2_X1 U432 ( .A1(G227GAT), .A2(G233GAT), .ZN(n368) );
  XNOR2_X1 U433 ( .A(n369), .B(n368), .ZN(n370) );
  XNOR2_X1 U434 ( .A(n371), .B(n370), .ZN(n372) );
  XNOR2_X1 U435 ( .A(n373), .B(n372), .ZN(n374) );
  XNOR2_X1 U436 ( .A(n375), .B(n374), .ZN(n546) );
  NAND2_X1 U437 ( .A1(n537), .A2(n546), .ZN(n376) );
  XNOR2_X1 U438 ( .A(n376), .B(KEYINPUT96), .ZN(n394) );
  XNOR2_X1 U439 ( .A(n377), .B(G218GAT), .ZN(n378) );
  XNOR2_X1 U440 ( .A(n378), .B(KEYINPUT85), .ZN(n382) );
  XOR2_X1 U441 ( .A(G155GAT), .B(KEYINPUT23), .Z(n380) );
  XNOR2_X1 U442 ( .A(KEYINPUT88), .B(KEYINPUT24), .ZN(n379) );
  XNOR2_X1 U443 ( .A(n380), .B(n379), .ZN(n381) );
  XOR2_X1 U444 ( .A(n382), .B(n381), .Z(n391) );
  XOR2_X1 U445 ( .A(G204GAT), .B(KEYINPUT89), .Z(n384) );
  XNOR2_X1 U446 ( .A(G22GAT), .B(KEYINPUT22), .ZN(n383) );
  XNOR2_X1 U447 ( .A(n384), .B(n383), .ZN(n389) );
  XOR2_X1 U448 ( .A(G50GAT), .B(KEYINPUT74), .Z(n423) );
  XOR2_X1 U449 ( .A(n423), .B(n385), .Z(n387) );
  NAND2_X1 U450 ( .A1(G228GAT), .A2(G233GAT), .ZN(n386) );
  XNOR2_X1 U451 ( .A(n387), .B(n386), .ZN(n388) );
  XNOR2_X1 U452 ( .A(n389), .B(n388), .ZN(n390) );
  XNOR2_X1 U453 ( .A(n391), .B(n390), .ZN(n392) );
  XNOR2_X1 U454 ( .A(n393), .B(n392), .ZN(n544) );
  NAND2_X1 U455 ( .A1(n394), .A2(n544), .ZN(n396) );
  XOR2_X1 U456 ( .A(KEYINPUT25), .B(KEYINPUT97), .Z(n395) );
  XNOR2_X1 U457 ( .A(n396), .B(n395), .ZN(n400) );
  XOR2_X1 U458 ( .A(n537), .B(KEYINPUT27), .Z(n403) );
  NOR2_X1 U459 ( .A1(n546), .A2(n544), .ZN(n398) );
  XNOR2_X1 U460 ( .A(KEYINPUT95), .B(KEYINPUT26), .ZN(n397) );
  XNOR2_X1 U461 ( .A(n398), .B(n397), .ZN(n526) );
  NOR2_X1 U462 ( .A1(n403), .A2(n526), .ZN(n399) );
  NOR2_X1 U463 ( .A1(n400), .A2(n399), .ZN(n401) );
  NOR2_X1 U464 ( .A1(n402), .A2(n401), .ZN(n406) );
  NOR2_X1 U465 ( .A1(n403), .A2(n479), .ZN(n506) );
  XNOR2_X1 U466 ( .A(KEYINPUT28), .B(n544), .ZN(n488) );
  NAND2_X1 U467 ( .A1(n506), .A2(n488), .ZN(n404) );
  NOR2_X1 U468 ( .A1(n404), .A2(n546), .ZN(n405) );
  NOR2_X1 U469 ( .A1(n406), .A2(n405), .ZN(n450) );
  XOR2_X1 U470 ( .A(KEYINPUT16), .B(KEYINPUT77), .Z(n439) );
  XOR2_X1 U471 ( .A(KEYINPUT12), .B(KEYINPUT15), .Z(n408) );
  XNOR2_X1 U472 ( .A(G64GAT), .B(KEYINPUT14), .ZN(n407) );
  XNOR2_X1 U473 ( .A(n408), .B(n407), .ZN(n412) );
  XNOR2_X1 U474 ( .A(n409), .B(G211GAT), .ZN(n410) );
  XNOR2_X1 U475 ( .A(n410), .B(G78GAT), .ZN(n411) );
  XOR2_X1 U476 ( .A(n412), .B(n411), .Z(n416) );
  XNOR2_X1 U477 ( .A(n414), .B(n413), .ZN(n415) );
  XNOR2_X1 U478 ( .A(n416), .B(n415), .ZN(n417) );
  XOR2_X1 U479 ( .A(n418), .B(n417), .Z(n420) );
  NAND2_X1 U480 ( .A1(G231GAT), .A2(G233GAT), .ZN(n419) );
  XNOR2_X1 U481 ( .A(n420), .B(n419), .ZN(n575) );
  INV_X1 U482 ( .A(n575), .ZN(n497) );
  XOR2_X1 U483 ( .A(KEYINPUT75), .B(G92GAT), .Z(n422) );
  XNOR2_X1 U484 ( .A(G162GAT), .B(G106GAT), .ZN(n421) );
  XNOR2_X1 U485 ( .A(n422), .B(n421), .ZN(n425) );
  XOR2_X1 U486 ( .A(n426), .B(KEYINPUT11), .Z(n433) );
  XNOR2_X1 U487 ( .A(n427), .B(KEYINPUT64), .ZN(n431) );
  XOR2_X1 U488 ( .A(KEYINPUT66), .B(KEYINPUT9), .Z(n429) );
  XNOR2_X1 U489 ( .A(G99GAT), .B(KEYINPUT10), .ZN(n428) );
  XOR2_X1 U490 ( .A(n429), .B(n428), .Z(n430) );
  XNOR2_X1 U491 ( .A(n435), .B(n434), .ZN(n436) );
  XNOR2_X1 U492 ( .A(n437), .B(n436), .ZN(n558) );
  INV_X1 U493 ( .A(n558), .ZN(n535) );
  NAND2_X1 U494 ( .A1(n497), .A2(n535), .ZN(n438) );
  XNOR2_X1 U495 ( .A(n439), .B(n438), .ZN(n440) );
  NOR2_X1 U496 ( .A1(n450), .A2(n440), .ZN(n467) );
  NAND2_X1 U497 ( .A1(n455), .A2(n467), .ZN(n448) );
  NOR2_X1 U498 ( .A1(n479), .A2(n448), .ZN(n441) );
  XOR2_X1 U499 ( .A(KEYINPUT34), .B(n441), .Z(n442) );
  XNOR2_X1 U500 ( .A(G1GAT), .B(n442), .ZN(G1324GAT) );
  INV_X1 U501 ( .A(n537), .ZN(n481) );
  NOR2_X1 U502 ( .A1(n481), .A2(n448), .ZN(n443) );
  XOR2_X1 U503 ( .A(G8GAT), .B(n443), .Z(G1325GAT) );
  INV_X1 U504 ( .A(n546), .ZN(n484) );
  NOR2_X1 U505 ( .A1(n448), .A2(n484), .ZN(n447) );
  XOR2_X1 U506 ( .A(KEYINPUT98), .B(KEYINPUT99), .Z(n445) );
  XNOR2_X1 U507 ( .A(G15GAT), .B(KEYINPUT35), .ZN(n444) );
  XNOR2_X1 U508 ( .A(n445), .B(n444), .ZN(n446) );
  XNOR2_X1 U509 ( .A(n447), .B(n446), .ZN(G1326GAT) );
  NOR2_X1 U510 ( .A1(n488), .A2(n448), .ZN(n449) );
  XOR2_X1 U511 ( .A(G22GAT), .B(n449), .Z(G1327GAT) );
  XOR2_X1 U512 ( .A(KEYINPUT38), .B(KEYINPUT102), .Z(n457) );
  NOR2_X1 U513 ( .A1(n450), .A2(n497), .ZN(n451) );
  XNOR2_X1 U514 ( .A(n451), .B(KEYINPUT100), .ZN(n452) );
  XNOR2_X1 U515 ( .A(KEYINPUT36), .B(n558), .ZN(n580) );
  NAND2_X1 U516 ( .A1(n452), .A2(n580), .ZN(n454) );
  XOR2_X1 U517 ( .A(KEYINPUT37), .B(KEYINPUT101), .Z(n453) );
  XNOR2_X1 U518 ( .A(n454), .B(n453), .ZN(n478) );
  NAND2_X1 U519 ( .A1(n455), .A2(n478), .ZN(n456) );
  XNOR2_X1 U520 ( .A(n457), .B(n456), .ZN(n464) );
  NAND2_X1 U521 ( .A1(n464), .A2(n543), .ZN(n460) );
  XNOR2_X1 U522 ( .A(G29GAT), .B(KEYINPUT103), .ZN(n458) );
  XNOR2_X1 U523 ( .A(n458), .B(KEYINPUT39), .ZN(n459) );
  XNOR2_X1 U524 ( .A(n460), .B(n459), .ZN(G1328GAT) );
  NAND2_X1 U525 ( .A1(n464), .A2(n537), .ZN(n461) );
  XNOR2_X1 U526 ( .A(n461), .B(G36GAT), .ZN(G1329GAT) );
  NAND2_X1 U527 ( .A1(n546), .A2(n464), .ZN(n462) );
  XNOR2_X1 U528 ( .A(n462), .B(KEYINPUT40), .ZN(n463) );
  XNOR2_X1 U529 ( .A(G43GAT), .B(n463), .ZN(G1330GAT) );
  XNOR2_X1 U530 ( .A(G50GAT), .B(KEYINPUT104), .ZN(n466) );
  INV_X1 U531 ( .A(n488), .ZN(n510) );
  NAND2_X1 U532 ( .A1(n464), .A2(n510), .ZN(n465) );
  XNOR2_X1 U533 ( .A(n466), .B(n465), .ZN(G1331GAT) );
  NOR2_X1 U534 ( .A1(n553), .A2(n511), .ZN(n477) );
  NAND2_X1 U535 ( .A1(n477), .A2(n467), .ZN(n473) );
  NOR2_X1 U536 ( .A1(n479), .A2(n473), .ZN(n468) );
  XOR2_X1 U537 ( .A(G57GAT), .B(n468), .Z(n469) );
  XNOR2_X1 U538 ( .A(KEYINPUT42), .B(n469), .ZN(G1332GAT) );
  NOR2_X1 U539 ( .A1(n481), .A2(n473), .ZN(n470) );
  XOR2_X1 U540 ( .A(G64GAT), .B(n470), .Z(G1333GAT) );
  NOR2_X1 U541 ( .A1(n484), .A2(n473), .ZN(n472) );
  XNOR2_X1 U542 ( .A(G71GAT), .B(KEYINPUT105), .ZN(n471) );
  XNOR2_X1 U543 ( .A(n472), .B(n471), .ZN(G1334GAT) );
  NOR2_X1 U544 ( .A1(n488), .A2(n473), .ZN(n475) );
  XNOR2_X1 U545 ( .A(KEYINPUT106), .B(KEYINPUT43), .ZN(n474) );
  XNOR2_X1 U546 ( .A(n475), .B(n474), .ZN(n476) );
  XNOR2_X1 U547 ( .A(G78GAT), .B(n476), .ZN(G1335GAT) );
  NAND2_X1 U548 ( .A1(n478), .A2(n477), .ZN(n487) );
  NOR2_X1 U549 ( .A1(n479), .A2(n487), .ZN(n480) );
  XOR2_X1 U550 ( .A(G85GAT), .B(n480), .Z(G1336GAT) );
  NOR2_X1 U551 ( .A1(n481), .A2(n487), .ZN(n483) );
  XNOR2_X1 U552 ( .A(G92GAT), .B(KEYINPUT107), .ZN(n482) );
  XNOR2_X1 U553 ( .A(n483), .B(n482), .ZN(G1337GAT) );
  NOR2_X1 U554 ( .A1(n484), .A2(n487), .ZN(n485) );
  XOR2_X1 U555 ( .A(KEYINPUT108), .B(n485), .Z(n486) );
  XNOR2_X1 U556 ( .A(G99GAT), .B(n486), .ZN(G1338GAT) );
  NOR2_X1 U557 ( .A1(n488), .A2(n487), .ZN(n490) );
  XNOR2_X1 U558 ( .A(KEYINPUT44), .B(KEYINPUT109), .ZN(n489) );
  XNOR2_X1 U559 ( .A(n490), .B(n489), .ZN(n491) );
  XNOR2_X1 U560 ( .A(G106GAT), .B(n491), .ZN(G1339GAT) );
  XOR2_X1 U561 ( .A(n575), .B(KEYINPUT110), .Z(n556) );
  NOR2_X1 U562 ( .A1(n558), .A2(n556), .ZN(n495) );
  XOR2_X1 U563 ( .A(KEYINPUT46), .B(KEYINPUT111), .Z(n493) );
  NOR2_X1 U564 ( .A1(n566), .A2(n553), .ZN(n492) );
  XOR2_X1 U565 ( .A(n493), .B(n492), .Z(n494) );
  NAND2_X1 U566 ( .A1(n495), .A2(n494), .ZN(n496) );
  XNOR2_X1 U567 ( .A(n496), .B(KEYINPUT47), .ZN(n504) );
  NAND2_X1 U568 ( .A1(n580), .A2(n497), .ZN(n499) );
  NAND2_X1 U569 ( .A1(n500), .A2(n570), .ZN(n501) );
  XNOR2_X1 U570 ( .A(KEYINPUT112), .B(n501), .ZN(n502) );
  NOR2_X1 U571 ( .A1(n511), .A2(n502), .ZN(n503) );
  NOR2_X1 U572 ( .A1(n504), .A2(n503), .ZN(n505) );
  XNOR2_X1 U573 ( .A(n505), .B(KEYINPUT48), .ZN(n539) );
  INV_X1 U574 ( .A(n506), .ZN(n507) );
  NOR2_X1 U575 ( .A1(n539), .A2(n507), .ZN(n527) );
  NAND2_X1 U576 ( .A1(n527), .A2(n546), .ZN(n508) );
  XOR2_X1 U577 ( .A(KEYINPUT113), .B(n508), .Z(n509) );
  NOR2_X1 U578 ( .A1(n510), .A2(n509), .ZN(n521) );
  NAND2_X1 U579 ( .A1(n511), .A2(n521), .ZN(n512) );
  XNOR2_X1 U580 ( .A(n512), .B(G113GAT), .ZN(G1340GAT) );
  XOR2_X1 U581 ( .A(G120GAT), .B(KEYINPUT114), .Z(n515) );
  INV_X1 U582 ( .A(n553), .ZN(n513) );
  NAND2_X1 U583 ( .A1(n521), .A2(n513), .ZN(n514) );
  XNOR2_X1 U584 ( .A(n515), .B(n514), .ZN(n517) );
  XOR2_X1 U585 ( .A(KEYINPUT115), .B(KEYINPUT49), .Z(n516) );
  XNOR2_X1 U586 ( .A(n517), .B(n516), .ZN(G1341GAT) );
  XOR2_X1 U587 ( .A(KEYINPUT116), .B(KEYINPUT50), .Z(n519) );
  NAND2_X1 U588 ( .A1(n521), .A2(n556), .ZN(n518) );
  XNOR2_X1 U589 ( .A(n519), .B(n518), .ZN(n520) );
  XOR2_X1 U590 ( .A(G127GAT), .B(n520), .Z(G1342GAT) );
  XOR2_X1 U591 ( .A(KEYINPUT118), .B(KEYINPUT51), .Z(n523) );
  NAND2_X1 U592 ( .A1(n521), .A2(n558), .ZN(n522) );
  XNOR2_X1 U593 ( .A(n523), .B(n522), .ZN(n525) );
  XOR2_X1 U594 ( .A(G134GAT), .B(KEYINPUT117), .Z(n524) );
  XNOR2_X1 U595 ( .A(n525), .B(n524), .ZN(G1343GAT) );
  INV_X1 U596 ( .A(n526), .ZN(n564) );
  NAND2_X1 U597 ( .A1(n527), .A2(n564), .ZN(n534) );
  NOR2_X1 U598 ( .A1(n566), .A2(n534), .ZN(n528) );
  XOR2_X1 U599 ( .A(G141GAT), .B(n528), .Z(G1344GAT) );
  NOR2_X1 U600 ( .A1(n534), .A2(n553), .ZN(n532) );
  XOR2_X1 U601 ( .A(KEYINPUT53), .B(KEYINPUT52), .Z(n530) );
  XNOR2_X1 U602 ( .A(G148GAT), .B(KEYINPUT119), .ZN(n529) );
  XNOR2_X1 U603 ( .A(n530), .B(n529), .ZN(n531) );
  XNOR2_X1 U604 ( .A(n532), .B(n531), .ZN(G1345GAT) );
  NOR2_X1 U605 ( .A1(n575), .A2(n534), .ZN(n533) );
  XOR2_X1 U606 ( .A(G155GAT), .B(n533), .Z(G1346GAT) );
  NOR2_X1 U607 ( .A1(n535), .A2(n534), .ZN(n536) );
  XOR2_X1 U608 ( .A(G162GAT), .B(n536), .Z(G1347GAT) );
  XOR2_X1 U609 ( .A(KEYINPUT120), .B(n537), .Z(n538) );
  NOR2_X1 U610 ( .A1(n539), .A2(n538), .ZN(n541) );
  NOR2_X1 U611 ( .A1(n543), .A2(n542), .ZN(n565) );
  NAND2_X1 U612 ( .A1(n565), .A2(n544), .ZN(n545) );
  XNOR2_X1 U613 ( .A(n545), .B(KEYINPUT55), .ZN(n547) );
  INV_X1 U614 ( .A(n559), .ZN(n552) );
  NOR2_X1 U615 ( .A1(n566), .A2(n552), .ZN(n549) );
  XNOR2_X1 U616 ( .A(G169GAT), .B(KEYINPUT121), .ZN(n548) );
  XNOR2_X1 U617 ( .A(n549), .B(n548), .ZN(G1348GAT) );
  XOR2_X1 U618 ( .A(KEYINPUT56), .B(KEYINPUT122), .Z(n551) );
  XNOR2_X1 U619 ( .A(G176GAT), .B(KEYINPUT57), .ZN(n550) );
  XNOR2_X1 U620 ( .A(n551), .B(n550), .ZN(n555) );
  NOR2_X1 U621 ( .A1(n553), .A2(n552), .ZN(n554) );
  XOR2_X1 U622 ( .A(n555), .B(n554), .Z(G1349GAT) );
  NAND2_X1 U623 ( .A1(n559), .A2(n556), .ZN(n557) );
  XNOR2_X1 U624 ( .A(n557), .B(G183GAT), .ZN(G1350GAT) );
  XNOR2_X1 U625 ( .A(G190GAT), .B(KEYINPUT123), .ZN(n563) );
  XOR2_X1 U626 ( .A(KEYINPUT58), .B(KEYINPUT124), .Z(n561) );
  NAND2_X1 U627 ( .A1(n559), .A2(n558), .ZN(n560) );
  XNOR2_X1 U628 ( .A(n561), .B(n560), .ZN(n562) );
  XNOR2_X1 U629 ( .A(n563), .B(n562), .ZN(G1351GAT) );
  NAND2_X1 U630 ( .A1(n565), .A2(n564), .ZN(n578) );
  NOR2_X1 U631 ( .A1(n566), .A2(n578), .ZN(n568) );
  XNOR2_X1 U632 ( .A(KEYINPUT60), .B(KEYINPUT59), .ZN(n567) );
  XNOR2_X1 U633 ( .A(n568), .B(n567), .ZN(n569) );
  XNOR2_X1 U634 ( .A(G197GAT), .B(n569), .ZN(G1352GAT) );
  NOR2_X1 U635 ( .A1(n578), .A2(n570), .ZN(n574) );
  XOR2_X1 U636 ( .A(KEYINPUT125), .B(KEYINPUT126), .Z(n572) );
  XNOR2_X1 U637 ( .A(G204GAT), .B(KEYINPUT61), .ZN(n571) );
  XNOR2_X1 U638 ( .A(n572), .B(n571), .ZN(n573) );
  XNOR2_X1 U639 ( .A(n574), .B(n573), .ZN(G1353GAT) );
  NOR2_X1 U640 ( .A1(n575), .A2(n578), .ZN(n577) );
  XNOR2_X1 U641 ( .A(G211GAT), .B(KEYINPUT127), .ZN(n576) );
  XNOR2_X1 U642 ( .A(n577), .B(n576), .ZN(G1354GAT) );
  INV_X1 U643 ( .A(n578), .ZN(n579) );
  NAND2_X1 U644 ( .A1(n580), .A2(n579), .ZN(n581) );
  XNOR2_X1 U645 ( .A(n581), .B(KEYINPUT62), .ZN(n582) );
  XNOR2_X1 U646 ( .A(G218GAT), .B(n582), .ZN(G1355GAT) );
endmodule

