//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 0 1 0 0 0 0 0 0 0 1 1 1 1 1 0 1 1 0 0 1 0 0 0 1 0 1 0 1 0 1 0 1 0 0 1 0 1 0 0 0 1 1 1 1 1 1 0 1 1 1 1 1 1 0 1 1 1 0 1 0 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:40:47 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n202, new_n203, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n227, new_n228, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n236, new_n237, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n244, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1257, new_n1258, new_n1259, new_n1260,
    new_n1261, new_n1262, new_n1263, new_n1264, new_n1265, new_n1267,
    new_n1268, new_n1269, new_n1270, new_n1271, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1338, new_n1339, new_n1340, new_n1341,
    new_n1342;
  NOR4_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .A4(G77), .ZN(G353));
  OAI21_X1  g0001(.A(G87), .B1(G97), .B2(G107), .ZN(new_n202));
  XNOR2_X1  g0002(.A(new_n202), .B(KEYINPUT64), .ZN(new_n203));
  INV_X1    g0003(.A(new_n203), .ZN(G355));
  INV_X1    g0004(.A(G1), .ZN(new_n205));
  INV_X1    g0005(.A(G20), .ZN(new_n206));
  NOR2_X1   g0006(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  INV_X1    g0007(.A(new_n207), .ZN(new_n208));
  NOR2_X1   g0008(.A1(new_n208), .A2(G13), .ZN(new_n209));
  OAI211_X1 g0009(.A(new_n209), .B(G250), .C1(G257), .C2(G264), .ZN(new_n210));
  XNOR2_X1  g0010(.A(new_n210), .B(KEYINPUT0), .ZN(new_n211));
  OAI21_X1  g0011(.A(G50), .B1(G58), .B2(G68), .ZN(new_n212));
  INV_X1    g0012(.A(new_n212), .ZN(new_n213));
  NAND2_X1  g0013(.A1(G1), .A2(G13), .ZN(new_n214));
  NOR2_X1   g0014(.A1(new_n214), .A2(new_n206), .ZN(new_n215));
  NAND2_X1  g0015(.A1(new_n213), .A2(new_n215), .ZN(new_n216));
  XNOR2_X1  g0016(.A(KEYINPUT65), .B(G244), .ZN(new_n217));
  AND2_X1   g0017(.A1(new_n217), .A2(G77), .ZN(new_n218));
  AOI22_X1  g0018(.A1(G58), .A2(G232), .B1(G87), .B2(G250), .ZN(new_n219));
  AOI22_X1  g0019(.A1(G50), .A2(G226), .B1(G107), .B2(G264), .ZN(new_n220));
  AOI22_X1  g0020(.A1(G68), .A2(G238), .B1(G97), .B2(G257), .ZN(new_n221));
  NAND2_X1  g0021(.A1(G116), .A2(G270), .ZN(new_n222));
  NAND4_X1  g0022(.A1(new_n219), .A2(new_n220), .A3(new_n221), .A4(new_n222), .ZN(new_n223));
  OAI21_X1  g0023(.A(new_n208), .B1(new_n218), .B2(new_n223), .ZN(new_n224));
  OAI211_X1 g0024(.A(new_n211), .B(new_n216), .C1(KEYINPUT1), .C2(new_n224), .ZN(new_n225));
  AOI21_X1  g0025(.A(new_n225), .B1(KEYINPUT1), .B2(new_n224), .ZN(G361));
  XNOR2_X1  g0026(.A(G238), .B(G244), .ZN(new_n227));
  INV_X1    g0027(.A(G232), .ZN(new_n228));
  XNOR2_X1  g0028(.A(new_n227), .B(new_n228), .ZN(new_n229));
  XNOR2_X1  g0029(.A(KEYINPUT2), .B(G226), .ZN(new_n230));
  XNOR2_X1  g0030(.A(new_n229), .B(new_n230), .ZN(new_n231));
  XNOR2_X1  g0031(.A(G250), .B(G257), .ZN(new_n232));
  XNOR2_X1  g0032(.A(G264), .B(G270), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n232), .B(new_n233), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n231), .B(new_n234), .ZN(G358));
  XNOR2_X1  g0035(.A(G68), .B(G77), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n236), .B(KEYINPUT66), .ZN(new_n237));
  XOR2_X1   g0037(.A(G50), .B(G58), .Z(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XNOR2_X1  g0039(.A(G87), .B(G97), .ZN(new_n240));
  XNOR2_X1  g0040(.A(G107), .B(G116), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n239), .B(new_n242), .ZN(G351));
  NAND2_X1  g0043(.A1(new_n205), .A2(G20), .ZN(new_n244));
  NAND2_X1  g0044(.A1(new_n244), .A2(G50), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n245), .B(KEYINPUT69), .ZN(new_n246));
  NAND3_X1  g0046(.A1(new_n205), .A2(G13), .A3(G20), .ZN(new_n247));
  NAND3_X1  g0047(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n248));
  NAND3_X1  g0048(.A1(new_n247), .A2(new_n214), .A3(new_n248), .ZN(new_n249));
  INV_X1    g0049(.A(new_n249), .ZN(new_n250));
  NAND2_X1  g0050(.A1(new_n246), .A2(new_n250), .ZN(new_n251));
  INV_X1    g0051(.A(new_n247), .ZN(new_n252));
  INV_X1    g0052(.A(G50), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n252), .A2(new_n253), .ZN(new_n254));
  NAND2_X1  g0054(.A1(new_n251), .A2(new_n254), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n248), .A2(new_n214), .ZN(new_n256));
  INV_X1    g0056(.A(new_n256), .ZN(new_n257));
  INV_X1    g0057(.A(G58), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n258), .A2(KEYINPUT8), .ZN(new_n259));
  INV_X1    g0059(.A(KEYINPUT8), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n260), .A2(G58), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n259), .A2(new_n261), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n262), .A2(KEYINPUT68), .ZN(new_n263));
  XNOR2_X1  g0063(.A(KEYINPUT8), .B(G58), .ZN(new_n264));
  INV_X1    g0064(.A(KEYINPUT68), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n206), .A2(G33), .ZN(new_n267));
  INV_X1    g0067(.A(new_n267), .ZN(new_n268));
  NAND3_X1  g0068(.A1(new_n263), .A2(new_n266), .A3(new_n268), .ZN(new_n269));
  INV_X1    g0069(.A(G68), .ZN(new_n270));
  NAND3_X1  g0070(.A1(new_n253), .A2(new_n258), .A3(new_n270), .ZN(new_n271));
  NOR2_X1   g0071(.A1(G20), .A2(G33), .ZN(new_n272));
  AOI22_X1  g0072(.A1(new_n271), .A2(G20), .B1(G150), .B2(new_n272), .ZN(new_n273));
  AOI21_X1  g0073(.A(new_n257), .B1(new_n269), .B2(new_n273), .ZN(new_n274));
  NOR2_X1   g0074(.A1(new_n255), .A2(new_n274), .ZN(new_n275));
  INV_X1    g0075(.A(G169), .ZN(new_n276));
  INV_X1    g0076(.A(new_n214), .ZN(new_n277));
  NAND2_X1  g0077(.A1(G33), .A2(G41), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  INV_X1    g0079(.A(G1698), .ZN(new_n280));
  OR2_X1    g0080(.A1(KEYINPUT3), .A2(G33), .ZN(new_n281));
  NAND2_X1  g0081(.A1(KEYINPUT3), .A2(G33), .ZN(new_n282));
  AOI21_X1  g0082(.A(new_n280), .B1(new_n281), .B2(new_n282), .ZN(new_n283));
  AND2_X1   g0083(.A1(KEYINPUT3), .A2(G33), .ZN(new_n284));
  NOR2_X1   g0084(.A1(KEYINPUT3), .A2(G33), .ZN(new_n285));
  NOR2_X1   g0085(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  AOI22_X1  g0086(.A1(new_n283), .A2(G223), .B1(new_n286), .B2(G77), .ZN(new_n287));
  AOI21_X1  g0087(.A(G1698), .B1(new_n281), .B2(new_n282), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n288), .A2(G222), .ZN(new_n289));
  AOI21_X1  g0089(.A(new_n279), .B1(new_n287), .B2(new_n289), .ZN(new_n290));
  INV_X1    g0090(.A(G41), .ZN(new_n291));
  INV_X1    g0091(.A(G45), .ZN(new_n292));
  AOI21_X1  g0092(.A(G1), .B1(new_n291), .B2(new_n292), .ZN(new_n293));
  INV_X1    g0093(.A(KEYINPUT67), .ZN(new_n294));
  AOI21_X1  g0094(.A(new_n214), .B1(new_n294), .B2(new_n278), .ZN(new_n295));
  NAND3_X1  g0095(.A1(KEYINPUT67), .A2(G33), .A3(G41), .ZN(new_n296));
  AOI21_X1  g0096(.A(new_n293), .B1(new_n295), .B2(new_n296), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n297), .A2(G226), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n278), .A2(new_n294), .ZN(new_n299));
  NAND3_X1  g0099(.A1(new_n299), .A2(new_n277), .A3(new_n296), .ZN(new_n300));
  NAND3_X1  g0100(.A1(new_n300), .A2(G274), .A3(new_n293), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n298), .A2(new_n301), .ZN(new_n302));
  OR2_X1    g0102(.A1(new_n290), .A2(new_n302), .ZN(new_n303));
  AOI21_X1  g0103(.A(new_n275), .B1(new_n276), .B2(new_n303), .ZN(new_n304));
  NOR2_X1   g0104(.A1(new_n290), .A2(new_n302), .ZN(new_n305));
  XNOR2_X1  g0105(.A(KEYINPUT70), .B(G179), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n305), .A2(new_n306), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n304), .A2(new_n307), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n281), .A2(new_n282), .ZN(new_n309));
  NOR2_X1   g0109(.A1(G232), .A2(G1698), .ZN(new_n310));
  NOR2_X1   g0110(.A1(new_n280), .A2(G238), .ZN(new_n311));
  OAI21_X1  g0111(.A(new_n309), .B1(new_n310), .B2(new_n311), .ZN(new_n312));
  INV_X1    g0112(.A(new_n279), .ZN(new_n313));
  OAI211_X1 g0113(.A(new_n312), .B(new_n313), .C1(G107), .C2(new_n309), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n297), .A2(new_n217), .ZN(new_n315));
  NAND3_X1  g0115(.A1(new_n314), .A2(new_n301), .A3(new_n315), .ZN(new_n316));
  INV_X1    g0116(.A(G190), .ZN(new_n317));
  NOR2_X1   g0117(.A1(new_n316), .A2(new_n317), .ZN(new_n318));
  AND2_X1   g0118(.A1(new_n262), .A2(new_n272), .ZN(new_n319));
  XNOR2_X1  g0119(.A(KEYINPUT15), .B(G87), .ZN(new_n320));
  INV_X1    g0120(.A(G77), .ZN(new_n321));
  OAI22_X1  g0121(.A1(new_n320), .A2(new_n267), .B1(new_n206), .B2(new_n321), .ZN(new_n322));
  OAI21_X1  g0122(.A(new_n256), .B1(new_n319), .B2(new_n322), .ZN(new_n323));
  AOI21_X1  g0123(.A(new_n321), .B1(new_n205), .B2(G20), .ZN(new_n324));
  AOI22_X1  g0124(.A1(new_n250), .A2(new_n324), .B1(new_n321), .B2(new_n252), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n323), .A2(new_n325), .ZN(new_n326));
  NOR2_X1   g0126(.A1(new_n318), .A2(new_n326), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n316), .A2(G200), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n327), .A2(new_n328), .ZN(new_n329));
  XOR2_X1   g0129(.A(KEYINPUT70), .B(G179), .Z(new_n330));
  OR2_X1    g0130(.A1(new_n316), .A2(new_n330), .ZN(new_n331));
  AOI22_X1  g0131(.A1(new_n316), .A2(new_n276), .B1(new_n323), .B2(new_n325), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n331), .A2(new_n332), .ZN(new_n333));
  AND2_X1   g0133(.A1(new_n329), .A2(new_n333), .ZN(new_n334));
  INV_X1    g0134(.A(KEYINPUT9), .ZN(new_n335));
  OAI21_X1  g0135(.A(new_n335), .B1(new_n255), .B2(new_n274), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n305), .A2(G190), .ZN(new_n337));
  AND2_X1   g0137(.A1(new_n336), .A2(new_n337), .ZN(new_n338));
  AOI22_X1  g0138(.A1(new_n275), .A2(KEYINPUT9), .B1(new_n303), .B2(G200), .ZN(new_n339));
  INV_X1    g0139(.A(KEYINPUT10), .ZN(new_n340));
  NAND3_X1  g0140(.A1(new_n338), .A2(new_n339), .A3(new_n340), .ZN(new_n341));
  INV_X1    g0141(.A(new_n341), .ZN(new_n342));
  AOI21_X1  g0142(.A(new_n340), .B1(new_n338), .B2(new_n339), .ZN(new_n343));
  OAI211_X1 g0143(.A(new_n308), .B(new_n334), .C1(new_n342), .C2(new_n343), .ZN(new_n344));
  OAI22_X1  g0144(.A1(new_n267), .A2(new_n321), .B1(new_n206), .B2(G68), .ZN(new_n345));
  INV_X1    g0145(.A(KEYINPUT71), .ZN(new_n346));
  OR2_X1    g0146(.A1(new_n345), .A2(new_n346), .ZN(new_n347));
  AOI22_X1  g0147(.A1(new_n345), .A2(new_n346), .B1(G50), .B2(new_n272), .ZN(new_n348));
  AOI21_X1  g0148(.A(new_n257), .B1(new_n347), .B2(new_n348), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n349), .A2(KEYINPUT11), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n252), .A2(new_n270), .ZN(new_n351));
  XNOR2_X1  g0151(.A(new_n351), .B(KEYINPUT12), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n244), .A2(G68), .ZN(new_n353));
  OAI211_X1 g0153(.A(new_n350), .B(new_n352), .C1(new_n249), .C2(new_n353), .ZN(new_n354));
  NOR2_X1   g0154(.A1(new_n349), .A2(KEYINPUT11), .ZN(new_n355));
  NOR2_X1   g0155(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  INV_X1    g0156(.A(KEYINPUT72), .ZN(new_n357));
  INV_X1    g0157(.A(new_n293), .ZN(new_n358));
  NAND3_X1  g0158(.A1(new_n300), .A2(new_n358), .A3(G238), .ZN(new_n359));
  NOR2_X1   g0159(.A1(G226), .A2(G1698), .ZN(new_n360));
  AOI21_X1  g0160(.A(new_n360), .B1(new_n228), .B2(G1698), .ZN(new_n361));
  AOI22_X1  g0161(.A1(new_n361), .A2(new_n309), .B1(G33), .B2(G97), .ZN(new_n362));
  OAI211_X1 g0162(.A(new_n359), .B(new_n301), .C1(new_n362), .C2(new_n279), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n363), .A2(KEYINPUT13), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n228), .A2(G1698), .ZN(new_n365));
  OAI21_X1  g0165(.A(new_n365), .B1(G226), .B2(G1698), .ZN(new_n366));
  INV_X1    g0166(.A(G33), .ZN(new_n367));
  INV_X1    g0167(.A(G97), .ZN(new_n368));
  OAI22_X1  g0168(.A1(new_n366), .A2(new_n286), .B1(new_n367), .B2(new_n368), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n369), .A2(new_n313), .ZN(new_n370));
  INV_X1    g0170(.A(KEYINPUT13), .ZN(new_n371));
  NAND4_X1  g0171(.A1(new_n370), .A2(new_n371), .A3(new_n359), .A4(new_n301), .ZN(new_n372));
  AND2_X1   g0172(.A1(new_n364), .A2(new_n372), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n373), .A2(G179), .ZN(new_n374));
  AOI21_X1  g0174(.A(new_n276), .B1(new_n364), .B2(new_n372), .ZN(new_n375));
  INV_X1    g0175(.A(KEYINPUT14), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n375), .A2(new_n376), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n374), .A2(new_n377), .ZN(new_n378));
  NOR2_X1   g0178(.A1(new_n375), .A2(new_n376), .ZN(new_n379));
  OAI21_X1  g0179(.A(new_n357), .B1(new_n378), .B2(new_n379), .ZN(new_n380));
  INV_X1    g0180(.A(new_n379), .ZN(new_n381));
  NAND4_X1  g0181(.A1(new_n381), .A2(KEYINPUT72), .A3(new_n374), .A4(new_n377), .ZN(new_n382));
  AOI21_X1  g0182(.A(new_n356), .B1(new_n380), .B2(new_n382), .ZN(new_n383));
  INV_X1    g0183(.A(G200), .ZN(new_n384));
  OR2_X1    g0184(.A1(new_n373), .A2(new_n384), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n373), .A2(G190), .ZN(new_n386));
  NAND3_X1  g0186(.A1(new_n385), .A2(new_n356), .A3(new_n386), .ZN(new_n387));
  INV_X1    g0187(.A(new_n387), .ZN(new_n388));
  NAND3_X1  g0188(.A1(new_n263), .A2(new_n266), .A3(new_n244), .ZN(new_n389));
  AOI21_X1  g0189(.A(new_n249), .B1(new_n389), .B2(KEYINPUT75), .ZN(new_n390));
  INV_X1    g0190(.A(KEYINPUT75), .ZN(new_n391));
  NAND4_X1  g0191(.A1(new_n263), .A2(new_n266), .A3(new_n391), .A4(new_n244), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n263), .A2(new_n266), .ZN(new_n393));
  AOI22_X1  g0193(.A1(new_n390), .A2(new_n392), .B1(new_n252), .B2(new_n393), .ZN(new_n394));
  XNOR2_X1  g0194(.A(KEYINPUT73), .B(KEYINPUT16), .ZN(new_n395));
  INV_X1    g0195(.A(new_n395), .ZN(new_n396));
  NAND3_X1  g0196(.A1(new_n281), .A2(new_n206), .A3(new_n282), .ZN(new_n397));
  INV_X1    g0197(.A(KEYINPUT7), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n397), .A2(new_n398), .ZN(new_n399));
  INV_X1    g0199(.A(KEYINPUT74), .ZN(new_n400));
  NAND4_X1  g0200(.A1(new_n281), .A2(KEYINPUT7), .A3(new_n206), .A4(new_n282), .ZN(new_n401));
  NAND3_X1  g0201(.A1(new_n399), .A2(new_n400), .A3(new_n401), .ZN(new_n402));
  NOR4_X1   g0202(.A1(new_n284), .A2(new_n285), .A3(new_n398), .A4(G20), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n403), .A2(KEYINPUT74), .ZN(new_n404));
  NAND3_X1  g0204(.A1(new_n402), .A2(G68), .A3(new_n404), .ZN(new_n405));
  NOR2_X1   g0205(.A1(new_n258), .A2(new_n270), .ZN(new_n406));
  NOR2_X1   g0206(.A1(G58), .A2(G68), .ZN(new_n407));
  OAI21_X1  g0207(.A(G20), .B1(new_n406), .B2(new_n407), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n272), .A2(G159), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n408), .A2(new_n409), .ZN(new_n410));
  INV_X1    g0210(.A(new_n410), .ZN(new_n411));
  AOI21_X1  g0211(.A(new_n396), .B1(new_n405), .B2(new_n411), .ZN(new_n412));
  AOI21_X1  g0212(.A(KEYINPUT7), .B1(new_n286), .B2(new_n206), .ZN(new_n413));
  OAI21_X1  g0213(.A(G68), .B1(new_n413), .B2(new_n403), .ZN(new_n414));
  NAND3_X1  g0214(.A1(new_n414), .A2(KEYINPUT16), .A3(new_n411), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n415), .A2(new_n256), .ZN(new_n416));
  OAI21_X1  g0216(.A(new_n394), .B1(new_n412), .B2(new_n416), .ZN(new_n417));
  NAND3_X1  g0217(.A1(new_n300), .A2(new_n358), .A3(G232), .ZN(new_n418));
  NOR2_X1   g0218(.A1(G223), .A2(G1698), .ZN(new_n419));
  INV_X1    g0219(.A(G226), .ZN(new_n420));
  AOI21_X1  g0220(.A(new_n419), .B1(new_n420), .B2(G1698), .ZN(new_n421));
  AOI22_X1  g0221(.A1(new_n421), .A2(new_n309), .B1(G33), .B2(G87), .ZN(new_n422));
  OAI211_X1 g0222(.A(new_n301), .B(new_n418), .C1(new_n422), .C2(new_n279), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n423), .A2(G169), .ZN(new_n424));
  OAI21_X1  g0224(.A(new_n424), .B1(new_n306), .B2(new_n423), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n417), .A2(new_n425), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n426), .A2(KEYINPUT18), .ZN(new_n427));
  NAND2_X1  g0227(.A1(G33), .A2(G87), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n420), .A2(G1698), .ZN(new_n429));
  OAI21_X1  g0229(.A(new_n429), .B1(G223), .B2(G1698), .ZN(new_n430));
  OAI21_X1  g0230(.A(new_n428), .B1(new_n430), .B2(new_n286), .ZN(new_n431));
  INV_X1    g0231(.A(G274), .ZN(new_n432));
  AOI21_X1  g0232(.A(new_n432), .B1(new_n295), .B2(new_n296), .ZN(new_n433));
  AOI22_X1  g0233(.A1(new_n431), .A2(new_n313), .B1(new_n433), .B2(new_n293), .ZN(new_n434));
  INV_X1    g0234(.A(KEYINPUT76), .ZN(new_n435));
  NAND4_X1  g0235(.A1(new_n434), .A2(new_n435), .A3(new_n317), .A4(new_n418), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n431), .A2(new_n313), .ZN(new_n437));
  NAND4_X1  g0237(.A1(new_n437), .A2(new_n317), .A3(new_n301), .A4(new_n418), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n438), .A2(KEYINPUT76), .ZN(new_n439));
  AOI21_X1  g0239(.A(G200), .B1(new_n434), .B2(new_n418), .ZN(new_n440));
  OAI21_X1  g0240(.A(new_n436), .B1(new_n439), .B2(new_n440), .ZN(new_n441));
  INV_X1    g0241(.A(new_n441), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n389), .A2(KEYINPUT75), .ZN(new_n443));
  NAND3_X1  g0243(.A1(new_n443), .A2(new_n250), .A3(new_n392), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n393), .A2(new_n252), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n444), .A2(new_n445), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n405), .A2(new_n411), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n447), .A2(new_n395), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n399), .A2(new_n401), .ZN(new_n449));
  AOI21_X1  g0249(.A(new_n410), .B1(new_n449), .B2(G68), .ZN(new_n450));
  AOI21_X1  g0250(.A(new_n257), .B1(new_n450), .B2(KEYINPUT16), .ZN(new_n451));
  AOI21_X1  g0251(.A(new_n446), .B1(new_n448), .B2(new_n451), .ZN(new_n452));
  NAND3_X1  g0252(.A1(new_n442), .A2(new_n452), .A3(KEYINPUT17), .ZN(new_n453));
  INV_X1    g0253(.A(KEYINPUT18), .ZN(new_n454));
  NAND3_X1  g0254(.A1(new_n417), .A2(new_n425), .A3(new_n454), .ZN(new_n455));
  INV_X1    g0255(.A(KEYINPUT17), .ZN(new_n456));
  OAI21_X1  g0256(.A(new_n456), .B1(new_n417), .B2(new_n441), .ZN(new_n457));
  NAND4_X1  g0257(.A1(new_n427), .A2(new_n453), .A3(new_n455), .A4(new_n457), .ZN(new_n458));
  NOR4_X1   g0258(.A1(new_n344), .A2(new_n383), .A3(new_n388), .A4(new_n458), .ZN(new_n459));
  INV_X1    g0259(.A(KEYINPUT79), .ZN(new_n460));
  OAI211_X1 g0260(.A(G244), .B(new_n280), .C1(new_n284), .C2(new_n285), .ZN(new_n461));
  INV_X1    g0261(.A(KEYINPUT78), .ZN(new_n462));
  NOR2_X1   g0262(.A1(new_n462), .A2(KEYINPUT4), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n461), .A2(new_n463), .ZN(new_n464));
  NAND2_X1  g0264(.A1(G33), .A2(G283), .ZN(new_n465));
  NAND3_X1  g0265(.A1(new_n309), .A2(G250), .A3(G1698), .ZN(new_n466));
  NAND3_X1  g0266(.A1(new_n464), .A2(new_n465), .A3(new_n466), .ZN(new_n467));
  INV_X1    g0267(.A(KEYINPUT4), .ZN(new_n468));
  AOI21_X1  g0268(.A(new_n468), .B1(new_n461), .B2(KEYINPUT78), .ZN(new_n469));
  OAI21_X1  g0269(.A(new_n313), .B1(new_n467), .B2(new_n469), .ZN(new_n470));
  XNOR2_X1  g0270(.A(KEYINPUT5), .B(G41), .ZN(new_n471));
  NOR2_X1   g0271(.A1(new_n292), .A2(G1), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  NAND3_X1  g0273(.A1(new_n473), .A2(G257), .A3(new_n300), .ZN(new_n474));
  NAND4_X1  g0274(.A1(new_n300), .A2(G274), .A3(new_n472), .A4(new_n471), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  INV_X1    g0276(.A(new_n476), .ZN(new_n477));
  NAND3_X1  g0277(.A1(new_n470), .A2(new_n306), .A3(new_n477), .ZN(new_n478));
  AOI22_X1  g0278(.A1(new_n283), .A2(G250), .B1(G33), .B2(G283), .ZN(new_n479));
  AOI21_X1  g0279(.A(new_n462), .B1(new_n288), .B2(G244), .ZN(new_n480));
  OAI211_X1 g0280(.A(new_n479), .B(new_n464), .C1(new_n480), .C2(new_n468), .ZN(new_n481));
  AOI21_X1  g0281(.A(new_n476), .B1(new_n481), .B2(new_n313), .ZN(new_n482));
  OAI21_X1  g0282(.A(new_n478), .B1(new_n482), .B2(G169), .ZN(new_n483));
  NOR2_X1   g0283(.A1(new_n247), .A2(G97), .ZN(new_n484));
  INV_X1    g0284(.A(KEYINPUT77), .ZN(new_n485));
  OAI21_X1  g0285(.A(new_n485), .B1(new_n367), .B2(G1), .ZN(new_n486));
  NAND3_X1  g0286(.A1(new_n205), .A2(KEYINPUT77), .A3(G33), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n486), .A2(new_n487), .ZN(new_n488));
  NOR2_X1   g0288(.A1(new_n249), .A2(new_n488), .ZN(new_n489));
  AOI21_X1  g0289(.A(new_n484), .B1(new_n489), .B2(G97), .ZN(new_n490));
  INV_X1    g0290(.A(new_n490), .ZN(new_n491));
  NAND3_X1  g0291(.A1(new_n402), .A2(G107), .A3(new_n404), .ZN(new_n492));
  INV_X1    g0292(.A(G107), .ZN(new_n493));
  NAND3_X1  g0293(.A1(new_n493), .A2(KEYINPUT6), .A3(G97), .ZN(new_n494));
  NOR2_X1   g0294(.A1(new_n368), .A2(new_n493), .ZN(new_n495));
  NOR2_X1   g0295(.A1(G97), .A2(G107), .ZN(new_n496));
  NOR2_X1   g0296(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  OAI21_X1  g0297(.A(new_n494), .B1(new_n497), .B2(KEYINPUT6), .ZN(new_n498));
  AOI22_X1  g0298(.A1(new_n498), .A2(G20), .B1(G77), .B2(new_n272), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n492), .A2(new_n499), .ZN(new_n500));
  AOI21_X1  g0300(.A(new_n491), .B1(new_n500), .B2(new_n256), .ZN(new_n501));
  OAI21_X1  g0301(.A(new_n460), .B1(new_n483), .B2(new_n501), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n500), .A2(new_n256), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n503), .A2(new_n490), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n470), .A2(new_n477), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n505), .A2(new_n276), .ZN(new_n506));
  NAND4_X1  g0306(.A1(new_n504), .A2(KEYINPUT79), .A3(new_n478), .A4(new_n506), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n505), .A2(G200), .ZN(new_n508));
  OAI211_X1 g0308(.A(new_n508), .B(new_n501), .C1(new_n317), .C2(new_n505), .ZN(new_n509));
  AND3_X1   g0309(.A1(new_n502), .A2(new_n507), .A3(new_n509), .ZN(new_n510));
  OAI211_X1 g0310(.A(G257), .B(G1698), .C1(new_n284), .C2(new_n285), .ZN(new_n511));
  OAI211_X1 g0311(.A(G250), .B(new_n280), .C1(new_n284), .C2(new_n285), .ZN(new_n512));
  NAND2_X1  g0312(.A1(G33), .A2(G294), .ZN(new_n513));
  NAND3_X1  g0313(.A1(new_n511), .A2(new_n512), .A3(new_n513), .ZN(new_n514));
  AOI22_X1  g0314(.A1(new_n296), .A2(new_n295), .B1(new_n471), .B2(new_n472), .ZN(new_n515));
  AOI22_X1  g0315(.A1(new_n313), .A2(new_n514), .B1(new_n515), .B2(G264), .ZN(new_n516));
  INV_X1    g0316(.A(KEYINPUT83), .ZN(new_n517));
  NAND3_X1  g0317(.A1(new_n516), .A2(new_n517), .A3(new_n475), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n514), .A2(new_n313), .ZN(new_n519));
  NAND3_X1  g0319(.A1(new_n473), .A2(G264), .A3(new_n300), .ZN(new_n520));
  NAND3_X1  g0320(.A1(new_n519), .A2(new_n475), .A3(new_n520), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n521), .A2(KEYINPUT83), .ZN(new_n522));
  NAND3_X1  g0322(.A1(new_n518), .A2(new_n522), .A3(G169), .ZN(new_n523));
  NAND3_X1  g0323(.A1(new_n516), .A2(G179), .A3(new_n475), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  OAI21_X1  g0325(.A(KEYINPUT82), .B1(new_n206), .B2(G107), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n526), .A2(KEYINPUT23), .ZN(new_n527));
  INV_X1    g0327(.A(KEYINPUT23), .ZN(new_n528));
  OAI211_X1 g0328(.A(KEYINPUT82), .B(new_n528), .C1(new_n206), .C2(G107), .ZN(new_n529));
  AOI22_X1  g0329(.A1(new_n527), .A2(new_n529), .B1(G116), .B2(new_n268), .ZN(new_n530));
  AND2_X1   g0330(.A1(KEYINPUT81), .A2(KEYINPUT22), .ZN(new_n531));
  NAND4_X1  g0331(.A1(new_n309), .A2(new_n206), .A3(G87), .A4(new_n531), .ZN(new_n532));
  OAI211_X1 g0332(.A(new_n206), .B(G87), .C1(new_n284), .C2(new_n285), .ZN(new_n533));
  NOR2_X1   g0333(.A1(KEYINPUT81), .A2(KEYINPUT22), .ZN(new_n534));
  NOR2_X1   g0334(.A1(new_n531), .A2(new_n534), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n533), .A2(new_n535), .ZN(new_n536));
  NAND3_X1  g0336(.A1(new_n530), .A2(new_n532), .A3(new_n536), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n537), .A2(KEYINPUT24), .ZN(new_n538));
  INV_X1    g0338(.A(KEYINPUT24), .ZN(new_n539));
  NAND4_X1  g0339(.A1(new_n530), .A2(new_n532), .A3(new_n539), .A4(new_n536), .ZN(new_n540));
  AOI21_X1  g0340(.A(new_n257), .B1(new_n538), .B2(new_n540), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n489), .A2(G107), .ZN(new_n542));
  AOI21_X1  g0342(.A(KEYINPUT25), .B1(new_n252), .B2(new_n493), .ZN(new_n543));
  INV_X1    g0343(.A(KEYINPUT25), .ZN(new_n544));
  NOR3_X1   g0344(.A1(new_n247), .A2(new_n544), .A3(G107), .ZN(new_n545));
  OAI21_X1  g0345(.A(new_n542), .B1(new_n543), .B2(new_n545), .ZN(new_n546));
  OR2_X1    g0346(.A1(new_n541), .A2(new_n546), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n525), .A2(new_n547), .ZN(new_n548));
  NOR2_X1   g0348(.A1(new_n541), .A2(new_n546), .ZN(new_n549));
  AOI21_X1  g0349(.A(G190), .B1(new_n518), .B2(new_n522), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n521), .A2(new_n384), .ZN(new_n551));
  INV_X1    g0351(.A(new_n551), .ZN(new_n552));
  OAI21_X1  g0352(.A(new_n549), .B1(new_n550), .B2(new_n552), .ZN(new_n553));
  AND2_X1   g0353(.A1(new_n548), .A2(new_n553), .ZN(new_n554));
  OAI211_X1 g0354(.A(G264), .B(G1698), .C1(new_n284), .C2(new_n285), .ZN(new_n555));
  OAI211_X1 g0355(.A(G257), .B(new_n280), .C1(new_n284), .C2(new_n285), .ZN(new_n556));
  INV_X1    g0356(.A(G303), .ZN(new_n557));
  OAI211_X1 g0357(.A(new_n555), .B(new_n556), .C1(new_n557), .C2(new_n309), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n558), .A2(new_n313), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n515), .A2(G270), .ZN(new_n560));
  NAND3_X1  g0360(.A1(new_n559), .A2(new_n475), .A3(new_n560), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n489), .A2(G116), .ZN(new_n562));
  INV_X1    g0362(.A(G116), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n252), .A2(new_n563), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n563), .A2(G20), .ZN(new_n565));
  AND2_X1   g0365(.A1(new_n256), .A2(new_n565), .ZN(new_n566));
  OAI211_X1 g0366(.A(new_n465), .B(new_n206), .C1(G33), .C2(new_n368), .ZN(new_n567));
  AOI21_X1  g0367(.A(KEYINPUT20), .B1(new_n566), .B2(new_n567), .ZN(new_n568));
  AND4_X1   g0368(.A1(KEYINPUT20), .A2(new_n567), .A3(new_n256), .A4(new_n565), .ZN(new_n569));
  OAI211_X1 g0369(.A(new_n562), .B(new_n564), .C1(new_n568), .C2(new_n569), .ZN(new_n570));
  NAND3_X1  g0370(.A1(new_n561), .A2(new_n570), .A3(G169), .ZN(new_n571));
  INV_X1    g0371(.A(KEYINPUT21), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  INV_X1    g0373(.A(G179), .ZN(new_n574));
  NOR2_X1   g0374(.A1(new_n561), .A2(new_n574), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n575), .A2(new_n570), .ZN(new_n576));
  NAND4_X1  g0376(.A1(new_n561), .A2(new_n570), .A3(KEYINPUT21), .A4(G169), .ZN(new_n577));
  NAND3_X1  g0377(.A1(new_n573), .A2(new_n576), .A3(new_n577), .ZN(new_n578));
  INV_X1    g0378(.A(new_n578), .ZN(new_n579));
  AOI21_X1  g0379(.A(new_n570), .B1(G200), .B2(new_n561), .ZN(new_n580));
  OAI21_X1  g0380(.A(new_n580), .B1(new_n317), .B2(new_n561), .ZN(new_n581));
  OAI211_X1 g0381(.A(G244), .B(G1698), .C1(new_n284), .C2(new_n285), .ZN(new_n582));
  OAI211_X1 g0382(.A(G238), .B(new_n280), .C1(new_n284), .C2(new_n285), .ZN(new_n583));
  NAND2_X1  g0383(.A1(G33), .A2(G116), .ZN(new_n584));
  NAND3_X1  g0384(.A1(new_n582), .A2(new_n583), .A3(new_n584), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n585), .A2(new_n313), .ZN(new_n586));
  AOI21_X1  g0386(.A(G250), .B1(new_n205), .B2(G45), .ZN(new_n587));
  AOI21_X1  g0387(.A(new_n587), .B1(new_n432), .B2(new_n472), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n588), .A2(new_n300), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n586), .A2(new_n589), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n590), .A2(new_n276), .ZN(new_n591));
  NAND3_X1  g0391(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n592));
  INV_X1    g0392(.A(KEYINPUT80), .ZN(new_n593));
  AND3_X1   g0393(.A1(new_n592), .A2(new_n593), .A3(new_n206), .ZN(new_n594));
  AOI21_X1  g0394(.A(new_n593), .B1(new_n592), .B2(new_n206), .ZN(new_n595));
  NOR3_X1   g0395(.A1(G87), .A2(G97), .A3(G107), .ZN(new_n596));
  NOR3_X1   g0396(.A1(new_n594), .A2(new_n595), .A3(new_n596), .ZN(new_n597));
  OAI211_X1 g0397(.A(new_n206), .B(G68), .C1(new_n284), .C2(new_n285), .ZN(new_n598));
  NOR2_X1   g0398(.A1(new_n267), .A2(new_n368), .ZN(new_n599));
  OAI21_X1  g0399(.A(new_n598), .B1(KEYINPUT19), .B2(new_n599), .ZN(new_n600));
  OAI21_X1  g0400(.A(new_n256), .B1(new_n597), .B2(new_n600), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n320), .A2(new_n252), .ZN(new_n602));
  INV_X1    g0402(.A(new_n320), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n489), .A2(new_n603), .ZN(new_n604));
  NAND3_X1  g0404(.A1(new_n601), .A2(new_n602), .A3(new_n604), .ZN(new_n605));
  AOI22_X1  g0405(.A1(new_n585), .A2(new_n313), .B1(new_n300), .B2(new_n588), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n606), .A2(new_n306), .ZN(new_n607));
  NAND3_X1  g0407(.A1(new_n591), .A2(new_n605), .A3(new_n607), .ZN(new_n608));
  NOR2_X1   g0408(.A1(new_n606), .A2(new_n384), .ZN(new_n609));
  NAND3_X1  g0409(.A1(new_n586), .A2(G190), .A3(new_n589), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n489), .A2(G87), .ZN(new_n611));
  NAND4_X1  g0411(.A1(new_n610), .A2(new_n602), .A3(new_n601), .A4(new_n611), .ZN(new_n612));
  OAI21_X1  g0412(.A(new_n608), .B1(new_n609), .B2(new_n612), .ZN(new_n613));
  INV_X1    g0413(.A(new_n613), .ZN(new_n614));
  AND3_X1   g0414(.A1(new_n579), .A2(new_n581), .A3(new_n614), .ZN(new_n615));
  AND4_X1   g0415(.A1(new_n459), .A2(new_n510), .A3(new_n554), .A4(new_n615), .ZN(G372));
  NAND2_X1  g0416(.A1(new_n453), .A2(new_n457), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n380), .A2(new_n382), .ZN(new_n618));
  INV_X1    g0418(.A(new_n356), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  AND2_X1   g0420(.A1(new_n331), .A2(new_n332), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n387), .A2(new_n621), .ZN(new_n622));
  AOI21_X1  g0422(.A(new_n617), .B1(new_n620), .B2(new_n622), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n427), .A2(new_n455), .ZN(new_n624));
  NOR2_X1   g0424(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n625), .A2(KEYINPUT85), .ZN(new_n626));
  INV_X1    g0426(.A(new_n343), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n627), .A2(new_n341), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n626), .A2(new_n628), .ZN(new_n629));
  NOR2_X1   g0429(.A1(new_n625), .A2(KEYINPUT85), .ZN(new_n630));
  OAI21_X1  g0430(.A(new_n308), .B1(new_n629), .B2(new_n630), .ZN(new_n631));
  INV_X1    g0431(.A(new_n631), .ZN(new_n632));
  AOI21_X1  g0432(.A(new_n613), .B1(new_n502), .B2(new_n507), .ZN(new_n633));
  INV_X1    g0433(.A(KEYINPUT26), .ZN(new_n634));
  NOR2_X1   g0434(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  AND3_X1   g0435(.A1(new_n470), .A2(new_n306), .A3(new_n477), .ZN(new_n636));
  AOI21_X1  g0436(.A(G169), .B1(new_n470), .B2(new_n477), .ZN(new_n637));
  NOR2_X1   g0437(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  AND3_X1   g0438(.A1(new_n601), .A2(new_n602), .A3(new_n611), .ZN(new_n639));
  INV_X1    g0439(.A(KEYINPUT84), .ZN(new_n640));
  NAND3_X1  g0440(.A1(new_n590), .A2(new_n640), .A3(G200), .ZN(new_n641));
  OAI21_X1  g0441(.A(KEYINPUT84), .B1(new_n606), .B2(new_n384), .ZN(new_n642));
  NAND4_X1  g0442(.A1(new_n639), .A2(new_n641), .A3(new_n642), .A4(new_n610), .ZN(new_n643));
  NAND4_X1  g0443(.A1(new_n638), .A2(new_n504), .A3(new_n608), .A4(new_n643), .ZN(new_n644));
  OAI21_X1  g0444(.A(new_n608), .B1(new_n644), .B2(KEYINPUT26), .ZN(new_n645));
  NOR2_X1   g0445(.A1(new_n635), .A2(new_n645), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n579), .A2(new_n548), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n641), .A2(new_n642), .ZN(new_n648));
  OAI21_X1  g0448(.A(new_n608), .B1(new_n648), .B2(new_n612), .ZN(new_n649));
  AOI21_X1  g0449(.A(new_n517), .B1(new_n516), .B2(new_n475), .ZN(new_n650));
  AND4_X1   g0450(.A1(new_n517), .A2(new_n519), .A3(new_n475), .A4(new_n520), .ZN(new_n651));
  OAI21_X1  g0451(.A(new_n317), .B1(new_n650), .B2(new_n651), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n652), .A2(new_n551), .ZN(new_n653));
  AOI21_X1  g0453(.A(new_n649), .B1(new_n653), .B2(new_n549), .ZN(new_n654));
  NAND3_X1  g0454(.A1(new_n510), .A2(new_n647), .A3(new_n654), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n646), .A2(new_n655), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n459), .A2(new_n656), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n632), .A2(new_n657), .ZN(G369));
  NAND3_X1  g0458(.A1(new_n205), .A2(new_n206), .A3(G13), .ZN(new_n659));
  AND3_X1   g0459(.A1(new_n659), .A2(KEYINPUT86), .A3(KEYINPUT27), .ZN(new_n660));
  AOI21_X1  g0460(.A(KEYINPUT86), .B1(new_n659), .B2(KEYINPUT27), .ZN(new_n661));
  OAI221_X1 g0461(.A(G213), .B1(KEYINPUT27), .B2(new_n659), .C1(new_n660), .C2(new_n661), .ZN(new_n662));
  INV_X1    g0462(.A(G343), .ZN(new_n663));
  NOR2_X1   g0463(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n664), .A2(new_n570), .ZN(new_n665));
  NAND3_X1  g0465(.A1(new_n579), .A2(new_n581), .A3(new_n665), .ZN(new_n666));
  NAND3_X1  g0466(.A1(new_n578), .A2(new_n570), .A3(new_n664), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n668), .A2(G330), .ZN(new_n669));
  INV_X1    g0469(.A(new_n669), .ZN(new_n670));
  INV_X1    g0470(.A(new_n664), .ZN(new_n671));
  OAI21_X1  g0471(.A(new_n554), .B1(new_n549), .B2(new_n671), .ZN(new_n672));
  NAND3_X1  g0472(.A1(new_n525), .A2(new_n547), .A3(new_n664), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n670), .A2(new_n674), .ZN(new_n675));
  NOR2_X1   g0475(.A1(new_n579), .A2(new_n664), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n554), .A2(new_n676), .ZN(new_n677));
  NAND3_X1  g0477(.A1(new_n525), .A2(new_n547), .A3(new_n671), .ZN(new_n678));
  AND2_X1   g0478(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n675), .A2(new_n679), .ZN(G399));
  INV_X1    g0480(.A(new_n209), .ZN(new_n681));
  NOR2_X1   g0481(.A1(new_n681), .A2(G41), .ZN(new_n682));
  INV_X1    g0482(.A(new_n682), .ZN(new_n683));
  AND2_X1   g0483(.A1(new_n596), .A2(new_n563), .ZN(new_n684));
  NAND3_X1  g0484(.A1(new_n683), .A2(G1), .A3(new_n684), .ZN(new_n685));
  OAI21_X1  g0485(.A(new_n685), .B1(new_n212), .B2(new_n683), .ZN(new_n686));
  XNOR2_X1  g0486(.A(new_n686), .B(KEYINPUT28), .ZN(new_n687));
  NAND4_X1  g0487(.A1(new_n615), .A2(new_n510), .A3(new_n554), .A4(new_n671), .ZN(new_n688));
  NAND4_X1  g0488(.A1(new_n575), .A2(new_n482), .A3(new_n516), .A4(new_n606), .ZN(new_n689));
  INV_X1    g0489(.A(KEYINPUT30), .ZN(new_n690));
  NOR2_X1   g0490(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n516), .A2(new_n606), .ZN(new_n692));
  NOR3_X1   g0492(.A1(new_n692), .A2(new_n561), .A3(new_n574), .ZN(new_n693));
  AOI21_X1  g0493(.A(KEYINPUT30), .B1(new_n693), .B2(new_n482), .ZN(new_n694));
  NOR2_X1   g0494(.A1(new_n691), .A2(new_n694), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n505), .A2(new_n521), .ZN(new_n696));
  NAND3_X1  g0496(.A1(new_n561), .A2(new_n306), .A3(new_n590), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n697), .A2(KEYINPUT87), .ZN(new_n698));
  INV_X1    g0498(.A(KEYINPUT87), .ZN(new_n699));
  NAND4_X1  g0499(.A1(new_n561), .A2(new_n699), .A3(new_n306), .A4(new_n590), .ZN(new_n700));
  AOI21_X1  g0500(.A(new_n696), .B1(new_n698), .B2(new_n700), .ZN(new_n701));
  INV_X1    g0501(.A(new_n701), .ZN(new_n702));
  AOI21_X1  g0502(.A(new_n671), .B1(new_n695), .B2(new_n702), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n703), .A2(KEYINPUT31), .ZN(new_n704));
  INV_X1    g0504(.A(KEYINPUT31), .ZN(new_n705));
  NOR3_X1   g0505(.A1(new_n691), .A2(new_n701), .A3(new_n694), .ZN(new_n706));
  OAI21_X1  g0506(.A(new_n705), .B1(new_n706), .B2(new_n671), .ZN(new_n707));
  NAND3_X1  g0507(.A1(new_n688), .A2(new_n704), .A3(new_n707), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n708), .A2(G330), .ZN(new_n709));
  INV_X1    g0509(.A(new_n709), .ZN(new_n710));
  INV_X1    g0510(.A(KEYINPUT89), .ZN(new_n711));
  NAND4_X1  g0511(.A1(new_n654), .A2(new_n502), .A3(new_n507), .A4(new_n509), .ZN(new_n712));
  AOI21_X1  g0512(.A(new_n578), .B1(new_n525), .B2(new_n547), .ZN(new_n713));
  OAI21_X1  g0513(.A(new_n711), .B1(new_n712), .B2(new_n713), .ZN(new_n714));
  NAND4_X1  g0514(.A1(new_n510), .A2(KEYINPUT89), .A3(new_n647), .A4(new_n654), .ZN(new_n715));
  AOI21_X1  g0515(.A(KEYINPUT79), .B1(new_n638), .B2(new_n504), .ZN(new_n716));
  NOR3_X1   g0516(.A1(new_n483), .A2(new_n460), .A3(new_n501), .ZN(new_n717));
  OAI211_X1 g0517(.A(new_n634), .B(new_n614), .C1(new_n716), .C2(new_n717), .ZN(new_n718));
  INV_X1    g0518(.A(new_n608), .ZN(new_n719));
  AOI21_X1  g0519(.A(new_n719), .B1(new_n644), .B2(KEYINPUT26), .ZN(new_n720));
  AND2_X1   g0520(.A1(new_n718), .A2(new_n720), .ZN(new_n721));
  NAND3_X1  g0521(.A1(new_n714), .A2(new_n715), .A3(new_n721), .ZN(new_n722));
  NAND3_X1  g0522(.A1(new_n722), .A2(KEYINPUT29), .A3(new_n671), .ZN(new_n723));
  INV_X1    g0523(.A(KEYINPUT90), .ZN(new_n724));
  NAND2_X1  g0524(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  NAND4_X1  g0525(.A1(new_n722), .A2(KEYINPUT90), .A3(KEYINPUT29), .A4(new_n671), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  AOI21_X1  g0527(.A(new_n664), .B1(new_n646), .B2(new_n655), .ZN(new_n728));
  INV_X1    g0528(.A(new_n728), .ZN(new_n729));
  XOR2_X1   g0529(.A(KEYINPUT88), .B(KEYINPUT29), .Z(new_n730));
  INV_X1    g0530(.A(new_n730), .ZN(new_n731));
  NAND2_X1  g0531(.A1(new_n729), .A2(new_n731), .ZN(new_n732));
  AOI21_X1  g0532(.A(new_n710), .B1(new_n727), .B2(new_n732), .ZN(new_n733));
  OAI21_X1  g0533(.A(new_n687), .B1(new_n733), .B2(G1), .ZN(G364));
  AND2_X1   g0534(.A1(new_n206), .A2(G13), .ZN(new_n735));
  AOI21_X1  g0535(.A(new_n205), .B1(new_n735), .B2(G45), .ZN(new_n736));
  INV_X1    g0536(.A(new_n736), .ZN(new_n737));
  NOR2_X1   g0537(.A1(new_n682), .A2(new_n737), .ZN(new_n738));
  NOR2_X1   g0538(.A1(new_n670), .A2(new_n738), .ZN(new_n739));
  OAI21_X1  g0539(.A(new_n739), .B1(G330), .B2(new_n668), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n209), .A2(new_n309), .ZN(new_n741));
  OAI22_X1  g0541(.A1(new_n741), .A2(new_n203), .B1(G116), .B2(new_n209), .ZN(new_n742));
  NAND2_X1  g0542(.A1(new_n209), .A2(new_n286), .ZN(new_n743));
  XOR2_X1   g0543(.A(new_n743), .B(KEYINPUT91), .Z(new_n744));
  INV_X1    g0544(.A(new_n744), .ZN(new_n745));
  AOI21_X1  g0545(.A(new_n745), .B1(new_n292), .B2(new_n213), .ZN(new_n746));
  NAND2_X1  g0546(.A1(new_n239), .A2(G45), .ZN(new_n747));
  AOI21_X1  g0547(.A(new_n742), .B1(new_n746), .B2(new_n747), .ZN(new_n748));
  NOR2_X1   g0548(.A1(G13), .A2(G33), .ZN(new_n749));
  INV_X1    g0549(.A(new_n749), .ZN(new_n750));
  NOR2_X1   g0550(.A1(new_n750), .A2(G20), .ZN(new_n751));
  XNOR2_X1  g0551(.A(new_n751), .B(KEYINPUT92), .ZN(new_n752));
  INV_X1    g0552(.A(new_n752), .ZN(new_n753));
  AOI21_X1  g0553(.A(new_n214), .B1(G20), .B2(new_n276), .ZN(new_n754));
  NOR2_X1   g0554(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  INV_X1    g0555(.A(new_n755), .ZN(new_n756));
  OAI21_X1  g0556(.A(new_n738), .B1(new_n748), .B2(new_n756), .ZN(new_n757));
  NOR2_X1   g0557(.A1(new_n206), .A2(G190), .ZN(new_n758));
  NOR2_X1   g0558(.A1(G179), .A2(G200), .ZN(new_n759));
  NAND2_X1  g0559(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  INV_X1    g0560(.A(new_n760), .ZN(new_n761));
  AOI21_X1  g0561(.A(new_n309), .B1(new_n761), .B2(G329), .ZN(new_n762));
  NOR2_X1   g0562(.A1(new_n206), .A2(new_n317), .ZN(new_n763));
  NAND3_X1  g0563(.A1(new_n763), .A2(new_n574), .A3(G200), .ZN(new_n764));
  OAI21_X1  g0564(.A(new_n762), .B1(new_n557), .B2(new_n764), .ZN(new_n765));
  AOI21_X1  g0565(.A(new_n206), .B1(new_n759), .B2(G190), .ZN(new_n766));
  INV_X1    g0566(.A(new_n766), .ZN(new_n767));
  AOI21_X1  g0567(.A(new_n765), .B1(G294), .B2(new_n767), .ZN(new_n768));
  NAND3_X1  g0568(.A1(new_n758), .A2(new_n574), .A3(G200), .ZN(new_n769));
  INV_X1    g0569(.A(KEYINPUT94), .ZN(new_n770));
  OR2_X1    g0570(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  NAND2_X1  g0571(.A1(new_n769), .A2(new_n770), .ZN(new_n772));
  AND2_X1   g0572(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  NAND3_X1  g0573(.A1(new_n330), .A2(new_n384), .A3(new_n758), .ZN(new_n774));
  INV_X1    g0574(.A(new_n774), .ZN(new_n775));
  AOI22_X1  g0575(.A1(new_n773), .A2(G283), .B1(G311), .B2(new_n775), .ZN(new_n776));
  NOR2_X1   g0576(.A1(new_n206), .A2(new_n384), .ZN(new_n777));
  NAND3_X1  g0577(.A1(new_n330), .A2(new_n317), .A3(new_n777), .ZN(new_n778));
  INV_X1    g0578(.A(KEYINPUT95), .ZN(new_n779));
  XNOR2_X1  g0579(.A(new_n778), .B(new_n779), .ZN(new_n780));
  XNOR2_X1  g0580(.A(KEYINPUT33), .B(G317), .ZN(new_n781));
  NAND2_X1  g0581(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  NOR3_X1   g0582(.A1(new_n306), .A2(new_n206), .A3(new_n384), .ZN(new_n783));
  AND2_X1   g0583(.A1(new_n783), .A2(G190), .ZN(new_n784));
  NAND3_X1  g0584(.A1(new_n330), .A2(new_n384), .A3(new_n763), .ZN(new_n785));
  INV_X1    g0585(.A(new_n785), .ZN(new_n786));
  AOI22_X1  g0586(.A1(new_n784), .A2(G326), .B1(new_n786), .B2(G322), .ZN(new_n787));
  NAND4_X1  g0587(.A1(new_n768), .A2(new_n776), .A3(new_n782), .A4(new_n787), .ZN(new_n788));
  NOR2_X1   g0588(.A1(new_n766), .A2(new_n368), .ZN(new_n789));
  INV_X1    g0589(.A(new_n764), .ZN(new_n790));
  NAND2_X1  g0590(.A1(new_n790), .A2(G87), .ZN(new_n791));
  INV_X1    g0591(.A(KEYINPUT32), .ZN(new_n792));
  INV_X1    g0592(.A(G159), .ZN(new_n793));
  NOR2_X1   g0593(.A1(new_n760), .A2(new_n793), .ZN(new_n794));
  OAI211_X1 g0594(.A(new_n791), .B(new_n309), .C1(new_n792), .C2(new_n794), .ZN(new_n795));
  AOI211_X1 g0595(.A(new_n789), .B(new_n795), .C1(new_n792), .C2(new_n794), .ZN(new_n796));
  NAND2_X1  g0596(.A1(new_n773), .A2(G107), .ZN(new_n797));
  XNOR2_X1  g0597(.A(new_n778), .B(KEYINPUT95), .ZN(new_n798));
  OAI211_X1 g0598(.A(new_n796), .B(new_n797), .C1(new_n270), .C2(new_n798), .ZN(new_n799));
  AOI22_X1  g0599(.A1(new_n786), .A2(G58), .B1(new_n775), .B2(G77), .ZN(new_n800));
  NAND2_X1  g0600(.A1(new_n783), .A2(G190), .ZN(new_n801));
  OAI21_X1  g0601(.A(new_n800), .B1(new_n253), .B2(new_n801), .ZN(new_n802));
  XNOR2_X1  g0602(.A(new_n802), .B(KEYINPUT93), .ZN(new_n803));
  OAI21_X1  g0603(.A(new_n788), .B1(new_n799), .B2(new_n803), .ZN(new_n804));
  AOI21_X1  g0604(.A(new_n757), .B1(new_n804), .B2(new_n754), .ZN(new_n805));
  OAI21_X1  g0605(.A(new_n805), .B1(new_n668), .B2(new_n752), .ZN(new_n806));
  AND2_X1   g0606(.A1(new_n740), .A2(new_n806), .ZN(new_n807));
  INV_X1    g0607(.A(new_n807), .ZN(G396));
  INV_X1    g0608(.A(KEYINPUT99), .ZN(new_n809));
  NAND2_X1  g0609(.A1(new_n621), .A2(new_n809), .ZN(new_n810));
  NAND2_X1  g0610(.A1(new_n333), .A2(KEYINPUT99), .ZN(new_n811));
  NAND2_X1  g0611(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  AOI21_X1  g0612(.A(new_n812), .B1(new_n328), .B2(new_n327), .ZN(new_n813));
  NOR3_X1   g0613(.A1(new_n649), .A2(new_n501), .A3(new_n483), .ZN(new_n814));
  NAND2_X1  g0614(.A1(new_n814), .A2(new_n634), .ZN(new_n815));
  OAI211_X1 g0615(.A(new_n815), .B(new_n608), .C1(new_n634), .C2(new_n633), .ZN(new_n816));
  NAND3_X1  g0616(.A1(new_n502), .A2(new_n507), .A3(new_n509), .ZN(new_n817));
  NAND3_X1  g0617(.A1(new_n553), .A2(new_n608), .A3(new_n643), .ZN(new_n818));
  NOR3_X1   g0618(.A1(new_n713), .A2(new_n817), .A3(new_n818), .ZN(new_n819));
  OAI211_X1 g0619(.A(new_n671), .B(new_n813), .C1(new_n816), .C2(new_n819), .ZN(new_n820));
  NAND2_X1  g0620(.A1(new_n664), .A2(new_n326), .ZN(new_n821));
  NAND4_X1  g0621(.A1(new_n810), .A2(new_n329), .A3(new_n821), .A4(new_n811), .ZN(new_n822));
  OAI21_X1  g0622(.A(new_n822), .B1(new_n333), .B2(new_n671), .ZN(new_n823));
  OAI21_X1  g0623(.A(new_n820), .B1(new_n728), .B2(new_n823), .ZN(new_n824));
  NOR2_X1   g0624(.A1(new_n824), .A2(new_n709), .ZN(new_n825));
  XOR2_X1   g0625(.A(new_n825), .B(KEYINPUT100), .Z(new_n826));
  AOI21_X1  g0626(.A(new_n738), .B1(new_n824), .B2(new_n709), .ZN(new_n827));
  NAND2_X1  g0627(.A1(new_n826), .A2(new_n827), .ZN(new_n828));
  NOR2_X1   g0628(.A1(new_n754), .A2(new_n749), .ZN(new_n829));
  INV_X1    g0629(.A(new_n829), .ZN(new_n830));
  NAND2_X1  g0630(.A1(new_n773), .A2(G87), .ZN(new_n831));
  INV_X1    g0631(.A(G311), .ZN(new_n832));
  OAI21_X1  g0632(.A(new_n831), .B1(new_n832), .B2(new_n760), .ZN(new_n833));
  XNOR2_X1  g0633(.A(new_n833), .B(KEYINPUT97), .ZN(new_n834));
  AOI211_X1 g0634(.A(new_n309), .B(new_n789), .C1(G107), .C2(new_n790), .ZN(new_n835));
  OAI21_X1  g0635(.A(new_n835), .B1(new_n557), .B2(new_n801), .ZN(new_n836));
  INV_X1    g0636(.A(G294), .ZN(new_n837));
  OAI22_X1  g0637(.A1(new_n563), .A2(new_n774), .B1(new_n785), .B2(new_n837), .ZN(new_n838));
  NOR3_X1   g0638(.A1(new_n834), .A2(new_n836), .A3(new_n838), .ZN(new_n839));
  NOR2_X1   g0639(.A1(new_n798), .A2(KEYINPUT96), .ZN(new_n840));
  INV_X1    g0640(.A(KEYINPUT96), .ZN(new_n841));
  NOR2_X1   g0641(.A1(new_n780), .A2(new_n841), .ZN(new_n842));
  NOR2_X1   g0642(.A1(new_n840), .A2(new_n842), .ZN(new_n843));
  INV_X1    g0643(.A(new_n843), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n844), .A2(G283), .ZN(new_n845));
  AOI22_X1  g0645(.A1(new_n784), .A2(G137), .B1(new_n786), .B2(G143), .ZN(new_n846));
  OAI21_X1  g0646(.A(new_n846), .B1(new_n793), .B2(new_n774), .ZN(new_n847));
  AOI21_X1  g0647(.A(new_n847), .B1(G150), .B2(new_n780), .ZN(new_n848));
  OR2_X1    g0648(.A1(new_n848), .A2(KEYINPUT34), .ZN(new_n849));
  NAND2_X1  g0649(.A1(new_n773), .A2(G68), .ZN(new_n850));
  OAI21_X1  g0650(.A(new_n309), .B1(new_n764), .B2(new_n253), .ZN(new_n851));
  AOI21_X1  g0651(.A(new_n851), .B1(G132), .B2(new_n761), .ZN(new_n852));
  OAI211_X1 g0652(.A(new_n850), .B(new_n852), .C1(new_n258), .C2(new_n766), .ZN(new_n853));
  AOI21_X1  g0653(.A(new_n853), .B1(new_n848), .B2(KEYINPUT34), .ZN(new_n854));
  AOI22_X1  g0654(.A1(new_n839), .A2(new_n845), .B1(new_n849), .B2(new_n854), .ZN(new_n855));
  INV_X1    g0655(.A(new_n754), .ZN(new_n856));
  OAI221_X1 g0656(.A(new_n738), .B1(G77), .B2(new_n830), .C1(new_n855), .C2(new_n856), .ZN(new_n857));
  XNOR2_X1  g0657(.A(new_n857), .B(KEYINPUT98), .ZN(new_n858));
  OAI21_X1  g0658(.A(new_n858), .B1(new_n750), .B2(new_n823), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n828), .A2(new_n859), .ZN(G384));
  OR2_X1    g0660(.A1(new_n498), .A2(KEYINPUT35), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n498), .A2(KEYINPUT35), .ZN(new_n862));
  NAND4_X1  g0662(.A1(new_n861), .A2(G116), .A3(new_n215), .A4(new_n862), .ZN(new_n863));
  XOR2_X1   g0663(.A(new_n863), .B(KEYINPUT36), .Z(new_n864));
  OAI211_X1 g0664(.A(new_n213), .B(G77), .C1(new_n258), .C2(new_n270), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n253), .A2(G68), .ZN(new_n866));
  AOI211_X1 g0666(.A(new_n205), .B(G13), .C1(new_n865), .C2(new_n866), .ZN(new_n867));
  NOR2_X1   g0667(.A1(new_n864), .A2(new_n867), .ZN(new_n868));
  INV_X1    g0668(.A(KEYINPUT39), .ZN(new_n869));
  OAI21_X1  g0669(.A(new_n451), .B1(new_n396), .B2(new_n450), .ZN(new_n870));
  AOI21_X1  g0670(.A(new_n662), .B1(new_n870), .B2(new_n394), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n458), .A2(new_n871), .ZN(new_n872));
  INV_X1    g0672(.A(new_n425), .ZN(new_n873));
  AOI22_X1  g0673(.A1(new_n873), .A2(new_n662), .B1(new_n870), .B2(new_n394), .ZN(new_n874));
  NOR2_X1   g0674(.A1(new_n417), .A2(new_n441), .ZN(new_n875));
  OAI21_X1  g0675(.A(KEYINPUT37), .B1(new_n874), .B2(new_n875), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n448), .A2(new_n451), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n423), .A2(new_n384), .ZN(new_n878));
  NAND3_X1  g0678(.A1(new_n878), .A2(KEYINPUT76), .A3(new_n438), .ZN(new_n879));
  NAND4_X1  g0679(.A1(new_n877), .A2(new_n394), .A3(new_n436), .A4(new_n879), .ZN(new_n880));
  XNOR2_X1  g0680(.A(new_n662), .B(KEYINPUT101), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n417), .A2(new_n881), .ZN(new_n882));
  INV_X1    g0682(.A(KEYINPUT37), .ZN(new_n883));
  NAND4_X1  g0683(.A1(new_n880), .A2(new_n426), .A3(new_n882), .A4(new_n883), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n876), .A2(new_n884), .ZN(new_n885));
  NAND3_X1  g0685(.A1(new_n872), .A2(KEYINPUT38), .A3(new_n885), .ZN(new_n886));
  NAND3_X1  g0686(.A1(new_n880), .A2(new_n426), .A3(new_n882), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n887), .A2(KEYINPUT37), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n888), .A2(new_n884), .ZN(new_n889));
  INV_X1    g0689(.A(new_n882), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n458), .A2(new_n890), .ZN(new_n891));
  AOI21_X1  g0691(.A(KEYINPUT38), .B1(new_n889), .B2(new_n891), .ZN(new_n892));
  OAI21_X1  g0692(.A(new_n886), .B1(new_n892), .B2(KEYINPUT102), .ZN(new_n893));
  AOI22_X1  g0693(.A1(new_n884), .A2(new_n888), .B1(new_n458), .B2(new_n890), .ZN(new_n894));
  INV_X1    g0694(.A(KEYINPUT102), .ZN(new_n895));
  NOR3_X1   g0695(.A1(new_n894), .A2(new_n895), .A3(KEYINPUT38), .ZN(new_n896));
  OAI21_X1  g0696(.A(new_n869), .B1(new_n893), .B2(new_n896), .ZN(new_n897));
  NOR2_X1   g0697(.A1(new_n620), .A2(new_n664), .ZN(new_n898));
  AND3_X1   g0698(.A1(new_n872), .A2(KEYINPUT38), .A3(new_n885), .ZN(new_n899));
  AOI21_X1  g0699(.A(KEYINPUT38), .B1(new_n872), .B2(new_n885), .ZN(new_n900));
  NOR3_X1   g0700(.A1(new_n899), .A2(new_n900), .A3(new_n869), .ZN(new_n901));
  INV_X1    g0701(.A(new_n901), .ZN(new_n902));
  NAND3_X1  g0702(.A1(new_n897), .A2(new_n898), .A3(new_n902), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n812), .A2(new_n671), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n619), .A2(new_n664), .ZN(new_n905));
  NAND3_X1  g0705(.A1(new_n620), .A2(new_n387), .A3(new_n905), .ZN(new_n906));
  OAI211_X1 g0706(.A(new_n619), .B(new_n664), .C1(new_n618), .C2(new_n388), .ZN(new_n907));
  AOI22_X1  g0707(.A1(new_n820), .A2(new_n904), .B1(new_n906), .B2(new_n907), .ZN(new_n908));
  OR2_X1    g0708(.A1(new_n899), .A2(new_n900), .ZN(new_n909));
  INV_X1    g0709(.A(new_n881), .ZN(new_n910));
  AOI22_X1  g0710(.A1(new_n908), .A2(new_n909), .B1(new_n624), .B2(new_n910), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n903), .A2(new_n911), .ZN(new_n912));
  XNOR2_X1  g0712(.A(new_n912), .B(KEYINPUT104), .ZN(new_n913));
  OAI21_X1  g0713(.A(new_n459), .B1(new_n728), .B2(new_n730), .ZN(new_n914));
  INV_X1    g0714(.A(new_n914), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n718), .A2(new_n720), .ZN(new_n916));
  AOI21_X1  g0716(.A(new_n916), .B1(new_n711), .B2(new_n655), .ZN(new_n917));
  AOI21_X1  g0717(.A(new_n664), .B1(new_n917), .B2(new_n715), .ZN(new_n918));
  AOI21_X1  g0718(.A(KEYINPUT90), .B1(new_n918), .B2(KEYINPUT29), .ZN(new_n919));
  INV_X1    g0719(.A(new_n726), .ZN(new_n920));
  OAI21_X1  g0720(.A(new_n915), .B1(new_n919), .B2(new_n920), .ZN(new_n921));
  INV_X1    g0721(.A(KEYINPUT103), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  NAND3_X1  g0723(.A1(new_n727), .A2(KEYINPUT103), .A3(new_n915), .ZN(new_n924));
  AOI21_X1  g0724(.A(new_n631), .B1(new_n923), .B2(new_n924), .ZN(new_n925));
  XNOR2_X1  g0725(.A(new_n913), .B(new_n925), .ZN(new_n926));
  INV_X1    g0726(.A(new_n823), .ZN(new_n927));
  AOI21_X1  g0727(.A(new_n927), .B1(new_n906), .B2(new_n907), .ZN(new_n928));
  OAI21_X1  g0728(.A(KEYINPUT105), .B1(new_n703), .B2(KEYINPUT31), .ZN(new_n929));
  INV_X1    g0729(.A(KEYINPUT105), .ZN(new_n930));
  OAI211_X1 g0730(.A(new_n930), .B(new_n705), .C1(new_n706), .C2(new_n671), .ZN(new_n931));
  NAND4_X1  g0731(.A1(new_n929), .A2(new_n704), .A3(new_n688), .A4(new_n931), .ZN(new_n932));
  AND2_X1   g0732(.A1(new_n928), .A2(new_n932), .ZN(new_n933));
  INV_X1    g0733(.A(KEYINPUT40), .ZN(new_n934));
  NAND3_X1  g0734(.A1(new_n933), .A2(new_n934), .A3(new_n909), .ZN(new_n935));
  NOR2_X1   g0735(.A1(new_n893), .A2(new_n896), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n928), .A2(new_n932), .ZN(new_n937));
  OAI21_X1  g0737(.A(KEYINPUT40), .B1(new_n936), .B2(new_n937), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n935), .A2(new_n938), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n932), .A2(new_n459), .ZN(new_n940));
  XOR2_X1   g0740(.A(new_n940), .B(KEYINPUT106), .Z(new_n941));
  OAI21_X1  g0741(.A(G330), .B1(new_n939), .B2(new_n941), .ZN(new_n942));
  OR2_X1    g0742(.A1(new_n942), .A2(KEYINPUT107), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n942), .A2(KEYINPUT107), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n939), .A2(new_n941), .ZN(new_n945));
  NAND3_X1  g0745(.A1(new_n943), .A2(new_n944), .A3(new_n945), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n926), .A2(new_n946), .ZN(new_n947));
  OAI21_X1  g0747(.A(new_n947), .B1(new_n205), .B2(new_n735), .ZN(new_n948));
  NOR2_X1   g0748(.A1(new_n926), .A2(new_n946), .ZN(new_n949));
  OAI21_X1  g0749(.A(new_n868), .B1(new_n948), .B2(new_n949), .ZN(G367));
  OAI21_X1  g0750(.A(new_n510), .B1(new_n501), .B2(new_n671), .ZN(new_n951));
  NAND3_X1  g0751(.A1(new_n638), .A2(new_n504), .A3(new_n664), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n951), .A2(new_n952), .ZN(new_n953));
  INV_X1    g0753(.A(new_n677), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n953), .A2(new_n954), .ZN(new_n955));
  INV_X1    g0755(.A(KEYINPUT42), .ZN(new_n956));
  XNOR2_X1  g0756(.A(new_n955), .B(new_n956), .ZN(new_n957));
  AND2_X1   g0757(.A1(new_n951), .A2(new_n952), .ZN(new_n958));
  NOR2_X1   g0758(.A1(new_n958), .A2(new_n548), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n502), .A2(new_n507), .ZN(new_n960));
  OAI21_X1  g0760(.A(new_n671), .B1(new_n959), .B2(new_n960), .ZN(new_n961));
  NOR2_X1   g0761(.A1(new_n639), .A2(new_n671), .ZN(new_n962));
  OR2_X1    g0762(.A1(new_n649), .A2(new_n962), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n719), .A2(new_n962), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n963), .A2(new_n964), .ZN(new_n965));
  AOI22_X1  g0765(.A1(new_n957), .A2(new_n961), .B1(KEYINPUT43), .B2(new_n965), .ZN(new_n966));
  OR2_X1    g0766(.A1(new_n965), .A2(KEYINPUT43), .ZN(new_n967));
  XNOR2_X1  g0767(.A(new_n966), .B(new_n967), .ZN(new_n968));
  NOR2_X1   g0768(.A1(new_n675), .A2(new_n958), .ZN(new_n969));
  XNOR2_X1  g0769(.A(new_n968), .B(new_n969), .ZN(new_n970));
  XOR2_X1   g0770(.A(new_n682), .B(KEYINPUT41), .Z(new_n971));
  OAI21_X1  g0771(.A(new_n732), .B1(new_n919), .B2(new_n920), .ZN(new_n972));
  OAI21_X1  g0772(.A(new_n677), .B1(new_n674), .B2(new_n676), .ZN(new_n973));
  XNOR2_X1  g0773(.A(new_n973), .B(new_n669), .ZN(new_n974));
  INV_X1    g0774(.A(new_n974), .ZN(new_n975));
  NAND3_X1  g0775(.A1(new_n972), .A2(new_n709), .A3(new_n975), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n976), .A2(KEYINPUT108), .ZN(new_n977));
  INV_X1    g0777(.A(KEYINPUT108), .ZN(new_n978));
  NAND3_X1  g0778(.A1(new_n733), .A2(new_n978), .A3(new_n975), .ZN(new_n979));
  INV_X1    g0779(.A(KEYINPUT45), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n677), .A2(new_n678), .ZN(new_n981));
  OAI21_X1  g0781(.A(new_n980), .B1(new_n958), .B2(new_n981), .ZN(new_n982));
  NAND3_X1  g0782(.A1(new_n679), .A2(new_n953), .A3(KEYINPUT45), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n982), .A2(new_n983), .ZN(new_n984));
  NAND3_X1  g0784(.A1(new_n958), .A2(KEYINPUT44), .A3(new_n981), .ZN(new_n985));
  INV_X1    g0785(.A(KEYINPUT44), .ZN(new_n986));
  OAI21_X1  g0786(.A(new_n986), .B1(new_n679), .B2(new_n953), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n985), .A2(new_n987), .ZN(new_n988));
  NAND2_X1  g0788(.A1(new_n984), .A2(new_n988), .ZN(new_n989));
  INV_X1    g0789(.A(new_n675), .ZN(new_n990));
  NAND2_X1  g0790(.A1(new_n989), .A2(new_n990), .ZN(new_n991));
  NAND3_X1  g0791(.A1(new_n984), .A2(new_n988), .A3(new_n675), .ZN(new_n992));
  NAND2_X1  g0792(.A1(new_n991), .A2(new_n992), .ZN(new_n993));
  INV_X1    g0793(.A(new_n993), .ZN(new_n994));
  NAND3_X1  g0794(.A1(new_n977), .A2(new_n979), .A3(new_n994), .ZN(new_n995));
  AOI21_X1  g0795(.A(new_n971), .B1(new_n995), .B2(new_n733), .ZN(new_n996));
  OAI21_X1  g0796(.A(new_n970), .B1(new_n996), .B2(new_n737), .ZN(new_n997));
  AND2_X1   g0797(.A1(new_n744), .A2(new_n234), .ZN(new_n998));
  OAI21_X1  g0798(.A(new_n755), .B1(new_n209), .B2(new_n320), .ZN(new_n999));
  INV_X1    g0799(.A(G137), .ZN(new_n1000));
  OAI221_X1 g0800(.A(new_n309), .B1(new_n760), .B2(new_n1000), .C1(new_n764), .C2(new_n258), .ZN(new_n1001));
  AOI22_X1  g0801(.A1(new_n784), .A2(G143), .B1(G50), .B2(new_n775), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n773), .A2(G77), .ZN(new_n1003));
  INV_X1    g0803(.A(G150), .ZN(new_n1004));
  OAI211_X1 g0804(.A(new_n1002), .B(new_n1003), .C1(new_n1004), .C2(new_n785), .ZN(new_n1005));
  AOI211_X1 g0805(.A(new_n1001), .B(new_n1005), .C1(G68), .C2(new_n767), .ZN(new_n1006));
  OAI21_X1  g0806(.A(new_n1006), .B1(new_n793), .B2(new_n843), .ZN(new_n1007));
  AOI22_X1  g0807(.A1(new_n784), .A2(G311), .B1(G283), .B2(new_n775), .ZN(new_n1008));
  NAND2_X1  g0808(.A1(new_n773), .A2(G97), .ZN(new_n1009));
  OAI211_X1 g0809(.A(new_n1008), .B(new_n1009), .C1(new_n557), .C2(new_n785), .ZN(new_n1010));
  AOI21_X1  g0810(.A(new_n309), .B1(new_n761), .B2(G317), .ZN(new_n1011));
  OAI21_X1  g0811(.A(new_n1011), .B1(new_n493), .B2(new_n766), .ZN(new_n1012));
  NOR2_X1   g0812(.A1(new_n764), .A2(new_n563), .ZN(new_n1013));
  XNOR2_X1  g0813(.A(new_n1013), .B(KEYINPUT46), .ZN(new_n1014));
  NOR3_X1   g0814(.A1(new_n1010), .A2(new_n1012), .A3(new_n1014), .ZN(new_n1015));
  OAI21_X1  g0815(.A(new_n1015), .B1(new_n837), .B2(new_n843), .ZN(new_n1016));
  NAND2_X1  g0816(.A1(new_n1007), .A2(new_n1016), .ZN(new_n1017));
  XOR2_X1   g0817(.A(new_n1017), .B(KEYINPUT47), .Z(new_n1018));
  OAI221_X1 g0818(.A(new_n738), .B1(new_n998), .B2(new_n999), .C1(new_n1018), .C2(new_n856), .ZN(new_n1019));
  XOR2_X1   g0819(.A(new_n1019), .B(KEYINPUT109), .Z(new_n1020));
  NAND3_X1  g0820(.A1(new_n963), .A2(new_n753), .A3(new_n964), .ZN(new_n1021));
  NAND2_X1  g0821(.A1(new_n1020), .A2(new_n1021), .ZN(new_n1022));
  XNOR2_X1  g0822(.A(new_n1022), .B(KEYINPUT110), .ZN(new_n1023));
  NAND2_X1  g0823(.A1(new_n997), .A2(new_n1023), .ZN(G387));
  AOI21_X1  g0824(.A(new_n978), .B1(new_n733), .B2(new_n975), .ZN(new_n1025));
  AOI22_X1  g0825(.A1(new_n725), .A2(new_n726), .B1(new_n729), .B2(new_n731), .ZN(new_n1026));
  NOR4_X1   g0826(.A1(new_n1026), .A2(KEYINPUT108), .A3(new_n710), .A4(new_n974), .ZN(new_n1027));
  OAI221_X1 g0827(.A(new_n682), .B1(new_n733), .B2(new_n975), .C1(new_n1025), .C2(new_n1027), .ZN(new_n1028));
  INV_X1    g0828(.A(new_n738), .ZN(new_n1029));
  NAND2_X1  g0829(.A1(new_n231), .A2(G45), .ZN(new_n1030));
  XNOR2_X1  g0830(.A(new_n1030), .B(KEYINPUT111), .ZN(new_n1031));
  NAND2_X1  g0831(.A1(new_n262), .A2(new_n253), .ZN(new_n1032));
  XNOR2_X1  g0832(.A(new_n1032), .B(KEYINPUT50), .ZN(new_n1033));
  OAI211_X1 g0833(.A(new_n684), .B(new_n292), .C1(new_n270), .C2(new_n321), .ZN(new_n1034));
  OAI211_X1 g0834(.A(new_n1031), .B(new_n744), .C1(new_n1033), .C2(new_n1034), .ZN(new_n1035));
  OAI221_X1 g0835(.A(new_n1035), .B1(G107), .B2(new_n209), .C1(new_n684), .C2(new_n741), .ZN(new_n1036));
  AOI21_X1  g0836(.A(new_n1029), .B1(new_n1036), .B2(new_n755), .ZN(new_n1037));
  OAI21_X1  g0837(.A(new_n1037), .B1(new_n674), .B2(new_n752), .ZN(new_n1038));
  AOI22_X1  g0838(.A1(new_n784), .A2(G159), .B1(G68), .B2(new_n775), .ZN(new_n1039));
  OAI211_X1 g0839(.A(new_n1039), .B(new_n1009), .C1(new_n253), .C2(new_n785), .ZN(new_n1040));
  NOR2_X1   g0840(.A1(new_n766), .A2(new_n320), .ZN(new_n1041));
  NAND2_X1  g0841(.A1(new_n790), .A2(G77), .ZN(new_n1042));
  OAI211_X1 g0842(.A(new_n1042), .B(new_n309), .C1(new_n1004), .C2(new_n760), .ZN(new_n1043));
  NOR3_X1   g0843(.A1(new_n1040), .A2(new_n1041), .A3(new_n1043), .ZN(new_n1044));
  OAI21_X1  g0844(.A(new_n1044), .B1(new_n393), .B2(new_n798), .ZN(new_n1045));
  INV_X1    g0845(.A(G322), .ZN(new_n1046));
  OAI22_X1  g0846(.A1(new_n801), .A2(new_n1046), .B1(new_n557), .B2(new_n774), .ZN(new_n1047));
  AOI21_X1  g0847(.A(new_n1047), .B1(G317), .B2(new_n786), .ZN(new_n1048));
  OAI21_X1  g0848(.A(new_n1048), .B1(new_n843), .B2(new_n832), .ZN(new_n1049));
  INV_X1    g0849(.A(KEYINPUT48), .ZN(new_n1050));
  OR2_X1    g0850(.A1(new_n1049), .A2(new_n1050), .ZN(new_n1051));
  NAND2_X1  g0851(.A1(new_n1049), .A2(new_n1050), .ZN(new_n1052));
  AOI22_X1  g0852(.A1(new_n790), .A2(G294), .B1(new_n767), .B2(G283), .ZN(new_n1053));
  NAND3_X1  g0853(.A1(new_n1051), .A2(new_n1052), .A3(new_n1053), .ZN(new_n1054));
  XOR2_X1   g0854(.A(new_n1054), .B(KEYINPUT49), .Z(new_n1055));
  AOI21_X1  g0855(.A(new_n309), .B1(new_n761), .B2(G326), .ZN(new_n1056));
  INV_X1    g0856(.A(new_n773), .ZN(new_n1057));
  OAI21_X1  g0857(.A(new_n1056), .B1(new_n1057), .B2(new_n563), .ZN(new_n1058));
  OAI21_X1  g0858(.A(new_n1045), .B1(new_n1055), .B2(new_n1058), .ZN(new_n1059));
  AOI21_X1  g0859(.A(new_n1038), .B1(new_n1059), .B2(new_n754), .ZN(new_n1060));
  XNOR2_X1  g0860(.A(new_n1060), .B(KEYINPUT112), .ZN(new_n1061));
  NOR2_X1   g0861(.A1(new_n974), .A2(new_n736), .ZN(new_n1062));
  INV_X1    g0862(.A(new_n1062), .ZN(new_n1063));
  NAND2_X1  g0863(.A1(new_n1061), .A2(new_n1063), .ZN(new_n1064));
  INV_X1    g0864(.A(new_n1064), .ZN(new_n1065));
  NAND2_X1  g0865(.A1(new_n1028), .A2(new_n1065), .ZN(G393));
  NAND3_X1  g0866(.A1(new_n991), .A2(new_n737), .A3(new_n992), .ZN(new_n1067));
  NAND2_X1  g0867(.A1(new_n958), .A2(new_n753), .ZN(new_n1068));
  XNOR2_X1  g0868(.A(new_n1068), .B(KEYINPUT113), .ZN(new_n1069));
  AOI21_X1  g0869(.A(new_n756), .B1(G97), .B2(new_n681), .ZN(new_n1070));
  NAND2_X1  g0870(.A1(new_n744), .A2(new_n242), .ZN(new_n1071));
  AOI21_X1  g0871(.A(new_n1029), .B1(new_n1070), .B2(new_n1071), .ZN(new_n1072));
  NAND2_X1  g0872(.A1(new_n844), .A2(G50), .ZN(new_n1073));
  OAI22_X1  g0873(.A1(new_n801), .A2(new_n1004), .B1(new_n793), .B2(new_n785), .ZN(new_n1074));
  XOR2_X1   g0874(.A(new_n1074), .B(KEYINPUT51), .Z(new_n1075));
  NAND2_X1  g0875(.A1(new_n767), .A2(G77), .ZN(new_n1076));
  OAI21_X1  g0876(.A(new_n309), .B1(new_n764), .B2(new_n270), .ZN(new_n1077));
  AOI21_X1  g0877(.A(new_n1077), .B1(G143), .B2(new_n761), .ZN(new_n1078));
  NAND2_X1  g0878(.A1(new_n775), .A2(new_n262), .ZN(new_n1079));
  NAND4_X1  g0879(.A1(new_n831), .A2(new_n1076), .A3(new_n1078), .A4(new_n1079), .ZN(new_n1080));
  NOR2_X1   g0880(.A1(new_n1075), .A2(new_n1080), .ZN(new_n1081));
  NAND2_X1  g0881(.A1(new_n844), .A2(G303), .ZN(new_n1082));
  INV_X1    g0882(.A(G283), .ZN(new_n1083));
  OAI221_X1 g0883(.A(new_n286), .B1(new_n760), .B2(new_n1046), .C1(new_n764), .C2(new_n1083), .ZN(new_n1084));
  AOI21_X1  g0884(.A(new_n1084), .B1(G116), .B2(new_n767), .ZN(new_n1085));
  OAI211_X1 g0885(.A(new_n1085), .B(new_n797), .C1(new_n837), .C2(new_n774), .ZN(new_n1086));
  AOI22_X1  g0886(.A1(new_n784), .A2(G317), .B1(new_n786), .B2(G311), .ZN(new_n1087));
  XOR2_X1   g0887(.A(KEYINPUT114), .B(KEYINPUT52), .Z(new_n1088));
  INV_X1    g0888(.A(new_n1088), .ZN(new_n1089));
  AND2_X1   g0889(.A1(new_n1087), .A2(new_n1089), .ZN(new_n1090));
  NOR2_X1   g0890(.A1(new_n1087), .A2(new_n1089), .ZN(new_n1091));
  NOR3_X1   g0891(.A1(new_n1086), .A2(new_n1090), .A3(new_n1091), .ZN(new_n1092));
  AOI22_X1  g0892(.A1(new_n1073), .A2(new_n1081), .B1(new_n1082), .B2(new_n1092), .ZN(new_n1093));
  OAI211_X1 g0893(.A(new_n1069), .B(new_n1072), .C1(new_n856), .C2(new_n1093), .ZN(new_n1094));
  AND3_X1   g0894(.A1(new_n1067), .A2(KEYINPUT115), .A3(new_n1094), .ZN(new_n1095));
  AOI21_X1  g0895(.A(KEYINPUT115), .B1(new_n1067), .B2(new_n1094), .ZN(new_n1096));
  NOR2_X1   g0896(.A1(new_n1095), .A2(new_n1096), .ZN(new_n1097));
  NOR2_X1   g0897(.A1(new_n1025), .A2(new_n1027), .ZN(new_n1098));
  AOI21_X1  g0898(.A(new_n683), .B1(new_n1098), .B2(new_n994), .ZN(new_n1099));
  OAI21_X1  g0899(.A(new_n993), .B1(new_n1025), .B2(new_n1027), .ZN(new_n1100));
  AOI21_X1  g0900(.A(new_n1097), .B1(new_n1099), .B2(new_n1100), .ZN(new_n1101));
  INV_X1    g0901(.A(new_n1101), .ZN(G390));
  NAND2_X1  g0902(.A1(new_n892), .A2(KEYINPUT102), .ZN(new_n1103));
  OAI21_X1  g0903(.A(new_n895), .B1(new_n894), .B2(KEYINPUT38), .ZN(new_n1104));
  NAND3_X1  g0904(.A1(new_n1103), .A2(new_n1104), .A3(new_n886), .ZN(new_n1105));
  AOI21_X1  g0905(.A(new_n901), .B1(new_n1105), .B2(new_n869), .ZN(new_n1106));
  NOR2_X1   g0906(.A1(new_n908), .A2(new_n898), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n906), .A2(new_n907), .ZN(new_n1108));
  INV_X1    g0908(.A(new_n1108), .ZN(new_n1109));
  NAND3_X1  g0909(.A1(new_n722), .A2(new_n671), .A3(new_n813), .ZN(new_n1110));
  AOI21_X1  g0910(.A(new_n1109), .B1(new_n1110), .B2(new_n904), .ZN(new_n1111));
  OAI22_X1  g0911(.A1(new_n893), .A2(new_n896), .B1(new_n620), .B2(new_n664), .ZN(new_n1112));
  OAI22_X1  g0912(.A1(new_n1106), .A2(new_n1107), .B1(new_n1111), .B2(new_n1112), .ZN(new_n1113));
  AND2_X1   g0913(.A1(new_n932), .A2(G330), .ZN(new_n1114));
  NAND3_X1  g0914(.A1(new_n1114), .A2(KEYINPUT116), .A3(new_n928), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n1113), .A2(new_n1115), .ZN(new_n1116));
  NAND2_X1  g0916(.A1(new_n889), .A2(new_n891), .ZN(new_n1117));
  INV_X1    g0917(.A(KEYINPUT38), .ZN(new_n1118));
  NAND2_X1  g0918(.A1(new_n1117), .A2(new_n1118), .ZN(new_n1119));
  AOI21_X1  g0919(.A(new_n899), .B1(new_n1119), .B2(new_n895), .ZN(new_n1120));
  AOI21_X1  g0920(.A(KEYINPUT39), .B1(new_n1120), .B2(new_n1103), .ZN(new_n1121));
  OAI22_X1  g0921(.A1(new_n1121), .A2(new_n901), .B1(new_n898), .B2(new_n908), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n1110), .A2(new_n904), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n1123), .A2(new_n1108), .ZN(new_n1124));
  AOI21_X1  g0924(.A(new_n898), .B1(new_n1120), .B2(new_n1103), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n1124), .A2(new_n1125), .ZN(new_n1126));
  NAND3_X1  g0926(.A1(new_n708), .A2(G330), .A3(new_n823), .ZN(new_n1127));
  NOR2_X1   g0927(.A1(new_n1127), .A2(new_n1109), .ZN(new_n1128));
  INV_X1    g0928(.A(KEYINPUT116), .ZN(new_n1129));
  NAND4_X1  g0929(.A1(new_n928), .A2(new_n1129), .A3(G330), .A4(new_n932), .ZN(new_n1130));
  AND2_X1   g0930(.A1(new_n1128), .A2(new_n1130), .ZN(new_n1131));
  NAND3_X1  g0931(.A1(new_n1122), .A2(new_n1126), .A3(new_n1131), .ZN(new_n1132));
  NAND2_X1  g0932(.A1(new_n1114), .A2(new_n459), .ZN(new_n1133));
  AOI21_X1  g0933(.A(KEYINPUT103), .B1(new_n727), .B2(new_n915), .ZN(new_n1134));
  AOI211_X1 g0934(.A(new_n922), .B(new_n914), .C1(new_n725), .C2(new_n726), .ZN(new_n1135));
  OAI211_X1 g0935(.A(new_n632), .B(new_n1133), .C1(new_n1134), .C2(new_n1135), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n820), .A2(new_n904), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n1114), .A2(new_n928), .ZN(new_n1138));
  NAND2_X1  g0938(.A1(new_n1127), .A2(new_n1109), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n1138), .A2(new_n1139), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n1114), .A2(new_n823), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n1141), .A2(new_n1109), .ZN(new_n1142));
  NOR2_X1   g0942(.A1(new_n1128), .A2(new_n1123), .ZN(new_n1143));
  AOI22_X1  g0943(.A1(new_n1137), .A2(new_n1140), .B1(new_n1142), .B2(new_n1143), .ZN(new_n1144));
  OAI211_X1 g0944(.A(new_n1116), .B(new_n1132), .C1(new_n1136), .C2(new_n1144), .ZN(new_n1145));
  NAND2_X1  g0945(.A1(new_n1116), .A2(new_n1132), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n1140), .A2(new_n1137), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n1142), .A2(new_n1143), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n1147), .A2(new_n1148), .ZN(new_n1149));
  NAND4_X1  g0949(.A1(new_n1146), .A2(new_n925), .A3(new_n1133), .A4(new_n1149), .ZN(new_n1150));
  NAND3_X1  g0950(.A1(new_n1145), .A2(new_n1150), .A3(new_n682), .ZN(new_n1151));
  NOR2_X1   g0951(.A1(new_n1106), .A2(new_n750), .ZN(new_n1152));
  AOI21_X1  g0952(.A(new_n1029), .B1(new_n393), .B2(new_n829), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n761), .A2(G294), .ZN(new_n1154));
  NAND4_X1  g0954(.A1(new_n791), .A2(new_n1154), .A3(new_n1076), .A4(new_n286), .ZN(new_n1155));
  AOI22_X1  g0955(.A1(new_n786), .A2(G116), .B1(new_n775), .B2(G97), .ZN(new_n1156));
  OAI211_X1 g0956(.A(new_n850), .B(new_n1156), .C1(new_n1083), .C2(new_n801), .ZN(new_n1157));
  AOI211_X1 g0957(.A(new_n1155), .B(new_n1157), .C1(new_n844), .C2(G107), .ZN(new_n1158));
  XNOR2_X1  g0958(.A(KEYINPUT54), .B(G143), .ZN(new_n1159));
  OAI22_X1  g0959(.A1(new_n843), .A2(new_n1000), .B1(new_n774), .B2(new_n1159), .ZN(new_n1160));
  NOR2_X1   g0960(.A1(new_n1160), .A2(KEYINPUT117), .ZN(new_n1161));
  AOI21_X1  g0961(.A(new_n286), .B1(new_n761), .B2(G125), .ZN(new_n1162));
  OAI221_X1 g0962(.A(new_n1162), .B1(new_n793), .B2(new_n766), .C1(new_n1057), .C2(new_n253), .ZN(new_n1163));
  NOR2_X1   g0963(.A1(new_n764), .A2(new_n1004), .ZN(new_n1164));
  XNOR2_X1  g0964(.A(new_n1164), .B(KEYINPUT53), .ZN(new_n1165));
  INV_X1    g0965(.A(G128), .ZN(new_n1166));
  INV_X1    g0966(.A(G132), .ZN(new_n1167));
  OAI221_X1 g0967(.A(new_n1165), .B1(new_n1166), .B2(new_n801), .C1(new_n1167), .C2(new_n785), .ZN(new_n1168));
  NOR3_X1   g0968(.A1(new_n1161), .A2(new_n1163), .A3(new_n1168), .ZN(new_n1169));
  NAND2_X1  g0969(.A1(new_n1160), .A2(KEYINPUT117), .ZN(new_n1170));
  AOI21_X1  g0970(.A(new_n1158), .B1(new_n1169), .B2(new_n1170), .ZN(new_n1171));
  OAI21_X1  g0971(.A(new_n1153), .B1(new_n1171), .B2(new_n856), .ZN(new_n1172));
  NOR2_X1   g0972(.A1(new_n1152), .A2(new_n1172), .ZN(new_n1173));
  AOI21_X1  g0973(.A(new_n1173), .B1(new_n1146), .B2(new_n737), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n1151), .A2(new_n1174), .ZN(G378));
  AND2_X1   g0975(.A1(new_n1116), .A2(new_n1132), .ZN(new_n1176));
  OAI211_X1 g0976(.A(new_n925), .B(new_n1133), .C1(new_n1176), .C2(new_n1144), .ZN(new_n1177));
  INV_X1    g0977(.A(G330), .ZN(new_n1178));
  AOI21_X1  g0978(.A(new_n1178), .B1(new_n935), .B2(new_n938), .ZN(new_n1179));
  NAND2_X1  g0979(.A1(new_n628), .A2(new_n308), .ZN(new_n1180));
  NOR2_X1   g0980(.A1(new_n275), .A2(new_n662), .ZN(new_n1181));
  INV_X1    g0981(.A(new_n1181), .ZN(new_n1182));
  XNOR2_X1  g0982(.A(new_n1180), .B(new_n1182), .ZN(new_n1183));
  XNOR2_X1  g0983(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1184));
  XNOR2_X1  g0984(.A(new_n1183), .B(new_n1184), .ZN(new_n1185));
  INV_X1    g0985(.A(new_n1185), .ZN(new_n1186));
  NAND2_X1  g0986(.A1(new_n912), .A2(new_n1186), .ZN(new_n1187));
  NAND3_X1  g0987(.A1(new_n903), .A2(new_n1185), .A3(new_n911), .ZN(new_n1188));
  AOI21_X1  g0988(.A(new_n1179), .B1(new_n1187), .B2(new_n1188), .ZN(new_n1189));
  INV_X1    g0989(.A(new_n1189), .ZN(new_n1190));
  NAND3_X1  g0990(.A1(new_n1187), .A2(new_n1179), .A3(new_n1188), .ZN(new_n1191));
  NAND2_X1  g0991(.A1(new_n1190), .A2(new_n1191), .ZN(new_n1192));
  AOI21_X1  g0992(.A(KEYINPUT57), .B1(new_n1177), .B2(new_n1192), .ZN(new_n1193));
  INV_X1    g0993(.A(new_n1188), .ZN(new_n1194));
  AOI21_X1  g0994(.A(new_n934), .B1(new_n933), .B2(new_n1105), .ZN(new_n1195));
  AND4_X1   g0995(.A1(new_n934), .A2(new_n909), .A3(new_n932), .A4(new_n928), .ZN(new_n1196));
  OAI21_X1  g0996(.A(G330), .B1(new_n1195), .B2(new_n1196), .ZN(new_n1197));
  AOI21_X1  g0997(.A(new_n1185), .B1(new_n903), .B2(new_n911), .ZN(new_n1198));
  NOR3_X1   g0998(.A1(new_n1194), .A2(new_n1197), .A3(new_n1198), .ZN(new_n1199));
  OAI21_X1  g0999(.A(KEYINPUT57), .B1(new_n1199), .B2(new_n1189), .ZN(new_n1200));
  AOI21_X1  g1000(.A(new_n1136), .B1(new_n1146), .B2(new_n1149), .ZN(new_n1201));
  OAI21_X1  g1001(.A(new_n682), .B1(new_n1200), .B2(new_n1201), .ZN(new_n1202));
  OR2_X1    g1002(.A1(new_n1193), .A2(new_n1202), .ZN(new_n1203));
  NAND2_X1  g1003(.A1(new_n1186), .A2(new_n749), .ZN(new_n1204));
  OAI21_X1  g1004(.A(new_n738), .B1(G50), .B2(new_n830), .ZN(new_n1205));
  XNOR2_X1  g1005(.A(new_n1205), .B(KEYINPUT121), .ZN(new_n1206));
  NOR2_X1   g1006(.A1(new_n309), .A2(G41), .ZN(new_n1207));
  OAI211_X1 g1007(.A(new_n1042), .B(new_n1207), .C1(new_n1083), .C2(new_n760), .ZN(new_n1208));
  NAND2_X1  g1008(.A1(new_n773), .A2(G58), .ZN(new_n1209));
  OAI221_X1 g1009(.A(new_n1209), .B1(new_n493), .B2(new_n785), .C1(new_n563), .C2(new_n801), .ZN(new_n1210));
  AOI211_X1 g1010(.A(new_n1208), .B(new_n1210), .C1(G68), .C2(new_n767), .ZN(new_n1211));
  AOI22_X1  g1011(.A1(new_n780), .A2(G97), .B1(new_n603), .B2(new_n775), .ZN(new_n1212));
  INV_X1    g1012(.A(KEYINPUT119), .ZN(new_n1213));
  AND2_X1   g1013(.A1(new_n1212), .A2(new_n1213), .ZN(new_n1214));
  NOR2_X1   g1014(.A1(new_n1212), .A2(new_n1213), .ZN(new_n1215));
  OAI21_X1  g1015(.A(new_n1211), .B1(new_n1214), .B2(new_n1215), .ZN(new_n1216));
  XOR2_X1   g1016(.A(KEYINPUT120), .B(KEYINPUT58), .Z(new_n1217));
  OR2_X1    g1017(.A1(new_n1216), .A2(new_n1217), .ZN(new_n1218));
  NAND2_X1  g1018(.A1(new_n1216), .A2(new_n1217), .ZN(new_n1219));
  AOI211_X1 g1019(.A(G50), .B(new_n1207), .C1(new_n367), .C2(new_n291), .ZN(new_n1220));
  XNOR2_X1  g1020(.A(new_n1220), .B(KEYINPUT118), .ZN(new_n1221));
  OAI22_X1  g1021(.A1(new_n764), .A2(new_n1159), .B1(new_n766), .B2(new_n1004), .ZN(new_n1222));
  AOI21_X1  g1022(.A(new_n1222), .B1(new_n784), .B2(G125), .ZN(new_n1223));
  AOI22_X1  g1023(.A1(new_n786), .A2(G128), .B1(new_n775), .B2(G137), .ZN(new_n1224));
  OAI211_X1 g1024(.A(new_n1223), .B(new_n1224), .C1(new_n798), .C2(new_n1167), .ZN(new_n1225));
  OR2_X1    g1025(.A1(new_n1225), .A2(KEYINPUT59), .ZN(new_n1226));
  AOI211_X1 g1026(.A(G33), .B(G41), .C1(new_n761), .C2(G124), .ZN(new_n1227));
  OAI21_X1  g1027(.A(new_n1227), .B1(new_n1057), .B2(new_n793), .ZN(new_n1228));
  AOI21_X1  g1028(.A(new_n1228), .B1(new_n1225), .B2(KEYINPUT59), .ZN(new_n1229));
  AOI21_X1  g1029(.A(new_n1221), .B1(new_n1226), .B2(new_n1229), .ZN(new_n1230));
  NAND3_X1  g1030(.A1(new_n1218), .A2(new_n1219), .A3(new_n1230), .ZN(new_n1231));
  AOI21_X1  g1031(.A(new_n1206), .B1(new_n1231), .B2(new_n754), .ZN(new_n1232));
  AOI22_X1  g1032(.A1(new_n1192), .A2(new_n737), .B1(new_n1204), .B2(new_n1232), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(new_n1203), .A2(new_n1233), .ZN(G375));
  NAND3_X1  g1034(.A1(new_n925), .A2(new_n1133), .A3(new_n1149), .ZN(new_n1235));
  NAND2_X1  g1035(.A1(new_n1136), .A2(new_n1144), .ZN(new_n1236));
  INV_X1    g1036(.A(new_n971), .ZN(new_n1237));
  NAND3_X1  g1037(.A1(new_n1235), .A2(new_n1236), .A3(new_n1237), .ZN(new_n1238));
  NAND2_X1  g1038(.A1(new_n1109), .A2(new_n749), .ZN(new_n1239));
  OAI21_X1  g1039(.A(new_n738), .B1(G68), .B2(new_n830), .ZN(new_n1240));
  NOR2_X1   g1040(.A1(new_n843), .A2(new_n563), .ZN(new_n1241));
  AOI22_X1  g1041(.A1(new_n784), .A2(G294), .B1(G107), .B2(new_n775), .ZN(new_n1242));
  OAI21_X1  g1042(.A(new_n286), .B1(new_n760), .B2(new_n557), .ZN(new_n1243));
  AOI211_X1 g1043(.A(new_n1041), .B(new_n1243), .C1(G97), .C2(new_n790), .ZN(new_n1244));
  NAND2_X1  g1044(.A1(new_n786), .A2(G283), .ZN(new_n1245));
  NAND4_X1  g1045(.A1(new_n1242), .A2(new_n1003), .A3(new_n1244), .A4(new_n1245), .ZN(new_n1246));
  NOR2_X1   g1046(.A1(new_n843), .A2(new_n1159), .ZN(new_n1247));
  AOI22_X1  g1047(.A1(new_n784), .A2(G132), .B1(G150), .B2(new_n775), .ZN(new_n1248));
  OAI221_X1 g1048(.A(new_n309), .B1(new_n760), .B2(new_n1166), .C1(new_n764), .C2(new_n793), .ZN(new_n1249));
  AOI21_X1  g1049(.A(new_n1249), .B1(G50), .B2(new_n767), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(new_n786), .A2(G137), .ZN(new_n1251));
  NAND4_X1  g1051(.A1(new_n1248), .A2(new_n1250), .A3(new_n1209), .A4(new_n1251), .ZN(new_n1252));
  OAI22_X1  g1052(.A1(new_n1241), .A2(new_n1246), .B1(new_n1247), .B2(new_n1252), .ZN(new_n1253));
  AOI21_X1  g1053(.A(new_n1240), .B1(new_n1253), .B2(new_n754), .ZN(new_n1254));
  AOI22_X1  g1054(.A1(new_n1149), .A2(new_n737), .B1(new_n1239), .B2(new_n1254), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(new_n1238), .A2(new_n1255), .ZN(G381));
  AND3_X1   g1056(.A1(new_n1028), .A2(new_n807), .A3(new_n1065), .ZN(new_n1257));
  INV_X1    g1057(.A(G384), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(new_n1257), .A2(new_n1258), .ZN(new_n1259));
  XNOR2_X1  g1059(.A(new_n1259), .B(KEYINPUT122), .ZN(new_n1260));
  NAND3_X1  g1060(.A1(new_n997), .A2(new_n1101), .A3(new_n1023), .ZN(new_n1261));
  INV_X1    g1061(.A(new_n1174), .ZN(new_n1262));
  AOI21_X1  g1062(.A(new_n683), .B1(new_n1235), .B2(new_n1176), .ZN(new_n1263));
  AOI21_X1  g1063(.A(new_n1262), .B1(new_n1263), .B2(new_n1150), .ZN(new_n1264));
  NAND3_X1  g1064(.A1(new_n1264), .A2(new_n1255), .A3(new_n1238), .ZN(new_n1265));
  OR4_X1    g1065(.A1(G375), .A2(new_n1260), .A3(new_n1261), .A4(new_n1265), .ZN(G407));
  INV_X1    g1066(.A(G213), .ZN(new_n1267));
  NOR2_X1   g1067(.A1(new_n1267), .A2(G343), .ZN(new_n1268));
  INV_X1    g1068(.A(new_n1268), .ZN(new_n1269));
  NOR3_X1   g1069(.A1(G375), .A2(G378), .A3(new_n1269), .ZN(new_n1270));
  XNOR2_X1  g1070(.A(new_n1270), .B(KEYINPUT123), .ZN(new_n1271));
  NAND3_X1  g1071(.A1(new_n1271), .A2(G213), .A3(G407), .ZN(G409));
  OAI211_X1 g1072(.A(G378), .B(new_n1233), .C1(new_n1193), .C2(new_n1202), .ZN(new_n1273));
  NOR2_X1   g1073(.A1(new_n1199), .A2(new_n1189), .ZN(new_n1274));
  NOR3_X1   g1074(.A1(new_n1274), .A2(new_n1201), .A3(new_n971), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(new_n1204), .A2(new_n1232), .ZN(new_n1276));
  OAI21_X1  g1076(.A(new_n1276), .B1(new_n1274), .B2(new_n736), .ZN(new_n1277));
  OAI21_X1  g1077(.A(new_n1264), .B1(new_n1275), .B2(new_n1277), .ZN(new_n1278));
  AOI21_X1  g1078(.A(new_n1268), .B1(new_n1273), .B2(new_n1278), .ZN(new_n1279));
  INV_X1    g1079(.A(new_n1279), .ZN(new_n1280));
  NAND2_X1  g1080(.A1(new_n1268), .A2(G2897), .ZN(new_n1281));
  NAND3_X1  g1081(.A1(new_n1136), .A2(KEYINPUT60), .A3(new_n1144), .ZN(new_n1282));
  NAND3_X1  g1082(.A1(new_n1282), .A2(new_n1235), .A3(new_n682), .ZN(new_n1283));
  AOI21_X1  g1083(.A(KEYINPUT60), .B1(new_n1136), .B2(new_n1144), .ZN(new_n1284));
  OAI211_X1 g1084(.A(G384), .B(new_n1255), .C1(new_n1283), .C2(new_n1284), .ZN(new_n1285));
  INV_X1    g1085(.A(new_n1285), .ZN(new_n1286));
  INV_X1    g1086(.A(KEYINPUT60), .ZN(new_n1287));
  NAND2_X1  g1087(.A1(new_n1236), .A2(new_n1287), .ZN(new_n1288));
  NAND4_X1  g1088(.A1(new_n1288), .A2(new_n682), .A3(new_n1235), .A4(new_n1282), .ZN(new_n1289));
  AOI21_X1  g1089(.A(G384), .B1(new_n1289), .B2(new_n1255), .ZN(new_n1290));
  OAI21_X1  g1090(.A(new_n1281), .B1(new_n1286), .B2(new_n1290), .ZN(new_n1291));
  INV_X1    g1091(.A(KEYINPUT124), .ZN(new_n1292));
  OAI21_X1  g1092(.A(new_n1255), .B1(new_n1283), .B2(new_n1284), .ZN(new_n1293));
  NAND2_X1  g1093(.A1(new_n1293), .A2(new_n1258), .ZN(new_n1294));
  INV_X1    g1094(.A(new_n1281), .ZN(new_n1295));
  NAND3_X1  g1095(.A1(new_n1294), .A2(new_n1285), .A3(new_n1295), .ZN(new_n1296));
  AND3_X1   g1096(.A1(new_n1291), .A2(new_n1292), .A3(new_n1296), .ZN(new_n1297));
  AOI21_X1  g1097(.A(new_n1292), .B1(new_n1291), .B2(new_n1296), .ZN(new_n1298));
  OAI21_X1  g1098(.A(new_n1280), .B1(new_n1297), .B2(new_n1298), .ZN(new_n1299));
  NAND2_X1  g1099(.A1(new_n1299), .A2(KEYINPUT125), .ZN(new_n1300));
  NOR2_X1   g1100(.A1(new_n1286), .A2(new_n1290), .ZN(new_n1301));
  AND3_X1   g1101(.A1(new_n1279), .A2(KEYINPUT63), .A3(new_n1301), .ZN(new_n1302));
  NAND3_X1  g1102(.A1(new_n1100), .A2(new_n995), .A3(new_n682), .ZN(new_n1303));
  OAI211_X1 g1103(.A(new_n1303), .B(KEYINPUT127), .C1(new_n1096), .C2(new_n1095), .ZN(new_n1304));
  INV_X1    g1104(.A(new_n969), .ZN(new_n1305));
  XNOR2_X1  g1105(.A(new_n968), .B(new_n1305), .ZN(new_n1306));
  NOR3_X1   g1106(.A1(new_n1025), .A2(new_n1027), .A3(new_n993), .ZN(new_n1307));
  INV_X1    g1107(.A(new_n733), .ZN(new_n1308));
  OAI21_X1  g1108(.A(new_n1237), .B1(new_n1307), .B2(new_n1308), .ZN(new_n1309));
  AOI21_X1  g1109(.A(new_n1306), .B1(new_n1309), .B2(new_n736), .ZN(new_n1310));
  XOR2_X1   g1110(.A(new_n1022), .B(KEYINPUT110), .Z(new_n1311));
  OAI21_X1  g1111(.A(new_n1304), .B1(new_n1310), .B2(new_n1311), .ZN(new_n1312));
  INV_X1    g1112(.A(KEYINPUT126), .ZN(new_n1313));
  AOI21_X1  g1113(.A(new_n807), .B1(new_n1028), .B2(new_n1065), .ZN(new_n1314));
  OR2_X1    g1114(.A1(new_n1257), .A2(new_n1314), .ZN(new_n1315));
  NAND4_X1  g1115(.A1(new_n1312), .A2(new_n1313), .A3(new_n1261), .A4(new_n1315), .ZN(new_n1316));
  NAND2_X1  g1116(.A1(new_n1261), .A2(new_n1313), .ZN(new_n1317));
  NOR2_X1   g1117(.A1(new_n1257), .A2(new_n1314), .ZN(new_n1318));
  NAND2_X1  g1118(.A1(new_n1317), .A2(new_n1318), .ZN(new_n1319));
  INV_X1    g1119(.A(KEYINPUT61), .ZN(new_n1320));
  INV_X1    g1120(.A(KEYINPUT127), .ZN(new_n1321));
  OAI211_X1 g1121(.A(G387), .B(G390), .C1(new_n1318), .C2(new_n1321), .ZN(new_n1322));
  NAND4_X1  g1122(.A1(new_n1316), .A2(new_n1319), .A3(new_n1320), .A4(new_n1322), .ZN(new_n1323));
  AOI21_X1  g1123(.A(KEYINPUT63), .B1(new_n1279), .B2(new_n1301), .ZN(new_n1324));
  NOR3_X1   g1124(.A1(new_n1302), .A2(new_n1323), .A3(new_n1324), .ZN(new_n1325));
  INV_X1    g1125(.A(KEYINPUT125), .ZN(new_n1326));
  OAI211_X1 g1126(.A(new_n1326), .B(new_n1280), .C1(new_n1297), .C2(new_n1298), .ZN(new_n1327));
  NAND3_X1  g1127(.A1(new_n1300), .A2(new_n1325), .A3(new_n1327), .ZN(new_n1328));
  NAND3_X1  g1128(.A1(new_n1316), .A2(new_n1319), .A3(new_n1322), .ZN(new_n1329));
  INV_X1    g1129(.A(new_n1301), .ZN(new_n1330));
  OAI21_X1  g1130(.A(KEYINPUT62), .B1(new_n1280), .B2(new_n1330), .ZN(new_n1331));
  NAND2_X1  g1131(.A1(new_n1291), .A2(new_n1296), .ZN(new_n1332));
  AOI21_X1  g1132(.A(KEYINPUT61), .B1(new_n1280), .B2(new_n1332), .ZN(new_n1333));
  NAND2_X1  g1133(.A1(new_n1331), .A2(new_n1333), .ZN(new_n1334));
  NOR3_X1   g1134(.A1(new_n1280), .A2(KEYINPUT62), .A3(new_n1330), .ZN(new_n1335));
  OAI21_X1  g1135(.A(new_n1329), .B1(new_n1334), .B2(new_n1335), .ZN(new_n1336));
  NAND2_X1  g1136(.A1(new_n1328), .A2(new_n1336), .ZN(G405));
  NAND2_X1  g1137(.A1(G375), .A2(new_n1264), .ZN(new_n1338));
  NAND2_X1  g1138(.A1(new_n1338), .A2(new_n1273), .ZN(new_n1339));
  NAND2_X1  g1139(.A1(new_n1339), .A2(new_n1301), .ZN(new_n1340));
  NAND3_X1  g1140(.A1(new_n1338), .A2(new_n1273), .A3(new_n1330), .ZN(new_n1341));
  NAND2_X1  g1141(.A1(new_n1340), .A2(new_n1341), .ZN(new_n1342));
  XNOR2_X1  g1142(.A(new_n1342), .B(new_n1329), .ZN(G402));
endmodule


