

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n622, n623, n624, n625, n626, n627, n628, n629, n630,
         n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641,
         n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652,
         n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663,
         n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674,
         n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685,
         n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696,
         n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707,
         n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718,
         n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729,
         n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740,
         n741, n742, n743, n744, n745, n746, n747;

  XNOR2_X1 U375 ( .A(n356), .B(n355), .ZN(n656) );
  AND2_X2 U376 ( .A1(n660), .A2(n659), .ZN(n706) );
  INV_X1 U377 ( .A(KEYINPUT79), .ZN(n355) );
  AND2_X1 U378 ( .A1(n386), .A2(n384), .ZN(n401) );
  NAND2_X1 U379 ( .A1(n539), .A2(n538), .ZN(n541) );
  BUF_X1 U380 ( .A(n625), .Z(n357) );
  XNOR2_X1 U381 ( .A(n530), .B(n364), .ZN(n421) );
  XNOR2_X1 U382 ( .A(n559), .B(n509), .ZN(n625) );
  XNOR2_X1 U383 ( .A(n428), .B(n390), .ZN(n676) );
  XNOR2_X1 U384 ( .A(n392), .B(n393), .ZN(n428) );
  NOR2_X2 U385 ( .A1(G953), .A2(G237), .ZN(n480) );
  INV_X1 U386 ( .A(G953), .ZN(n733) );
  NAND2_X2 U387 ( .A1(n606), .A2(n605), .ZN(n660) );
  XNOR2_X2 U388 ( .A(n429), .B(KEYINPUT84), .ZN(n369) );
  XNOR2_X2 U389 ( .A(n446), .B(n383), .ZN(n731) );
  XNOR2_X2 U390 ( .A(n493), .B(KEYINPUT4), .ZN(n383) );
  NAND2_X1 U391 ( .A1(n620), .A2(n659), .ZN(n356) );
  XNOR2_X1 U392 ( .A(G119), .B(G116), .ZN(n447) );
  NOR2_X1 U393 ( .A1(n537), .A2(n523), .ZN(n626) );
  NOR2_X1 U394 ( .A1(n663), .A2(G902), .ZN(n455) );
  NAND2_X1 U395 ( .A1(n607), .A2(n732), .ZN(n659) );
  AND2_X1 U396 ( .A1(n720), .A2(KEYINPUT2), .ZN(n607) );
  AND2_X1 U397 ( .A1(n539), .A2(n373), .ZN(n682) );
  OR2_X1 U398 ( .A1(n601), .A2(n697), .ZN(n571) );
  XNOR2_X1 U399 ( .A(n369), .B(n468), .ZN(n578) );
  XNOR2_X1 U400 ( .A(G137), .B(G134), .ZN(n445) );
  XNOR2_X2 U401 ( .A(n498), .B(n399), .ZN(n398) );
  NOR2_X1 U402 ( .A1(n592), .A2(n369), .ZN(n575) );
  XNOR2_X1 U403 ( .A(n731), .B(G146), .ZN(n507) );
  NOR2_X1 U404 ( .A1(n547), .A2(n546), .ZN(n441) );
  INV_X1 U405 ( .A(n741), .ZN(n430) );
  NAND2_X1 U406 ( .A1(n547), .A2(n546), .ZN(n440) );
  XNOR2_X1 U407 ( .A(n371), .B(n370), .ZN(n535) );
  INV_X1 U408 ( .A(KEYINPUT102), .ZN(n370) );
  NAND2_X1 U409 ( .A1(n375), .A2(n372), .ZN(n371) );
  NAND2_X1 U410 ( .A1(n377), .A2(n376), .ZN(n375) );
  AND2_X1 U411 ( .A1(n380), .A2(n362), .ZN(n406) );
  XNOR2_X1 U412 ( .A(n488), .B(n436), .ZN(n513) );
  INV_X1 U413 ( .A(KEYINPUT8), .ZN(n436) );
  XNOR2_X1 U414 ( .A(G125), .B(G146), .ZN(n476) );
  XNOR2_X1 U415 ( .A(n476), .B(n462), .ZN(n368) );
  XNOR2_X1 U416 ( .A(KEYINPUT18), .B(KEYINPUT17), .ZN(n462) );
  XNOR2_X1 U417 ( .A(n432), .B(n431), .ZN(n444) );
  INV_X1 U418 ( .A(KEYINPUT70), .ZN(n431) );
  NAND2_X1 U419 ( .A1(n625), .A2(n626), .ZN(n432) );
  XNOR2_X1 U420 ( .A(n507), .B(n358), .ZN(n663) );
  XNOR2_X1 U421 ( .A(n397), .B(G110), .ZN(n512) );
  INV_X1 U422 ( .A(G119), .ZN(n397) );
  XNOR2_X1 U423 ( .A(G128), .B(G137), .ZN(n510) );
  NAND2_X1 U424 ( .A1(n513), .A2(G221), .ZN(n417) );
  XNOR2_X1 U425 ( .A(n512), .B(n416), .ZN(n415) );
  INV_X1 U426 ( .A(KEYINPUT89), .ZN(n416) );
  XNOR2_X1 U427 ( .A(G122), .B(G134), .ZN(n490) );
  NAND2_X1 U428 ( .A1(n513), .A2(G217), .ZN(n435) );
  XNOR2_X1 U429 ( .A(n476), .B(n477), .ZN(n730) );
  XNOR2_X1 U430 ( .A(G140), .B(KEYINPUT10), .ZN(n477) );
  NOR2_X1 U431 ( .A1(n616), .A2(KEYINPUT2), .ZN(n617) );
  NAND2_X1 U432 ( .A1(n701), .A2(n433), .ZN(n592) );
  AND2_X1 U433 ( .A1(n574), .A2(n573), .ZN(n433) );
  INV_X1 U434 ( .A(KEYINPUT22), .ZN(n399) );
  AND2_X1 U435 ( .A1(n497), .A2(n438), .ZN(n437) );
  XNOR2_X1 U436 ( .A(n536), .B(KEYINPUT103), .ZN(n563) );
  BUF_X1 U437 ( .A(n706), .Z(n714) );
  XNOR2_X1 U438 ( .A(n507), .B(n405), .ZN(n707) );
  XNOR2_X1 U439 ( .A(KEYINPUT68), .B(G140), .ZN(n506) );
  NAND2_X1 U440 ( .A1(n379), .A2(n378), .ZN(n377) );
  INV_X1 U441 ( .A(n688), .ZN(n378) );
  INV_X1 U442 ( .A(n645), .ZN(n376) );
  INV_X1 U443 ( .A(n682), .ZN(n372) );
  INV_X1 U444 ( .A(KEYINPUT48), .ZN(n411) );
  AND2_X1 U445 ( .A1(n535), .A2(n361), .ZN(n439) );
  NAND2_X1 U446 ( .A1(G237), .A2(G234), .ZN(n469) );
  INV_X1 U447 ( .A(n523), .ZN(n438) );
  XNOR2_X1 U448 ( .A(n525), .B(n524), .ZN(n636) );
  XNOR2_X1 U449 ( .A(G902), .B(KEYINPUT15), .ZN(n603) );
  NAND2_X1 U450 ( .A1(n707), .A2(n508), .ZN(n404) );
  XNOR2_X1 U451 ( .A(n452), .B(n451), .ZN(n461) );
  INV_X1 U452 ( .A(G101), .ZN(n451) );
  XOR2_X1 U453 ( .A(KEYINPUT11), .B(KEYINPUT12), .Z(n479) );
  XNOR2_X1 U454 ( .A(G143), .B(G113), .ZN(n478) );
  XNOR2_X1 U455 ( .A(n426), .B(G104), .ZN(n422) );
  INV_X1 U456 ( .A(G122), .ZN(n426) );
  XNOR2_X1 U457 ( .A(G107), .B(G101), .ZN(n499) );
  XOR2_X1 U458 ( .A(G110), .B(G104), .Z(n500) );
  XNOR2_X1 U459 ( .A(n463), .B(n464), .ZN(n395) );
  INV_X1 U460 ( .A(n567), .ZN(n583) );
  INV_X1 U461 ( .A(KEYINPUT19), .ZN(n468) );
  XNOR2_X1 U462 ( .A(n382), .B(n381), .ZN(n521) );
  XNOR2_X1 U463 ( .A(n487), .B(G475), .ZN(n381) );
  OR2_X1 U464 ( .A1(n669), .A2(G902), .ZN(n382) );
  XNOR2_X1 U465 ( .A(n536), .B(n456), .ZN(n573) );
  XNOR2_X1 U466 ( .A(n512), .B(n422), .ZN(n393) );
  XNOR2_X1 U467 ( .A(n394), .B(n461), .ZN(n392) );
  XNOR2_X1 U468 ( .A(n424), .B(n396), .ZN(n394) );
  XNOR2_X1 U469 ( .A(n418), .B(n414), .ZN(n715) );
  XNOR2_X1 U470 ( .A(n730), .B(n514), .ZN(n418) );
  XNOR2_X1 U471 ( .A(n417), .B(n415), .ZN(n414) );
  XNOR2_X1 U472 ( .A(n495), .B(n494), .ZN(n608) );
  XNOR2_X1 U473 ( .A(n435), .B(n434), .ZN(n495) );
  AND2_X1 U474 ( .A1(n654), .A2(n443), .ZN(n655) );
  INV_X1 U475 ( .A(n653), .ZN(n419) );
  NAND2_X1 U476 ( .A1(n408), .A2(n582), .ZN(n533) );
  XNOR2_X1 U477 ( .A(n409), .B(n365), .ZN(n408) );
  INV_X1 U478 ( .A(KEYINPUT104), .ZN(n540) );
  XNOR2_X1 U479 ( .A(n520), .B(KEYINPUT98), .ZN(n701) );
  AND2_X1 U480 ( .A1(n531), .A2(n521), .ZN(n520) );
  NOR2_X1 U481 ( .A1(n573), .A2(n374), .ZN(n373) );
  INV_X1 U482 ( .A(n622), .ZN(n374) );
  XNOR2_X1 U483 ( .A(n712), .B(n711), .ZN(n713) );
  XOR2_X1 U484 ( .A(n454), .B(n453), .Z(n358) );
  XOR2_X1 U485 ( .A(n544), .B(KEYINPUT75), .Z(n359) );
  AND2_X1 U486 ( .A1(n467), .A2(G210), .ZN(n360) );
  AND2_X1 U487 ( .A1(n534), .A2(n440), .ZN(n361) );
  AND2_X1 U488 ( .A1(n614), .A2(n548), .ZN(n362) );
  NOR2_X1 U489 ( .A1(n648), .A2(n420), .ZN(n363) );
  XOR2_X1 U490 ( .A(KEYINPUT105), .B(KEYINPUT33), .Z(n364) );
  XOR2_X1 U491 ( .A(KEYINPUT74), .B(KEYINPUT34), .Z(n365) );
  XOR2_X1 U492 ( .A(KEYINPUT82), .B(KEYINPUT46), .Z(n366) );
  XNOR2_X1 U493 ( .A(n391), .B(n395), .ZN(n390) );
  XNOR2_X2 U494 ( .A(n367), .B(KEYINPUT45), .ZN(n616) );
  NAND2_X1 U495 ( .A1(n401), .A2(n439), .ZN(n367) );
  XNOR2_X1 U496 ( .A(n600), .B(n599), .ZN(n380) );
  XNOR2_X1 U497 ( .A(n383), .B(n368), .ZN(n391) );
  XNOR2_X2 U498 ( .A(G143), .B(G128), .ZN(n493) );
  INV_X1 U499 ( .A(n700), .ZN(n379) );
  AND2_X1 U500 ( .A1(n380), .A2(n614), .ZN(n732) );
  NAND2_X1 U501 ( .A1(n385), .A2(n441), .ZN(n384) );
  INV_X1 U502 ( .A(n387), .ZN(n385) );
  NAND2_X1 U503 ( .A1(n388), .A2(n387), .ZN(n386) );
  NOR2_X2 U504 ( .A1(n400), .A2(n746), .ZN(n387) );
  NAND2_X1 U505 ( .A1(n389), .A2(KEYINPUT64), .ZN(n388) );
  NAND2_X1 U506 ( .A1(n430), .A2(n546), .ZN(n389) );
  INV_X1 U507 ( .A(KEYINPUT16), .ZN(n396) );
  AND2_X2 U508 ( .A1(n398), .A2(n543), .ZN(n539) );
  AND2_X1 U509 ( .A1(n398), .A2(n359), .ZN(n545) );
  XNOR2_X1 U510 ( .A(n400), .B(n742), .ZN(G12) );
  XNOR2_X2 U511 ( .A(n541), .B(n540), .ZN(n400) );
  INV_X2 U512 ( .A(G116), .ZN(n427) );
  XNOR2_X1 U513 ( .A(n407), .B(KEYINPUT78), .ZN(n606) );
  XNOR2_X1 U514 ( .A(n402), .B(n658), .ZN(G75) );
  NAND2_X1 U515 ( .A1(n657), .A2(n733), .ZN(n402) );
  NAND2_X1 U516 ( .A1(n403), .A2(n413), .ZN(n412) );
  AND2_X1 U517 ( .A1(n591), .A2(n590), .ZN(n403) );
  XNOR2_X2 U518 ( .A(n404), .B(G469), .ZN(n559) );
  XNOR2_X1 U519 ( .A(n505), .B(n506), .ZN(n405) );
  NAND2_X1 U520 ( .A1(n406), .A2(n616), .ZN(n407) );
  NAND2_X1 U521 ( .A1(n421), .A2(n529), .ZN(n409) );
  NAND2_X1 U522 ( .A1(n410), .A2(n598), .ZN(n600) );
  XNOR2_X1 U523 ( .A(n412), .B(n411), .ZN(n410) );
  XNOR2_X1 U524 ( .A(n572), .B(n366), .ZN(n413) );
  NAND2_X1 U525 ( .A1(n626), .A2(n566), .ZN(n567) );
  NAND2_X1 U526 ( .A1(n421), .A2(n419), .ZN(n443) );
  INV_X1 U527 ( .A(n421), .ZN(n420) );
  XNOR2_X2 U528 ( .A(n425), .B(KEYINPUT0), .ZN(n529) );
  XNOR2_X1 U529 ( .A(n422), .B(n730), .ZN(n486) );
  INV_X1 U530 ( .A(n423), .ZN(n596) );
  NAND2_X1 U531 ( .A1(n423), .A2(n640), .ZN(n429) );
  XNOR2_X2 U532 ( .A(n466), .B(n360), .ZN(n423) );
  XNOR2_X1 U533 ( .A(n596), .B(KEYINPUT38), .ZN(n641) );
  NAND2_X1 U534 ( .A1(n584), .A2(n423), .ZN(n586) );
  XNOR2_X1 U535 ( .A(n424), .B(n489), .ZN(n434) );
  XNOR2_X2 U536 ( .A(n427), .B(G107), .ZN(n424) );
  NOR2_X2 U537 ( .A1(n578), .A2(n475), .ZN(n425) );
  NAND2_X1 U538 ( .A1(n428), .A2(n719), .ZN(n729) );
  XNOR2_X2 U539 ( .A(n533), .B(KEYINPUT35), .ZN(n741) );
  NAND2_X1 U540 ( .A1(n444), .A2(n573), .ZN(n530) );
  NAND2_X1 U541 ( .A1(n529), .A2(n437), .ZN(n498) );
  AND2_X1 U542 ( .A1(n568), .A2(n641), .ZN(n442) );
  INV_X1 U543 ( .A(KEYINPUT64), .ZN(n547) );
  INV_X1 U544 ( .A(KEYINPUT73), .ZN(n501) );
  XNOR2_X1 U545 ( .A(n502), .B(n501), .ZN(n503) );
  XNOR2_X1 U546 ( .A(n504), .B(n503), .ZN(n505) );
  INV_X1 U547 ( .A(KEYINPUT94), .ZN(n524) );
  BUF_X1 U548 ( .A(n616), .Z(n720) );
  NAND2_X1 U549 ( .A1(n563), .A2(n640), .ZN(n565) );
  NAND2_X1 U550 ( .A1(n587), .A2(n442), .ZN(n570) );
  XNOR2_X1 U551 ( .A(n707), .B(n710), .ZN(n711) );
  AND2_X1 U552 ( .A1(n656), .A2(n655), .ZN(n657) );
  INV_X1 U553 ( .A(KEYINPUT123), .ZN(n612) );
  XNOR2_X2 U554 ( .A(KEYINPUT67), .B(G131), .ZN(n482) );
  XNOR2_X1 U555 ( .A(n482), .B(n445), .ZN(n446) );
  NAND2_X1 U556 ( .A1(n480), .A2(G210), .ZN(n448) );
  XNOR2_X1 U557 ( .A(n448), .B(n447), .ZN(n450) );
  XNOR2_X1 U558 ( .A(KEYINPUT72), .B(KEYINPUT5), .ZN(n449) );
  XNOR2_X1 U559 ( .A(n450), .B(n449), .ZN(n454) );
  XNOR2_X1 U560 ( .A(KEYINPUT3), .B(G113), .ZN(n452) );
  INV_X1 U561 ( .A(n461), .ZN(n453) );
  XNOR2_X2 U562 ( .A(n455), .B(G472), .ZN(n536) );
  XNOR2_X1 U563 ( .A(KEYINPUT100), .B(KEYINPUT6), .ZN(n456) );
  XOR2_X1 U564 ( .A(KEYINPUT92), .B(KEYINPUT21), .Z(n460) );
  XOR2_X1 U565 ( .A(KEYINPUT20), .B(KEYINPUT91), .Z(n458) );
  NAND2_X1 U566 ( .A1(G234), .A2(n603), .ZN(n457) );
  XNOR2_X1 U567 ( .A(n458), .B(n457), .ZN(n515) );
  NAND2_X1 U568 ( .A1(n515), .A2(G221), .ZN(n459) );
  XNOR2_X1 U569 ( .A(n460), .B(n459), .ZN(n623) );
  XNOR2_X1 U570 ( .A(n623), .B(KEYINPUT93), .ZN(n523) );
  XOR2_X1 U571 ( .A(KEYINPUT68), .B(KEYINPUT85), .Z(n463) );
  NAND2_X1 U572 ( .A1(G224), .A2(n733), .ZN(n464) );
  NAND2_X1 U573 ( .A1(n676), .A2(n603), .ZN(n466) );
  NOR2_X1 U574 ( .A1(G237), .A2(G902), .ZN(n465) );
  XNOR2_X1 U575 ( .A(KEYINPUT71), .B(n465), .ZN(n467) );
  NAND2_X1 U576 ( .A1(n467), .A2(G214), .ZN(n640) );
  XOR2_X1 U577 ( .A(KEYINPUT69), .B(KEYINPUT14), .Z(n470) );
  XNOR2_X1 U578 ( .A(n470), .B(n469), .ZN(n472) );
  NAND2_X1 U579 ( .A1(n472), .A2(G952), .ZN(n471) );
  XNOR2_X1 U580 ( .A(n471), .B(KEYINPUT87), .ZN(n651) );
  NAND2_X1 U581 ( .A1(n651), .A2(n733), .ZN(n554) );
  INV_X1 U582 ( .A(n554), .ZN(n474) );
  NAND2_X1 U583 ( .A1(G902), .A2(n472), .ZN(n551) );
  XOR2_X1 U584 ( .A(KEYINPUT88), .B(G898), .Z(n723) );
  NAND2_X1 U585 ( .A1(G953), .A2(n723), .ZN(n719) );
  NOR2_X1 U586 ( .A1(n551), .A2(n719), .ZN(n473) );
  NOR2_X1 U587 ( .A1(n474), .A2(n473), .ZN(n475) );
  XNOR2_X1 U588 ( .A(n479), .B(n478), .ZN(n484) );
  NAND2_X1 U589 ( .A1(n480), .A2(G214), .ZN(n481) );
  XNOR2_X1 U590 ( .A(n482), .B(n481), .ZN(n483) );
  XNOR2_X1 U591 ( .A(n484), .B(n483), .ZN(n485) );
  XNOR2_X1 U592 ( .A(n486), .B(n485), .ZN(n669) );
  XNOR2_X1 U593 ( .A(KEYINPUT13), .B(KEYINPUT95), .ZN(n487) );
  INV_X1 U594 ( .A(n521), .ZN(n532) );
  XOR2_X1 U595 ( .A(KEYINPUT96), .B(KEYINPUT97), .Z(n489) );
  NAND2_X1 U596 ( .A1(G234), .A2(n733), .ZN(n488) );
  XOR2_X1 U597 ( .A(KEYINPUT9), .B(KEYINPUT7), .Z(n491) );
  XNOR2_X1 U598 ( .A(n491), .B(n490), .ZN(n492) );
  XNOR2_X1 U599 ( .A(n493), .B(n492), .ZN(n494) );
  NOR2_X1 U600 ( .A1(n608), .A2(G902), .ZN(n496) );
  XNOR2_X1 U601 ( .A(G478), .B(n496), .ZN(n531) );
  NAND2_X1 U602 ( .A1(n532), .A2(n531), .ZN(n643) );
  INV_X1 U603 ( .A(n643), .ZN(n497) );
  XNOR2_X1 U604 ( .A(n500), .B(n499), .ZN(n504) );
  NAND2_X1 U605 ( .A1(G227), .A2(n733), .ZN(n502) );
  INV_X1 U606 ( .A(G902), .ZN(n508) );
  XOR2_X1 U607 ( .A(KEYINPUT1), .B(KEYINPUT65), .Z(n509) );
  XOR2_X1 U608 ( .A(KEYINPUT24), .B(KEYINPUT23), .Z(n511) );
  XNOR2_X1 U609 ( .A(n511), .B(n510), .ZN(n514) );
  NOR2_X1 U610 ( .A1(G902), .A2(n715), .ZN(n519) );
  XOR2_X1 U611 ( .A(KEYINPUT90), .B(KEYINPUT25), .Z(n517) );
  NAND2_X1 U612 ( .A1(n515), .A2(G217), .ZN(n516) );
  XNOR2_X1 U613 ( .A(n517), .B(n516), .ZN(n518) );
  XNOR2_X1 U614 ( .A(n519), .B(n518), .ZN(n537) );
  XNOR2_X1 U615 ( .A(KEYINPUT101), .B(n537), .ZN(n622) );
  OR2_X1 U616 ( .A1(n531), .A2(n521), .ZN(n522) );
  XNOR2_X1 U617 ( .A(KEYINPUT99), .B(n522), .ZN(n703) );
  NOR2_X1 U618 ( .A1(n701), .A2(n703), .ZN(n645) );
  INV_X1 U619 ( .A(n536), .ZN(n632) );
  NAND2_X1 U620 ( .A1(n444), .A2(n632), .ZN(n525) );
  NAND2_X1 U621 ( .A1(n636), .A2(n529), .ZN(n526) );
  XNOR2_X1 U622 ( .A(n526), .B(KEYINPUT31), .ZN(n700) );
  NAND2_X1 U623 ( .A1(n626), .A2(n536), .ZN(n527) );
  INV_X1 U624 ( .A(n559), .ZN(n585) );
  NOR2_X1 U625 ( .A1(n527), .A2(n585), .ZN(n528) );
  AND2_X1 U626 ( .A1(n529), .A2(n528), .ZN(n688) );
  NOR2_X1 U627 ( .A1(n532), .A2(n531), .ZN(n582) );
  NAND2_X1 U628 ( .A1(KEYINPUT44), .A2(n741), .ZN(n534) );
  INV_X1 U629 ( .A(n537), .ZN(n556) );
  NOR2_X1 U630 ( .A1(n563), .A2(n556), .ZN(n538) );
  INV_X1 U631 ( .A(n357), .ZN(n543) );
  OR2_X1 U632 ( .A1(n573), .A2(n622), .ZN(n542) );
  NOR2_X1 U633 ( .A1(n543), .A2(n542), .ZN(n544) );
  XNOR2_X1 U634 ( .A(KEYINPUT32), .B(n545), .ZN(n746) );
  INV_X1 U635 ( .A(KEYINPUT44), .ZN(n546) );
  INV_X1 U636 ( .A(n603), .ZN(n548) );
  NAND2_X1 U637 ( .A1(n641), .A2(n640), .ZN(n644) );
  NOR2_X1 U638 ( .A1(n644), .A2(n643), .ZN(n550) );
  XNOR2_X1 U639 ( .A(KEYINPUT41), .B(KEYINPUT108), .ZN(n549) );
  XNOR2_X1 U640 ( .A(n550), .B(n549), .ZN(n653) );
  NOR2_X1 U641 ( .A1(G900), .A2(n551), .ZN(n552) );
  NAND2_X1 U642 ( .A1(n552), .A2(G953), .ZN(n553) );
  NAND2_X1 U643 ( .A1(n554), .A2(n553), .ZN(n566) );
  NAND2_X1 U644 ( .A1(n623), .A2(n566), .ZN(n555) );
  NOR2_X1 U645 ( .A1(n556), .A2(n555), .ZN(n574) );
  NAND2_X1 U646 ( .A1(n563), .A2(n574), .ZN(n558) );
  INV_X1 U647 ( .A(KEYINPUT28), .ZN(n557) );
  XNOR2_X1 U648 ( .A(n558), .B(n557), .ZN(n560) );
  NAND2_X1 U649 ( .A1(n560), .A2(n559), .ZN(n579) );
  NOR2_X1 U650 ( .A1(n653), .A2(n579), .ZN(n562) );
  INV_X1 U651 ( .A(KEYINPUT42), .ZN(n561) );
  XNOR2_X1 U652 ( .A(n562), .B(n561), .ZN(n747) );
  XNOR2_X1 U653 ( .A(KEYINPUT107), .B(KEYINPUT30), .ZN(n564) );
  XNOR2_X1 U654 ( .A(n565), .B(n564), .ZN(n587) );
  NOR2_X1 U655 ( .A1(n567), .A2(n585), .ZN(n568) );
  INV_X1 U656 ( .A(KEYINPUT39), .ZN(n569) );
  XNOR2_X1 U657 ( .A(n570), .B(n569), .ZN(n601) );
  INV_X1 U658 ( .A(n701), .ZN(n697) );
  XNOR2_X2 U659 ( .A(n571), .B(KEYINPUT40), .ZN(n615) );
  NAND2_X1 U660 ( .A1(n747), .A2(n615), .ZN(n572) );
  XNOR2_X1 U661 ( .A(KEYINPUT36), .B(n575), .ZN(n576) );
  NAND2_X1 U662 ( .A1(n576), .A2(n357), .ZN(n577) );
  XNOR2_X2 U663 ( .A(n577), .B(KEYINPUT109), .ZN(n743) );
  XNOR2_X1 U664 ( .A(n743), .B(KEYINPUT83), .ZN(n591) );
  OR2_X1 U665 ( .A1(n579), .A2(n578), .ZN(n696) );
  NOR2_X1 U666 ( .A1(n696), .A2(n645), .ZN(n581) );
  INV_X1 U667 ( .A(KEYINPUT47), .ZN(n580) );
  XNOR2_X1 U668 ( .A(n581), .B(n580), .ZN(n589) );
  AND2_X1 U669 ( .A1(n583), .A2(n582), .ZN(n584) );
  NOR2_X1 U670 ( .A1(n586), .A2(n585), .ZN(n588) );
  AND2_X1 U671 ( .A1(n588), .A2(n587), .ZN(n694) );
  NOR2_X1 U672 ( .A1(n589), .A2(n694), .ZN(n590) );
  NOR2_X1 U673 ( .A1(n357), .A2(n592), .ZN(n593) );
  AND2_X1 U674 ( .A1(n593), .A2(n640), .ZN(n595) );
  XOR2_X1 U675 ( .A(KEYINPUT106), .B(KEYINPUT43), .Z(n594) );
  XNOR2_X1 U676 ( .A(n595), .B(n594), .ZN(n597) );
  AND2_X1 U677 ( .A1(n597), .A2(n596), .ZN(n705) );
  INV_X1 U678 ( .A(n705), .ZN(n598) );
  INV_X1 U679 ( .A(KEYINPUT80), .ZN(n599) );
  INV_X1 U680 ( .A(n703), .ZN(n691) );
  OR2_X1 U681 ( .A1(n601), .A2(n691), .ZN(n614) );
  INV_X1 U682 ( .A(KEYINPUT2), .ZN(n602) );
  OR2_X1 U683 ( .A1(n603), .A2(n602), .ZN(n604) );
  XNOR2_X1 U684 ( .A(n604), .B(KEYINPUT66), .ZN(n605) );
  NAND2_X1 U685 ( .A1(n706), .A2(G478), .ZN(n609) );
  XNOR2_X1 U686 ( .A(n609), .B(n608), .ZN(n611) );
  INV_X1 U687 ( .A(G952), .ZN(n610) );
  AND2_X1 U688 ( .A1(n610), .A2(G953), .ZN(n718) );
  NOR2_X2 U689 ( .A1(n611), .A2(n718), .ZN(n613) );
  XNOR2_X1 U690 ( .A(n613), .B(n612), .ZN(G63) );
  XNOR2_X1 U691 ( .A(n614), .B(G134), .ZN(G36) );
  XNOR2_X1 U692 ( .A(n615), .B(G131), .ZN(G33) );
  INV_X1 U693 ( .A(KEYINPUT53), .ZN(n658) );
  XNOR2_X1 U694 ( .A(n617), .B(KEYINPUT77), .ZN(n619) );
  OR2_X1 U695 ( .A1(n732), .A2(KEYINPUT2), .ZN(n618) );
  AND2_X1 U696 ( .A1(n619), .A2(n618), .ZN(n620) );
  NOR2_X1 U697 ( .A1(n623), .A2(n622), .ZN(n624) );
  XNOR2_X1 U698 ( .A(KEYINPUT49), .B(n624), .ZN(n631) );
  NOR2_X1 U699 ( .A1(n626), .A2(n357), .ZN(n628) );
  XNOR2_X1 U700 ( .A(KEYINPUT118), .B(KEYINPUT50), .ZN(n627) );
  XNOR2_X1 U701 ( .A(n628), .B(n627), .ZN(n629) );
  XNOR2_X1 U702 ( .A(KEYINPUT117), .B(n629), .ZN(n630) );
  NAND2_X1 U703 ( .A1(n631), .A2(n630), .ZN(n633) );
  NOR2_X1 U704 ( .A1(n633), .A2(n632), .ZN(n634) );
  XOR2_X1 U705 ( .A(KEYINPUT119), .B(n634), .Z(n635) );
  NOR2_X1 U706 ( .A1(n636), .A2(n635), .ZN(n637) );
  XOR2_X1 U707 ( .A(KEYINPUT51), .B(n637), .Z(n638) );
  NOR2_X1 U708 ( .A1(n653), .A2(n638), .ZN(n639) );
  XNOR2_X1 U709 ( .A(n639), .B(KEYINPUT120), .ZN(n649) );
  NOR2_X1 U710 ( .A1(n641), .A2(n640), .ZN(n642) );
  NOR2_X1 U711 ( .A1(n643), .A2(n642), .ZN(n647) );
  NOR2_X1 U712 ( .A1(n645), .A2(n644), .ZN(n646) );
  NOR2_X1 U713 ( .A1(n647), .A2(n646), .ZN(n648) );
  NOR2_X1 U714 ( .A1(n649), .A2(n363), .ZN(n650) );
  XOR2_X1 U715 ( .A(KEYINPUT52), .B(n650), .Z(n652) );
  NAND2_X1 U716 ( .A1(n652), .A2(n651), .ZN(n654) );
  NAND2_X1 U717 ( .A1(n660), .A2(n659), .ZN(n662) );
  INV_X1 U718 ( .A(G472), .ZN(n661) );
  NOR2_X1 U719 ( .A1(n662), .A2(n661), .ZN(n665) );
  XOR2_X1 U720 ( .A(KEYINPUT62), .B(n663), .Z(n664) );
  XNOR2_X1 U721 ( .A(n665), .B(n664), .ZN(n666) );
  NOR2_X1 U722 ( .A1(n666), .A2(n718), .ZN(n668) );
  XOR2_X1 U723 ( .A(KEYINPUT86), .B(KEYINPUT63), .Z(n667) );
  XNOR2_X1 U724 ( .A(n668), .B(n667), .ZN(G57) );
  NAND2_X1 U725 ( .A1(n706), .A2(G475), .ZN(n671) );
  XOR2_X1 U726 ( .A(n669), .B(KEYINPUT59), .Z(n670) );
  XNOR2_X1 U727 ( .A(n671), .B(n670), .ZN(n672) );
  NOR2_X2 U728 ( .A1(n672), .A2(n718), .ZN(n673) );
  XNOR2_X1 U729 ( .A(n673), .B(KEYINPUT60), .ZN(G60) );
  NAND2_X1 U730 ( .A1(n706), .A2(G210), .ZN(n678) );
  XNOR2_X1 U731 ( .A(KEYINPUT76), .B(KEYINPUT54), .ZN(n674) );
  XNOR2_X1 U732 ( .A(n674), .B(KEYINPUT55), .ZN(n675) );
  XNOR2_X1 U733 ( .A(n676), .B(n675), .ZN(n677) );
  XNOR2_X1 U734 ( .A(n678), .B(n677), .ZN(n679) );
  NOR2_X2 U735 ( .A1(n679), .A2(n718), .ZN(n681) );
  XOR2_X1 U736 ( .A(KEYINPUT81), .B(KEYINPUT56), .Z(n680) );
  XNOR2_X1 U737 ( .A(n681), .B(n680), .ZN(G51) );
  XOR2_X1 U738 ( .A(G101), .B(n682), .Z(G3) );
  NAND2_X1 U739 ( .A1(n701), .A2(n688), .ZN(n683) );
  XNOR2_X1 U740 ( .A(n683), .B(KEYINPUT110), .ZN(n684) );
  XNOR2_X1 U741 ( .A(G104), .B(n684), .ZN(G6) );
  XOR2_X1 U742 ( .A(KEYINPUT27), .B(KEYINPUT112), .Z(n686) );
  XNOR2_X1 U743 ( .A(G107), .B(KEYINPUT111), .ZN(n685) );
  XNOR2_X1 U744 ( .A(n686), .B(n685), .ZN(n687) );
  XOR2_X1 U745 ( .A(KEYINPUT26), .B(n687), .Z(n690) );
  NAND2_X1 U746 ( .A1(n688), .A2(n703), .ZN(n689) );
  XNOR2_X1 U747 ( .A(n690), .B(n689), .ZN(G9) );
  NOR2_X1 U748 ( .A1(n691), .A2(n696), .ZN(n693) );
  XNOR2_X1 U749 ( .A(G128), .B(KEYINPUT29), .ZN(n692) );
  XNOR2_X1 U750 ( .A(n693), .B(n692), .ZN(G30) );
  XOR2_X1 U751 ( .A(G143), .B(n694), .Z(n695) );
  XNOR2_X1 U752 ( .A(KEYINPUT114), .B(n695), .ZN(G45) );
  NOR2_X1 U753 ( .A1(n697), .A2(n696), .ZN(n699) );
  XNOR2_X1 U754 ( .A(G146), .B(KEYINPUT115), .ZN(n698) );
  XNOR2_X1 U755 ( .A(n699), .B(n698), .ZN(G48) );
  NAND2_X1 U756 ( .A1(n701), .A2(n700), .ZN(n702) );
  XNOR2_X1 U757 ( .A(n702), .B(G113), .ZN(G15) );
  NAND2_X1 U758 ( .A1(n700), .A2(n703), .ZN(n704) );
  XNOR2_X1 U759 ( .A(n704), .B(G116), .ZN(G18) );
  XOR2_X1 U760 ( .A(G140), .B(n705), .Z(G42) );
  NAND2_X1 U761 ( .A1(n714), .A2(G469), .ZN(n712) );
  XOR2_X1 U762 ( .A(KEYINPUT58), .B(KEYINPUT57), .Z(n709) );
  XNOR2_X1 U763 ( .A(KEYINPUT122), .B(KEYINPUT121), .ZN(n708) );
  XNOR2_X1 U764 ( .A(n709), .B(n708), .ZN(n710) );
  NOR2_X1 U765 ( .A1(n718), .A2(n713), .ZN(G54) );
  NAND2_X1 U766 ( .A1(n714), .A2(G217), .ZN(n716) );
  XNOR2_X1 U767 ( .A(n716), .B(n715), .ZN(n717) );
  NOR2_X1 U768 ( .A1(n718), .A2(n717), .ZN(G66) );
  NAND2_X1 U769 ( .A1(n733), .A2(n720), .ZN(n726) );
  NAND2_X1 U770 ( .A1(G953), .A2(G224), .ZN(n721) );
  XOR2_X1 U771 ( .A(KEYINPUT61), .B(n721), .Z(n722) );
  NOR2_X1 U772 ( .A1(n723), .A2(n722), .ZN(n724) );
  XOR2_X1 U773 ( .A(KEYINPUT124), .B(n724), .Z(n725) );
  NAND2_X1 U774 ( .A1(n726), .A2(n725), .ZN(n727) );
  XNOR2_X1 U775 ( .A(n727), .B(KEYINPUT125), .ZN(n728) );
  XNOR2_X1 U776 ( .A(n729), .B(n728), .ZN(G69) );
  XOR2_X1 U777 ( .A(n731), .B(n730), .Z(n735) );
  XNOR2_X1 U778 ( .A(n732), .B(n735), .ZN(n734) );
  NAND2_X1 U779 ( .A1(n734), .A2(n733), .ZN(n740) );
  XOR2_X1 U780 ( .A(G227), .B(n735), .Z(n736) );
  NAND2_X1 U781 ( .A1(n736), .A2(G900), .ZN(n737) );
  XNOR2_X1 U782 ( .A(KEYINPUT126), .B(n737), .ZN(n738) );
  NAND2_X1 U783 ( .A1(n738), .A2(G953), .ZN(n739) );
  NAND2_X1 U784 ( .A1(n740), .A2(n739), .ZN(G72) );
  XOR2_X1 U785 ( .A(n741), .B(G122), .Z(G24) );
  XNOR2_X1 U786 ( .A(G110), .B(KEYINPUT113), .ZN(n742) );
  XNOR2_X1 U787 ( .A(n743), .B(KEYINPUT116), .ZN(n744) );
  XNOR2_X1 U788 ( .A(n744), .B(KEYINPUT37), .ZN(n745) );
  XNOR2_X1 U789 ( .A(G125), .B(n745), .ZN(G27) );
  XOR2_X1 U790 ( .A(n746), .B(G119), .Z(G21) );
  XNOR2_X1 U791 ( .A(G137), .B(n747), .ZN(G39) );
endmodule

