//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 0 0 0 1 0 0 1 0 0 0 0 0 0 0 0 1 0 0 1 0 1 0 0 0 1 0 0 1 1 0 1 1 0 0 1 0 1 1 0 0 0 0 0 0 0 1 0 1 1 0 1 1 1 1 0 1 0 0 0 1 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:37:50 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n587, new_n588, new_n589, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n597, new_n598,
    new_n599, new_n600, new_n601, new_n602, new_n603, new_n604, new_n605,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n986, new_n987, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1018, new_n1019, new_n1020, new_n1021, new_n1022,
    new_n1023, new_n1024, new_n1025, new_n1026, new_n1027, new_n1028,
    new_n1029, new_n1030, new_n1031, new_n1032, new_n1033, new_n1034,
    new_n1035, new_n1036, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1051, new_n1052, new_n1053,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1108,
    new_n1109, new_n1110, new_n1111, new_n1112, new_n1113, new_n1114,
    new_n1115, new_n1116, new_n1117, new_n1118, new_n1119, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1182, new_n1183, new_n1184, new_n1185, new_n1186, new_n1187,
    new_n1188, new_n1189, new_n1190, new_n1191, new_n1192, new_n1193,
    new_n1194, new_n1195, new_n1196, new_n1197, new_n1198, new_n1199,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1207, new_n1208,
    new_n1209, new_n1210, new_n1211, new_n1212, new_n1213, new_n1214,
    new_n1215, new_n1216, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1260, new_n1261, new_n1262, new_n1263,
    new_n1264, new_n1265, new_n1266, new_n1267, new_n1268, new_n1269,
    new_n1270, new_n1271;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  AOI22_X1  g0005(.A1(G50), .A2(G226), .B1(G77), .B2(G244), .ZN(new_n206));
  INV_X1    g0006(.A(G116), .ZN(new_n207));
  INV_X1    g0007(.A(G270), .ZN(new_n208));
  OAI21_X1  g0008(.A(new_n206), .B1(new_n207), .B2(new_n208), .ZN(new_n209));
  AOI22_X1  g0009(.A1(G87), .A2(G250), .B1(G107), .B2(G264), .ZN(new_n210));
  INV_X1    g0010(.A(G68), .ZN(new_n211));
  INV_X1    g0011(.A(G238), .ZN(new_n212));
  INV_X1    g0012(.A(G97), .ZN(new_n213));
  INV_X1    g0013(.A(G257), .ZN(new_n214));
  OAI221_X1 g0014(.A(new_n210), .B1(new_n211), .B2(new_n212), .C1(new_n213), .C2(new_n214), .ZN(new_n215));
  AOI211_X1 g0015(.A(new_n209), .B(new_n215), .C1(G58), .C2(G232), .ZN(new_n216));
  INV_X1    g0016(.A(G1), .ZN(new_n217));
  INV_X1    g0017(.A(G20), .ZN(new_n218));
  NOR2_X1   g0018(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  NOR2_X1   g0019(.A1(new_n216), .A2(new_n219), .ZN(new_n220));
  XOR2_X1   g0020(.A(new_n220), .B(KEYINPUT1), .Z(new_n221));
  INV_X1    g0021(.A(new_n201), .ZN(new_n222));
  NAND2_X1  g0022(.A1(new_n222), .A2(G50), .ZN(new_n223));
  INV_X1    g0023(.A(G13), .ZN(new_n224));
  NOR2_X1   g0024(.A1(new_n217), .A2(new_n224), .ZN(new_n225));
  INV_X1    g0025(.A(new_n225), .ZN(new_n226));
  NOR3_X1   g0026(.A1(new_n223), .A2(new_n226), .A3(new_n218), .ZN(new_n227));
  NAND2_X1  g0027(.A1(new_n219), .A2(new_n224), .ZN(new_n228));
  INV_X1    g0028(.A(new_n228), .ZN(new_n229));
  OAI211_X1 g0029(.A(new_n229), .B(G250), .C1(G257), .C2(G264), .ZN(new_n230));
  XOR2_X1   g0030(.A(new_n230), .B(KEYINPUT0), .Z(new_n231));
  NOR3_X1   g0031(.A1(new_n221), .A2(new_n227), .A3(new_n231), .ZN(G361));
  XOR2_X1   g0032(.A(KEYINPUT64), .B(KEYINPUT2), .Z(new_n233));
  XNOR2_X1  g0033(.A(G238), .B(G244), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XNOR2_X1  g0035(.A(G226), .B(G232), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XOR2_X1   g0037(.A(new_n237), .B(KEYINPUT65), .Z(new_n238));
  XNOR2_X1  g0038(.A(G250), .B(G257), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n239), .B(G264), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n240), .B(new_n208), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n238), .B(new_n241), .ZN(G358));
  XNOR2_X1  g0042(.A(G50), .B(G68), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n243), .B(G58), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n244), .B(G77), .ZN(new_n245));
  XNOR2_X1  g0045(.A(G87), .B(G97), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n246), .B(G107), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n247), .B(new_n207), .ZN(new_n248));
  XOR2_X1   g0048(.A(new_n245), .B(new_n248), .Z(G351));
  NAND2_X1  g0049(.A1(KEYINPUT71), .A2(KEYINPUT10), .ZN(new_n250));
  OR2_X1    g0050(.A1(KEYINPUT3), .A2(G33), .ZN(new_n251));
  NAND2_X1  g0051(.A1(KEYINPUT3), .A2(G33), .ZN(new_n252));
  NAND2_X1  g0052(.A1(new_n251), .A2(new_n252), .ZN(new_n253));
  AND2_X1   g0053(.A1(new_n253), .A2(G1698), .ZN(new_n254));
  XNOR2_X1  g0054(.A(KEYINPUT66), .B(G1698), .ZN(new_n255));
  NAND3_X1  g0055(.A1(new_n253), .A2(new_n255), .A3(G222), .ZN(new_n256));
  AOI22_X1  g0056(.A1(new_n254), .A2(G223), .B1(new_n256), .B2(KEYINPUT67), .ZN(new_n257));
  INV_X1    g0057(.A(G77), .ZN(new_n258));
  OAI221_X1 g0058(.A(new_n257), .B1(KEYINPUT67), .B2(new_n256), .C1(new_n258), .C2(new_n253), .ZN(new_n259));
  INV_X1    g0059(.A(G33), .ZN(new_n260));
  INV_X1    g0060(.A(G41), .ZN(new_n261));
  OAI211_X1 g0061(.A(G1), .B(G13), .C1(new_n260), .C2(new_n261), .ZN(new_n262));
  INV_X1    g0062(.A(new_n262), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n259), .A2(new_n263), .ZN(new_n264));
  OAI21_X1  g0064(.A(new_n217), .B1(G41), .B2(G45), .ZN(new_n265));
  INV_X1    g0065(.A(G274), .ZN(new_n266));
  NOR2_X1   g0066(.A1(new_n265), .A2(new_n266), .ZN(new_n267));
  INV_X1    g0067(.A(new_n267), .ZN(new_n268));
  AND2_X1   g0068(.A1(new_n262), .A2(new_n265), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n269), .A2(G226), .ZN(new_n270));
  NAND3_X1  g0070(.A1(new_n264), .A2(new_n268), .A3(new_n270), .ZN(new_n271));
  INV_X1    g0071(.A(G190), .ZN(new_n272));
  OAI21_X1  g0072(.A(new_n250), .B1(new_n271), .B2(new_n272), .ZN(new_n273));
  INV_X1    g0073(.A(KEYINPUT70), .ZN(new_n274));
  AOI21_X1  g0074(.A(new_n274), .B1(new_n271), .B2(G200), .ZN(new_n275));
  NOR2_X1   g0075(.A1(new_n273), .A2(new_n275), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n203), .A2(G20), .ZN(new_n277));
  INV_X1    g0077(.A(G150), .ZN(new_n278));
  NOR2_X1   g0078(.A1(G20), .A2(G33), .ZN(new_n279));
  INV_X1    g0079(.A(new_n279), .ZN(new_n280));
  INV_X1    g0080(.A(KEYINPUT68), .ZN(new_n281));
  OAI21_X1  g0081(.A(new_n281), .B1(new_n260), .B2(G20), .ZN(new_n282));
  NAND3_X1  g0082(.A1(new_n218), .A2(KEYINPUT68), .A3(G33), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  XNOR2_X1  g0084(.A(KEYINPUT8), .B(G58), .ZN(new_n285));
  OAI221_X1 g0085(.A(new_n277), .B1(new_n278), .B2(new_n280), .C1(new_n284), .C2(new_n285), .ZN(new_n286));
  AOI21_X1  g0086(.A(new_n225), .B1(G33), .B2(new_n219), .ZN(new_n287));
  INV_X1    g0087(.A(new_n287), .ZN(new_n288));
  NAND3_X1  g0088(.A1(new_n217), .A2(G13), .A3(G20), .ZN(new_n289));
  INV_X1    g0089(.A(new_n289), .ZN(new_n290));
  AOI22_X1  g0090(.A1(new_n286), .A2(new_n288), .B1(new_n202), .B2(new_n290), .ZN(new_n291));
  OAI21_X1  g0091(.A(new_n287), .B1(G1), .B2(new_n218), .ZN(new_n292));
  OAI21_X1  g0092(.A(new_n291), .B1(new_n202), .B2(new_n292), .ZN(new_n293));
  XNOR2_X1  g0093(.A(new_n293), .B(KEYINPUT9), .ZN(new_n294));
  NAND3_X1  g0094(.A1(new_n271), .A2(new_n274), .A3(G200), .ZN(new_n295));
  NAND3_X1  g0095(.A1(new_n276), .A2(new_n294), .A3(new_n295), .ZN(new_n296));
  NOR2_X1   g0096(.A1(KEYINPUT71), .A2(KEYINPUT10), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n296), .A2(new_n297), .ZN(new_n298));
  INV_X1    g0098(.A(new_n297), .ZN(new_n299));
  NAND4_X1  g0099(.A1(new_n276), .A2(new_n299), .A3(new_n294), .A4(new_n295), .ZN(new_n300));
  INV_X1    g0100(.A(G169), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n271), .A2(new_n301), .ZN(new_n302));
  XOR2_X1   g0102(.A(KEYINPUT69), .B(G179), .Z(new_n303));
  INV_X1    g0103(.A(new_n303), .ZN(new_n304));
  OAI211_X1 g0104(.A(new_n302), .B(new_n293), .C1(new_n304), .C2(new_n271), .ZN(new_n305));
  NAND3_X1  g0105(.A1(new_n298), .A2(new_n300), .A3(new_n305), .ZN(new_n306));
  INV_X1    g0106(.A(KEYINPUT14), .ZN(new_n307));
  AOI22_X1  g0107(.A1(new_n255), .A2(G226), .B1(G232), .B2(G1698), .ZN(new_n308));
  AND2_X1   g0108(.A1(KEYINPUT3), .A2(G33), .ZN(new_n309));
  NOR2_X1   g0109(.A1(KEYINPUT3), .A2(G33), .ZN(new_n310));
  NOR2_X1   g0110(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  OAI22_X1  g0111(.A1(new_n308), .A2(new_n311), .B1(new_n260), .B2(new_n213), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n312), .A2(new_n263), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n269), .A2(G238), .ZN(new_n314));
  NAND3_X1  g0114(.A1(new_n313), .A2(new_n268), .A3(new_n314), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n315), .A2(KEYINPUT13), .ZN(new_n316));
  INV_X1    g0116(.A(KEYINPUT13), .ZN(new_n317));
  NAND4_X1  g0117(.A1(new_n313), .A2(new_n317), .A3(new_n268), .A4(new_n314), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n316), .A2(new_n318), .ZN(new_n319));
  AOI21_X1  g0119(.A(new_n307), .B1(new_n319), .B2(G169), .ZN(new_n320));
  AOI211_X1 g0120(.A(KEYINPUT14), .B(new_n301), .C1(new_n316), .C2(new_n318), .ZN(new_n321));
  INV_X1    g0121(.A(G179), .ZN(new_n322));
  NOR2_X1   g0122(.A1(new_n319), .A2(new_n322), .ZN(new_n323));
  NOR3_X1   g0123(.A1(new_n320), .A2(new_n321), .A3(new_n323), .ZN(new_n324));
  INV_X1    g0124(.A(new_n324), .ZN(new_n325));
  OAI22_X1  g0125(.A1(new_n284), .A2(new_n258), .B1(new_n202), .B2(new_n280), .ZN(new_n326));
  NOR2_X1   g0126(.A1(new_n218), .A2(G68), .ZN(new_n327));
  OAI21_X1  g0127(.A(new_n288), .B1(new_n326), .B2(new_n327), .ZN(new_n328));
  INV_X1    g0128(.A(KEYINPUT11), .ZN(new_n329));
  OAI22_X1  g0129(.A1(new_n328), .A2(new_n329), .B1(new_n211), .B2(new_n292), .ZN(new_n330));
  AND2_X1   g0130(.A1(new_n328), .A2(new_n329), .ZN(new_n331));
  NOR2_X1   g0131(.A1(new_n224), .A2(G1), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n327), .A2(new_n332), .ZN(new_n333));
  XOR2_X1   g0133(.A(new_n333), .B(KEYINPUT12), .Z(new_n334));
  OR3_X1    g0134(.A1(new_n330), .A2(new_n331), .A3(new_n334), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n325), .A2(new_n335), .ZN(new_n336));
  AOI21_X1  g0136(.A(new_n335), .B1(G200), .B2(new_n319), .ZN(new_n337));
  OAI21_X1  g0137(.A(new_n337), .B1(new_n272), .B2(new_n319), .ZN(new_n338));
  NAND2_X1  g0138(.A1(G20), .A2(G77), .ZN(new_n339));
  XNOR2_X1  g0139(.A(KEYINPUT15), .B(G87), .ZN(new_n340));
  OAI221_X1 g0140(.A(new_n339), .B1(new_n285), .B2(new_n280), .C1(new_n284), .C2(new_n340), .ZN(new_n341));
  AOI22_X1  g0141(.A1(new_n341), .A2(new_n288), .B1(new_n258), .B2(new_n290), .ZN(new_n342));
  OAI21_X1  g0142(.A(new_n342), .B1(new_n258), .B2(new_n292), .ZN(new_n343));
  AOI22_X1  g0143(.A1(new_n254), .A2(G238), .B1(G107), .B2(new_n311), .ZN(new_n344));
  INV_X1    g0144(.A(G232), .ZN(new_n345));
  AND2_X1   g0145(.A1(KEYINPUT66), .A2(G1698), .ZN(new_n346));
  NOR2_X1   g0146(.A1(KEYINPUT66), .A2(G1698), .ZN(new_n347));
  OAI22_X1  g0147(.A1(new_n309), .A2(new_n310), .B1(new_n346), .B2(new_n347), .ZN(new_n348));
  OAI21_X1  g0148(.A(new_n344), .B1(new_n345), .B2(new_n348), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n349), .A2(new_n263), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n269), .A2(G244), .ZN(new_n351));
  NAND3_X1  g0151(.A1(new_n350), .A2(new_n268), .A3(new_n351), .ZN(new_n352));
  AOI21_X1  g0152(.A(new_n343), .B1(new_n352), .B2(G200), .ZN(new_n353));
  OAI21_X1  g0153(.A(new_n353), .B1(new_n272), .B2(new_n352), .ZN(new_n354));
  NAND3_X1  g0154(.A1(new_n336), .A2(new_n338), .A3(new_n354), .ZN(new_n355));
  INV_X1    g0155(.A(KEYINPUT16), .ZN(new_n356));
  NAND2_X1  g0156(.A1(G58), .A2(G68), .ZN(new_n357));
  AOI21_X1  g0157(.A(new_n218), .B1(new_n222), .B2(new_n357), .ZN(new_n358));
  NAND3_X1  g0158(.A1(new_n251), .A2(new_n218), .A3(new_n252), .ZN(new_n359));
  INV_X1    g0159(.A(KEYINPUT7), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n359), .A2(new_n360), .ZN(new_n361));
  NAND4_X1  g0161(.A1(new_n251), .A2(KEYINPUT7), .A3(new_n218), .A4(new_n252), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n361), .A2(new_n362), .ZN(new_n363));
  AOI21_X1  g0163(.A(new_n358), .B1(new_n363), .B2(G68), .ZN(new_n364));
  INV_X1    g0164(.A(G159), .ZN(new_n365));
  NOR2_X1   g0165(.A1(new_n280), .A2(new_n365), .ZN(new_n366));
  INV_X1    g0166(.A(new_n366), .ZN(new_n367));
  AOI21_X1  g0167(.A(new_n356), .B1(new_n364), .B2(new_n367), .ZN(new_n368));
  AOI21_X1  g0168(.A(new_n211), .B1(new_n361), .B2(new_n362), .ZN(new_n369));
  NOR4_X1   g0169(.A1(new_n369), .A2(KEYINPUT16), .A3(new_n366), .A4(new_n358), .ZN(new_n370));
  OAI21_X1  g0170(.A(new_n288), .B1(new_n368), .B2(new_n370), .ZN(new_n371));
  NOR2_X1   g0171(.A1(new_n292), .A2(new_n285), .ZN(new_n372));
  INV_X1    g0172(.A(new_n372), .ZN(new_n373));
  INV_X1    g0173(.A(new_n285), .ZN(new_n374));
  NOR2_X1   g0174(.A1(new_n374), .A2(new_n289), .ZN(new_n375));
  INV_X1    g0175(.A(new_n375), .ZN(new_n376));
  NAND3_X1  g0176(.A1(new_n371), .A2(new_n373), .A3(new_n376), .ZN(new_n377));
  NAND3_X1  g0177(.A1(new_n253), .A2(new_n255), .A3(G223), .ZN(new_n378));
  NAND3_X1  g0178(.A1(new_n253), .A2(G226), .A3(G1698), .ZN(new_n379));
  NAND2_X1  g0179(.A1(G33), .A2(G87), .ZN(new_n380));
  NAND3_X1  g0180(.A1(new_n378), .A2(new_n379), .A3(new_n380), .ZN(new_n381));
  INV_X1    g0181(.A(KEYINPUT72), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n381), .A2(new_n382), .ZN(new_n383));
  NAND4_X1  g0183(.A1(new_n378), .A2(new_n379), .A3(KEYINPUT72), .A4(new_n380), .ZN(new_n384));
  NAND3_X1  g0184(.A1(new_n383), .A2(new_n263), .A3(new_n384), .ZN(new_n385));
  AOI21_X1  g0185(.A(new_n267), .B1(new_n269), .B2(G232), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n385), .A2(new_n386), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n387), .A2(new_n301), .ZN(new_n388));
  NAND3_X1  g0188(.A1(new_n385), .A2(new_n386), .A3(new_n303), .ZN(new_n389));
  NAND3_X1  g0189(.A1(new_n377), .A2(new_n388), .A3(new_n389), .ZN(new_n390));
  INV_X1    g0190(.A(KEYINPUT18), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n390), .A2(new_n391), .ZN(new_n392));
  NAND4_X1  g0192(.A1(new_n377), .A2(KEYINPUT18), .A3(new_n388), .A4(new_n389), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n392), .A2(new_n393), .ZN(new_n394));
  AOI21_X1  g0194(.A(KEYINPUT7), .B1(new_n311), .B2(new_n218), .ZN(new_n395));
  NOR4_X1   g0195(.A1(new_n309), .A2(new_n310), .A3(new_n360), .A4(G20), .ZN(new_n396));
  OAI21_X1  g0196(.A(G68), .B1(new_n395), .B2(new_n396), .ZN(new_n397));
  INV_X1    g0197(.A(new_n358), .ZN(new_n398));
  NAND3_X1  g0198(.A1(new_n397), .A2(new_n367), .A3(new_n398), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n399), .A2(KEYINPUT16), .ZN(new_n400));
  NAND3_X1  g0200(.A1(new_n364), .A2(new_n356), .A3(new_n367), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n400), .A2(new_n401), .ZN(new_n402));
  AOI211_X1 g0202(.A(new_n372), .B(new_n375), .C1(new_n402), .C2(new_n288), .ZN(new_n403));
  INV_X1    g0203(.A(KEYINPUT17), .ZN(new_n404));
  XOR2_X1   g0204(.A(KEYINPUT73), .B(G190), .Z(new_n405));
  NAND3_X1  g0205(.A1(new_n385), .A2(new_n405), .A3(new_n386), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n387), .A2(G200), .ZN(new_n407));
  NAND4_X1  g0207(.A1(new_n403), .A2(new_n404), .A3(new_n406), .A4(new_n407), .ZN(new_n408));
  NAND4_X1  g0208(.A1(new_n407), .A2(new_n371), .A3(new_n373), .A4(new_n376), .ZN(new_n409));
  INV_X1    g0209(.A(new_n406), .ZN(new_n410));
  OAI21_X1  g0210(.A(KEYINPUT17), .B1(new_n409), .B2(new_n410), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n408), .A2(new_n411), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n394), .A2(new_n412), .ZN(new_n413));
  AND3_X1   g0213(.A1(new_n350), .A2(new_n268), .A3(new_n351), .ZN(new_n414));
  NOR2_X1   g0214(.A1(new_n414), .A2(G169), .ZN(new_n415));
  OAI21_X1  g0215(.A(new_n343), .B1(new_n352), .B2(new_n304), .ZN(new_n416));
  NOR2_X1   g0216(.A1(new_n415), .A2(new_n416), .ZN(new_n417));
  NOR4_X1   g0217(.A1(new_n306), .A2(new_n355), .A3(new_n413), .A4(new_n417), .ZN(new_n418));
  NAND2_X1  g0218(.A1(G33), .A2(G294), .ZN(new_n419));
  OAI211_X1 g0219(.A(G257), .B(G1698), .C1(new_n309), .C2(new_n310), .ZN(new_n420));
  INV_X1    g0220(.A(G250), .ZN(new_n421));
  OAI211_X1 g0221(.A(new_n419), .B(new_n420), .C1(new_n348), .C2(new_n421), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n422), .A2(KEYINPUT83), .ZN(new_n423));
  NAND3_X1  g0223(.A1(new_n253), .A2(new_n255), .A3(G250), .ZN(new_n424));
  INV_X1    g0224(.A(KEYINPUT83), .ZN(new_n425));
  NAND4_X1  g0225(.A1(new_n424), .A2(new_n425), .A3(new_n419), .A4(new_n420), .ZN(new_n426));
  NAND3_X1  g0226(.A1(new_n423), .A2(new_n263), .A3(new_n426), .ZN(new_n427));
  INV_X1    g0227(.A(G45), .ZN(new_n428));
  NOR2_X1   g0228(.A1(new_n428), .A2(G1), .ZN(new_n429));
  AND2_X1   g0229(.A1(KEYINPUT5), .A2(G41), .ZN(new_n430));
  NOR2_X1   g0230(.A1(KEYINPUT5), .A2(G41), .ZN(new_n431));
  OAI21_X1  g0231(.A(new_n429), .B1(new_n430), .B2(new_n431), .ZN(new_n432));
  OR2_X1    g0232(.A1(new_n432), .A2(new_n266), .ZN(new_n433));
  NAND3_X1  g0233(.A1(new_n432), .A2(G264), .A3(new_n262), .ZN(new_n434));
  NAND3_X1  g0234(.A1(new_n427), .A2(new_n433), .A3(new_n434), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n435), .A2(G169), .ZN(new_n436));
  INV_X1    g0236(.A(KEYINPUT84), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n436), .A2(new_n437), .ZN(new_n438));
  OR2_X1    g0238(.A1(new_n435), .A2(new_n322), .ZN(new_n439));
  NAND3_X1  g0239(.A1(new_n435), .A2(KEYINPUT84), .A3(G169), .ZN(new_n440));
  NAND3_X1  g0240(.A1(new_n438), .A2(new_n439), .A3(new_n440), .ZN(new_n441));
  NAND3_X1  g0241(.A1(new_n218), .A2(G33), .A3(G116), .ZN(new_n442));
  NOR2_X1   g0242(.A1(new_n218), .A2(G107), .ZN(new_n443));
  XNOR2_X1  g0243(.A(new_n443), .B(KEYINPUT23), .ZN(new_n444));
  NAND3_X1  g0244(.A1(new_n253), .A2(new_n218), .A3(G87), .ZN(new_n445));
  AND2_X1   g0245(.A1(new_n445), .A2(KEYINPUT22), .ZN(new_n446));
  NOR2_X1   g0246(.A1(new_n445), .A2(KEYINPUT22), .ZN(new_n447));
  OAI211_X1 g0247(.A(new_n442), .B(new_n444), .C1(new_n446), .C2(new_n447), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n448), .A2(KEYINPUT81), .ZN(new_n449));
  XNOR2_X1  g0249(.A(new_n445), .B(KEYINPUT22), .ZN(new_n450));
  INV_X1    g0250(.A(KEYINPUT81), .ZN(new_n451));
  NAND4_X1  g0251(.A1(new_n450), .A2(new_n451), .A3(new_n442), .A4(new_n444), .ZN(new_n452));
  NAND3_X1  g0252(.A1(new_n449), .A2(new_n452), .A3(KEYINPUT24), .ZN(new_n453));
  INV_X1    g0253(.A(KEYINPUT24), .ZN(new_n454));
  NAND3_X1  g0254(.A1(new_n448), .A2(KEYINPUT81), .A3(new_n454), .ZN(new_n455));
  NAND3_X1  g0255(.A1(new_n453), .A2(new_n288), .A3(new_n455), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n332), .A2(new_n443), .ZN(new_n457));
  XNOR2_X1  g0257(.A(new_n457), .B(KEYINPUT25), .ZN(new_n458));
  OAI211_X1 g0258(.A(new_n287), .B(new_n289), .C1(G1), .C2(new_n260), .ZN(new_n459));
  INV_X1    g0259(.A(new_n459), .ZN(new_n460));
  AOI21_X1  g0260(.A(new_n458), .B1(new_n460), .B2(G107), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n456), .A2(new_n461), .ZN(new_n462));
  INV_X1    g0262(.A(KEYINPUT82), .ZN(new_n463));
  NOR2_X1   g0263(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  AOI21_X1  g0264(.A(KEYINPUT82), .B1(new_n456), .B2(new_n461), .ZN(new_n465));
  OAI21_X1  g0265(.A(new_n441), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  INV_X1    g0266(.A(new_n433), .ZN(new_n467));
  INV_X1    g0267(.A(KEYINPUT4), .ZN(new_n468));
  INV_X1    g0268(.A(G244), .ZN(new_n469));
  OAI21_X1  g0269(.A(new_n468), .B1(new_n348), .B2(new_n469), .ZN(new_n470));
  NAND2_X1  g0270(.A1(G33), .A2(G283), .ZN(new_n471));
  NAND3_X1  g0271(.A1(new_n253), .A2(G250), .A3(G1698), .ZN(new_n472));
  NAND4_X1  g0272(.A1(new_n253), .A2(new_n255), .A3(KEYINPUT4), .A4(G244), .ZN(new_n473));
  NAND4_X1  g0273(.A1(new_n470), .A2(new_n471), .A3(new_n472), .A4(new_n473), .ZN(new_n474));
  AOI21_X1  g0274(.A(new_n467), .B1(new_n474), .B2(new_n263), .ZN(new_n475));
  NAND3_X1  g0275(.A1(new_n432), .A2(G257), .A3(new_n262), .ZN(new_n476));
  INV_X1    g0276(.A(KEYINPUT76), .ZN(new_n477));
  XNOR2_X1  g0277(.A(new_n476), .B(new_n477), .ZN(new_n478));
  NAND3_X1  g0278(.A1(new_n475), .A2(new_n272), .A3(new_n478), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n474), .A2(new_n263), .ZN(new_n480));
  AND3_X1   g0280(.A1(new_n480), .A2(new_n433), .A3(new_n478), .ZN(new_n481));
  OAI21_X1  g0281(.A(new_n479), .B1(new_n481), .B2(G200), .ZN(new_n482));
  INV_X1    g0282(.A(KEYINPUT75), .ZN(new_n483));
  OAI21_X1  g0283(.A(G107), .B1(new_n395), .B2(new_n396), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n484), .A2(KEYINPUT74), .ZN(new_n485));
  INV_X1    g0285(.A(G107), .ZN(new_n486));
  NAND3_X1  g0286(.A1(new_n486), .A2(KEYINPUT6), .A3(G97), .ZN(new_n487));
  NOR2_X1   g0287(.A1(new_n213), .A2(new_n486), .ZN(new_n488));
  NOR2_X1   g0288(.A1(G97), .A2(G107), .ZN(new_n489));
  NOR2_X1   g0289(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  OAI21_X1  g0290(.A(new_n487), .B1(new_n490), .B2(KEYINPUT6), .ZN(new_n491));
  AOI22_X1  g0291(.A1(new_n491), .A2(G20), .B1(G77), .B2(new_n279), .ZN(new_n492));
  INV_X1    g0292(.A(KEYINPUT74), .ZN(new_n493));
  NAND3_X1  g0293(.A1(new_n363), .A2(new_n493), .A3(G107), .ZN(new_n494));
  NAND3_X1  g0294(.A1(new_n485), .A2(new_n492), .A3(new_n494), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n495), .A2(new_n288), .ZN(new_n496));
  NOR2_X1   g0296(.A1(new_n289), .A2(G97), .ZN(new_n497));
  INV_X1    g0297(.A(new_n497), .ZN(new_n498));
  OAI21_X1  g0298(.A(new_n498), .B1(new_n459), .B2(new_n213), .ZN(new_n499));
  INV_X1    g0299(.A(new_n499), .ZN(new_n500));
  AOI21_X1  g0300(.A(new_n483), .B1(new_n496), .B2(new_n500), .ZN(new_n501));
  AOI211_X1 g0301(.A(KEYINPUT75), .B(new_n499), .C1(new_n495), .C2(new_n288), .ZN(new_n502));
  OAI21_X1  g0302(.A(new_n482), .B1(new_n501), .B2(new_n502), .ZN(new_n503));
  AND2_X1   g0303(.A1(new_n340), .A2(new_n290), .ZN(new_n504));
  NAND3_X1  g0304(.A1(new_n282), .A2(G97), .A3(new_n283), .ZN(new_n505));
  INV_X1    g0305(.A(KEYINPUT19), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  NAND3_X1  g0307(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n508), .A2(new_n218), .ZN(new_n509));
  INV_X1    g0309(.A(G87), .ZN(new_n510));
  NAND3_X1  g0310(.A1(new_n510), .A2(new_n213), .A3(new_n486), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n509), .A2(new_n511), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n512), .A2(KEYINPUT77), .ZN(new_n513));
  NAND3_X1  g0313(.A1(new_n253), .A2(new_n218), .A3(G68), .ZN(new_n514));
  INV_X1    g0314(.A(KEYINPUT77), .ZN(new_n515));
  NAND3_X1  g0315(.A1(new_n509), .A2(new_n515), .A3(new_n511), .ZN(new_n516));
  NAND4_X1  g0316(.A1(new_n507), .A2(new_n513), .A3(new_n514), .A4(new_n516), .ZN(new_n517));
  AOI21_X1  g0317(.A(new_n504), .B1(new_n517), .B2(new_n288), .ZN(new_n518));
  NAND2_X1  g0318(.A1(G33), .A2(G116), .ZN(new_n519));
  OAI211_X1 g0319(.A(G244), .B(G1698), .C1(new_n309), .C2(new_n310), .ZN(new_n520));
  OAI211_X1 g0320(.A(new_n519), .B(new_n520), .C1(new_n348), .C2(new_n212), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n521), .A2(new_n263), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n217), .A2(G45), .ZN(new_n523));
  NAND3_X1  g0323(.A1(new_n262), .A2(G250), .A3(new_n523), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n429), .A2(G274), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  INV_X1    g0326(.A(new_n526), .ZN(new_n527));
  NAND3_X1  g0327(.A1(new_n522), .A2(G190), .A3(new_n527), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n460), .A2(G87), .ZN(new_n529));
  AND3_X1   g0329(.A1(new_n518), .A2(new_n528), .A3(new_n529), .ZN(new_n530));
  INV_X1    g0330(.A(G200), .ZN(new_n531));
  AOI21_X1  g0331(.A(new_n526), .B1(new_n521), .B2(new_n263), .ZN(new_n532));
  OAI21_X1  g0332(.A(new_n530), .B1(new_n531), .B2(new_n532), .ZN(new_n533));
  OR2_X1    g0333(.A1(new_n459), .A2(new_n340), .ZN(new_n534));
  AOI22_X1  g0334(.A1(new_n518), .A2(new_n534), .B1(new_n303), .B2(new_n532), .ZN(new_n535));
  OAI21_X1  g0335(.A(new_n535), .B1(G169), .B2(new_n532), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n533), .A2(new_n536), .ZN(new_n537));
  INV_X1    g0337(.A(new_n537), .ZN(new_n538));
  AND3_X1   g0338(.A1(new_n475), .A2(new_n303), .A3(new_n478), .ZN(new_n539));
  AOI21_X1  g0339(.A(G169), .B1(new_n475), .B2(new_n478), .ZN(new_n540));
  NOR2_X1   g0340(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  AOI21_X1  g0341(.A(new_n499), .B1(new_n495), .B2(new_n288), .ZN(new_n542));
  INV_X1    g0342(.A(new_n542), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n541), .A2(new_n543), .ZN(new_n544));
  AND3_X1   g0344(.A1(new_n503), .A2(new_n538), .A3(new_n544), .ZN(new_n545));
  OR2_X1    g0345(.A1(KEYINPUT79), .A2(G303), .ZN(new_n546));
  NAND2_X1  g0346(.A1(KEYINPUT79), .A2(G303), .ZN(new_n547));
  NAND4_X1  g0347(.A1(new_n546), .A2(new_n251), .A3(new_n252), .A4(new_n547), .ZN(new_n548));
  OAI211_X1 g0348(.A(G264), .B(G1698), .C1(new_n309), .C2(new_n310), .ZN(new_n549));
  OAI211_X1 g0349(.A(new_n548), .B(new_n549), .C1(new_n348), .C2(new_n214), .ZN(new_n550));
  INV_X1    g0350(.A(KEYINPUT80), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  NAND3_X1  g0352(.A1(new_n253), .A2(new_n255), .A3(G257), .ZN(new_n553));
  NAND4_X1  g0353(.A1(new_n553), .A2(KEYINPUT80), .A3(new_n548), .A4(new_n549), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n552), .A2(new_n554), .ZN(new_n555));
  AOI21_X1  g0355(.A(new_n467), .B1(new_n555), .B2(new_n263), .ZN(new_n556));
  NAND3_X1  g0356(.A1(new_n432), .A2(G270), .A3(new_n262), .ZN(new_n557));
  XOR2_X1   g0357(.A(new_n557), .B(KEYINPUT78), .Z(new_n558));
  AOI21_X1  g0358(.A(new_n301), .B1(new_n556), .B2(new_n558), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n460), .A2(G116), .ZN(new_n560));
  NOR2_X1   g0360(.A1(new_n218), .A2(G116), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n332), .A2(new_n561), .ZN(new_n562));
  NOR2_X1   g0362(.A1(new_n287), .A2(new_n561), .ZN(new_n563));
  OAI211_X1 g0363(.A(new_n471), .B(new_n218), .C1(G33), .C2(new_n213), .ZN(new_n564));
  AND3_X1   g0364(.A1(new_n563), .A2(KEYINPUT20), .A3(new_n564), .ZN(new_n565));
  AOI21_X1  g0365(.A(KEYINPUT20), .B1(new_n563), .B2(new_n564), .ZN(new_n566));
  OAI211_X1 g0366(.A(new_n560), .B(new_n562), .C1(new_n565), .C2(new_n566), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n559), .A2(new_n567), .ZN(new_n568));
  INV_X1    g0368(.A(KEYINPUT21), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n555), .A2(new_n263), .ZN(new_n571));
  NAND3_X1  g0371(.A1(new_n571), .A2(new_n433), .A3(new_n558), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n572), .A2(G200), .ZN(new_n573));
  INV_X1    g0373(.A(new_n567), .ZN(new_n574));
  INV_X1    g0374(.A(new_n405), .ZN(new_n575));
  OAI211_X1 g0375(.A(new_n573), .B(new_n574), .C1(new_n575), .C2(new_n572), .ZN(new_n576));
  NAND4_X1  g0376(.A1(new_n567), .A2(new_n556), .A3(G179), .A4(new_n558), .ZN(new_n577));
  NAND4_X1  g0377(.A1(new_n572), .A2(KEYINPUT21), .A3(G169), .A4(new_n567), .ZN(new_n578));
  AND4_X1   g0378(.A1(new_n570), .A2(new_n576), .A3(new_n577), .A4(new_n578), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n435), .A2(new_n531), .ZN(new_n580));
  NAND4_X1  g0380(.A1(new_n427), .A2(new_n272), .A3(new_n433), .A4(new_n434), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  NAND3_X1  g0382(.A1(new_n456), .A2(new_n582), .A3(new_n461), .ZN(new_n583));
  NAND4_X1  g0383(.A1(new_n466), .A2(new_n545), .A3(new_n579), .A4(new_n583), .ZN(new_n584));
  INV_X1    g0384(.A(new_n584), .ZN(new_n585));
  AND2_X1   g0385(.A1(new_n418), .A2(new_n585), .ZN(G372));
  AND3_X1   g0386(.A1(new_n392), .A2(KEYINPUT87), .A3(new_n393), .ZN(new_n587));
  AOI21_X1  g0387(.A(KEYINPUT87), .B1(new_n392), .B2(new_n393), .ZN(new_n588));
  OR2_X1    g0388(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  AOI22_X1  g0389(.A1(new_n325), .A2(new_n335), .B1(new_n417), .B2(new_n338), .ZN(new_n590));
  INV_X1    g0390(.A(new_n412), .ZN(new_n591));
  OAI21_X1  g0391(.A(new_n589), .B1(new_n590), .B2(new_n591), .ZN(new_n592));
  NAND3_X1  g0392(.A1(new_n592), .A2(new_n298), .A3(new_n300), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n593), .A2(new_n305), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n594), .A2(KEYINPUT88), .ZN(new_n595));
  INV_X1    g0395(.A(KEYINPUT88), .ZN(new_n596));
  NAND3_X1  g0396(.A1(new_n593), .A2(new_n596), .A3(new_n305), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n595), .A2(new_n597), .ZN(new_n598));
  INV_X1    g0398(.A(KEYINPUT85), .ZN(new_n599));
  XNOR2_X1  g0399(.A(new_n526), .B(new_n599), .ZN(new_n600));
  INV_X1    g0400(.A(new_n522), .ZN(new_n601));
  OAI21_X1  g0401(.A(new_n301), .B1(new_n600), .B2(new_n601), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n535), .A2(new_n602), .ZN(new_n603));
  INV_X1    g0403(.A(new_n603), .ZN(new_n604));
  OAI21_X1  g0404(.A(G200), .B1(new_n600), .B2(new_n601), .ZN(new_n605));
  AOI22_X1  g0405(.A1(new_n530), .A2(new_n605), .B1(new_n535), .B2(new_n602), .ZN(new_n606));
  AND4_X1   g0406(.A1(new_n583), .A2(new_n503), .A3(new_n544), .A4(new_n606), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n578), .A2(new_n577), .ZN(new_n608));
  AOI21_X1  g0408(.A(KEYINPUT21), .B1(new_n559), .B2(new_n567), .ZN(new_n609));
  NOR2_X1   g0409(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n441), .A2(new_n462), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  AOI21_X1  g0412(.A(new_n604), .B1(new_n607), .B2(new_n612), .ZN(new_n613));
  NOR3_X1   g0413(.A1(new_n539), .A2(new_n542), .A3(new_n540), .ZN(new_n614));
  NAND4_X1  g0414(.A1(new_n538), .A2(KEYINPUT86), .A3(KEYINPUT26), .A4(new_n614), .ZN(new_n615));
  INV_X1    g0415(.A(KEYINPUT86), .ZN(new_n616));
  AOI21_X1  g0416(.A(new_n493), .B1(new_n363), .B2(G107), .ZN(new_n617));
  AOI211_X1 g0417(.A(KEYINPUT74), .B(new_n486), .C1(new_n361), .C2(new_n362), .ZN(new_n618));
  NOR2_X1   g0418(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  AOI21_X1  g0419(.A(new_n287), .B1(new_n619), .B2(new_n492), .ZN(new_n620));
  OAI21_X1  g0420(.A(KEYINPUT75), .B1(new_n620), .B2(new_n499), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n542), .A2(new_n483), .ZN(new_n622));
  NAND4_X1  g0422(.A1(new_n606), .A2(new_n541), .A3(new_n621), .A4(new_n622), .ZN(new_n623));
  INV_X1    g0423(.A(KEYINPUT26), .ZN(new_n624));
  AOI21_X1  g0424(.A(new_n616), .B1(new_n623), .B2(new_n624), .ZN(new_n625));
  NOR3_X1   g0425(.A1(new_n544), .A2(new_n537), .A3(new_n624), .ZN(new_n626));
  OAI21_X1  g0426(.A(new_n615), .B1(new_n625), .B2(new_n626), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n613), .A2(new_n627), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n418), .A2(new_n628), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n598), .A2(new_n629), .ZN(G369));
  XOR2_X1   g0430(.A(new_n579), .B(KEYINPUT90), .Z(new_n631));
  NAND2_X1  g0431(.A1(new_n332), .A2(new_n218), .ZN(new_n632));
  NOR2_X1   g0432(.A1(new_n632), .A2(KEYINPUT27), .ZN(new_n633));
  XNOR2_X1  g0433(.A(new_n633), .B(KEYINPUT89), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n632), .A2(KEYINPUT27), .ZN(new_n635));
  NAND3_X1  g0435(.A1(new_n634), .A2(G213), .A3(new_n635), .ZN(new_n636));
  INV_X1    g0436(.A(G343), .ZN(new_n637));
  NOR2_X1   g0437(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n638), .A2(new_n567), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n631), .A2(new_n639), .ZN(new_n640));
  INV_X1    g0440(.A(new_n610), .ZN(new_n641));
  OAI21_X1  g0441(.A(new_n640), .B1(new_n641), .B2(new_n639), .ZN(new_n642));
  INV_X1    g0442(.A(G330), .ZN(new_n643));
  OR2_X1    g0443(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  INV_X1    g0444(.A(new_n466), .ZN(new_n645));
  NAND3_X1  g0445(.A1(new_n645), .A2(KEYINPUT91), .A3(new_n638), .ZN(new_n646));
  INV_X1    g0446(.A(KEYINPUT91), .ZN(new_n647));
  INV_X1    g0447(.A(new_n638), .ZN(new_n648));
  OAI21_X1  g0448(.A(new_n647), .B1(new_n466), .B2(new_n648), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n646), .A2(new_n649), .ZN(new_n650));
  AND2_X1   g0450(.A1(new_n466), .A2(new_n583), .ZN(new_n651));
  OAI21_X1  g0451(.A(new_n638), .B1(new_n464), .B2(new_n465), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  AND2_X1   g0453(.A1(new_n650), .A2(new_n653), .ZN(new_n654));
  NOR2_X1   g0454(.A1(new_n644), .A2(new_n654), .ZN(new_n655));
  NOR2_X1   g0455(.A1(new_n611), .A2(new_n638), .ZN(new_n656));
  INV_X1    g0456(.A(new_n656), .ZN(new_n657));
  NOR2_X1   g0457(.A1(new_n610), .A2(new_n638), .ZN(new_n658));
  INV_X1    g0458(.A(new_n658), .ZN(new_n659));
  OAI21_X1  g0459(.A(new_n657), .B1(new_n654), .B2(new_n659), .ZN(new_n660));
  OR2_X1    g0460(.A1(new_n655), .A2(new_n660), .ZN(G399));
  NAND3_X1  g0461(.A1(new_n229), .A2(KEYINPUT92), .A3(new_n261), .ZN(new_n662));
  INV_X1    g0462(.A(KEYINPUT92), .ZN(new_n663));
  OAI21_X1  g0463(.A(new_n663), .B1(new_n228), .B2(G41), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n662), .A2(new_n664), .ZN(new_n665));
  INV_X1    g0465(.A(new_n665), .ZN(new_n666));
  NOR2_X1   g0466(.A1(new_n511), .A2(G116), .ZN(new_n667));
  INV_X1    g0467(.A(new_n667), .ZN(new_n668));
  NOR3_X1   g0468(.A1(new_n666), .A2(new_n217), .A3(new_n668), .ZN(new_n669));
  INV_X1    g0469(.A(new_n223), .ZN(new_n670));
  AOI21_X1  g0470(.A(new_n669), .B1(new_n670), .B2(new_n666), .ZN(new_n671));
  XOR2_X1   g0471(.A(new_n671), .B(KEYINPUT28), .Z(new_n672));
  NAND3_X1  g0472(.A1(new_n556), .A2(G179), .A3(new_n558), .ZN(new_n673));
  OR2_X1    g0473(.A1(new_n673), .A2(KEYINPUT93), .ZN(new_n674));
  AND3_X1   g0474(.A1(new_n481), .A2(new_n434), .A3(new_n427), .ZN(new_n675));
  INV_X1    g0475(.A(new_n532), .ZN(new_n676));
  AOI21_X1  g0476(.A(new_n676), .B1(new_n673), .B2(KEYINPUT93), .ZN(new_n677));
  NAND3_X1  g0477(.A1(new_n674), .A2(new_n675), .A3(new_n677), .ZN(new_n678));
  INV_X1    g0478(.A(KEYINPUT30), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  NAND4_X1  g0480(.A1(new_n674), .A2(new_n677), .A3(KEYINPUT30), .A4(new_n675), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  NOR2_X1   g0482(.A1(new_n600), .A2(new_n601), .ZN(new_n683));
  NOR3_X1   g0483(.A1(new_n481), .A2(new_n304), .A3(new_n683), .ZN(new_n684));
  NAND3_X1  g0484(.A1(new_n684), .A2(new_n435), .A3(new_n572), .ZN(new_n685));
  INV_X1    g0485(.A(new_n685), .ZN(new_n686));
  OAI21_X1  g0486(.A(new_n638), .B1(new_n682), .B2(new_n686), .ZN(new_n687));
  OAI211_X1 g0487(.A(new_n687), .B(KEYINPUT31), .C1(new_n584), .C2(new_n638), .ZN(new_n688));
  INV_X1    g0488(.A(KEYINPUT31), .ZN(new_n689));
  OAI211_X1 g0489(.A(new_n689), .B(new_n638), .C1(new_n682), .C2(new_n686), .ZN(new_n690));
  AND2_X1   g0490(.A1(new_n688), .A2(new_n690), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n691), .A2(G330), .ZN(new_n692));
  AOI21_X1  g0492(.A(new_n638), .B1(new_n613), .B2(new_n627), .ZN(new_n693));
  OR2_X1    g0493(.A1(new_n693), .A2(KEYINPUT29), .ZN(new_n694));
  OAI21_X1  g0494(.A(new_n607), .B1(new_n645), .B2(new_n641), .ZN(new_n695));
  NAND3_X1  g0495(.A1(new_n538), .A2(new_n624), .A3(new_n614), .ZN(new_n696));
  AOI21_X1  g0496(.A(new_n604), .B1(new_n623), .B2(KEYINPUT26), .ZN(new_n697));
  NAND3_X1  g0497(.A1(new_n695), .A2(new_n696), .A3(new_n697), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n698), .A2(new_n648), .ZN(new_n699));
  INV_X1    g0499(.A(KEYINPUT29), .ZN(new_n700));
  OAI21_X1  g0500(.A(new_n694), .B1(new_n699), .B2(new_n700), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n692), .A2(new_n701), .ZN(new_n702));
  INV_X1    g0502(.A(new_n702), .ZN(new_n703));
  OAI21_X1  g0503(.A(new_n672), .B1(new_n703), .B2(G1), .ZN(G364));
  NOR2_X1   g0504(.A1(new_n224), .A2(G20), .ZN(new_n705));
  AOI21_X1  g0505(.A(new_n217), .B1(new_n705), .B2(G45), .ZN(new_n706));
  INV_X1    g0506(.A(new_n706), .ZN(new_n707));
  NOR2_X1   g0507(.A1(new_n666), .A2(new_n707), .ZN(new_n708));
  INV_X1    g0508(.A(new_n708), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n642), .A2(new_n643), .ZN(new_n710));
  NAND3_X1  g0510(.A1(new_n644), .A2(new_n709), .A3(new_n710), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n245), .A2(G45), .ZN(new_n712));
  NOR2_X1   g0512(.A1(new_n228), .A2(new_n253), .ZN(new_n713));
  OAI211_X1 g0513(.A(new_n712), .B(new_n713), .C1(G45), .C2(new_n223), .ZN(new_n714));
  NAND3_X1  g0514(.A1(new_n229), .A2(G355), .A3(new_n253), .ZN(new_n715));
  OAI211_X1 g0515(.A(new_n714), .B(new_n715), .C1(G116), .C2(new_n229), .ZN(new_n716));
  OAI21_X1  g0516(.A(new_n225), .B1(new_n218), .B2(G169), .ZN(new_n717));
  OR2_X1    g0517(.A1(new_n717), .A2(KEYINPUT95), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n717), .A2(KEYINPUT95), .ZN(new_n719));
  NAND2_X1  g0519(.A1(new_n718), .A2(new_n719), .ZN(new_n720));
  NOR2_X1   g0520(.A1(G13), .A2(G33), .ZN(new_n721));
  XOR2_X1   g0521(.A(new_n721), .B(KEYINPUT94), .Z(new_n722));
  NOR2_X1   g0522(.A1(new_n722), .A2(G20), .ZN(new_n723));
  NOR2_X1   g0523(.A1(new_n720), .A2(new_n723), .ZN(new_n724));
  NAND2_X1  g0524(.A1(new_n716), .A2(new_n724), .ZN(new_n725));
  NOR2_X1   g0525(.A1(new_n218), .A2(G190), .ZN(new_n726));
  NOR2_X1   g0526(.A1(new_n531), .A2(G179), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  XOR2_X1   g0528(.A(new_n728), .B(KEYINPUT99), .Z(new_n729));
  INV_X1    g0529(.A(G283), .ZN(new_n730));
  NOR2_X1   g0530(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  INV_X1    g0531(.A(G294), .ZN(new_n732));
  NOR2_X1   g0532(.A1(G179), .A2(G200), .ZN(new_n733));
  AOI21_X1  g0533(.A(new_n218), .B1(new_n733), .B2(G190), .ZN(new_n734));
  NAND3_X1  g0534(.A1(new_n727), .A2(G20), .A3(G190), .ZN(new_n735));
  INV_X1    g0535(.A(KEYINPUT98), .ZN(new_n736));
  OR2_X1    g0536(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  NAND2_X1  g0537(.A1(new_n735), .A2(new_n736), .ZN(new_n738));
  NAND2_X1  g0538(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  INV_X1    g0539(.A(G303), .ZN(new_n740));
  OAI221_X1 g0540(.A(new_n311), .B1(new_n732), .B2(new_n734), .C1(new_n739), .C2(new_n740), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n726), .A2(new_n733), .ZN(new_n742));
  INV_X1    g0542(.A(new_n742), .ZN(new_n743));
  AOI211_X1 g0543(.A(new_n731), .B(new_n741), .C1(G329), .C2(new_n743), .ZN(new_n744));
  NOR2_X1   g0544(.A1(new_n303), .A2(new_n218), .ZN(new_n745));
  NAND2_X1  g0545(.A1(new_n745), .A2(G200), .ZN(new_n746));
  NOR2_X1   g0546(.A1(new_n746), .A2(new_n575), .ZN(new_n747));
  NOR2_X1   g0547(.A1(new_n746), .A2(G190), .ZN(new_n748));
  XNOR2_X1  g0548(.A(KEYINPUT33), .B(G317), .ZN(new_n749));
  AOI22_X1  g0549(.A1(G326), .A2(new_n747), .B1(new_n748), .B2(new_n749), .ZN(new_n750));
  INV_X1    g0550(.A(G322), .ZN(new_n751));
  NAND2_X1  g0551(.A1(new_n745), .A2(new_n531), .ZN(new_n752));
  NOR2_X1   g0552(.A1(new_n752), .A2(new_n575), .ZN(new_n753));
  AND2_X1   g0553(.A1(new_n753), .A2(KEYINPUT96), .ZN(new_n754));
  NOR2_X1   g0554(.A1(new_n753), .A2(KEYINPUT96), .ZN(new_n755));
  NOR2_X1   g0555(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  OAI211_X1 g0556(.A(new_n744), .B(new_n750), .C1(new_n751), .C2(new_n756), .ZN(new_n757));
  NOR2_X1   g0557(.A1(new_n752), .A2(G190), .ZN(new_n758));
  AOI21_X1  g0558(.A(new_n757), .B1(G311), .B2(new_n758), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n729), .A2(new_n486), .ZN(new_n760));
  NOR2_X1   g0560(.A1(new_n742), .A2(new_n365), .ZN(new_n761));
  INV_X1    g0561(.A(KEYINPUT32), .ZN(new_n762));
  OAI22_X1  g0562(.A1(new_n761), .A2(new_n762), .B1(new_n213), .B2(new_n734), .ZN(new_n763));
  INV_X1    g0563(.A(G58), .ZN(new_n764));
  INV_X1    g0564(.A(new_n758), .ZN(new_n765));
  OAI22_X1  g0565(.A1(new_n756), .A2(new_n764), .B1(new_n258), .B2(new_n765), .ZN(new_n766));
  INV_X1    g0566(.A(new_n747), .ZN(new_n767));
  NOR2_X1   g0567(.A1(new_n767), .A2(new_n202), .ZN(new_n768));
  NOR2_X1   g0568(.A1(new_n766), .A2(new_n768), .ZN(new_n769));
  INV_X1    g0569(.A(new_n769), .ZN(new_n770));
  AOI211_X1 g0570(.A(new_n760), .B(new_n763), .C1(new_n770), .C2(KEYINPUT97), .ZN(new_n771));
  AOI21_X1  g0571(.A(new_n311), .B1(new_n761), .B2(new_n762), .ZN(new_n772));
  INV_X1    g0572(.A(new_n748), .ZN(new_n773));
  OAI221_X1 g0573(.A(new_n772), .B1(new_n510), .B2(new_n739), .C1(new_n773), .C2(new_n211), .ZN(new_n774));
  INV_X1    g0574(.A(KEYINPUT97), .ZN(new_n775));
  AOI21_X1  g0575(.A(new_n774), .B1(new_n769), .B2(new_n775), .ZN(new_n776));
  AOI21_X1  g0576(.A(new_n759), .B1(new_n771), .B2(new_n776), .ZN(new_n777));
  INV_X1    g0577(.A(new_n720), .ZN(new_n778));
  OAI21_X1  g0578(.A(new_n725), .B1(new_n777), .B2(new_n778), .ZN(new_n779));
  AOI21_X1  g0579(.A(new_n779), .B1(new_n642), .B2(new_n723), .ZN(new_n780));
  NAND2_X1  g0580(.A1(new_n780), .A2(new_n708), .ZN(new_n781));
  AND2_X1   g0581(.A1(new_n711), .A2(new_n781), .ZN(new_n782));
  INV_X1    g0582(.A(new_n782), .ZN(G396));
  INV_X1    g0583(.A(G137), .ZN(new_n784));
  OAI22_X1  g0584(.A1(new_n784), .A2(new_n767), .B1(new_n773), .B2(new_n278), .ZN(new_n785));
  INV_X1    g0585(.A(new_n756), .ZN(new_n786));
  AOI21_X1  g0586(.A(new_n785), .B1(new_n786), .B2(G143), .ZN(new_n787));
  OAI21_X1  g0587(.A(new_n787), .B1(new_n365), .B2(new_n765), .ZN(new_n788));
  XNOR2_X1  g0588(.A(new_n788), .B(KEYINPUT34), .ZN(new_n789));
  INV_X1    g0589(.A(new_n739), .ZN(new_n790));
  NAND2_X1  g0590(.A1(new_n790), .A2(G50), .ZN(new_n791));
  AOI21_X1  g0591(.A(new_n311), .B1(new_n743), .B2(G132), .ZN(new_n792));
  NOR2_X1   g0592(.A1(new_n729), .A2(new_n211), .ZN(new_n793));
  INV_X1    g0593(.A(new_n734), .ZN(new_n794));
  AOI21_X1  g0594(.A(new_n793), .B1(G58), .B2(new_n794), .ZN(new_n795));
  NAND4_X1  g0595(.A1(new_n789), .A2(new_n791), .A3(new_n792), .A4(new_n795), .ZN(new_n796));
  AOI22_X1  g0596(.A1(new_n786), .A2(G294), .B1(G97), .B2(new_n794), .ZN(new_n797));
  AOI22_X1  g0597(.A1(G116), .A2(new_n758), .B1(new_n747), .B2(G303), .ZN(new_n798));
  OAI21_X1  g0598(.A(new_n798), .B1(new_n730), .B2(new_n773), .ZN(new_n799));
  OR2_X1    g0599(.A1(new_n799), .A2(KEYINPUT100), .ZN(new_n800));
  NAND2_X1  g0600(.A1(new_n799), .A2(KEYINPUT100), .ZN(new_n801));
  INV_X1    g0601(.A(G311), .ZN(new_n802));
  OAI21_X1  g0602(.A(new_n311), .B1(new_n742), .B2(new_n802), .ZN(new_n803));
  NOR2_X1   g0603(.A1(new_n729), .A2(new_n510), .ZN(new_n804));
  AOI211_X1 g0604(.A(new_n803), .B(new_n804), .C1(G107), .C2(new_n790), .ZN(new_n805));
  NAND4_X1  g0605(.A1(new_n797), .A2(new_n800), .A3(new_n801), .A4(new_n805), .ZN(new_n806));
  AOI21_X1  g0606(.A(new_n778), .B1(new_n796), .B2(new_n806), .ZN(new_n807));
  NAND2_X1  g0607(.A1(new_n638), .A2(new_n343), .ZN(new_n808));
  NAND2_X1  g0608(.A1(new_n354), .A2(new_n808), .ZN(new_n809));
  OAI21_X1  g0609(.A(new_n809), .B1(new_n415), .B2(new_n416), .ZN(new_n810));
  NAND2_X1  g0610(.A1(new_n417), .A2(new_n648), .ZN(new_n811));
  AND2_X1   g0611(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  NOR2_X1   g0612(.A1(new_n812), .A2(new_n722), .ZN(new_n813));
  INV_X1    g0613(.A(new_n722), .ZN(new_n814));
  NOR2_X1   g0614(.A1(new_n720), .A2(new_n814), .ZN(new_n815));
  INV_X1    g0615(.A(new_n815), .ZN(new_n816));
  NOR2_X1   g0616(.A1(new_n816), .A2(G77), .ZN(new_n817));
  NOR4_X1   g0617(.A1(new_n807), .A2(new_n709), .A3(new_n813), .A4(new_n817), .ZN(new_n818));
  INV_X1    g0618(.A(new_n818), .ZN(new_n819));
  NAND3_X1  g0619(.A1(new_n628), .A2(new_n648), .A3(new_n812), .ZN(new_n820));
  INV_X1    g0620(.A(KEYINPUT101), .ZN(new_n821));
  NAND2_X1  g0621(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  NAND3_X1  g0622(.A1(new_n693), .A2(KEYINPUT101), .A3(new_n812), .ZN(new_n823));
  NAND2_X1  g0623(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  OAI21_X1  g0624(.A(new_n824), .B1(new_n693), .B2(new_n812), .ZN(new_n825));
  XNOR2_X1  g0625(.A(new_n825), .B(new_n692), .ZN(new_n826));
  OAI21_X1  g0626(.A(new_n819), .B1(new_n826), .B2(new_n708), .ZN(G384));
  OAI211_X1 g0627(.A(G20), .B(new_n225), .C1(new_n491), .C2(KEYINPUT35), .ZN(new_n828));
  AOI211_X1 g0628(.A(new_n207), .B(new_n828), .C1(KEYINPUT35), .C2(new_n491), .ZN(new_n829));
  XOR2_X1   g0629(.A(new_n829), .B(KEYINPUT36), .Z(new_n830));
  NAND2_X1  g0630(.A1(new_n357), .A2(G77), .ZN(new_n831));
  OAI22_X1  g0631(.A1(new_n223), .A2(new_n831), .B1(G50), .B2(new_n211), .ZN(new_n832));
  NAND3_X1  g0632(.A1(new_n832), .A2(G1), .A3(new_n224), .ZN(new_n833));
  INV_X1    g0633(.A(KEYINPUT40), .ZN(new_n834));
  INV_X1    g0634(.A(new_n636), .ZN(new_n835));
  NAND2_X1  g0635(.A1(new_n377), .A2(new_n835), .ZN(new_n836));
  AOI21_X1  g0636(.A(new_n836), .B1(new_n394), .B2(new_n412), .ZN(new_n837));
  AOI21_X1  g0637(.A(new_n372), .B1(new_n402), .B2(new_n288), .ZN(new_n838));
  NAND4_X1  g0638(.A1(new_n838), .A2(new_n406), .A3(new_n407), .A4(new_n376), .ZN(new_n839));
  NAND4_X1  g0639(.A1(new_n390), .A2(new_n839), .A3(KEYINPUT37), .A4(new_n836), .ZN(new_n840));
  INV_X1    g0640(.A(new_n840), .ZN(new_n841));
  NOR2_X1   g0641(.A1(new_n837), .A2(new_n841), .ZN(new_n842));
  INV_X1    g0642(.A(KEYINPUT103), .ZN(new_n843));
  XNOR2_X1  g0643(.A(new_n636), .B(new_n843), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n377), .A2(new_n844), .ZN(new_n845));
  NAND3_X1  g0645(.A1(new_n390), .A2(new_n839), .A3(new_n845), .ZN(new_n846));
  INV_X1    g0646(.A(new_n846), .ZN(new_n847));
  OR2_X1    g0647(.A1(new_n847), .A2(KEYINPUT37), .ZN(new_n848));
  AOI21_X1  g0648(.A(KEYINPUT38), .B1(new_n842), .B2(new_n848), .ZN(new_n849));
  NOR2_X1   g0649(.A1(new_n847), .A2(KEYINPUT37), .ZN(new_n850));
  INV_X1    g0650(.A(KEYINPUT38), .ZN(new_n851));
  NOR4_X1   g0651(.A1(new_n837), .A2(new_n850), .A3(new_n851), .A4(new_n841), .ZN(new_n852));
  OAI21_X1  g0652(.A(KEYINPUT104), .B1(new_n849), .B2(new_n852), .ZN(new_n853));
  INV_X1    g0653(.A(new_n836), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n413), .A2(new_n854), .ZN(new_n855));
  NAND3_X1  g0655(.A1(new_n855), .A2(new_n848), .A3(new_n840), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n856), .A2(new_n851), .ZN(new_n857));
  INV_X1    g0657(.A(KEYINPUT104), .ZN(new_n858));
  NAND3_X1  g0658(.A1(new_n842), .A2(KEYINPUT38), .A3(new_n848), .ZN(new_n859));
  NAND3_X1  g0659(.A1(new_n857), .A2(new_n858), .A3(new_n859), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n853), .A2(new_n860), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n335), .A2(new_n638), .ZN(new_n862));
  NAND4_X1  g0662(.A1(new_n336), .A2(KEYINPUT102), .A3(new_n338), .A4(new_n862), .ZN(new_n863));
  INV_X1    g0663(.A(new_n335), .ZN(new_n864));
  OAI211_X1 g0664(.A(KEYINPUT102), .B(new_n338), .C1(new_n324), .C2(new_n864), .ZN(new_n865));
  NAND3_X1  g0665(.A1(new_n865), .A2(new_n335), .A3(new_n638), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n863), .A2(new_n866), .ZN(new_n867));
  NAND4_X1  g0667(.A1(new_n688), .A2(new_n690), .A3(new_n867), .A4(new_n812), .ZN(new_n868));
  OAI21_X1  g0668(.A(new_n834), .B1(new_n861), .B2(new_n868), .ZN(new_n869));
  INV_X1    g0669(.A(new_n868), .ZN(new_n870));
  NAND3_X1  g0670(.A1(new_n839), .A2(new_n845), .A3(KEYINPUT87), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n871), .A2(KEYINPUT37), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n872), .A2(new_n846), .ZN(new_n873));
  AND2_X1   g0673(.A1(new_n839), .A2(new_n845), .ZN(new_n874));
  NAND4_X1  g0674(.A1(new_n874), .A2(KEYINPUT37), .A3(new_n871), .A4(new_n390), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n873), .A2(new_n875), .ZN(new_n876));
  OAI21_X1  g0676(.A(new_n412), .B1(new_n587), .B2(new_n588), .ZN(new_n877));
  INV_X1    g0677(.A(new_n845), .ZN(new_n878));
  AOI21_X1  g0678(.A(new_n876), .B1(new_n877), .B2(new_n878), .ZN(new_n879));
  OAI21_X1  g0679(.A(new_n859), .B1(new_n879), .B2(KEYINPUT38), .ZN(new_n880));
  NAND3_X1  g0680(.A1(new_n870), .A2(KEYINPUT40), .A3(new_n880), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n869), .A2(new_n881), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n691), .A2(new_n418), .ZN(new_n883));
  XOR2_X1   g0683(.A(new_n882), .B(new_n883), .Z(new_n884));
  NAND2_X1  g0684(.A1(new_n884), .A2(G330), .ZN(new_n885));
  OAI21_X1  g0685(.A(KEYINPUT39), .B1(new_n849), .B2(new_n852), .ZN(new_n886));
  INV_X1    g0686(.A(KEYINPUT39), .ZN(new_n887));
  OAI211_X1 g0687(.A(new_n887), .B(new_n859), .C1(new_n879), .C2(KEYINPUT38), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n886), .A2(new_n888), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n889), .A2(KEYINPUT105), .ZN(new_n890));
  NOR2_X1   g0690(.A1(new_n336), .A2(new_n638), .ZN(new_n891));
  INV_X1    g0691(.A(KEYINPUT105), .ZN(new_n892));
  NAND3_X1  g0692(.A1(new_n886), .A2(new_n888), .A3(new_n892), .ZN(new_n893));
  NAND3_X1  g0693(.A1(new_n890), .A2(new_n891), .A3(new_n893), .ZN(new_n894));
  OR2_X1    g0694(.A1(new_n589), .A2(new_n844), .ZN(new_n895));
  INV_X1    g0695(.A(new_n811), .ZN(new_n896));
  AOI21_X1  g0696(.A(new_n896), .B1(new_n822), .B2(new_n823), .ZN(new_n897));
  INV_X1    g0697(.A(new_n897), .ZN(new_n898));
  NAND4_X1  g0698(.A1(new_n898), .A2(new_n853), .A3(new_n860), .A4(new_n867), .ZN(new_n899));
  NAND3_X1  g0699(.A1(new_n894), .A2(new_n895), .A3(new_n899), .ZN(new_n900));
  OAI211_X1 g0700(.A(new_n418), .B(new_n694), .C1(new_n699), .C2(new_n700), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n598), .A2(new_n901), .ZN(new_n902));
  XNOR2_X1  g0702(.A(new_n900), .B(new_n902), .ZN(new_n903));
  OAI22_X1  g0703(.A1(new_n885), .A2(new_n903), .B1(new_n217), .B2(new_n705), .ZN(new_n904));
  XOR2_X1   g0704(.A(new_n904), .B(KEYINPUT106), .Z(new_n905));
  AND2_X1   g0705(.A1(new_n885), .A2(new_n903), .ZN(new_n906));
  OAI211_X1 g0706(.A(new_n830), .B(new_n833), .C1(new_n905), .C2(new_n906), .ZN(G367));
  NOR2_X1   g0707(.A1(new_n501), .A2(new_n502), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n908), .A2(new_n638), .ZN(new_n909));
  NAND3_X1  g0709(.A1(new_n909), .A2(new_n544), .A3(new_n503), .ZN(new_n910));
  NAND3_X1  g0710(.A1(new_n908), .A2(new_n541), .A3(new_n638), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n655), .A2(new_n912), .ZN(new_n913));
  INV_X1    g0713(.A(new_n654), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n914), .A2(new_n658), .ZN(new_n915));
  INV_X1    g0715(.A(new_n912), .ZN(new_n916));
  OAI21_X1  g0716(.A(KEYINPUT42), .B1(new_n915), .B2(new_n916), .ZN(new_n917));
  OAI21_X1  g0717(.A(new_n544), .B1(new_n916), .B2(new_n466), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n918), .A2(new_n648), .ZN(new_n919));
  NOR2_X1   g0719(.A1(new_n654), .A2(new_n659), .ZN(new_n920));
  INV_X1    g0720(.A(KEYINPUT42), .ZN(new_n921));
  NAND3_X1  g0721(.A1(new_n920), .A2(new_n921), .A3(new_n912), .ZN(new_n922));
  NAND3_X1  g0722(.A1(new_n917), .A2(new_n919), .A3(new_n922), .ZN(new_n923));
  AOI21_X1  g0723(.A(new_n648), .B1(new_n518), .B2(new_n529), .ZN(new_n924));
  MUX2_X1   g0724(.A(new_n606), .B(new_n604), .S(new_n924), .Z(new_n925));
  NAND2_X1  g0725(.A1(new_n925), .A2(KEYINPUT43), .ZN(new_n926));
  AND3_X1   g0726(.A1(new_n913), .A2(new_n923), .A3(new_n926), .ZN(new_n927));
  AOI21_X1  g0727(.A(new_n913), .B1(new_n923), .B2(new_n926), .ZN(new_n928));
  NOR2_X1   g0728(.A1(new_n925), .A2(KEYINPUT43), .ZN(new_n929));
  INV_X1    g0729(.A(new_n929), .ZN(new_n930));
  OR3_X1    g0730(.A1(new_n927), .A2(new_n928), .A3(new_n930), .ZN(new_n931));
  OAI21_X1  g0731(.A(new_n930), .B1(new_n927), .B2(new_n928), .ZN(new_n932));
  XOR2_X1   g0732(.A(new_n665), .B(KEYINPUT41), .Z(new_n933));
  INV_X1    g0733(.A(new_n933), .ZN(new_n934));
  OAI211_X1 g0734(.A(new_n657), .B(new_n912), .C1(new_n654), .C2(new_n659), .ZN(new_n935));
  XOR2_X1   g0735(.A(new_n935), .B(KEYINPUT45), .Z(new_n936));
  INV_X1    g0736(.A(KEYINPUT44), .ZN(new_n937));
  INV_X1    g0737(.A(new_n660), .ZN(new_n938));
  OAI21_X1  g0738(.A(new_n937), .B1(new_n938), .B2(new_n912), .ZN(new_n939));
  NAND3_X1  g0739(.A1(new_n660), .A2(KEYINPUT44), .A3(new_n916), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n939), .A2(new_n940), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n936), .A2(new_n941), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n942), .A2(new_n655), .ZN(new_n943));
  INV_X1    g0743(.A(new_n644), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n944), .A2(new_n914), .ZN(new_n945));
  NAND3_X1  g0745(.A1(new_n936), .A2(new_n941), .A3(new_n945), .ZN(new_n946));
  INV_X1    g0746(.A(KEYINPUT107), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n644), .A2(new_n947), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n654), .A2(new_n659), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n915), .A2(new_n949), .ZN(new_n950));
  OR2_X1    g0750(.A1(new_n948), .A2(new_n950), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n948), .A2(new_n950), .ZN(new_n952));
  AOI21_X1  g0752(.A(new_n702), .B1(new_n951), .B2(new_n952), .ZN(new_n953));
  NAND3_X1  g0753(.A1(new_n943), .A2(new_n946), .A3(new_n953), .ZN(new_n954));
  AOI21_X1  g0754(.A(new_n934), .B1(new_n954), .B2(new_n703), .ZN(new_n955));
  OAI211_X1 g0755(.A(new_n931), .B(new_n932), .C1(new_n955), .C2(new_n707), .ZN(new_n956));
  OAI22_X1  g0756(.A1(new_n756), .A2(new_n278), .B1(new_n211), .B2(new_n734), .ZN(new_n957));
  XNOR2_X1  g0757(.A(new_n957), .B(KEYINPUT108), .ZN(new_n958));
  OAI221_X1 g0758(.A(new_n253), .B1(new_n258), .B2(new_n728), .C1(new_n739), .C2(new_n764), .ZN(new_n959));
  OAI22_X1  g0759(.A1(new_n202), .A2(new_n765), .B1(new_n773), .B2(new_n365), .ZN(new_n960));
  AOI211_X1 g0760(.A(new_n959), .B(new_n960), .C1(G143), .C2(new_n747), .ZN(new_n961));
  OAI211_X1 g0761(.A(new_n958), .B(new_n961), .C1(new_n784), .C2(new_n742), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n546), .A2(new_n547), .ZN(new_n963));
  INV_X1    g0763(.A(new_n963), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n786), .A2(new_n964), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n790), .A2(G116), .ZN(new_n966));
  INV_X1    g0766(.A(KEYINPUT46), .ZN(new_n967));
  OAI22_X1  g0767(.A1(new_n966), .A2(new_n967), .B1(new_n767), .B2(new_n802), .ZN(new_n968));
  AOI21_X1  g0768(.A(new_n968), .B1(G283), .B2(new_n758), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n966), .A2(new_n967), .ZN(new_n970));
  INV_X1    g0770(.A(G317), .ZN(new_n971));
  NOR2_X1   g0771(.A1(new_n742), .A2(new_n971), .ZN(new_n972));
  OAI221_X1 g0772(.A(new_n311), .B1(new_n734), .B2(new_n486), .C1(new_n728), .C2(new_n213), .ZN(new_n973));
  AOI211_X1 g0773(.A(new_n972), .B(new_n973), .C1(new_n748), .C2(G294), .ZN(new_n974));
  NAND4_X1  g0774(.A1(new_n965), .A2(new_n969), .A3(new_n970), .A4(new_n974), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n962), .A2(new_n975), .ZN(new_n976));
  XOR2_X1   g0776(.A(new_n976), .B(KEYINPUT47), .Z(new_n977));
  NOR2_X1   g0777(.A1(new_n977), .A2(new_n778), .ZN(new_n978));
  INV_X1    g0778(.A(new_n713), .ZN(new_n979));
  OAI221_X1 g0779(.A(new_n724), .B1(new_n229), .B2(new_n340), .C1(new_n241), .C2(new_n979), .ZN(new_n980));
  INV_X1    g0780(.A(new_n723), .ZN(new_n981));
  OAI211_X1 g0781(.A(new_n708), .B(new_n980), .C1(new_n925), .C2(new_n981), .ZN(new_n982));
  NOR2_X1   g0782(.A1(new_n978), .A2(new_n982), .ZN(new_n983));
  INV_X1    g0783(.A(new_n983), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n956), .A2(new_n984), .ZN(G387));
  NAND2_X1  g0785(.A1(new_n951), .A2(new_n952), .ZN(new_n986));
  NAND2_X1  g0786(.A1(new_n986), .A2(new_n707), .ZN(new_n987));
  AOI22_X1  g0787(.A1(G311), .A2(new_n748), .B1(new_n747), .B2(G322), .ZN(new_n988));
  OAI221_X1 g0788(.A(new_n988), .B1(new_n963), .B2(new_n765), .C1(new_n756), .C2(new_n971), .ZN(new_n989));
  XNOR2_X1  g0789(.A(new_n989), .B(KEYINPUT48), .ZN(new_n990));
  OAI221_X1 g0790(.A(new_n990), .B1(new_n730), .B2(new_n734), .C1(new_n732), .C2(new_n739), .ZN(new_n991));
  INV_X1    g0791(.A(KEYINPUT49), .ZN(new_n992));
  OR2_X1    g0792(.A1(new_n991), .A2(new_n992), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n743), .A2(G326), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n991), .A2(new_n992), .ZN(new_n995));
  INV_X1    g0795(.A(new_n728), .ZN(new_n996));
  AOI21_X1  g0796(.A(new_n253), .B1(new_n996), .B2(G116), .ZN(new_n997));
  NAND4_X1  g0797(.A1(new_n993), .A2(new_n994), .A3(new_n995), .A4(new_n997), .ZN(new_n998));
  OAI22_X1  g0798(.A1(new_n365), .A2(new_n767), .B1(new_n773), .B2(new_n285), .ZN(new_n999));
  OAI221_X1 g0799(.A(new_n253), .B1(new_n742), .B2(new_n278), .C1(new_n340), .C2(new_n734), .ZN(new_n1000));
  OAI22_X1  g0800(.A1(new_n729), .A2(new_n213), .B1(new_n739), .B2(new_n258), .ZN(new_n1001));
  NOR3_X1   g0801(.A1(new_n999), .A2(new_n1000), .A3(new_n1001), .ZN(new_n1002));
  OAI221_X1 g0802(.A(new_n1002), .B1(new_n202), .B2(new_n756), .C1(new_n211), .C2(new_n765), .ZN(new_n1003));
  AOI21_X1  g0803(.A(new_n778), .B1(new_n998), .B2(new_n1003), .ZN(new_n1004));
  AOI21_X1  g0804(.A(new_n668), .B1(G68), .B2(G77), .ZN(new_n1005));
  XOR2_X1   g0805(.A(KEYINPUT109), .B(KEYINPUT50), .Z(new_n1006));
  OR3_X1    g0806(.A1(new_n1006), .A2(G50), .A3(new_n285), .ZN(new_n1007));
  OAI21_X1  g0807(.A(new_n1006), .B1(G50), .B2(new_n285), .ZN(new_n1008));
  NAND4_X1  g0808(.A1(new_n1005), .A2(new_n428), .A3(new_n1007), .A4(new_n1008), .ZN(new_n1009));
  AOI21_X1  g0809(.A(new_n979), .B1(new_n237), .B2(G45), .ZN(new_n1010));
  NOR3_X1   g0810(.A1(new_n667), .A2(new_n228), .A3(new_n311), .ZN(new_n1011));
  OAI21_X1  g0811(.A(new_n1009), .B1(new_n1010), .B2(new_n1011), .ZN(new_n1012));
  OAI21_X1  g0812(.A(new_n1012), .B1(G107), .B2(new_n229), .ZN(new_n1013));
  AOI21_X1  g0813(.A(new_n1004), .B1(new_n724), .B2(new_n1013), .ZN(new_n1014));
  OAI211_X1 g0814(.A(new_n1014), .B(new_n708), .C1(new_n914), .C2(new_n981), .ZN(new_n1015));
  OAI21_X1  g0815(.A(new_n666), .B1(new_n986), .B2(new_n703), .ZN(new_n1016));
  OAI211_X1 g0816(.A(new_n987), .B(new_n1015), .C1(new_n1016), .C2(new_n953), .ZN(G393));
  NAND2_X1  g0817(.A1(new_n943), .A2(new_n946), .ZN(new_n1018));
  INV_X1    g0818(.A(new_n953), .ZN(new_n1019));
  AOI21_X1  g0819(.A(new_n665), .B1(new_n1018), .B2(new_n1019), .ZN(new_n1020));
  NAND2_X1  g0820(.A1(new_n1020), .A2(new_n954), .ZN(new_n1021));
  NAND3_X1  g0821(.A1(new_n943), .A2(new_n707), .A3(new_n946), .ZN(new_n1022));
  OAI221_X1 g0822(.A(new_n724), .B1(new_n213), .B2(new_n229), .C1(new_n248), .C2(new_n979), .ZN(new_n1023));
  OAI22_X1  g0823(.A1(new_n756), .A2(new_n365), .B1(new_n278), .B2(new_n767), .ZN(new_n1024));
  XOR2_X1   g0824(.A(new_n1024), .B(KEYINPUT110), .Z(new_n1025));
  XNOR2_X1  g0825(.A(new_n1025), .B(KEYINPUT51), .ZN(new_n1026));
  NOR2_X1   g0826(.A1(new_n773), .A2(new_n202), .ZN(new_n1027));
  AOI21_X1  g0827(.A(new_n311), .B1(new_n743), .B2(G143), .ZN(new_n1028));
  OAI21_X1  g0828(.A(new_n1028), .B1(new_n258), .B2(new_n734), .ZN(new_n1029));
  NOR2_X1   g0829(.A1(new_n739), .A2(new_n211), .ZN(new_n1030));
  NOR4_X1   g0830(.A1(new_n1027), .A2(new_n804), .A3(new_n1029), .A4(new_n1030), .ZN(new_n1031));
  OAI211_X1 g0831(.A(new_n1026), .B(new_n1031), .C1(new_n285), .C2(new_n765), .ZN(new_n1032));
  AOI22_X1  g0832(.A1(G294), .A2(new_n758), .B1(new_n748), .B2(new_n964), .ZN(new_n1033));
  OAI21_X1  g0833(.A(new_n1033), .B1(new_n207), .B2(new_n734), .ZN(new_n1034));
  NOR2_X1   g0834(.A1(new_n1034), .A2(KEYINPUT111), .ZN(new_n1035));
  AOI211_X1 g0835(.A(new_n760), .B(new_n1035), .C1(G283), .C2(new_n790), .ZN(new_n1036));
  OAI21_X1  g0836(.A(new_n311), .B1(new_n742), .B2(new_n751), .ZN(new_n1037));
  AOI21_X1  g0837(.A(new_n1037), .B1(new_n1034), .B2(KEYINPUT111), .ZN(new_n1038));
  AOI22_X1  g0838(.A1(new_n786), .A2(G311), .B1(G317), .B2(new_n747), .ZN(new_n1039));
  INV_X1    g0839(.A(KEYINPUT52), .ZN(new_n1040));
  AND2_X1   g0840(.A1(new_n1039), .A2(new_n1040), .ZN(new_n1041));
  NOR2_X1   g0841(.A1(new_n1039), .A2(new_n1040), .ZN(new_n1042));
  OAI211_X1 g0842(.A(new_n1036), .B(new_n1038), .C1(new_n1041), .C2(new_n1042), .ZN(new_n1043));
  AND2_X1   g0843(.A1(new_n1032), .A2(new_n1043), .ZN(new_n1044));
  OAI211_X1 g0844(.A(new_n708), .B(new_n1023), .C1(new_n1044), .C2(new_n778), .ZN(new_n1045));
  XNOR2_X1  g0845(.A(new_n1045), .B(KEYINPUT112), .ZN(new_n1046));
  OAI21_X1  g0846(.A(new_n1046), .B1(new_n981), .B2(new_n912), .ZN(new_n1047));
  AOI21_X1  g0847(.A(KEYINPUT113), .B1(new_n1022), .B2(new_n1047), .ZN(new_n1048));
  AND3_X1   g0848(.A1(new_n1022), .A2(KEYINPUT113), .A3(new_n1047), .ZN(new_n1049));
  OAI21_X1  g0849(.A(new_n1021), .B1(new_n1048), .B2(new_n1049), .ZN(G390));
  NAND4_X1  g0850(.A1(new_n688), .A2(G330), .A3(new_n690), .A4(new_n812), .ZN(new_n1051));
  INV_X1    g0851(.A(new_n867), .ZN(new_n1052));
  AND2_X1   g0852(.A1(new_n1051), .A2(new_n1052), .ZN(new_n1053));
  NOR2_X1   g0853(.A1(new_n1051), .A2(new_n1052), .ZN(new_n1054));
  NOR2_X1   g0854(.A1(new_n1053), .A2(new_n1054), .ZN(new_n1055));
  NAND3_X1  g0855(.A1(new_n698), .A2(new_n648), .A3(new_n810), .ZN(new_n1056));
  AND2_X1   g0856(.A1(new_n1056), .A2(new_n811), .ZN(new_n1057));
  NAND2_X1  g0857(.A1(new_n1055), .A2(new_n1057), .ZN(new_n1058));
  OAI21_X1  g0858(.A(new_n898), .B1(new_n1053), .B2(new_n1054), .ZN(new_n1059));
  NAND2_X1  g0859(.A1(new_n1058), .A2(new_n1059), .ZN(new_n1060));
  INV_X1    g0860(.A(new_n902), .ZN(new_n1061));
  NAND3_X1  g0861(.A1(new_n691), .A2(new_n418), .A3(G330), .ZN(new_n1062));
  NAND3_X1  g0862(.A1(new_n1060), .A2(new_n1061), .A3(new_n1062), .ZN(new_n1063));
  INV_X1    g0863(.A(new_n891), .ZN(new_n1064));
  OAI21_X1  g0864(.A(new_n1064), .B1(new_n897), .B2(new_n1052), .ZN(new_n1065));
  INV_X1    g0865(.A(KEYINPUT114), .ZN(new_n1066));
  NAND2_X1  g0866(.A1(new_n1065), .A2(new_n1066), .ZN(new_n1067));
  NAND2_X1  g0867(.A1(new_n890), .A2(new_n893), .ZN(new_n1068));
  OAI211_X1 g0868(.A(KEYINPUT114), .B(new_n1064), .C1(new_n897), .C2(new_n1052), .ZN(new_n1069));
  NAND3_X1  g0869(.A1(new_n1067), .A2(new_n1068), .A3(new_n1069), .ZN(new_n1070));
  OAI211_X1 g0870(.A(new_n1064), .B(new_n880), .C1(new_n1057), .C2(new_n1052), .ZN(new_n1071));
  INV_X1    g0871(.A(new_n1054), .ZN(new_n1072));
  AND3_X1   g0872(.A1(new_n1070), .A2(new_n1071), .A3(new_n1072), .ZN(new_n1073));
  AOI21_X1  g0873(.A(new_n1072), .B1(new_n1070), .B2(new_n1071), .ZN(new_n1074));
  OAI21_X1  g0874(.A(new_n1063), .B1(new_n1073), .B2(new_n1074), .ZN(new_n1075));
  NAND2_X1  g0875(.A1(new_n1070), .A2(new_n1071), .ZN(new_n1076));
  NAND2_X1  g0876(.A1(new_n1076), .A2(new_n1054), .ZN(new_n1077));
  NAND3_X1  g0877(.A1(new_n1070), .A2(new_n1071), .A3(new_n1072), .ZN(new_n1078));
  NAND3_X1  g0878(.A1(new_n598), .A2(new_n901), .A3(new_n1062), .ZN(new_n1079));
  AOI21_X1  g0879(.A(new_n1079), .B1(new_n1059), .B2(new_n1058), .ZN(new_n1080));
  NAND3_X1  g0880(.A1(new_n1077), .A2(new_n1078), .A3(new_n1080), .ZN(new_n1081));
  NAND3_X1  g0881(.A1(new_n1075), .A2(new_n1081), .A3(new_n666), .ZN(new_n1082));
  NAND3_X1  g0882(.A1(new_n1077), .A2(new_n707), .A3(new_n1078), .ZN(new_n1083));
  NAND2_X1  g0883(.A1(new_n1068), .A2(new_n814), .ZN(new_n1084));
  OAI21_X1  g0884(.A(new_n708), .B1(new_n816), .B2(new_n374), .ZN(new_n1085));
  XNOR2_X1  g0885(.A(new_n1085), .B(KEYINPUT115), .ZN(new_n1086));
  OAI22_X1  g0886(.A1(new_n486), .A2(new_n773), .B1(new_n767), .B2(new_n730), .ZN(new_n1087));
  NOR2_X1   g0887(.A1(new_n739), .A2(new_n510), .ZN(new_n1088));
  OAI221_X1 g0888(.A(new_n311), .B1(new_n734), .B2(new_n258), .C1(new_n732), .C2(new_n742), .ZN(new_n1089));
  NOR4_X1   g0889(.A1(new_n1087), .A2(new_n793), .A3(new_n1088), .A4(new_n1089), .ZN(new_n1090));
  OAI221_X1 g0890(.A(new_n1090), .B1(new_n213), .B2(new_n765), .C1(new_n207), .C2(new_n756), .ZN(new_n1091));
  NAND2_X1  g0891(.A1(new_n786), .A2(G132), .ZN(new_n1092));
  NAND2_X1  g0892(.A1(new_n748), .A2(G137), .ZN(new_n1093));
  NOR2_X1   g0893(.A1(new_n728), .A2(new_n202), .ZN(new_n1094));
  AOI21_X1  g0894(.A(new_n311), .B1(new_n743), .B2(G125), .ZN(new_n1095));
  OAI21_X1  g0895(.A(new_n1095), .B1(new_n365), .B2(new_n734), .ZN(new_n1096));
  NOR2_X1   g0896(.A1(new_n739), .A2(new_n278), .ZN(new_n1097));
  XOR2_X1   g0897(.A(KEYINPUT116), .B(KEYINPUT53), .Z(new_n1098));
  AOI211_X1 g0898(.A(new_n1094), .B(new_n1096), .C1(new_n1097), .C2(new_n1098), .ZN(new_n1099));
  INV_X1    g0899(.A(G128), .ZN(new_n1100));
  OAI22_X1  g0900(.A1(new_n767), .A2(new_n1100), .B1(new_n1097), .B2(new_n1098), .ZN(new_n1101));
  XOR2_X1   g0901(.A(KEYINPUT54), .B(G143), .Z(new_n1102));
  AOI21_X1  g0902(.A(new_n1101), .B1(new_n758), .B2(new_n1102), .ZN(new_n1103));
  NAND4_X1  g0903(.A1(new_n1092), .A2(new_n1093), .A3(new_n1099), .A4(new_n1103), .ZN(new_n1104));
  AND2_X1   g0904(.A1(new_n1091), .A2(new_n1104), .ZN(new_n1105));
  OAI211_X1 g0905(.A(new_n1084), .B(new_n1086), .C1(new_n778), .C2(new_n1105), .ZN(new_n1106));
  NAND3_X1  g0906(.A1(new_n1082), .A2(new_n1083), .A3(new_n1106), .ZN(G378));
  AOI22_X1  g0907(.A1(G132), .A2(new_n748), .B1(new_n758), .B2(G137), .ZN(new_n1108));
  AOI22_X1  g0908(.A1(new_n747), .A2(G125), .B1(new_n790), .B2(new_n1102), .ZN(new_n1109));
  OAI211_X1 g0909(.A(new_n1108), .B(new_n1109), .C1(new_n756), .C2(new_n1100), .ZN(new_n1110));
  AOI21_X1  g0910(.A(new_n1110), .B1(G150), .B2(new_n794), .ZN(new_n1111));
  XNOR2_X1  g0911(.A(new_n1111), .B(KEYINPUT59), .ZN(new_n1112));
  AOI21_X1  g0912(.A(G41), .B1(new_n996), .B2(G159), .ZN(new_n1113));
  INV_X1    g0913(.A(G124), .ZN(new_n1114));
  AOI21_X1  g0914(.A(new_n742), .B1(KEYINPUT118), .B2(new_n1114), .ZN(new_n1115));
  OAI21_X1  g0915(.A(new_n1115), .B1(KEYINPUT118), .B2(new_n1114), .ZN(new_n1116));
  NAND4_X1  g0916(.A1(new_n1112), .A2(new_n260), .A3(new_n1113), .A4(new_n1116), .ZN(new_n1117));
  OAI21_X1  g0917(.A(new_n202), .B1(new_n309), .B2(G41), .ZN(new_n1118));
  OAI22_X1  g0918(.A1(new_n207), .A2(new_n767), .B1(new_n765), .B2(new_n340), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n996), .A2(G58), .ZN(new_n1120));
  XNOR2_X1  g0920(.A(new_n1120), .B(KEYINPUT117), .ZN(new_n1121));
  OAI211_X1 g0921(.A(new_n1121), .B(new_n311), .C1(new_n730), .C2(new_n742), .ZN(new_n1122));
  OAI221_X1 g0922(.A(new_n261), .B1(new_n211), .B2(new_n734), .C1(new_n739), .C2(new_n258), .ZN(new_n1123));
  NOR3_X1   g0923(.A1(new_n1119), .A2(new_n1122), .A3(new_n1123), .ZN(new_n1124));
  OAI221_X1 g0924(.A(new_n1124), .B1(new_n213), .B2(new_n773), .C1(new_n486), .C2(new_n756), .ZN(new_n1125));
  XNOR2_X1  g0925(.A(new_n1125), .B(KEYINPUT58), .ZN(new_n1126));
  NAND3_X1  g0926(.A1(new_n1117), .A2(new_n1118), .A3(new_n1126), .ZN(new_n1127));
  AOI21_X1  g0927(.A(new_n709), .B1(new_n1127), .B2(new_n720), .ZN(new_n1128));
  INV_X1    g0928(.A(KEYINPUT56), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n835), .A2(new_n293), .ZN(new_n1130));
  INV_X1    g0930(.A(new_n1130), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n306), .A2(new_n1131), .ZN(new_n1132));
  INV_X1    g0932(.A(KEYINPUT55), .ZN(new_n1133));
  NAND4_X1  g0933(.A1(new_n298), .A2(new_n300), .A3(new_n305), .A4(new_n1130), .ZN(new_n1134));
  AND3_X1   g0934(.A1(new_n1132), .A2(new_n1133), .A3(new_n1134), .ZN(new_n1135));
  AOI21_X1  g0935(.A(new_n1133), .B1(new_n1132), .B2(new_n1134), .ZN(new_n1136));
  OAI21_X1  g0936(.A(new_n1129), .B1(new_n1135), .B2(new_n1136), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n1132), .A2(new_n1134), .ZN(new_n1138));
  NAND2_X1  g0938(.A1(new_n1138), .A2(KEYINPUT55), .ZN(new_n1139));
  NAND3_X1  g0939(.A1(new_n1132), .A2(new_n1133), .A3(new_n1134), .ZN(new_n1140));
  NAND3_X1  g0940(.A1(new_n1139), .A2(KEYINPUT56), .A3(new_n1140), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n1137), .A2(new_n1141), .ZN(new_n1142));
  OAI221_X1 g0942(.A(new_n1128), .B1(G50), .B2(new_n816), .C1(new_n1142), .C2(new_n722), .ZN(new_n1143));
  XOR2_X1   g0943(.A(new_n1143), .B(KEYINPUT119), .Z(new_n1144));
  NAND3_X1  g0944(.A1(new_n869), .A2(G330), .A3(new_n881), .ZN(new_n1145));
  NAND2_X1  g0945(.A1(new_n1145), .A2(new_n1142), .ZN(new_n1146));
  AND2_X1   g0946(.A1(new_n1137), .A2(new_n1141), .ZN(new_n1147));
  NAND4_X1  g0947(.A1(new_n1147), .A2(new_n869), .A3(G330), .A4(new_n881), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n1146), .A2(new_n1148), .ZN(new_n1149));
  INV_X1    g0949(.A(new_n900), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n1149), .A2(new_n1150), .ZN(new_n1151));
  INV_X1    g0951(.A(KEYINPUT120), .ZN(new_n1152));
  NAND3_X1  g0952(.A1(new_n1146), .A2(new_n1148), .A3(new_n900), .ZN(new_n1153));
  NAND3_X1  g0953(.A1(new_n1151), .A2(new_n1152), .A3(new_n1153), .ZN(new_n1154));
  NAND4_X1  g0954(.A1(new_n1146), .A2(new_n1148), .A3(new_n900), .A4(KEYINPUT120), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n1154), .A2(new_n1155), .ZN(new_n1156));
  INV_X1    g0956(.A(new_n1156), .ZN(new_n1157));
  AOI21_X1  g0957(.A(new_n1144), .B1(new_n1157), .B2(new_n707), .ZN(new_n1158));
  INV_X1    g0958(.A(KEYINPUT123), .ZN(new_n1159));
  NAND3_X1  g0959(.A1(new_n1151), .A2(new_n1159), .A3(new_n1153), .ZN(new_n1160));
  NAND4_X1  g0960(.A1(new_n1146), .A2(new_n1148), .A3(new_n900), .A4(KEYINPUT123), .ZN(new_n1161));
  AND3_X1   g0961(.A1(new_n1160), .A2(KEYINPUT57), .A3(new_n1161), .ZN(new_n1162));
  XNOR2_X1  g0962(.A(new_n1079), .B(KEYINPUT121), .ZN(new_n1163));
  INV_X1    g0963(.A(new_n1163), .ZN(new_n1164));
  AND3_X1   g0964(.A1(new_n1081), .A2(KEYINPUT122), .A3(new_n1164), .ZN(new_n1165));
  AOI21_X1  g0965(.A(KEYINPUT122), .B1(new_n1081), .B2(new_n1164), .ZN(new_n1166));
  OAI21_X1  g0966(.A(new_n1162), .B1(new_n1165), .B2(new_n1166), .ZN(new_n1167));
  NAND2_X1  g0967(.A1(new_n1167), .A2(new_n666), .ZN(new_n1168));
  INV_X1    g0968(.A(KEYINPUT122), .ZN(new_n1169));
  NOR3_X1   g0969(.A1(new_n1073), .A2(new_n1074), .A3(new_n1063), .ZN(new_n1170));
  OAI21_X1  g0970(.A(new_n1169), .B1(new_n1170), .B2(new_n1163), .ZN(new_n1171));
  NAND3_X1  g0971(.A1(new_n1081), .A2(KEYINPUT122), .A3(new_n1164), .ZN(new_n1172));
  NAND2_X1  g0972(.A1(new_n1171), .A2(new_n1172), .ZN(new_n1173));
  AOI21_X1  g0973(.A(KEYINPUT57), .B1(new_n1173), .B2(new_n1157), .ZN(new_n1174));
  OAI21_X1  g0974(.A(new_n1158), .B1(new_n1168), .B2(new_n1174), .ZN(new_n1175));
  INV_X1    g0975(.A(KEYINPUT124), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n1175), .A2(new_n1176), .ZN(new_n1177));
  AOI21_X1  g0977(.A(new_n1156), .B1(new_n1171), .B2(new_n1172), .ZN(new_n1178));
  OAI211_X1 g0978(.A(new_n1167), .B(new_n666), .C1(new_n1178), .C2(KEYINPUT57), .ZN(new_n1179));
  NAND3_X1  g0979(.A1(new_n1179), .A2(KEYINPUT124), .A3(new_n1158), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n1177), .A2(new_n1180), .ZN(G375));
  NOR2_X1   g0981(.A1(new_n867), .A2(new_n722), .ZN(new_n1182));
  OAI21_X1  g0982(.A(new_n253), .B1(new_n734), .B2(new_n202), .ZN(new_n1183));
  OAI21_X1  g0983(.A(new_n1121), .B1(new_n1100), .B2(new_n742), .ZN(new_n1184));
  AOI211_X1 g0984(.A(new_n1183), .B(new_n1184), .C1(G159), .C2(new_n790), .ZN(new_n1185));
  AOI22_X1  g0985(.A1(G132), .A2(new_n747), .B1(new_n748), .B2(new_n1102), .ZN(new_n1186));
  AND2_X1   g0986(.A1(new_n1185), .A2(new_n1186), .ZN(new_n1187));
  OAI221_X1 g0987(.A(new_n1187), .B1(new_n784), .B2(new_n756), .C1(new_n278), .C2(new_n765), .ZN(new_n1188));
  OAI22_X1  g0988(.A1(new_n486), .A2(new_n765), .B1(new_n767), .B2(new_n732), .ZN(new_n1189));
  OAI22_X1  g0989(.A1(new_n739), .A2(new_n213), .B1(new_n340), .B2(new_n734), .ZN(new_n1190));
  OAI221_X1 g0990(.A(new_n311), .B1(new_n740), .B2(new_n742), .C1(new_n729), .C2(new_n258), .ZN(new_n1191));
  NOR3_X1   g0991(.A1(new_n1189), .A2(new_n1190), .A3(new_n1191), .ZN(new_n1192));
  OAI221_X1 g0992(.A(new_n1192), .B1(new_n207), .B2(new_n773), .C1(new_n730), .C2(new_n756), .ZN(new_n1193));
  AOI21_X1  g0993(.A(new_n778), .B1(new_n1188), .B2(new_n1193), .ZN(new_n1194));
  NOR2_X1   g0994(.A1(new_n816), .A2(G68), .ZN(new_n1195));
  NOR4_X1   g0995(.A1(new_n1182), .A2(new_n709), .A3(new_n1194), .A4(new_n1195), .ZN(new_n1196));
  AOI21_X1  g0996(.A(new_n1196), .B1(new_n1060), .B2(new_n707), .ZN(new_n1197));
  NAND3_X1  g0997(.A1(new_n1079), .A2(new_n1058), .A3(new_n1059), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(new_n1198), .A2(new_n933), .ZN(new_n1199));
  OAI21_X1  g0999(.A(new_n1197), .B1(new_n1199), .B2(new_n1080), .ZN(G381));
  INV_X1    g1000(.A(G378), .ZN(new_n1201));
  NAND3_X1  g1001(.A1(new_n1177), .A2(new_n1201), .A3(new_n1180), .ZN(new_n1202));
  OR3_X1    g1002(.A1(new_n1202), .A2(G384), .A3(G381), .ZN(new_n1203));
  OR4_X1    g1003(.A1(G396), .A2(G387), .A3(G393), .A4(G390), .ZN(new_n1204));
  OR2_X1    g1004(.A1(new_n1203), .A2(new_n1204), .ZN(G407));
  OAI221_X1 g1005(.A(G213), .B1(G343), .B2(new_n1202), .C1(new_n1203), .C2(new_n1204), .ZN(G409));
  INV_X1    g1006(.A(KEYINPUT60), .ZN(new_n1207));
  AOI21_X1  g1007(.A(new_n665), .B1(new_n1198), .B2(new_n1207), .ZN(new_n1208));
  OAI211_X1 g1008(.A(new_n1208), .B(new_n1063), .C1(new_n1207), .C2(new_n1198), .ZN(new_n1209));
  AND3_X1   g1009(.A1(new_n1209), .A2(G384), .A3(new_n1197), .ZN(new_n1210));
  AOI21_X1  g1010(.A(G384), .B1(new_n1209), .B2(new_n1197), .ZN(new_n1211));
  NOR2_X1   g1011(.A1(new_n1210), .A2(new_n1211), .ZN(new_n1212));
  NAND3_X1  g1012(.A1(new_n637), .A2(G213), .A3(G2897), .ZN(new_n1213));
  XOR2_X1   g1013(.A(new_n1213), .B(KEYINPUT125), .Z(new_n1214));
  XOR2_X1   g1014(.A(new_n1212), .B(new_n1214), .Z(new_n1215));
  NAND2_X1  g1015(.A1(new_n1175), .A2(G378), .ZN(new_n1216));
  AND2_X1   g1016(.A1(new_n1201), .A2(new_n1143), .ZN(new_n1217));
  AND3_X1   g1017(.A1(new_n1160), .A2(new_n707), .A3(new_n1161), .ZN(new_n1218));
  AOI21_X1  g1018(.A(new_n1218), .B1(new_n1178), .B2(new_n933), .ZN(new_n1219));
  AOI22_X1  g1019(.A1(new_n1217), .A2(new_n1219), .B1(G213), .B2(new_n637), .ZN(new_n1220));
  AOI21_X1  g1020(.A(new_n1215), .B1(new_n1216), .B2(new_n1220), .ZN(new_n1221));
  NOR2_X1   g1021(.A1(new_n1221), .A2(KEYINPUT61), .ZN(new_n1222));
  NAND3_X1  g1022(.A1(new_n1216), .A2(new_n1220), .A3(new_n1212), .ZN(new_n1223));
  XOR2_X1   g1023(.A(KEYINPUT126), .B(KEYINPUT62), .Z(new_n1224));
  NAND2_X1  g1024(.A1(new_n1223), .A2(new_n1224), .ZN(new_n1225));
  NOR2_X1   g1025(.A1(KEYINPUT126), .A2(KEYINPUT62), .ZN(new_n1226));
  NAND4_X1  g1026(.A1(new_n1216), .A2(new_n1220), .A3(new_n1212), .A4(new_n1226), .ZN(new_n1227));
  NAND3_X1  g1027(.A1(new_n1222), .A2(new_n1225), .A3(new_n1227), .ZN(new_n1228));
  INV_X1    g1028(.A(KEYINPUT127), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n1022), .A2(new_n1047), .ZN(new_n1230));
  INV_X1    g1030(.A(KEYINPUT113), .ZN(new_n1231));
  NAND2_X1  g1031(.A1(new_n1230), .A2(new_n1231), .ZN(new_n1232));
  NAND3_X1  g1032(.A1(new_n1022), .A2(KEYINPUT113), .A3(new_n1047), .ZN(new_n1233));
  AOI22_X1  g1033(.A1(new_n1232), .A2(new_n1233), .B1(new_n954), .B2(new_n1020), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n931), .A2(new_n932), .ZN(new_n1235));
  NAND2_X1  g1035(.A1(new_n954), .A2(new_n703), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n1236), .A2(new_n933), .ZN(new_n1237));
  AOI21_X1  g1037(.A(new_n1235), .B1(new_n1237), .B2(new_n706), .ZN(new_n1238));
  OAI21_X1  g1038(.A(new_n1234), .B1(new_n1238), .B2(new_n983), .ZN(new_n1239));
  XNOR2_X1  g1039(.A(G393), .B(new_n782), .ZN(new_n1240));
  NAND3_X1  g1040(.A1(G390), .A2(new_n984), .A3(new_n956), .ZN(new_n1241));
  AND3_X1   g1041(.A1(new_n1239), .A2(new_n1240), .A3(new_n1241), .ZN(new_n1242));
  AOI21_X1  g1042(.A(new_n1240), .B1(new_n1239), .B2(new_n1241), .ZN(new_n1243));
  OAI21_X1  g1043(.A(new_n1229), .B1(new_n1242), .B2(new_n1243), .ZN(new_n1244));
  NAND2_X1  g1044(.A1(new_n1239), .A2(new_n1241), .ZN(new_n1245));
  INV_X1    g1045(.A(new_n1240), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(new_n1245), .A2(new_n1246), .ZN(new_n1247));
  NAND3_X1  g1047(.A1(new_n1239), .A2(new_n1241), .A3(new_n1240), .ZN(new_n1248));
  NAND3_X1  g1048(.A1(new_n1247), .A2(KEYINPUT127), .A3(new_n1248), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n1244), .A2(new_n1249), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(new_n1228), .A2(new_n1250), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n1247), .A2(new_n1248), .ZN(new_n1252));
  INV_X1    g1052(.A(new_n1223), .ZN(new_n1253));
  AOI21_X1  g1053(.A(new_n1252), .B1(new_n1253), .B2(KEYINPUT63), .ZN(new_n1254));
  INV_X1    g1054(.A(KEYINPUT61), .ZN(new_n1255));
  INV_X1    g1055(.A(KEYINPUT63), .ZN(new_n1256));
  OAI21_X1  g1056(.A(new_n1223), .B1(new_n1221), .B2(new_n1256), .ZN(new_n1257));
  NAND3_X1  g1057(.A1(new_n1254), .A2(new_n1255), .A3(new_n1257), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(new_n1251), .A2(new_n1258), .ZN(G405));
  INV_X1    g1059(.A(new_n1212), .ZN(new_n1260));
  AND3_X1   g1060(.A1(new_n1202), .A2(new_n1216), .A3(new_n1260), .ZN(new_n1261));
  AOI21_X1  g1061(.A(new_n1260), .B1(new_n1202), .B2(new_n1216), .ZN(new_n1262));
  NOR3_X1   g1062(.A1(new_n1261), .A2(new_n1262), .A3(new_n1250), .ZN(new_n1263));
  AND2_X1   g1063(.A1(new_n1244), .A2(new_n1249), .ZN(new_n1264));
  AND3_X1   g1064(.A1(new_n1179), .A2(KEYINPUT124), .A3(new_n1158), .ZN(new_n1265));
  AOI21_X1  g1065(.A(KEYINPUT124), .B1(new_n1179), .B2(new_n1158), .ZN(new_n1266));
  NOR3_X1   g1066(.A1(new_n1265), .A2(new_n1266), .A3(G378), .ZN(new_n1267));
  INV_X1    g1067(.A(new_n1216), .ZN(new_n1268));
  OAI21_X1  g1068(.A(new_n1212), .B1(new_n1267), .B2(new_n1268), .ZN(new_n1269));
  NAND3_X1  g1069(.A1(new_n1202), .A2(new_n1216), .A3(new_n1260), .ZN(new_n1270));
  AOI21_X1  g1070(.A(new_n1264), .B1(new_n1269), .B2(new_n1270), .ZN(new_n1271));
  NOR2_X1   g1071(.A1(new_n1263), .A2(new_n1271), .ZN(G402));
endmodule


