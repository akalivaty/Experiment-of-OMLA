//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 0 0 1 1 1 1 0 1 1 1 0 0 1 0 0 0 1 0 1 1 0 0 0 1 1 0 1 1 1 0 1 0 0 1 0 0 1 1 1 1 0 1 0 0 1 1 1 1 1 1 0 0 0 1 0 1 1 1 0 1 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:33:43 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n447, new_n448, new_n452, new_n453, new_n454, new_n455,
    new_n456, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n521, new_n522, new_n523, new_n524, new_n525,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n531, new_n532,
    new_n534, new_n535, new_n536, new_n537, new_n538, new_n539, new_n540,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n551, new_n552, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n571, new_n572, new_n573, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n581, new_n582, new_n583, new_n584,
    new_n585, new_n586, new_n587, new_n588, new_n589, new_n591, new_n592,
    new_n593, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n608, new_n609,
    new_n612, new_n613, new_n615, new_n616, new_n617, new_n619, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1217, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  XOR2_X1   g005(.A(KEYINPUT64), .B(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  AND2_X1   g016(.A1(G2072), .A2(G2078), .ZN(new_n442));
  NAND3_X1  g017(.A1(new_n442), .A2(G2084), .A3(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XNOR2_X1  g022(.A(new_n447), .B(KEYINPUT65), .ZN(new_n448));
  XNOR2_X1  g023(.A(new_n448), .B(KEYINPUT1), .ZN(G223));
  NAND3_X1  g024(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g025(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g026(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n452));
  XNOR2_X1  g027(.A(new_n452), .B(KEYINPUT2), .ZN(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NOR4_X1   g029(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n455));
  INV_X1    g030(.A(new_n455), .ZN(new_n456));
  NOR2_X1   g031(.A1(new_n454), .A2(new_n456), .ZN(G325));
  INV_X1    g032(.A(G325), .ZN(G261));
  AOI22_X1  g033(.A1(new_n454), .A2(G2106), .B1(G567), .B2(new_n456), .ZN(G319));
  INV_X1    g034(.A(G125), .ZN(new_n460));
  INV_X1    g035(.A(KEYINPUT3), .ZN(new_n461));
  INV_X1    g036(.A(G2104), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  NAND2_X1  g038(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n464));
  AOI21_X1  g039(.A(new_n460), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  AND2_X1   g040(.A1(G113), .A2(G2104), .ZN(new_n466));
  OAI21_X1  g041(.A(G2105), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  INV_X1    g042(.A(G2105), .ZN(new_n468));
  INV_X1    g043(.A(G137), .ZN(new_n469));
  AOI21_X1  g044(.A(new_n469), .B1(new_n463), .B2(new_n464), .ZN(new_n470));
  AND2_X1   g045(.A1(G101), .A2(G2104), .ZN(new_n471));
  OAI21_X1  g046(.A(new_n468), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  AND2_X1   g047(.A1(new_n467), .A2(new_n472), .ZN(G160));
  AOI21_X1  g048(.A(new_n468), .B1(new_n463), .B2(new_n464), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n474), .A2(G124), .ZN(new_n475));
  XOR2_X1   g050(.A(new_n475), .B(KEYINPUT66), .Z(new_n476));
  AOI21_X1  g051(.A(G2105), .B1(new_n463), .B2(new_n464), .ZN(new_n477));
  OR2_X1    g052(.A1(G100), .A2(G2105), .ZN(new_n478));
  INV_X1    g053(.A(G112), .ZN(new_n479));
  AOI21_X1  g054(.A(new_n462), .B1(new_n479), .B2(G2105), .ZN(new_n480));
  AOI22_X1  g055(.A1(new_n477), .A2(G136), .B1(new_n478), .B2(new_n480), .ZN(new_n481));
  AND2_X1   g056(.A1(new_n476), .A2(new_n481), .ZN(G162));
  INV_X1    g057(.A(G114), .ZN(new_n483));
  AOI21_X1  g058(.A(new_n462), .B1(new_n483), .B2(G2105), .ZN(new_n484));
  NOR2_X1   g059(.A1(G102), .A2(G2105), .ZN(new_n485));
  INV_X1    g060(.A(new_n485), .ZN(new_n486));
  NAND3_X1  g061(.A1(new_n484), .A2(KEYINPUT67), .A3(new_n486), .ZN(new_n487));
  INV_X1    g062(.A(KEYINPUT67), .ZN(new_n488));
  OAI21_X1  g063(.A(G2104), .B1(new_n468), .B2(G114), .ZN(new_n489));
  OAI21_X1  g064(.A(new_n488), .B1(new_n489), .B2(new_n485), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n487), .A2(new_n490), .ZN(new_n491));
  NAND2_X1  g066(.A1(new_n474), .A2(G126), .ZN(new_n492));
  AND2_X1   g067(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n493));
  NOR2_X1   g068(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n494));
  OAI211_X1 g069(.A(G138), .B(new_n468), .C1(new_n493), .C2(new_n494), .ZN(new_n495));
  INV_X1    g070(.A(KEYINPUT4), .ZN(new_n496));
  NAND2_X1  g071(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  XNOR2_X1  g072(.A(KEYINPUT3), .B(G2104), .ZN(new_n498));
  NAND4_X1  g073(.A1(new_n498), .A2(KEYINPUT4), .A3(G138), .A4(new_n468), .ZN(new_n499));
  NAND4_X1  g074(.A1(new_n491), .A2(new_n492), .A3(new_n497), .A4(new_n499), .ZN(new_n500));
  INV_X1    g075(.A(new_n500), .ZN(G164));
  XNOR2_X1  g076(.A(KEYINPUT5), .B(G543), .ZN(new_n502));
  INV_X1    g077(.A(G651), .ZN(new_n503));
  NAND2_X1  g078(.A1(new_n503), .A2(KEYINPUT6), .ZN(new_n504));
  INV_X1    g079(.A(KEYINPUT6), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n505), .A2(G651), .ZN(new_n506));
  NAND3_X1  g081(.A1(new_n502), .A2(new_n504), .A3(new_n506), .ZN(new_n507));
  NOR2_X1   g082(.A1(new_n507), .A2(KEYINPUT69), .ZN(new_n508));
  INV_X1    g083(.A(KEYINPUT69), .ZN(new_n509));
  AND2_X1   g084(.A1(new_n504), .A2(new_n506), .ZN(new_n510));
  AOI21_X1  g085(.A(new_n509), .B1(new_n510), .B2(new_n502), .ZN(new_n511));
  NOR2_X1   g086(.A1(new_n508), .A2(new_n511), .ZN(new_n512));
  XNOR2_X1  g087(.A(KEYINPUT70), .B(G88), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  AOI22_X1  g089(.A1(new_n502), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n515));
  OR2_X1    g090(.A1(new_n515), .A2(new_n503), .ZN(new_n516));
  NAND3_X1  g091(.A1(new_n510), .A2(G50), .A3(G543), .ZN(new_n517));
  XNOR2_X1  g092(.A(new_n517), .B(KEYINPUT68), .ZN(new_n518));
  NAND3_X1  g093(.A1(new_n514), .A2(new_n516), .A3(new_n518), .ZN(new_n519));
  INV_X1    g094(.A(new_n519), .ZN(G166));
  NAND3_X1  g095(.A1(new_n502), .A2(G63), .A3(G651), .ZN(new_n521));
  XNOR2_X1  g096(.A(new_n521), .B(KEYINPUT71), .ZN(new_n522));
  NAND3_X1  g097(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n523));
  XOR2_X1   g098(.A(new_n523), .B(KEYINPUT7), .Z(new_n524));
  AND3_X1   g099(.A1(new_n504), .A2(new_n506), .A3(G543), .ZN(new_n525));
  AOI21_X1  g100(.A(new_n524), .B1(G51), .B2(new_n525), .ZN(new_n526));
  NAND2_X1  g101(.A1(new_n522), .A2(new_n526), .ZN(new_n527));
  NAND2_X1  g102(.A1(new_n507), .A2(KEYINPUT69), .ZN(new_n528));
  NAND3_X1  g103(.A1(new_n510), .A2(new_n509), .A3(new_n502), .ZN(new_n529));
  NAND2_X1  g104(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  XNOR2_X1  g105(.A(KEYINPUT72), .B(G89), .ZN(new_n531));
  NOR2_X1   g106(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  NOR2_X1   g107(.A1(new_n527), .A2(new_n532), .ZN(G168));
  XNOR2_X1  g108(.A(KEYINPUT73), .B(G90), .ZN(new_n534));
  NAND2_X1  g109(.A1(new_n512), .A2(new_n534), .ZN(new_n535));
  NAND2_X1  g110(.A1(G77), .A2(G543), .ZN(new_n536));
  INV_X1    g111(.A(new_n502), .ZN(new_n537));
  INV_X1    g112(.A(G64), .ZN(new_n538));
  OAI21_X1  g113(.A(new_n536), .B1(new_n537), .B2(new_n538), .ZN(new_n539));
  AOI22_X1  g114(.A1(new_n539), .A2(G651), .B1(G52), .B2(new_n525), .ZN(new_n540));
  AND2_X1   g115(.A1(new_n535), .A2(new_n540), .ZN(G171));
  NAND2_X1  g116(.A1(new_n512), .A2(G81), .ZN(new_n542));
  NAND2_X1  g117(.A1(G68), .A2(G543), .ZN(new_n543));
  INV_X1    g118(.A(G56), .ZN(new_n544));
  OAI21_X1  g119(.A(new_n543), .B1(new_n537), .B2(new_n544), .ZN(new_n545));
  AOI22_X1  g120(.A1(new_n545), .A2(G651), .B1(G43), .B2(new_n525), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n542), .A2(new_n546), .ZN(new_n547));
  INV_X1    g122(.A(new_n547), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n548), .A2(G860), .ZN(G153));
  NAND4_X1  g124(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g125(.A1(G1), .A2(G3), .ZN(new_n551));
  XNOR2_X1  g126(.A(new_n551), .B(KEYINPUT8), .ZN(new_n552));
  NAND4_X1  g127(.A1(G319), .A2(G483), .A3(G661), .A4(new_n552), .ZN(G188));
  NAND2_X1  g128(.A1(new_n525), .A2(G53), .ZN(new_n554));
  OR2_X1    g129(.A1(new_n554), .A2(KEYINPUT9), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n554), .A2(KEYINPUT9), .ZN(new_n556));
  NAND2_X1  g131(.A1(G78), .A2(G543), .ZN(new_n557));
  INV_X1    g132(.A(G65), .ZN(new_n558));
  OAI21_X1  g133(.A(new_n557), .B1(new_n537), .B2(new_n558), .ZN(new_n559));
  AOI22_X1  g134(.A1(new_n555), .A2(new_n556), .B1(G651), .B2(new_n559), .ZN(new_n560));
  INV_X1    g135(.A(new_n560), .ZN(new_n561));
  INV_X1    g136(.A(G91), .ZN(new_n562));
  INV_X1    g137(.A(KEYINPUT74), .ZN(new_n563));
  OAI21_X1  g138(.A(new_n563), .B1(new_n508), .B2(new_n511), .ZN(new_n564));
  NAND3_X1  g139(.A1(new_n528), .A2(KEYINPUT74), .A3(new_n529), .ZN(new_n565));
  AOI21_X1  g140(.A(new_n562), .B1(new_n564), .B2(new_n565), .ZN(new_n566));
  NOR2_X1   g141(.A1(new_n561), .A2(new_n566), .ZN(new_n567));
  INV_X1    g142(.A(new_n567), .ZN(G299));
  NAND2_X1  g143(.A1(new_n535), .A2(new_n540), .ZN(G301));
  INV_X1    g144(.A(G168), .ZN(G286));
  INV_X1    g145(.A(KEYINPUT75), .ZN(new_n571));
  NAND2_X1  g146(.A1(new_n519), .A2(new_n571), .ZN(new_n572));
  NAND4_X1  g147(.A1(new_n514), .A2(new_n518), .A3(KEYINPUT75), .A4(new_n516), .ZN(new_n573));
  AND2_X1   g148(.A1(new_n572), .A2(new_n573), .ZN(G303));
  AND3_X1   g149(.A1(new_n528), .A2(KEYINPUT74), .A3(new_n529), .ZN(new_n575));
  AOI21_X1  g150(.A(KEYINPUT74), .B1(new_n528), .B2(new_n529), .ZN(new_n576));
  OAI21_X1  g151(.A(G87), .B1(new_n575), .B2(new_n576), .ZN(new_n577));
  OR2_X1    g152(.A1(new_n502), .A2(G74), .ZN(new_n578));
  AOI22_X1  g153(.A1(new_n578), .A2(G651), .B1(new_n525), .B2(G49), .ZN(new_n579));
  NAND2_X1  g154(.A1(new_n577), .A2(new_n579), .ZN(G288));
  INV_X1    g155(.A(G86), .ZN(new_n581));
  AOI21_X1  g156(.A(new_n581), .B1(new_n564), .B2(new_n565), .ZN(new_n582));
  NAND2_X1  g157(.A1(G73), .A2(G543), .ZN(new_n583));
  INV_X1    g158(.A(G61), .ZN(new_n584));
  OAI21_X1  g159(.A(new_n583), .B1(new_n537), .B2(new_n584), .ZN(new_n585));
  NAND2_X1  g160(.A1(new_n585), .A2(G651), .ZN(new_n586));
  NAND2_X1  g161(.A1(new_n525), .A2(G48), .ZN(new_n587));
  NAND2_X1  g162(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  NOR2_X1   g163(.A1(new_n582), .A2(new_n588), .ZN(new_n589));
  INV_X1    g164(.A(new_n589), .ZN(G305));
  NAND2_X1  g165(.A1(new_n525), .A2(G47), .ZN(new_n591));
  AOI22_X1  g166(.A1(new_n502), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n592));
  INV_X1    g167(.A(G85), .ZN(new_n593));
  OAI221_X1 g168(.A(new_n591), .B1(new_n503), .B2(new_n592), .C1(new_n530), .C2(new_n593), .ZN(G290));
  NAND2_X1  g169(.A1(G301), .A2(G868), .ZN(new_n595));
  NAND2_X1  g170(.A1(new_n525), .A2(G54), .ZN(new_n596));
  XOR2_X1   g171(.A(KEYINPUT76), .B(G66), .Z(new_n597));
  AOI22_X1  g172(.A1(new_n597), .A2(new_n502), .B1(G79), .B2(G543), .ZN(new_n598));
  OAI21_X1  g173(.A(new_n596), .B1(new_n598), .B2(new_n503), .ZN(new_n599));
  INV_X1    g174(.A(KEYINPUT10), .ZN(new_n600));
  NOR2_X1   g175(.A1(new_n575), .A2(new_n576), .ZN(new_n601));
  INV_X1    g176(.A(G92), .ZN(new_n602));
  OAI21_X1  g177(.A(new_n600), .B1(new_n601), .B2(new_n602), .ZN(new_n603));
  OAI211_X1 g178(.A(KEYINPUT10), .B(G92), .C1(new_n575), .C2(new_n576), .ZN(new_n604));
  AOI21_X1  g179(.A(new_n599), .B1(new_n603), .B2(new_n604), .ZN(new_n605));
  OAI21_X1  g180(.A(new_n595), .B1(new_n605), .B2(G868), .ZN(G284));
  OAI21_X1  g181(.A(new_n595), .B1(new_n605), .B2(G868), .ZN(G321));
  NAND2_X1  g182(.A1(G286), .A2(G868), .ZN(new_n608));
  XOR2_X1   g183(.A(new_n608), .B(KEYINPUT77), .Z(new_n609));
  OAI21_X1  g184(.A(new_n609), .B1(G868), .B2(new_n567), .ZN(G297));
  OAI21_X1  g185(.A(new_n609), .B1(G868), .B2(new_n567), .ZN(G280));
  INV_X1    g186(.A(G559), .ZN(new_n612));
  OAI21_X1  g187(.A(new_n605), .B1(new_n612), .B2(G860), .ZN(new_n613));
  XNOR2_X1  g188(.A(new_n613), .B(KEYINPUT78), .ZN(G148));
  NOR2_X1   g189(.A1(new_n548), .A2(G868), .ZN(new_n615));
  NAND2_X1  g190(.A1(new_n605), .A2(new_n612), .ZN(new_n616));
  AOI21_X1  g191(.A(new_n615), .B1(new_n616), .B2(G868), .ZN(new_n617));
  XNOR2_X1  g192(.A(new_n617), .B(KEYINPUT79), .ZN(G323));
  XNOR2_X1  g193(.A(G323), .B(KEYINPUT80), .ZN(new_n619));
  XOR2_X1   g194(.A(new_n619), .B(KEYINPUT11), .Z(G282));
  NAND2_X1  g195(.A1(new_n477), .A2(G2104), .ZN(new_n621));
  XNOR2_X1  g196(.A(new_n621), .B(KEYINPUT12), .ZN(new_n622));
  XNOR2_X1  g197(.A(new_n622), .B(KEYINPUT13), .ZN(new_n623));
  INV_X1    g198(.A(G2100), .ZN(new_n624));
  OR2_X1    g199(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  NAND2_X1  g200(.A1(new_n623), .A2(new_n624), .ZN(new_n626));
  NAND2_X1  g201(.A1(new_n477), .A2(G135), .ZN(new_n627));
  NAND2_X1  g202(.A1(new_n474), .A2(G123), .ZN(new_n628));
  NOR2_X1   g203(.A1(G99), .A2(G2105), .ZN(new_n629));
  OAI21_X1  g204(.A(G2104), .B1(new_n468), .B2(G111), .ZN(new_n630));
  OAI211_X1 g205(.A(new_n627), .B(new_n628), .C1(new_n629), .C2(new_n630), .ZN(new_n631));
  INV_X1    g206(.A(G2096), .ZN(new_n632));
  XNOR2_X1  g207(.A(new_n631), .B(new_n632), .ZN(new_n633));
  NAND3_X1  g208(.A1(new_n625), .A2(new_n626), .A3(new_n633), .ZN(G156));
  XOR2_X1   g209(.A(G2451), .B(G2454), .Z(new_n635));
  XNOR2_X1  g210(.A(new_n635), .B(KEYINPUT16), .ZN(new_n636));
  XNOR2_X1  g211(.A(G1341), .B(G1348), .ZN(new_n637));
  XNOR2_X1  g212(.A(new_n636), .B(new_n637), .ZN(new_n638));
  XNOR2_X1  g213(.A(G2443), .B(G2446), .ZN(new_n639));
  XNOR2_X1  g214(.A(new_n638), .B(new_n639), .ZN(new_n640));
  XNOR2_X1  g215(.A(G2427), .B(G2438), .ZN(new_n641));
  XNOR2_X1  g216(.A(new_n641), .B(G2430), .ZN(new_n642));
  XNOR2_X1  g217(.A(KEYINPUT15), .B(G2435), .ZN(new_n643));
  OR2_X1    g218(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  NAND2_X1  g219(.A1(new_n642), .A2(new_n643), .ZN(new_n645));
  NAND3_X1  g220(.A1(new_n644), .A2(new_n645), .A3(KEYINPUT14), .ZN(new_n646));
  INV_X1    g221(.A(new_n646), .ZN(new_n647));
  OR2_X1    g222(.A1(new_n640), .A2(new_n647), .ZN(new_n648));
  NAND2_X1  g223(.A1(new_n640), .A2(new_n647), .ZN(new_n649));
  NAND3_X1  g224(.A1(new_n648), .A2(new_n649), .A3(G14), .ZN(new_n650));
  XNOR2_X1  g225(.A(new_n650), .B(KEYINPUT81), .ZN(G401));
  XOR2_X1   g226(.A(G2084), .B(G2090), .Z(new_n652));
  XNOR2_X1  g227(.A(G2072), .B(G2078), .ZN(new_n653));
  XNOR2_X1  g228(.A(G2067), .B(G2678), .ZN(new_n654));
  NAND3_X1  g229(.A1(new_n652), .A2(new_n653), .A3(new_n654), .ZN(new_n655));
  XOR2_X1   g230(.A(new_n655), .B(KEYINPUT18), .Z(new_n656));
  OR2_X1    g231(.A1(new_n653), .A2(KEYINPUT82), .ZN(new_n657));
  NAND2_X1  g232(.A1(new_n653), .A2(KEYINPUT82), .ZN(new_n658));
  INV_X1    g233(.A(new_n654), .ZN(new_n659));
  NAND3_X1  g234(.A1(new_n657), .A2(new_n658), .A3(new_n659), .ZN(new_n660));
  INV_X1    g235(.A(new_n652), .ZN(new_n661));
  XOR2_X1   g236(.A(new_n653), .B(KEYINPUT17), .Z(new_n662));
  OAI211_X1 g237(.A(new_n660), .B(new_n661), .C1(new_n662), .C2(new_n659), .ZN(new_n663));
  NAND3_X1  g238(.A1(new_n662), .A2(new_n659), .A3(new_n652), .ZN(new_n664));
  NAND3_X1  g239(.A1(new_n656), .A2(new_n663), .A3(new_n664), .ZN(new_n665));
  XNOR2_X1  g240(.A(new_n665), .B(new_n632), .ZN(new_n666));
  XNOR2_X1  g241(.A(new_n666), .B(G2100), .ZN(G227));
  XOR2_X1   g242(.A(G1971), .B(G1976), .Z(new_n668));
  XNOR2_X1  g243(.A(new_n668), .B(KEYINPUT19), .ZN(new_n669));
  XNOR2_X1  g244(.A(G1956), .B(G2474), .ZN(new_n670));
  XNOR2_X1  g245(.A(G1961), .B(G1966), .ZN(new_n671));
  NOR2_X1   g246(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  AND2_X1   g247(.A1(new_n670), .A2(new_n671), .ZN(new_n673));
  NOR3_X1   g248(.A1(new_n669), .A2(new_n672), .A3(new_n673), .ZN(new_n674));
  NAND2_X1  g249(.A1(new_n669), .A2(new_n672), .ZN(new_n675));
  XOR2_X1   g250(.A(new_n675), .B(KEYINPUT20), .Z(new_n676));
  AOI211_X1 g251(.A(new_n674), .B(new_n676), .C1(new_n669), .C2(new_n673), .ZN(new_n677));
  XOR2_X1   g252(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n678));
  XNOR2_X1  g253(.A(new_n678), .B(KEYINPUT83), .ZN(new_n679));
  INV_X1    g254(.A(new_n679), .ZN(new_n680));
  XNOR2_X1  g255(.A(new_n677), .B(new_n680), .ZN(new_n681));
  XOR2_X1   g256(.A(G1981), .B(G1986), .Z(new_n682));
  XNOR2_X1  g257(.A(new_n681), .B(new_n682), .ZN(new_n683));
  XNOR2_X1  g258(.A(G1991), .B(G1996), .ZN(new_n684));
  XNOR2_X1  g259(.A(new_n683), .B(new_n684), .ZN(new_n685));
  INV_X1    g260(.A(new_n685), .ZN(G229));
  INV_X1    g261(.A(G16), .ZN(new_n687));
  NAND2_X1  g262(.A1(new_n687), .A2(G22), .ZN(new_n688));
  OAI21_X1  g263(.A(new_n688), .B1(G166), .B2(new_n687), .ZN(new_n689));
  XNOR2_X1  g264(.A(new_n689), .B(G1971), .ZN(new_n690));
  NAND2_X1  g265(.A1(new_n687), .A2(G23), .ZN(new_n691));
  INV_X1    g266(.A(G288), .ZN(new_n692));
  OAI21_X1  g267(.A(new_n691), .B1(new_n692), .B2(new_n687), .ZN(new_n693));
  XOR2_X1   g268(.A(KEYINPUT33), .B(G1976), .Z(new_n694));
  AOI21_X1  g269(.A(new_n690), .B1(new_n693), .B2(new_n694), .ZN(new_n695));
  NAND2_X1  g270(.A1(new_n687), .A2(G6), .ZN(new_n696));
  OAI21_X1  g271(.A(new_n696), .B1(new_n589), .B2(new_n687), .ZN(new_n697));
  XOR2_X1   g272(.A(KEYINPUT32), .B(G1981), .Z(new_n698));
  XNOR2_X1  g273(.A(new_n697), .B(new_n698), .ZN(new_n699));
  OAI211_X1 g274(.A(new_n695), .B(new_n699), .C1(new_n693), .C2(new_n694), .ZN(new_n700));
  OR2_X1    g275(.A1(new_n700), .A2(KEYINPUT34), .ZN(new_n701));
  NAND2_X1  g276(.A1(new_n700), .A2(KEYINPUT34), .ZN(new_n702));
  NAND2_X1  g277(.A1(new_n477), .A2(G131), .ZN(new_n703));
  NAND2_X1  g278(.A1(new_n474), .A2(G119), .ZN(new_n704));
  NOR2_X1   g279(.A1(G95), .A2(G2105), .ZN(new_n705));
  OAI21_X1  g280(.A(G2104), .B1(new_n468), .B2(G107), .ZN(new_n706));
  OAI211_X1 g281(.A(new_n703), .B(new_n704), .C1(new_n705), .C2(new_n706), .ZN(new_n707));
  XOR2_X1   g282(.A(KEYINPUT84), .B(G29), .Z(new_n708));
  INV_X1    g283(.A(new_n708), .ZN(new_n709));
  MUX2_X1   g284(.A(G25), .B(new_n707), .S(new_n709), .Z(new_n710));
  XNOR2_X1  g285(.A(KEYINPUT35), .B(G1991), .ZN(new_n711));
  XOR2_X1   g286(.A(new_n710), .B(new_n711), .Z(new_n712));
  MUX2_X1   g287(.A(G24), .B(G290), .S(G16), .Z(new_n713));
  INV_X1    g288(.A(G1986), .ZN(new_n714));
  XNOR2_X1  g289(.A(new_n713), .B(new_n714), .ZN(new_n715));
  INV_X1    g290(.A(new_n715), .ZN(new_n716));
  OAI21_X1  g291(.A(new_n712), .B1(new_n716), .B2(KEYINPUT85), .ZN(new_n717));
  AOI21_X1  g292(.A(new_n717), .B1(KEYINPUT85), .B2(new_n716), .ZN(new_n718));
  NAND3_X1  g293(.A1(new_n701), .A2(new_n702), .A3(new_n718), .ZN(new_n719));
  XOR2_X1   g294(.A(new_n719), .B(KEYINPUT36), .Z(new_n720));
  NAND3_X1  g295(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n721));
  XNOR2_X1  g296(.A(new_n721), .B(KEYINPUT88), .ZN(new_n722));
  INV_X1    g297(.A(KEYINPUT26), .ZN(new_n723));
  XNOR2_X1  g298(.A(new_n722), .B(new_n723), .ZN(new_n724));
  NAND2_X1  g299(.A1(new_n477), .A2(G141), .ZN(new_n725));
  NAND2_X1  g300(.A1(new_n474), .A2(G129), .ZN(new_n726));
  NAND3_X1  g301(.A1(new_n468), .A2(G105), .A3(G2104), .ZN(new_n727));
  NAND3_X1  g302(.A1(new_n725), .A2(new_n726), .A3(new_n727), .ZN(new_n728));
  OR3_X1    g303(.A1(new_n724), .A2(KEYINPUT89), .A3(new_n728), .ZN(new_n729));
  OAI21_X1  g304(.A(KEYINPUT89), .B1(new_n724), .B2(new_n728), .ZN(new_n730));
  AND2_X1   g305(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  INV_X1    g306(.A(G29), .ZN(new_n732));
  NOR2_X1   g307(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  AOI21_X1  g308(.A(new_n733), .B1(new_n732), .B2(G32), .ZN(new_n734));
  XNOR2_X1  g309(.A(KEYINPUT27), .B(G1996), .ZN(new_n735));
  NAND2_X1  g310(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  XNOR2_X1  g311(.A(new_n736), .B(KEYINPUT90), .ZN(new_n737));
  NAND2_X1  g312(.A1(new_n687), .A2(G4), .ZN(new_n738));
  OAI21_X1  g313(.A(new_n738), .B1(new_n605), .B2(new_n687), .ZN(new_n739));
  OR2_X1    g314(.A1(new_n739), .A2(G1348), .ZN(new_n740));
  NAND2_X1  g315(.A1(new_n739), .A2(G1348), .ZN(new_n741));
  NAND3_X1  g316(.A1(new_n737), .A2(new_n740), .A3(new_n741), .ZN(new_n742));
  NAND2_X1  g317(.A1(G168), .A2(G16), .ZN(new_n743));
  XOR2_X1   g318(.A(new_n743), .B(KEYINPUT91), .Z(new_n744));
  OAI21_X1  g319(.A(new_n744), .B1(G16), .B2(G21), .ZN(new_n745));
  XNOR2_X1  g320(.A(new_n745), .B(G1966), .ZN(new_n746));
  INV_X1    g321(.A(G2090), .ZN(new_n747));
  NOR2_X1   g322(.A1(new_n709), .A2(G35), .ZN(new_n748));
  AOI21_X1  g323(.A(new_n748), .B1(G162), .B2(new_n709), .ZN(new_n749));
  XOR2_X1   g324(.A(new_n749), .B(KEYINPUT29), .Z(new_n750));
  OAI221_X1 g325(.A(new_n746), .B1(new_n747), .B2(new_n750), .C1(new_n734), .C2(new_n735), .ZN(new_n751));
  NOR2_X1   g326(.A1(G171), .A2(new_n687), .ZN(new_n752));
  AOI21_X1  g327(.A(new_n752), .B1(G5), .B2(new_n687), .ZN(new_n753));
  INV_X1    g328(.A(G1961), .ZN(new_n754));
  NOR2_X1   g329(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  XOR2_X1   g330(.A(new_n755), .B(KEYINPUT94), .Z(new_n756));
  NAND2_X1  g331(.A1(new_n687), .A2(G20), .ZN(new_n757));
  XOR2_X1   g332(.A(new_n757), .B(KEYINPUT23), .Z(new_n758));
  AOI21_X1  g333(.A(new_n758), .B1(G299), .B2(G16), .ZN(new_n759));
  XNOR2_X1  g334(.A(new_n759), .B(G1956), .ZN(new_n760));
  NOR2_X1   g335(.A1(new_n709), .A2(G27), .ZN(new_n761));
  AOI21_X1  g336(.A(new_n761), .B1(G164), .B2(new_n709), .ZN(new_n762));
  XOR2_X1   g337(.A(new_n762), .B(G2078), .Z(new_n763));
  XNOR2_X1  g338(.A(KEYINPUT24), .B(G34), .ZN(new_n764));
  NAND2_X1  g339(.A1(new_n708), .A2(new_n764), .ZN(new_n765));
  XOR2_X1   g340(.A(new_n765), .B(KEYINPUT86), .Z(new_n766));
  INV_X1    g341(.A(G160), .ZN(new_n767));
  OAI21_X1  g342(.A(new_n766), .B1(new_n767), .B2(new_n732), .ZN(new_n768));
  INV_X1    g343(.A(new_n768), .ZN(new_n769));
  NAND2_X1  g344(.A1(new_n769), .A2(G2084), .ZN(new_n770));
  XOR2_X1   g345(.A(new_n770), .B(KEYINPUT87), .Z(new_n771));
  NAND2_X1  g346(.A1(new_n732), .A2(G33), .ZN(new_n772));
  NAND3_X1  g347(.A1(new_n468), .A2(G103), .A3(G2104), .ZN(new_n773));
  XOR2_X1   g348(.A(new_n773), .B(KEYINPUT25), .Z(new_n774));
  NAND2_X1  g349(.A1(new_n477), .A2(G139), .ZN(new_n775));
  NAND2_X1  g350(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  NAND2_X1  g351(.A1(new_n498), .A2(G127), .ZN(new_n777));
  NAND2_X1  g352(.A1(G115), .A2(G2104), .ZN(new_n778));
  AOI21_X1  g353(.A(new_n468), .B1(new_n777), .B2(new_n778), .ZN(new_n779));
  NOR2_X1   g354(.A1(new_n776), .A2(new_n779), .ZN(new_n780));
  OAI21_X1  g355(.A(new_n772), .B1(new_n780), .B2(new_n732), .ZN(new_n781));
  OAI22_X1  g356(.A1(new_n769), .A2(G2084), .B1(new_n781), .B2(G2072), .ZN(new_n782));
  AOI21_X1  g357(.A(new_n782), .B1(G2072), .B2(new_n781), .ZN(new_n783));
  NAND2_X1  g358(.A1(new_n687), .A2(G19), .ZN(new_n784));
  OAI21_X1  g359(.A(new_n784), .B1(new_n548), .B2(new_n687), .ZN(new_n785));
  INV_X1    g360(.A(G1341), .ZN(new_n786));
  XNOR2_X1  g361(.A(new_n785), .B(new_n786), .ZN(new_n787));
  AND4_X1   g362(.A1(new_n763), .A2(new_n771), .A3(new_n783), .A4(new_n787), .ZN(new_n788));
  NAND2_X1  g363(.A1(new_n708), .A2(G26), .ZN(new_n789));
  XNOR2_X1  g364(.A(new_n789), .B(KEYINPUT28), .ZN(new_n790));
  NAND2_X1  g365(.A1(new_n477), .A2(G140), .ZN(new_n791));
  NAND2_X1  g366(.A1(new_n474), .A2(G128), .ZN(new_n792));
  OR2_X1    g367(.A1(G104), .A2(G2105), .ZN(new_n793));
  OAI211_X1 g368(.A(new_n793), .B(G2104), .C1(G116), .C2(new_n468), .ZN(new_n794));
  NAND3_X1  g369(.A1(new_n791), .A2(new_n792), .A3(new_n794), .ZN(new_n795));
  INV_X1    g370(.A(new_n795), .ZN(new_n796));
  OAI21_X1  g371(.A(new_n790), .B1(new_n796), .B2(new_n732), .ZN(new_n797));
  INV_X1    g372(.A(G2067), .ZN(new_n798));
  XNOR2_X1  g373(.A(new_n797), .B(new_n798), .ZN(new_n799));
  XOR2_X1   g374(.A(KEYINPUT93), .B(G28), .Z(new_n800));
  AOI21_X1  g375(.A(G29), .B1(new_n800), .B2(KEYINPUT30), .ZN(new_n801));
  OAI21_X1  g376(.A(new_n801), .B1(KEYINPUT30), .B2(new_n800), .ZN(new_n802));
  XNOR2_X1  g377(.A(KEYINPUT31), .B(G11), .ZN(new_n803));
  NAND2_X1  g378(.A1(new_n802), .A2(new_n803), .ZN(new_n804));
  OR2_X1    g379(.A1(new_n631), .A2(new_n708), .ZN(new_n805));
  INV_X1    g380(.A(KEYINPUT92), .ZN(new_n806));
  AOI21_X1  g381(.A(new_n804), .B1(new_n805), .B2(new_n806), .ZN(new_n807));
  OAI211_X1 g382(.A(new_n799), .B(new_n807), .C1(new_n806), .C2(new_n805), .ZN(new_n808));
  AOI21_X1  g383(.A(new_n808), .B1(new_n754), .B2(new_n753), .ZN(new_n809));
  NAND4_X1  g384(.A1(new_n756), .A2(new_n760), .A3(new_n788), .A4(new_n809), .ZN(new_n810));
  NAND2_X1  g385(.A1(new_n750), .A2(new_n747), .ZN(new_n811));
  XNOR2_X1  g386(.A(new_n811), .B(KEYINPUT95), .ZN(new_n812));
  OR4_X1    g387(.A1(new_n742), .A2(new_n751), .A3(new_n810), .A4(new_n812), .ZN(new_n813));
  NOR2_X1   g388(.A1(new_n720), .A2(new_n813), .ZN(G311));
  OR2_X1    g389(.A1(new_n720), .A2(new_n813), .ZN(G150));
  NAND2_X1  g390(.A1(new_n525), .A2(G55), .ZN(new_n816));
  INV_X1    g391(.A(G93), .ZN(new_n817));
  OAI21_X1  g392(.A(new_n816), .B1(new_n530), .B2(new_n817), .ZN(new_n818));
  INV_X1    g393(.A(KEYINPUT96), .ZN(new_n819));
  XNOR2_X1  g394(.A(new_n818), .B(new_n819), .ZN(new_n820));
  AOI22_X1  g395(.A1(new_n502), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n821));
  OR2_X1    g396(.A1(new_n821), .A2(new_n503), .ZN(new_n822));
  NAND2_X1  g397(.A1(new_n820), .A2(new_n822), .ZN(new_n823));
  NAND2_X1  g398(.A1(new_n823), .A2(G860), .ZN(new_n824));
  XOR2_X1   g399(.A(new_n824), .B(KEYINPUT37), .Z(new_n825));
  NAND2_X1  g400(.A1(new_n823), .A2(new_n547), .ZN(new_n826));
  NAND3_X1  g401(.A1(new_n820), .A2(new_n548), .A3(new_n822), .ZN(new_n827));
  NAND2_X1  g402(.A1(new_n826), .A2(new_n827), .ZN(new_n828));
  XOR2_X1   g403(.A(new_n828), .B(KEYINPUT38), .Z(new_n829));
  INV_X1    g404(.A(new_n605), .ZN(new_n830));
  NOR2_X1   g405(.A1(new_n830), .A2(new_n612), .ZN(new_n831));
  NAND2_X1  g406(.A1(new_n829), .A2(new_n831), .ZN(new_n832));
  XNOR2_X1  g407(.A(new_n828), .B(KEYINPUT38), .ZN(new_n833));
  OAI21_X1  g408(.A(new_n833), .B1(new_n612), .B2(new_n830), .ZN(new_n834));
  NAND2_X1  g409(.A1(new_n832), .A2(new_n834), .ZN(new_n835));
  INV_X1    g410(.A(KEYINPUT39), .ZN(new_n836));
  AOI21_X1  g411(.A(G860), .B1(new_n835), .B2(new_n836), .ZN(new_n837));
  NAND3_X1  g412(.A1(new_n832), .A2(new_n834), .A3(KEYINPUT39), .ZN(new_n838));
  AND3_X1   g413(.A1(new_n837), .A2(KEYINPUT97), .A3(new_n838), .ZN(new_n839));
  AOI21_X1  g414(.A(KEYINPUT97), .B1(new_n837), .B2(new_n838), .ZN(new_n840));
  OAI21_X1  g415(.A(new_n825), .B1(new_n839), .B2(new_n840), .ZN(new_n841));
  INV_X1    g416(.A(KEYINPUT98), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  OAI211_X1 g418(.A(KEYINPUT98), .B(new_n825), .C1(new_n839), .C2(new_n840), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n843), .A2(new_n844), .ZN(G145));
  NAND2_X1  g420(.A1(new_n731), .A2(new_n796), .ZN(new_n846));
  NAND2_X1  g421(.A1(new_n729), .A2(new_n730), .ZN(new_n847));
  NAND2_X1  g422(.A1(new_n847), .A2(new_n795), .ZN(new_n848));
  NAND2_X1  g423(.A1(new_n846), .A2(new_n848), .ZN(new_n849));
  AOI21_X1  g424(.A(KEYINPUT4), .B1(new_n477), .B2(G138), .ZN(new_n850));
  NOR2_X1   g425(.A1(new_n495), .A2(new_n496), .ZN(new_n851));
  OAI21_X1  g426(.A(KEYINPUT99), .B1(new_n850), .B2(new_n851), .ZN(new_n852));
  AOI22_X1  g427(.A1(new_n487), .A2(new_n490), .B1(new_n474), .B2(G126), .ZN(new_n853));
  INV_X1    g428(.A(KEYINPUT99), .ZN(new_n854));
  NAND3_X1  g429(.A1(new_n497), .A2(new_n499), .A3(new_n854), .ZN(new_n855));
  NAND3_X1  g430(.A1(new_n852), .A2(new_n853), .A3(new_n855), .ZN(new_n856));
  NAND2_X1  g431(.A1(new_n856), .A2(KEYINPUT100), .ZN(new_n857));
  AOI21_X1  g432(.A(new_n854), .B1(new_n497), .B2(new_n499), .ZN(new_n858));
  AOI21_X1  g433(.A(KEYINPUT67), .B1(new_n484), .B2(new_n486), .ZN(new_n859));
  NOR3_X1   g434(.A1(new_n489), .A2(new_n488), .A3(new_n485), .ZN(new_n860));
  OAI21_X1  g435(.A(new_n492), .B1(new_n859), .B2(new_n860), .ZN(new_n861));
  NOR2_X1   g436(.A1(new_n858), .A2(new_n861), .ZN(new_n862));
  INV_X1    g437(.A(KEYINPUT100), .ZN(new_n863));
  NAND3_X1  g438(.A1(new_n862), .A2(new_n863), .A3(new_n855), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n857), .A2(new_n864), .ZN(new_n865));
  INV_X1    g440(.A(new_n865), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n849), .A2(new_n866), .ZN(new_n867));
  NAND3_X1  g442(.A1(new_n846), .A2(new_n865), .A3(new_n848), .ZN(new_n868));
  NAND2_X1  g443(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  INV_X1    g444(.A(new_n780), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n477), .A2(G142), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n474), .A2(G130), .ZN(new_n873));
  NOR2_X1   g448(.A1(G106), .A2(G2105), .ZN(new_n874));
  OAI21_X1  g449(.A(G2104), .B1(new_n468), .B2(G118), .ZN(new_n875));
  OAI211_X1 g450(.A(new_n872), .B(new_n873), .C1(new_n874), .C2(new_n875), .ZN(new_n876));
  XOR2_X1   g451(.A(new_n622), .B(new_n876), .Z(new_n877));
  XNOR2_X1  g452(.A(new_n877), .B(new_n707), .ZN(new_n878));
  NAND3_X1  g453(.A1(new_n867), .A2(new_n780), .A3(new_n868), .ZN(new_n879));
  NAND3_X1  g454(.A1(new_n871), .A2(new_n878), .A3(new_n879), .ZN(new_n880));
  XOR2_X1   g455(.A(G160), .B(new_n631), .Z(new_n881));
  XOR2_X1   g456(.A(new_n881), .B(G162), .Z(new_n882));
  INV_X1    g457(.A(new_n882), .ZN(new_n883));
  AND2_X1   g458(.A1(new_n880), .A2(new_n883), .ZN(new_n884));
  INV_X1    g459(.A(new_n878), .ZN(new_n885));
  INV_X1    g460(.A(new_n879), .ZN(new_n886));
  AOI21_X1  g461(.A(new_n780), .B1(new_n867), .B2(new_n868), .ZN(new_n887));
  OAI21_X1  g462(.A(new_n885), .B1(new_n886), .B2(new_n887), .ZN(new_n888));
  INV_X1    g463(.A(KEYINPUT102), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  OAI211_X1 g465(.A(KEYINPUT102), .B(new_n885), .C1(new_n886), .C2(new_n887), .ZN(new_n891));
  NAND3_X1  g466(.A1(new_n884), .A2(new_n890), .A3(new_n891), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n892), .A2(KEYINPUT103), .ZN(new_n893));
  INV_X1    g468(.A(KEYINPUT103), .ZN(new_n894));
  NAND4_X1  g469(.A1(new_n884), .A2(new_n890), .A3(new_n894), .A4(new_n891), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n893), .A2(new_n895), .ZN(new_n896));
  XOR2_X1   g471(.A(KEYINPUT101), .B(G37), .Z(new_n897));
  NAND2_X1  g472(.A1(new_n888), .A2(new_n880), .ZN(new_n898));
  AOI21_X1  g473(.A(new_n897), .B1(new_n898), .B2(new_n882), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n896), .A2(new_n899), .ZN(new_n900));
  XNOR2_X1  g475(.A(new_n900), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g476(.A1(new_n830), .A2(new_n567), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n605), .A2(G299), .ZN(new_n903));
  AND2_X1   g478(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  XOR2_X1   g479(.A(KEYINPUT104), .B(KEYINPUT41), .Z(new_n905));
  INV_X1    g480(.A(new_n905), .ZN(new_n906));
  NAND3_X1  g481(.A1(new_n904), .A2(KEYINPUT105), .A3(new_n906), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n902), .A2(new_n903), .ZN(new_n908));
  INV_X1    g483(.A(KEYINPUT41), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  INV_X1    g485(.A(KEYINPUT105), .ZN(new_n911));
  OAI21_X1  g486(.A(new_n911), .B1(new_n908), .B2(new_n905), .ZN(new_n912));
  NAND3_X1  g487(.A1(new_n907), .A2(new_n910), .A3(new_n912), .ZN(new_n913));
  XNOR2_X1  g488(.A(new_n828), .B(new_n616), .ZN(new_n914));
  INV_X1    g489(.A(new_n914), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n913), .A2(new_n915), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n914), .A2(new_n908), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  INV_X1    g493(.A(KEYINPUT106), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  XOR2_X1   g495(.A(G288), .B(G290), .Z(new_n921));
  XNOR2_X1  g496(.A(new_n589), .B(new_n519), .ZN(new_n922));
  XNOR2_X1  g497(.A(new_n921), .B(new_n922), .ZN(new_n923));
  XNOR2_X1  g498(.A(new_n923), .B(KEYINPUT42), .ZN(new_n924));
  AND2_X1   g499(.A1(new_n920), .A2(new_n924), .ZN(new_n925));
  NAND3_X1  g500(.A1(new_n916), .A2(KEYINPUT106), .A3(new_n917), .ZN(new_n926));
  AOI21_X1  g501(.A(new_n924), .B1(new_n920), .B2(new_n926), .ZN(new_n927));
  OAI21_X1  g502(.A(G868), .B1(new_n925), .B2(new_n927), .ZN(new_n928));
  INV_X1    g503(.A(new_n823), .ZN(new_n929));
  OAI21_X1  g504(.A(new_n928), .B1(G868), .B2(new_n929), .ZN(G295));
  OAI21_X1  g505(.A(new_n928), .B1(G868), .B2(new_n929), .ZN(G331));
  INV_X1    g506(.A(KEYINPUT43), .ZN(new_n932));
  INV_X1    g507(.A(KEYINPUT107), .ZN(new_n933));
  NAND2_X1  g508(.A1(G171), .A2(new_n933), .ZN(new_n934));
  NAND2_X1  g509(.A1(G301), .A2(KEYINPUT107), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n936), .A2(G286), .ZN(new_n937));
  NAND3_X1  g512(.A1(new_n934), .A2(G168), .A3(new_n935), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  OR2_X1    g514(.A1(new_n828), .A2(new_n939), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n828), .A2(new_n939), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n913), .A2(new_n942), .ZN(new_n943));
  INV_X1    g518(.A(KEYINPUT108), .ZN(new_n944));
  NAND3_X1  g519(.A1(new_n828), .A2(new_n939), .A3(new_n944), .ZN(new_n945));
  INV_X1    g520(.A(new_n945), .ZN(new_n946));
  AOI21_X1  g521(.A(new_n944), .B1(new_n828), .B2(new_n939), .ZN(new_n947));
  NOR2_X1   g522(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  NOR2_X1   g523(.A1(new_n828), .A2(new_n939), .ZN(new_n949));
  NOR2_X1   g524(.A1(new_n949), .A2(new_n904), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n948), .A2(new_n950), .ZN(new_n951));
  NAND3_X1  g526(.A1(new_n943), .A2(new_n951), .A3(new_n923), .ZN(new_n952));
  INV_X1    g527(.A(G37), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n952), .A2(new_n953), .ZN(new_n954));
  AOI22_X1  g529(.A1(new_n913), .A2(new_n942), .B1(new_n948), .B2(new_n950), .ZN(new_n955));
  NOR2_X1   g530(.A1(new_n955), .A2(new_n923), .ZN(new_n956));
  OAI21_X1  g531(.A(new_n932), .B1(new_n954), .B2(new_n956), .ZN(new_n957));
  AOI21_X1  g532(.A(new_n897), .B1(new_n955), .B2(new_n923), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n941), .A2(KEYINPUT108), .ZN(new_n959));
  NAND3_X1  g534(.A1(new_n959), .A2(new_n940), .A3(new_n945), .ZN(new_n960));
  AOI21_X1  g535(.A(new_n905), .B1(new_n902), .B2(new_n903), .ZN(new_n961));
  AOI21_X1  g536(.A(new_n961), .B1(new_n909), .B2(new_n904), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n960), .A2(new_n962), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n950), .A2(new_n941), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n963), .A2(new_n964), .ZN(new_n965));
  INV_X1    g540(.A(new_n923), .ZN(new_n966));
  AOI21_X1  g541(.A(KEYINPUT109), .B1(new_n965), .B2(new_n966), .ZN(new_n967));
  INV_X1    g542(.A(KEYINPUT109), .ZN(new_n968));
  AOI211_X1 g543(.A(new_n968), .B(new_n923), .C1(new_n963), .C2(new_n964), .ZN(new_n969));
  OAI21_X1  g544(.A(new_n958), .B1(new_n967), .B2(new_n969), .ZN(new_n970));
  OAI21_X1  g545(.A(new_n957), .B1(new_n970), .B2(new_n932), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n971), .A2(KEYINPUT44), .ZN(new_n972));
  OAI211_X1 g547(.A(new_n958), .B(new_n932), .C1(new_n967), .C2(new_n969), .ZN(new_n973));
  OAI21_X1  g548(.A(KEYINPUT43), .B1(new_n954), .B2(new_n956), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n973), .A2(new_n974), .ZN(new_n975));
  INV_X1    g550(.A(KEYINPUT44), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n975), .A2(new_n976), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n972), .A2(new_n977), .ZN(G397));
  INV_X1    g553(.A(G1384), .ZN(new_n979));
  NAND3_X1  g554(.A1(new_n857), .A2(new_n979), .A3(new_n864), .ZN(new_n980));
  INV_X1    g555(.A(KEYINPUT45), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n980), .A2(new_n981), .ZN(new_n982));
  INV_X1    g557(.A(new_n982), .ZN(new_n983));
  NAND3_X1  g558(.A1(new_n467), .A2(new_n472), .A3(G40), .ZN(new_n984));
  INV_X1    g559(.A(KEYINPUT110), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n984), .A2(new_n985), .ZN(new_n986));
  NAND4_X1  g561(.A1(new_n467), .A2(new_n472), .A3(KEYINPUT110), .A4(G40), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n986), .A2(new_n987), .ZN(new_n988));
  NAND2_X1  g563(.A1(new_n983), .A2(new_n988), .ZN(new_n989));
  NOR2_X1   g564(.A1(new_n989), .A2(G1996), .ZN(new_n990));
  OR2_X1    g565(.A1(new_n990), .A2(KEYINPUT46), .ZN(new_n991));
  INV_X1    g566(.A(new_n989), .ZN(new_n992));
  XNOR2_X1  g567(.A(new_n795), .B(G2067), .ZN(new_n993));
  OAI21_X1  g568(.A(new_n992), .B1(new_n847), .B2(new_n993), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n991), .A2(new_n994), .ZN(new_n995));
  AOI21_X1  g570(.A(new_n995), .B1(KEYINPUT46), .B2(new_n990), .ZN(new_n996));
  AND2_X1   g571(.A1(new_n996), .A2(KEYINPUT47), .ZN(new_n997));
  NOR2_X1   g572(.A1(new_n996), .A2(KEYINPUT47), .ZN(new_n998));
  INV_X1    g573(.A(KEYINPUT48), .ZN(new_n999));
  OR3_X1    g574(.A1(new_n989), .A2(G1986), .A3(G290), .ZN(new_n1000));
  OR2_X1    g575(.A1(new_n731), .A2(G1996), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n731), .A2(G1996), .ZN(new_n1002));
  AOI21_X1  g577(.A(new_n993), .B1(new_n1001), .B2(new_n1002), .ZN(new_n1003));
  XOR2_X1   g578(.A(new_n707), .B(new_n711), .Z(new_n1004));
  NAND2_X1  g579(.A1(new_n1003), .A2(new_n1004), .ZN(new_n1005));
  AOI22_X1  g580(.A1(new_n999), .A2(new_n1000), .B1(new_n1005), .B2(new_n992), .ZN(new_n1006));
  OAI21_X1  g581(.A(new_n1006), .B1(new_n999), .B2(new_n1000), .ZN(new_n1007));
  NOR2_X1   g582(.A1(new_n707), .A2(new_n711), .ZN(new_n1008));
  AOI22_X1  g583(.A1(new_n1003), .A2(new_n1008), .B1(new_n798), .B2(new_n796), .ZN(new_n1009));
  OAI21_X1  g584(.A(new_n1007), .B1(new_n989), .B2(new_n1009), .ZN(new_n1010));
  NOR3_X1   g585(.A1(new_n997), .A2(new_n998), .A3(new_n1010), .ZN(new_n1011));
  INV_X1    g586(.A(KEYINPUT53), .ZN(new_n1012));
  NOR2_X1   g587(.A1(new_n981), .A2(G1384), .ZN(new_n1013));
  NAND3_X1  g588(.A1(new_n857), .A2(new_n864), .A3(new_n1013), .ZN(new_n1014));
  INV_X1    g589(.A(KEYINPUT111), .ZN(new_n1015));
  NOR2_X1   g590(.A1(new_n850), .A2(new_n851), .ZN(new_n1016));
  AOI21_X1  g591(.A(G1384), .B1(new_n1016), .B2(new_n853), .ZN(new_n1017));
  OAI21_X1  g592(.A(new_n1015), .B1(new_n1017), .B2(KEYINPUT45), .ZN(new_n1018));
  AOI21_X1  g593(.A(KEYINPUT45), .B1(new_n500), .B2(new_n979), .ZN(new_n1019));
  AOI22_X1  g594(.A1(new_n1019), .A2(KEYINPUT111), .B1(new_n986), .B2(new_n987), .ZN(new_n1020));
  NAND3_X1  g595(.A1(new_n1014), .A2(new_n1018), .A3(new_n1020), .ZN(new_n1021));
  OAI21_X1  g596(.A(new_n1012), .B1(new_n1021), .B2(G2078), .ZN(new_n1022));
  INV_X1    g597(.A(new_n984), .ZN(new_n1023));
  NOR2_X1   g598(.A1(new_n1012), .A2(G2078), .ZN(new_n1024));
  NAND4_X1  g599(.A1(new_n982), .A2(new_n1023), .A3(new_n1014), .A4(new_n1024), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n497), .A2(new_n499), .ZN(new_n1026));
  OAI21_X1  g601(.A(new_n979), .B1(new_n861), .B2(new_n1026), .ZN(new_n1027));
  AOI22_X1  g602(.A1(new_n987), .A2(new_n986), .B1(new_n1027), .B2(KEYINPUT50), .ZN(new_n1028));
  INV_X1    g603(.A(KEYINPUT50), .ZN(new_n1029));
  NAND3_X1  g604(.A1(new_n856), .A2(new_n1029), .A3(new_n979), .ZN(new_n1030));
  NAND2_X1  g605(.A1(new_n1028), .A2(new_n1030), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n1031), .A2(new_n754), .ZN(new_n1032));
  NAND3_X1  g607(.A1(new_n1022), .A2(new_n1025), .A3(new_n1032), .ZN(new_n1033));
  OR3_X1    g608(.A1(new_n1033), .A2(KEYINPUT124), .A3(G171), .ZN(new_n1034));
  OAI21_X1  g609(.A(KEYINPUT124), .B1(new_n1033), .B2(G171), .ZN(new_n1035));
  AOI21_X1  g610(.A(G1384), .B1(new_n862), .B2(new_n855), .ZN(new_n1036));
  NOR2_X1   g611(.A1(new_n1036), .A2(KEYINPUT45), .ZN(new_n1037));
  OAI21_X1  g612(.A(new_n988), .B1(new_n981), .B2(new_n1027), .ZN(new_n1038));
  NOR2_X1   g613(.A1(new_n1037), .A2(new_n1038), .ZN(new_n1039));
  AOI22_X1  g614(.A1(new_n1039), .A2(new_n1024), .B1(new_n754), .B2(new_n1031), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n1040), .A2(new_n1022), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n1041), .A2(G171), .ZN(new_n1042));
  NAND3_X1  g617(.A1(new_n1034), .A2(new_n1035), .A3(new_n1042), .ZN(new_n1043));
  INV_X1    g618(.A(KEYINPUT54), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n1043), .A2(new_n1044), .ZN(new_n1045));
  INV_X1    g620(.A(KEYINPUT51), .ZN(new_n1046));
  INV_X1    g621(.A(G1966), .ZN(new_n1047));
  OAI21_X1  g622(.A(new_n1047), .B1(new_n1037), .B2(new_n1038), .ZN(new_n1048));
  XOR2_X1   g623(.A(KEYINPUT114), .B(G2084), .Z(new_n1049));
  NAND3_X1  g624(.A1(new_n1028), .A2(new_n1030), .A3(new_n1049), .ZN(new_n1050));
  NAND2_X1  g625(.A1(new_n1048), .A2(new_n1050), .ZN(new_n1051));
  OAI211_X1 g626(.A(new_n1046), .B(G8), .C1(new_n1051), .C2(G286), .ZN(new_n1052));
  INV_X1    g627(.A(new_n1050), .ZN(new_n1053));
  AND3_X1   g628(.A1(new_n497), .A2(new_n499), .A3(new_n854), .ZN(new_n1054));
  NOR3_X1   g629(.A1(new_n1054), .A2(new_n858), .A3(new_n861), .ZN(new_n1055));
  OAI21_X1  g630(.A(new_n981), .B1(new_n1055), .B2(G1384), .ZN(new_n1056));
  AOI22_X1  g631(.A1(new_n1017), .A2(KEYINPUT45), .B1(new_n986), .B2(new_n987), .ZN(new_n1057));
  AOI21_X1  g632(.A(G1966), .B1(new_n1056), .B2(new_n1057), .ZN(new_n1058));
  OAI21_X1  g633(.A(G8), .B1(new_n1053), .B2(new_n1058), .ZN(new_n1059));
  INV_X1    g634(.A(G8), .ZN(new_n1060));
  NOR2_X1   g635(.A1(G168), .A2(new_n1060), .ZN(new_n1061));
  INV_X1    g636(.A(new_n1061), .ZN(new_n1062));
  NAND3_X1  g637(.A1(new_n1059), .A2(KEYINPUT51), .A3(new_n1062), .ZN(new_n1063));
  INV_X1    g638(.A(KEYINPUT123), .ZN(new_n1064));
  AOI21_X1  g639(.A(new_n1064), .B1(new_n1051), .B2(new_n1061), .ZN(new_n1065));
  AOI211_X1 g640(.A(KEYINPUT123), .B(new_n1062), .C1(new_n1048), .C2(new_n1050), .ZN(new_n1066));
  OAI211_X1 g641(.A(new_n1052), .B(new_n1063), .C1(new_n1065), .C2(new_n1066), .ZN(new_n1067));
  INV_X1    g642(.A(KEYINPUT49), .ZN(new_n1068));
  NOR3_X1   g643(.A1(new_n582), .A2(G1981), .A3(new_n588), .ZN(new_n1069));
  INV_X1    g644(.A(G1981), .ZN(new_n1070));
  AND2_X1   g645(.A1(new_n586), .A2(new_n587), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n512), .A2(G86), .ZN(new_n1072));
  AOI21_X1  g647(.A(new_n1070), .B1(new_n1071), .B2(new_n1072), .ZN(new_n1073));
  OAI21_X1  g648(.A(new_n1068), .B1(new_n1069), .B2(new_n1073), .ZN(new_n1074));
  AOI21_X1  g649(.A(new_n1060), .B1(new_n1036), .B2(new_n988), .ZN(new_n1075));
  OAI211_X1 g650(.A(new_n1070), .B(new_n1071), .C1(new_n601), .C2(new_n581), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n1071), .A2(new_n1072), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n1077), .A2(G1981), .ZN(new_n1078));
  NAND3_X1  g653(.A1(new_n1076), .A2(new_n1078), .A3(KEYINPUT49), .ZN(new_n1079));
  NAND3_X1  g654(.A1(new_n1074), .A2(new_n1075), .A3(new_n1079), .ZN(new_n1080));
  INV_X1    g655(.A(G1976), .ZN(new_n1081));
  AOI21_X1  g656(.A(KEYINPUT52), .B1(G288), .B2(new_n1081), .ZN(new_n1082));
  OAI211_X1 g657(.A(new_n1082), .B(new_n1075), .C1(new_n1081), .C2(G288), .ZN(new_n1083));
  OAI21_X1  g658(.A(new_n1075), .B1(new_n1081), .B2(G288), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n1084), .A2(KEYINPUT52), .ZN(new_n1085));
  NAND3_X1  g660(.A1(new_n1080), .A2(new_n1083), .A3(new_n1085), .ZN(new_n1086));
  NAND3_X1  g661(.A1(new_n500), .A2(new_n1029), .A3(new_n979), .ZN(new_n1087));
  NAND2_X1  g662(.A1(new_n988), .A2(new_n1087), .ZN(new_n1088));
  AOI21_X1  g663(.A(new_n1029), .B1(new_n856), .B2(new_n979), .ZN(new_n1089));
  OAI21_X1  g664(.A(KEYINPUT113), .B1(new_n1088), .B2(new_n1089), .ZN(new_n1090));
  OAI21_X1  g665(.A(KEYINPUT50), .B1(new_n1055), .B2(G1384), .ZN(new_n1091));
  AOI22_X1  g666(.A1(new_n1017), .A2(new_n1029), .B1(new_n986), .B2(new_n987), .ZN(new_n1092));
  INV_X1    g667(.A(KEYINPUT113), .ZN(new_n1093));
  NAND3_X1  g668(.A1(new_n1091), .A2(new_n1092), .A3(new_n1093), .ZN(new_n1094));
  NAND3_X1  g669(.A1(new_n1090), .A2(new_n1094), .A3(new_n747), .ZN(new_n1095));
  INV_X1    g670(.A(G1971), .ZN(new_n1096));
  AND3_X1   g671(.A1(new_n857), .A2(new_n864), .A3(new_n1013), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n1019), .A2(KEYINPUT111), .ZN(new_n1098));
  NAND3_X1  g673(.A1(new_n1018), .A2(new_n988), .A3(new_n1098), .ZN(new_n1099));
  OAI21_X1  g674(.A(new_n1096), .B1(new_n1097), .B2(new_n1099), .ZN(new_n1100));
  NAND2_X1  g675(.A1(new_n1095), .A2(new_n1100), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n1101), .A2(G8), .ZN(new_n1102));
  NAND3_X1  g677(.A1(new_n572), .A2(G8), .A3(new_n573), .ZN(new_n1103));
  XNOR2_X1  g678(.A(new_n1103), .B(KEYINPUT55), .ZN(new_n1104));
  AOI21_X1  g679(.A(new_n1086), .B1(new_n1102), .B2(new_n1104), .ZN(new_n1105));
  INV_X1    g680(.A(KEYINPUT55), .ZN(new_n1106));
  XNOR2_X1  g681(.A(new_n1103), .B(new_n1106), .ZN(new_n1107));
  INV_X1    g682(.A(KEYINPUT112), .ZN(new_n1108));
  OAI22_X1  g683(.A1(new_n1100), .A2(new_n1108), .B1(G2090), .B2(new_n1031), .ZN(new_n1109));
  AOI21_X1  g684(.A(KEYINPUT112), .B1(new_n1021), .B2(new_n1096), .ZN(new_n1110));
  OAI211_X1 g685(.A(new_n1107), .B(G8), .C1(new_n1109), .C2(new_n1110), .ZN(new_n1111));
  NAND3_X1  g686(.A1(new_n1067), .A2(new_n1105), .A3(new_n1111), .ZN(new_n1112));
  NAND3_X1  g687(.A1(new_n1040), .A2(new_n1022), .A3(G301), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n1113), .A2(KEYINPUT54), .ZN(new_n1114));
  INV_X1    g689(.A(KEYINPUT125), .ZN(new_n1115));
  AOI21_X1  g690(.A(G301), .B1(new_n1033), .B2(new_n1115), .ZN(new_n1116));
  NAND4_X1  g691(.A1(new_n1022), .A2(new_n1025), .A3(KEYINPUT125), .A4(new_n1032), .ZN(new_n1117));
  AOI21_X1  g692(.A(new_n1114), .B1(new_n1116), .B2(new_n1117), .ZN(new_n1118));
  NOR2_X1   g693(.A1(new_n1112), .A2(new_n1118), .ZN(new_n1119));
  AOI21_X1  g694(.A(G1956), .B1(new_n1091), .B2(new_n1092), .ZN(new_n1120));
  XNOR2_X1  g695(.A(KEYINPUT56), .B(G2072), .ZN(new_n1121));
  NAND4_X1  g696(.A1(new_n1014), .A2(new_n1018), .A3(new_n1020), .A4(new_n1121), .ZN(new_n1122));
  AOI21_X1  g697(.A(new_n1120), .B1(new_n1122), .B2(KEYINPUT116), .ZN(new_n1123));
  AND2_X1   g698(.A1(new_n1020), .A2(new_n1018), .ZN(new_n1124));
  INV_X1    g699(.A(KEYINPUT116), .ZN(new_n1125));
  NAND4_X1  g700(.A1(new_n1124), .A2(new_n1125), .A3(new_n1014), .A4(new_n1121), .ZN(new_n1126));
  NAND2_X1  g701(.A1(new_n1123), .A2(new_n1126), .ZN(new_n1127));
  INV_X1    g702(.A(KEYINPUT57), .ZN(new_n1128));
  INV_X1    g703(.A(new_n566), .ZN(new_n1129));
  AOI21_X1  g704(.A(new_n1128), .B1(new_n1129), .B2(new_n560), .ZN(new_n1130));
  NOR3_X1   g705(.A1(new_n561), .A2(new_n566), .A3(KEYINPUT57), .ZN(new_n1131));
  OAI21_X1  g706(.A(KEYINPUT117), .B1(new_n1130), .B2(new_n1131), .ZN(new_n1132));
  OAI21_X1  g707(.A(KEYINPUT57), .B1(new_n561), .B2(new_n566), .ZN(new_n1133));
  NAND3_X1  g708(.A1(new_n1129), .A2(new_n1128), .A3(new_n560), .ZN(new_n1134));
  INV_X1    g709(.A(KEYINPUT117), .ZN(new_n1135));
  NAND3_X1  g710(.A1(new_n1133), .A2(new_n1134), .A3(new_n1135), .ZN(new_n1136));
  AND2_X1   g711(.A1(new_n1132), .A2(new_n1136), .ZN(new_n1137));
  NAND2_X1  g712(.A1(new_n1127), .A2(new_n1137), .ZN(new_n1138));
  NOR2_X1   g713(.A1(new_n1130), .A2(new_n1131), .ZN(new_n1139));
  NAND3_X1  g714(.A1(new_n1123), .A2(new_n1126), .A3(new_n1139), .ZN(new_n1140));
  NAND3_X1  g715(.A1(new_n1138), .A2(KEYINPUT61), .A3(new_n1140), .ZN(new_n1141));
  INV_X1    g716(.A(KEYINPUT61), .ZN(new_n1142));
  NAND2_X1  g717(.A1(new_n1122), .A2(KEYINPUT116), .ZN(new_n1143));
  INV_X1    g718(.A(new_n1120), .ZN(new_n1144));
  AND4_X1   g719(.A1(new_n1126), .A2(new_n1143), .A3(new_n1144), .A4(new_n1139), .ZN(new_n1145));
  AOI21_X1  g720(.A(new_n1139), .B1(new_n1123), .B2(new_n1126), .ZN(new_n1146));
  OAI21_X1  g721(.A(new_n1142), .B1(new_n1145), .B2(new_n1146), .ZN(new_n1147));
  NAND2_X1  g722(.A1(new_n1036), .A2(new_n988), .ZN(new_n1148));
  XNOR2_X1  g723(.A(KEYINPUT119), .B(KEYINPUT58), .ZN(new_n1149));
  XNOR2_X1  g724(.A(new_n1149), .B(new_n786), .ZN(new_n1150));
  NAND2_X1  g725(.A1(new_n1148), .A2(new_n1150), .ZN(new_n1151));
  OAI21_X1  g726(.A(new_n1151), .B1(new_n1021), .B2(G1996), .ZN(new_n1152));
  INV_X1    g727(.A(KEYINPUT121), .ZN(new_n1153));
  AOI21_X1  g728(.A(new_n547), .B1(new_n1153), .B2(KEYINPUT59), .ZN(new_n1154));
  NAND2_X1  g729(.A1(new_n1152), .A2(new_n1154), .ZN(new_n1155));
  INV_X1    g730(.A(KEYINPUT120), .ZN(new_n1156));
  AOI21_X1  g731(.A(new_n1153), .B1(new_n1156), .B2(KEYINPUT59), .ZN(new_n1157));
  INV_X1    g732(.A(new_n1157), .ZN(new_n1158));
  NAND2_X1  g733(.A1(new_n1155), .A2(new_n1158), .ZN(new_n1159));
  NAND3_X1  g734(.A1(new_n1152), .A2(new_n1157), .A3(new_n1154), .ZN(new_n1160));
  NAND2_X1  g735(.A1(new_n1159), .A2(new_n1160), .ZN(new_n1161));
  INV_X1    g736(.A(G1348), .ZN(new_n1162));
  AND3_X1   g737(.A1(new_n856), .A2(new_n1029), .A3(new_n979), .ZN(new_n1163));
  NAND2_X1  g738(.A1(new_n1027), .A2(KEYINPUT50), .ZN(new_n1164));
  NAND2_X1  g739(.A1(new_n988), .A2(new_n1164), .ZN(new_n1165));
  OAI21_X1  g740(.A(new_n1162), .B1(new_n1163), .B2(new_n1165), .ZN(new_n1166));
  NAND3_X1  g741(.A1(new_n1036), .A2(new_n798), .A3(new_n988), .ZN(new_n1167));
  NAND2_X1  g742(.A1(new_n1166), .A2(new_n1167), .ZN(new_n1168));
  INV_X1    g743(.A(KEYINPUT60), .ZN(new_n1169));
  AOI21_X1  g744(.A(new_n830), .B1(new_n1168), .B2(new_n1169), .ZN(new_n1170));
  AOI21_X1  g745(.A(G1348), .B1(new_n1028), .B2(new_n1030), .ZN(new_n1171));
  AND3_X1   g746(.A1(new_n1036), .A2(new_n798), .A3(new_n988), .ZN(new_n1172));
  NOR2_X1   g747(.A1(new_n1171), .A2(new_n1172), .ZN(new_n1173));
  AOI21_X1  g748(.A(KEYINPUT122), .B1(new_n1173), .B2(KEYINPUT60), .ZN(new_n1174));
  INV_X1    g749(.A(KEYINPUT122), .ZN(new_n1175));
  NOR4_X1   g750(.A1(new_n1171), .A2(new_n1172), .A3(new_n1175), .A4(new_n1169), .ZN(new_n1176));
  OAI21_X1  g751(.A(new_n1170), .B1(new_n1174), .B2(new_n1176), .ZN(new_n1177));
  OAI21_X1  g752(.A(new_n1175), .B1(new_n1168), .B2(new_n1169), .ZN(new_n1178));
  OAI21_X1  g753(.A(new_n1169), .B1(new_n1171), .B2(new_n1172), .ZN(new_n1179));
  NAND2_X1  g754(.A1(new_n1179), .A2(new_n605), .ZN(new_n1180));
  NAND3_X1  g755(.A1(new_n1173), .A2(KEYINPUT122), .A3(KEYINPUT60), .ZN(new_n1181));
  NAND3_X1  g756(.A1(new_n1178), .A2(new_n1180), .A3(new_n1181), .ZN(new_n1182));
  NAND2_X1  g757(.A1(new_n1177), .A2(new_n1182), .ZN(new_n1183));
  AND4_X1   g758(.A1(new_n1141), .A2(new_n1147), .A3(new_n1161), .A4(new_n1183), .ZN(new_n1184));
  NOR2_X1   g759(.A1(new_n1173), .A2(new_n830), .ZN(new_n1185));
  AOI21_X1  g760(.A(new_n1185), .B1(new_n1127), .B2(new_n1137), .ZN(new_n1186));
  OAI21_X1  g761(.A(KEYINPUT118), .B1(new_n1186), .B2(new_n1145), .ZN(new_n1187));
  INV_X1    g762(.A(KEYINPUT118), .ZN(new_n1188));
  NAND2_X1  g763(.A1(new_n1132), .A2(new_n1136), .ZN(new_n1189));
  AOI21_X1  g764(.A(new_n1189), .B1(new_n1123), .B2(new_n1126), .ZN(new_n1190));
  OAI211_X1 g765(.A(new_n1188), .B(new_n1140), .C1(new_n1190), .C2(new_n1185), .ZN(new_n1191));
  NAND2_X1  g766(.A1(new_n1187), .A2(new_n1191), .ZN(new_n1192));
  OAI211_X1 g767(.A(new_n1045), .B(new_n1119), .C1(new_n1184), .C2(new_n1192), .ZN(new_n1193));
  AND3_X1   g768(.A1(new_n1080), .A2(new_n1081), .A3(new_n692), .ZN(new_n1194));
  OAI21_X1  g769(.A(new_n1075), .B1(new_n1194), .B2(new_n1069), .ZN(new_n1195));
  OAI21_X1  g770(.A(new_n1195), .B1(new_n1111), .B2(new_n1086), .ZN(new_n1196));
  INV_X1    g771(.A(KEYINPUT115), .ZN(new_n1197));
  OAI21_X1  g772(.A(new_n1197), .B1(new_n1059), .B2(G286), .ZN(new_n1198));
  NAND4_X1  g773(.A1(new_n1051), .A2(KEYINPUT115), .A3(G8), .A4(G168), .ZN(new_n1199));
  NAND2_X1  g774(.A1(new_n1198), .A2(new_n1199), .ZN(new_n1200));
  NAND3_X1  g775(.A1(new_n1105), .A2(new_n1111), .A3(new_n1200), .ZN(new_n1201));
  INV_X1    g776(.A(KEYINPUT63), .ZN(new_n1202));
  NAND2_X1  g777(.A1(new_n1201), .A2(new_n1202), .ZN(new_n1203));
  OAI21_X1  g778(.A(G8), .B1(new_n1109), .B2(new_n1110), .ZN(new_n1204));
  NAND2_X1  g779(.A1(new_n1204), .A2(new_n1104), .ZN(new_n1205));
  NOR2_X1   g780(.A1(new_n1086), .A2(new_n1202), .ZN(new_n1206));
  NAND4_X1  g781(.A1(new_n1205), .A2(new_n1111), .A3(new_n1200), .A4(new_n1206), .ZN(new_n1207));
  AOI21_X1  g782(.A(new_n1196), .B1(new_n1203), .B2(new_n1207), .ZN(new_n1208));
  AND3_X1   g783(.A1(new_n1193), .A2(KEYINPUT126), .A3(new_n1208), .ZN(new_n1209));
  AOI21_X1  g784(.A(KEYINPUT126), .B1(new_n1193), .B2(new_n1208), .ZN(new_n1210));
  NAND2_X1  g785(.A1(new_n1105), .A2(new_n1111), .ZN(new_n1211));
  OAI211_X1 g786(.A(G171), .B(new_n1041), .C1(new_n1067), .C2(KEYINPUT62), .ZN(new_n1212));
  AOI211_X1 g787(.A(new_n1211), .B(new_n1212), .C1(KEYINPUT62), .C2(new_n1067), .ZN(new_n1213));
  NOR3_X1   g788(.A1(new_n1209), .A2(new_n1210), .A3(new_n1213), .ZN(new_n1214));
  INV_X1    g789(.A(new_n1005), .ZN(new_n1215));
  XNOR2_X1  g790(.A(G290), .B(new_n714), .ZN(new_n1216));
  AOI21_X1  g791(.A(new_n989), .B1(new_n1215), .B2(new_n1216), .ZN(new_n1217));
  OAI21_X1  g792(.A(new_n1011), .B1(new_n1214), .B2(new_n1217), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g793(.A(G401), .ZN(new_n1220));
  INV_X1    g794(.A(G319), .ZN(new_n1221));
  NOR2_X1   g795(.A1(G227), .A2(new_n1221), .ZN(new_n1222));
  XOR2_X1   g796(.A(new_n1222), .B(KEYINPUT127), .Z(new_n1223));
  AND3_X1   g797(.A1(new_n685), .A2(new_n1220), .A3(new_n1223), .ZN(new_n1224));
  NAND3_X1  g798(.A1(new_n975), .A2(new_n900), .A3(new_n1224), .ZN(G225));
  INV_X1    g799(.A(G225), .ZN(G308));
endmodule


