

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n522, n523, n524, n525,
         n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536,
         n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547,
         n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558,
         n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569,
         n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580,
         n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591,
         n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602,
         n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613,
         n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624,
         n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635,
         n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646,
         n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657,
         n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668,
         n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679,
         n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690,
         n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701,
         n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712,
         n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723,
         n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734,
         n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745,
         n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756,
         n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n767,
         n768, n769, n770, n771, n772, n773, n774, n775, n776, n777, n778,
         n779, n780, n781, n782, n783, n784, n785, n786, n787, n788, n789,
         n790, n791, n792, n793, n794, n795, n796, n797, n798, n799, n800,
         n801, n802, n803, n804, n805, n806, n807, n808, n809, n810, n811,
         n812, n813, n814, n815, n816, n817, n818, n819, n820, n821, n822,
         n823, n824, n825, n826, n827, n828, n829, n830, n831, n832, n833,
         n834, n835, n836, n837, n838, n839, n840, n841, n842, n843, n844,
         n845, n846, n847, n848, n849, n850, n851, n852, n853, n854, n855,
         n856, n857, n858, n859, n860, n861, n862, n863, n864, n865, n866,
         n867, n868, n869, n870, n871, n872, n873, n874, n875, n876, n877,
         n878, n879, n880, n881, n882, n883, n884, n885, n886, n887, n888,
         n889, n890, n891, n892, n893, n894, n895, n896, n897, n898, n899,
         n900, n901, n902, n903, n904, n905, n906, n907, n908, n909, n910,
         n911, n912, n913, n914, n915, n916, n917, n918, n919, n920, n921,
         n922, n923, n924, n925, n926, n927, n928, n929, n930, n931, n932,
         n933, n934, n935, n936, n937, n938, n939, n940, n941, n942, n943,
         n944, n945, n946, n947, n948, n949, n950, n951, n952, n953, n954,
         n955, n956, n957, n958, n959, n960, n961, n962, n963, n964, n965,
         n966, n967, n968, n969, n970, n971, n972, n973, n974, n975, n976,
         n977, n978, n979, n980, n981, n982, n983, n984, n985, n986, n987,
         n988, n989, n990, n991, n992, n993, n994, n995, n996, n997, n998,
         n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008,
         n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018,
         n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028,
         n1029, n1030, n1031, n1032, n1033;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  AND2_X1 U554 ( .A1(n745), .A2(n522), .ZN(n746) );
  NOR2_X2 U555 ( .A1(n702), .A2(n701), .ZN(n709) );
  OR2_X1 U556 ( .A1(n679), .A2(n656), .ZN(n657) );
  NOR2_X1 U557 ( .A1(n803), .A2(n647), .ZN(n648) );
  NOR2_X1 U558 ( .A1(n593), .A2(n711), .ZN(n639) );
  NOR2_X1 U559 ( .A1(n766), .A2(G1384), .ZN(n712) );
  XNOR2_X1 U560 ( .A(n710), .B(KEYINPUT104), .ZN(n745) );
  AND2_X1 U561 ( .A1(n756), .A2(n749), .ZN(n522) );
  NOR2_X1 U562 ( .A1(n707), .A2(n689), .ZN(n523) );
  INV_X1 U563 ( .A(KEYINPUT26), .ZN(n618) );
  XNOR2_X1 U564 ( .A(KEYINPUT97), .B(KEYINPUT27), .ZN(n640) );
  XNOR2_X1 U565 ( .A(n641), .B(n640), .ZN(n644) );
  INV_X1 U566 ( .A(n639), .ZN(n664) );
  NAND2_X1 U567 ( .A1(n889), .A2(G138), .ZN(n585) );
  INV_X1 U568 ( .A(KEYINPUT17), .ZN(n524) );
  NOR2_X1 U569 ( .A1(G651), .A2(G543), .ZN(n792) );
  XNOR2_X1 U570 ( .A(n530), .B(KEYINPUT65), .ZN(n895) );
  NOR2_X1 U571 ( .A1(G651), .A2(n564), .ZN(n797) );
  NOR2_X1 U572 ( .A1(n534), .A2(n533), .ZN(G160) );
  NOR2_X1 U573 ( .A1(G2104), .A2(G2105), .ZN(n525) );
  XNOR2_X2 U574 ( .A(n525), .B(n524), .ZN(n889) );
  NAND2_X1 U575 ( .A1(n889), .A2(G137), .ZN(n528) );
  XOR2_X1 U576 ( .A(G2104), .B(KEYINPUT64), .Z(n529) );
  NOR2_X1 U577 ( .A1(n529), .A2(G2105), .ZN(n713) );
  NAND2_X1 U578 ( .A1(G101), .A2(n713), .ZN(n526) );
  XOR2_X1 U579 ( .A(KEYINPUT23), .B(n526), .Z(n527) );
  NAND2_X1 U580 ( .A1(n528), .A2(n527), .ZN(n534) );
  AND2_X1 U581 ( .A1(G2105), .A2(n529), .ZN(n893) );
  NAND2_X1 U582 ( .A1(G125), .A2(n893), .ZN(n532) );
  NAND2_X1 U583 ( .A1(G2105), .A2(G2104), .ZN(n530) );
  NAND2_X1 U584 ( .A1(G113), .A2(n895), .ZN(n531) );
  NAND2_X1 U585 ( .A1(n532), .A2(n531), .ZN(n533) );
  XNOR2_X1 U586 ( .A(KEYINPUT67), .B(KEYINPUT9), .ZN(n538) );
  NAND2_X1 U587 ( .A1(G90), .A2(n792), .ZN(n536) );
  XOR2_X1 U588 ( .A(KEYINPUT0), .B(G543), .Z(n564) );
  INV_X1 U589 ( .A(G651), .ZN(n539) );
  NOR2_X1 U590 ( .A1(n564), .A2(n539), .ZN(n793) );
  NAND2_X1 U591 ( .A1(G77), .A2(n793), .ZN(n535) );
  NAND2_X1 U592 ( .A1(n536), .A2(n535), .ZN(n537) );
  XNOR2_X1 U593 ( .A(n538), .B(n537), .ZN(n543) );
  NOR2_X1 U594 ( .A1(G543), .A2(n539), .ZN(n540) );
  XOR2_X1 U595 ( .A(KEYINPUT1), .B(n540), .Z(n796) );
  NAND2_X1 U596 ( .A1(n796), .A2(G64), .ZN(n541) );
  XOR2_X1 U597 ( .A(KEYINPUT66), .B(n541), .Z(n542) );
  NOR2_X1 U598 ( .A1(n543), .A2(n542), .ZN(n545) );
  NAND2_X1 U599 ( .A1(n797), .A2(G52), .ZN(n544) );
  NAND2_X1 U600 ( .A1(n545), .A2(n544), .ZN(G301) );
  INV_X1 U601 ( .A(G301), .ZN(G171) );
  NAND2_X1 U602 ( .A1(n792), .A2(G89), .ZN(n546) );
  XNOR2_X1 U603 ( .A(n546), .B(KEYINPUT4), .ZN(n548) );
  NAND2_X1 U604 ( .A1(G76), .A2(n793), .ZN(n547) );
  NAND2_X1 U605 ( .A1(n548), .A2(n547), .ZN(n549) );
  XNOR2_X1 U606 ( .A(n549), .B(KEYINPUT5), .ZN(n554) );
  NAND2_X1 U607 ( .A1(G63), .A2(n796), .ZN(n551) );
  NAND2_X1 U608 ( .A1(G51), .A2(n797), .ZN(n550) );
  NAND2_X1 U609 ( .A1(n551), .A2(n550), .ZN(n552) );
  XOR2_X1 U610 ( .A(KEYINPUT6), .B(n552), .Z(n553) );
  NAND2_X1 U611 ( .A1(n554), .A2(n553), .ZN(n555) );
  XNOR2_X1 U612 ( .A(n555), .B(KEYINPUT7), .ZN(G168) );
  NAND2_X1 U613 ( .A1(G88), .A2(n792), .ZN(n556) );
  XNOR2_X1 U614 ( .A(n556), .B(KEYINPUT82), .ZN(n563) );
  NAND2_X1 U615 ( .A1(G75), .A2(n793), .ZN(n558) );
  NAND2_X1 U616 ( .A1(G62), .A2(n796), .ZN(n557) );
  NAND2_X1 U617 ( .A1(n558), .A2(n557), .ZN(n561) );
  NAND2_X1 U618 ( .A1(G50), .A2(n797), .ZN(n559) );
  XNOR2_X1 U619 ( .A(KEYINPUT81), .B(n559), .ZN(n560) );
  NOR2_X1 U620 ( .A1(n561), .A2(n560), .ZN(n562) );
  NAND2_X1 U621 ( .A1(n563), .A2(n562), .ZN(G303) );
  XOR2_X1 U622 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U623 ( .A1(G74), .A2(G651), .ZN(n569) );
  NAND2_X1 U624 ( .A1(G49), .A2(n797), .ZN(n566) );
  NAND2_X1 U625 ( .A1(G87), .A2(n564), .ZN(n565) );
  NAND2_X1 U626 ( .A1(n566), .A2(n565), .ZN(n567) );
  NOR2_X1 U627 ( .A1(n796), .A2(n567), .ZN(n568) );
  NAND2_X1 U628 ( .A1(n569), .A2(n568), .ZN(n570) );
  XNOR2_X1 U629 ( .A(n570), .B(KEYINPUT80), .ZN(G288) );
  NAND2_X1 U630 ( .A1(G86), .A2(n792), .ZN(n572) );
  NAND2_X1 U631 ( .A1(G61), .A2(n796), .ZN(n571) );
  NAND2_X1 U632 ( .A1(n572), .A2(n571), .ZN(n575) );
  NAND2_X1 U633 ( .A1(n793), .A2(G73), .ZN(n573) );
  XOR2_X1 U634 ( .A(KEYINPUT2), .B(n573), .Z(n574) );
  NOR2_X1 U635 ( .A1(n575), .A2(n574), .ZN(n577) );
  NAND2_X1 U636 ( .A1(n797), .A2(G48), .ZN(n576) );
  NAND2_X1 U637 ( .A1(n577), .A2(n576), .ZN(G305) );
  NAND2_X1 U638 ( .A1(G85), .A2(n792), .ZN(n579) );
  NAND2_X1 U639 ( .A1(G72), .A2(n793), .ZN(n578) );
  NAND2_X1 U640 ( .A1(n579), .A2(n578), .ZN(n583) );
  NAND2_X1 U641 ( .A1(G60), .A2(n796), .ZN(n581) );
  NAND2_X1 U642 ( .A1(G47), .A2(n797), .ZN(n580) );
  NAND2_X1 U643 ( .A1(n581), .A2(n580), .ZN(n582) );
  OR2_X1 U644 ( .A1(n583), .A2(n582), .ZN(G290) );
  NAND2_X1 U645 ( .A1(n713), .A2(G102), .ZN(n584) );
  NAND2_X1 U646 ( .A1(n585), .A2(n584), .ZN(n587) );
  INV_X1 U647 ( .A(KEYINPUT86), .ZN(n586) );
  XNOR2_X1 U648 ( .A(n587), .B(n586), .ZN(n589) );
  NAND2_X1 U649 ( .A1(n895), .A2(G114), .ZN(n588) );
  NAND2_X1 U650 ( .A1(n589), .A2(n588), .ZN(n592) );
  NAND2_X1 U651 ( .A1(G126), .A2(n893), .ZN(n590) );
  XNOR2_X1 U652 ( .A(KEYINPUT85), .B(n590), .ZN(n591) );
  NOR2_X1 U653 ( .A1(n592), .A2(n591), .ZN(n766) );
  INV_X1 U654 ( .A(n712), .ZN(n593) );
  NAND2_X1 U655 ( .A1(G160), .A2(G40), .ZN(n711) );
  INV_X1 U656 ( .A(n664), .ZN(n642) );
  NOR2_X1 U657 ( .A1(n642), .A2(G1961), .ZN(n594) );
  XOR2_X1 U658 ( .A(KEYINPUT96), .B(n594), .Z(n596) );
  XNOR2_X1 U659 ( .A(G2078), .B(KEYINPUT25), .ZN(n954) );
  NAND2_X1 U660 ( .A1(n642), .A2(n954), .ZN(n595) );
  NAND2_X1 U661 ( .A1(n596), .A2(n595), .ZN(n654) );
  NAND2_X1 U662 ( .A1(n654), .A2(G171), .ZN(n653) );
  NAND2_X1 U663 ( .A1(G66), .A2(n796), .ZN(n605) );
  NAND2_X1 U664 ( .A1(G79), .A2(n793), .ZN(n597) );
  XNOR2_X1 U665 ( .A(n597), .B(KEYINPUT74), .ZN(n600) );
  NAND2_X1 U666 ( .A1(G54), .A2(n797), .ZN(n598) );
  XOR2_X1 U667 ( .A(KEYINPUT75), .B(n598), .Z(n599) );
  NAND2_X1 U668 ( .A1(n600), .A2(n599), .ZN(n603) );
  NAND2_X1 U669 ( .A1(G92), .A2(n792), .ZN(n601) );
  XNOR2_X1 U670 ( .A(KEYINPUT73), .B(n601), .ZN(n602) );
  NOR2_X1 U671 ( .A1(n603), .A2(n602), .ZN(n604) );
  NAND2_X1 U672 ( .A1(n605), .A2(n604), .ZN(n606) );
  XNOR2_X1 U673 ( .A(n606), .B(KEYINPUT15), .ZN(n991) );
  NAND2_X1 U674 ( .A1(n792), .A2(G81), .ZN(n607) );
  XNOR2_X1 U675 ( .A(KEYINPUT12), .B(n607), .ZN(n610) );
  NAND2_X1 U676 ( .A1(n793), .A2(G68), .ZN(n608) );
  XOR2_X1 U677 ( .A(KEYINPUT71), .B(n608), .Z(n609) );
  NAND2_X1 U678 ( .A1(n610), .A2(n609), .ZN(n611) );
  XNOR2_X1 U679 ( .A(KEYINPUT13), .B(n611), .ZN(n617) );
  NAND2_X1 U680 ( .A1(G56), .A2(n796), .ZN(n612) );
  XOR2_X1 U681 ( .A(KEYINPUT14), .B(n612), .Z(n615) );
  NAND2_X1 U682 ( .A1(n797), .A2(G43), .ZN(n613) );
  XOR2_X1 U683 ( .A(KEYINPUT72), .B(n613), .Z(n614) );
  NOR2_X1 U684 ( .A1(n615), .A2(n614), .ZN(n616) );
  NAND2_X1 U685 ( .A1(n617), .A2(n616), .ZN(n975) );
  INV_X1 U686 ( .A(G1996), .ZN(n861) );
  NOR2_X1 U687 ( .A1(n664), .A2(n861), .ZN(n619) );
  XNOR2_X1 U688 ( .A(n619), .B(n618), .ZN(n621) );
  NAND2_X1 U689 ( .A1(n664), .A2(G1341), .ZN(n620) );
  NAND2_X1 U690 ( .A1(n621), .A2(n620), .ZN(n622) );
  NOR2_X1 U691 ( .A1(n975), .A2(n622), .ZN(n628) );
  NAND2_X1 U692 ( .A1(n991), .A2(n628), .ZN(n627) );
  NAND2_X1 U693 ( .A1(n664), .A2(G1348), .ZN(n623) );
  XNOR2_X1 U694 ( .A(n623), .B(KEYINPUT98), .ZN(n625) );
  NAND2_X1 U695 ( .A1(n642), .A2(G2067), .ZN(n624) );
  NAND2_X1 U696 ( .A1(n625), .A2(n624), .ZN(n626) );
  NAND2_X1 U697 ( .A1(n627), .A2(n626), .ZN(n630) );
  OR2_X1 U698 ( .A1(n991), .A2(n628), .ZN(n629) );
  NAND2_X1 U699 ( .A1(n630), .A2(n629), .ZN(n646) );
  NAND2_X1 U700 ( .A1(G91), .A2(n792), .ZN(n632) );
  NAND2_X1 U701 ( .A1(G78), .A2(n793), .ZN(n631) );
  NAND2_X1 U702 ( .A1(n632), .A2(n631), .ZN(n637) );
  NAND2_X1 U703 ( .A1(G65), .A2(n796), .ZN(n634) );
  NAND2_X1 U704 ( .A1(G53), .A2(n797), .ZN(n633) );
  NAND2_X1 U705 ( .A1(n634), .A2(n633), .ZN(n635) );
  XNOR2_X1 U706 ( .A(KEYINPUT68), .B(n635), .ZN(n636) );
  NOR2_X1 U707 ( .A1(n637), .A2(n636), .ZN(n638) );
  XOR2_X1 U708 ( .A(n638), .B(KEYINPUT69), .Z(n803) );
  AND2_X1 U709 ( .A1(G2072), .A2(n639), .ZN(n641) );
  INV_X1 U710 ( .A(G1956), .ZN(n860) );
  NOR2_X1 U711 ( .A1(n642), .A2(n860), .ZN(n643) );
  NOR2_X1 U712 ( .A1(n644), .A2(n643), .ZN(n647) );
  NAND2_X1 U713 ( .A1(n803), .A2(n647), .ZN(n645) );
  NAND2_X1 U714 ( .A1(n646), .A2(n645), .ZN(n650) );
  XOR2_X1 U715 ( .A(n648), .B(KEYINPUT28), .Z(n649) );
  NAND2_X1 U716 ( .A1(n650), .A2(n649), .ZN(n651) );
  XOR2_X1 U717 ( .A(KEYINPUT29), .B(n651), .Z(n652) );
  NAND2_X1 U718 ( .A1(n653), .A2(n652), .ZN(n677) );
  NOR2_X1 U719 ( .A1(G171), .A2(n654), .ZN(n660) );
  NAND2_X1 U720 ( .A1(G8), .A2(n664), .ZN(n707) );
  NOR2_X1 U721 ( .A1(G1966), .A2(n707), .ZN(n679) );
  NOR2_X1 U722 ( .A1(G2084), .A2(n664), .ZN(n680) );
  INV_X1 U723 ( .A(G8), .ZN(n655) );
  OR2_X1 U724 ( .A1(n680), .A2(n655), .ZN(n656) );
  XNOR2_X1 U725 ( .A(KEYINPUT30), .B(n657), .ZN(n658) );
  NOR2_X1 U726 ( .A1(G168), .A2(n658), .ZN(n659) );
  NOR2_X1 U727 ( .A1(n660), .A2(n659), .ZN(n663) );
  XNOR2_X1 U728 ( .A(KEYINPUT99), .B(KEYINPUT100), .ZN(n661) );
  XNOR2_X1 U729 ( .A(n661), .B(KEYINPUT31), .ZN(n662) );
  XNOR2_X1 U730 ( .A(n663), .B(n662), .ZN(n676) );
  NOR2_X1 U731 ( .A1(G1971), .A2(n707), .ZN(n666) );
  NOR2_X1 U732 ( .A1(G2090), .A2(n664), .ZN(n665) );
  NOR2_X1 U733 ( .A1(n666), .A2(n665), .ZN(n667) );
  NAND2_X1 U734 ( .A1(n667), .A2(G303), .ZN(n668) );
  OR2_X1 U735 ( .A1(n655), .A2(n668), .ZN(n670) );
  AND2_X1 U736 ( .A1(n676), .A2(n670), .ZN(n669) );
  NAND2_X1 U737 ( .A1(n677), .A2(n669), .ZN(n673) );
  INV_X1 U738 ( .A(n670), .ZN(n671) );
  OR2_X1 U739 ( .A1(n671), .A2(G286), .ZN(n672) );
  NAND2_X1 U740 ( .A1(n673), .A2(n672), .ZN(n675) );
  XOR2_X1 U741 ( .A(KEYINPUT32), .B(KEYINPUT101), .Z(n674) );
  XNOR2_X1 U742 ( .A(n675), .B(n674), .ZN(n684) );
  AND2_X1 U743 ( .A1(n677), .A2(n676), .ZN(n678) );
  NOR2_X1 U744 ( .A1(n679), .A2(n678), .ZN(n682) );
  NAND2_X1 U745 ( .A1(G8), .A2(n680), .ZN(n681) );
  NAND2_X1 U746 ( .A1(n682), .A2(n681), .ZN(n683) );
  NAND2_X1 U747 ( .A1(n684), .A2(n683), .ZN(n705) );
  NOR2_X1 U748 ( .A1(G1976), .A2(G288), .ZN(n980) );
  NOR2_X1 U749 ( .A1(G1971), .A2(G303), .ZN(n979) );
  XNOR2_X1 U750 ( .A(KEYINPUT102), .B(n979), .ZN(n685) );
  NOR2_X1 U751 ( .A1(n980), .A2(n685), .ZN(n687) );
  INV_X1 U752 ( .A(KEYINPUT33), .ZN(n686) );
  AND2_X1 U753 ( .A1(n687), .A2(n686), .ZN(n688) );
  NAND2_X1 U754 ( .A1(n705), .A2(n688), .ZN(n695) );
  NAND2_X1 U755 ( .A1(G1976), .A2(G288), .ZN(n977) );
  INV_X1 U756 ( .A(n977), .ZN(n689) );
  OR2_X1 U757 ( .A1(KEYINPUT33), .A2(n523), .ZN(n692) );
  NAND2_X1 U758 ( .A1(n980), .A2(KEYINPUT33), .ZN(n690) );
  OR2_X1 U759 ( .A1(n690), .A2(n707), .ZN(n691) );
  AND2_X1 U760 ( .A1(n692), .A2(n691), .ZN(n693) );
  XOR2_X1 U761 ( .A(G1981), .B(G305), .Z(n972) );
  AND2_X1 U762 ( .A1(n693), .A2(n972), .ZN(n694) );
  NAND2_X1 U763 ( .A1(n695), .A2(n694), .ZN(n696) );
  XNOR2_X1 U764 ( .A(n696), .B(KEYINPUT103), .ZN(n702) );
  NOR2_X1 U765 ( .A1(G1981), .A2(G305), .ZN(n699) );
  XNOR2_X1 U766 ( .A(KEYINPUT24), .B(KEYINPUT95), .ZN(n697) );
  XNOR2_X1 U767 ( .A(n697), .B(KEYINPUT94), .ZN(n698) );
  XNOR2_X1 U768 ( .A(n699), .B(n698), .ZN(n700) );
  NOR2_X1 U769 ( .A1(n707), .A2(n700), .ZN(n701) );
  NOR2_X1 U770 ( .A1(G2090), .A2(G303), .ZN(n703) );
  NAND2_X1 U771 ( .A1(G8), .A2(n703), .ZN(n704) );
  NAND2_X1 U772 ( .A1(n705), .A2(n704), .ZN(n706) );
  NAND2_X1 U773 ( .A1(n707), .A2(n706), .ZN(n708) );
  NAND2_X1 U774 ( .A1(n709), .A2(n708), .ZN(n710) );
  NOR2_X1 U775 ( .A1(n712), .A2(n711), .ZN(n761) );
  NAND2_X1 U776 ( .A1(G140), .A2(n889), .ZN(n715) );
  BUF_X1 U777 ( .A(n713), .Z(n890) );
  NAND2_X1 U778 ( .A1(G104), .A2(n890), .ZN(n714) );
  NAND2_X1 U779 ( .A1(n715), .A2(n714), .ZN(n717) );
  XOR2_X1 U780 ( .A(KEYINPUT34), .B(KEYINPUT87), .Z(n716) );
  XNOR2_X1 U781 ( .A(n717), .B(n716), .ZN(n722) );
  NAND2_X1 U782 ( .A1(G128), .A2(n893), .ZN(n719) );
  NAND2_X1 U783 ( .A1(G116), .A2(n895), .ZN(n718) );
  NAND2_X1 U784 ( .A1(n719), .A2(n718), .ZN(n720) );
  XOR2_X1 U785 ( .A(KEYINPUT35), .B(n720), .Z(n721) );
  NOR2_X1 U786 ( .A1(n722), .A2(n721), .ZN(n723) );
  XNOR2_X1 U787 ( .A(n723), .B(KEYINPUT36), .ZN(n724) );
  XNOR2_X1 U788 ( .A(n724), .B(KEYINPUT88), .ZN(n907) );
  XNOR2_X1 U789 ( .A(G2067), .B(KEYINPUT37), .ZN(n759) );
  NOR2_X1 U790 ( .A1(n907), .A2(n759), .ZN(n935) );
  NAND2_X1 U791 ( .A1(n761), .A2(n935), .ZN(n756) );
  NAND2_X1 U792 ( .A1(G141), .A2(n889), .ZN(n726) );
  NAND2_X1 U793 ( .A1(G129), .A2(n893), .ZN(n725) );
  NAND2_X1 U794 ( .A1(n726), .A2(n725), .ZN(n729) );
  NAND2_X1 U795 ( .A1(n890), .A2(G105), .ZN(n727) );
  XOR2_X1 U796 ( .A(KEYINPUT38), .B(n727), .Z(n728) );
  NOR2_X1 U797 ( .A1(n729), .A2(n728), .ZN(n731) );
  NAND2_X1 U798 ( .A1(n895), .A2(G117), .ZN(n730) );
  NAND2_X1 U799 ( .A1(n731), .A2(n730), .ZN(n877) );
  NAND2_X1 U800 ( .A1(G1996), .A2(n877), .ZN(n732) );
  XNOR2_X1 U801 ( .A(KEYINPUT93), .B(n732), .ZN(n743) );
  NAND2_X1 U802 ( .A1(G95), .A2(n890), .ZN(n733) );
  XOR2_X1 U803 ( .A(KEYINPUT90), .B(n733), .Z(n738) );
  NAND2_X1 U804 ( .A1(G119), .A2(n893), .ZN(n735) );
  NAND2_X1 U805 ( .A1(G107), .A2(n895), .ZN(n734) );
  NAND2_X1 U806 ( .A1(n735), .A2(n734), .ZN(n736) );
  XOR2_X1 U807 ( .A(KEYINPUT89), .B(n736), .Z(n737) );
  NOR2_X1 U808 ( .A1(n738), .A2(n737), .ZN(n740) );
  NAND2_X1 U809 ( .A1(n889), .A2(G131), .ZN(n739) );
  AND2_X1 U810 ( .A1(n740), .A2(n739), .ZN(n902) );
  XNOR2_X1 U811 ( .A(KEYINPUT91), .B(G1991), .ZN(n955) );
  NOR2_X1 U812 ( .A1(n902), .A2(n955), .ZN(n741) );
  XNOR2_X1 U813 ( .A(n741), .B(KEYINPUT92), .ZN(n742) );
  NOR2_X1 U814 ( .A1(n743), .A2(n742), .ZN(n944) );
  INV_X1 U815 ( .A(n944), .ZN(n744) );
  NAND2_X1 U816 ( .A1(n744), .A2(n761), .ZN(n749) );
  XOR2_X1 U817 ( .A(KEYINPUT105), .B(n746), .Z(n748) );
  XNOR2_X1 U818 ( .A(G1986), .B(G290), .ZN(n978) );
  NAND2_X1 U819 ( .A1(n978), .A2(n761), .ZN(n747) );
  NAND2_X1 U820 ( .A1(n748), .A2(n747), .ZN(n764) );
  NOR2_X1 U821 ( .A1(G1996), .A2(n877), .ZN(n924) );
  INV_X1 U822 ( .A(n749), .ZN(n752) );
  AND2_X1 U823 ( .A1(n955), .A2(n902), .ZN(n930) );
  NOR2_X1 U824 ( .A1(G1986), .A2(G290), .ZN(n750) );
  NOR2_X1 U825 ( .A1(n930), .A2(n750), .ZN(n751) );
  NOR2_X1 U826 ( .A1(n752), .A2(n751), .ZN(n753) );
  NOR2_X1 U827 ( .A1(n924), .A2(n753), .ZN(n754) );
  XNOR2_X1 U828 ( .A(KEYINPUT39), .B(n754), .ZN(n755) );
  XNOR2_X1 U829 ( .A(n755), .B(KEYINPUT106), .ZN(n757) );
  NAND2_X1 U830 ( .A1(n757), .A2(n756), .ZN(n758) );
  XOR2_X1 U831 ( .A(KEYINPUT107), .B(n758), .Z(n760) );
  NAND2_X1 U832 ( .A1(n907), .A2(n759), .ZN(n927) );
  NAND2_X1 U833 ( .A1(n760), .A2(n927), .ZN(n762) );
  NAND2_X1 U834 ( .A1(n762), .A2(n761), .ZN(n763) );
  NAND2_X1 U835 ( .A1(n764), .A2(n763), .ZN(n765) );
  XNOR2_X1 U836 ( .A(n765), .B(KEYINPUT40), .ZN(G329) );
  AND2_X1 U837 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U838 ( .A(G57), .ZN(G237) );
  INV_X1 U839 ( .A(G132), .ZN(G219) );
  INV_X1 U840 ( .A(G82), .ZN(G220) );
  BUF_X1 U841 ( .A(n766), .Z(G164) );
  NAND2_X1 U842 ( .A1(G7), .A2(G661), .ZN(n767) );
  XNOR2_X1 U843 ( .A(n767), .B(KEYINPUT10), .ZN(G223) );
  XOR2_X1 U844 ( .A(G223), .B(KEYINPUT70), .Z(n829) );
  NAND2_X1 U845 ( .A1(n829), .A2(G567), .ZN(n768) );
  XOR2_X1 U846 ( .A(KEYINPUT11), .B(n768), .Z(G234) );
  INV_X1 U847 ( .A(G860), .ZN(n791) );
  OR2_X1 U848 ( .A1(n975), .A2(n791), .ZN(G153) );
  NAND2_X1 U849 ( .A1(G868), .A2(G301), .ZN(n770) );
  OR2_X1 U850 ( .A1(n991), .A2(G868), .ZN(n769) );
  NAND2_X1 U851 ( .A1(n770), .A2(n769), .ZN(G284) );
  INV_X1 U852 ( .A(n803), .ZN(G299) );
  INV_X1 U853 ( .A(G868), .ZN(n813) );
  NOR2_X1 U854 ( .A1(G286), .A2(n813), .ZN(n771) );
  XNOR2_X1 U855 ( .A(n771), .B(KEYINPUT76), .ZN(n773) );
  NOR2_X1 U856 ( .A1(G299), .A2(G868), .ZN(n772) );
  NOR2_X1 U857 ( .A1(n773), .A2(n772), .ZN(G297) );
  NAND2_X1 U858 ( .A1(G559), .A2(n791), .ZN(n774) );
  XOR2_X1 U859 ( .A(KEYINPUT77), .B(n774), .Z(n775) );
  NAND2_X1 U860 ( .A1(n775), .A2(n991), .ZN(n776) );
  XNOR2_X1 U861 ( .A(n776), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U862 ( .A1(G868), .A2(n975), .ZN(n779) );
  NAND2_X1 U863 ( .A1(G868), .A2(n991), .ZN(n777) );
  NOR2_X1 U864 ( .A1(G559), .A2(n777), .ZN(n778) );
  NOR2_X1 U865 ( .A1(n779), .A2(n778), .ZN(G282) );
  NAND2_X1 U866 ( .A1(G123), .A2(n893), .ZN(n780) );
  XNOR2_X1 U867 ( .A(n780), .B(KEYINPUT18), .ZN(n782) );
  NAND2_X1 U868 ( .A1(n890), .A2(G99), .ZN(n781) );
  NAND2_X1 U869 ( .A1(n782), .A2(n781), .ZN(n786) );
  NAND2_X1 U870 ( .A1(G135), .A2(n889), .ZN(n784) );
  NAND2_X1 U871 ( .A1(G111), .A2(n895), .ZN(n783) );
  NAND2_X1 U872 ( .A1(n784), .A2(n783), .ZN(n785) );
  NOR2_X1 U873 ( .A1(n786), .A2(n785), .ZN(n929) );
  XNOR2_X1 U874 ( .A(n929), .B(G2096), .ZN(n787) );
  XNOR2_X1 U875 ( .A(n787), .B(KEYINPUT78), .ZN(n788) );
  INV_X1 U876 ( .A(G2100), .ZN(n853) );
  NAND2_X1 U877 ( .A1(n788), .A2(n853), .ZN(G156) );
  XNOR2_X1 U878 ( .A(n975), .B(KEYINPUT79), .ZN(n790) );
  NAND2_X1 U879 ( .A1(n991), .A2(G559), .ZN(n789) );
  XNOR2_X1 U880 ( .A(n790), .B(n789), .ZN(n810) );
  NAND2_X1 U881 ( .A1(n791), .A2(n810), .ZN(n802) );
  NAND2_X1 U882 ( .A1(G93), .A2(n792), .ZN(n795) );
  NAND2_X1 U883 ( .A1(G80), .A2(n793), .ZN(n794) );
  NAND2_X1 U884 ( .A1(n795), .A2(n794), .ZN(n801) );
  NAND2_X1 U885 ( .A1(G67), .A2(n796), .ZN(n799) );
  NAND2_X1 U886 ( .A1(G55), .A2(n797), .ZN(n798) );
  NAND2_X1 U887 ( .A1(n799), .A2(n798), .ZN(n800) );
  NOR2_X1 U888 ( .A1(n801), .A2(n800), .ZN(n812) );
  XOR2_X1 U889 ( .A(n802), .B(n812), .Z(G145) );
  XOR2_X1 U890 ( .A(G303), .B(n812), .Z(n809) );
  XOR2_X1 U891 ( .A(G288), .B(n803), .Z(n804) );
  XNOR2_X1 U892 ( .A(n804), .B(G305), .ZN(n805) );
  XNOR2_X1 U893 ( .A(KEYINPUT83), .B(n805), .ZN(n807) );
  XNOR2_X1 U894 ( .A(G290), .B(KEYINPUT19), .ZN(n806) );
  XNOR2_X1 U895 ( .A(n807), .B(n806), .ZN(n808) );
  XNOR2_X1 U896 ( .A(n809), .B(n808), .ZN(n912) );
  XOR2_X1 U897 ( .A(n912), .B(n810), .Z(n811) );
  NOR2_X1 U898 ( .A1(n813), .A2(n811), .ZN(n815) );
  AND2_X1 U899 ( .A1(n813), .A2(n812), .ZN(n814) );
  NOR2_X1 U900 ( .A1(n815), .A2(n814), .ZN(G295) );
  NAND2_X1 U901 ( .A1(G2084), .A2(G2078), .ZN(n816) );
  XOR2_X1 U902 ( .A(KEYINPUT20), .B(n816), .Z(n817) );
  NAND2_X1 U903 ( .A1(G2090), .A2(n817), .ZN(n818) );
  XNOR2_X1 U904 ( .A(KEYINPUT21), .B(n818), .ZN(n819) );
  NAND2_X1 U905 ( .A1(n819), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U906 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U907 ( .A1(G220), .A2(G219), .ZN(n820) );
  XOR2_X1 U908 ( .A(KEYINPUT22), .B(n820), .Z(n821) );
  NOR2_X1 U909 ( .A1(G218), .A2(n821), .ZN(n822) );
  NAND2_X1 U910 ( .A1(G96), .A2(n822), .ZN(n833) );
  NAND2_X1 U911 ( .A1(n833), .A2(G2106), .ZN(n826) );
  NAND2_X1 U912 ( .A1(G69), .A2(G120), .ZN(n823) );
  NOR2_X1 U913 ( .A1(G237), .A2(n823), .ZN(n824) );
  NAND2_X1 U914 ( .A1(G108), .A2(n824), .ZN(n834) );
  NAND2_X1 U915 ( .A1(n834), .A2(G567), .ZN(n825) );
  NAND2_X1 U916 ( .A1(n826), .A2(n825), .ZN(n922) );
  NAND2_X1 U917 ( .A1(G483), .A2(G661), .ZN(n827) );
  NOR2_X1 U918 ( .A1(n922), .A2(n827), .ZN(n832) );
  NAND2_X1 U919 ( .A1(n832), .A2(G36), .ZN(n828) );
  XNOR2_X1 U920 ( .A(KEYINPUT84), .B(n828), .ZN(G176) );
  INV_X1 U921 ( .A(G303), .ZN(G166) );
  NAND2_X1 U922 ( .A1(G2106), .A2(n829), .ZN(G217) );
  AND2_X1 U923 ( .A1(G15), .A2(G2), .ZN(n830) );
  NAND2_X1 U924 ( .A1(G661), .A2(n830), .ZN(G259) );
  NAND2_X1 U925 ( .A1(G3), .A2(G1), .ZN(n831) );
  NAND2_X1 U926 ( .A1(n832), .A2(n831), .ZN(G188) );
  INV_X1 U928 ( .A(G120), .ZN(G236) );
  INV_X1 U929 ( .A(G96), .ZN(G221) );
  INV_X1 U930 ( .A(G69), .ZN(G235) );
  NOR2_X1 U931 ( .A1(n834), .A2(n833), .ZN(G325) );
  INV_X1 U932 ( .A(G325), .ZN(G261) );
  XNOR2_X1 U933 ( .A(G1348), .B(G1341), .ZN(n835) );
  XNOR2_X1 U934 ( .A(n835), .B(G2427), .ZN(n845) );
  XOR2_X1 U935 ( .A(G2446), .B(G2430), .Z(n837) );
  XNOR2_X1 U936 ( .A(KEYINPUT108), .B(G2451), .ZN(n836) );
  XNOR2_X1 U937 ( .A(n837), .B(n836), .ZN(n841) );
  XOR2_X1 U938 ( .A(G2438), .B(G2435), .Z(n839) );
  XNOR2_X1 U939 ( .A(KEYINPUT109), .B(G2454), .ZN(n838) );
  XNOR2_X1 U940 ( .A(n839), .B(n838), .ZN(n840) );
  XOR2_X1 U941 ( .A(n841), .B(n840), .Z(n843) );
  XNOR2_X1 U942 ( .A(KEYINPUT110), .B(G2443), .ZN(n842) );
  XNOR2_X1 U943 ( .A(n843), .B(n842), .ZN(n844) );
  XNOR2_X1 U944 ( .A(n845), .B(n844), .ZN(n846) );
  NAND2_X1 U945 ( .A1(n846), .A2(G14), .ZN(n847) );
  XNOR2_X1 U946 ( .A(n847), .B(KEYINPUT111), .ZN(G401) );
  XOR2_X1 U947 ( .A(G2096), .B(KEYINPUT43), .Z(n849) );
  XNOR2_X1 U948 ( .A(G2072), .B(G2678), .ZN(n848) );
  XNOR2_X1 U949 ( .A(n849), .B(n848), .ZN(n850) );
  XOR2_X1 U950 ( .A(n850), .B(KEYINPUT42), .Z(n852) );
  XNOR2_X1 U951 ( .A(G2067), .B(G2090), .ZN(n851) );
  XNOR2_X1 U952 ( .A(n852), .B(n851), .ZN(n857) );
  XNOR2_X1 U953 ( .A(KEYINPUT112), .B(n853), .ZN(n855) );
  XNOR2_X1 U954 ( .A(G2084), .B(G2078), .ZN(n854) );
  XNOR2_X1 U955 ( .A(n855), .B(n854), .ZN(n856) );
  XNOR2_X1 U956 ( .A(n857), .B(n856), .ZN(G227) );
  XOR2_X1 U957 ( .A(G1971), .B(G1961), .Z(n859) );
  XNOR2_X1 U958 ( .A(G1986), .B(G1966), .ZN(n858) );
  XNOR2_X1 U959 ( .A(n859), .B(n858), .ZN(n865) );
  XNOR2_X1 U960 ( .A(G1976), .B(n860), .ZN(n863) );
  XOR2_X1 U961 ( .A(n861), .B(G1991), .Z(n862) );
  XNOR2_X1 U962 ( .A(n863), .B(n862), .ZN(n864) );
  XOR2_X1 U963 ( .A(n865), .B(n864), .Z(n867) );
  XNOR2_X1 U964 ( .A(KEYINPUT113), .B(G2474), .ZN(n866) );
  XNOR2_X1 U965 ( .A(n867), .B(n866), .ZN(n869) );
  XOR2_X1 U966 ( .A(G1981), .B(KEYINPUT41), .Z(n868) );
  XNOR2_X1 U967 ( .A(n869), .B(n868), .ZN(G229) );
  NAND2_X1 U968 ( .A1(G124), .A2(n893), .ZN(n870) );
  XNOR2_X1 U969 ( .A(n870), .B(KEYINPUT44), .ZN(n872) );
  NAND2_X1 U970 ( .A1(n890), .A2(G100), .ZN(n871) );
  NAND2_X1 U971 ( .A1(n872), .A2(n871), .ZN(n876) );
  NAND2_X1 U972 ( .A1(G136), .A2(n889), .ZN(n874) );
  NAND2_X1 U973 ( .A1(G112), .A2(n895), .ZN(n873) );
  NAND2_X1 U974 ( .A1(n874), .A2(n873), .ZN(n875) );
  NOR2_X1 U975 ( .A1(n876), .A2(n875), .ZN(G162) );
  XNOR2_X1 U976 ( .A(KEYINPUT48), .B(KEYINPUT46), .ZN(n879) );
  XNOR2_X1 U977 ( .A(n877), .B(KEYINPUT116), .ZN(n878) );
  XNOR2_X1 U978 ( .A(n879), .B(n878), .ZN(n880) );
  XNOR2_X1 U979 ( .A(G164), .B(n880), .ZN(n906) );
  NAND2_X1 U980 ( .A1(G130), .A2(n893), .ZN(n882) );
  NAND2_X1 U981 ( .A1(G118), .A2(n895), .ZN(n881) );
  NAND2_X1 U982 ( .A1(n882), .A2(n881), .ZN(n888) );
  NAND2_X1 U983 ( .A1(n889), .A2(G142), .ZN(n883) );
  XNOR2_X1 U984 ( .A(n883), .B(KEYINPUT114), .ZN(n885) );
  NAND2_X1 U985 ( .A1(G106), .A2(n890), .ZN(n884) );
  NAND2_X1 U986 ( .A1(n885), .A2(n884), .ZN(n886) );
  XOR2_X1 U987 ( .A(KEYINPUT45), .B(n886), .Z(n887) );
  NOR2_X1 U988 ( .A1(n888), .A2(n887), .ZN(n901) );
  NAND2_X1 U989 ( .A1(G139), .A2(n889), .ZN(n892) );
  NAND2_X1 U990 ( .A1(G103), .A2(n890), .ZN(n891) );
  NAND2_X1 U991 ( .A1(n892), .A2(n891), .ZN(n900) );
  NAND2_X1 U992 ( .A1(n893), .A2(G127), .ZN(n894) );
  XOR2_X1 U993 ( .A(KEYINPUT115), .B(n894), .Z(n897) );
  NAND2_X1 U994 ( .A1(n895), .A2(G115), .ZN(n896) );
  NAND2_X1 U995 ( .A1(n897), .A2(n896), .ZN(n898) );
  XOR2_X1 U996 ( .A(KEYINPUT47), .B(n898), .Z(n899) );
  NOR2_X1 U997 ( .A1(n900), .A2(n899), .ZN(n937) );
  XOR2_X1 U998 ( .A(n901), .B(n937), .Z(n904) );
  XNOR2_X1 U999 ( .A(G160), .B(n902), .ZN(n903) );
  XNOR2_X1 U1000 ( .A(n904), .B(n903), .ZN(n905) );
  XNOR2_X1 U1001 ( .A(n906), .B(n905), .ZN(n910) );
  XOR2_X1 U1002 ( .A(n907), .B(n929), .Z(n908) );
  XNOR2_X1 U1003 ( .A(G162), .B(n908), .ZN(n909) );
  XOR2_X1 U1004 ( .A(n910), .B(n909), .Z(n911) );
  NOR2_X1 U1005 ( .A1(G37), .A2(n911), .ZN(G395) );
  XOR2_X1 U1006 ( .A(n912), .B(G286), .Z(n914) );
  XOR2_X1 U1007 ( .A(G301), .B(n991), .Z(n913) );
  XNOR2_X1 U1008 ( .A(n914), .B(n913), .ZN(n915) );
  XNOR2_X1 U1009 ( .A(n915), .B(n975), .ZN(n916) );
  NOR2_X1 U1010 ( .A1(G37), .A2(n916), .ZN(G397) );
  OR2_X1 U1011 ( .A1(n922), .A2(G401), .ZN(n919) );
  NOR2_X1 U1012 ( .A1(G227), .A2(G229), .ZN(n917) );
  XNOR2_X1 U1013 ( .A(KEYINPUT49), .B(n917), .ZN(n918) );
  NOR2_X1 U1014 ( .A1(n919), .A2(n918), .ZN(n921) );
  NOR2_X1 U1015 ( .A1(G395), .A2(G397), .ZN(n920) );
  NAND2_X1 U1016 ( .A1(n921), .A2(n920), .ZN(G225) );
  INV_X1 U1017 ( .A(G225), .ZN(G308) );
  INV_X1 U1018 ( .A(n922), .ZN(G319) );
  INV_X1 U1019 ( .A(G108), .ZN(G238) );
  XOR2_X1 U1020 ( .A(G2090), .B(G162), .Z(n923) );
  NOR2_X1 U1021 ( .A1(n924), .A2(n923), .ZN(n925) );
  XNOR2_X1 U1022 ( .A(KEYINPUT51), .B(n925), .ZN(n926) );
  XNOR2_X1 U1023 ( .A(n926), .B(KEYINPUT119), .ZN(n928) );
  NAND2_X1 U1024 ( .A1(n928), .A2(n927), .ZN(n946) );
  NOR2_X1 U1025 ( .A1(n930), .A2(n929), .ZN(n931) );
  XOR2_X1 U1026 ( .A(KEYINPUT117), .B(n931), .Z(n933) );
  XNOR2_X1 U1027 ( .A(G160), .B(G2084), .ZN(n932) );
  NAND2_X1 U1028 ( .A1(n933), .A2(n932), .ZN(n934) );
  NOR2_X1 U1029 ( .A1(n935), .A2(n934), .ZN(n936) );
  XOR2_X1 U1030 ( .A(KEYINPUT118), .B(n936), .Z(n942) );
  XOR2_X1 U1031 ( .A(G2072), .B(n937), .Z(n939) );
  XOR2_X1 U1032 ( .A(G164), .B(G2078), .Z(n938) );
  NOR2_X1 U1033 ( .A1(n939), .A2(n938), .ZN(n940) );
  XOR2_X1 U1034 ( .A(KEYINPUT50), .B(n940), .Z(n941) );
  NOR2_X1 U1035 ( .A1(n942), .A2(n941), .ZN(n943) );
  NAND2_X1 U1036 ( .A1(n944), .A2(n943), .ZN(n945) );
  NOR2_X1 U1037 ( .A1(n946), .A2(n945), .ZN(n947) );
  XNOR2_X1 U1038 ( .A(KEYINPUT52), .B(n947), .ZN(n949) );
  INV_X1 U1039 ( .A(KEYINPUT55), .ZN(n948) );
  NAND2_X1 U1040 ( .A1(n949), .A2(n948), .ZN(n950) );
  NAND2_X1 U1041 ( .A1(n950), .A2(G29), .ZN(n1031) );
  XNOR2_X1 U1042 ( .A(G2090), .B(G35), .ZN(n964) );
  XOR2_X1 U1043 ( .A(G32), .B(G1996), .Z(n951) );
  NAND2_X1 U1044 ( .A1(n951), .A2(G28), .ZN(n961) );
  XNOR2_X1 U1045 ( .A(G2067), .B(G26), .ZN(n953) );
  XNOR2_X1 U1046 ( .A(G33), .B(G2072), .ZN(n952) );
  NOR2_X1 U1047 ( .A1(n953), .A2(n952), .ZN(n959) );
  XOR2_X1 U1048 ( .A(n954), .B(G27), .Z(n957) );
  XOR2_X1 U1049 ( .A(n955), .B(G25), .Z(n956) );
  NOR2_X1 U1050 ( .A1(n957), .A2(n956), .ZN(n958) );
  NAND2_X1 U1051 ( .A1(n959), .A2(n958), .ZN(n960) );
  NOR2_X1 U1052 ( .A1(n961), .A2(n960), .ZN(n962) );
  XNOR2_X1 U1053 ( .A(KEYINPUT53), .B(n962), .ZN(n963) );
  NOR2_X1 U1054 ( .A1(n964), .A2(n963), .ZN(n967) );
  XOR2_X1 U1055 ( .A(G2084), .B(G34), .Z(n965) );
  XNOR2_X1 U1056 ( .A(KEYINPUT54), .B(n965), .ZN(n966) );
  NAND2_X1 U1057 ( .A1(n967), .A2(n966), .ZN(n968) );
  XOR2_X1 U1058 ( .A(KEYINPUT55), .B(n968), .Z(n970) );
  INV_X1 U1059 ( .A(G29), .ZN(n969) );
  NAND2_X1 U1060 ( .A1(n970), .A2(n969), .ZN(n971) );
  NAND2_X1 U1061 ( .A1(G11), .A2(n971), .ZN(n1029) );
  INV_X1 U1062 ( .A(G16), .ZN(n1025) );
  XOR2_X1 U1063 ( .A(n1025), .B(KEYINPUT56), .Z(n1000) );
  XNOR2_X1 U1064 ( .A(G1966), .B(G168), .ZN(n973) );
  NAND2_X1 U1065 ( .A1(n973), .A2(n972), .ZN(n974) );
  XNOR2_X1 U1066 ( .A(n974), .B(KEYINPUT57), .ZN(n998) );
  XNOR2_X1 U1067 ( .A(n975), .B(G1341), .ZN(n996) );
  NAND2_X1 U1068 ( .A1(G1971), .A2(G303), .ZN(n976) );
  NAND2_X1 U1069 ( .A1(n977), .A2(n976), .ZN(n986) );
  NOR2_X1 U1070 ( .A1(n979), .A2(n978), .ZN(n984) );
  XOR2_X1 U1071 ( .A(n980), .B(KEYINPUT121), .Z(n982) );
  XNOR2_X1 U1072 ( .A(G299), .B(G1956), .ZN(n981) );
  NOR2_X1 U1073 ( .A1(n982), .A2(n981), .ZN(n983) );
  NAND2_X1 U1074 ( .A1(n984), .A2(n983), .ZN(n985) );
  NOR2_X1 U1075 ( .A1(n986), .A2(n985), .ZN(n987) );
  XNOR2_X1 U1076 ( .A(KEYINPUT122), .B(n987), .ZN(n990) );
  XOR2_X1 U1077 ( .A(G301), .B(G1961), .Z(n988) );
  XNOR2_X1 U1078 ( .A(n988), .B(KEYINPUT120), .ZN(n989) );
  NAND2_X1 U1079 ( .A1(n990), .A2(n989), .ZN(n993) );
  XOR2_X1 U1080 ( .A(G1348), .B(n991), .Z(n992) );
  NOR2_X1 U1081 ( .A1(n993), .A2(n992), .ZN(n994) );
  XNOR2_X1 U1082 ( .A(KEYINPUT123), .B(n994), .ZN(n995) );
  NOR2_X1 U1083 ( .A1(n996), .A2(n995), .ZN(n997) );
  NAND2_X1 U1084 ( .A1(n998), .A2(n997), .ZN(n999) );
  NAND2_X1 U1085 ( .A1(n1000), .A2(n999), .ZN(n1027) );
  XNOR2_X1 U1086 ( .A(G1971), .B(G22), .ZN(n1002) );
  XNOR2_X1 U1087 ( .A(G23), .B(G1976), .ZN(n1001) );
  NOR2_X1 U1088 ( .A1(n1002), .A2(n1001), .ZN(n1004) );
  XOR2_X1 U1089 ( .A(G1986), .B(G24), .Z(n1003) );
  NAND2_X1 U1090 ( .A1(n1004), .A2(n1003), .ZN(n1006) );
  XOR2_X1 U1091 ( .A(KEYINPUT126), .B(KEYINPUT58), .Z(n1005) );
  XNOR2_X1 U1092 ( .A(n1006), .B(n1005), .ZN(n1020) );
  XOR2_X1 U1093 ( .A(KEYINPUT124), .B(G4), .Z(n1008) );
  XNOR2_X1 U1094 ( .A(G1348), .B(KEYINPUT59), .ZN(n1007) );
  XNOR2_X1 U1095 ( .A(n1008), .B(n1007), .ZN(n1014) );
  XOR2_X1 U1096 ( .A(G20), .B(G1956), .Z(n1012) );
  XNOR2_X1 U1097 ( .A(G1341), .B(G19), .ZN(n1010) );
  XNOR2_X1 U1098 ( .A(G6), .B(G1981), .ZN(n1009) );
  NOR2_X1 U1099 ( .A1(n1010), .A2(n1009), .ZN(n1011) );
  NAND2_X1 U1100 ( .A1(n1012), .A2(n1011), .ZN(n1013) );
  NOR2_X1 U1101 ( .A1(n1014), .A2(n1013), .ZN(n1015) );
  XOR2_X1 U1102 ( .A(KEYINPUT60), .B(n1015), .Z(n1016) );
  XOR2_X1 U1103 ( .A(KEYINPUT125), .B(n1016), .Z(n1018) );
  XNOR2_X1 U1104 ( .A(G1966), .B(G21), .ZN(n1017) );
  NOR2_X1 U1105 ( .A1(n1018), .A2(n1017), .ZN(n1019) );
  NAND2_X1 U1106 ( .A1(n1020), .A2(n1019), .ZN(n1022) );
  XNOR2_X1 U1107 ( .A(G5), .B(G1961), .ZN(n1021) );
  NOR2_X1 U1108 ( .A1(n1022), .A2(n1021), .ZN(n1023) );
  XNOR2_X1 U1109 ( .A(KEYINPUT61), .B(n1023), .ZN(n1024) );
  NAND2_X1 U1110 ( .A1(n1025), .A2(n1024), .ZN(n1026) );
  NAND2_X1 U1111 ( .A1(n1027), .A2(n1026), .ZN(n1028) );
  NOR2_X1 U1112 ( .A1(n1029), .A2(n1028), .ZN(n1030) );
  NAND2_X1 U1113 ( .A1(n1031), .A2(n1030), .ZN(n1032) );
  XNOR2_X1 U1114 ( .A(n1032), .B(KEYINPUT62), .ZN(n1033) );
  XOR2_X1 U1115 ( .A(KEYINPUT127), .B(n1033), .Z(G150) );
  INV_X1 U1116 ( .A(G150), .ZN(G311) );
endmodule

