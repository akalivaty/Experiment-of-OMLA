//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 1 0 0 0 0 1 1 0 1 1 0 1 0 0 0 1 1 0 0 1 0 0 1 0 1 1 0 0 1 0 0 1 0 0 1 0 1 1 1 0 1 0 0 1 0 0 1 1 1 0 0 1 0 0 0 0 0 0 0 1 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:40:24 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n209, new_n210, new_n211, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n236, new_n237,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n244, new_n245,
    new_n246, new_n248, new_n249, new_n250, new_n251, new_n252, new_n253,
    new_n254, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n605,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n812, new_n813,
    new_n814, new_n815, new_n816, new_n817, new_n818, new_n819, new_n820,
    new_n821, new_n822, new_n823, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n883, new_n884,
    new_n885, new_n886, new_n887, new_n888, new_n889, new_n890, new_n891,
    new_n892, new_n893, new_n894, new_n895, new_n896, new_n897, new_n898,
    new_n899, new_n900, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n946, new_n947, new_n948,
    new_n949, new_n950, new_n951, new_n952, new_n953, new_n954, new_n955,
    new_n956, new_n957, new_n958, new_n959, new_n960, new_n961, new_n962,
    new_n963, new_n964, new_n965, new_n966, new_n967, new_n968, new_n969,
    new_n970, new_n971, new_n972, new_n973, new_n974, new_n975, new_n976,
    new_n977, new_n979, new_n980, new_n981, new_n982, new_n983, new_n984,
    new_n985, new_n986, new_n987, new_n988, new_n989, new_n990, new_n991,
    new_n992, new_n993, new_n994, new_n995, new_n996, new_n997, new_n998,
    new_n999, new_n1000, new_n1001, new_n1002, new_n1003, new_n1005,
    new_n1006, new_n1007, new_n1008, new_n1009, new_n1010, new_n1011,
    new_n1012, new_n1013, new_n1014, new_n1015, new_n1016, new_n1017,
    new_n1018, new_n1019, new_n1020, new_n1021, new_n1022, new_n1023,
    new_n1024, new_n1025, new_n1026, new_n1027, new_n1028, new_n1029,
    new_n1030, new_n1031, new_n1032, new_n1033, new_n1034, new_n1035,
    new_n1036, new_n1037, new_n1038, new_n1039, new_n1040, new_n1041,
    new_n1042, new_n1043, new_n1044, new_n1045, new_n1046, new_n1047,
    new_n1048, new_n1049, new_n1050, new_n1051, new_n1052, new_n1053,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1079, new_n1080, new_n1081, new_n1082, new_n1083, new_n1084,
    new_n1085, new_n1086, new_n1087, new_n1088, new_n1089, new_n1090,
    new_n1091, new_n1092, new_n1093, new_n1094, new_n1095, new_n1096,
    new_n1097, new_n1098, new_n1099, new_n1100, new_n1101, new_n1102,
    new_n1103, new_n1104, new_n1105, new_n1106, new_n1107, new_n1108,
    new_n1109, new_n1110, new_n1111, new_n1112, new_n1113, new_n1114,
    new_n1115, new_n1116, new_n1117, new_n1118, new_n1119, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1160, new_n1161, new_n1162, new_n1163,
    new_n1164, new_n1165, new_n1166, new_n1167, new_n1168, new_n1169,
    new_n1170, new_n1171, new_n1172, new_n1173, new_n1174, new_n1175,
    new_n1176, new_n1177, new_n1178, new_n1179, new_n1180, new_n1181,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1189,
    new_n1191, new_n1192, new_n1193, new_n1194, new_n1195, new_n1196,
    new_n1197, new_n1198, new_n1199, new_n1200, new_n1201, new_n1202,
    new_n1203, new_n1204, new_n1205, new_n1206, new_n1207, new_n1208,
    new_n1209, new_n1210, new_n1211, new_n1212, new_n1213, new_n1214,
    new_n1215, new_n1216, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1239,
    new_n1240, new_n1241, new_n1242, new_n1243, new_n1244, new_n1245,
    new_n1246;
  XNOR2_X1  g0000(.A(KEYINPUT64), .B(G50), .ZN(new_n201));
  INV_X1    g0001(.A(G58), .ZN(new_n202));
  INV_X1    g0002(.A(G68), .ZN(new_n203));
  NAND2_X1  g0003(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  NOR2_X1   g0004(.A1(new_n201), .A2(new_n204), .ZN(new_n205));
  INV_X1    g0005(.A(G77), .ZN(new_n206));
  NAND2_X1  g0006(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  XOR2_X1   g0007(.A(new_n207), .B(KEYINPUT65), .Z(G353));
  NOR2_X1   g0008(.A1(G97), .A2(G107), .ZN(new_n209));
  INV_X1    g0009(.A(new_n209), .ZN(new_n210));
  NAND2_X1  g0010(.A1(new_n210), .A2(G87), .ZN(new_n211));
  XNOR2_X1  g0011(.A(new_n211), .B(KEYINPUT66), .ZN(G355));
  INV_X1    g0012(.A(G244), .ZN(new_n213));
  NOR2_X1   g0013(.A1(new_n206), .A2(new_n213), .ZN(new_n214));
  AOI22_X1  g0014(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n215));
  INV_X1    g0015(.A(G238), .ZN(new_n216));
  INV_X1    g0016(.A(G107), .ZN(new_n217));
  INV_X1    g0017(.A(G264), .ZN(new_n218));
  OAI221_X1 g0018(.A(new_n215), .B1(new_n203), .B2(new_n216), .C1(new_n217), .C2(new_n218), .ZN(new_n219));
  AOI211_X1 g0019(.A(new_n214), .B(new_n219), .C1(G116), .C2(G270), .ZN(new_n220));
  NAND2_X1  g0020(.A1(G50), .A2(G226), .ZN(new_n221));
  INV_X1    g0021(.A(G232), .ZN(new_n222));
  OAI211_X1 g0022(.A(new_n220), .B(new_n221), .C1(new_n202), .C2(new_n222), .ZN(new_n223));
  INV_X1    g0023(.A(G1), .ZN(new_n224));
  INV_X1    g0024(.A(G20), .ZN(new_n225));
  NOR2_X1   g0025(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  INV_X1    g0026(.A(new_n226), .ZN(new_n227));
  NAND2_X1  g0027(.A1(KEYINPUT67), .A2(KEYINPUT1), .ZN(new_n228));
  NAND3_X1  g0028(.A1(new_n223), .A2(new_n227), .A3(new_n228), .ZN(new_n229));
  NOR2_X1   g0029(.A1(KEYINPUT67), .A2(KEYINPUT1), .ZN(new_n230));
  XOR2_X1   g0030(.A(new_n229), .B(new_n230), .Z(new_n231));
  NAND2_X1  g0031(.A1(new_n204), .A2(G50), .ZN(new_n232));
  NAND2_X1  g0032(.A1(G1), .A2(G13), .ZN(new_n233));
  NOR3_X1   g0033(.A1(new_n232), .A2(new_n225), .A3(new_n233), .ZN(new_n234));
  NOR2_X1   g0034(.A1(new_n227), .A2(G13), .ZN(new_n235));
  OAI211_X1 g0035(.A(new_n235), .B(G250), .C1(G257), .C2(G264), .ZN(new_n236));
  XOR2_X1   g0036(.A(new_n236), .B(KEYINPUT0), .Z(new_n237));
  NOR3_X1   g0037(.A1(new_n231), .A2(new_n234), .A3(new_n237), .ZN(G361));
  XOR2_X1   g0038(.A(G238), .B(G244), .Z(new_n239));
  XNOR2_X1  g0039(.A(KEYINPUT68), .B(KEYINPUT2), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XNOR2_X1  g0041(.A(G226), .B(G232), .ZN(new_n242));
  XOR2_X1   g0042(.A(new_n241), .B(new_n242), .Z(new_n243));
  XNOR2_X1  g0043(.A(G250), .B(G257), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n244), .B(new_n218), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n245), .B(G270), .ZN(new_n246));
  XOR2_X1   g0046(.A(new_n243), .B(new_n246), .Z(G358));
  XNOR2_X1  g0047(.A(G68), .B(G77), .ZN(new_n248));
  INV_X1    g0048(.A(G50), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n248), .B(new_n249), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n250), .B(G58), .ZN(new_n251));
  XOR2_X1   g0051(.A(G97), .B(G107), .Z(new_n252));
  XNOR2_X1  g0052(.A(G87), .B(G116), .ZN(new_n253));
  XNOR2_X1  g0053(.A(new_n252), .B(new_n253), .ZN(new_n254));
  XNOR2_X1  g0054(.A(new_n251), .B(new_n254), .ZN(G351));
  AOI21_X1  g0055(.A(new_n233), .B1(G33), .B2(G41), .ZN(new_n256));
  INV_X1    g0056(.A(new_n256), .ZN(new_n257));
  OAI21_X1  g0057(.A(new_n224), .B1(G41), .B2(G45), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  INV_X1    g0059(.A(new_n259), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n260), .A2(G226), .ZN(new_n261));
  INV_X1    g0061(.A(G274), .ZN(new_n262));
  INV_X1    g0062(.A(KEYINPUT69), .ZN(new_n263));
  INV_X1    g0063(.A(G41), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  NAND2_X1  g0065(.A1(KEYINPUT69), .A2(G41), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n265), .A2(new_n266), .ZN(new_n267));
  INV_X1    g0067(.A(G45), .ZN(new_n268));
  AOI211_X1 g0068(.A(G1), .B(new_n262), .C1(new_n267), .C2(new_n268), .ZN(new_n269));
  INV_X1    g0069(.A(new_n269), .ZN(new_n270));
  XNOR2_X1  g0070(.A(KEYINPUT3), .B(G33), .ZN(new_n271));
  INV_X1    g0071(.A(G1698), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n272), .A2(G222), .ZN(new_n273));
  NAND2_X1  g0073(.A1(G223), .A2(G1698), .ZN(new_n274));
  NAND3_X1  g0074(.A1(new_n271), .A2(new_n273), .A3(new_n274), .ZN(new_n275));
  OAI211_X1 g0075(.A(new_n275), .B(new_n256), .C1(G77), .C2(new_n271), .ZN(new_n276));
  NAND3_X1  g0076(.A1(new_n261), .A2(new_n270), .A3(new_n276), .ZN(new_n277));
  INV_X1    g0077(.A(new_n277), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n278), .A2(G190), .ZN(new_n279));
  AOI21_X1  g0079(.A(KEYINPUT73), .B1(new_n277), .B2(G200), .ZN(new_n280));
  XOR2_X1   g0080(.A(KEYINPUT8), .B(G58), .Z(new_n281));
  INV_X1    g0081(.A(G33), .ZN(new_n282));
  NOR2_X1   g0082(.A1(new_n282), .A2(G20), .ZN(new_n283));
  NOR2_X1   g0083(.A1(G20), .A2(G33), .ZN(new_n284));
  AOI22_X1  g0084(.A1(new_n281), .A2(new_n283), .B1(G150), .B2(new_n284), .ZN(new_n285));
  OAI21_X1  g0085(.A(new_n285), .B1(new_n225), .B2(new_n205), .ZN(new_n286));
  NAND3_X1  g0086(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n287), .A2(new_n233), .ZN(new_n288));
  AOI21_X1  g0088(.A(new_n288), .B1(new_n224), .B2(G20), .ZN(new_n289));
  AOI22_X1  g0089(.A1(new_n286), .A2(new_n288), .B1(G50), .B2(new_n289), .ZN(new_n290));
  NAND3_X1  g0090(.A1(new_n224), .A2(G13), .A3(G20), .ZN(new_n291));
  OAI21_X1  g0091(.A(new_n290), .B1(G50), .B2(new_n291), .ZN(new_n292));
  INV_X1    g0092(.A(KEYINPUT72), .ZN(new_n293));
  INV_X1    g0093(.A(KEYINPUT9), .ZN(new_n294));
  NAND3_X1  g0094(.A1(new_n292), .A2(new_n293), .A3(new_n294), .ZN(new_n295));
  INV_X1    g0095(.A(new_n295), .ZN(new_n296));
  AOI21_X1  g0096(.A(new_n293), .B1(new_n292), .B2(new_n294), .ZN(new_n297));
  OAI211_X1 g0097(.A(new_n279), .B(new_n280), .C1(new_n296), .C2(new_n297), .ZN(new_n298));
  NOR2_X1   g0098(.A1(new_n292), .A2(new_n294), .ZN(new_n299));
  OAI21_X1  g0099(.A(KEYINPUT10), .B1(new_n298), .B2(new_n299), .ZN(new_n300));
  INV_X1    g0100(.A(new_n280), .ZN(new_n301));
  INV_X1    g0101(.A(new_n297), .ZN(new_n302));
  AOI21_X1  g0102(.A(new_n301), .B1(new_n302), .B2(new_n295), .ZN(new_n303));
  INV_X1    g0103(.A(KEYINPUT10), .ZN(new_n304));
  INV_X1    g0104(.A(new_n299), .ZN(new_n305));
  NAND4_X1  g0105(.A1(new_n303), .A2(new_n304), .A3(new_n305), .A4(new_n279), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n300), .A2(new_n306), .ZN(new_n307));
  INV_X1    g0107(.A(G179), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n278), .A2(new_n308), .ZN(new_n309));
  INV_X1    g0109(.A(G169), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n277), .A2(new_n310), .ZN(new_n311));
  NAND3_X1  g0111(.A1(new_n309), .A2(new_n292), .A3(new_n311), .ZN(new_n312));
  AND2_X1   g0112(.A1(KEYINPUT75), .A2(KEYINPUT14), .ZN(new_n313));
  INV_X1    g0113(.A(KEYINPUT13), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n222), .A2(G1698), .ZN(new_n315));
  OAI211_X1 g0115(.A(new_n271), .B(new_n315), .C1(G226), .C2(G1698), .ZN(new_n316));
  NAND2_X1  g0116(.A1(G33), .A2(G97), .ZN(new_n317));
  AOI21_X1  g0117(.A(new_n257), .B1(new_n316), .B2(new_n317), .ZN(new_n318));
  NOR2_X1   g0118(.A1(new_n318), .A2(new_n269), .ZN(new_n319));
  NOR2_X1   g0119(.A1(new_n259), .A2(new_n216), .ZN(new_n320));
  INV_X1    g0120(.A(new_n320), .ZN(new_n321));
  AOI21_X1  g0121(.A(new_n314), .B1(new_n319), .B2(new_n321), .ZN(new_n322));
  NOR4_X1   g0122(.A1(new_n318), .A2(new_n320), .A3(KEYINPUT13), .A4(new_n269), .ZN(new_n323));
  NOR2_X1   g0123(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  OAI21_X1  g0124(.A(new_n313), .B1(new_n324), .B2(new_n310), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n324), .A2(G179), .ZN(new_n326));
  NAND2_X1  g0126(.A1(KEYINPUT75), .A2(KEYINPUT14), .ZN(new_n327));
  OAI211_X1 g0127(.A(G169), .B(new_n327), .C1(new_n322), .C2(new_n323), .ZN(new_n328));
  NAND3_X1  g0128(.A1(new_n325), .A2(new_n326), .A3(new_n328), .ZN(new_n329));
  INV_X1    g0129(.A(new_n288), .ZN(new_n330));
  AOI22_X1  g0130(.A1(new_n283), .A2(G77), .B1(G20), .B2(new_n203), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n284), .A2(G50), .ZN(new_n332));
  AOI21_X1  g0132(.A(new_n330), .B1(new_n331), .B2(new_n332), .ZN(new_n333));
  XOR2_X1   g0133(.A(new_n333), .B(KEYINPUT11), .Z(new_n334));
  NAND2_X1  g0134(.A1(new_n289), .A2(G68), .ZN(new_n335));
  OAI21_X1  g0135(.A(KEYINPUT74), .B1(new_n291), .B2(G68), .ZN(new_n336));
  XOR2_X1   g0136(.A(new_n336), .B(KEYINPUT12), .Z(new_n337));
  NAND3_X1  g0137(.A1(new_n334), .A2(new_n335), .A3(new_n337), .ZN(new_n338));
  OAI21_X1  g0138(.A(G200), .B1(new_n322), .B2(new_n323), .ZN(new_n339));
  AOI21_X1  g0139(.A(new_n338), .B1(new_n324), .B2(G190), .ZN(new_n340));
  AOI22_X1  g0140(.A1(new_n329), .A2(new_n338), .B1(new_n339), .B2(new_n340), .ZN(new_n341));
  XNOR2_X1  g0141(.A(KEYINPUT8), .B(G58), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n225), .A2(new_n282), .ZN(new_n343));
  OAI22_X1  g0143(.A1(new_n342), .A2(new_n343), .B1(new_n225), .B2(new_n206), .ZN(new_n344));
  XNOR2_X1  g0144(.A(new_n344), .B(KEYINPUT70), .ZN(new_n345));
  INV_X1    g0145(.A(new_n283), .ZN(new_n346));
  XNOR2_X1  g0146(.A(KEYINPUT15), .B(G87), .ZN(new_n347));
  OR2_X1    g0147(.A1(new_n347), .A2(KEYINPUT71), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n347), .A2(KEYINPUT71), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n348), .A2(new_n349), .ZN(new_n350));
  OAI21_X1  g0150(.A(new_n345), .B1(new_n346), .B2(new_n350), .ZN(new_n351));
  INV_X1    g0151(.A(new_n291), .ZN(new_n352));
  AOI22_X1  g0152(.A1(new_n351), .A2(new_n288), .B1(new_n206), .B2(new_n352), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n289), .A2(G77), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  INV_X1    g0155(.A(new_n355), .ZN(new_n356));
  NAND2_X1  g0156(.A1(G238), .A2(G1698), .ZN(new_n357));
  OAI211_X1 g0157(.A(new_n271), .B(new_n357), .C1(new_n222), .C2(G1698), .ZN(new_n358));
  OAI211_X1 g0158(.A(new_n358), .B(new_n256), .C1(G107), .C2(new_n271), .ZN(new_n359));
  OAI211_X1 g0159(.A(new_n359), .B(new_n270), .C1(new_n213), .C2(new_n259), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n360), .A2(G200), .ZN(new_n361));
  INV_X1    g0161(.A(G190), .ZN(new_n362));
  OAI211_X1 g0162(.A(new_n356), .B(new_n361), .C1(new_n362), .C2(new_n360), .ZN(new_n363));
  AND4_X1   g0163(.A1(new_n307), .A2(new_n312), .A3(new_n341), .A4(new_n363), .ZN(new_n364));
  INV_X1    g0164(.A(KEYINPUT7), .ZN(new_n365));
  OAI21_X1  g0165(.A(new_n365), .B1(new_n271), .B2(G20), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n225), .A2(KEYINPUT7), .ZN(new_n367));
  OAI21_X1  g0167(.A(KEYINPUT76), .B1(new_n271), .B2(new_n367), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n282), .A2(KEYINPUT3), .ZN(new_n369));
  INV_X1    g0169(.A(KEYINPUT3), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n370), .A2(G33), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n369), .A2(new_n371), .ZN(new_n372));
  INV_X1    g0172(.A(KEYINPUT76), .ZN(new_n373));
  INV_X1    g0173(.A(new_n367), .ZN(new_n374));
  NAND3_X1  g0174(.A1(new_n372), .A2(new_n373), .A3(new_n374), .ZN(new_n375));
  NAND3_X1  g0175(.A1(new_n366), .A2(new_n368), .A3(new_n375), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n376), .A2(G68), .ZN(new_n377));
  NAND2_X1  g0177(.A1(G58), .A2(G68), .ZN(new_n378));
  AOI21_X1  g0178(.A(new_n225), .B1(new_n204), .B2(new_n378), .ZN(new_n379));
  INV_X1    g0179(.A(G159), .ZN(new_n380));
  NOR2_X1   g0180(.A1(new_n343), .A2(new_n380), .ZN(new_n381));
  OAI21_X1  g0181(.A(KEYINPUT77), .B1(new_n379), .B2(new_n381), .ZN(new_n382));
  INV_X1    g0182(.A(new_n378), .ZN(new_n383));
  NOR2_X1   g0183(.A1(G58), .A2(G68), .ZN(new_n384));
  OAI21_X1  g0184(.A(G20), .B1(new_n383), .B2(new_n384), .ZN(new_n385));
  INV_X1    g0185(.A(KEYINPUT77), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n284), .A2(G159), .ZN(new_n387));
  NAND3_X1  g0187(.A1(new_n385), .A2(new_n386), .A3(new_n387), .ZN(new_n388));
  AND2_X1   g0188(.A1(new_n382), .A2(new_n388), .ZN(new_n389));
  NAND3_X1  g0189(.A1(new_n377), .A2(KEYINPUT16), .A3(new_n389), .ZN(new_n390));
  INV_X1    g0190(.A(KEYINPUT16), .ZN(new_n391));
  OAI21_X1  g0191(.A(KEYINPUT78), .B1(new_n282), .B2(KEYINPUT3), .ZN(new_n392));
  INV_X1    g0192(.A(KEYINPUT78), .ZN(new_n393));
  NAND3_X1  g0193(.A1(new_n393), .A2(new_n370), .A3(G33), .ZN(new_n394));
  NAND3_X1  g0194(.A1(new_n392), .A2(new_n394), .A3(new_n369), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n395), .A2(new_n374), .ZN(new_n396));
  AOI21_X1  g0196(.A(new_n203), .B1(new_n396), .B2(new_n366), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n382), .A2(new_n388), .ZN(new_n398));
  OAI21_X1  g0198(.A(new_n391), .B1(new_n397), .B2(new_n398), .ZN(new_n399));
  NAND3_X1  g0199(.A1(new_n390), .A2(new_n288), .A3(new_n399), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n400), .A2(KEYINPUT79), .ZN(new_n401));
  NOR2_X1   g0201(.A1(new_n281), .A2(new_n291), .ZN(new_n402));
  AOI21_X1  g0202(.A(new_n402), .B1(new_n289), .B2(new_n281), .ZN(new_n403));
  INV_X1    g0203(.A(KEYINPUT79), .ZN(new_n404));
  NAND4_X1  g0204(.A1(new_n390), .A2(new_n399), .A3(new_n404), .A4(new_n288), .ZN(new_n405));
  AND3_X1   g0205(.A1(new_n401), .A2(new_n403), .A3(new_n405), .ZN(new_n406));
  OAI21_X1  g0206(.A(new_n271), .B1(G226), .B2(new_n272), .ZN(new_n407));
  NOR2_X1   g0207(.A1(G223), .A2(G1698), .ZN(new_n408));
  INV_X1    g0208(.A(G87), .ZN(new_n409));
  OAI22_X1  g0209(.A1(new_n407), .A2(new_n408), .B1(new_n282), .B2(new_n409), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n410), .A2(new_n256), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n260), .A2(G232), .ZN(new_n412));
  NAND3_X1  g0212(.A1(new_n411), .A2(new_n270), .A3(new_n412), .ZN(new_n413));
  INV_X1    g0213(.A(new_n413), .ZN(new_n414));
  INV_X1    g0214(.A(G200), .ZN(new_n415));
  NOR2_X1   g0215(.A1(new_n414), .A2(new_n415), .ZN(new_n416));
  INV_X1    g0216(.A(new_n416), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n414), .A2(G190), .ZN(new_n418));
  NAND4_X1  g0218(.A1(new_n406), .A2(KEYINPUT17), .A3(new_n417), .A4(new_n418), .ZN(new_n419));
  INV_X1    g0219(.A(KEYINPUT17), .ZN(new_n420));
  NAND4_X1  g0220(.A1(new_n401), .A2(new_n418), .A3(new_n403), .A4(new_n405), .ZN(new_n421));
  OAI21_X1  g0221(.A(new_n420), .B1(new_n421), .B2(new_n416), .ZN(new_n422));
  AND2_X1   g0222(.A1(new_n419), .A2(new_n422), .ZN(new_n423));
  NAND3_X1  g0223(.A1(new_n401), .A2(new_n403), .A3(new_n405), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n414), .A2(G179), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n413), .A2(G169), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n425), .A2(new_n426), .ZN(new_n427));
  AND3_X1   g0227(.A1(new_n424), .A2(KEYINPUT18), .A3(new_n427), .ZN(new_n428));
  AOI21_X1  g0228(.A(KEYINPUT18), .B1(new_n424), .B2(new_n427), .ZN(new_n429));
  OR2_X1    g0229(.A1(new_n428), .A2(new_n429), .ZN(new_n430));
  NOR2_X1   g0230(.A1(new_n360), .A2(G179), .ZN(new_n431));
  AOI21_X1  g0231(.A(new_n431), .B1(new_n310), .B2(new_n360), .ZN(new_n432));
  AND2_X1   g0232(.A1(new_n355), .A2(new_n432), .ZN(new_n433));
  INV_X1    g0233(.A(new_n433), .ZN(new_n434));
  AND4_X1   g0234(.A1(new_n364), .A2(new_n423), .A3(new_n430), .A4(new_n434), .ZN(new_n435));
  INV_X1    g0235(.A(new_n435), .ZN(new_n436));
  INV_X1    g0236(.A(KEYINPUT19), .ZN(new_n437));
  INV_X1    g0237(.A(G97), .ZN(new_n438));
  OAI21_X1  g0238(.A(new_n437), .B1(new_n346), .B2(new_n438), .ZN(new_n439));
  NAND3_X1  g0239(.A1(new_n271), .A2(new_n225), .A3(G68), .ZN(new_n440));
  XOR2_X1   g0240(.A(KEYINPUT84), .B(G87), .Z(new_n441));
  NOR2_X1   g0241(.A1(new_n441), .A2(new_n210), .ZN(new_n442));
  NOR2_X1   g0242(.A1(new_n317), .A2(new_n437), .ZN(new_n443));
  NOR2_X1   g0243(.A1(new_n443), .A2(G20), .ZN(new_n444));
  OAI211_X1 g0244(.A(new_n439), .B(new_n440), .C1(new_n442), .C2(new_n444), .ZN(new_n445));
  AOI22_X1  g0245(.A1(new_n445), .A2(new_n288), .B1(new_n352), .B2(new_n350), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n224), .A2(G33), .ZN(new_n447));
  NAND3_X1  g0247(.A1(new_n330), .A2(new_n291), .A3(new_n447), .ZN(new_n448));
  OR2_X1    g0248(.A1(new_n350), .A2(new_n448), .ZN(new_n449));
  INV_X1    g0249(.A(G250), .ZN(new_n450));
  OAI21_X1  g0250(.A(new_n450), .B1(new_n268), .B2(G1), .ZN(new_n451));
  NOR2_X1   g0251(.A1(new_n268), .A2(G1), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n452), .A2(new_n262), .ZN(new_n453));
  NAND3_X1  g0253(.A1(new_n257), .A2(new_n451), .A3(new_n453), .ZN(new_n454));
  INV_X1    g0254(.A(G116), .ZN(new_n455));
  NOR2_X1   g0255(.A1(new_n282), .A2(new_n455), .ZN(new_n456));
  NOR2_X1   g0256(.A1(G238), .A2(G1698), .ZN(new_n457));
  AOI21_X1  g0257(.A(new_n457), .B1(new_n213), .B2(G1698), .ZN(new_n458));
  AOI21_X1  g0258(.A(new_n456), .B1(new_n458), .B2(new_n271), .ZN(new_n459));
  OAI21_X1  g0259(.A(new_n454), .B1(new_n459), .B2(new_n257), .ZN(new_n460));
  AOI22_X1  g0260(.A1(new_n446), .A2(new_n449), .B1(new_n460), .B2(new_n310), .ZN(new_n461));
  OAI211_X1 g0261(.A(new_n454), .B(new_n308), .C1(new_n459), .C2(new_n257), .ZN(new_n462));
  INV_X1    g0262(.A(KEYINPUT83), .ZN(new_n463));
  XNOR2_X1  g0263(.A(new_n462), .B(new_n463), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n461), .A2(new_n464), .ZN(new_n465));
  OAI211_X1 g0265(.A(new_n454), .B(G190), .C1(new_n459), .C2(new_n257), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n445), .A2(new_n288), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n350), .A2(new_n352), .ZN(new_n468));
  OAI21_X1  g0268(.A(KEYINPUT85), .B1(new_n448), .B2(new_n409), .ZN(new_n469));
  AOI21_X1  g0269(.A(new_n288), .B1(new_n224), .B2(G33), .ZN(new_n470));
  INV_X1    g0270(.A(KEYINPUT85), .ZN(new_n471));
  NAND4_X1  g0271(.A1(new_n470), .A2(new_n471), .A3(G87), .A4(new_n291), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n469), .A2(new_n472), .ZN(new_n473));
  AND4_X1   g0273(.A1(new_n466), .A2(new_n467), .A3(new_n468), .A4(new_n473), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n460), .A2(G200), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n465), .A2(new_n476), .ZN(new_n477));
  INV_X1    g0277(.A(KEYINPUT20), .ZN(new_n478));
  OAI21_X1  g0278(.A(new_n225), .B1(new_n438), .B2(G33), .ZN(new_n479));
  INV_X1    g0279(.A(KEYINPUT81), .ZN(new_n480));
  NAND3_X1  g0280(.A1(new_n480), .A2(G33), .A3(G283), .ZN(new_n481));
  NAND2_X1  g0281(.A1(G33), .A2(G283), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n482), .A2(KEYINPUT81), .ZN(new_n483));
  AOI21_X1  g0283(.A(new_n479), .B1(new_n481), .B2(new_n483), .ZN(new_n484));
  AOI22_X1  g0284(.A1(new_n287), .A2(new_n233), .B1(G20), .B2(new_n455), .ZN(new_n485));
  INV_X1    g0285(.A(new_n485), .ZN(new_n486));
  OAI21_X1  g0286(.A(new_n478), .B1(new_n484), .B2(new_n486), .ZN(new_n487));
  AND2_X1   g0287(.A1(new_n483), .A2(new_n481), .ZN(new_n488));
  OAI211_X1 g0288(.A(KEYINPUT20), .B(new_n485), .C1(new_n488), .C2(new_n479), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n487), .A2(new_n489), .ZN(new_n490));
  NAND3_X1  g0290(.A1(new_n470), .A2(G116), .A3(new_n291), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n352), .A2(new_n455), .ZN(new_n492));
  NAND3_X1  g0292(.A1(new_n490), .A2(new_n491), .A3(new_n492), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n272), .A2(G257), .ZN(new_n494));
  OAI211_X1 g0294(.A(new_n271), .B(new_n494), .C1(new_n218), .C2(new_n272), .ZN(new_n495));
  OAI211_X1 g0295(.A(new_n495), .B(new_n256), .C1(G303), .C2(new_n271), .ZN(new_n496));
  INV_X1    g0296(.A(KEYINPUT5), .ZN(new_n497));
  NAND3_X1  g0297(.A1(new_n265), .A2(new_n497), .A3(new_n266), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n264), .A2(KEYINPUT5), .ZN(new_n499));
  NAND3_X1  g0299(.A1(new_n498), .A2(new_n499), .A3(new_n452), .ZN(new_n500));
  NAND3_X1  g0300(.A1(new_n500), .A2(G270), .A3(new_n257), .ZN(new_n501));
  NAND4_X1  g0301(.A1(new_n498), .A2(G274), .A3(new_n499), .A4(new_n452), .ZN(new_n502));
  NAND3_X1  g0302(.A1(new_n496), .A2(new_n501), .A3(new_n502), .ZN(new_n503));
  NAND3_X1  g0303(.A1(new_n493), .A2(G169), .A3(new_n503), .ZN(new_n504));
  INV_X1    g0304(.A(KEYINPUT21), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  INV_X1    g0306(.A(new_n493), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n503), .A2(G200), .ZN(new_n508));
  NAND4_X1  g0308(.A1(new_n496), .A2(new_n501), .A3(G190), .A4(new_n502), .ZN(new_n509));
  NAND3_X1  g0309(.A1(new_n507), .A2(new_n508), .A3(new_n509), .ZN(new_n510));
  NOR2_X1   g0310(.A1(new_n503), .A2(new_n308), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n511), .A2(new_n493), .ZN(new_n512));
  NAND4_X1  g0312(.A1(new_n493), .A2(KEYINPUT21), .A3(new_n503), .A4(G169), .ZN(new_n513));
  NAND4_X1  g0313(.A1(new_n506), .A2(new_n510), .A3(new_n512), .A4(new_n513), .ZN(new_n514));
  NOR2_X1   g0314(.A1(new_n477), .A2(new_n514), .ZN(new_n515));
  NAND3_X1  g0315(.A1(new_n500), .A2(G257), .A3(new_n257), .ZN(new_n516));
  AND2_X1   g0316(.A1(new_n516), .A2(new_n502), .ZN(new_n517));
  AND2_X1   g0317(.A1(G250), .A2(G1698), .ZN(new_n518));
  AND3_X1   g0318(.A1(new_n369), .A2(new_n371), .A3(new_n518), .ZN(new_n519));
  NAND4_X1  g0319(.A1(new_n369), .A2(new_n371), .A3(G244), .A4(new_n272), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n520), .A2(KEYINPUT4), .ZN(new_n521));
  INV_X1    g0321(.A(KEYINPUT4), .ZN(new_n522));
  NAND4_X1  g0322(.A1(new_n271), .A2(new_n522), .A3(G244), .A4(new_n272), .ZN(new_n523));
  AOI211_X1 g0323(.A(new_n488), .B(new_n519), .C1(new_n521), .C2(new_n523), .ZN(new_n524));
  OAI211_X1 g0324(.A(new_n517), .B(G190), .C1(new_n257), .C2(new_n524), .ZN(new_n525));
  INV_X1    g0325(.A(KEYINPUT82), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  NOR2_X1   g0327(.A1(new_n291), .A2(G97), .ZN(new_n528));
  NOR2_X1   g0328(.A1(new_n448), .A2(new_n438), .ZN(new_n529));
  INV_X1    g0329(.A(KEYINPUT6), .ZN(new_n530));
  NOR2_X1   g0330(.A1(new_n438), .A2(new_n217), .ZN(new_n531));
  OAI21_X1  g0331(.A(new_n530), .B1(new_n531), .B2(new_n209), .ZN(new_n532));
  NAND3_X1  g0332(.A1(new_n217), .A2(KEYINPUT6), .A3(G97), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n534), .A2(G20), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n284), .A2(G77), .ZN(new_n536));
  XOR2_X1   g0336(.A(new_n536), .B(KEYINPUT80), .Z(new_n537));
  NOR2_X1   g0337(.A1(new_n370), .A2(G33), .ZN(new_n538));
  NOR2_X1   g0338(.A1(new_n282), .A2(KEYINPUT3), .ZN(new_n539));
  OAI21_X1  g0339(.A(new_n225), .B1(new_n538), .B2(new_n539), .ZN(new_n540));
  AOI22_X1  g0340(.A1(new_n365), .A2(new_n540), .B1(new_n395), .B2(new_n374), .ZN(new_n541));
  OAI211_X1 g0341(.A(new_n535), .B(new_n537), .C1(new_n541), .C2(new_n217), .ZN(new_n542));
  AOI211_X1 g0342(.A(new_n528), .B(new_n529), .C1(new_n542), .C2(new_n288), .ZN(new_n543));
  AOI21_X1  g0343(.A(new_n519), .B1(new_n521), .B2(new_n523), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n483), .A2(new_n481), .ZN(new_n545));
  AOI21_X1  g0345(.A(new_n257), .B1(new_n544), .B2(new_n545), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n516), .A2(new_n502), .ZN(new_n547));
  OAI21_X1  g0347(.A(G200), .B1(new_n546), .B2(new_n547), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n521), .A2(new_n523), .ZN(new_n549));
  INV_X1    g0349(.A(new_n519), .ZN(new_n550));
  NAND3_X1  g0350(.A1(new_n549), .A2(new_n545), .A3(new_n550), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n551), .A2(new_n256), .ZN(new_n552));
  NAND4_X1  g0352(.A1(new_n552), .A2(KEYINPUT82), .A3(G190), .A4(new_n517), .ZN(new_n553));
  NAND4_X1  g0353(.A1(new_n527), .A2(new_n543), .A3(new_n548), .A4(new_n553), .ZN(new_n554));
  AOI21_X1  g0354(.A(new_n528), .B1(new_n542), .B2(new_n288), .ZN(new_n555));
  INV_X1    g0355(.A(new_n529), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  OAI21_X1  g0357(.A(new_n310), .B1(new_n546), .B2(new_n547), .ZN(new_n558));
  NAND3_X1  g0358(.A1(new_n552), .A2(new_n308), .A3(new_n517), .ZN(new_n559));
  NAND3_X1  g0359(.A1(new_n557), .A2(new_n558), .A3(new_n559), .ZN(new_n560));
  AND2_X1   g0360(.A1(new_n554), .A2(new_n560), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n450), .A2(new_n272), .ZN(new_n562));
  OAI211_X1 g0362(.A(new_n271), .B(new_n562), .C1(G257), .C2(new_n272), .ZN(new_n563));
  NAND2_X1  g0363(.A1(G33), .A2(G294), .ZN(new_n564));
  AOI21_X1  g0364(.A(new_n257), .B1(new_n563), .B2(new_n564), .ZN(new_n565));
  NAND3_X1  g0365(.A1(new_n500), .A2(G264), .A3(new_n257), .ZN(new_n566));
  INV_X1    g0366(.A(KEYINPUT87), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  NAND4_X1  g0368(.A1(new_n500), .A2(KEYINPUT87), .A3(G264), .A4(new_n257), .ZN(new_n569));
  AOI21_X1  g0369(.A(new_n565), .B1(new_n568), .B2(new_n569), .ZN(new_n570));
  NAND3_X1  g0370(.A1(new_n570), .A2(new_n362), .A3(new_n502), .ZN(new_n571));
  INV_X1    g0371(.A(new_n502), .ZN(new_n572));
  AOI211_X1 g0372(.A(new_n572), .B(new_n565), .C1(new_n568), .C2(new_n569), .ZN(new_n573));
  OAI211_X1 g0373(.A(new_n571), .B(KEYINPUT88), .C1(new_n573), .C2(G200), .ZN(new_n574));
  NOR2_X1   g0374(.A1(new_n225), .A2(G107), .ZN(new_n575));
  NAND3_X1  g0375(.A1(new_n575), .A2(new_n224), .A3(G13), .ZN(new_n576));
  XOR2_X1   g0376(.A(new_n576), .B(KEYINPUT25), .Z(new_n577));
  OAI21_X1  g0377(.A(new_n577), .B1(new_n217), .B2(new_n448), .ZN(new_n578));
  NAND2_X1  g0378(.A1(KEYINPUT86), .A2(KEYINPUT24), .ZN(new_n579));
  NAND4_X1  g0379(.A1(new_n369), .A2(new_n371), .A3(new_n225), .A4(G87), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n580), .A2(KEYINPUT22), .ZN(new_n581));
  INV_X1    g0381(.A(KEYINPUT22), .ZN(new_n582));
  NAND4_X1  g0382(.A1(new_n271), .A2(new_n582), .A3(new_n225), .A4(G87), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n581), .A2(new_n583), .ZN(new_n584));
  XNOR2_X1  g0384(.A(new_n575), .B(KEYINPUT23), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n456), .A2(new_n225), .ZN(new_n586));
  NAND3_X1  g0386(.A1(new_n584), .A2(new_n585), .A3(new_n586), .ZN(new_n587));
  NOR2_X1   g0387(.A1(KEYINPUT86), .A2(KEYINPUT24), .ZN(new_n588));
  NOR2_X1   g0388(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  INV_X1    g0389(.A(new_n588), .ZN(new_n590));
  AOI22_X1  g0390(.A1(new_n581), .A2(new_n583), .B1(new_n225), .B2(new_n456), .ZN(new_n591));
  AOI21_X1  g0391(.A(new_n590), .B1(new_n591), .B2(new_n585), .ZN(new_n592));
  OAI21_X1  g0392(.A(new_n579), .B1(new_n589), .B2(new_n592), .ZN(new_n593));
  AOI21_X1  g0393(.A(new_n578), .B1(new_n593), .B2(new_n288), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n570), .A2(new_n502), .ZN(new_n595));
  INV_X1    g0395(.A(KEYINPUT88), .ZN(new_n596));
  NAND3_X1  g0396(.A1(new_n595), .A2(new_n596), .A3(new_n415), .ZN(new_n597));
  NAND3_X1  g0397(.A1(new_n574), .A2(new_n594), .A3(new_n597), .ZN(new_n598));
  NAND3_X1  g0398(.A1(new_n570), .A2(new_n308), .A3(new_n502), .ZN(new_n599));
  OAI21_X1  g0399(.A(new_n599), .B1(new_n573), .B2(G169), .ZN(new_n600));
  OR2_X1    g0400(.A1(new_n594), .A2(new_n600), .ZN(new_n601));
  NAND4_X1  g0401(.A1(new_n515), .A2(new_n561), .A3(new_n598), .A4(new_n601), .ZN(new_n602));
  NOR2_X1   g0402(.A1(new_n436), .A2(new_n602), .ZN(new_n603));
  XOR2_X1   g0403(.A(new_n603), .B(KEYINPUT89), .Z(G372));
  NAND2_X1  g0404(.A1(new_n329), .A2(new_n338), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n605), .A2(new_n434), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n340), .A2(new_n339), .ZN(new_n607));
  NAND4_X1  g0407(.A1(new_n606), .A2(new_n607), .A3(new_n422), .A4(new_n419), .ZN(new_n608));
  AND2_X1   g0408(.A1(new_n608), .A2(new_n430), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n609), .A2(KEYINPUT91), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n610), .A2(new_n307), .ZN(new_n611));
  NOR2_X1   g0411(.A1(new_n609), .A2(KEYINPUT91), .ZN(new_n612));
  OAI21_X1  g0412(.A(new_n312), .B1(new_n611), .B2(new_n612), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n613), .A2(KEYINPUT92), .ZN(new_n614));
  INV_X1    g0414(.A(KEYINPUT92), .ZN(new_n615));
  OAI211_X1 g0415(.A(new_n615), .B(new_n312), .C1(new_n611), .C2(new_n612), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n614), .A2(new_n616), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n461), .A2(new_n462), .ZN(new_n618));
  INV_X1    g0418(.A(new_n618), .ZN(new_n619));
  INV_X1    g0419(.A(KEYINPUT26), .ZN(new_n620));
  INV_X1    g0420(.A(KEYINPUT90), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n475), .A2(new_n621), .ZN(new_n622));
  NAND3_X1  g0422(.A1(new_n460), .A2(KEYINPUT90), .A3(G200), .ZN(new_n623));
  NAND3_X1  g0423(.A1(new_n474), .A2(new_n622), .A3(new_n623), .ZN(new_n624));
  AND2_X1   g0424(.A1(new_n559), .A2(new_n558), .ZN(new_n625));
  NAND3_X1  g0425(.A1(new_n624), .A2(new_n625), .A3(new_n557), .ZN(new_n626));
  NOR2_X1   g0426(.A1(new_n594), .A2(new_n600), .ZN(new_n627));
  NAND3_X1  g0427(.A1(new_n506), .A2(new_n512), .A3(new_n513), .ZN(new_n628));
  OAI21_X1  g0428(.A(new_n598), .B1(new_n627), .B2(new_n628), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n554), .A2(new_n624), .ZN(new_n630));
  OAI211_X1 g0430(.A(new_n620), .B(new_n626), .C1(new_n629), .C2(new_n630), .ZN(new_n631));
  INV_X1    g0431(.A(new_n560), .ZN(new_n632));
  AOI22_X1  g0432(.A1(new_n464), .A2(new_n461), .B1(new_n474), .B2(new_n475), .ZN(new_n633));
  NAND3_X1  g0433(.A1(new_n632), .A2(KEYINPUT26), .A3(new_n633), .ZN(new_n634));
  AOI21_X1  g0434(.A(new_n619), .B1(new_n631), .B2(new_n634), .ZN(new_n635));
  OAI21_X1  g0435(.A(new_n617), .B1(new_n436), .B2(new_n635), .ZN(new_n636));
  XOR2_X1   g0436(.A(new_n636), .B(KEYINPUT93), .Z(G369));
  NAND3_X1  g0437(.A1(new_n224), .A2(new_n225), .A3(G13), .ZN(new_n638));
  OR2_X1    g0438(.A1(new_n638), .A2(KEYINPUT27), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n638), .A2(KEYINPUT27), .ZN(new_n640));
  NAND3_X1  g0440(.A1(new_n639), .A2(G213), .A3(new_n640), .ZN(new_n641));
  INV_X1    g0441(.A(G343), .ZN(new_n642));
  NOR2_X1   g0442(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  AND2_X1   g0443(.A1(new_n593), .A2(new_n288), .ZN(new_n644));
  OAI21_X1  g0444(.A(new_n643), .B1(new_n644), .B2(new_n578), .ZN(new_n645));
  AOI21_X1  g0445(.A(new_n627), .B1(new_n645), .B2(new_n598), .ZN(new_n646));
  NOR2_X1   g0446(.A1(new_n601), .A2(new_n643), .ZN(new_n647));
  OR2_X1    g0447(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  INV_X1    g0448(.A(new_n643), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n628), .A2(new_n649), .ZN(new_n650));
  NOR2_X1   g0450(.A1(new_n648), .A2(new_n650), .ZN(new_n651));
  NOR2_X1   g0451(.A1(new_n651), .A2(new_n647), .ZN(new_n652));
  NOR2_X1   g0452(.A1(new_n507), .A2(new_n649), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n628), .A2(new_n653), .ZN(new_n654));
  OAI21_X1  g0454(.A(new_n654), .B1(new_n514), .B2(new_n653), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n655), .A2(G330), .ZN(new_n656));
  NOR2_X1   g0456(.A1(new_n648), .A2(new_n656), .ZN(new_n657));
  INV_X1    g0457(.A(new_n657), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n652), .A2(new_n658), .ZN(G399));
  INV_X1    g0459(.A(new_n235), .ZN(new_n660));
  INV_X1    g0460(.A(new_n267), .ZN(new_n661));
  NOR2_X1   g0461(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  INV_X1    g0462(.A(new_n662), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n663), .A2(G1), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n442), .A2(new_n455), .ZN(new_n665));
  OAI22_X1  g0465(.A1(new_n664), .A2(new_n665), .B1(new_n232), .B2(new_n663), .ZN(new_n666));
  XNOR2_X1  g0466(.A(new_n666), .B(KEYINPUT28), .ZN(new_n667));
  NOR2_X1   g0467(.A1(new_n546), .A2(new_n547), .ZN(new_n668));
  INV_X1    g0468(.A(new_n460), .ZN(new_n669));
  NAND4_X1  g0469(.A1(new_n668), .A2(new_n511), .A3(new_n570), .A4(new_n669), .ZN(new_n670));
  INV_X1    g0470(.A(KEYINPUT30), .ZN(new_n671));
  XNOR2_X1  g0471(.A(new_n670), .B(new_n671), .ZN(new_n672));
  NOR2_X1   g0472(.A1(new_n573), .A2(new_n668), .ZN(new_n673));
  AND4_X1   g0473(.A1(new_n308), .A2(new_n673), .A3(new_n460), .A4(new_n503), .ZN(new_n674));
  OAI21_X1  g0474(.A(new_n643), .B1(new_n672), .B2(new_n674), .ZN(new_n675));
  INV_X1    g0475(.A(KEYINPUT31), .ZN(new_n676));
  AND2_X1   g0476(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  OAI21_X1  g0477(.A(new_n675), .B1(new_n602), .B2(new_n643), .ZN(new_n678));
  AOI21_X1  g0478(.A(new_n677), .B1(new_n678), .B2(KEYINPUT31), .ZN(new_n679));
  INV_X1    g0479(.A(G330), .ZN(new_n680));
  NOR2_X1   g0480(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  NAND3_X1  g0481(.A1(new_n632), .A2(new_n620), .A3(new_n633), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n626), .A2(KEYINPUT26), .ZN(new_n683));
  NAND3_X1  g0483(.A1(new_n682), .A2(new_n683), .A3(new_n618), .ZN(new_n684));
  INV_X1    g0484(.A(new_n624), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n554), .A2(new_n560), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n686), .A2(KEYINPUT95), .ZN(new_n687));
  INV_X1    g0487(.A(KEYINPUT95), .ZN(new_n688));
  NAND3_X1  g0488(.A1(new_n554), .A2(new_n560), .A3(new_n688), .ZN(new_n689));
  AOI21_X1  g0489(.A(new_n685), .B1(new_n687), .B2(new_n689), .ZN(new_n690));
  INV_X1    g0490(.A(new_n629), .ZN(new_n691));
  AOI21_X1  g0491(.A(new_n684), .B1(new_n690), .B2(new_n691), .ZN(new_n692));
  OAI21_X1  g0492(.A(KEYINPUT96), .B1(new_n692), .B2(new_n643), .ZN(new_n693));
  AND3_X1   g0493(.A1(new_n682), .A2(new_n683), .A3(new_n618), .ZN(new_n694));
  AND3_X1   g0494(.A1(new_n554), .A2(new_n560), .A3(new_n688), .ZN(new_n695));
  AOI21_X1  g0495(.A(new_n688), .B1(new_n554), .B2(new_n560), .ZN(new_n696));
  OAI21_X1  g0496(.A(new_n624), .B1(new_n695), .B2(new_n696), .ZN(new_n697));
  OAI21_X1  g0497(.A(new_n694), .B1(new_n697), .B2(new_n629), .ZN(new_n698));
  INV_X1    g0498(.A(KEYINPUT96), .ZN(new_n699));
  NAND3_X1  g0499(.A1(new_n698), .A2(new_n699), .A3(new_n649), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n693), .A2(new_n700), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n701), .A2(KEYINPUT29), .ZN(new_n702));
  OR2_X1    g0502(.A1(new_n635), .A2(new_n643), .ZN(new_n703));
  XOR2_X1   g0503(.A(KEYINPUT94), .B(KEYINPUT29), .Z(new_n704));
  NAND2_X1  g0504(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  AOI21_X1  g0505(.A(new_n681), .B1(new_n702), .B2(new_n705), .ZN(new_n706));
  OAI21_X1  g0506(.A(new_n667), .B1(new_n706), .B2(G1), .ZN(G364));
  AOI21_X1  g0507(.A(new_n233), .B1(G20), .B2(new_n310), .ZN(new_n708));
  INV_X1    g0508(.A(new_n708), .ZN(new_n709));
  NOR2_X1   g0509(.A1(new_n225), .A2(G190), .ZN(new_n710));
  NAND3_X1  g0510(.A1(new_n710), .A2(new_n308), .A3(new_n415), .ZN(new_n711));
  INV_X1    g0511(.A(KEYINPUT98), .ZN(new_n712));
  OR2_X1    g0512(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n711), .A2(new_n712), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  INV_X1    g0515(.A(new_n715), .ZN(new_n716));
  NAND3_X1  g0516(.A1(new_n710), .A2(new_n308), .A3(G200), .ZN(new_n717));
  INV_X1    g0517(.A(new_n717), .ZN(new_n718));
  AOI22_X1  g0518(.A1(new_n716), .A2(G329), .B1(G283), .B2(new_n718), .ZN(new_n719));
  XOR2_X1   g0519(.A(new_n719), .B(KEYINPUT100), .Z(new_n720));
  NOR3_X1   g0520(.A1(new_n362), .A2(G179), .A3(G200), .ZN(new_n721));
  NOR2_X1   g0521(.A1(new_n721), .A2(new_n225), .ZN(new_n722));
  INV_X1    g0522(.A(new_n722), .ZN(new_n723));
  NAND3_X1  g0523(.A1(new_n710), .A2(G179), .A3(new_n415), .ZN(new_n724));
  INV_X1    g0524(.A(new_n724), .ZN(new_n725));
  AOI22_X1  g0525(.A1(new_n723), .A2(G294), .B1(new_n725), .B2(G311), .ZN(new_n726));
  INV_X1    g0526(.A(G322), .ZN(new_n727));
  NOR2_X1   g0527(.A1(new_n225), .A2(new_n362), .ZN(new_n728));
  NAND2_X1  g0528(.A1(new_n728), .A2(G179), .ZN(new_n729));
  NOR2_X1   g0529(.A1(new_n729), .A2(G200), .ZN(new_n730));
  INV_X1    g0530(.A(new_n730), .ZN(new_n731));
  OAI21_X1  g0531(.A(new_n726), .B1(new_n727), .B2(new_n731), .ZN(new_n732));
  NOR3_X1   g0532(.A1(new_n720), .A2(new_n271), .A3(new_n732), .ZN(new_n733));
  NAND3_X1  g0533(.A1(new_n710), .A2(G179), .A3(G200), .ZN(new_n734));
  INV_X1    g0534(.A(new_n734), .ZN(new_n735));
  XNOR2_X1  g0535(.A(KEYINPUT33), .B(G317), .ZN(new_n736));
  NAND2_X1  g0536(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  NOR2_X1   g0537(.A1(new_n729), .A2(new_n415), .ZN(new_n738));
  NAND2_X1  g0538(.A1(new_n738), .A2(G326), .ZN(new_n739));
  NAND3_X1  g0539(.A1(new_n728), .A2(new_n308), .A3(G200), .ZN(new_n740));
  INV_X1    g0540(.A(new_n740), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n741), .A2(G303), .ZN(new_n742));
  NAND4_X1  g0542(.A1(new_n733), .A2(new_n737), .A3(new_n739), .A4(new_n742), .ZN(new_n743));
  NAND2_X1  g0543(.A1(new_n716), .A2(G159), .ZN(new_n744));
  XNOR2_X1  g0544(.A(new_n744), .B(KEYINPUT99), .ZN(new_n745));
  XNOR2_X1  g0545(.A(new_n745), .B(KEYINPUT32), .ZN(new_n746));
  OAI22_X1  g0546(.A1(new_n731), .A2(new_n202), .B1(new_n438), .B2(new_n722), .ZN(new_n747));
  AOI21_X1  g0547(.A(new_n372), .B1(new_n735), .B2(G68), .ZN(new_n748));
  INV_X1    g0548(.A(new_n738), .ZN(new_n749));
  OAI221_X1 g0549(.A(new_n748), .B1(new_n217), .B2(new_n717), .C1(new_n749), .C2(new_n249), .ZN(new_n750));
  AOI211_X1 g0550(.A(new_n747), .B(new_n750), .C1(new_n441), .C2(new_n741), .ZN(new_n751));
  OAI211_X1 g0551(.A(new_n746), .B(new_n751), .C1(new_n206), .C2(new_n724), .ZN(new_n752));
  AOI21_X1  g0552(.A(new_n709), .B1(new_n743), .B2(new_n752), .ZN(new_n753));
  NOR2_X1   g0553(.A1(G13), .A2(G33), .ZN(new_n754));
  INV_X1    g0554(.A(new_n754), .ZN(new_n755));
  NOR2_X1   g0555(.A1(new_n755), .A2(G20), .ZN(new_n756));
  NOR2_X1   g0556(.A1(new_n756), .A2(new_n708), .ZN(new_n757));
  NOR2_X1   g0557(.A1(new_n660), .A2(new_n372), .ZN(new_n758));
  AOI22_X1  g0558(.A1(new_n758), .A2(G355), .B1(new_n455), .B2(new_n660), .ZN(new_n759));
  XNOR2_X1  g0559(.A(new_n759), .B(KEYINPUT97), .ZN(new_n760));
  NAND3_X1  g0560(.A1(new_n204), .A2(new_n268), .A3(G50), .ZN(new_n761));
  NOR2_X1   g0561(.A1(new_n660), .A2(new_n271), .ZN(new_n762));
  OAI211_X1 g0562(.A(new_n761), .B(new_n762), .C1(new_n251), .C2(new_n268), .ZN(new_n763));
  NAND2_X1  g0563(.A1(new_n760), .A2(new_n763), .ZN(new_n764));
  AOI21_X1  g0564(.A(new_n753), .B1(new_n757), .B2(new_n764), .ZN(new_n765));
  INV_X1    g0565(.A(G13), .ZN(new_n766));
  NOR2_X1   g0566(.A1(new_n766), .A2(G20), .ZN(new_n767));
  AOI21_X1  g0567(.A(new_n664), .B1(G45), .B2(new_n767), .ZN(new_n768));
  INV_X1    g0568(.A(new_n756), .ZN(new_n769));
  OAI211_X1 g0569(.A(new_n765), .B(new_n768), .C1(new_n655), .C2(new_n769), .ZN(new_n770));
  AOI21_X1  g0570(.A(new_n768), .B1(new_n655), .B2(G330), .ZN(new_n771));
  OAI21_X1  g0571(.A(new_n771), .B1(G330), .B2(new_n655), .ZN(new_n772));
  NAND2_X1  g0572(.A1(new_n770), .A2(new_n772), .ZN(G396));
  XNOR2_X1  g0573(.A(new_n433), .B(KEYINPUT101), .ZN(new_n774));
  NAND2_X1  g0574(.A1(new_n355), .A2(new_n643), .ZN(new_n775));
  AND2_X1   g0575(.A1(new_n363), .A2(new_n775), .ZN(new_n776));
  NAND2_X1  g0576(.A1(new_n774), .A2(new_n776), .ZN(new_n777));
  NOR3_X1   g0577(.A1(new_n635), .A2(new_n643), .A3(new_n777), .ZN(new_n778));
  AOI22_X1  g0578(.A1(new_n774), .A2(new_n776), .B1(new_n433), .B2(new_n643), .ZN(new_n779));
  AOI21_X1  g0579(.A(new_n778), .B1(new_n703), .B2(new_n779), .ZN(new_n780));
  XOR2_X1   g0580(.A(new_n780), .B(new_n681), .Z(new_n781));
  INV_X1    g0581(.A(new_n768), .ZN(new_n782));
  NAND2_X1  g0582(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  INV_X1    g0583(.A(new_n779), .ZN(new_n784));
  NOR2_X1   g0584(.A1(new_n784), .A2(new_n755), .ZN(new_n785));
  NAND2_X1  g0585(.A1(new_n730), .A2(G143), .ZN(new_n786));
  NAND2_X1  g0586(.A1(new_n735), .A2(G150), .ZN(new_n787));
  AND2_X1   g0587(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  INV_X1    g0588(.A(G137), .ZN(new_n789));
  OAI221_X1 g0589(.A(new_n788), .B1(new_n789), .B2(new_n749), .C1(new_n380), .C2(new_n724), .ZN(new_n790));
  INV_X1    g0590(.A(KEYINPUT34), .ZN(new_n791));
  OAI21_X1  g0591(.A(new_n271), .B1(new_n790), .B2(new_n791), .ZN(new_n792));
  INV_X1    g0592(.A(new_n790), .ZN(new_n793));
  OAI22_X1  g0593(.A1(new_n793), .A2(KEYINPUT34), .B1(new_n203), .B2(new_n717), .ZN(new_n794));
  AOI211_X1 g0594(.A(new_n792), .B(new_n794), .C1(G58), .C2(new_n723), .ZN(new_n795));
  INV_X1    g0595(.A(G132), .ZN(new_n796));
  OAI221_X1 g0596(.A(new_n795), .B1(new_n249), .B2(new_n740), .C1(new_n796), .C2(new_n715), .ZN(new_n797));
  INV_X1    g0597(.A(G294), .ZN(new_n798));
  OAI22_X1  g0598(.A1(new_n731), .A2(new_n798), .B1(new_n217), .B2(new_n740), .ZN(new_n799));
  AOI21_X1  g0599(.A(new_n799), .B1(G283), .B2(new_n735), .ZN(new_n800));
  OAI221_X1 g0600(.A(new_n372), .B1(new_n724), .B2(new_n455), .C1(new_n722), .C2(new_n438), .ZN(new_n801));
  AOI21_X1  g0601(.A(new_n801), .B1(new_n716), .B2(G311), .ZN(new_n802));
  AND2_X1   g0602(.A1(new_n800), .A2(new_n802), .ZN(new_n803));
  INV_X1    g0603(.A(G303), .ZN(new_n804));
  OAI221_X1 g0604(.A(new_n803), .B1(new_n409), .B2(new_n717), .C1(new_n804), .C2(new_n749), .ZN(new_n805));
  AOI21_X1  g0605(.A(new_n709), .B1(new_n797), .B2(new_n805), .ZN(new_n806));
  NOR3_X1   g0606(.A1(new_n785), .A2(new_n782), .A3(new_n806), .ZN(new_n807));
  NOR2_X1   g0607(.A1(new_n708), .A2(new_n754), .ZN(new_n808));
  INV_X1    g0608(.A(new_n808), .ZN(new_n809));
  OAI21_X1  g0609(.A(new_n807), .B1(G77), .B2(new_n809), .ZN(new_n810));
  NAND2_X1  g0610(.A1(new_n783), .A2(new_n810), .ZN(G384));
  NAND3_X1  g0611(.A1(new_n702), .A2(new_n435), .A3(new_n705), .ZN(new_n812));
  AND2_X1   g0612(.A1(new_n617), .A2(new_n812), .ZN(new_n813));
  INV_X1    g0613(.A(new_n641), .ZN(new_n814));
  NOR2_X1   g0614(.A1(new_n430), .A2(new_n814), .ZN(new_n815));
  INV_X1    g0615(.A(new_n815), .ZN(new_n816));
  NAND2_X1  g0616(.A1(new_n338), .A2(new_n643), .ZN(new_n817));
  AND3_X1   g0617(.A1(new_n341), .A2(KEYINPUT102), .A3(new_n817), .ZN(new_n818));
  AOI21_X1  g0618(.A(new_n817), .B1(new_n341), .B2(KEYINPUT102), .ZN(new_n819));
  NOR2_X1   g0619(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  INV_X1    g0620(.A(new_n820), .ZN(new_n821));
  NOR2_X1   g0621(.A1(new_n774), .A2(new_n643), .ZN(new_n822));
  OAI21_X1  g0622(.A(new_n821), .B1(new_n778), .B2(new_n822), .ZN(new_n823));
  OAI211_X1 g0623(.A(new_n419), .B(new_n422), .C1(new_n428), .C2(new_n429), .ZN(new_n824));
  NAND2_X1  g0624(.A1(new_n390), .A2(new_n288), .ZN(new_n825));
  AOI21_X1  g0625(.A(KEYINPUT16), .B1(new_n377), .B2(new_n389), .ZN(new_n826));
  OAI21_X1  g0626(.A(new_n403), .B1(new_n825), .B2(new_n826), .ZN(new_n827));
  NAND3_X1  g0627(.A1(new_n824), .A2(new_n814), .A3(new_n827), .ZN(new_n828));
  NAND3_X1  g0628(.A1(new_n425), .A2(new_n426), .A3(new_n641), .ZN(new_n829));
  NAND2_X1  g0629(.A1(new_n424), .A2(new_n829), .ZN(new_n830));
  INV_X1    g0630(.A(KEYINPUT37), .ZN(new_n831));
  OAI211_X1 g0631(.A(new_n830), .B(new_n831), .C1(new_n416), .C2(new_n421), .ZN(new_n832));
  NOR2_X1   g0632(.A1(new_n421), .A2(new_n416), .ZN(new_n833));
  AOI21_X1  g0633(.A(new_n833), .B1(new_n829), .B2(new_n827), .ZN(new_n834));
  OAI21_X1  g0634(.A(new_n832), .B1(new_n834), .B2(new_n831), .ZN(new_n835));
  NAND3_X1  g0635(.A1(new_n828), .A2(KEYINPUT38), .A3(new_n835), .ZN(new_n836));
  INV_X1    g0636(.A(new_n836), .ZN(new_n837));
  AOI21_X1  g0637(.A(KEYINPUT38), .B1(new_n828), .B2(new_n835), .ZN(new_n838));
  NOR2_X1   g0638(.A1(new_n837), .A2(new_n838), .ZN(new_n839));
  OAI21_X1  g0639(.A(new_n816), .B1(new_n823), .B2(new_n839), .ZN(new_n840));
  INV_X1    g0640(.A(new_n840), .ZN(new_n841));
  INV_X1    g0641(.A(new_n829), .ZN(new_n842));
  OAI22_X1  g0642(.A1(new_n406), .A2(new_n842), .B1(new_n421), .B2(new_n416), .ZN(new_n843));
  NAND2_X1  g0643(.A1(new_n843), .A2(KEYINPUT37), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n844), .A2(new_n832), .ZN(new_n845));
  INV_X1    g0645(.A(KEYINPUT103), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  NAND3_X1  g0647(.A1(new_n824), .A2(new_n424), .A3(new_n814), .ZN(new_n848));
  NAND3_X1  g0648(.A1(new_n844), .A2(KEYINPUT103), .A3(new_n832), .ZN(new_n849));
  NAND3_X1  g0649(.A1(new_n847), .A2(new_n848), .A3(new_n849), .ZN(new_n850));
  INV_X1    g0650(.A(KEYINPUT38), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  AOI21_X1  g0652(.A(KEYINPUT39), .B1(new_n852), .B2(new_n836), .ZN(new_n853));
  INV_X1    g0653(.A(KEYINPUT39), .ZN(new_n854));
  NOR3_X1   g0654(.A1(new_n837), .A2(new_n838), .A3(new_n854), .ZN(new_n855));
  NOR2_X1   g0655(.A1(new_n853), .A2(new_n855), .ZN(new_n856));
  INV_X1    g0656(.A(new_n856), .ZN(new_n857));
  NOR2_X1   g0657(.A1(new_n605), .A2(new_n643), .ZN(new_n858));
  INV_X1    g0658(.A(new_n858), .ZN(new_n859));
  OAI21_X1  g0659(.A(new_n841), .B1(new_n857), .B2(new_n859), .ZN(new_n860));
  XNOR2_X1  g0660(.A(new_n813), .B(new_n860), .ZN(new_n861));
  INV_X1    g0661(.A(KEYINPUT40), .ZN(new_n862));
  AOI21_X1  g0662(.A(new_n862), .B1(new_n852), .B2(new_n836), .ZN(new_n863));
  NOR3_X1   g0663(.A1(new_n679), .A2(new_n820), .A3(new_n779), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n678), .A2(KEYINPUT31), .ZN(new_n865));
  INV_X1    g0665(.A(new_n677), .ZN(new_n866));
  AOI21_X1  g0666(.A(new_n779), .B1(new_n865), .B2(new_n866), .ZN(new_n867));
  OAI211_X1 g0667(.A(new_n867), .B(new_n821), .C1(new_n837), .C2(new_n838), .ZN(new_n868));
  AOI22_X1  g0668(.A1(new_n863), .A2(new_n864), .B1(new_n868), .B2(new_n862), .ZN(new_n869));
  NOR2_X1   g0669(.A1(new_n436), .A2(new_n679), .ZN(new_n870));
  XOR2_X1   g0670(.A(new_n869), .B(new_n870), .Z(new_n871));
  NAND2_X1  g0671(.A1(new_n871), .A2(G330), .ZN(new_n872));
  XNOR2_X1  g0672(.A(new_n861), .B(new_n872), .ZN(new_n873));
  OAI21_X1  g0673(.A(new_n873), .B1(new_n224), .B2(new_n767), .ZN(new_n874));
  AOI21_X1  g0674(.A(new_n455), .B1(new_n534), .B2(KEYINPUT35), .ZN(new_n875));
  NOR2_X1   g0675(.A1(new_n233), .A2(new_n225), .ZN(new_n876));
  OAI211_X1 g0676(.A(new_n875), .B(new_n876), .C1(KEYINPUT35), .C2(new_n534), .ZN(new_n877));
  XNOR2_X1  g0677(.A(new_n877), .B(KEYINPUT36), .ZN(new_n878));
  NOR3_X1   g0678(.A1(new_n232), .A2(new_n206), .A3(new_n383), .ZN(new_n879));
  NOR2_X1   g0679(.A1(new_n201), .A2(new_n203), .ZN(new_n880));
  OAI211_X1 g0680(.A(G1), .B(new_n766), .C1(new_n879), .C2(new_n880), .ZN(new_n881));
  NAND3_X1  g0681(.A1(new_n874), .A2(new_n878), .A3(new_n881), .ZN(G367));
  NAND2_X1  g0682(.A1(new_n687), .A2(new_n689), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n557), .A2(new_n643), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  OAI21_X1  g0685(.A(new_n885), .B1(new_n560), .B2(new_n649), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n651), .A2(new_n886), .ZN(new_n887));
  XNOR2_X1  g0687(.A(new_n887), .B(KEYINPUT42), .ZN(new_n888));
  NAND3_X1  g0688(.A1(new_n883), .A2(new_n627), .A3(new_n884), .ZN(new_n889));
  AOI21_X1  g0689(.A(new_n643), .B1(new_n889), .B2(new_n560), .ZN(new_n890));
  OR2_X1    g0690(.A1(new_n888), .A2(new_n890), .ZN(new_n891));
  AOI21_X1  g0691(.A(new_n649), .B1(new_n446), .B2(new_n473), .ZN(new_n892));
  INV_X1    g0692(.A(new_n892), .ZN(new_n893));
  NAND3_X1  g0693(.A1(new_n624), .A2(new_n618), .A3(new_n893), .ZN(new_n894));
  OAI21_X1  g0694(.A(new_n894), .B1(new_n618), .B2(new_n893), .ZN(new_n895));
  NOR3_X1   g0695(.A1(new_n891), .A2(KEYINPUT43), .A3(new_n895), .ZN(new_n896));
  XNOR2_X1  g0696(.A(new_n896), .B(KEYINPUT104), .ZN(new_n897));
  XOR2_X1   g0697(.A(new_n895), .B(KEYINPUT43), .Z(new_n898));
  NAND2_X1  g0698(.A1(new_n891), .A2(new_n898), .ZN(new_n899));
  XNOR2_X1  g0699(.A(new_n899), .B(KEYINPUT105), .ZN(new_n900));
  NOR2_X1   g0700(.A1(new_n897), .A2(new_n900), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n657), .A2(new_n886), .ZN(new_n902));
  XOR2_X1   g0702(.A(new_n901), .B(new_n902), .Z(new_n903));
  AOI21_X1  g0703(.A(new_n224), .B1(new_n767), .B2(G45), .ZN(new_n904));
  INV_X1    g0704(.A(new_n904), .ZN(new_n905));
  NOR2_X1   g0705(.A1(new_n652), .A2(new_n886), .ZN(new_n906));
  XOR2_X1   g0706(.A(new_n906), .B(KEYINPUT44), .Z(new_n907));
  NAND2_X1  g0707(.A1(new_n652), .A2(new_n886), .ZN(new_n908));
  XNOR2_X1  g0708(.A(new_n908), .B(KEYINPUT45), .ZN(new_n909));
  NOR2_X1   g0709(.A1(new_n907), .A2(new_n909), .ZN(new_n910));
  XNOR2_X1  g0710(.A(new_n910), .B(new_n658), .ZN(new_n911));
  XOR2_X1   g0711(.A(new_n648), .B(new_n650), .Z(new_n912));
  XNOR2_X1  g0712(.A(new_n912), .B(new_n656), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n913), .A2(new_n706), .ZN(new_n914));
  OR2_X1    g0714(.A1(new_n911), .A2(new_n914), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n915), .A2(new_n706), .ZN(new_n916));
  XNOR2_X1  g0716(.A(new_n662), .B(KEYINPUT41), .ZN(new_n917));
  AOI21_X1  g0717(.A(new_n905), .B1(new_n916), .B2(new_n917), .ZN(new_n918));
  NOR2_X1   g0718(.A1(new_n895), .A2(new_n769), .ZN(new_n919));
  INV_X1    g0719(.A(new_n762), .ZN(new_n920));
  OAI221_X1 g0720(.A(new_n757), .B1(new_n235), .B2(new_n350), .C1(new_n246), .C2(new_n920), .ZN(new_n921));
  XNOR2_X1  g0721(.A(new_n921), .B(KEYINPUT106), .ZN(new_n922));
  AOI22_X1  g0722(.A1(new_n723), .A2(G68), .B1(new_n725), .B2(new_n201), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n738), .A2(G143), .ZN(new_n924));
  INV_X1    g0724(.A(G150), .ZN(new_n925));
  OAI211_X1 g0725(.A(new_n923), .B(new_n924), .C1(new_n925), .C2(new_n731), .ZN(new_n926));
  AOI22_X1  g0726(.A1(G58), .A2(new_n741), .B1(new_n718), .B2(G77), .ZN(new_n927));
  OAI211_X1 g0727(.A(new_n271), .B(new_n927), .C1(new_n715), .C2(new_n789), .ZN(new_n928));
  AOI211_X1 g0728(.A(new_n926), .B(new_n928), .C1(G159), .C2(new_n735), .ZN(new_n929));
  XNOR2_X1  g0729(.A(new_n929), .B(KEYINPUT108), .ZN(new_n930));
  AND2_X1   g0730(.A1(new_n716), .A2(G317), .ZN(new_n931));
  INV_X1    g0731(.A(KEYINPUT107), .ZN(new_n932));
  OAI21_X1  g0732(.A(new_n932), .B1(new_n740), .B2(new_n455), .ZN(new_n933));
  OAI221_X1 g0733(.A(new_n372), .B1(new_n933), .B2(KEYINPUT46), .C1(new_n804), .C2(new_n731), .ZN(new_n934));
  AOI21_X1  g0734(.A(new_n934), .B1(G107), .B2(new_n723), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n738), .A2(G311), .ZN(new_n936));
  AOI22_X1  g0736(.A1(new_n735), .A2(G294), .B1(new_n718), .B2(G97), .ZN(new_n937));
  INV_X1    g0737(.A(G283), .ZN(new_n938));
  OAI21_X1  g0738(.A(new_n937), .B1(new_n938), .B2(new_n724), .ZN(new_n939));
  AOI21_X1  g0739(.A(new_n939), .B1(KEYINPUT46), .B2(new_n933), .ZN(new_n940));
  NAND3_X1  g0740(.A1(new_n935), .A2(new_n936), .A3(new_n940), .ZN(new_n941));
  OAI21_X1  g0741(.A(new_n930), .B1(new_n931), .B2(new_n941), .ZN(new_n942));
  XOR2_X1   g0742(.A(new_n942), .B(KEYINPUT47), .Z(new_n943));
  OAI211_X1 g0743(.A(new_n768), .B(new_n922), .C1(new_n943), .C2(new_n709), .ZN(new_n944));
  OAI22_X1  g0744(.A1(new_n903), .A2(new_n918), .B1(new_n919), .B2(new_n944), .ZN(G387));
  NAND2_X1  g0745(.A1(new_n913), .A2(new_n905), .ZN(new_n946));
  OAI21_X1  g0746(.A(new_n271), .B1(new_n734), .B2(new_n342), .ZN(new_n947));
  AOI21_X1  g0747(.A(new_n947), .B1(new_n716), .B2(G150), .ZN(new_n948));
  NOR2_X1   g0748(.A1(new_n740), .A2(new_n206), .ZN(new_n949));
  OAI22_X1  g0749(.A1(new_n203), .A2(new_n724), .B1(new_n717), .B2(new_n438), .ZN(new_n950));
  AOI211_X1 g0750(.A(new_n949), .B(new_n950), .C1(G159), .C2(new_n738), .ZN(new_n951));
  NAND3_X1  g0751(.A1(new_n348), .A2(new_n723), .A3(new_n349), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n730), .A2(G50), .ZN(new_n953));
  NAND4_X1  g0753(.A1(new_n948), .A2(new_n951), .A3(new_n952), .A4(new_n953), .ZN(new_n954));
  AOI22_X1  g0754(.A1(new_n730), .A2(G317), .B1(new_n735), .B2(G311), .ZN(new_n955));
  OAI221_X1 g0755(.A(new_n955), .B1(new_n804), .B2(new_n724), .C1(new_n727), .C2(new_n749), .ZN(new_n956));
  XNOR2_X1  g0756(.A(new_n956), .B(KEYINPUT48), .ZN(new_n957));
  OAI221_X1 g0757(.A(new_n957), .B1(new_n938), .B2(new_n722), .C1(new_n798), .C2(new_n740), .ZN(new_n958));
  XOR2_X1   g0758(.A(new_n958), .B(KEYINPUT49), .Z(new_n959));
  INV_X1    g0759(.A(G326), .ZN(new_n960));
  OAI221_X1 g0760(.A(new_n372), .B1(new_n455), .B2(new_n717), .C1(new_n715), .C2(new_n960), .ZN(new_n961));
  OAI21_X1  g0761(.A(new_n954), .B1(new_n959), .B2(new_n961), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n962), .A2(new_n708), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n281), .A2(new_n249), .ZN(new_n964));
  XNOR2_X1  g0764(.A(new_n964), .B(KEYINPUT50), .ZN(new_n965));
  NOR2_X1   g0765(.A1(new_n203), .A2(new_n206), .ZN(new_n966));
  NOR4_X1   g0766(.A1(new_n965), .A2(G45), .A3(new_n966), .A4(new_n665), .ZN(new_n967));
  INV_X1    g0767(.A(new_n243), .ZN(new_n968));
  OAI21_X1  g0768(.A(new_n762), .B1(new_n968), .B2(new_n268), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n758), .A2(new_n665), .ZN(new_n970));
  AOI21_X1  g0770(.A(new_n967), .B1(new_n969), .B2(new_n970), .ZN(new_n971));
  NOR2_X1   g0771(.A1(new_n235), .A2(G107), .ZN(new_n972));
  OAI21_X1  g0772(.A(new_n757), .B1(new_n971), .B2(new_n972), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n648), .A2(new_n756), .ZN(new_n974));
  NAND4_X1  g0774(.A1(new_n963), .A2(new_n768), .A3(new_n973), .A4(new_n974), .ZN(new_n975));
  INV_X1    g0775(.A(new_n914), .ZN(new_n976));
  OAI21_X1  g0776(.A(new_n662), .B1(new_n913), .B2(new_n706), .ZN(new_n977));
  OAI211_X1 g0777(.A(new_n946), .B(new_n975), .C1(new_n976), .C2(new_n977), .ZN(G393));
  AOI21_X1  g0778(.A(new_n663), .B1(new_n911), .B2(new_n914), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n915), .A2(new_n979), .ZN(new_n980));
  AOI22_X1  g0780(.A1(G311), .A2(new_n730), .B1(new_n738), .B2(G317), .ZN(new_n981));
  XNOR2_X1  g0781(.A(new_n981), .B(KEYINPUT110), .ZN(new_n982));
  XNOR2_X1  g0782(.A(new_n982), .B(KEYINPUT52), .ZN(new_n983));
  AOI22_X1  g0783(.A1(new_n723), .A2(G116), .B1(new_n741), .B2(G283), .ZN(new_n984));
  OAI21_X1  g0784(.A(new_n984), .B1(new_n798), .B2(new_n724), .ZN(new_n985));
  AOI21_X1  g0785(.A(new_n985), .B1(G322), .B2(new_n716), .ZN(new_n986));
  OAI211_X1 g0786(.A(new_n983), .B(new_n986), .C1(new_n804), .C2(new_n734), .ZN(new_n987));
  AOI211_X1 g0787(.A(new_n271), .B(new_n987), .C1(G107), .C2(new_n718), .ZN(new_n988));
  AOI22_X1  g0788(.A1(G150), .A2(new_n738), .B1(new_n730), .B2(G159), .ZN(new_n989));
  XOR2_X1   g0789(.A(new_n989), .B(KEYINPUT51), .Z(new_n990));
  NAND2_X1  g0790(.A1(new_n723), .A2(G77), .ZN(new_n991));
  NAND2_X1  g0791(.A1(new_n716), .A2(G143), .ZN(new_n992));
  NAND4_X1  g0792(.A1(new_n990), .A2(new_n271), .A3(new_n991), .A4(new_n992), .ZN(new_n993));
  NOR2_X1   g0793(.A1(new_n724), .A2(new_n342), .ZN(new_n994));
  NOR2_X1   g0794(.A1(new_n740), .A2(new_n203), .ZN(new_n995));
  INV_X1    g0795(.A(new_n201), .ZN(new_n996));
  OAI22_X1  g0796(.A1(new_n996), .A2(new_n734), .B1(new_n717), .B2(new_n409), .ZN(new_n997));
  NOR4_X1   g0797(.A1(new_n993), .A2(new_n994), .A3(new_n995), .A4(new_n997), .ZN(new_n998));
  OAI21_X1  g0798(.A(new_n708), .B1(new_n988), .B2(new_n998), .ZN(new_n999));
  OAI221_X1 g0799(.A(new_n757), .B1(new_n438), .B2(new_n235), .C1(new_n920), .C2(new_n254), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n768), .A2(new_n1000), .ZN(new_n1001));
  XOR2_X1   g0801(.A(new_n1001), .B(KEYINPUT109), .Z(new_n1002));
  OAI211_X1 g0802(.A(new_n999), .B(new_n1002), .C1(new_n886), .C2(new_n769), .ZN(new_n1003));
  OAI211_X1 g0803(.A(new_n980), .B(new_n1003), .C1(new_n904), .C2(new_n911), .ZN(G390));
  AND3_X1   g0804(.A1(new_n844), .A2(KEYINPUT103), .A3(new_n832), .ZN(new_n1005));
  AOI21_X1  g0805(.A(KEYINPUT103), .B1(new_n844), .B2(new_n832), .ZN(new_n1006));
  NOR2_X1   g0806(.A1(new_n1005), .A2(new_n1006), .ZN(new_n1007));
  AOI21_X1  g0807(.A(KEYINPUT38), .B1(new_n1007), .B2(new_n848), .ZN(new_n1008));
  OAI21_X1  g0808(.A(new_n854), .B1(new_n1008), .B2(new_n837), .ZN(new_n1009));
  INV_X1    g0809(.A(new_n838), .ZN(new_n1010));
  NAND3_X1  g0810(.A1(new_n1010), .A2(KEYINPUT39), .A3(new_n836), .ZN(new_n1011));
  AOI22_X1  g0811(.A1(new_n1009), .A2(new_n1011), .B1(new_n859), .B2(new_n823), .ZN(new_n1012));
  INV_X1    g0812(.A(KEYINPUT111), .ZN(new_n1013));
  NOR3_X1   g0813(.A1(new_n692), .A2(KEYINPUT96), .A3(new_n643), .ZN(new_n1014));
  AOI21_X1  g0814(.A(new_n699), .B1(new_n698), .B2(new_n649), .ZN(new_n1015));
  OAI21_X1  g0815(.A(new_n784), .B1(new_n1014), .B2(new_n1015), .ZN(new_n1016));
  INV_X1    g0816(.A(new_n822), .ZN(new_n1017));
  AOI21_X1  g0817(.A(new_n820), .B1(new_n1016), .B2(new_n1017), .ZN(new_n1018));
  OAI21_X1  g0818(.A(new_n859), .B1(new_n1008), .B2(new_n837), .ZN(new_n1019));
  OAI21_X1  g0819(.A(new_n1013), .B1(new_n1018), .B2(new_n1019), .ZN(new_n1020));
  AOI21_X1  g0820(.A(new_n779), .B1(new_n693), .B2(new_n700), .ZN(new_n1021));
  OAI21_X1  g0821(.A(new_n821), .B1(new_n1021), .B2(new_n822), .ZN(new_n1022));
  AOI21_X1  g0822(.A(new_n858), .B1(new_n852), .B2(new_n836), .ZN(new_n1023));
  NAND3_X1  g0823(.A1(new_n1022), .A2(KEYINPUT111), .A3(new_n1023), .ZN(new_n1024));
  AOI21_X1  g0824(.A(new_n1012), .B1(new_n1020), .B2(new_n1024), .ZN(new_n1025));
  NAND2_X1  g0825(.A1(new_n681), .A2(new_n784), .ZN(new_n1026));
  NOR2_X1   g0826(.A1(new_n1026), .A2(new_n820), .ZN(new_n1027));
  INV_X1    g0827(.A(new_n1027), .ZN(new_n1028));
  OAI21_X1  g0828(.A(KEYINPUT112), .B1(new_n1025), .B2(new_n1028), .ZN(new_n1029));
  NAND2_X1  g0829(.A1(new_n823), .A2(new_n859), .ZN(new_n1030));
  OAI21_X1  g0830(.A(new_n1030), .B1(new_n853), .B2(new_n855), .ZN(new_n1031));
  AND3_X1   g0831(.A1(new_n1022), .A2(KEYINPUT111), .A3(new_n1023), .ZN(new_n1032));
  AOI21_X1  g0832(.A(KEYINPUT111), .B1(new_n1022), .B2(new_n1023), .ZN(new_n1033));
  OAI21_X1  g0833(.A(new_n1031), .B1(new_n1032), .B2(new_n1033), .ZN(new_n1034));
  INV_X1    g0834(.A(KEYINPUT112), .ZN(new_n1035));
  NAND3_X1  g0835(.A1(new_n1034), .A2(new_n1035), .A3(new_n1027), .ZN(new_n1036));
  NAND2_X1  g0836(.A1(new_n1029), .A2(new_n1036), .ZN(new_n1037));
  INV_X1    g0837(.A(KEYINPUT113), .ZN(new_n1038));
  OAI21_X1  g0838(.A(new_n1038), .B1(new_n1034), .B2(new_n1027), .ZN(new_n1039));
  NAND3_X1  g0839(.A1(new_n1025), .A2(KEYINPUT113), .A3(new_n1028), .ZN(new_n1040));
  NAND4_X1  g0840(.A1(new_n1037), .A2(new_n905), .A3(new_n1039), .A4(new_n1040), .ZN(new_n1041));
  XNOR2_X1  g0841(.A(new_n1041), .B(KEYINPUT114), .ZN(new_n1042));
  NAND3_X1  g0842(.A1(new_n1037), .A2(new_n1039), .A3(new_n1040), .ZN(new_n1043));
  NAND2_X1  g0843(.A1(new_n870), .A2(G330), .ZN(new_n1044));
  NAND3_X1  g0844(.A1(new_n617), .A2(new_n812), .A3(new_n1044), .ZN(new_n1045));
  NAND2_X1  g0845(.A1(new_n1026), .A2(new_n820), .ZN(new_n1046));
  NAND2_X1  g0846(.A1(new_n1028), .A2(new_n1046), .ZN(new_n1047));
  OAI21_X1  g0847(.A(new_n1047), .B1(new_n778), .B2(new_n822), .ZN(new_n1048));
  NAND4_X1  g0848(.A1(new_n1046), .A2(new_n1017), .A3(new_n1028), .A4(new_n1016), .ZN(new_n1049));
  AOI21_X1  g0849(.A(new_n1045), .B1(new_n1048), .B2(new_n1049), .ZN(new_n1050));
  INV_X1    g0850(.A(new_n1050), .ZN(new_n1051));
  NAND2_X1  g0851(.A1(new_n1043), .A2(new_n1051), .ZN(new_n1052));
  NAND4_X1  g0852(.A1(new_n1037), .A2(new_n1050), .A3(new_n1039), .A4(new_n1040), .ZN(new_n1053));
  NAND3_X1  g0853(.A1(new_n1052), .A2(new_n662), .A3(new_n1053), .ZN(new_n1054));
  NAND2_X1  g0854(.A1(new_n857), .A2(new_n754), .ZN(new_n1055));
  NAND2_X1  g0855(.A1(new_n808), .A2(new_n342), .ZN(new_n1056));
  AOI21_X1  g0856(.A(new_n271), .B1(new_n716), .B2(G294), .ZN(new_n1057));
  AOI22_X1  g0857(.A1(new_n723), .A2(G77), .B1(new_n725), .B2(G97), .ZN(new_n1058));
  OAI211_X1 g0858(.A(new_n1057), .B(new_n1058), .C1(new_n217), .C2(new_n734), .ZN(new_n1059));
  NOR2_X1   g0859(.A1(new_n749), .A2(new_n938), .ZN(new_n1060));
  NOR2_X1   g0860(.A1(new_n740), .A2(new_n409), .ZN(new_n1061));
  OAI22_X1  g0861(.A1(new_n731), .A2(new_n455), .B1(new_n717), .B2(new_n203), .ZN(new_n1062));
  NOR4_X1   g0862(.A1(new_n1059), .A2(new_n1060), .A3(new_n1061), .A4(new_n1062), .ZN(new_n1063));
  NAND2_X1  g0863(.A1(new_n716), .A2(G125), .ZN(new_n1064));
  NAND2_X1  g0864(.A1(new_n738), .A2(G128), .ZN(new_n1065));
  NAND2_X1  g0865(.A1(new_n741), .A2(G150), .ZN(new_n1066));
  XOR2_X1   g0866(.A(KEYINPUT115), .B(KEYINPUT53), .Z(new_n1067));
  NAND2_X1  g0867(.A1(new_n1066), .A2(new_n1067), .ZN(new_n1068));
  XOR2_X1   g0868(.A(KEYINPUT54), .B(G143), .Z(new_n1069));
  AOI22_X1  g0869(.A1(new_n735), .A2(G137), .B1(new_n725), .B2(new_n1069), .ZN(new_n1070));
  NAND4_X1  g0870(.A1(new_n1064), .A2(new_n1065), .A3(new_n1068), .A4(new_n1070), .ZN(new_n1071));
  NOR2_X1   g0871(.A1(new_n731), .A2(new_n796), .ZN(new_n1072));
  NOR2_X1   g0872(.A1(new_n996), .A2(new_n717), .ZN(new_n1073));
  OAI221_X1 g0873(.A(new_n271), .B1(new_n380), .B2(new_n722), .C1(new_n1066), .C2(new_n1067), .ZN(new_n1074));
  NOR4_X1   g0874(.A1(new_n1071), .A2(new_n1072), .A3(new_n1073), .A4(new_n1074), .ZN(new_n1075));
  OAI21_X1  g0875(.A(new_n708), .B1(new_n1063), .B2(new_n1075), .ZN(new_n1076));
  NAND4_X1  g0876(.A1(new_n1055), .A2(new_n768), .A3(new_n1056), .A4(new_n1076), .ZN(new_n1077));
  NAND3_X1  g0877(.A1(new_n1042), .A2(new_n1054), .A3(new_n1077), .ZN(G378));
  INV_X1    g0878(.A(KEYINPUT57), .ZN(new_n1079));
  INV_X1    g0879(.A(new_n1045), .ZN(new_n1080));
  AND2_X1   g0880(.A1(new_n1053), .A2(new_n1080), .ZN(new_n1081));
  XOR2_X1   g0881(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1082));
  INV_X1    g0882(.A(new_n1082), .ZN(new_n1083));
  AOI21_X1  g0883(.A(new_n1083), .B1(new_n307), .B2(new_n312), .ZN(new_n1084));
  INV_X1    g0884(.A(new_n1084), .ZN(new_n1085));
  NAND2_X1  g0885(.A1(new_n292), .A2(new_n814), .ZN(new_n1086));
  INV_X1    g0886(.A(new_n1086), .ZN(new_n1087));
  NAND3_X1  g0887(.A1(new_n307), .A2(new_n312), .A3(new_n1083), .ZN(new_n1088));
  NAND3_X1  g0888(.A1(new_n1085), .A2(new_n1087), .A3(new_n1088), .ZN(new_n1089));
  INV_X1    g0889(.A(new_n312), .ZN(new_n1090));
  AOI211_X1 g0890(.A(new_n1090), .B(new_n1082), .C1(new_n300), .C2(new_n306), .ZN(new_n1091));
  OAI21_X1  g0891(.A(new_n1086), .B1(new_n1084), .B2(new_n1091), .ZN(new_n1092));
  INV_X1    g0892(.A(KEYINPUT117), .ZN(new_n1093));
  AND3_X1   g0893(.A1(new_n1089), .A2(new_n1092), .A3(new_n1093), .ZN(new_n1094));
  AOI21_X1  g0894(.A(new_n1093), .B1(new_n1089), .B2(new_n1092), .ZN(new_n1095));
  NOR2_X1   g0895(.A1(new_n1094), .A2(new_n1095), .ZN(new_n1096));
  AOI21_X1  g0896(.A(new_n1096), .B1(new_n869), .B2(G330), .ZN(new_n1097));
  NAND2_X1  g0897(.A1(new_n868), .A2(new_n862), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n1089), .A2(new_n1092), .ZN(new_n1099));
  NAND2_X1  g0899(.A1(new_n1099), .A2(KEYINPUT117), .ZN(new_n1100));
  OAI211_X1 g0900(.A(new_n864), .B(KEYINPUT40), .C1(new_n1008), .C2(new_n837), .ZN(new_n1101));
  NAND4_X1  g0901(.A1(new_n1098), .A2(new_n1100), .A3(new_n1101), .A4(G330), .ZN(new_n1102));
  INV_X1    g0902(.A(new_n1102), .ZN(new_n1103));
  OAI21_X1  g0903(.A(new_n860), .B1(new_n1097), .B2(new_n1103), .ZN(new_n1104));
  NAND3_X1  g0904(.A1(new_n1098), .A2(new_n1101), .A3(G330), .ZN(new_n1105));
  NAND3_X1  g0905(.A1(new_n1089), .A2(new_n1092), .A3(new_n1093), .ZN(new_n1106));
  NAND2_X1  g0906(.A1(new_n1100), .A2(new_n1106), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n1105), .A2(new_n1107), .ZN(new_n1108));
  AOI21_X1  g0908(.A(new_n840), .B1(new_n856), .B2(new_n858), .ZN(new_n1109));
  NAND3_X1  g0909(.A1(new_n1108), .A2(new_n1109), .A3(new_n1102), .ZN(new_n1110));
  AOI21_X1  g0910(.A(KEYINPUT118), .B1(new_n1104), .B2(new_n1110), .ZN(new_n1111));
  AOI21_X1  g0911(.A(new_n1109), .B1(new_n1108), .B2(new_n1102), .ZN(new_n1112));
  INV_X1    g0912(.A(KEYINPUT118), .ZN(new_n1113));
  NOR2_X1   g0913(.A1(new_n1112), .A2(new_n1113), .ZN(new_n1114));
  OAI21_X1  g0914(.A(KEYINPUT119), .B1(new_n1111), .B2(new_n1114), .ZN(new_n1115));
  AND3_X1   g0915(.A1(new_n1108), .A2(new_n1109), .A3(new_n1102), .ZN(new_n1116));
  OAI21_X1  g0916(.A(new_n1113), .B1(new_n1116), .B2(new_n1112), .ZN(new_n1117));
  INV_X1    g0917(.A(KEYINPUT119), .ZN(new_n1118));
  NAND2_X1  g0918(.A1(new_n1104), .A2(KEYINPUT118), .ZN(new_n1119));
  NAND3_X1  g0919(.A1(new_n1117), .A2(new_n1118), .A3(new_n1119), .ZN(new_n1120));
  NAND2_X1  g0920(.A1(new_n1115), .A2(new_n1120), .ZN(new_n1121));
  OAI21_X1  g0921(.A(new_n1079), .B1(new_n1081), .B2(new_n1121), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n1122), .A2(KEYINPUT120), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n1053), .A2(new_n1080), .ZN(new_n1124));
  NAND2_X1  g0924(.A1(new_n1104), .A2(new_n1110), .ZN(new_n1125));
  NAND3_X1  g0925(.A1(new_n1124), .A2(KEYINPUT57), .A3(new_n1125), .ZN(new_n1126));
  INV_X1    g0926(.A(KEYINPUT120), .ZN(new_n1127));
  OAI211_X1 g0927(.A(new_n1127), .B(new_n1079), .C1(new_n1081), .C2(new_n1121), .ZN(new_n1128));
  NAND4_X1  g0928(.A1(new_n1123), .A2(new_n662), .A3(new_n1126), .A4(new_n1128), .ZN(new_n1129));
  AOI21_X1  g0929(.A(new_n755), .B1(new_n1089), .B2(new_n1092), .ZN(new_n1130));
  AOI21_X1  g0930(.A(new_n949), .B1(G97), .B2(new_n735), .ZN(new_n1131));
  OAI221_X1 g0931(.A(new_n1131), .B1(new_n203), .B2(new_n722), .C1(new_n217), .C2(new_n731), .ZN(new_n1132));
  NAND2_X1  g0932(.A1(new_n372), .A2(new_n267), .ZN(new_n1133));
  NOR2_X1   g0933(.A1(new_n717), .A2(new_n202), .ZN(new_n1134));
  NOR2_X1   g0934(.A1(new_n749), .A2(new_n455), .ZN(new_n1135));
  NOR4_X1   g0935(.A1(new_n1132), .A2(new_n1133), .A3(new_n1134), .A4(new_n1135), .ZN(new_n1136));
  OAI221_X1 g0936(.A(new_n1136), .B1(new_n938), .B2(new_n715), .C1(new_n350), .C2(new_n724), .ZN(new_n1137));
  XNOR2_X1  g0937(.A(new_n1137), .B(KEYINPUT58), .ZN(new_n1138));
  NOR2_X1   g0938(.A1(G33), .A2(G41), .ZN(new_n1139));
  AOI211_X1 g0939(.A(G50), .B(new_n1139), .C1(new_n372), .C2(new_n267), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n741), .A2(new_n1069), .ZN(new_n1141));
  XOR2_X1   g0941(.A(new_n1141), .B(KEYINPUT116), .Z(new_n1142));
  NAND2_X1  g0942(.A1(new_n730), .A2(G128), .ZN(new_n1143));
  AOI22_X1  g0943(.A1(new_n723), .A2(G150), .B1(new_n725), .B2(G137), .ZN(new_n1144));
  AOI22_X1  g0944(.A1(new_n738), .A2(G125), .B1(new_n735), .B2(G132), .ZN(new_n1145));
  NAND4_X1  g0945(.A1(new_n1142), .A2(new_n1143), .A3(new_n1144), .A4(new_n1145), .ZN(new_n1146));
  XOR2_X1   g0946(.A(new_n1146), .B(KEYINPUT59), .Z(new_n1147));
  INV_X1    g0947(.A(G124), .ZN(new_n1148));
  OAI21_X1  g0948(.A(new_n1139), .B1(new_n715), .B2(new_n1148), .ZN(new_n1149));
  AOI21_X1  g0949(.A(new_n1149), .B1(G159), .B2(new_n718), .ZN(new_n1150));
  AOI21_X1  g0950(.A(new_n1140), .B1(new_n1147), .B2(new_n1150), .ZN(new_n1151));
  AOI21_X1  g0951(.A(new_n709), .B1(new_n1138), .B2(new_n1151), .ZN(new_n1152));
  NOR2_X1   g0952(.A1(new_n809), .A2(new_n201), .ZN(new_n1153));
  NOR4_X1   g0953(.A1(new_n1130), .A2(new_n782), .A3(new_n1152), .A4(new_n1153), .ZN(new_n1154));
  NOR3_X1   g0954(.A1(new_n1111), .A2(new_n1114), .A3(KEYINPUT119), .ZN(new_n1155));
  AOI21_X1  g0955(.A(new_n1118), .B1(new_n1117), .B2(new_n1119), .ZN(new_n1156));
  NOR2_X1   g0956(.A1(new_n1155), .A2(new_n1156), .ZN(new_n1157));
  AOI21_X1  g0957(.A(new_n1154), .B1(new_n1157), .B2(new_n905), .ZN(new_n1158));
  NAND2_X1  g0958(.A1(new_n1129), .A2(new_n1158), .ZN(G375));
  NAND2_X1  g0959(.A1(new_n1048), .A2(new_n1049), .ZN(new_n1160));
  NOR2_X1   g0960(.A1(new_n1080), .A2(new_n1160), .ZN(new_n1161));
  INV_X1    g0961(.A(new_n1161), .ZN(new_n1162));
  NAND3_X1  g0962(.A1(new_n1162), .A2(new_n917), .A3(new_n1051), .ZN(new_n1163));
  AOI22_X1  g0963(.A1(new_n716), .A2(G128), .B1(new_n735), .B2(new_n1069), .ZN(new_n1164));
  AOI21_X1  g0964(.A(new_n1134), .B1(G132), .B2(new_n738), .ZN(new_n1165));
  OAI211_X1 g0965(.A(new_n1164), .B(new_n1165), .C1(new_n925), .C2(new_n724), .ZN(new_n1166));
  NOR2_X1   g0966(.A1(new_n731), .A2(new_n789), .ZN(new_n1167));
  NOR2_X1   g0967(.A1(new_n740), .A2(new_n380), .ZN(new_n1168));
  OAI21_X1  g0968(.A(new_n271), .B1(new_n722), .B2(new_n249), .ZN(new_n1169));
  NOR4_X1   g0969(.A1(new_n1166), .A2(new_n1167), .A3(new_n1168), .A4(new_n1169), .ZN(new_n1170));
  OAI22_X1  g0970(.A1(new_n724), .A2(new_n217), .B1(new_n734), .B2(new_n455), .ZN(new_n1171));
  XNOR2_X1  g0971(.A(new_n1171), .B(KEYINPUT121), .ZN(new_n1172));
  OAI221_X1 g0972(.A(new_n1172), .B1(new_n206), .B2(new_n717), .C1(new_n938), .C2(new_n731), .ZN(new_n1173));
  NOR2_X1   g0973(.A1(new_n749), .A2(new_n798), .ZN(new_n1174));
  NOR2_X1   g0974(.A1(new_n740), .A2(new_n438), .ZN(new_n1175));
  OAI211_X1 g0975(.A(new_n372), .B(new_n952), .C1(new_n715), .C2(new_n804), .ZN(new_n1176));
  NOR4_X1   g0976(.A1(new_n1173), .A2(new_n1174), .A3(new_n1175), .A4(new_n1176), .ZN(new_n1177));
  OAI21_X1  g0977(.A(new_n708), .B1(new_n1170), .B2(new_n1177), .ZN(new_n1178));
  OAI211_X1 g0978(.A(new_n768), .B(new_n1178), .C1(new_n821), .C2(new_n755), .ZN(new_n1179));
  AOI21_X1  g0979(.A(new_n1179), .B1(new_n203), .B2(new_n808), .ZN(new_n1180));
  AOI21_X1  g0980(.A(new_n1180), .B1(new_n1160), .B2(new_n905), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n1163), .A2(new_n1181), .ZN(G381));
  OR2_X1    g0982(.A1(G387), .A2(G390), .ZN(new_n1183));
  INV_X1    g0983(.A(G384), .ZN(new_n1184));
  NAND3_X1  g0984(.A1(new_n1163), .A2(new_n1184), .A3(new_n1181), .ZN(new_n1185));
  NOR4_X1   g0985(.A1(new_n1183), .A2(G396), .A3(G393), .A4(new_n1185), .ZN(new_n1186));
  NOR2_X1   g0986(.A1(G375), .A2(G378), .ZN(new_n1187));
  NAND2_X1  g0987(.A1(new_n1186), .A2(new_n1187), .ZN(G407));
  OAI21_X1  g0988(.A(new_n1187), .B1(new_n1186), .B2(new_n642), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n1189), .A2(G213), .ZN(G409));
  NAND2_X1  g0990(.A1(G387), .A2(G390), .ZN(new_n1191));
  NAND2_X1  g0991(.A1(new_n1183), .A2(new_n1191), .ZN(new_n1192));
  XOR2_X1   g0992(.A(G393), .B(G396), .Z(new_n1193));
  NAND2_X1  g0993(.A1(new_n1192), .A2(new_n1193), .ZN(new_n1194));
  INV_X1    g0994(.A(new_n1193), .ZN(new_n1195));
  NAND3_X1  g0995(.A1(new_n1183), .A2(new_n1195), .A3(new_n1191), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(new_n1194), .A2(new_n1196), .ZN(new_n1197));
  NAND3_X1  g0997(.A1(new_n1129), .A2(G378), .A3(new_n1158), .ZN(new_n1198));
  NAND4_X1  g0998(.A1(new_n1124), .A2(new_n917), .A3(new_n1115), .A4(new_n1120), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n1199), .A2(KEYINPUT122), .ZN(new_n1200));
  OR2_X1    g1000(.A1(new_n1125), .A2(KEYINPUT123), .ZN(new_n1201));
  AOI21_X1  g1001(.A(new_n904), .B1(new_n1125), .B2(KEYINPUT123), .ZN(new_n1202));
  AOI21_X1  g1002(.A(new_n1154), .B1(new_n1201), .B2(new_n1202), .ZN(new_n1203));
  INV_X1    g1003(.A(KEYINPUT122), .ZN(new_n1204));
  NAND4_X1  g1004(.A1(new_n1157), .A2(new_n1204), .A3(new_n917), .A4(new_n1124), .ZN(new_n1205));
  NAND3_X1  g1005(.A1(new_n1200), .A2(new_n1203), .A3(new_n1205), .ZN(new_n1206));
  INV_X1    g1006(.A(G378), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n1206), .A2(new_n1207), .ZN(new_n1208));
  NAND2_X1  g1008(.A1(new_n1208), .A2(KEYINPUT124), .ZN(new_n1209));
  INV_X1    g1009(.A(KEYINPUT124), .ZN(new_n1210));
  NAND3_X1  g1010(.A1(new_n1206), .A2(new_n1207), .A3(new_n1210), .ZN(new_n1211));
  NAND3_X1  g1011(.A1(new_n1198), .A2(new_n1209), .A3(new_n1211), .ZN(new_n1212));
  NAND2_X1  g1012(.A1(new_n642), .A2(G213), .ZN(new_n1213));
  AOI21_X1  g1013(.A(new_n663), .B1(new_n1161), .B2(KEYINPUT60), .ZN(new_n1214));
  OAI211_X1 g1014(.A(new_n1214), .B(new_n1051), .C1(KEYINPUT60), .C2(new_n1161), .ZN(new_n1215));
  INV_X1    g1015(.A(KEYINPUT125), .ZN(new_n1216));
  AOI22_X1  g1016(.A1(new_n1215), .A2(new_n1181), .B1(new_n1216), .B2(G384), .ZN(new_n1217));
  NOR2_X1   g1017(.A1(G384), .A2(new_n1216), .ZN(new_n1218));
  INV_X1    g1018(.A(new_n1218), .ZN(new_n1219));
  XNOR2_X1  g1019(.A(new_n1217), .B(new_n1219), .ZN(new_n1220));
  NAND3_X1  g1020(.A1(new_n1212), .A2(new_n1213), .A3(new_n1220), .ZN(new_n1221));
  INV_X1    g1021(.A(KEYINPUT126), .ZN(new_n1222));
  NAND2_X1  g1022(.A1(new_n1221), .A2(new_n1222), .ZN(new_n1223));
  NAND4_X1  g1023(.A1(new_n1212), .A2(KEYINPUT126), .A3(new_n1213), .A4(new_n1220), .ZN(new_n1224));
  AOI21_X1  g1024(.A(KEYINPUT62), .B1(new_n1223), .B2(new_n1224), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(new_n1212), .A2(new_n1213), .ZN(new_n1226));
  AND3_X1   g1026(.A1(new_n642), .A2(G213), .A3(G2897), .ZN(new_n1227));
  XNOR2_X1  g1027(.A(new_n1220), .B(new_n1227), .ZN(new_n1228));
  AOI21_X1  g1028(.A(KEYINPUT61), .B1(new_n1226), .B2(new_n1228), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n1221), .A2(KEYINPUT62), .ZN(new_n1230));
  NAND2_X1  g1030(.A1(new_n1229), .A2(new_n1230), .ZN(new_n1231));
  OAI21_X1  g1031(.A(new_n1197), .B1(new_n1225), .B2(new_n1231), .ZN(new_n1232));
  INV_X1    g1032(.A(KEYINPUT63), .ZN(new_n1233));
  NAND3_X1  g1033(.A1(new_n1223), .A2(new_n1233), .A3(new_n1224), .ZN(new_n1234));
  AND2_X1   g1034(.A1(new_n1194), .A2(new_n1196), .ZN(new_n1235));
  OR2_X1    g1035(.A1(new_n1221), .A2(new_n1233), .ZN(new_n1236));
  NAND4_X1  g1036(.A1(new_n1234), .A2(new_n1235), .A3(new_n1229), .A4(new_n1236), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(new_n1232), .A2(new_n1237), .ZN(G405));
  INV_X1    g1038(.A(KEYINPUT127), .ZN(new_n1239));
  AOI21_X1  g1039(.A(new_n1207), .B1(new_n1129), .B2(new_n1158), .ZN(new_n1240));
  NOR2_X1   g1040(.A1(new_n1187), .A2(new_n1240), .ZN(new_n1241));
  OAI21_X1  g1041(.A(new_n1235), .B1(new_n1239), .B2(new_n1241), .ZN(new_n1242));
  OAI211_X1 g1042(.A(new_n1197), .B(KEYINPUT127), .C1(new_n1187), .C2(new_n1240), .ZN(new_n1243));
  AOI21_X1  g1043(.A(new_n1220), .B1(new_n1241), .B2(new_n1239), .ZN(new_n1244));
  AND3_X1   g1044(.A1(new_n1242), .A2(new_n1243), .A3(new_n1244), .ZN(new_n1245));
  AOI21_X1  g1045(.A(new_n1244), .B1(new_n1242), .B2(new_n1243), .ZN(new_n1246));
  NOR2_X1   g1046(.A1(new_n1245), .A2(new_n1246), .ZN(G402));
endmodule


