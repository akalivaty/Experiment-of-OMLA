

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359,
         n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370,
         n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381,
         n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392,
         n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403,
         n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414,
         n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425,
         n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436,
         n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447,
         n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458,
         n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469,
         n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480,
         n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491,
         n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502,
         n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513,
         n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601,
         n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612,
         n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623,
         n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634,
         n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645,
         n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656,
         n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667,
         n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678,
         n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689,
         n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700,
         n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711,
         n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722,
         n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733,
         n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744,
         n745, n746, n747, n748;

  OR2_X2 U372 ( .A1(n598), .A2(n616), .ZN(n546) );
  XNOR2_X2 U373 ( .A(n529), .B(KEYINPUT33), .ZN(n619) );
  NAND2_X2 U374 ( .A1(n626), .A2(n625), .ZN(n627) );
  XNOR2_X2 U375 ( .A(n624), .B(KEYINPUT35), .ZN(n625) );
  XNOR2_X2 U376 ( .A(n555), .B(n517), .ZN(n373) );
  AND2_X1 U377 ( .A1(n700), .A2(n362), .ZN(n694) );
  NAND2_X1 U378 ( .A1(n657), .A2(n728), .ZN(n701) );
  NAND2_X1 U379 ( .A1(n659), .A2(n658), .ZN(n700) );
  NOR2_X1 U380 ( .A1(n654), .A2(n653), .ZN(n656) );
  XNOR2_X1 U381 ( .A(n419), .B(n418), .ZN(n593) );
  BUF_X1 U382 ( .A(n528), .Z(n637) );
  XNOR2_X1 U383 ( .A(n450), .B(KEYINPUT66), .ZN(n480) );
  XNOR2_X1 U384 ( .A(G131), .B(KEYINPUT67), .ZN(n450) );
  XOR2_X1 U385 ( .A(G146), .B(G125), .Z(n466) );
  OR2_X1 U386 ( .A1(n654), .A2(n653), .ZN(n735) );
  OR2_X1 U387 ( .A1(G237), .A2(G902), .ZN(n475) );
  XNOR2_X1 U388 ( .A(n489), .B(n488), .ZN(n528) );
  NOR2_X1 U389 ( .A1(G902), .A2(n662), .ZN(n489) );
  XNOR2_X1 U390 ( .A(G902), .B(KEYINPUT15), .ZN(n708) );
  XNOR2_X1 U391 ( .A(n385), .B(n384), .ZN(n586) );
  INV_X1 U392 ( .A(KEYINPUT46), .ZN(n384) );
  NAND2_X1 U393 ( .A1(n377), .A2(n376), .ZN(n385) );
  AND2_X1 U394 ( .A1(n378), .A2(n383), .ZN(n377) );
  INV_X1 U395 ( .A(n551), .ZN(n421) );
  XNOR2_X1 U396 ( .A(n528), .B(n527), .ZN(n562) );
  AND2_X1 U397 ( .A1(n410), .A2(n409), .ZN(n414) );
  NAND2_X1 U398 ( .A1(n413), .A2(n412), .ZN(n411) );
  AND2_X1 U399 ( .A1(n549), .A2(n577), .ZN(n550) );
  XNOR2_X1 U400 ( .A(n474), .B(KEYINPUT91), .ZN(n418) );
  NAND2_X1 U401 ( .A1(n695), .A2(n708), .ZN(n419) );
  XNOR2_X1 U402 ( .A(n399), .B(KEYINPUT72), .ZN(n573) );
  OR2_X1 U403 ( .A1(n639), .A2(n400), .ZN(n399) );
  INV_X1 U404 ( .A(KEYINPUT47), .ZN(n401) );
  INV_X1 U405 ( .A(n690), .ZN(n584) );
  XNOR2_X1 U406 ( .A(n404), .B(n455), .ZN(n709) );
  XNOR2_X1 U407 ( .A(n734), .B(n405), .ZN(n404) );
  NOR2_X1 U408 ( .A1(G902), .A2(n703), .ZN(n516) );
  XNOR2_X1 U409 ( .A(n371), .B(n487), .ZN(n662) );
  XOR2_X1 U410 ( .A(KEYINPUT23), .B(KEYINPUT24), .Z(n492) );
  AND2_X1 U411 ( .A1(n428), .A2(n431), .ZN(n427) );
  AND2_X1 U412 ( .A1(n710), .A2(n363), .ZN(n428) );
  NAND2_X1 U413 ( .A1(n701), .A2(n700), .ZN(n396) );
  INV_X1 U414 ( .A(n722), .ZN(n431) );
  NAND2_X1 U415 ( .A1(n565), .A2(n568), .ZN(n588) );
  XNOR2_X1 U416 ( .A(n499), .B(KEYINPUT25), .ZN(n392) );
  OR2_X2 U417 ( .A1(n718), .A2(G902), .ZN(n393) );
  INV_X1 U418 ( .A(n562), .ZN(n631) );
  NOR2_X1 U419 ( .A1(n615), .A2(n614), .ZN(n629) );
  AND2_X1 U420 ( .A1(n700), .A2(n361), .ZN(n661) );
  XNOR2_X1 U421 ( .A(n723), .B(n372), .ZN(n695) );
  XNOR2_X1 U422 ( .A(n473), .B(n467), .ZN(n372) );
  XNOR2_X1 U423 ( .A(n466), .B(n465), .ZN(n467) );
  NOR2_X1 U424 ( .A1(G952), .A2(n736), .ZN(n722) );
  XNOR2_X1 U425 ( .A(n735), .B(KEYINPUT82), .ZN(n389) );
  AND2_X1 U426 ( .A1(n646), .A2(n388), .ZN(n387) );
  NOR2_X1 U427 ( .A1(n648), .A2(n352), .ZN(n388) );
  NAND2_X1 U428 ( .A1(n381), .A2(n380), .ZN(n376) );
  NAND2_X1 U429 ( .A1(n397), .A2(n575), .ZN(n682) );
  INV_X1 U430 ( .A(n574), .ZN(n397) );
  INV_X1 U431 ( .A(n681), .ZN(n402) );
  XNOR2_X1 U432 ( .A(n532), .B(n403), .ZN(n639) );
  INV_X1 U433 ( .A(KEYINPUT102), .ZN(n403) );
  XNOR2_X1 U434 ( .A(n458), .B(n406), .ZN(n405) );
  XNOR2_X1 U435 ( .A(n354), .B(n454), .ZN(n406) );
  NOR2_X1 U436 ( .A1(G953), .A2(G237), .ZN(n485) );
  XNOR2_X1 U437 ( .A(G119), .B(G146), .ZN(n483) );
  XNOR2_X1 U438 ( .A(n368), .B(n359), .ZN(n654) );
  INV_X1 U439 ( .A(KEYINPUT105), .ZN(n375) );
  NOR2_X1 U440 ( .A1(n373), .A2(n546), .ZN(n526) );
  XNOR2_X1 U441 ( .A(KEYINPUT69), .B(n463), .ZN(n486) );
  XNOR2_X1 U442 ( .A(G143), .B(G128), .ZN(n468) );
  XNOR2_X1 U443 ( .A(G116), .B(G134), .ZN(n441) );
  XOR2_X1 U444 ( .A(G122), .B(G107), .Z(n442) );
  XNOR2_X1 U445 ( .A(n511), .B(G140), .ZN(n513) );
  XOR2_X1 U446 ( .A(G101), .B(G104), .Z(n512) );
  XNOR2_X1 U447 ( .A(n507), .B(n433), .ZN(n733) );
  INV_X1 U448 ( .A(KEYINPUT94), .ZN(n433) );
  XNOR2_X1 U449 ( .A(n468), .B(KEYINPUT4), .ZN(n479) );
  XOR2_X1 U450 ( .A(KEYINPUT17), .B(KEYINPUT18), .Z(n470) );
  AND2_X1 U451 ( .A1(n420), .A2(n351), .ZN(n577) );
  XNOR2_X1 U452 ( .A(n390), .B(n547), .ZN(n420) );
  INV_X1 U453 ( .A(KEYINPUT28), .ZN(n365) );
  XNOR2_X1 U454 ( .A(n457), .B(n398), .ZN(n574) );
  XNOR2_X1 U455 ( .A(n456), .B(G475), .ZN(n398) );
  NOR2_X1 U456 ( .A1(n546), .A2(n555), .ZN(n635) );
  XNOR2_X1 U457 ( .A(n408), .B(n407), .ZN(n634) );
  INV_X1 U458 ( .A(KEYINPUT0), .ZN(n407) );
  XNOR2_X1 U459 ( .A(G128), .B(G137), .ZN(n495) );
  AND2_X1 U460 ( .A1(n426), .A2(n425), .ZN(n424) );
  NAND2_X1 U461 ( .A1(n349), .A2(n431), .ZN(n425) );
  XNOR2_X1 U462 ( .A(n733), .B(n432), .ZN(n703) );
  XNOR2_X1 U463 ( .A(n510), .B(n514), .ZN(n432) );
  XNOR2_X1 U464 ( .A(n513), .B(n512), .ZN(n514) );
  XNOR2_X1 U465 ( .A(n509), .B(G110), .ZN(n510) );
  XNOR2_X1 U466 ( .A(n591), .B(n590), .ZN(n592) );
  XNOR2_X1 U467 ( .A(KEYINPUT43), .B(KEYINPUT108), .ZN(n590) );
  AND2_X1 U468 ( .A1(n370), .A2(n369), .ZN(n690) );
  INV_X1 U469 ( .A(n609), .ZN(n369) );
  NOR2_X1 U470 ( .A1(n631), .A2(n610), .ZN(n611) );
  NOR2_X1 U471 ( .A1(n637), .A2(n617), .ZN(n677) );
  INV_X1 U472 ( .A(n682), .ZN(n684) );
  NOR2_X1 U473 ( .A1(n667), .A2(n722), .ZN(n366) );
  NOR2_X1 U474 ( .A1(n698), .A2(n722), .ZN(n699) );
  XNOR2_X1 U475 ( .A(n695), .B(n434), .ZN(n696) );
  XNOR2_X1 U476 ( .A(n386), .B(n652), .ZN(G75) );
  NAND2_X1 U477 ( .A1(n647), .A2(n387), .ZN(n386) );
  NAND2_X1 U478 ( .A1(n357), .A2(n376), .ZN(n744) );
  NOR2_X1 U479 ( .A1(n710), .A2(n363), .ZN(n349) );
  AND2_X1 U480 ( .A1(n701), .A2(n394), .ZN(n350) );
  XOR2_X1 U481 ( .A(KEYINPUT30), .B(n548), .Z(n351) );
  OR2_X1 U482 ( .A1(G953), .A2(n651), .ZN(n352) );
  XOR2_X1 U483 ( .A(n484), .B(n483), .Z(n353) );
  XOR2_X1 U484 ( .A(G113), .B(G143), .Z(n354) );
  AND2_X1 U485 ( .A1(n396), .A2(n430), .ZN(n355) );
  AND2_X1 U486 ( .A1(n627), .A2(n642), .ZN(n356) );
  AND2_X1 U487 ( .A1(n383), .A2(n382), .ZN(n357) );
  XOR2_X1 U488 ( .A(KEYINPUT112), .B(KEYINPUT40), .Z(n358) );
  XOR2_X1 U489 ( .A(KEYINPUT48), .B(KEYINPUT83), .Z(n359) );
  XNOR2_X1 U490 ( .A(KEYINPUT59), .B(KEYINPUT89), .ZN(n360) );
  NOR2_X1 U491 ( .A1(n660), .A2(n708), .ZN(n361) );
  NOR2_X1 U492 ( .A1(n693), .A2(n708), .ZN(n362) );
  NOR2_X1 U493 ( .A1(n708), .A2(n707), .ZN(n363) );
  AND2_X1 U494 ( .A1(n626), .A2(KEYINPUT84), .ZN(n364) );
  XNOR2_X1 U495 ( .A(n554), .B(n365), .ZN(n557) );
  XNOR2_X1 U496 ( .A(n507), .B(n353), .ZN(n371) );
  XNOR2_X1 U497 ( .A(n697), .B(n696), .ZN(n698) );
  NAND2_X1 U498 ( .A1(n402), .A2(n401), .ZN(n400) );
  INV_X1 U499 ( .A(n367), .ZN(n415) );
  NAND2_X1 U500 ( .A1(n416), .A2(n641), .ZN(n367) );
  XNOR2_X1 U501 ( .A(n366), .B(n668), .ZN(G57) );
  NAND2_X1 U502 ( .A1(n619), .A2(n634), .ZN(n621) );
  XNOR2_X1 U503 ( .A(n618), .B(n364), .ZN(n417) );
  NAND2_X1 U504 ( .A1(n367), .A2(n642), .ZN(n409) );
  NAND2_X1 U505 ( .A1(n585), .A2(n586), .ZN(n368) );
  XNOR2_X1 U506 ( .A(n567), .B(KEYINPUT36), .ZN(n370) );
  NAND2_X1 U507 ( .A1(n429), .A2(n427), .ZN(n426) );
  NOR2_X1 U508 ( .A1(n745), .A2(n379), .ZN(n378) );
  NAND2_X1 U509 ( .A1(n374), .A2(n631), .ZN(n529) );
  XNOR2_X1 U510 ( .A(n526), .B(n375), .ZN(n374) );
  XNOR2_X1 U511 ( .A(n481), .B(n482), .ZN(n507) );
  INV_X1 U512 ( .A(n382), .ZN(n379) );
  NOR2_X1 U513 ( .A1(n682), .A2(n358), .ZN(n380) );
  INV_X1 U514 ( .A(n594), .ZN(n381) );
  NAND2_X1 U515 ( .A1(n682), .A2(n358), .ZN(n382) );
  NAND2_X1 U516 ( .A1(n594), .A2(n358), .ZN(n383) );
  NOR2_X1 U517 ( .A1(n389), .A2(KEYINPUT2), .ZN(n643) );
  NAND2_X1 U518 ( .A1(n391), .A2(n421), .ZN(n390) );
  XNOR2_X1 U519 ( .A(n635), .B(n422), .ZN(n391) );
  XNOR2_X2 U520 ( .A(n393), .B(n392), .ZN(n616) );
  AND2_X1 U521 ( .A1(n700), .A2(n395), .ZN(n394) );
  INV_X1 U522 ( .A(n708), .ZN(n395) );
  INV_X1 U523 ( .A(n396), .ZN(n429) );
  XNOR2_X2 U524 ( .A(n550), .B(KEYINPUT39), .ZN(n594) );
  XNOR2_X2 U525 ( .A(n449), .B(G140), .ZN(n734) );
  NAND2_X1 U526 ( .A1(n350), .A2(G478), .ZN(n715) );
  NAND2_X1 U527 ( .A1(n350), .A2(G217), .ZN(n719) );
  NAND2_X1 U528 ( .A1(n350), .A2(G469), .ZN(n705) );
  NAND2_X1 U529 ( .A1(n634), .A2(n607), .ZN(n608) );
  NAND2_X1 U530 ( .A1(n606), .A2(n605), .ZN(n408) );
  XNOR2_X1 U531 ( .A(n570), .B(n569), .ZN(n606) );
  NAND2_X1 U532 ( .A1(n417), .A2(n356), .ZN(n410) );
  NAND2_X2 U533 ( .A1(n414), .A2(n411), .ZN(n658) );
  NAND2_X1 U534 ( .A1(n417), .A2(n627), .ZN(n412) );
  AND2_X1 U535 ( .A1(n415), .A2(KEYINPUT45), .ZN(n413) );
  NAND2_X1 U536 ( .A1(n625), .A2(n627), .ZN(n416) );
  INV_X1 U537 ( .A(KEYINPUT109), .ZN(n422) );
  NAND2_X1 U538 ( .A1(n424), .A2(n423), .ZN(n713) );
  NAND2_X1 U539 ( .A1(n355), .A2(n431), .ZN(n423) );
  INV_X1 U540 ( .A(n710), .ZN(n430) );
  XNOR2_X1 U541 ( .A(n479), .B(n472), .ZN(n473) );
  AND2_X1 U542 ( .A1(n584), .A2(n583), .ZN(n585) );
  XNOR2_X1 U543 ( .A(KEYINPUT54), .B(KEYINPUT55), .ZN(n434) );
  AND2_X1 U544 ( .A1(n485), .A2(G210), .ZN(n435) );
  XNOR2_X1 U545 ( .A(n486), .B(n435), .ZN(n487) );
  INV_X1 U546 ( .A(G475), .ZN(n707) );
  INV_X1 U547 ( .A(KEYINPUT107), .ZN(n587) );
  XNOR2_X1 U548 ( .A(KEYINPUT1), .B(KEYINPUT64), .ZN(n517) );
  OR2_X1 U549 ( .A1(n692), .A2(n596), .ZN(n653) );
  XNOR2_X1 U550 ( .A(n476), .B(KEYINPUT113), .ZN(n477) );
  XNOR2_X1 U551 ( .A(n664), .B(n663), .ZN(n665) );
  XNOR2_X1 U552 ( .A(n709), .B(n360), .ZN(n710) );
  XNOR2_X1 U553 ( .A(n478), .B(n477), .ZN(n649) );
  XNOR2_X1 U554 ( .A(n666), .B(n665), .ZN(n667) );
  XNOR2_X1 U555 ( .A(KEYINPUT85), .B(KEYINPUT63), .ZN(n668) );
  NAND2_X1 U556 ( .A1(G234), .A2(G237), .ZN(n436) );
  XNOR2_X1 U557 ( .A(n436), .B(KEYINPUT14), .ZN(n542) );
  NAND2_X1 U558 ( .A1(G952), .A2(n542), .ZN(n541) );
  XOR2_X1 U559 ( .A(KEYINPUT100), .B(KEYINPUT7), .Z(n440) );
  INV_X2 U560 ( .A(G953), .ZN(n736) );
  NAND2_X1 U561 ( .A1(n736), .A2(G234), .ZN(n438) );
  XNOR2_X1 U562 ( .A(KEYINPUT81), .B(KEYINPUT8), .ZN(n437) );
  XNOR2_X1 U563 ( .A(n438), .B(n437), .ZN(n490) );
  NAND2_X1 U564 ( .A1(G217), .A2(n490), .ZN(n439) );
  XNOR2_X1 U565 ( .A(n440), .B(n439), .ZN(n446) );
  XNOR2_X1 U566 ( .A(n442), .B(n441), .ZN(n443) );
  XNOR2_X1 U567 ( .A(KEYINPUT9), .B(n443), .ZN(n444) );
  XNOR2_X1 U568 ( .A(n468), .B(n444), .ZN(n445) );
  XNOR2_X1 U569 ( .A(n446), .B(n445), .ZN(n714) );
  NOR2_X1 U570 ( .A1(G902), .A2(n714), .ZN(n447) );
  XOR2_X1 U571 ( .A(G478), .B(n447), .Z(n448) );
  XNOR2_X1 U572 ( .A(KEYINPUT101), .B(n448), .ZN(n575) );
  XNOR2_X1 U573 ( .A(n466), .B(KEYINPUT10), .ZN(n449) );
  XOR2_X1 U574 ( .A(KEYINPUT98), .B(KEYINPUT12), .Z(n452) );
  XNOR2_X1 U575 ( .A(KEYINPUT11), .B(KEYINPUT97), .ZN(n451) );
  XNOR2_X1 U576 ( .A(n452), .B(n451), .ZN(n453) );
  XOR2_X1 U577 ( .A(n480), .B(n453), .Z(n455) );
  NAND2_X1 U578 ( .A1(G214), .A2(n485), .ZN(n454) );
  XOR2_X1 U579 ( .A(G122), .B(G104), .Z(n458) );
  NOR2_X1 U580 ( .A1(G902), .A2(n709), .ZN(n457) );
  XNOR2_X1 U581 ( .A(KEYINPUT13), .B(KEYINPUT99), .ZN(n456) );
  NAND2_X1 U582 ( .A1(n575), .A2(n574), .ZN(n597) );
  XNOR2_X1 U583 ( .A(G119), .B(G110), .ZN(n494) );
  XNOR2_X1 U584 ( .A(KEYINPUT16), .B(n494), .ZN(n460) );
  XOR2_X1 U585 ( .A(G107), .B(KEYINPUT74), .Z(n508) );
  XNOR2_X1 U586 ( .A(n458), .B(n508), .ZN(n459) );
  XNOR2_X1 U587 ( .A(n460), .B(n459), .ZN(n464) );
  XOR2_X1 U588 ( .A(KEYINPUT3), .B(G116), .Z(n462) );
  XNOR2_X1 U589 ( .A(G113), .B(G101), .ZN(n461) );
  XNOR2_X1 U590 ( .A(n462), .B(n461), .ZN(n463) );
  XNOR2_X1 U591 ( .A(n464), .B(n486), .ZN(n723) );
  XOR2_X1 U592 ( .A(KEYINPUT90), .B(KEYINPUT78), .Z(n465) );
  NAND2_X1 U593 ( .A1(G224), .A2(n736), .ZN(n469) );
  XNOR2_X1 U594 ( .A(n470), .B(n469), .ZN(n471) );
  XNOR2_X1 U595 ( .A(KEYINPUT86), .B(n471), .ZN(n472) );
  NAND2_X1 U596 ( .A1(G210), .A2(n475), .ZN(n474) );
  XOR2_X1 U597 ( .A(KEYINPUT38), .B(n593), .Z(n549) );
  NAND2_X1 U598 ( .A1(G214), .A2(n475), .ZN(n568) );
  NAND2_X1 U599 ( .A1(n549), .A2(n568), .ZN(n533) );
  NOR2_X1 U600 ( .A1(n597), .A2(n533), .ZN(n478) );
  INV_X1 U601 ( .A(KEYINPUT41), .ZN(n476) );
  XNOR2_X1 U602 ( .A(n479), .B(G134), .ZN(n482) );
  XOR2_X1 U603 ( .A(G137), .B(n480), .Z(n481) );
  XOR2_X1 U604 ( .A(KEYINPUT73), .B(KEYINPUT5), .Z(n484) );
  XNOR2_X1 U605 ( .A(G472), .B(KEYINPUT71), .ZN(n488) );
  NAND2_X1 U606 ( .A1(G221), .A2(n490), .ZN(n491) );
  XNOR2_X1 U607 ( .A(n492), .B(n491), .ZN(n493) );
  XNOR2_X1 U608 ( .A(n734), .B(n493), .ZN(n497) );
  XNOR2_X1 U609 ( .A(n495), .B(n494), .ZN(n496) );
  XNOR2_X1 U610 ( .A(n497), .B(n496), .ZN(n718) );
  NAND2_X1 U611 ( .A1(G234), .A2(n708), .ZN(n498) );
  XNOR2_X1 U612 ( .A(KEYINPUT20), .B(n498), .ZN(n500) );
  NAND2_X1 U613 ( .A1(G217), .A2(n500), .ZN(n499) );
  XOR2_X1 U614 ( .A(KEYINPUT95), .B(KEYINPUT21), .Z(n502) );
  NAND2_X1 U615 ( .A1(G221), .A2(n500), .ZN(n501) );
  XNOR2_X1 U616 ( .A(n502), .B(n501), .ZN(n598) );
  NAND2_X1 U617 ( .A1(n616), .A2(n598), .ZN(n503) );
  XNOR2_X1 U618 ( .A(n503), .B(KEYINPUT120), .ZN(n504) );
  XNOR2_X1 U619 ( .A(n504), .B(KEYINPUT49), .ZN(n505) );
  NOR2_X1 U620 ( .A1(n637), .A2(n505), .ZN(n506) );
  XNOR2_X1 U621 ( .A(KEYINPUT121), .B(n506), .ZN(n520) );
  XOR2_X1 U622 ( .A(n508), .B(G146), .Z(n509) );
  AND2_X1 U623 ( .A1(G227), .A2(n736), .ZN(n511) );
  XNOR2_X1 U624 ( .A(KEYINPUT68), .B(G469), .ZN(n515) );
  XNOR2_X2 U625 ( .A(n516), .B(n515), .ZN(n555) );
  NAND2_X1 U626 ( .A1(n373), .A2(n546), .ZN(n518) );
  XOR2_X1 U627 ( .A(KEYINPUT50), .B(n518), .Z(n519) );
  NOR2_X1 U628 ( .A1(n520), .A2(n519), .ZN(n522) );
  NAND2_X1 U629 ( .A1(n526), .A2(n637), .ZN(n521) );
  XOR2_X1 U630 ( .A(KEYINPUT96), .B(n521), .Z(n632) );
  NOR2_X1 U631 ( .A1(n522), .A2(n632), .ZN(n523) );
  XOR2_X1 U632 ( .A(KEYINPUT51), .B(n523), .Z(n524) );
  NOR2_X1 U633 ( .A1(n649), .A2(n524), .ZN(n525) );
  XNOR2_X1 U634 ( .A(n525), .B(KEYINPUT122), .ZN(n538) );
  XOR2_X1 U635 ( .A(KEYINPUT6), .B(KEYINPUT103), .Z(n527) );
  INV_X1 U636 ( .A(n619), .ZN(n650) );
  NOR2_X1 U637 ( .A1(n549), .A2(n568), .ZN(n530) );
  NOR2_X1 U638 ( .A1(n597), .A2(n530), .ZN(n535) );
  INV_X1 U639 ( .A(n575), .ZN(n531) );
  NAND2_X1 U640 ( .A1(n531), .A2(n574), .ZN(n678) );
  NAND2_X1 U641 ( .A1(n682), .A2(n678), .ZN(n532) );
  NOR2_X1 U642 ( .A1(n533), .A2(n639), .ZN(n534) );
  NOR2_X1 U643 ( .A1(n535), .A2(n534), .ZN(n536) );
  NOR2_X1 U644 ( .A1(n650), .A2(n536), .ZN(n537) );
  NOR2_X1 U645 ( .A1(n538), .A2(n537), .ZN(n539) );
  XNOR2_X1 U646 ( .A(n539), .B(KEYINPUT52), .ZN(n540) );
  NOR2_X1 U647 ( .A1(n541), .A2(n540), .ZN(n648) );
  INV_X1 U648 ( .A(KEYINPUT76), .ZN(n547) );
  NOR2_X1 U649 ( .A1(G953), .A2(n541), .ZN(n601) );
  NAND2_X1 U650 ( .A1(n542), .A2(G902), .ZN(n543) );
  XOR2_X1 U651 ( .A(KEYINPUT92), .B(n543), .Z(n600) );
  NAND2_X1 U652 ( .A1(n600), .A2(G953), .ZN(n544) );
  NOR2_X1 U653 ( .A1(G900), .A2(n544), .ZN(n545) );
  NOR2_X1 U654 ( .A1(n601), .A2(n545), .ZN(n551) );
  NAND2_X1 U655 ( .A1(n637), .A2(n568), .ZN(n548) );
  INV_X1 U656 ( .A(n637), .ZN(n553) );
  NOR2_X1 U657 ( .A1(n598), .A2(n551), .ZN(n552) );
  NAND2_X1 U658 ( .A1(n616), .A2(n552), .ZN(n561) );
  NOR2_X1 U659 ( .A1(n553), .A2(n561), .ZN(n554) );
  XOR2_X1 U660 ( .A(n555), .B(KEYINPUT111), .Z(n556) );
  NOR2_X1 U661 ( .A1(n557), .A2(n556), .ZN(n571) );
  INV_X1 U662 ( .A(n571), .ZN(n558) );
  NOR2_X1 U663 ( .A1(n649), .A2(n558), .ZN(n560) );
  XNOR2_X1 U664 ( .A(KEYINPUT114), .B(KEYINPUT42), .ZN(n559) );
  XNOR2_X1 U665 ( .A(n560), .B(n559), .ZN(n745) );
  XNOR2_X1 U666 ( .A(n373), .B(KEYINPUT88), .ZN(n609) );
  INV_X1 U667 ( .A(n593), .ZN(n566) );
  NOR2_X1 U668 ( .A1(n562), .A2(n561), .ZN(n563) );
  XOR2_X1 U669 ( .A(KEYINPUT106), .B(n563), .Z(n564) );
  NOR2_X1 U670 ( .A1(n682), .A2(n564), .ZN(n565) );
  NOR2_X1 U671 ( .A1(n566), .A2(n588), .ZN(n567) );
  NAND2_X1 U672 ( .A1(n593), .A2(n568), .ZN(n570) );
  XOR2_X1 U673 ( .A(KEYINPUT77), .B(KEYINPUT19), .Z(n569) );
  NAND2_X1 U674 ( .A1(n606), .A2(n571), .ZN(n681) );
  NAND2_X1 U675 ( .A1(n681), .A2(KEYINPUT47), .ZN(n572) );
  NAND2_X1 U676 ( .A1(n573), .A2(n572), .ZN(n582) );
  NOR2_X1 U677 ( .A1(n575), .A2(n574), .ZN(n622) );
  AND2_X1 U678 ( .A1(n622), .A2(n593), .ZN(n576) );
  NAND2_X1 U679 ( .A1(n577), .A2(n576), .ZN(n578) );
  XNOR2_X1 U680 ( .A(KEYINPUT110), .B(n578), .ZN(n747) );
  NAND2_X1 U681 ( .A1(KEYINPUT47), .A2(n639), .ZN(n579) );
  NAND2_X1 U682 ( .A1(n747), .A2(n579), .ZN(n580) );
  XNOR2_X1 U683 ( .A(KEYINPUT80), .B(n580), .ZN(n581) );
  NOR2_X1 U684 ( .A1(n582), .A2(n581), .ZN(n583) );
  INV_X1 U685 ( .A(n373), .ZN(n614) );
  XNOR2_X1 U686 ( .A(n588), .B(n587), .ZN(n589) );
  NOR2_X1 U687 ( .A1(n614), .A2(n589), .ZN(n591) );
  NOR2_X1 U688 ( .A1(n593), .A2(n592), .ZN(n692) );
  NOR2_X1 U689 ( .A1(n594), .A2(n678), .ZN(n595) );
  XNOR2_X1 U690 ( .A(n595), .B(KEYINPUT115), .ZN(n743) );
  INV_X1 U691 ( .A(n743), .ZN(n596) );
  NOR2_X1 U692 ( .A1(n598), .A2(n597), .ZN(n599) );
  XNOR2_X1 U693 ( .A(KEYINPUT104), .B(n599), .ZN(n607) );
  NOR2_X1 U694 ( .A1(G898), .A2(n736), .ZN(n724) );
  NAND2_X1 U695 ( .A1(n724), .A2(n600), .ZN(n603) );
  INV_X1 U696 ( .A(n601), .ZN(n602) );
  NAND2_X1 U697 ( .A1(n603), .A2(n602), .ZN(n604) );
  XOR2_X1 U698 ( .A(KEYINPUT93), .B(n604), .Z(n605) );
  XNOR2_X1 U699 ( .A(n608), .B(KEYINPUT22), .ZN(n615) );
  INV_X1 U700 ( .A(n616), .ZN(n628) );
  OR2_X1 U701 ( .A1(n628), .A2(n609), .ZN(n610) );
  XNOR2_X1 U702 ( .A(n611), .B(KEYINPUT79), .ZN(n612) );
  NOR2_X1 U703 ( .A1(n615), .A2(n612), .ZN(n613) );
  XNOR2_X1 U704 ( .A(KEYINPUT32), .B(n613), .ZN(n748) );
  NAND2_X1 U705 ( .A1(n616), .A2(n629), .ZN(n617) );
  NOR2_X1 U706 ( .A1(n748), .A2(n677), .ZN(n618) );
  INV_X1 U707 ( .A(KEYINPUT44), .ZN(n626) );
  XOR2_X1 U708 ( .A(KEYINPUT70), .B(KEYINPUT34), .Z(n620) );
  XNOR2_X1 U709 ( .A(n621), .B(n620), .ZN(n623) );
  NAND2_X1 U710 ( .A1(n623), .A2(n622), .ZN(n624) );
  INV_X1 U711 ( .A(n625), .ZN(n746) );
  NAND2_X1 U712 ( .A1(n629), .A2(n628), .ZN(n630) );
  NOR2_X1 U713 ( .A1(n631), .A2(n630), .ZN(n669) );
  NAND2_X1 U714 ( .A1(n632), .A2(n634), .ZN(n633) );
  XNOR2_X1 U715 ( .A(n633), .B(KEYINPUT31), .ZN(n687) );
  NAND2_X1 U716 ( .A1(n635), .A2(n634), .ZN(n636) );
  NOR2_X1 U717 ( .A1(n637), .A2(n636), .ZN(n672) );
  NOR2_X1 U718 ( .A1(n687), .A2(n672), .ZN(n638) );
  NOR2_X1 U719 ( .A1(n639), .A2(n638), .ZN(n640) );
  NOR2_X1 U720 ( .A1(n669), .A2(n640), .ZN(n641) );
  INV_X1 U721 ( .A(KEYINPUT45), .ZN(n642) );
  INV_X1 U722 ( .A(n658), .ZN(n728) );
  NAND2_X1 U723 ( .A1(n643), .A2(n728), .ZN(n647) );
  INV_X1 U724 ( .A(KEYINPUT2), .ZN(n659) );
  NOR2_X1 U725 ( .A1(n658), .A2(n735), .ZN(n644) );
  NOR2_X1 U726 ( .A1(n659), .A2(n644), .ZN(n645) );
  NAND2_X1 U727 ( .A1(KEYINPUT82), .A2(n645), .ZN(n646) );
  NOR2_X1 U728 ( .A1(n650), .A2(n649), .ZN(n651) );
  XNOR2_X1 U729 ( .A(KEYINPUT123), .B(KEYINPUT53), .ZN(n652) );
  OR2_X1 U730 ( .A1(KEYINPUT2), .A2(KEYINPUT75), .ZN(n655) );
  XNOR2_X1 U731 ( .A(n656), .B(n655), .ZN(n657) );
  INV_X1 U732 ( .A(G472), .ZN(n660) );
  NAND2_X1 U733 ( .A1(n701), .A2(n661), .ZN(n666) );
  XNOR2_X1 U734 ( .A(n662), .B(KEYINPUT116), .ZN(n664) );
  XOR2_X1 U735 ( .A(KEYINPUT62), .B(KEYINPUT87), .Z(n663) );
  XOR2_X1 U736 ( .A(G101), .B(n669), .Z(G3) );
  XOR2_X1 U737 ( .A(G104), .B(KEYINPUT117), .Z(n671) );
  NAND2_X1 U738 ( .A1(n672), .A2(n684), .ZN(n670) );
  XNOR2_X1 U739 ( .A(n671), .B(n670), .ZN(G6) );
  XNOR2_X1 U740 ( .A(G107), .B(KEYINPUT27), .ZN(n676) );
  XOR2_X1 U741 ( .A(KEYINPUT118), .B(KEYINPUT26), .Z(n674) );
  INV_X1 U742 ( .A(n678), .ZN(n686) );
  NAND2_X1 U743 ( .A1(n672), .A2(n686), .ZN(n673) );
  XNOR2_X1 U744 ( .A(n674), .B(n673), .ZN(n675) );
  XNOR2_X1 U745 ( .A(n676), .B(n675), .ZN(G9) );
  XOR2_X1 U746 ( .A(G110), .B(n677), .Z(G12) );
  NOR2_X1 U747 ( .A1(n678), .A2(n681), .ZN(n680) );
  XNOR2_X1 U748 ( .A(G128), .B(KEYINPUT29), .ZN(n679) );
  XNOR2_X1 U749 ( .A(n680), .B(n679), .ZN(G30) );
  NOR2_X1 U750 ( .A1(n682), .A2(n681), .ZN(n683) );
  XOR2_X1 U751 ( .A(G146), .B(n683), .Z(G48) );
  NAND2_X1 U752 ( .A1(n684), .A2(n687), .ZN(n685) );
  XNOR2_X1 U753 ( .A(G113), .B(n685), .ZN(G15) );
  XOR2_X1 U754 ( .A(G116), .B(KEYINPUT119), .Z(n689) );
  NAND2_X1 U755 ( .A1(n687), .A2(n686), .ZN(n688) );
  XNOR2_X1 U756 ( .A(n689), .B(n688), .ZN(G18) );
  XNOR2_X1 U757 ( .A(n690), .B(G125), .ZN(n691) );
  XNOR2_X1 U758 ( .A(n691), .B(KEYINPUT37), .ZN(G27) );
  XOR2_X1 U759 ( .A(G140), .B(n692), .Z(G42) );
  INV_X1 U760 ( .A(G210), .ZN(n693) );
  NAND2_X1 U761 ( .A1(n701), .A2(n694), .ZN(n697) );
  XNOR2_X1 U762 ( .A(KEYINPUT56), .B(n699), .ZN(G51) );
  XOR2_X1 U763 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n702) );
  XNOR2_X1 U764 ( .A(n703), .B(n702), .ZN(n704) );
  XNOR2_X1 U765 ( .A(n705), .B(n704), .ZN(n706) );
  NOR2_X1 U766 ( .A1(n722), .A2(n706), .ZN(G54) );
  XOR2_X1 U767 ( .A(KEYINPUT124), .B(KEYINPUT60), .Z(n711) );
  XNOR2_X1 U768 ( .A(KEYINPUT65), .B(n711), .ZN(n712) );
  XNOR2_X1 U769 ( .A(n713), .B(n712), .ZN(G60) );
  XOR2_X1 U770 ( .A(n714), .B(KEYINPUT125), .Z(n716) );
  XNOR2_X1 U771 ( .A(n716), .B(n715), .ZN(n717) );
  NOR2_X1 U772 ( .A1(n722), .A2(n717), .ZN(G63) );
  XNOR2_X1 U773 ( .A(n718), .B(KEYINPUT126), .ZN(n720) );
  XNOR2_X1 U774 ( .A(n720), .B(n719), .ZN(n721) );
  NOR2_X1 U775 ( .A1(n722), .A2(n721), .ZN(G66) );
  NOR2_X1 U776 ( .A1(n724), .A2(n723), .ZN(n732) );
  XOR2_X1 U777 ( .A(KEYINPUT61), .B(KEYINPUT127), .Z(n726) );
  NAND2_X1 U778 ( .A1(G224), .A2(G953), .ZN(n725) );
  XNOR2_X1 U779 ( .A(n726), .B(n725), .ZN(n727) );
  NAND2_X1 U780 ( .A1(n727), .A2(G898), .ZN(n730) );
  NAND2_X1 U781 ( .A1(n728), .A2(n736), .ZN(n729) );
  NAND2_X1 U782 ( .A1(n730), .A2(n729), .ZN(n731) );
  XNOR2_X1 U783 ( .A(n732), .B(n731), .ZN(G69) );
  XOR2_X1 U784 ( .A(n733), .B(n734), .Z(n738) );
  XNOR2_X1 U785 ( .A(n735), .B(n738), .ZN(n737) );
  NAND2_X1 U786 ( .A1(n737), .A2(n736), .ZN(n742) );
  XNOR2_X1 U787 ( .A(G227), .B(n738), .ZN(n739) );
  NAND2_X1 U788 ( .A1(n739), .A2(G900), .ZN(n740) );
  NAND2_X1 U789 ( .A1(n740), .A2(G953), .ZN(n741) );
  NAND2_X1 U790 ( .A1(n742), .A2(n741), .ZN(G72) );
  XNOR2_X1 U791 ( .A(G134), .B(n743), .ZN(G36) );
  XOR2_X1 U792 ( .A(n744), .B(G131), .Z(G33) );
  XOR2_X1 U793 ( .A(G137), .B(n745), .Z(G39) );
  XNOR2_X1 U794 ( .A(n746), .B(G122), .ZN(G24) );
  XNOR2_X1 U795 ( .A(G143), .B(n747), .ZN(G45) );
  XOR2_X1 U796 ( .A(G119), .B(n748), .Z(G21) );
endmodule

