

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n514, n515, n516, n517,
         n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583,
         n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594,
         n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605,
         n606, n607, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
         n1023, n1024, n1025, n1026, n1027, n1028;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NOR2_X2 U550 ( .A1(n676), .A2(n675), .ZN(n698) );
  NOR2_X1 U551 ( .A1(n537), .A2(n536), .ZN(G160) );
  BUF_X1 U552 ( .A(n880), .Z(n514) );
  XNOR2_X1 U553 ( .A(n531), .B(n530), .ZN(n880) );
  NOR2_X1 U554 ( .A1(n641), .A2(n640), .ZN(n643) );
  NOR2_X1 U555 ( .A1(G543), .A2(n518), .ZN(n519) );
  NOR2_X1 U556 ( .A1(n522), .A2(n521), .ZN(n523) );
  NOR2_X1 U557 ( .A1(n690), .A2(n684), .ZN(n515) );
  INV_X1 U558 ( .A(KEYINPUT91), .ZN(n615) );
  XNOR2_X1 U559 ( .A(n616), .B(n615), .ZN(n617) );
  INV_X1 U560 ( .A(KEYINPUT28), .ZN(n632) );
  NOR2_X1 U561 ( .A1(n652), .A2(n651), .ZN(n653) );
  INV_X1 U562 ( .A(n979), .ZN(n680) );
  INV_X1 U563 ( .A(KEYINPUT32), .ZN(n666) );
  AND2_X1 U564 ( .A1(n681), .A2(n680), .ZN(n682) );
  NOR2_X1 U565 ( .A1(G1384), .A2(G164), .ZN(n609) );
  NAND2_X1 U566 ( .A1(n880), .A2(G138), .ZN(n541) );
  INV_X1 U567 ( .A(KEYINPUT17), .ZN(n530) );
  AND2_X1 U568 ( .A1(G2105), .A2(G2104), .ZN(n883) );
  NOR2_X1 U569 ( .A1(n577), .A2(G651), .ZN(n791) );
  NOR2_X1 U570 ( .A1(n545), .A2(n544), .ZN(G164) );
  XNOR2_X1 U571 ( .A(n525), .B(KEYINPUT70), .ZN(G299) );
  XOR2_X1 U572 ( .A(KEYINPUT0), .B(G543), .Z(n577) );
  NAND2_X1 U573 ( .A1(G53), .A2(n791), .ZN(n524) );
  NOR2_X1 U574 ( .A1(G543), .A2(G651), .ZN(n786) );
  NAND2_X1 U575 ( .A1(G91), .A2(n786), .ZN(n517) );
  XNOR2_X1 U576 ( .A(KEYINPUT67), .B(G651), .ZN(n518) );
  NOR2_X1 U577 ( .A1(n577), .A2(n518), .ZN(n787) );
  NAND2_X1 U578 ( .A1(G78), .A2(n787), .ZN(n516) );
  NAND2_X1 U579 ( .A1(n517), .A2(n516), .ZN(n522) );
  XOR2_X1 U580 ( .A(KEYINPUT1), .B(n519), .Z(n792) );
  NAND2_X1 U581 ( .A1(G65), .A2(n792), .ZN(n520) );
  XNOR2_X1 U582 ( .A(KEYINPUT69), .B(n520), .ZN(n521) );
  NAND2_X1 U583 ( .A1(n524), .A2(n523), .ZN(n525) );
  INV_X1 U584 ( .A(G2105), .ZN(n534) );
  NAND2_X1 U585 ( .A1(G113), .A2(n883), .ZN(n526) );
  XOR2_X1 U586 ( .A(KEYINPUT66), .B(n526), .Z(n529) );
  AND2_X1 U587 ( .A1(n534), .A2(G2104), .ZN(n879) );
  NAND2_X1 U588 ( .A1(G101), .A2(n879), .ZN(n527) );
  XNOR2_X1 U589 ( .A(KEYINPUT23), .B(n527), .ZN(n528) );
  NOR2_X1 U590 ( .A1(n529), .A2(n528), .ZN(n533) );
  NOR2_X1 U591 ( .A1(G2104), .A2(G2105), .ZN(n531) );
  NAND2_X1 U592 ( .A1(n514), .A2(G137), .ZN(n532) );
  NAND2_X1 U593 ( .A1(n533), .A2(n532), .ZN(n537) );
  NOR2_X1 U594 ( .A1(n534), .A2(G2104), .ZN(n885) );
  NAND2_X1 U595 ( .A1(G125), .A2(n885), .ZN(n535) );
  XNOR2_X1 U596 ( .A(KEYINPUT65), .B(n535), .ZN(n536) );
  NAND2_X1 U597 ( .A1(G114), .A2(n883), .ZN(n539) );
  NAND2_X1 U598 ( .A1(G126), .A2(n885), .ZN(n538) );
  NAND2_X1 U599 ( .A1(n539), .A2(n538), .ZN(n545) );
  INV_X1 U600 ( .A(KEYINPUT81), .ZN(n543) );
  NAND2_X1 U601 ( .A1(G102), .A2(n879), .ZN(n540) );
  NAND2_X1 U602 ( .A1(n541), .A2(n540), .ZN(n542) );
  XNOR2_X1 U603 ( .A(n543), .B(n542), .ZN(n544) );
  NAND2_X1 U604 ( .A1(n787), .A2(G73), .ZN(n546) );
  XNOR2_X1 U605 ( .A(n546), .B(KEYINPUT2), .ZN(n553) );
  NAND2_X1 U606 ( .A1(G86), .A2(n786), .ZN(n548) );
  NAND2_X1 U607 ( .A1(G48), .A2(n791), .ZN(n547) );
  NAND2_X1 U608 ( .A1(n548), .A2(n547), .ZN(n551) );
  NAND2_X1 U609 ( .A1(G61), .A2(n792), .ZN(n549) );
  XNOR2_X1 U610 ( .A(KEYINPUT77), .B(n549), .ZN(n550) );
  NOR2_X1 U611 ( .A1(n551), .A2(n550), .ZN(n552) );
  NAND2_X1 U612 ( .A1(n553), .A2(n552), .ZN(G305) );
  NAND2_X1 U613 ( .A1(G90), .A2(n786), .ZN(n555) );
  NAND2_X1 U614 ( .A1(G77), .A2(n787), .ZN(n554) );
  NAND2_X1 U615 ( .A1(n555), .A2(n554), .ZN(n556) );
  XNOR2_X1 U616 ( .A(KEYINPUT9), .B(n556), .ZN(n560) );
  NAND2_X1 U617 ( .A1(n792), .A2(G64), .ZN(n558) );
  NAND2_X1 U618 ( .A1(n791), .A2(G52), .ZN(n557) );
  AND2_X1 U619 ( .A1(n558), .A2(n557), .ZN(n559) );
  NAND2_X1 U620 ( .A1(n560), .A2(n559), .ZN(G301) );
  NAND2_X1 U621 ( .A1(n786), .A2(G89), .ZN(n561) );
  XNOR2_X1 U622 ( .A(n561), .B(KEYINPUT4), .ZN(n563) );
  NAND2_X1 U623 ( .A1(G76), .A2(n787), .ZN(n562) );
  NAND2_X1 U624 ( .A1(n563), .A2(n562), .ZN(n564) );
  XNOR2_X1 U625 ( .A(n564), .B(KEYINPUT5), .ZN(n569) );
  NAND2_X1 U626 ( .A1(n791), .A2(G51), .ZN(n566) );
  NAND2_X1 U627 ( .A1(G63), .A2(n792), .ZN(n565) );
  NAND2_X1 U628 ( .A1(n566), .A2(n565), .ZN(n567) );
  XOR2_X1 U629 ( .A(KEYINPUT6), .B(n567), .Z(n568) );
  NAND2_X1 U630 ( .A1(n569), .A2(n568), .ZN(n570) );
  XNOR2_X1 U631 ( .A(n570), .B(KEYINPUT7), .ZN(G168) );
  NAND2_X1 U632 ( .A1(G88), .A2(n786), .ZN(n572) );
  NAND2_X1 U633 ( .A1(G75), .A2(n787), .ZN(n571) );
  NAND2_X1 U634 ( .A1(n572), .A2(n571), .ZN(n576) );
  NAND2_X1 U635 ( .A1(n791), .A2(G50), .ZN(n574) );
  NAND2_X1 U636 ( .A1(G62), .A2(n792), .ZN(n573) );
  NAND2_X1 U637 ( .A1(n574), .A2(n573), .ZN(n575) );
  NOR2_X1 U638 ( .A1(n576), .A2(n575), .ZN(G166) );
  INV_X1 U639 ( .A(G166), .ZN(G303) );
  XOR2_X1 U640 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U641 ( .A1(G74), .A2(G651), .ZN(n579) );
  NAND2_X1 U642 ( .A1(G87), .A2(n577), .ZN(n578) );
  NAND2_X1 U643 ( .A1(n579), .A2(n578), .ZN(n580) );
  NOR2_X1 U644 ( .A1(n792), .A2(n580), .ZN(n582) );
  NAND2_X1 U645 ( .A1(n791), .A2(G49), .ZN(n581) );
  NAND2_X1 U646 ( .A1(n582), .A2(n581), .ZN(G288) );
  NAND2_X1 U647 ( .A1(n791), .A2(G47), .ZN(n584) );
  NAND2_X1 U648 ( .A1(G60), .A2(n792), .ZN(n583) );
  NAND2_X1 U649 ( .A1(n584), .A2(n583), .ZN(n585) );
  XOR2_X1 U650 ( .A(KEYINPUT68), .B(n585), .Z(n589) );
  NAND2_X1 U651 ( .A1(n787), .A2(G72), .ZN(n587) );
  NAND2_X1 U652 ( .A1(G85), .A2(n786), .ZN(n586) );
  AND2_X1 U653 ( .A1(n587), .A2(n586), .ZN(n588) );
  NAND2_X1 U654 ( .A1(n589), .A2(n588), .ZN(G290) );
  XNOR2_X1 U655 ( .A(G1981), .B(G305), .ZN(n975) );
  NAND2_X1 U656 ( .A1(n787), .A2(G79), .ZN(n596) );
  NAND2_X1 U657 ( .A1(n786), .A2(G92), .ZN(n591) );
  NAND2_X1 U658 ( .A1(G66), .A2(n792), .ZN(n590) );
  NAND2_X1 U659 ( .A1(n591), .A2(n590), .ZN(n594) );
  NAND2_X1 U660 ( .A1(n791), .A2(G54), .ZN(n592) );
  XOR2_X1 U661 ( .A(KEYINPUT72), .B(n592), .Z(n593) );
  NOR2_X1 U662 ( .A1(n594), .A2(n593), .ZN(n595) );
  NAND2_X1 U663 ( .A1(n596), .A2(n595), .ZN(n597) );
  XNOR2_X1 U664 ( .A(n597), .B(KEYINPUT15), .ZN(n966) );
  NAND2_X1 U665 ( .A1(n786), .A2(G81), .ZN(n598) );
  XNOR2_X1 U666 ( .A(n598), .B(KEYINPUT12), .ZN(n600) );
  NAND2_X1 U667 ( .A1(G68), .A2(n787), .ZN(n599) );
  NAND2_X1 U668 ( .A1(n600), .A2(n599), .ZN(n601) );
  XOR2_X1 U669 ( .A(KEYINPUT13), .B(n601), .Z(n605) );
  NAND2_X1 U670 ( .A1(n792), .A2(G56), .ZN(n602) );
  XNOR2_X1 U671 ( .A(n602), .B(KEYINPUT14), .ZN(n603) );
  XNOR2_X1 U672 ( .A(n603), .B(KEYINPUT71), .ZN(n604) );
  NOR2_X1 U673 ( .A1(n605), .A2(n604), .ZN(n607) );
  NAND2_X1 U674 ( .A1(n791), .A2(G43), .ZN(n606) );
  NAND2_X1 U675 ( .A1(n607), .A2(n606), .ZN(n967) );
  XNOR2_X1 U676 ( .A(G1996), .B(KEYINPUT90), .ZN(n942) );
  NAND2_X1 U677 ( .A1(G160), .A2(G40), .ZN(n706) );
  INV_X1 U678 ( .A(n706), .ZN(n612) );
  AND2_X1 U679 ( .A1(n942), .A2(n612), .ZN(n610) );
  XNOR2_X1 U680 ( .A(n609), .B(KEYINPUT64), .ZN(n705) );
  NAND2_X1 U681 ( .A1(n610), .A2(n705), .ZN(n611) );
  XNOR2_X1 U682 ( .A(n611), .B(KEYINPUT26), .ZN(n614) );
  NAND2_X1 U683 ( .A1(n705), .A2(n612), .ZN(n644) );
  NAND2_X1 U684 ( .A1(G1341), .A2(n644), .ZN(n613) );
  NAND2_X1 U685 ( .A1(n614), .A2(n613), .ZN(n616) );
  NOR2_X1 U686 ( .A1(n967), .A2(n617), .ZN(n618) );
  OR2_X1 U687 ( .A1(n966), .A2(n618), .ZN(n624) );
  NAND2_X1 U688 ( .A1(n966), .A2(n618), .ZN(n622) );
  INV_X1 U689 ( .A(n644), .ZN(n637) );
  NOR2_X1 U690 ( .A1(n637), .A2(G1348), .ZN(n620) );
  INV_X1 U691 ( .A(n637), .ZN(n654) );
  NOR2_X1 U692 ( .A1(G2067), .A2(n654), .ZN(n619) );
  NOR2_X1 U693 ( .A1(n620), .A2(n619), .ZN(n621) );
  NAND2_X1 U694 ( .A1(n622), .A2(n621), .ZN(n623) );
  NAND2_X1 U695 ( .A1(n624), .A2(n623), .ZN(n629) );
  NAND2_X1 U696 ( .A1(n637), .A2(G2072), .ZN(n625) );
  XNOR2_X1 U697 ( .A(n625), .B(KEYINPUT27), .ZN(n627) );
  INV_X1 U698 ( .A(G1956), .ZN(n916) );
  NOR2_X1 U699 ( .A1(n916), .A2(n637), .ZN(n626) );
  NOR2_X1 U700 ( .A1(n627), .A2(n626), .ZN(n631) );
  INV_X1 U701 ( .A(G299), .ZN(n630) );
  NAND2_X1 U702 ( .A1(n631), .A2(n630), .ZN(n628) );
  NAND2_X1 U703 ( .A1(n629), .A2(n628), .ZN(n635) );
  NOR2_X1 U704 ( .A1(n631), .A2(n630), .ZN(n633) );
  XNOR2_X1 U705 ( .A(n633), .B(n632), .ZN(n634) );
  NAND2_X1 U706 ( .A1(n635), .A2(n634), .ZN(n636) );
  XNOR2_X1 U707 ( .A(n636), .B(KEYINPUT29), .ZN(n641) );
  XOR2_X1 U708 ( .A(KEYINPUT25), .B(G2078), .Z(n948) );
  NOR2_X1 U709 ( .A1(n948), .A2(n654), .ZN(n639) );
  XOR2_X1 U710 ( .A(G1961), .B(KEYINPUT89), .Z(n926) );
  NOR2_X1 U711 ( .A1(n637), .A2(n926), .ZN(n638) );
  NOR2_X1 U712 ( .A1(n639), .A2(n638), .ZN(n650) );
  NOR2_X1 U713 ( .A1(G301), .A2(n650), .ZN(n640) );
  INV_X1 U714 ( .A(KEYINPUT92), .ZN(n642) );
  XNOR2_X1 U715 ( .A(n643), .B(n642), .ZN(n669) );
  NOR2_X1 U716 ( .A1(G2084), .A2(n654), .ZN(n670) );
  NAND2_X1 U717 ( .A1(G8), .A2(n644), .ZN(n690) );
  NOR2_X1 U718 ( .A1(G1966), .A2(n690), .ZN(n646) );
  INV_X1 U719 ( .A(KEYINPUT88), .ZN(n645) );
  XNOR2_X1 U720 ( .A(n646), .B(n645), .ZN(n672) );
  NAND2_X1 U721 ( .A1(n672), .A2(G8), .ZN(n647) );
  NOR2_X1 U722 ( .A1(n670), .A2(n647), .ZN(n648) );
  XOR2_X1 U723 ( .A(n648), .B(KEYINPUT30), .Z(n649) );
  NOR2_X1 U724 ( .A1(G168), .A2(n649), .ZN(n652) );
  AND2_X1 U725 ( .A1(G301), .A2(n650), .ZN(n651) );
  XOR2_X1 U726 ( .A(KEYINPUT31), .B(n653), .Z(n668) );
  INV_X1 U727 ( .A(G8), .ZN(n659) );
  NOR2_X1 U728 ( .A1(G1971), .A2(n690), .ZN(n656) );
  NOR2_X1 U729 ( .A1(G2090), .A2(n654), .ZN(n655) );
  NOR2_X1 U730 ( .A1(n656), .A2(n655), .ZN(n657) );
  NAND2_X1 U731 ( .A1(n657), .A2(G303), .ZN(n658) );
  OR2_X1 U732 ( .A1(n659), .A2(n658), .ZN(n661) );
  AND2_X1 U733 ( .A1(n668), .A2(n661), .ZN(n660) );
  NAND2_X1 U734 ( .A1(n669), .A2(n660), .ZN(n665) );
  INV_X1 U735 ( .A(n661), .ZN(n663) );
  AND2_X1 U736 ( .A1(G286), .A2(G8), .ZN(n662) );
  OR2_X1 U737 ( .A1(n663), .A2(n662), .ZN(n664) );
  NAND2_X1 U738 ( .A1(n665), .A2(n664), .ZN(n667) );
  XNOR2_X1 U739 ( .A(n667), .B(n666), .ZN(n676) );
  AND2_X1 U740 ( .A1(n669), .A2(n668), .ZN(n674) );
  NAND2_X1 U741 ( .A1(G8), .A2(n670), .ZN(n671) );
  NAND2_X1 U742 ( .A1(n672), .A2(n671), .ZN(n673) );
  NOR2_X1 U743 ( .A1(n674), .A2(n673), .ZN(n675) );
  INV_X1 U744 ( .A(n698), .ZN(n683) );
  NOR2_X1 U745 ( .A1(G1971), .A2(G303), .ZN(n677) );
  XNOR2_X1 U746 ( .A(n677), .B(KEYINPUT93), .ZN(n679) );
  INV_X1 U747 ( .A(KEYINPUT33), .ZN(n678) );
  AND2_X1 U748 ( .A1(n679), .A2(n678), .ZN(n681) );
  NOR2_X1 U749 ( .A1(G1976), .A2(G288), .ZN(n979) );
  NAND2_X1 U750 ( .A1(n683), .A2(n682), .ZN(n686) );
  NAND2_X1 U751 ( .A1(G1976), .A2(G288), .ZN(n980) );
  INV_X1 U752 ( .A(n980), .ZN(n684) );
  OR2_X1 U753 ( .A1(KEYINPUT33), .A2(n515), .ZN(n685) );
  NAND2_X1 U754 ( .A1(n686), .A2(n685), .ZN(n687) );
  XNOR2_X1 U755 ( .A(n687), .B(KEYINPUT94), .ZN(n688) );
  NOR2_X1 U756 ( .A1(n975), .A2(n688), .ZN(n693) );
  NAND2_X1 U757 ( .A1(n979), .A2(KEYINPUT33), .ZN(n689) );
  XNOR2_X1 U758 ( .A(KEYINPUT95), .B(n689), .ZN(n691) );
  INV_X1 U759 ( .A(n690), .ZN(n699) );
  NAND2_X1 U760 ( .A1(n691), .A2(n699), .ZN(n692) );
  AND2_X1 U761 ( .A1(n693), .A2(n692), .ZN(n704) );
  NOR2_X1 U762 ( .A1(G1981), .A2(G305), .ZN(n694) );
  XNOR2_X1 U763 ( .A(n694), .B(KEYINPUT24), .ZN(n695) );
  NAND2_X1 U764 ( .A1(n695), .A2(n699), .ZN(n702) );
  NAND2_X1 U765 ( .A1(G166), .A2(G8), .ZN(n696) );
  NOR2_X1 U766 ( .A1(G2090), .A2(n696), .ZN(n697) );
  NOR2_X1 U767 ( .A1(n698), .A2(n697), .ZN(n700) );
  OR2_X1 U768 ( .A1(n700), .A2(n699), .ZN(n701) );
  NAND2_X1 U769 ( .A1(n702), .A2(n701), .ZN(n703) );
  NOR2_X1 U770 ( .A1(n704), .A2(n703), .ZN(n738) );
  NOR2_X1 U771 ( .A1(n706), .A2(n705), .ZN(n751) );
  NAND2_X1 U772 ( .A1(G116), .A2(n883), .ZN(n708) );
  NAND2_X1 U773 ( .A1(G128), .A2(n885), .ZN(n707) );
  NAND2_X1 U774 ( .A1(n708), .A2(n707), .ZN(n709) );
  XNOR2_X1 U775 ( .A(n709), .B(KEYINPUT35), .ZN(n714) );
  NAND2_X1 U776 ( .A1(G104), .A2(n879), .ZN(n711) );
  NAND2_X1 U777 ( .A1(G140), .A2(n514), .ZN(n710) );
  NAND2_X1 U778 ( .A1(n711), .A2(n710), .ZN(n712) );
  XOR2_X1 U779 ( .A(KEYINPUT34), .B(n712), .Z(n713) );
  NAND2_X1 U780 ( .A1(n714), .A2(n713), .ZN(n715) );
  XOR2_X1 U781 ( .A(n715), .B(KEYINPUT36), .Z(n898) );
  XNOR2_X1 U782 ( .A(G2067), .B(KEYINPUT37), .ZN(n748) );
  NOR2_X1 U783 ( .A1(n898), .A2(n748), .ZN(n1006) );
  NAND2_X1 U784 ( .A1(n751), .A2(n1006), .ZN(n746) );
  NAND2_X1 U785 ( .A1(G117), .A2(n883), .ZN(n717) );
  NAND2_X1 U786 ( .A1(G141), .A2(n514), .ZN(n716) );
  NAND2_X1 U787 ( .A1(n717), .A2(n716), .ZN(n720) );
  NAND2_X1 U788 ( .A1(n879), .A2(G105), .ZN(n718) );
  XOR2_X1 U789 ( .A(KEYINPUT38), .B(n718), .Z(n719) );
  NOR2_X1 U790 ( .A1(n720), .A2(n719), .ZN(n722) );
  NAND2_X1 U791 ( .A1(n885), .A2(G129), .ZN(n721) );
  NAND2_X1 U792 ( .A1(n722), .A2(n721), .ZN(n897) );
  NAND2_X1 U793 ( .A1(n897), .A2(G1996), .ZN(n733) );
  XNOR2_X1 U794 ( .A(KEYINPUT84), .B(G1991), .ZN(n941) );
  NAND2_X1 U795 ( .A1(G119), .A2(n885), .ZN(n723) );
  XNOR2_X1 U796 ( .A(n723), .B(KEYINPUT82), .ZN(n730) );
  NAND2_X1 U797 ( .A1(G95), .A2(n879), .ZN(n725) );
  NAND2_X1 U798 ( .A1(G131), .A2(n514), .ZN(n724) );
  NAND2_X1 U799 ( .A1(n725), .A2(n724), .ZN(n728) );
  NAND2_X1 U800 ( .A1(G107), .A2(n883), .ZN(n726) );
  XNOR2_X1 U801 ( .A(KEYINPUT83), .B(n726), .ZN(n727) );
  NOR2_X1 U802 ( .A1(n728), .A2(n727), .ZN(n729) );
  NAND2_X1 U803 ( .A1(n730), .A2(n729), .ZN(n877) );
  NAND2_X1 U804 ( .A1(n941), .A2(n877), .ZN(n731) );
  XOR2_X1 U805 ( .A(KEYINPUT85), .B(n731), .Z(n732) );
  NAND2_X1 U806 ( .A1(n733), .A2(n732), .ZN(n734) );
  XNOR2_X1 U807 ( .A(n734), .B(KEYINPUT86), .ZN(n1010) );
  NAND2_X1 U808 ( .A1(n1010), .A2(n751), .ZN(n735) );
  XNOR2_X1 U809 ( .A(n735), .B(KEYINPUT87), .ZN(n743) );
  INV_X1 U810 ( .A(n743), .ZN(n736) );
  NAND2_X1 U811 ( .A1(n746), .A2(n736), .ZN(n737) );
  NOR2_X1 U812 ( .A1(n738), .A2(n737), .ZN(n740) );
  XNOR2_X1 U813 ( .A(G1986), .B(G290), .ZN(n971) );
  NAND2_X1 U814 ( .A1(n971), .A2(n751), .ZN(n739) );
  NAND2_X1 U815 ( .A1(n740), .A2(n739), .ZN(n754) );
  NOR2_X1 U816 ( .A1(G1996), .A2(n897), .ZN(n1014) );
  NOR2_X1 U817 ( .A1(G1986), .A2(G290), .ZN(n741) );
  NOR2_X1 U818 ( .A1(n941), .A2(n877), .ZN(n1003) );
  NOR2_X1 U819 ( .A1(n741), .A2(n1003), .ZN(n742) );
  NOR2_X1 U820 ( .A1(n743), .A2(n742), .ZN(n744) );
  NOR2_X1 U821 ( .A1(n1014), .A2(n744), .ZN(n745) );
  XNOR2_X1 U822 ( .A(KEYINPUT39), .B(n745), .ZN(n747) );
  NAND2_X1 U823 ( .A1(n747), .A2(n746), .ZN(n750) );
  AND2_X1 U824 ( .A1(n898), .A2(n748), .ZN(n749) );
  XOR2_X1 U825 ( .A(KEYINPUT96), .B(n749), .Z(n1012) );
  NAND2_X1 U826 ( .A1(n750), .A2(n1012), .ZN(n752) );
  NAND2_X1 U827 ( .A1(n752), .A2(n751), .ZN(n753) );
  NAND2_X1 U828 ( .A1(n754), .A2(n753), .ZN(n755) );
  XNOR2_X1 U829 ( .A(n755), .B(KEYINPUT40), .ZN(G329) );
  XOR2_X1 U830 ( .A(G2443), .B(G2446), .Z(n757) );
  XNOR2_X1 U831 ( .A(G2427), .B(G2451), .ZN(n756) );
  XNOR2_X1 U832 ( .A(n757), .B(n756), .ZN(n763) );
  XOR2_X1 U833 ( .A(G2430), .B(G2454), .Z(n759) );
  XNOR2_X1 U834 ( .A(G1348), .B(G1341), .ZN(n758) );
  XNOR2_X1 U835 ( .A(n759), .B(n758), .ZN(n761) );
  XOR2_X1 U836 ( .A(G2435), .B(G2438), .Z(n760) );
  XNOR2_X1 U837 ( .A(n761), .B(n760), .ZN(n762) );
  XOR2_X1 U838 ( .A(n763), .B(n762), .Z(n764) );
  AND2_X1 U839 ( .A1(G14), .A2(n764), .ZN(G401) );
  AND2_X1 U840 ( .A1(G452), .A2(G94), .ZN(G173) );
  NAND2_X1 U841 ( .A1(G111), .A2(n883), .ZN(n766) );
  NAND2_X1 U842 ( .A1(G135), .A2(n514), .ZN(n765) );
  NAND2_X1 U843 ( .A1(n766), .A2(n765), .ZN(n769) );
  NAND2_X1 U844 ( .A1(n885), .A2(G123), .ZN(n767) );
  XOR2_X1 U845 ( .A(KEYINPUT18), .B(n767), .Z(n768) );
  NOR2_X1 U846 ( .A1(n769), .A2(n768), .ZN(n771) );
  NAND2_X1 U847 ( .A1(n879), .A2(G99), .ZN(n770) );
  NAND2_X1 U848 ( .A1(n771), .A2(n770), .ZN(n1004) );
  XNOR2_X1 U849 ( .A(G2096), .B(n1004), .ZN(n772) );
  OR2_X1 U850 ( .A1(G2100), .A2(n772), .ZN(G156) );
  INV_X1 U851 ( .A(G57), .ZN(G237) );
  INV_X1 U852 ( .A(G132), .ZN(G219) );
  INV_X1 U853 ( .A(G82), .ZN(G220) );
  NAND2_X1 U854 ( .A1(G7), .A2(G661), .ZN(n773) );
  XNOR2_X1 U855 ( .A(n773), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U856 ( .A(G223), .ZN(n827) );
  NAND2_X1 U857 ( .A1(n827), .A2(G567), .ZN(n774) );
  XOR2_X1 U858 ( .A(KEYINPUT11), .B(n774), .Z(G234) );
  INV_X1 U859 ( .A(G860), .ZN(n779) );
  OR2_X1 U860 ( .A1(n967), .A2(n779), .ZN(G153) );
  NAND2_X1 U861 ( .A1(G868), .A2(G301), .ZN(n776) );
  OR2_X1 U862 ( .A1(n966), .A2(G868), .ZN(n775) );
  NAND2_X1 U863 ( .A1(n776), .A2(n775), .ZN(G284) );
  INV_X1 U864 ( .A(G868), .ZN(n809) );
  NOR2_X1 U865 ( .A1(G286), .A2(n809), .ZN(n778) );
  NOR2_X1 U866 ( .A1(G299), .A2(G868), .ZN(n777) );
  NOR2_X1 U867 ( .A1(n778), .A2(n777), .ZN(G297) );
  NAND2_X1 U868 ( .A1(n779), .A2(G559), .ZN(n780) );
  NAND2_X1 U869 ( .A1(n780), .A2(n966), .ZN(n781) );
  XNOR2_X1 U870 ( .A(n781), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U871 ( .A1(G559), .A2(n809), .ZN(n782) );
  NAND2_X1 U872 ( .A1(n966), .A2(n782), .ZN(n783) );
  XNOR2_X1 U873 ( .A(n783), .B(KEYINPUT73), .ZN(n785) );
  NOR2_X1 U874 ( .A1(n967), .A2(G868), .ZN(n784) );
  NOR2_X1 U875 ( .A1(n785), .A2(n784), .ZN(G282) );
  NAND2_X1 U876 ( .A1(G93), .A2(n786), .ZN(n789) );
  NAND2_X1 U877 ( .A1(G80), .A2(n787), .ZN(n788) );
  NAND2_X1 U878 ( .A1(n789), .A2(n788), .ZN(n790) );
  XNOR2_X1 U879 ( .A(KEYINPUT76), .B(n790), .ZN(n796) );
  NAND2_X1 U880 ( .A1(n791), .A2(G55), .ZN(n794) );
  NAND2_X1 U881 ( .A1(G67), .A2(n792), .ZN(n793) );
  NAND2_X1 U882 ( .A1(n794), .A2(n793), .ZN(n795) );
  OR2_X1 U883 ( .A1(n796), .A2(n795), .ZN(n808) );
  XNOR2_X1 U884 ( .A(n967), .B(KEYINPUT74), .ZN(n798) );
  NAND2_X1 U885 ( .A1(n966), .A2(G559), .ZN(n797) );
  XNOR2_X1 U886 ( .A(n798), .B(n797), .ZN(n806) );
  NOR2_X1 U887 ( .A1(n806), .A2(G860), .ZN(n799) );
  XOR2_X1 U888 ( .A(KEYINPUT75), .B(n799), .Z(n800) );
  XOR2_X1 U889 ( .A(n808), .B(n800), .Z(G145) );
  XNOR2_X1 U890 ( .A(KEYINPUT19), .B(G305), .ZN(n801) );
  XNOR2_X1 U891 ( .A(n801), .B(G288), .ZN(n802) );
  XNOR2_X1 U892 ( .A(n802), .B(n808), .ZN(n804) );
  XNOR2_X1 U893 ( .A(G299), .B(G166), .ZN(n803) );
  XNOR2_X1 U894 ( .A(n804), .B(n803), .ZN(n805) );
  XNOR2_X1 U895 ( .A(n805), .B(G290), .ZN(n901) );
  XNOR2_X1 U896 ( .A(n806), .B(n901), .ZN(n807) );
  NAND2_X1 U897 ( .A1(n807), .A2(G868), .ZN(n811) );
  NAND2_X1 U898 ( .A1(n809), .A2(n808), .ZN(n810) );
  NAND2_X1 U899 ( .A1(n811), .A2(n810), .ZN(G295) );
  NAND2_X1 U900 ( .A1(G2084), .A2(G2078), .ZN(n812) );
  XOR2_X1 U901 ( .A(KEYINPUT20), .B(n812), .Z(n813) );
  NAND2_X1 U902 ( .A1(G2090), .A2(n813), .ZN(n814) );
  XNOR2_X1 U903 ( .A(KEYINPUT21), .B(n814), .ZN(n815) );
  NAND2_X1 U904 ( .A1(n815), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U905 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NAND2_X1 U906 ( .A1(G483), .A2(G661), .ZN(n825) );
  NOR2_X1 U907 ( .A1(G220), .A2(G219), .ZN(n816) );
  XOR2_X1 U908 ( .A(KEYINPUT22), .B(n816), .Z(n817) );
  NOR2_X1 U909 ( .A1(G218), .A2(n817), .ZN(n818) );
  NAND2_X1 U910 ( .A1(G96), .A2(n818), .ZN(n834) );
  NAND2_X1 U911 ( .A1(n834), .A2(G2106), .ZN(n824) );
  NAND2_X1 U912 ( .A1(G120), .A2(G69), .ZN(n819) );
  NOR2_X1 U913 ( .A1(G237), .A2(n819), .ZN(n820) );
  XNOR2_X1 U914 ( .A(KEYINPUT78), .B(n820), .ZN(n821) );
  NAND2_X1 U915 ( .A1(n821), .A2(G108), .ZN(n822) );
  XOR2_X1 U916 ( .A(KEYINPUT79), .B(n822), .Z(n833) );
  NAND2_X1 U917 ( .A1(n833), .A2(G567), .ZN(n823) );
  NAND2_X1 U918 ( .A1(n824), .A2(n823), .ZN(n856) );
  NOR2_X1 U919 ( .A1(n825), .A2(n856), .ZN(n826) );
  XNOR2_X1 U920 ( .A(n826), .B(KEYINPUT80), .ZN(n832) );
  NAND2_X1 U921 ( .A1(G36), .A2(n832), .ZN(G176) );
  NAND2_X1 U922 ( .A1(G2106), .A2(n827), .ZN(G217) );
  NAND2_X1 U923 ( .A1(G15), .A2(G2), .ZN(n829) );
  INV_X1 U924 ( .A(G661), .ZN(n828) );
  NOR2_X1 U925 ( .A1(n829), .A2(n828), .ZN(n830) );
  XNOR2_X1 U926 ( .A(n830), .B(KEYINPUT97), .ZN(G259) );
  NAND2_X1 U927 ( .A1(G3), .A2(G1), .ZN(n831) );
  NAND2_X1 U928 ( .A1(n832), .A2(n831), .ZN(G188) );
  XOR2_X1 U929 ( .A(G96), .B(KEYINPUT98), .Z(G221) );
  XNOR2_X1 U930 ( .A(G108), .B(KEYINPUT113), .ZN(G238) );
  INV_X1 U932 ( .A(G120), .ZN(G236) );
  INV_X1 U933 ( .A(G69), .ZN(G235) );
  NOR2_X1 U934 ( .A1(n834), .A2(n833), .ZN(n835) );
  XNOR2_X1 U935 ( .A(n835), .B(KEYINPUT99), .ZN(G261) );
  INV_X1 U936 ( .A(G261), .ZN(G325) );
  XOR2_X1 U937 ( .A(KEYINPUT41), .B(G1961), .Z(n837) );
  XNOR2_X1 U938 ( .A(G1996), .B(G1991), .ZN(n836) );
  XNOR2_X1 U939 ( .A(n837), .B(n836), .ZN(n838) );
  XOR2_X1 U940 ( .A(n838), .B(KEYINPUT102), .Z(n840) );
  XNOR2_X1 U941 ( .A(G1956), .B(G1971), .ZN(n839) );
  XNOR2_X1 U942 ( .A(n840), .B(n839), .ZN(n844) );
  XOR2_X1 U943 ( .A(G1976), .B(G1981), .Z(n842) );
  XNOR2_X1 U944 ( .A(G1986), .B(G1966), .ZN(n841) );
  XNOR2_X1 U945 ( .A(n842), .B(n841), .ZN(n843) );
  XOR2_X1 U946 ( .A(n844), .B(n843), .Z(n846) );
  XNOR2_X1 U947 ( .A(G2474), .B(KEYINPUT101), .ZN(n845) );
  XNOR2_X1 U948 ( .A(n846), .B(n845), .ZN(G229) );
  XOR2_X1 U949 ( .A(G2096), .B(KEYINPUT43), .Z(n848) );
  XNOR2_X1 U950 ( .A(G2090), .B(KEYINPUT42), .ZN(n847) );
  XNOR2_X1 U951 ( .A(n848), .B(n847), .ZN(n849) );
  XOR2_X1 U952 ( .A(n849), .B(G2678), .Z(n851) );
  XNOR2_X1 U953 ( .A(G2067), .B(G2072), .ZN(n850) );
  XNOR2_X1 U954 ( .A(n851), .B(n850), .ZN(n855) );
  XOR2_X1 U955 ( .A(KEYINPUT100), .B(G2100), .Z(n853) );
  XNOR2_X1 U956 ( .A(G2084), .B(G2078), .ZN(n852) );
  XNOR2_X1 U957 ( .A(n853), .B(n852), .ZN(n854) );
  XNOR2_X1 U958 ( .A(n855), .B(n854), .ZN(G227) );
  INV_X1 U959 ( .A(n856), .ZN(G319) );
  NAND2_X1 U960 ( .A1(G112), .A2(n883), .ZN(n858) );
  NAND2_X1 U961 ( .A1(G100), .A2(n879), .ZN(n857) );
  NAND2_X1 U962 ( .A1(n858), .A2(n857), .ZN(n865) );
  NAND2_X1 U963 ( .A1(G136), .A2(n514), .ZN(n859) );
  XNOR2_X1 U964 ( .A(n859), .B(KEYINPUT104), .ZN(n863) );
  XOR2_X1 U965 ( .A(KEYINPUT44), .B(KEYINPUT103), .Z(n861) );
  NAND2_X1 U966 ( .A1(G124), .A2(n885), .ZN(n860) );
  XNOR2_X1 U967 ( .A(n861), .B(n860), .ZN(n862) );
  NAND2_X1 U968 ( .A1(n863), .A2(n862), .ZN(n864) );
  NOR2_X1 U969 ( .A1(n865), .A2(n864), .ZN(G162) );
  XOR2_X1 U970 ( .A(KEYINPUT46), .B(KEYINPUT48), .Z(n876) );
  NAND2_X1 U971 ( .A1(G118), .A2(n883), .ZN(n867) );
  NAND2_X1 U972 ( .A1(G130), .A2(n885), .ZN(n866) );
  NAND2_X1 U973 ( .A1(n867), .A2(n866), .ZN(n873) );
  NAND2_X1 U974 ( .A1(G106), .A2(n879), .ZN(n869) );
  NAND2_X1 U975 ( .A1(G142), .A2(n514), .ZN(n868) );
  NAND2_X1 U976 ( .A1(n869), .A2(n868), .ZN(n870) );
  XNOR2_X1 U977 ( .A(KEYINPUT105), .B(n870), .ZN(n871) );
  XNOR2_X1 U978 ( .A(KEYINPUT45), .B(n871), .ZN(n872) );
  NOR2_X1 U979 ( .A1(n873), .A2(n872), .ZN(n874) );
  XNOR2_X1 U980 ( .A(KEYINPUT107), .B(n874), .ZN(n875) );
  XNOR2_X1 U981 ( .A(n876), .B(n875), .ZN(n895) );
  XNOR2_X1 U982 ( .A(G164), .B(n877), .ZN(n878) );
  XNOR2_X1 U983 ( .A(n878), .B(n1004), .ZN(n891) );
  NAND2_X1 U984 ( .A1(G103), .A2(n879), .ZN(n882) );
  NAND2_X1 U985 ( .A1(G139), .A2(n514), .ZN(n881) );
  NAND2_X1 U986 ( .A1(n882), .A2(n881), .ZN(n890) );
  NAND2_X1 U987 ( .A1(n883), .A2(G115), .ZN(n884) );
  XNOR2_X1 U988 ( .A(n884), .B(KEYINPUT106), .ZN(n887) );
  NAND2_X1 U989 ( .A1(G127), .A2(n885), .ZN(n886) );
  NAND2_X1 U990 ( .A1(n887), .A2(n886), .ZN(n888) );
  XOR2_X1 U991 ( .A(KEYINPUT47), .B(n888), .Z(n889) );
  NOR2_X1 U992 ( .A1(n890), .A2(n889), .ZN(n997) );
  XOR2_X1 U993 ( .A(n891), .B(n997), .Z(n893) );
  XNOR2_X1 U994 ( .A(G160), .B(G162), .ZN(n892) );
  XNOR2_X1 U995 ( .A(n893), .B(n892), .ZN(n894) );
  XOR2_X1 U996 ( .A(n895), .B(n894), .Z(n896) );
  XNOR2_X1 U997 ( .A(n897), .B(n896), .ZN(n899) );
  XOR2_X1 U998 ( .A(n899), .B(n898), .Z(n900) );
  NOR2_X1 U999 ( .A1(G37), .A2(n900), .ZN(G395) );
  XOR2_X1 U1000 ( .A(KEYINPUT108), .B(KEYINPUT109), .Z(n903) );
  XNOR2_X1 U1001 ( .A(n966), .B(n901), .ZN(n902) );
  XNOR2_X1 U1002 ( .A(n903), .B(n902), .ZN(n904) );
  XNOR2_X1 U1003 ( .A(n904), .B(G301), .ZN(n905) );
  XNOR2_X1 U1004 ( .A(n905), .B(n967), .ZN(n906) );
  XNOR2_X1 U1005 ( .A(n906), .B(G286), .ZN(n907) );
  NOR2_X1 U1006 ( .A1(G37), .A2(n907), .ZN(G397) );
  NOR2_X1 U1007 ( .A1(G229), .A2(G227), .ZN(n908) );
  XOR2_X1 U1008 ( .A(KEYINPUT49), .B(n908), .Z(n909) );
  XNOR2_X1 U1009 ( .A(KEYINPUT110), .B(n909), .ZN(n910) );
  NAND2_X1 U1010 ( .A1(n910), .A2(G319), .ZN(n911) );
  NOR2_X1 U1011 ( .A1(G401), .A2(n911), .ZN(n912) );
  XOR2_X1 U1012 ( .A(KEYINPUT111), .B(n912), .Z(n915) );
  NOR2_X1 U1013 ( .A1(G395), .A2(G397), .ZN(n913) );
  XNOR2_X1 U1014 ( .A(KEYINPUT112), .B(n913), .ZN(n914) );
  NAND2_X1 U1015 ( .A1(n915), .A2(n914), .ZN(G225) );
  INV_X1 U1016 ( .A(G225), .ZN(G308) );
  XNOR2_X1 U1017 ( .A(G20), .B(n916), .ZN(n920) );
  XNOR2_X1 U1018 ( .A(G1341), .B(G19), .ZN(n918) );
  XNOR2_X1 U1019 ( .A(G6), .B(G1981), .ZN(n917) );
  NOR2_X1 U1020 ( .A1(n918), .A2(n917), .ZN(n919) );
  NAND2_X1 U1021 ( .A1(n920), .A2(n919), .ZN(n923) );
  XOR2_X1 U1022 ( .A(KEYINPUT59), .B(G1348), .Z(n921) );
  XNOR2_X1 U1023 ( .A(G4), .B(n921), .ZN(n922) );
  NOR2_X1 U1024 ( .A1(n923), .A2(n922), .ZN(n924) );
  XNOR2_X1 U1025 ( .A(KEYINPUT124), .B(n924), .ZN(n925) );
  XNOR2_X1 U1026 ( .A(n925), .B(KEYINPUT60), .ZN(n930) );
  XNOR2_X1 U1027 ( .A(G1966), .B(G21), .ZN(n928) );
  XNOR2_X1 U1028 ( .A(n926), .B(G5), .ZN(n927) );
  NOR2_X1 U1029 ( .A1(n928), .A2(n927), .ZN(n929) );
  NAND2_X1 U1030 ( .A1(n930), .A2(n929), .ZN(n937) );
  XNOR2_X1 U1031 ( .A(G1971), .B(G22), .ZN(n932) );
  XNOR2_X1 U1032 ( .A(G23), .B(G1976), .ZN(n931) );
  NOR2_X1 U1033 ( .A1(n932), .A2(n931), .ZN(n934) );
  XOR2_X1 U1034 ( .A(G1986), .B(G24), .Z(n933) );
  NAND2_X1 U1035 ( .A1(n934), .A2(n933), .ZN(n935) );
  XNOR2_X1 U1036 ( .A(KEYINPUT58), .B(n935), .ZN(n936) );
  NOR2_X1 U1037 ( .A1(n937), .A2(n936), .ZN(n938) );
  XOR2_X1 U1038 ( .A(KEYINPUT61), .B(n938), .Z(n939) );
  NOR2_X1 U1039 ( .A1(G16), .A2(n939), .ZN(n940) );
  XOR2_X1 U1040 ( .A(KEYINPUT125), .B(n940), .Z(n995) );
  XNOR2_X1 U1041 ( .A(n941), .B(G25), .ZN(n953) );
  XNOR2_X1 U1042 ( .A(n942), .B(G32), .ZN(n944) );
  XNOR2_X1 U1043 ( .A(G26), .B(G2067), .ZN(n943) );
  NOR2_X1 U1044 ( .A1(n944), .A2(n943), .ZN(n947) );
  XOR2_X1 U1045 ( .A(G2072), .B(KEYINPUT118), .Z(n945) );
  XNOR2_X1 U1046 ( .A(G33), .B(n945), .ZN(n946) );
  NAND2_X1 U1047 ( .A1(n947), .A2(n946), .ZN(n950) );
  XNOR2_X1 U1048 ( .A(G27), .B(n948), .ZN(n949) );
  NOR2_X1 U1049 ( .A1(n950), .A2(n949), .ZN(n951) );
  XNOR2_X1 U1050 ( .A(KEYINPUT119), .B(n951), .ZN(n952) );
  NOR2_X1 U1051 ( .A1(n953), .A2(n952), .ZN(n954) );
  NAND2_X1 U1052 ( .A1(G28), .A2(n954), .ZN(n955) );
  XNOR2_X1 U1053 ( .A(n955), .B(KEYINPUT53), .ZN(n958) );
  XOR2_X1 U1054 ( .A(G2084), .B(G34), .Z(n956) );
  XNOR2_X1 U1055 ( .A(KEYINPUT54), .B(n956), .ZN(n957) );
  NAND2_X1 U1056 ( .A1(n958), .A2(n957), .ZN(n960) );
  XNOR2_X1 U1057 ( .A(G35), .B(G2090), .ZN(n959) );
  NOR2_X1 U1058 ( .A1(n960), .A2(n959), .ZN(n961) );
  XNOR2_X1 U1059 ( .A(KEYINPUT55), .B(n961), .ZN(n963) );
  INV_X1 U1060 ( .A(G29), .ZN(n962) );
  NAND2_X1 U1061 ( .A1(n963), .A2(n962), .ZN(n964) );
  NAND2_X1 U1062 ( .A1(n964), .A2(G11), .ZN(n965) );
  XOR2_X1 U1063 ( .A(KEYINPUT120), .B(n965), .Z(n993) );
  XNOR2_X1 U1064 ( .A(G16), .B(KEYINPUT56), .ZN(n991) );
  XOR2_X1 U1065 ( .A(G1348), .B(n966), .Z(n969) );
  XNOR2_X1 U1066 ( .A(n967), .B(G1341), .ZN(n968) );
  NOR2_X1 U1067 ( .A1(n969), .A2(n968), .ZN(n973) );
  XNOR2_X1 U1068 ( .A(G1961), .B(G301), .ZN(n970) );
  NOR2_X1 U1069 ( .A1(n971), .A2(n970), .ZN(n972) );
  NAND2_X1 U1070 ( .A1(n973), .A2(n972), .ZN(n988) );
  XOR2_X1 U1071 ( .A(G168), .B(G1966), .Z(n974) );
  NOR2_X1 U1072 ( .A1(n975), .A2(n974), .ZN(n976) );
  XOR2_X1 U1073 ( .A(KEYINPUT57), .B(n976), .Z(n986) );
  XNOR2_X1 U1074 ( .A(G166), .B(G1971), .ZN(n977) );
  XNOR2_X1 U1075 ( .A(n977), .B(KEYINPUT121), .ZN(n983) );
  XNOR2_X1 U1076 ( .A(G299), .B(G1956), .ZN(n978) );
  NOR2_X1 U1077 ( .A1(n979), .A2(n978), .ZN(n981) );
  NAND2_X1 U1078 ( .A1(n981), .A2(n980), .ZN(n982) );
  NOR2_X1 U1079 ( .A1(n983), .A2(n982), .ZN(n984) );
  XNOR2_X1 U1080 ( .A(n984), .B(KEYINPUT122), .ZN(n985) );
  NAND2_X1 U1081 ( .A1(n986), .A2(n985), .ZN(n987) );
  NOR2_X1 U1082 ( .A1(n988), .A2(n987), .ZN(n989) );
  XNOR2_X1 U1083 ( .A(KEYINPUT123), .B(n989), .ZN(n990) );
  NAND2_X1 U1084 ( .A1(n991), .A2(n990), .ZN(n992) );
  NAND2_X1 U1085 ( .A1(n993), .A2(n992), .ZN(n994) );
  NOR2_X1 U1086 ( .A1(n995), .A2(n994), .ZN(n996) );
  XNOR2_X1 U1087 ( .A(n996), .B(KEYINPUT126), .ZN(n1027) );
  XOR2_X1 U1088 ( .A(n997), .B(KEYINPUT117), .Z(n998) );
  XOR2_X1 U1089 ( .A(G2072), .B(n998), .Z(n1000) );
  XOR2_X1 U1090 ( .A(G164), .B(G2078), .Z(n999) );
  NOR2_X1 U1091 ( .A1(n1000), .A2(n999), .ZN(n1001) );
  XOR2_X1 U1092 ( .A(KEYINPUT50), .B(n1001), .Z(n1021) );
  XOR2_X1 U1093 ( .A(G160), .B(G2084), .Z(n1002) );
  NOR2_X1 U1094 ( .A1(n1003), .A2(n1002), .ZN(n1005) );
  NAND2_X1 U1095 ( .A1(n1005), .A2(n1004), .ZN(n1007) );
  NOR2_X1 U1096 ( .A1(n1007), .A2(n1006), .ZN(n1008) );
  XOR2_X1 U1097 ( .A(KEYINPUT114), .B(n1008), .Z(n1009) );
  NOR2_X1 U1098 ( .A1(n1010), .A2(n1009), .ZN(n1011) );
  NAND2_X1 U1099 ( .A1(n1012), .A2(n1011), .ZN(n1018) );
  XOR2_X1 U1100 ( .A(G2090), .B(G162), .Z(n1013) );
  NOR2_X1 U1101 ( .A1(n1014), .A2(n1013), .ZN(n1015) );
  XOR2_X1 U1102 ( .A(KEYINPUT51), .B(n1015), .Z(n1016) );
  XNOR2_X1 U1103 ( .A(n1016), .B(KEYINPUT115), .ZN(n1017) );
  NOR2_X1 U1104 ( .A1(n1018), .A2(n1017), .ZN(n1019) );
  XOR2_X1 U1105 ( .A(KEYINPUT116), .B(n1019), .Z(n1020) );
  NOR2_X1 U1106 ( .A1(n1021), .A2(n1020), .ZN(n1022) );
  XNOR2_X1 U1107 ( .A(KEYINPUT52), .B(n1022), .ZN(n1024) );
  INV_X1 U1108 ( .A(KEYINPUT55), .ZN(n1023) );
  NAND2_X1 U1109 ( .A1(n1024), .A2(n1023), .ZN(n1025) );
  NAND2_X1 U1110 ( .A1(n1025), .A2(G29), .ZN(n1026) );
  NAND2_X1 U1111 ( .A1(n1027), .A2(n1026), .ZN(n1028) );
  XOR2_X1 U1112 ( .A(KEYINPUT62), .B(n1028), .Z(G311) );
  INV_X1 U1113 ( .A(G311), .ZN(G150) );
  INV_X1 U1114 ( .A(G301), .ZN(G171) );
endmodule

