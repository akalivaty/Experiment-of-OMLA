//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 1 0 1 0 1 0 1 0 0 0 1 1 1 0 0 0 1 1 1 0 1 1 1 1 1 1 0 1 0 1 1 1 0 0 1 1 1 0 0 0 1 0 0 1 1 0 0 1 1 0 1 1 1 1 0 1 1 0 0 0 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:22:20 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n592, new_n593, new_n594,
    new_n595, new_n596, new_n597, new_n599, new_n600, new_n601, new_n602,
    new_n603, new_n604, new_n605, new_n607, new_n608, new_n609, new_n610,
    new_n611, new_n612, new_n613, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n632, new_n633,
    new_n634, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n649,
    new_n651, new_n652, new_n653, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n663, new_n664, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n694, new_n695, new_n696,
    new_n697, new_n698, new_n699, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n860, new_n861, new_n862, new_n863,
    new_n864, new_n865, new_n866, new_n868, new_n869, new_n870, new_n871,
    new_n872, new_n873, new_n874, new_n875, new_n876, new_n877, new_n878,
    new_n879, new_n880, new_n881, new_n882, new_n883, new_n884, new_n885,
    new_n886, new_n887, new_n888, new_n889, new_n890, new_n891, new_n892,
    new_n893, new_n894, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n935, new_n936, new_n937, new_n938,
    new_n939, new_n940, new_n941, new_n942;
  INV_X1    g000(.A(G953), .ZN(new_n187));
  NAND3_X1  g001(.A1(new_n187), .A2(G221), .A3(G234), .ZN(new_n188));
  XNOR2_X1  g002(.A(new_n188), .B(KEYINPUT77), .ZN(new_n189));
  XOR2_X1   g003(.A(KEYINPUT22), .B(G137), .Z(new_n190));
  XNOR2_X1  g004(.A(new_n189), .B(new_n190), .ZN(new_n191));
  INV_X1    g005(.A(G146), .ZN(new_n192));
  INV_X1    g006(.A(G140), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n193), .A2(G125), .ZN(new_n194));
  NOR2_X1   g008(.A1(new_n194), .A2(KEYINPUT16), .ZN(new_n195));
  INV_X1    g009(.A(G125), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n196), .A2(G140), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n194), .A2(new_n197), .ZN(new_n198));
  INV_X1    g012(.A(new_n198), .ZN(new_n199));
  AOI211_X1 g013(.A(new_n192), .B(new_n195), .C1(new_n199), .C2(KEYINPUT16), .ZN(new_n200));
  INV_X1    g014(.A(new_n200), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n199), .A2(new_n192), .ZN(new_n202));
  INV_X1    g016(.A(G128), .ZN(new_n203));
  NOR2_X1   g017(.A1(new_n203), .A2(G119), .ZN(new_n204));
  XNOR2_X1  g018(.A(KEYINPUT69), .B(G128), .ZN(new_n205));
  AOI21_X1  g019(.A(new_n204), .B1(new_n205), .B2(G119), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n206), .A2(KEYINPUT23), .ZN(new_n207));
  INV_X1    g021(.A(G119), .ZN(new_n208));
  OR3_X1    g022(.A1(new_n208), .A2(KEYINPUT23), .A3(G128), .ZN(new_n209));
  AOI21_X1  g023(.A(G110), .B1(new_n207), .B2(new_n209), .ZN(new_n210));
  XOR2_X1   g024(.A(KEYINPUT24), .B(G110), .Z(new_n211));
  NOR2_X1   g025(.A1(new_n206), .A2(new_n211), .ZN(new_n212));
  OAI211_X1 g026(.A(new_n201), .B(new_n202), .C1(new_n210), .C2(new_n212), .ZN(new_n213));
  NAND3_X1  g027(.A1(new_n207), .A2(G110), .A3(new_n209), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n206), .A2(new_n211), .ZN(new_n215));
  AOI21_X1  g029(.A(new_n195), .B1(new_n199), .B2(KEYINPUT16), .ZN(new_n216));
  NOR2_X1   g030(.A1(new_n216), .A2(G146), .ZN(new_n217));
  OAI211_X1 g031(.A(new_n214), .B(new_n215), .C1(new_n217), .C2(new_n200), .ZN(new_n218));
  AOI21_X1  g032(.A(new_n191), .B1(new_n213), .B2(new_n218), .ZN(new_n219));
  INV_X1    g033(.A(new_n219), .ZN(new_n220));
  NAND3_X1  g034(.A1(new_n213), .A2(new_n218), .A3(new_n191), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  XOR2_X1   g036(.A(KEYINPUT75), .B(G902), .Z(new_n223));
  INV_X1    g037(.A(new_n223), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n222), .A2(new_n224), .ZN(new_n225));
  INV_X1    g039(.A(KEYINPUT79), .ZN(new_n226));
  XOR2_X1   g040(.A(KEYINPUT78), .B(KEYINPUT25), .Z(new_n227));
  NAND3_X1  g041(.A1(new_n225), .A2(new_n226), .A3(new_n227), .ZN(new_n228));
  AOI21_X1  g042(.A(new_n223), .B1(new_n220), .B2(new_n221), .ZN(new_n229));
  INV_X1    g043(.A(new_n227), .ZN(new_n230));
  OAI21_X1  g044(.A(KEYINPUT79), .B1(new_n229), .B2(new_n230), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n229), .A2(KEYINPUT25), .ZN(new_n232));
  NAND3_X1  g046(.A1(new_n228), .A2(new_n231), .A3(new_n232), .ZN(new_n233));
  INV_X1    g047(.A(G234), .ZN(new_n234));
  OAI21_X1  g048(.A(G217), .B1(new_n223), .B2(new_n234), .ZN(new_n235));
  XOR2_X1   g049(.A(new_n235), .B(KEYINPUT76), .Z(new_n236));
  NAND2_X1  g050(.A1(new_n233), .A2(new_n236), .ZN(new_n237));
  NOR2_X1   g051(.A1(new_n236), .A2(G902), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n222), .A2(new_n238), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n237), .A2(new_n239), .ZN(new_n240));
  XNOR2_X1  g054(.A(new_n240), .B(KEYINPUT80), .ZN(new_n241));
  XOR2_X1   g055(.A(G116), .B(G119), .Z(new_n242));
  XNOR2_X1  g056(.A(KEYINPUT2), .B(G113), .ZN(new_n243));
  XNOR2_X1  g057(.A(new_n242), .B(new_n243), .ZN(new_n244));
  INV_X1    g058(.A(new_n244), .ZN(new_n245));
  XNOR2_X1  g059(.A(G134), .B(G137), .ZN(new_n246));
  INV_X1    g060(.A(G131), .ZN(new_n247));
  OAI21_X1  g061(.A(KEYINPUT68), .B1(new_n246), .B2(new_n247), .ZN(new_n248));
  INV_X1    g062(.A(KEYINPUT68), .ZN(new_n249));
  INV_X1    g063(.A(G137), .ZN(new_n250));
  NOR2_X1   g064(.A1(new_n250), .A2(G134), .ZN(new_n251));
  INV_X1    g065(.A(G134), .ZN(new_n252));
  NOR2_X1   g066(.A1(new_n252), .A2(G137), .ZN(new_n253));
  OAI211_X1 g067(.A(new_n249), .B(G131), .C1(new_n251), .C2(new_n253), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n248), .A2(new_n254), .ZN(new_n255));
  INV_X1    g069(.A(KEYINPUT66), .ZN(new_n256));
  INV_X1    g070(.A(KEYINPUT11), .ZN(new_n257));
  AOI22_X1  g071(.A1(new_n256), .A2(new_n257), .B1(new_n252), .B2(G137), .ZN(new_n258));
  OAI22_X1  g072(.A1(new_n256), .A2(new_n257), .B1(new_n252), .B2(G137), .ZN(new_n259));
  NAND4_X1  g073(.A1(new_n250), .A2(KEYINPUT66), .A3(KEYINPUT11), .A4(G134), .ZN(new_n260));
  NAND4_X1  g074(.A1(new_n258), .A2(new_n259), .A3(new_n247), .A4(new_n260), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n255), .A2(new_n261), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n192), .A2(G143), .ZN(new_n263));
  INV_X1    g077(.A(G143), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n264), .A2(G146), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n263), .A2(new_n265), .ZN(new_n266));
  INV_X1    g080(.A(KEYINPUT1), .ZN(new_n267));
  AOI21_X1  g081(.A(new_n267), .B1(G143), .B2(new_n192), .ZN(new_n268));
  OAI21_X1  g082(.A(new_n266), .B1(new_n205), .B2(new_n268), .ZN(new_n269));
  NAND3_X1  g083(.A1(new_n192), .A2(KEYINPUT64), .A3(G143), .ZN(new_n270));
  NOR2_X1   g084(.A1(new_n203), .A2(KEYINPUT1), .ZN(new_n271));
  INV_X1    g085(.A(KEYINPUT64), .ZN(new_n272));
  AOI21_X1  g086(.A(new_n272), .B1(new_n264), .B2(G146), .ZN(new_n273));
  NOR2_X1   g087(.A1(new_n264), .A2(G146), .ZN(new_n274));
  OAI211_X1 g088(.A(new_n270), .B(new_n271), .C1(new_n273), .C2(new_n274), .ZN(new_n275));
  AND2_X1   g089(.A1(new_n269), .A2(new_n275), .ZN(new_n276));
  OAI21_X1  g090(.A(KEYINPUT70), .B1(new_n262), .B2(new_n276), .ZN(new_n277));
  AND3_X1   g091(.A1(new_n258), .A2(new_n259), .A3(new_n260), .ZN(new_n278));
  AOI22_X1  g092(.A1(new_n278), .A2(new_n247), .B1(new_n248), .B2(new_n254), .ZN(new_n279));
  INV_X1    g093(.A(KEYINPUT70), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n269), .A2(new_n275), .ZN(new_n281));
  NAND3_X1  g095(.A1(new_n279), .A2(new_n280), .A3(new_n281), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n277), .A2(new_n282), .ZN(new_n283));
  INV_X1    g097(.A(KEYINPUT0), .ZN(new_n284));
  NOR2_X1   g098(.A1(new_n284), .A2(new_n203), .ZN(new_n285));
  INV_X1    g099(.A(new_n285), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n284), .A2(new_n203), .ZN(new_n287));
  NAND3_X1  g101(.A1(new_n286), .A2(new_n266), .A3(new_n287), .ZN(new_n288));
  OAI211_X1 g102(.A(new_n285), .B(new_n270), .C1(new_n273), .C2(new_n274), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  INV_X1    g104(.A(KEYINPUT65), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  NAND3_X1  g106(.A1(new_n258), .A2(new_n259), .A3(new_n260), .ZN(new_n293));
  INV_X1    g107(.A(KEYINPUT67), .ZN(new_n294));
  NAND3_X1  g108(.A1(new_n293), .A2(new_n294), .A3(G131), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n294), .A2(G131), .ZN(new_n296));
  NAND4_X1  g110(.A1(new_n258), .A2(new_n259), .A3(new_n296), .A4(new_n260), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n295), .A2(new_n297), .ZN(new_n298));
  NAND3_X1  g112(.A1(new_n288), .A2(new_n289), .A3(KEYINPUT65), .ZN(new_n299));
  NAND3_X1  g113(.A1(new_n292), .A2(new_n298), .A3(new_n299), .ZN(new_n300));
  AOI21_X1  g114(.A(new_n245), .B1(new_n283), .B2(new_n300), .ZN(new_n301));
  AND3_X1   g115(.A1(new_n269), .A2(new_n275), .A3(KEYINPUT71), .ZN(new_n302));
  AOI21_X1  g116(.A(KEYINPUT71), .B1(new_n269), .B2(new_n275), .ZN(new_n303));
  OAI21_X1  g117(.A(new_n279), .B1(new_n302), .B2(new_n303), .ZN(new_n304));
  INV_X1    g118(.A(new_n290), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n298), .A2(new_n305), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n304), .A2(new_n306), .ZN(new_n307));
  NOR2_X1   g121(.A1(new_n307), .A2(new_n244), .ZN(new_n308));
  OAI21_X1  g122(.A(KEYINPUT28), .B1(new_n301), .B2(new_n308), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n309), .A2(KEYINPUT74), .ZN(new_n310));
  NOR2_X1   g124(.A1(new_n308), .A2(KEYINPUT28), .ZN(new_n311));
  INV_X1    g125(.A(new_n311), .ZN(new_n312));
  INV_X1    g126(.A(KEYINPUT74), .ZN(new_n313));
  OAI211_X1 g127(.A(new_n313), .B(KEYINPUT28), .C1(new_n301), .C2(new_n308), .ZN(new_n314));
  NAND3_X1  g128(.A1(new_n310), .A2(new_n312), .A3(new_n314), .ZN(new_n315));
  XNOR2_X1  g129(.A(KEYINPUT73), .B(G237), .ZN(new_n316));
  NAND3_X1  g130(.A1(new_n316), .A2(G210), .A3(new_n187), .ZN(new_n317));
  INV_X1    g131(.A(G101), .ZN(new_n318));
  XNOR2_X1  g132(.A(new_n317), .B(new_n318), .ZN(new_n319));
  XNOR2_X1  g133(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n320));
  XOR2_X1   g134(.A(new_n319), .B(new_n320), .Z(new_n321));
  INV_X1    g135(.A(new_n321), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n315), .A2(new_n322), .ZN(new_n323));
  INV_X1    g137(.A(KEYINPUT30), .ZN(new_n324));
  NOR2_X1   g138(.A1(new_n307), .A2(new_n324), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n325), .A2(KEYINPUT72), .ZN(new_n326));
  INV_X1    g140(.A(KEYINPUT72), .ZN(new_n327));
  AOI21_X1  g141(.A(new_n280), .B1(new_n279), .B2(new_n281), .ZN(new_n328));
  AND4_X1   g142(.A1(new_n280), .A2(new_n281), .A3(new_n255), .A4(new_n261), .ZN(new_n329));
  OAI21_X1  g143(.A(new_n300), .B1(new_n328), .B2(new_n329), .ZN(new_n330));
  AOI21_X1  g144(.A(new_n327), .B1(new_n330), .B2(new_n324), .ZN(new_n331));
  OAI211_X1 g145(.A(new_n326), .B(new_n244), .C1(new_n331), .C2(new_n325), .ZN(new_n332));
  INV_X1    g146(.A(new_n308), .ZN(new_n333));
  NAND3_X1  g147(.A1(new_n332), .A2(new_n321), .A3(new_n333), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n334), .A2(KEYINPUT31), .ZN(new_n335));
  INV_X1    g149(.A(KEYINPUT31), .ZN(new_n336));
  NAND4_X1  g150(.A1(new_n332), .A2(new_n336), .A3(new_n321), .A4(new_n333), .ZN(new_n337));
  NAND3_X1  g151(.A1(new_n323), .A2(new_n335), .A3(new_n337), .ZN(new_n338));
  NOR2_X1   g152(.A1(G472), .A2(G902), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n338), .A2(new_n339), .ZN(new_n340));
  INV_X1    g154(.A(KEYINPUT32), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n340), .A2(new_n341), .ZN(new_n342));
  NAND3_X1  g156(.A1(new_n338), .A2(KEYINPUT32), .A3(new_n339), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n315), .A2(new_n321), .ZN(new_n344));
  NAND3_X1  g158(.A1(new_n332), .A2(new_n322), .A3(new_n333), .ZN(new_n345));
  AOI21_X1  g159(.A(KEYINPUT29), .B1(new_n344), .B2(new_n345), .ZN(new_n346));
  XNOR2_X1  g160(.A(new_n307), .B(new_n244), .ZN(new_n347));
  AOI21_X1  g161(.A(new_n311), .B1(new_n347), .B2(KEYINPUT28), .ZN(new_n348));
  NAND3_X1  g162(.A1(new_n348), .A2(KEYINPUT29), .A3(new_n321), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n349), .A2(new_n224), .ZN(new_n350));
  OAI21_X1  g164(.A(G472), .B1(new_n346), .B2(new_n350), .ZN(new_n351));
  NAND3_X1  g165(.A1(new_n342), .A2(new_n343), .A3(new_n351), .ZN(new_n352));
  INV_X1    g166(.A(G902), .ZN(new_n353));
  XNOR2_X1  g167(.A(G110), .B(G140), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n187), .A2(G227), .ZN(new_n355));
  XNOR2_X1  g169(.A(new_n354), .B(new_n355), .ZN(new_n356));
  INV_X1    g170(.A(G104), .ZN(new_n357));
  OAI21_X1  g171(.A(KEYINPUT3), .B1(new_n357), .B2(G107), .ZN(new_n358));
  INV_X1    g172(.A(KEYINPUT3), .ZN(new_n359));
  INV_X1    g173(.A(G107), .ZN(new_n360));
  NAND3_X1  g174(.A1(new_n359), .A2(new_n360), .A3(G104), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n357), .A2(G107), .ZN(new_n362));
  NAND4_X1  g176(.A1(new_n358), .A2(new_n361), .A3(new_n318), .A4(new_n362), .ZN(new_n363));
  NOR2_X1   g177(.A1(new_n357), .A2(G107), .ZN(new_n364));
  NOR2_X1   g178(.A1(new_n360), .A2(G104), .ZN(new_n365));
  OAI21_X1  g179(.A(G101), .B1(new_n364), .B2(new_n365), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n363), .A2(new_n366), .ZN(new_n367));
  NAND3_X1  g181(.A1(new_n367), .A2(new_n269), .A3(new_n275), .ZN(new_n368));
  INV_X1    g182(.A(new_n368), .ZN(new_n369));
  OAI21_X1  g183(.A(new_n270), .B1(new_n273), .B2(new_n274), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n263), .A2(KEYINPUT1), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n371), .A2(G128), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n370), .A2(new_n372), .ZN(new_n373));
  AOI21_X1  g187(.A(new_n367), .B1(new_n373), .B2(new_n275), .ZN(new_n374));
  OAI211_X1 g188(.A(KEYINPUT12), .B(new_n298), .C1(new_n369), .C2(new_n374), .ZN(new_n375));
  INV_X1    g189(.A(KEYINPUT82), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n375), .A2(new_n376), .ZN(new_n377));
  OAI21_X1  g191(.A(new_n298), .B1(new_n369), .B2(new_n374), .ZN(new_n378));
  INV_X1    g192(.A(KEYINPUT12), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n378), .A2(new_n379), .ZN(new_n380));
  AND2_X1   g194(.A1(new_n363), .A2(new_n366), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n265), .A2(KEYINPUT64), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n382), .A2(new_n263), .ZN(new_n383));
  AOI22_X1  g197(.A1(new_n383), .A2(new_n270), .B1(G128), .B2(new_n371), .ZN(new_n384));
  INV_X1    g198(.A(new_n275), .ZN(new_n385));
  OAI21_X1  g199(.A(new_n381), .B1(new_n384), .B2(new_n385), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n386), .A2(new_n368), .ZN(new_n387));
  NAND4_X1  g201(.A1(new_n387), .A2(KEYINPUT82), .A3(KEYINPUT12), .A4(new_n298), .ZN(new_n388));
  NAND3_X1  g202(.A1(new_n377), .A2(new_n380), .A3(new_n388), .ZN(new_n389));
  OAI211_X1 g203(.A(KEYINPUT10), .B(new_n381), .C1(new_n302), .C2(new_n303), .ZN(new_n390));
  INV_X1    g204(.A(KEYINPUT10), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n386), .A2(new_n391), .ZN(new_n392));
  NAND3_X1  g206(.A1(new_n358), .A2(new_n361), .A3(new_n362), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n393), .A2(G101), .ZN(new_n394));
  INV_X1    g208(.A(KEYINPUT81), .ZN(new_n395));
  NAND4_X1  g209(.A1(new_n394), .A2(new_n395), .A3(KEYINPUT4), .A4(new_n363), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n395), .A2(KEYINPUT4), .ZN(new_n397));
  NAND3_X1  g211(.A1(new_n393), .A2(G101), .A3(new_n397), .ZN(new_n398));
  NAND3_X1  g212(.A1(new_n305), .A2(new_n396), .A3(new_n398), .ZN(new_n399));
  INV_X1    g213(.A(new_n298), .ZN(new_n400));
  NAND4_X1  g214(.A1(new_n390), .A2(new_n392), .A3(new_n399), .A4(new_n400), .ZN(new_n401));
  AOI21_X1  g215(.A(new_n356), .B1(new_n389), .B2(new_n401), .ZN(new_n402));
  NAND3_X1  g216(.A1(new_n390), .A2(new_n392), .A3(new_n399), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n403), .A2(new_n298), .ZN(new_n404));
  AND3_X1   g218(.A1(new_n404), .A2(new_n401), .A3(new_n356), .ZN(new_n405));
  OAI21_X1  g219(.A(new_n353), .B1(new_n402), .B2(new_n405), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n406), .A2(G469), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n404), .A2(new_n401), .ZN(new_n408));
  INV_X1    g222(.A(new_n356), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n408), .A2(new_n409), .ZN(new_n410));
  NAND3_X1  g224(.A1(new_n389), .A2(new_n401), .A3(new_n356), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n410), .A2(new_n411), .ZN(new_n412));
  INV_X1    g226(.A(G469), .ZN(new_n413));
  NAND3_X1  g227(.A1(new_n412), .A2(new_n413), .A3(new_n224), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n407), .A2(new_n414), .ZN(new_n415));
  INV_X1    g229(.A(KEYINPUT83), .ZN(new_n416));
  NOR2_X1   g230(.A1(new_n415), .A2(new_n416), .ZN(new_n417));
  XOR2_X1   g231(.A(KEYINPUT9), .B(G234), .Z(new_n418));
  INV_X1    g232(.A(new_n418), .ZN(new_n419));
  OAI21_X1  g233(.A(G221), .B1(new_n419), .B2(G902), .ZN(new_n420));
  OAI21_X1  g234(.A(new_n420), .B1(new_n407), .B2(KEYINPUT83), .ZN(new_n421));
  NOR2_X1   g235(.A1(new_n417), .A2(new_n421), .ZN(new_n422));
  NAND3_X1  g236(.A1(new_n316), .A2(G214), .A3(new_n187), .ZN(new_n423));
  NOR2_X1   g237(.A1(new_n423), .A2(new_n264), .ZN(new_n424));
  INV_X1    g238(.A(new_n424), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n423), .A2(new_n264), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n425), .A2(new_n426), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n427), .A2(G131), .ZN(new_n428));
  INV_X1    g242(.A(KEYINPUT17), .ZN(new_n429));
  NAND3_X1  g243(.A1(new_n425), .A2(new_n247), .A3(new_n426), .ZN(new_n430));
  NAND3_X1  g244(.A1(new_n428), .A2(new_n429), .A3(new_n430), .ZN(new_n431));
  NOR2_X1   g245(.A1(new_n217), .A2(new_n200), .ZN(new_n432));
  AOI21_X1  g246(.A(new_n247), .B1(new_n425), .B2(new_n426), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n433), .A2(KEYINPUT17), .ZN(new_n434));
  NAND3_X1  g248(.A1(new_n431), .A2(new_n432), .A3(new_n434), .ZN(new_n435));
  NAND3_X1  g249(.A1(new_n427), .A2(KEYINPUT18), .A3(G131), .ZN(new_n436));
  INV_X1    g250(.A(KEYINPUT87), .ZN(new_n437));
  OAI21_X1  g251(.A(new_n437), .B1(new_n199), .B2(new_n192), .ZN(new_n438));
  NAND3_X1  g252(.A1(new_n198), .A2(KEYINPUT87), .A3(G146), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n438), .A2(new_n439), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n202), .A2(KEYINPUT86), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n440), .A2(new_n441), .ZN(new_n442));
  INV_X1    g256(.A(KEYINPUT18), .ZN(new_n443));
  OAI211_X1 g257(.A(new_n425), .B(new_n426), .C1(new_n443), .C2(new_n247), .ZN(new_n444));
  OR2_X1    g258(.A1(new_n440), .A2(new_n441), .ZN(new_n445));
  NAND4_X1  g259(.A1(new_n436), .A2(new_n442), .A3(new_n444), .A4(new_n445), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n435), .A2(new_n446), .ZN(new_n447));
  XNOR2_X1  g261(.A(G113), .B(G122), .ZN(new_n448));
  XNOR2_X1  g262(.A(new_n448), .B(new_n357), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n447), .A2(new_n449), .ZN(new_n450));
  INV_X1    g264(.A(KEYINPUT20), .ZN(new_n451));
  INV_X1    g265(.A(KEYINPUT88), .ZN(new_n452));
  OR2_X1    g266(.A1(new_n198), .A2(KEYINPUT19), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n198), .A2(KEYINPUT19), .ZN(new_n454));
  NAND3_X1  g268(.A1(new_n453), .A2(new_n192), .A3(new_n454), .ZN(new_n455));
  AOI21_X1  g269(.A(new_n200), .B1(new_n452), .B2(new_n455), .ZN(new_n456));
  AND2_X1   g270(.A1(new_n453), .A2(new_n454), .ZN(new_n457));
  NAND3_X1  g271(.A1(new_n457), .A2(KEYINPUT88), .A3(new_n192), .ZN(new_n458));
  INV_X1    g272(.A(new_n426), .ZN(new_n459));
  NOR3_X1   g273(.A1(new_n459), .A2(new_n424), .A3(G131), .ZN(new_n460));
  OAI211_X1 g274(.A(new_n456), .B(new_n458), .C1(new_n433), .C2(new_n460), .ZN(new_n461));
  INV_X1    g275(.A(new_n449), .ZN(new_n462));
  NAND3_X1  g276(.A1(new_n446), .A2(new_n461), .A3(new_n462), .ZN(new_n463));
  NOR2_X1   g277(.A1(G475), .A2(G902), .ZN(new_n464));
  INV_X1    g278(.A(new_n464), .ZN(new_n465));
  OR2_X1    g279(.A1(new_n465), .A2(KEYINPUT89), .ZN(new_n466));
  NAND4_X1  g280(.A1(new_n450), .A2(new_n451), .A3(new_n463), .A4(new_n466), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n465), .A2(KEYINPUT89), .ZN(new_n468));
  INV_X1    g282(.A(new_n468), .ZN(new_n469));
  AOI21_X1  g283(.A(new_n462), .B1(new_n435), .B2(new_n446), .ZN(new_n470));
  AND3_X1   g284(.A1(new_n446), .A2(new_n462), .A3(new_n461), .ZN(new_n471));
  NOR3_X1   g285(.A1(new_n470), .A2(new_n471), .A3(new_n465), .ZN(new_n472));
  XOR2_X1   g286(.A(KEYINPUT85), .B(KEYINPUT20), .Z(new_n473));
  INV_X1    g287(.A(new_n473), .ZN(new_n474));
  OAI22_X1  g288(.A1(new_n467), .A2(new_n469), .B1(new_n472), .B2(new_n474), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n462), .A2(KEYINPUT90), .ZN(new_n476));
  AOI21_X1  g290(.A(G902), .B1(new_n447), .B2(new_n476), .ZN(new_n477));
  OAI21_X1  g291(.A(new_n477), .B1(new_n447), .B2(new_n476), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n478), .A2(G475), .ZN(new_n479));
  AND2_X1   g293(.A1(new_n475), .A2(new_n479), .ZN(new_n480));
  OAI21_X1  g294(.A(G214), .B1(G237), .B2(G902), .ZN(new_n481));
  INV_X1    g295(.A(new_n481), .ZN(new_n482));
  NAND3_X1  g296(.A1(new_n396), .A2(new_n244), .A3(new_n398), .ZN(new_n483));
  INV_X1    g297(.A(KEYINPUT84), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  INV_X1    g299(.A(KEYINPUT5), .ZN(new_n486));
  NAND3_X1  g300(.A1(new_n486), .A2(new_n208), .A3(G116), .ZN(new_n487));
  OAI211_X1 g301(.A(G113), .B(new_n487), .C1(new_n242), .C2(new_n486), .ZN(new_n488));
  OAI21_X1  g302(.A(new_n488), .B1(new_n243), .B2(new_n242), .ZN(new_n489));
  OR2_X1    g303(.A1(new_n489), .A2(new_n367), .ZN(new_n490));
  NAND4_X1  g304(.A1(new_n396), .A2(new_n244), .A3(KEYINPUT84), .A4(new_n398), .ZN(new_n491));
  NAND3_X1  g305(.A1(new_n485), .A2(new_n490), .A3(new_n491), .ZN(new_n492));
  XNOR2_X1  g306(.A(G110), .B(G122), .ZN(new_n493));
  INV_X1    g307(.A(new_n493), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n492), .A2(new_n494), .ZN(new_n495));
  NAND4_X1  g309(.A1(new_n485), .A2(new_n490), .A3(new_n493), .A4(new_n491), .ZN(new_n496));
  NAND3_X1  g310(.A1(new_n495), .A2(KEYINPUT6), .A3(new_n496), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n290), .A2(G125), .ZN(new_n498));
  OAI21_X1  g312(.A(new_n498), .B1(G125), .B2(new_n281), .ZN(new_n499));
  NAND3_X1  g313(.A1(new_n499), .A2(G224), .A3(new_n187), .ZN(new_n500));
  INV_X1    g314(.A(new_n500), .ZN(new_n501));
  AOI21_X1  g315(.A(new_n499), .B1(G224), .B2(new_n187), .ZN(new_n502));
  OR2_X1    g316(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  INV_X1    g317(.A(KEYINPUT6), .ZN(new_n504));
  NAND3_X1  g318(.A1(new_n492), .A2(new_n504), .A3(new_n494), .ZN(new_n505));
  NAND3_X1  g319(.A1(new_n497), .A2(new_n503), .A3(new_n505), .ZN(new_n506));
  XOR2_X1   g320(.A(new_n493), .B(KEYINPUT8), .Z(new_n507));
  NAND2_X1  g321(.A1(new_n489), .A2(new_n367), .ZN(new_n508));
  AOI21_X1  g322(.A(new_n507), .B1(new_n490), .B2(new_n508), .ZN(new_n509));
  INV_X1    g323(.A(KEYINPUT7), .ZN(new_n510));
  AOI21_X1  g324(.A(new_n509), .B1(new_n510), .B2(new_n499), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n502), .A2(KEYINPUT7), .ZN(new_n512));
  NAND4_X1  g326(.A1(new_n511), .A2(new_n500), .A3(new_n496), .A4(new_n512), .ZN(new_n513));
  NAND3_X1  g327(.A1(new_n506), .A2(new_n353), .A3(new_n513), .ZN(new_n514));
  OAI21_X1  g328(.A(G210), .B1(G237), .B2(G902), .ZN(new_n515));
  INV_X1    g329(.A(new_n515), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n514), .A2(new_n516), .ZN(new_n517));
  NAND4_X1  g331(.A1(new_n506), .A2(new_n513), .A3(new_n353), .A4(new_n515), .ZN(new_n518));
  AOI21_X1  g332(.A(new_n482), .B1(new_n517), .B2(new_n518), .ZN(new_n519));
  NAND2_X1  g333(.A1(G234), .A2(G237), .ZN(new_n520));
  AND3_X1   g334(.A1(new_n520), .A2(G952), .A3(new_n187), .ZN(new_n521));
  AND3_X1   g335(.A1(new_n223), .A2(G953), .A3(new_n520), .ZN(new_n522));
  XOR2_X1   g336(.A(KEYINPUT21), .B(G898), .Z(new_n523));
  INV_X1    g337(.A(new_n523), .ZN(new_n524));
  AOI21_X1  g338(.A(new_n521), .B1(new_n522), .B2(new_n524), .ZN(new_n525));
  INV_X1    g339(.A(new_n525), .ZN(new_n526));
  XNOR2_X1  g340(.A(KEYINPUT91), .B(G122), .ZN(new_n527));
  INV_X1    g341(.A(G116), .ZN(new_n528));
  NOR2_X1   g342(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  INV_X1    g343(.A(KEYINPUT14), .ZN(new_n530));
  NOR3_X1   g344(.A1(new_n529), .A2(new_n530), .A3(new_n360), .ZN(new_n531));
  NOR2_X1   g345(.A1(new_n203), .A2(G143), .ZN(new_n532));
  AOI211_X1 g346(.A(G134), .B(new_n532), .C1(new_n205), .C2(G143), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n205), .A2(G143), .ZN(new_n534));
  INV_X1    g348(.A(new_n532), .ZN(new_n535));
  AOI21_X1  g349(.A(new_n252), .B1(new_n534), .B2(new_n535), .ZN(new_n536));
  OAI21_X1  g350(.A(new_n531), .B1(new_n533), .B2(new_n536), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n528), .A2(G122), .ZN(new_n538));
  INV_X1    g352(.A(new_n538), .ZN(new_n539));
  OAI21_X1  g353(.A(new_n360), .B1(new_n529), .B2(new_n539), .ZN(new_n540));
  OAI211_X1 g354(.A(G107), .B(new_n538), .C1(new_n527), .C2(new_n528), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  INV_X1    g356(.A(new_n542), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n532), .A2(KEYINPUT13), .ZN(new_n544));
  XOR2_X1   g358(.A(new_n544), .B(KEYINPUT92), .Z(new_n545));
  NAND2_X1  g359(.A1(new_n534), .A2(KEYINPUT13), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n546), .A2(new_n535), .ZN(new_n547));
  AOI21_X1  g361(.A(new_n252), .B1(new_n545), .B2(new_n547), .ZN(new_n548));
  OAI211_X1 g362(.A(new_n537), .B(new_n543), .C1(new_n548), .C2(new_n533), .ZN(new_n549));
  NOR2_X1   g363(.A1(new_n536), .A2(new_n533), .ZN(new_n550));
  OAI21_X1  g364(.A(new_n542), .B1(new_n550), .B2(new_n531), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n549), .A2(new_n551), .ZN(new_n552));
  NAND3_X1  g366(.A1(new_n418), .A2(G217), .A3(new_n187), .ZN(new_n553));
  INV_X1    g367(.A(new_n553), .ZN(new_n554));
  XNOR2_X1  g368(.A(new_n552), .B(new_n554), .ZN(new_n555));
  INV_X1    g369(.A(KEYINPUT15), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n556), .A2(G478), .ZN(new_n557));
  NAND3_X1  g371(.A1(new_n555), .A2(new_n224), .A3(new_n557), .ZN(new_n558));
  INV_X1    g372(.A(new_n558), .ZN(new_n559));
  AOI21_X1  g373(.A(new_n557), .B1(new_n555), .B2(new_n224), .ZN(new_n560));
  NOR2_X1   g374(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  NAND4_X1  g375(.A1(new_n480), .A2(new_n519), .A3(new_n526), .A4(new_n561), .ZN(new_n562));
  INV_X1    g376(.A(new_n562), .ZN(new_n563));
  NAND4_X1  g377(.A1(new_n241), .A2(new_n352), .A3(new_n422), .A4(new_n563), .ZN(new_n564));
  XNOR2_X1  g378(.A(new_n564), .B(G101), .ZN(G3));
  INV_X1    g379(.A(G472), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n338), .A2(new_n224), .ZN(new_n567));
  INV_X1    g381(.A(KEYINPUT93), .ZN(new_n568));
  AOI21_X1  g382(.A(new_n566), .B1(new_n567), .B2(new_n568), .ZN(new_n569));
  NAND3_X1  g383(.A1(new_n338), .A2(KEYINPUT93), .A3(new_n224), .ZN(new_n570));
  AOI22_X1  g384(.A1(new_n569), .A2(new_n570), .B1(new_n339), .B2(new_n338), .ZN(new_n571));
  NAND3_X1  g385(.A1(new_n571), .A2(new_n241), .A3(new_n422), .ZN(new_n572));
  INV_X1    g386(.A(new_n572), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n519), .A2(new_n526), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n475), .A2(new_n479), .ZN(new_n575));
  INV_X1    g389(.A(KEYINPUT33), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n555), .A2(new_n576), .ZN(new_n577));
  NOR2_X1   g391(.A1(new_n552), .A2(new_n554), .ZN(new_n578));
  AOI21_X1  g392(.A(new_n553), .B1(new_n549), .B2(new_n551), .ZN(new_n579));
  NOR2_X1   g393(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n580), .A2(KEYINPUT33), .ZN(new_n581));
  NAND4_X1  g395(.A1(new_n577), .A2(new_n581), .A3(G478), .A4(new_n224), .ZN(new_n582));
  XNOR2_X1  g396(.A(KEYINPUT94), .B(G478), .ZN(new_n583));
  OAI21_X1  g397(.A(new_n583), .B1(new_n580), .B2(new_n223), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n582), .A2(new_n584), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n575), .A2(new_n585), .ZN(new_n586));
  NOR2_X1   g400(.A1(new_n574), .A2(new_n586), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n573), .A2(new_n587), .ZN(new_n588));
  XNOR2_X1  g402(.A(new_n588), .B(KEYINPUT95), .ZN(new_n589));
  XOR2_X1   g403(.A(KEYINPUT34), .B(G104), .Z(new_n590));
  XNOR2_X1  g404(.A(new_n589), .B(new_n590), .ZN(G6));
  AND2_X1   g405(.A1(new_n472), .A2(new_n474), .ZN(new_n592));
  NOR2_X1   g406(.A1(new_n472), .A2(new_n474), .ZN(new_n593));
  OAI21_X1  g407(.A(new_n479), .B1(new_n592), .B2(new_n593), .ZN(new_n594));
  NOR3_X1   g408(.A1(new_n574), .A2(new_n561), .A3(new_n594), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n573), .A2(new_n595), .ZN(new_n596));
  XOR2_X1   g410(.A(KEYINPUT35), .B(G107), .Z(new_n597));
  XNOR2_X1  g411(.A(new_n596), .B(new_n597), .ZN(G9));
  NAND2_X1  g412(.A1(new_n213), .A2(new_n218), .ZN(new_n599));
  NOR2_X1   g413(.A1(new_n191), .A2(KEYINPUT36), .ZN(new_n600));
  XNOR2_X1  g414(.A(new_n599), .B(new_n600), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n601), .A2(new_n238), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n237), .A2(new_n602), .ZN(new_n603));
  NAND4_X1  g417(.A1(new_n571), .A2(new_n422), .A3(new_n563), .A4(new_n603), .ZN(new_n604));
  XOR2_X1   g418(.A(KEYINPUT37), .B(G110), .Z(new_n605));
  XNOR2_X1  g419(.A(new_n604), .B(new_n605), .ZN(G12));
  INV_X1    g420(.A(new_n603), .ZN(new_n607));
  INV_X1    g421(.A(new_n519), .ZN(new_n608));
  NOR2_X1   g422(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  INV_X1    g423(.A(G900), .ZN(new_n610));
  AOI21_X1  g424(.A(new_n521), .B1(new_n522), .B2(new_n610), .ZN(new_n611));
  NOR3_X1   g425(.A1(new_n594), .A2(new_n561), .A3(new_n611), .ZN(new_n612));
  NAND4_X1  g426(.A1(new_n352), .A2(new_n609), .A3(new_n422), .A4(new_n612), .ZN(new_n613));
  XNOR2_X1  g427(.A(new_n613), .B(G128), .ZN(G30));
  XNOR2_X1  g428(.A(new_n611), .B(KEYINPUT39), .ZN(new_n615));
  NOR3_X1   g429(.A1(new_n417), .A2(new_n421), .A3(new_n615), .ZN(new_n616));
  XNOR2_X1  g430(.A(new_n616), .B(KEYINPUT96), .ZN(new_n617));
  XNOR2_X1  g431(.A(new_n617), .B(KEYINPUT40), .ZN(new_n618));
  AOI21_X1  g432(.A(new_n322), .B1(new_n332), .B2(new_n333), .ZN(new_n619));
  OAI21_X1  g433(.A(new_n353), .B1(new_n347), .B2(new_n321), .ZN(new_n620));
  OAI21_X1  g434(.A(G472), .B1(new_n619), .B2(new_n620), .ZN(new_n621));
  NAND3_X1  g435(.A1(new_n342), .A2(new_n343), .A3(new_n621), .ZN(new_n622));
  INV_X1    g436(.A(new_n622), .ZN(new_n623));
  NOR2_X1   g437(.A1(new_n623), .A2(new_n603), .ZN(new_n624));
  AOI21_X1  g438(.A(new_n482), .B1(new_n475), .B2(new_n479), .ZN(new_n625));
  INV_X1    g439(.A(new_n561), .ZN(new_n626));
  AND2_X1   g440(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n517), .A2(new_n518), .ZN(new_n628));
  XNOR2_X1  g442(.A(new_n628), .B(KEYINPUT38), .ZN(new_n629));
  NAND4_X1  g443(.A1(new_n618), .A2(new_n624), .A3(new_n627), .A4(new_n629), .ZN(new_n630));
  XNOR2_X1  g444(.A(new_n630), .B(G143), .ZN(G45));
  NOR2_X1   g445(.A1(new_n586), .A2(new_n611), .ZN(new_n632));
  NAND4_X1  g446(.A1(new_n352), .A2(new_n609), .A3(new_n422), .A4(new_n632), .ZN(new_n633));
  XNOR2_X1  g447(.A(KEYINPUT97), .B(G146), .ZN(new_n634));
  XNOR2_X1  g448(.A(new_n633), .B(new_n634), .ZN(G48));
  NAND2_X1  g449(.A1(new_n241), .A2(new_n352), .ZN(new_n636));
  INV_X1    g450(.A(new_n636), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n412), .A2(new_n224), .ZN(new_n638));
  NOR2_X1   g452(.A1(new_n413), .A2(KEYINPUT98), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  OAI211_X1 g454(.A(new_n412), .B(new_n224), .C1(KEYINPUT98), .C2(new_n413), .ZN(new_n641));
  AND2_X1   g455(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n642), .A2(new_n420), .ZN(new_n643));
  INV_X1    g457(.A(new_n643), .ZN(new_n644));
  NAND3_X1  g458(.A1(new_n637), .A2(new_n587), .A3(new_n644), .ZN(new_n645));
  XNOR2_X1  g459(.A(new_n645), .B(KEYINPUT99), .ZN(new_n646));
  XOR2_X1   g460(.A(KEYINPUT41), .B(G113), .Z(new_n647));
  XNOR2_X1  g461(.A(new_n646), .B(new_n647), .ZN(G15));
  NAND3_X1  g462(.A1(new_n637), .A2(new_n595), .A3(new_n644), .ZN(new_n649));
  XNOR2_X1  g463(.A(new_n649), .B(G116), .ZN(G18));
  NAND2_X1  g464(.A1(new_n480), .A2(new_n561), .ZN(new_n651));
  NOR2_X1   g465(.A1(new_n651), .A2(new_n643), .ZN(new_n652));
  NAND4_X1  g466(.A1(new_n352), .A2(new_n652), .A3(new_n526), .A4(new_n609), .ZN(new_n653));
  XNOR2_X1  g467(.A(new_n653), .B(G119), .ZN(G21));
  OAI211_X1 g468(.A(new_n335), .B(new_n337), .C1(new_n321), .C2(new_n348), .ZN(new_n655));
  AOI22_X1  g469(.A1(new_n567), .A2(G472), .B1(new_n339), .B2(new_n655), .ZN(new_n656));
  INV_X1    g470(.A(new_n656), .ZN(new_n657));
  NOR2_X1   g471(.A1(new_n657), .A2(new_n240), .ZN(new_n658));
  NAND3_X1  g472(.A1(new_n625), .A2(new_n626), .A3(new_n628), .ZN(new_n659));
  INV_X1    g473(.A(new_n659), .ZN(new_n660));
  NAND4_X1  g474(.A1(new_n658), .A2(new_n526), .A3(new_n644), .A4(new_n660), .ZN(new_n661));
  XNOR2_X1  g475(.A(new_n661), .B(G122), .ZN(G24));
  NOR2_X1   g476(.A1(new_n643), .A2(new_n608), .ZN(new_n663));
  NAND4_X1  g477(.A1(new_n663), .A2(new_n656), .A3(new_n632), .A4(new_n603), .ZN(new_n664));
  XNOR2_X1  g478(.A(new_n664), .B(G125), .ZN(G27));
  INV_X1    g479(.A(new_n632), .ZN(new_n666));
  INV_X1    g480(.A(KEYINPUT100), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n415), .A2(new_n667), .ZN(new_n668));
  NAND3_X1  g482(.A1(new_n407), .A2(KEYINPUT100), .A3(new_n414), .ZN(new_n669));
  NAND3_X1  g483(.A1(new_n668), .A2(new_n420), .A3(new_n669), .ZN(new_n670));
  NAND2_X1  g484(.A1(new_n670), .A2(KEYINPUT101), .ZN(new_n671));
  NOR2_X1   g485(.A1(new_n628), .A2(new_n482), .ZN(new_n672));
  INV_X1    g486(.A(KEYINPUT101), .ZN(new_n673));
  NAND4_X1  g487(.A1(new_n668), .A2(new_n669), .A3(new_n673), .A4(new_n420), .ZN(new_n674));
  NAND3_X1  g488(.A1(new_n671), .A2(new_n672), .A3(new_n674), .ZN(new_n675));
  INV_X1    g489(.A(KEYINPUT102), .ZN(new_n676));
  NAND2_X1  g490(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  NAND4_X1  g491(.A1(new_n671), .A2(KEYINPUT102), .A3(new_n672), .A4(new_n674), .ZN(new_n678));
  AOI21_X1  g492(.A(new_n666), .B1(new_n677), .B2(new_n678), .ZN(new_n679));
  NAND2_X1  g493(.A1(new_n343), .A2(KEYINPUT103), .ZN(new_n680));
  INV_X1    g494(.A(KEYINPUT103), .ZN(new_n681));
  NAND4_X1  g495(.A1(new_n338), .A2(new_n681), .A3(KEYINPUT32), .A4(new_n339), .ZN(new_n682));
  NAND4_X1  g496(.A1(new_n680), .A2(new_n342), .A3(new_n351), .A4(new_n682), .ZN(new_n683));
  INV_X1    g497(.A(new_n240), .ZN(new_n684));
  NAND2_X1  g498(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  INV_X1    g499(.A(KEYINPUT42), .ZN(new_n686));
  NOR2_X1   g500(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  NAND2_X1  g501(.A1(new_n679), .A2(new_n687), .ZN(new_n688));
  INV_X1    g502(.A(new_n688), .ZN(new_n689));
  AOI21_X1  g503(.A(new_n636), .B1(new_n677), .B2(new_n678), .ZN(new_n690));
  AOI21_X1  g504(.A(KEYINPUT42), .B1(new_n690), .B2(new_n632), .ZN(new_n691));
  NOR2_X1   g505(.A1(new_n689), .A2(new_n691), .ZN(new_n692));
  XNOR2_X1  g506(.A(new_n692), .B(new_n247), .ZN(G33));
  NAND2_X1  g507(.A1(new_n677), .A2(new_n678), .ZN(new_n694));
  NAND3_X1  g508(.A1(new_n694), .A2(new_n637), .A3(new_n612), .ZN(new_n695));
  INV_X1    g509(.A(KEYINPUT104), .ZN(new_n696));
  NAND2_X1  g510(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  NAND3_X1  g511(.A1(new_n690), .A2(KEYINPUT104), .A3(new_n612), .ZN(new_n698));
  NAND2_X1  g512(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  XNOR2_X1  g513(.A(new_n699), .B(G134), .ZN(G36));
  NOR2_X1   g514(.A1(new_n571), .A2(new_n607), .ZN(new_n701));
  XOR2_X1   g515(.A(new_n701), .B(KEYINPUT107), .Z(new_n702));
  INV_X1    g516(.A(new_n585), .ZN(new_n703));
  NOR3_X1   g517(.A1(new_n703), .A2(KEYINPUT43), .A3(new_n575), .ZN(new_n704));
  XNOR2_X1  g518(.A(new_n480), .B(KEYINPUT106), .ZN(new_n705));
  NAND2_X1  g519(.A1(new_n705), .A2(new_n585), .ZN(new_n706));
  AOI21_X1  g520(.A(new_n704), .B1(new_n706), .B2(KEYINPUT43), .ZN(new_n707));
  NAND2_X1  g521(.A1(new_n702), .A2(new_n707), .ZN(new_n708));
  XNOR2_X1  g522(.A(new_n708), .B(KEYINPUT44), .ZN(new_n709));
  NAND2_X1  g523(.A1(new_n709), .A2(new_n672), .ZN(new_n710));
  NOR2_X1   g524(.A1(new_n402), .A2(new_n405), .ZN(new_n711));
  OAI21_X1  g525(.A(G469), .B1(new_n711), .B2(KEYINPUT45), .ZN(new_n712));
  XNOR2_X1  g526(.A(new_n712), .B(KEYINPUT105), .ZN(new_n713));
  NAND2_X1  g527(.A1(new_n711), .A2(KEYINPUT45), .ZN(new_n714));
  NAND2_X1  g528(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  NOR2_X1   g529(.A1(new_n413), .A2(new_n353), .ZN(new_n716));
  INV_X1    g530(.A(new_n716), .ZN(new_n717));
  NAND3_X1  g531(.A1(new_n715), .A2(KEYINPUT46), .A3(new_n717), .ZN(new_n718));
  NAND2_X1  g532(.A1(new_n718), .A2(new_n414), .ZN(new_n719));
  AOI21_X1  g533(.A(KEYINPUT46), .B1(new_n715), .B2(new_n717), .ZN(new_n720));
  OR2_X1    g534(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  INV_X1    g535(.A(new_n615), .ZN(new_n722));
  NAND3_X1  g536(.A1(new_n721), .A2(new_n420), .A3(new_n722), .ZN(new_n723));
  OR2_X1    g537(.A1(new_n710), .A2(new_n723), .ZN(new_n724));
  XOR2_X1   g538(.A(KEYINPUT108), .B(G137), .Z(new_n725));
  XNOR2_X1  g539(.A(new_n724), .B(new_n725), .ZN(G39));
  INV_X1    g540(.A(KEYINPUT47), .ZN(new_n727));
  NAND3_X1  g541(.A1(new_n721), .A2(new_n727), .A3(new_n420), .ZN(new_n728));
  INV_X1    g542(.A(new_n728), .ZN(new_n729));
  AOI21_X1  g543(.A(new_n727), .B1(new_n721), .B2(new_n420), .ZN(new_n730));
  NOR2_X1   g544(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  NOR4_X1   g545(.A1(new_n352), .A2(new_n241), .A3(new_n482), .A4(new_n628), .ZN(new_n732));
  AND3_X1   g546(.A1(new_n731), .A2(new_n632), .A3(new_n732), .ZN(new_n733));
  XNOR2_X1  g547(.A(new_n733), .B(new_n193), .ZN(G42));
  INV_X1    g548(.A(KEYINPUT53), .ZN(new_n735));
  NAND4_X1  g549(.A1(new_n645), .A2(new_n649), .A3(new_n653), .A4(new_n661), .ZN(new_n736));
  NAND2_X1  g550(.A1(new_n690), .A2(new_n632), .ZN(new_n737));
  NAND2_X1  g551(.A1(new_n737), .A2(new_n686), .ZN(new_n738));
  AOI21_X1  g552(.A(new_n736), .B1(new_n738), .B2(new_n688), .ZN(new_n739));
  NAND2_X1  g553(.A1(new_n703), .A2(new_n575), .ZN(new_n740));
  AND4_X1   g554(.A1(new_n526), .A2(new_n740), .A3(new_n651), .A4(new_n519), .ZN(new_n741));
  NAND4_X1  g555(.A1(new_n741), .A2(new_n571), .A3(new_n241), .A4(new_n422), .ZN(new_n742));
  NAND3_X1  g556(.A1(new_n742), .A2(new_n604), .A3(new_n564), .ZN(new_n743));
  INV_X1    g557(.A(KEYINPUT109), .ZN(new_n744));
  NAND2_X1  g558(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  NAND4_X1  g559(.A1(new_n742), .A2(new_n604), .A3(KEYINPUT109), .A4(new_n564), .ZN(new_n746));
  NAND2_X1  g560(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  AOI211_X1 g561(.A(new_n666), .B(new_n657), .C1(new_n677), .C2(new_n678), .ZN(new_n748));
  NAND3_X1  g562(.A1(new_n352), .A2(new_n422), .A3(new_n672), .ZN(new_n749));
  NOR4_X1   g563(.A1(new_n749), .A2(new_n626), .A3(new_n594), .A4(new_n611), .ZN(new_n750));
  OAI21_X1  g564(.A(new_n603), .B1(new_n748), .B2(new_n750), .ZN(new_n751));
  NAND4_X1  g565(.A1(new_n739), .A2(new_n699), .A3(new_n747), .A4(new_n751), .ZN(new_n752));
  AND2_X1   g566(.A1(new_n633), .A2(new_n664), .ZN(new_n753));
  INV_X1    g567(.A(KEYINPUT110), .ZN(new_n754));
  NOR2_X1   g568(.A1(new_n659), .A2(new_n670), .ZN(new_n755));
  INV_X1    g569(.A(new_n611), .ZN(new_n756));
  NAND4_X1  g570(.A1(new_n755), .A2(new_n622), .A3(new_n607), .A4(new_n756), .ZN(new_n757));
  NAND4_X1  g571(.A1(new_n753), .A2(new_n754), .A3(new_n613), .A4(new_n757), .ZN(new_n758));
  INV_X1    g572(.A(KEYINPUT52), .ZN(new_n759));
  NAND4_X1  g573(.A1(new_n757), .A2(new_n613), .A3(new_n633), .A4(new_n664), .ZN(new_n760));
  NAND2_X1  g574(.A1(new_n760), .A2(KEYINPUT110), .ZN(new_n761));
  AND3_X1   g575(.A1(new_n758), .A2(new_n759), .A3(new_n761), .ZN(new_n762));
  AOI21_X1  g576(.A(new_n759), .B1(new_n758), .B2(new_n761), .ZN(new_n763));
  OR2_X1    g577(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  OAI21_X1  g578(.A(new_n735), .B1(new_n752), .B2(new_n764), .ZN(new_n765));
  INV_X1    g579(.A(KEYINPUT113), .ZN(new_n766));
  AOI21_X1  g580(.A(new_n735), .B1(new_n739), .B2(new_n766), .ZN(new_n767));
  AND2_X1   g581(.A1(new_n760), .A2(KEYINPUT52), .ZN(new_n768));
  NOR2_X1   g582(.A1(new_n762), .A2(new_n768), .ZN(new_n769));
  AND3_X1   g583(.A1(new_n699), .A2(new_n747), .A3(new_n751), .ZN(new_n770));
  AND4_X1   g584(.A1(new_n645), .A2(new_n649), .A3(new_n653), .A4(new_n661), .ZN(new_n771));
  OAI21_X1  g585(.A(new_n771), .B1(new_n689), .B2(new_n691), .ZN(new_n772));
  NAND2_X1  g586(.A1(new_n772), .A2(KEYINPUT113), .ZN(new_n773));
  NAND4_X1  g587(.A1(new_n767), .A2(new_n769), .A3(new_n770), .A4(new_n773), .ZN(new_n774));
  INV_X1    g588(.A(KEYINPUT54), .ZN(new_n775));
  NAND3_X1  g589(.A1(new_n765), .A2(new_n774), .A3(new_n775), .ZN(new_n776));
  NAND2_X1  g590(.A1(new_n776), .A2(KEYINPUT114), .ZN(new_n777));
  INV_X1    g591(.A(KEYINPUT114), .ZN(new_n778));
  NAND4_X1  g592(.A1(new_n765), .A2(new_n774), .A3(new_n778), .A4(new_n775), .ZN(new_n779));
  NAND2_X1  g593(.A1(new_n777), .A2(new_n779), .ZN(new_n780));
  AND3_X1   g594(.A1(new_n644), .A2(new_n521), .A3(new_n672), .ZN(new_n781));
  AND2_X1   g595(.A1(new_n707), .A2(new_n781), .ZN(new_n782));
  INV_X1    g596(.A(new_n685), .ZN(new_n783));
  NAND2_X1  g597(.A1(new_n782), .A2(new_n783), .ZN(new_n784));
  XOR2_X1   g598(.A(new_n784), .B(KEYINPUT48), .Z(new_n785));
  NAND3_X1  g599(.A1(new_n707), .A2(new_n521), .A3(new_n658), .ZN(new_n786));
  INV_X1    g600(.A(new_n786), .ZN(new_n787));
  NAND2_X1  g601(.A1(new_n787), .A2(new_n663), .ZN(new_n788));
  INV_X1    g602(.A(G952), .ZN(new_n789));
  AND3_X1   g603(.A1(new_n781), .A2(new_n623), .A3(new_n241), .ZN(new_n790));
  INV_X1    g604(.A(new_n586), .ZN(new_n791));
  AOI211_X1 g605(.A(new_n789), .B(G953), .C1(new_n790), .C2(new_n791), .ZN(new_n792));
  NAND2_X1  g606(.A1(new_n788), .A2(new_n792), .ZN(new_n793));
  XNOR2_X1  g607(.A(new_n793), .B(KEYINPUT118), .ZN(new_n794));
  OR3_X1    g608(.A1(new_n629), .A2(new_n481), .A3(new_n643), .ZN(new_n795));
  INV_X1    g609(.A(new_n795), .ZN(new_n796));
  NAND3_X1  g610(.A1(new_n787), .A2(KEYINPUT50), .A3(new_n796), .ZN(new_n797));
  INV_X1    g611(.A(KEYINPUT50), .ZN(new_n798));
  OAI21_X1  g612(.A(new_n798), .B1(new_n786), .B2(new_n795), .ZN(new_n799));
  NOR2_X1   g613(.A1(new_n657), .A2(new_n607), .ZN(new_n800));
  AOI22_X1  g614(.A1(new_n797), .A2(new_n799), .B1(new_n800), .B2(new_n782), .ZN(new_n801));
  NAND3_X1  g615(.A1(new_n790), .A2(new_n480), .A3(new_n703), .ZN(new_n802));
  XNOR2_X1  g616(.A(new_n802), .B(KEYINPUT116), .ZN(new_n803));
  NAND2_X1  g617(.A1(new_n801), .A2(new_n803), .ZN(new_n804));
  NAND2_X1  g618(.A1(new_n804), .A2(KEYINPUT117), .ZN(new_n805));
  INV_X1    g619(.A(KEYINPUT117), .ZN(new_n806));
  OAI211_X1 g620(.A(new_n801), .B(new_n803), .C1(new_n806), .C2(KEYINPUT51), .ZN(new_n807));
  INV_X1    g621(.A(new_n642), .ZN(new_n808));
  OAI22_X1  g622(.A1(new_n729), .A2(new_n730), .B1(new_n420), .B2(new_n808), .ZN(new_n809));
  NAND3_X1  g623(.A1(new_n809), .A2(new_n672), .A3(new_n787), .ZN(new_n810));
  NAND2_X1  g624(.A1(new_n810), .A2(KEYINPUT115), .ZN(new_n811));
  INV_X1    g625(.A(KEYINPUT115), .ZN(new_n812));
  NAND4_X1  g626(.A1(new_n809), .A2(new_n812), .A3(new_n672), .A4(new_n787), .ZN(new_n813));
  NAND4_X1  g627(.A1(new_n805), .A2(new_n807), .A3(new_n811), .A4(new_n813), .ZN(new_n814));
  INV_X1    g628(.A(new_n810), .ZN(new_n815));
  OAI21_X1  g629(.A(KEYINPUT51), .B1(new_n807), .B2(new_n815), .ZN(new_n816));
  AOI211_X1 g630(.A(new_n785), .B(new_n794), .C1(new_n814), .C2(new_n816), .ZN(new_n817));
  NOR2_X1   g631(.A1(new_n762), .A2(new_n763), .ZN(new_n818));
  NAND4_X1  g632(.A1(new_n770), .A2(KEYINPUT53), .A3(new_n818), .A4(new_n739), .ZN(new_n819));
  NAND2_X1  g633(.A1(new_n819), .A2(KEYINPUT111), .ZN(new_n820));
  INV_X1    g634(.A(new_n769), .ZN(new_n821));
  OAI21_X1  g635(.A(new_n735), .B1(new_n821), .B2(new_n752), .ZN(new_n822));
  NAND3_X1  g636(.A1(new_n699), .A2(new_n747), .A3(new_n751), .ZN(new_n823));
  NOR2_X1   g637(.A1(new_n823), .A2(new_n772), .ZN(new_n824));
  INV_X1    g638(.A(KEYINPUT111), .ZN(new_n825));
  NAND4_X1  g639(.A1(new_n824), .A2(new_n825), .A3(KEYINPUT53), .A4(new_n818), .ZN(new_n826));
  NAND3_X1  g640(.A1(new_n820), .A2(new_n822), .A3(new_n826), .ZN(new_n827));
  AND3_X1   g641(.A1(new_n827), .A2(KEYINPUT112), .A3(KEYINPUT54), .ZN(new_n828));
  AOI21_X1  g642(.A(KEYINPUT112), .B1(new_n827), .B2(KEYINPUT54), .ZN(new_n829));
  OAI211_X1 g643(.A(new_n780), .B(new_n817), .C1(new_n828), .C2(new_n829), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n789), .A2(new_n187), .ZN(new_n831));
  NAND2_X1  g645(.A1(new_n830), .A2(new_n831), .ZN(new_n832));
  OR2_X1    g646(.A1(new_n808), .A2(KEYINPUT49), .ZN(new_n833));
  NAND2_X1  g647(.A1(new_n808), .A2(KEYINPUT49), .ZN(new_n834));
  NAND3_X1  g648(.A1(new_n833), .A2(new_n684), .A3(new_n834), .ZN(new_n835));
  NOR3_X1   g649(.A1(new_n706), .A2(new_n835), .A3(new_n629), .ZN(new_n836));
  NAND4_X1  g650(.A1(new_n836), .A2(new_n420), .A3(new_n623), .A4(new_n481), .ZN(new_n837));
  NAND2_X1  g651(.A1(new_n832), .A2(new_n837), .ZN(new_n838));
  NAND2_X1  g652(.A1(new_n838), .A2(KEYINPUT119), .ZN(new_n839));
  INV_X1    g653(.A(KEYINPUT119), .ZN(new_n840));
  NAND3_X1  g654(.A1(new_n832), .A2(new_n840), .A3(new_n837), .ZN(new_n841));
  NAND2_X1  g655(.A1(new_n839), .A2(new_n841), .ZN(G75));
  AOI21_X1  g656(.A(new_n224), .B1(new_n765), .B2(new_n774), .ZN(new_n843));
  AOI21_X1  g657(.A(KEYINPUT56), .B1(new_n843), .B2(new_n516), .ZN(new_n844));
  NAND2_X1  g658(.A1(new_n497), .A2(new_n505), .ZN(new_n845));
  XNOR2_X1  g659(.A(new_n845), .B(new_n503), .ZN(new_n846));
  XNOR2_X1  g660(.A(new_n846), .B(KEYINPUT55), .ZN(new_n847));
  XNOR2_X1  g661(.A(new_n844), .B(new_n847), .ZN(new_n848));
  NOR2_X1   g662(.A1(new_n187), .A2(G952), .ZN(new_n849));
  NOR2_X1   g663(.A1(new_n848), .A2(new_n849), .ZN(G51));
  AND3_X1   g664(.A1(new_n765), .A2(new_n774), .A3(new_n775), .ZN(new_n851));
  AOI21_X1  g665(.A(new_n775), .B1(new_n765), .B2(new_n774), .ZN(new_n852));
  NOR2_X1   g666(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  XOR2_X1   g667(.A(new_n716), .B(KEYINPUT57), .Z(new_n854));
  OR3_X1    g668(.A1(new_n853), .A2(KEYINPUT120), .A3(new_n854), .ZN(new_n855));
  OAI21_X1  g669(.A(KEYINPUT120), .B1(new_n853), .B2(new_n854), .ZN(new_n856));
  NAND3_X1  g670(.A1(new_n855), .A2(new_n412), .A3(new_n856), .ZN(new_n857));
  NAND3_X1  g671(.A1(new_n843), .A2(new_n714), .A3(new_n713), .ZN(new_n858));
  AOI21_X1  g672(.A(new_n849), .B1(new_n857), .B2(new_n858), .ZN(G54));
  AND3_X1   g673(.A1(new_n843), .A2(KEYINPUT58), .A3(G475), .ZN(new_n860));
  NOR2_X1   g674(.A1(new_n470), .A2(new_n471), .ZN(new_n861));
  OR2_X1    g675(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  INV_X1    g676(.A(new_n849), .ZN(new_n863));
  NAND2_X1  g677(.A1(new_n860), .A2(new_n861), .ZN(new_n864));
  NAND3_X1  g678(.A1(new_n862), .A2(new_n863), .A3(new_n864), .ZN(new_n865));
  INV_X1    g679(.A(KEYINPUT121), .ZN(new_n866));
  XNOR2_X1  g680(.A(new_n865), .B(new_n866), .ZN(G60));
  NAND2_X1  g681(.A1(new_n577), .A2(new_n581), .ZN(new_n868));
  INV_X1    g682(.A(new_n868), .ZN(new_n869));
  OAI21_X1  g683(.A(new_n780), .B1(new_n828), .B2(new_n829), .ZN(new_n870));
  NAND2_X1  g684(.A1(G478), .A2(G902), .ZN(new_n871));
  XOR2_X1   g685(.A(new_n871), .B(KEYINPUT59), .Z(new_n872));
  INV_X1    g686(.A(new_n872), .ZN(new_n873));
  AOI21_X1  g687(.A(new_n869), .B1(new_n870), .B2(new_n873), .ZN(new_n874));
  INV_X1    g688(.A(KEYINPUT122), .ZN(new_n875));
  NAND2_X1  g689(.A1(new_n765), .A2(new_n774), .ZN(new_n876));
  NAND2_X1  g690(.A1(new_n876), .A2(KEYINPUT54), .ZN(new_n877));
  AOI21_X1  g691(.A(new_n868), .B1(new_n877), .B2(new_n776), .ZN(new_n878));
  AOI21_X1  g692(.A(new_n875), .B1(new_n878), .B2(new_n873), .ZN(new_n879));
  OAI211_X1 g693(.A(new_n869), .B(new_n873), .C1(new_n851), .C2(new_n852), .ZN(new_n880));
  NOR2_X1   g694(.A1(new_n880), .A2(KEYINPUT122), .ZN(new_n881));
  OAI21_X1  g695(.A(new_n863), .B1(new_n879), .B2(new_n881), .ZN(new_n882));
  OAI21_X1  g696(.A(KEYINPUT123), .B1(new_n874), .B2(new_n882), .ZN(new_n883));
  INV_X1    g697(.A(KEYINPUT123), .ZN(new_n884));
  NAND3_X1  g698(.A1(new_n878), .A2(new_n875), .A3(new_n873), .ZN(new_n885));
  NAND2_X1  g699(.A1(new_n880), .A2(KEYINPUT122), .ZN(new_n886));
  AOI21_X1  g700(.A(new_n849), .B1(new_n885), .B2(new_n886), .ZN(new_n887));
  NAND2_X1  g701(.A1(new_n827), .A2(KEYINPUT54), .ZN(new_n888));
  INV_X1    g702(.A(KEYINPUT112), .ZN(new_n889));
  NAND2_X1  g703(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  NAND3_X1  g704(.A1(new_n827), .A2(KEYINPUT112), .A3(KEYINPUT54), .ZN(new_n891));
  NAND2_X1  g705(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  AOI21_X1  g706(.A(new_n872), .B1(new_n892), .B2(new_n780), .ZN(new_n893));
  OAI211_X1 g707(.A(new_n884), .B(new_n887), .C1(new_n893), .C2(new_n869), .ZN(new_n894));
  NAND2_X1  g708(.A1(new_n883), .A2(new_n894), .ZN(G63));
  NAND2_X1  g709(.A1(G217), .A2(G902), .ZN(new_n896));
  XOR2_X1   g710(.A(new_n896), .B(KEYINPUT124), .Z(new_n897));
  XNOR2_X1  g711(.A(new_n897), .B(KEYINPUT60), .ZN(new_n898));
  AOI21_X1  g712(.A(new_n898), .B1(new_n765), .B2(new_n774), .ZN(new_n899));
  NAND2_X1  g713(.A1(new_n899), .A2(new_n601), .ZN(new_n900));
  OAI211_X1 g714(.A(new_n900), .B(new_n863), .C1(new_n222), .C2(new_n899), .ZN(new_n901));
  AOI21_X1  g715(.A(KEYINPUT61), .B1(new_n900), .B2(KEYINPUT125), .ZN(new_n902));
  XNOR2_X1  g716(.A(new_n901), .B(new_n902), .ZN(G66));
  NAND2_X1  g717(.A1(new_n747), .A2(new_n771), .ZN(new_n904));
  NAND2_X1  g718(.A1(new_n904), .A2(new_n187), .ZN(new_n905));
  AOI21_X1  g719(.A(new_n187), .B1(new_n523), .B2(G224), .ZN(new_n906));
  INV_X1    g720(.A(KEYINPUT126), .ZN(new_n907));
  OR2_X1    g721(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  NAND2_X1  g722(.A1(new_n906), .A2(new_n907), .ZN(new_n909));
  NAND3_X1  g723(.A1(new_n905), .A2(new_n908), .A3(new_n909), .ZN(new_n910));
  OAI21_X1  g724(.A(new_n845), .B1(G898), .B2(new_n187), .ZN(new_n911));
  XNOR2_X1  g725(.A(new_n910), .B(new_n911), .ZN(G69));
  NAND2_X1  g726(.A1(new_n753), .A2(new_n613), .ZN(new_n913));
  INV_X1    g727(.A(new_n913), .ZN(new_n914));
  INV_X1    g728(.A(KEYINPUT62), .ZN(new_n915));
  OAI211_X1 g729(.A(new_n630), .B(new_n914), .C1(KEYINPUT127), .C2(new_n915), .ZN(new_n916));
  AND2_X1   g730(.A1(new_n740), .A2(new_n651), .ZN(new_n917));
  NAND4_X1  g731(.A1(new_n637), .A2(new_n617), .A3(new_n672), .A4(new_n917), .ZN(new_n918));
  NAND2_X1  g732(.A1(new_n630), .A2(new_n914), .ZN(new_n919));
  XOR2_X1   g733(.A(KEYINPUT127), .B(KEYINPUT62), .Z(new_n920));
  AOI21_X1  g734(.A(new_n733), .B1(new_n919), .B2(new_n920), .ZN(new_n921));
  NAND4_X1  g735(.A1(new_n724), .A2(new_n916), .A3(new_n918), .A4(new_n921), .ZN(new_n922));
  NAND2_X1  g736(.A1(new_n922), .A2(new_n187), .ZN(new_n923));
  OAI21_X1  g737(.A(new_n326), .B1(new_n331), .B2(new_n325), .ZN(new_n924));
  XNOR2_X1  g738(.A(new_n924), .B(new_n457), .ZN(new_n925));
  NAND2_X1  g739(.A1(new_n923), .A2(new_n925), .ZN(new_n926));
  NOR2_X1   g740(.A1(new_n187), .A2(G900), .ZN(new_n927));
  NOR3_X1   g741(.A1(new_n733), .A2(new_n692), .A3(new_n913), .ZN(new_n928));
  AOI22_X1  g742(.A1(new_n709), .A2(new_n672), .B1(new_n660), .B2(new_n783), .ZN(new_n929));
  OAI211_X1 g743(.A(new_n699), .B(new_n928), .C1(new_n929), .C2(new_n723), .ZN(new_n930));
  AOI21_X1  g744(.A(new_n927), .B1(new_n930), .B2(new_n187), .ZN(new_n931));
  OAI21_X1  g745(.A(new_n926), .B1(new_n931), .B2(new_n925), .ZN(new_n932));
  AOI21_X1  g746(.A(new_n187), .B1(G227), .B2(G900), .ZN(new_n933));
  XNOR2_X1  g747(.A(new_n932), .B(new_n933), .ZN(G72));
  NAND2_X1  g748(.A1(G472), .A2(G902), .ZN(new_n935));
  XOR2_X1   g749(.A(new_n935), .B(KEYINPUT63), .Z(new_n936));
  OAI21_X1  g750(.A(new_n936), .B1(new_n922), .B2(new_n904), .ZN(new_n937));
  AOI21_X1  g751(.A(new_n849), .B1(new_n937), .B2(new_n619), .ZN(new_n938));
  NAND3_X1  g752(.A1(new_n827), .A2(new_n345), .A3(new_n936), .ZN(new_n939));
  OAI21_X1  g753(.A(new_n938), .B1(new_n619), .B2(new_n939), .ZN(new_n940));
  INV_X1    g754(.A(new_n345), .ZN(new_n941));
  OAI21_X1  g755(.A(new_n936), .B1(new_n930), .B2(new_n904), .ZN(new_n942));
  AOI21_X1  g756(.A(new_n940), .B1(new_n941), .B2(new_n942), .ZN(G57));
endmodule


