//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 1 1 0 1 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 0 1 0 0 0 0 1 0 0 1 0 0 1 0 1 1 1 0 1 1 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 0 1 1 0 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:30:06 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n440, new_n448, new_n452, new_n453, new_n454, new_n455,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n538, new_n539, new_n540, new_n541, new_n542,
    new_n543, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n554, new_n556, new_n557, new_n559, new_n560,
    new_n561, new_n562, new_n563, new_n564, new_n565, new_n566, new_n567,
    new_n568, new_n569, new_n570, new_n572, new_n573, new_n575, new_n576,
    new_n577, new_n579, new_n580, new_n581, new_n582, new_n583, new_n584,
    new_n585, new_n586, new_n587, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n609,
    new_n610, new_n613, new_n614, new_n616, new_n617, new_n618, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n835, new_n836,
    new_n837, new_n838, new_n839, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1199, new_n1200, new_n1201, new_n1202,
    new_n1203, new_n1204, new_n1205, new_n1207, new_n1208, new_n1209,
    new_n1210;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  XNOR2_X1  g002(.A(KEYINPUT64), .B(G452), .ZN(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  XNOR2_X1  g005(.A(KEYINPUT65), .B(G2066), .ZN(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  XNOR2_X1  g014(.A(KEYINPUT66), .B(G120), .ZN(new_n440));
  INV_X1    g015(.A(new_n440), .ZN(G236));
  INV_X1    g016(.A(G57), .ZN(G237));
  INV_X1    g017(.A(G108), .ZN(G238));
  NAND4_X1  g018(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g019(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g020(.A(G452), .Z(G391));
  AND2_X1   g021(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XOR2_X1   g023(.A(new_n448), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g024(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g025(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NAND4_X1  g026(.A1(new_n436), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n452));
  XNOR2_X1  g027(.A(new_n452), .B(KEYINPUT2), .ZN(new_n453));
  NAND4_X1  g028(.A1(new_n440), .A2(G57), .A3(G69), .A4(G108), .ZN(new_n454));
  XNOR2_X1  g029(.A(new_n454), .B(KEYINPUT67), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n453), .A2(new_n455), .ZN(G325));
  INV_X1    g031(.A(G325), .ZN(G261));
  AOI22_X1  g032(.A1(new_n453), .A2(G2106), .B1(new_n455), .B2(G567), .ZN(G319));
  XNOR2_X1  g033(.A(KEYINPUT68), .B(G2105), .ZN(new_n459));
  XNOR2_X1  g034(.A(KEYINPUT3), .B(G2104), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n460), .A2(G125), .ZN(new_n461));
  NAND2_X1  g036(.A1(G113), .A2(G2104), .ZN(new_n462));
  AOI21_X1  g037(.A(new_n459), .B1(new_n461), .B2(new_n462), .ZN(new_n463));
  INV_X1    g038(.A(G2104), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n464), .A2(KEYINPUT3), .ZN(new_n465));
  INV_X1    g040(.A(KEYINPUT3), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n466), .A2(G2104), .ZN(new_n467));
  AND2_X1   g042(.A1(KEYINPUT68), .A2(G2105), .ZN(new_n468));
  NOR2_X1   g043(.A1(KEYINPUT68), .A2(G2105), .ZN(new_n469));
  OAI211_X1 g044(.A(new_n465), .B(new_n467), .C1(new_n468), .C2(new_n469), .ZN(new_n470));
  INV_X1    g045(.A(G137), .ZN(new_n471));
  INV_X1    g046(.A(G101), .ZN(new_n472));
  INV_X1    g047(.A(G2105), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n473), .A2(G2104), .ZN(new_n474));
  OAI22_X1  g049(.A1(new_n470), .A2(new_n471), .B1(new_n472), .B2(new_n474), .ZN(new_n475));
  NOR2_X1   g050(.A1(new_n463), .A2(new_n475), .ZN(G160));
  NAND2_X1  g051(.A1(new_n465), .A2(new_n467), .ZN(new_n477));
  NOR2_X1   g052(.A1(new_n477), .A2(G2105), .ZN(new_n478));
  NAND3_X1  g053(.A1(new_n478), .A2(KEYINPUT69), .A3(G136), .ZN(new_n479));
  INV_X1    g054(.A(KEYINPUT69), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n460), .A2(new_n473), .ZN(new_n481));
  INV_X1    g056(.A(G136), .ZN(new_n482));
  OAI21_X1  g057(.A(new_n480), .B1(new_n481), .B2(new_n482), .ZN(new_n483));
  NOR2_X1   g058(.A1(new_n477), .A2(new_n459), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n484), .A2(G124), .ZN(new_n485));
  OAI221_X1 g060(.A(G2104), .B1(G100), .B2(G2105), .C1(new_n459), .C2(G112), .ZN(new_n486));
  NAND4_X1  g061(.A1(new_n479), .A2(new_n483), .A3(new_n485), .A4(new_n486), .ZN(new_n487));
  INV_X1    g062(.A(new_n487), .ZN(G162));
  INV_X1    g063(.A(KEYINPUT4), .ZN(new_n489));
  INV_X1    g064(.A(G138), .ZN(new_n490));
  OAI21_X1  g065(.A(new_n489), .B1(new_n470), .B2(new_n490), .ZN(new_n491));
  INV_X1    g066(.A(KEYINPUT70), .ZN(new_n492));
  OAI21_X1  g067(.A(G2104), .B1(new_n473), .B2(G114), .ZN(new_n493));
  NOR2_X1   g068(.A1(G102), .A2(G2105), .ZN(new_n494));
  OAI21_X1  g069(.A(new_n492), .B1(new_n493), .B2(new_n494), .ZN(new_n495));
  OR2_X1    g070(.A1(G102), .A2(G2105), .ZN(new_n496));
  INV_X1    g071(.A(G114), .ZN(new_n497));
  NAND2_X1  g072(.A1(new_n497), .A2(G2105), .ZN(new_n498));
  NAND4_X1  g073(.A1(new_n496), .A2(new_n498), .A3(KEYINPUT70), .A4(G2104), .ZN(new_n499));
  NAND2_X1  g074(.A1(new_n495), .A2(new_n499), .ZN(new_n500));
  NAND3_X1  g075(.A1(new_n460), .A2(G126), .A3(G2105), .ZN(new_n501));
  NAND4_X1  g076(.A1(new_n459), .A2(new_n460), .A3(KEYINPUT4), .A4(G138), .ZN(new_n502));
  NAND4_X1  g077(.A1(new_n491), .A2(new_n500), .A3(new_n501), .A4(new_n502), .ZN(new_n503));
  INV_X1    g078(.A(new_n503), .ZN(G164));
  NAND2_X1  g079(.A1(G75), .A2(G543), .ZN(new_n505));
  INV_X1    g080(.A(G543), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n506), .A2(KEYINPUT5), .ZN(new_n507));
  INV_X1    g082(.A(KEYINPUT5), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n508), .A2(G543), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n507), .A2(new_n509), .ZN(new_n510));
  INV_X1    g085(.A(G62), .ZN(new_n511));
  OAI21_X1  g086(.A(new_n505), .B1(new_n510), .B2(new_n511), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n512), .A2(G651), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n513), .A2(KEYINPUT72), .ZN(new_n514));
  XNOR2_X1  g089(.A(KEYINPUT6), .B(G651), .ZN(new_n515));
  AND2_X1   g090(.A1(new_n515), .A2(G543), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n516), .A2(G50), .ZN(new_n517));
  AND2_X1   g092(.A1(KEYINPUT6), .A2(G651), .ZN(new_n518));
  NOR2_X1   g093(.A1(KEYINPUT6), .A2(G651), .ZN(new_n519));
  OAI211_X1 g094(.A(new_n507), .B(new_n509), .C1(new_n518), .C2(new_n519), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n520), .A2(KEYINPUT71), .ZN(new_n521));
  XNOR2_X1  g096(.A(KEYINPUT5), .B(G543), .ZN(new_n522));
  INV_X1    g097(.A(KEYINPUT71), .ZN(new_n523));
  NAND3_X1  g098(.A1(new_n515), .A2(new_n522), .A3(new_n523), .ZN(new_n524));
  NAND3_X1  g099(.A1(new_n521), .A2(G88), .A3(new_n524), .ZN(new_n525));
  INV_X1    g100(.A(KEYINPUT72), .ZN(new_n526));
  NAND3_X1  g101(.A1(new_n512), .A2(new_n526), .A3(G651), .ZN(new_n527));
  NAND4_X1  g102(.A1(new_n514), .A2(new_n517), .A3(new_n525), .A4(new_n527), .ZN(G303));
  INV_X1    g103(.A(G303), .ZN(G166));
  NAND3_X1  g104(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n530));
  XNOR2_X1  g105(.A(new_n530), .B(KEYINPUT7), .ZN(new_n531));
  NAND3_X1  g106(.A1(new_n522), .A2(G63), .A3(G651), .ZN(new_n532));
  NAND3_X1  g107(.A1(new_n515), .A2(G51), .A3(G543), .ZN(new_n533));
  AND3_X1   g108(.A1(new_n531), .A2(new_n532), .A3(new_n533), .ZN(new_n534));
  NAND3_X1  g109(.A1(new_n521), .A2(G89), .A3(new_n524), .ZN(new_n535));
  NAND2_X1  g110(.A1(new_n534), .A2(new_n535), .ZN(G286));
  INV_X1    g111(.A(G286), .ZN(G168));
  AOI22_X1  g112(.A1(new_n522), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n538));
  INV_X1    g113(.A(G651), .ZN(new_n539));
  INV_X1    g114(.A(G52), .ZN(new_n540));
  NAND2_X1  g115(.A1(new_n515), .A2(G543), .ZN(new_n541));
  OAI22_X1  g116(.A1(new_n538), .A2(new_n539), .B1(new_n540), .B2(new_n541), .ZN(new_n542));
  AND2_X1   g117(.A1(new_n521), .A2(new_n524), .ZN(new_n543));
  AOI21_X1  g118(.A(new_n542), .B1(G90), .B2(new_n543), .ZN(G171));
  AOI22_X1  g119(.A1(new_n522), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n545));
  OR2_X1    g120(.A1(new_n545), .A2(new_n539), .ZN(new_n546));
  NAND3_X1  g121(.A1(new_n521), .A2(G81), .A3(new_n524), .ZN(new_n547));
  NAND2_X1  g122(.A1(new_n516), .A2(G43), .ZN(new_n548));
  AND3_X1   g123(.A1(new_n547), .A2(KEYINPUT73), .A3(new_n548), .ZN(new_n549));
  AOI21_X1  g124(.A(KEYINPUT73), .B1(new_n547), .B2(new_n548), .ZN(new_n550));
  OAI21_X1  g125(.A(new_n546), .B1(new_n549), .B2(new_n550), .ZN(new_n551));
  INV_X1    g126(.A(new_n551), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n552), .A2(G860), .ZN(G153));
  AND3_X1   g128(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n554), .A2(G36), .ZN(G176));
  NAND2_X1  g130(.A1(G1), .A2(G3), .ZN(new_n556));
  XNOR2_X1  g131(.A(new_n556), .B(KEYINPUT8), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n554), .A2(new_n557), .ZN(G188));
  NAND2_X1  g133(.A1(new_n521), .A2(new_n524), .ZN(new_n559));
  INV_X1    g134(.A(G91), .ZN(new_n560));
  OAI21_X1  g135(.A(KEYINPUT74), .B1(new_n559), .B2(new_n560), .ZN(new_n561));
  INV_X1    g136(.A(KEYINPUT74), .ZN(new_n562));
  NAND4_X1  g137(.A1(new_n521), .A2(new_n524), .A3(new_n562), .A4(G91), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n561), .A2(new_n563), .ZN(new_n564));
  NAND2_X1  g139(.A1(new_n516), .A2(G53), .ZN(new_n565));
  XNOR2_X1  g140(.A(new_n565), .B(KEYINPUT9), .ZN(new_n566));
  NAND2_X1  g141(.A1(G78), .A2(G543), .ZN(new_n567));
  INV_X1    g142(.A(G65), .ZN(new_n568));
  OAI21_X1  g143(.A(new_n567), .B1(new_n510), .B2(new_n568), .ZN(new_n569));
  NAND2_X1  g144(.A1(new_n569), .A2(G651), .ZN(new_n570));
  NAND3_X1  g145(.A1(new_n564), .A2(new_n566), .A3(new_n570), .ZN(G299));
  NAND2_X1  g146(.A1(new_n516), .A2(G52), .ZN(new_n572));
  INV_X1    g147(.A(G90), .ZN(new_n573));
  OAI221_X1 g148(.A(new_n572), .B1(new_n539), .B2(new_n538), .C1(new_n559), .C2(new_n573), .ZN(G301));
  OAI21_X1  g149(.A(G651), .B1(new_n522), .B2(G74), .ZN(new_n575));
  NAND2_X1  g150(.A1(new_n516), .A2(G49), .ZN(new_n576));
  INV_X1    g151(.A(G87), .ZN(new_n577));
  OAI211_X1 g152(.A(new_n575), .B(new_n576), .C1(new_n559), .C2(new_n577), .ZN(G288));
  INV_X1    g153(.A(KEYINPUT75), .ZN(new_n579));
  AOI22_X1  g154(.A1(new_n522), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n580));
  OAI21_X1  g155(.A(new_n579), .B1(new_n580), .B2(new_n539), .ZN(new_n581));
  NAND3_X1  g156(.A1(new_n521), .A2(G86), .A3(new_n524), .ZN(new_n582));
  NAND2_X1  g157(.A1(new_n516), .A2(G48), .ZN(new_n583));
  NAND3_X1  g158(.A1(new_n507), .A2(new_n509), .A3(G61), .ZN(new_n584));
  NAND2_X1  g159(.A1(G73), .A2(G543), .ZN(new_n585));
  NAND2_X1  g160(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  NAND3_X1  g161(.A1(new_n586), .A2(KEYINPUT75), .A3(G651), .ZN(new_n587));
  NAND4_X1  g162(.A1(new_n581), .A2(new_n582), .A3(new_n583), .A4(new_n587), .ZN(G305));
  NAND2_X1  g163(.A1(new_n516), .A2(G47), .ZN(new_n589));
  INV_X1    g164(.A(G85), .ZN(new_n590));
  OAI21_X1  g165(.A(new_n589), .B1(new_n559), .B2(new_n590), .ZN(new_n591));
  XNOR2_X1  g166(.A(new_n591), .B(KEYINPUT76), .ZN(new_n592));
  AOI22_X1  g167(.A1(new_n522), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n593));
  OR2_X1    g168(.A1(new_n593), .A2(new_n539), .ZN(new_n594));
  NAND2_X1  g169(.A1(new_n592), .A2(new_n594), .ZN(G290));
  NAND2_X1  g170(.A1(G301), .A2(G868), .ZN(new_n596));
  XNOR2_X1  g171(.A(new_n541), .B(KEYINPUT77), .ZN(new_n597));
  NAND2_X1  g172(.A1(G79), .A2(G543), .ZN(new_n598));
  INV_X1    g173(.A(G66), .ZN(new_n599));
  OAI21_X1  g174(.A(new_n598), .B1(new_n510), .B2(new_n599), .ZN(new_n600));
  AOI22_X1  g175(.A1(new_n597), .A2(G54), .B1(G651), .B2(new_n600), .ZN(new_n601));
  INV_X1    g176(.A(G92), .ZN(new_n602));
  OR3_X1    g177(.A1(new_n559), .A2(KEYINPUT10), .A3(new_n602), .ZN(new_n603));
  OAI21_X1  g178(.A(KEYINPUT10), .B1(new_n559), .B2(new_n602), .ZN(new_n604));
  NAND3_X1  g179(.A1(new_n601), .A2(new_n603), .A3(new_n604), .ZN(new_n605));
  INV_X1    g180(.A(new_n605), .ZN(new_n606));
  OAI21_X1  g181(.A(new_n596), .B1(new_n606), .B2(G868), .ZN(G284));
  OAI21_X1  g182(.A(new_n596), .B1(new_n606), .B2(G868), .ZN(G321));
  NAND2_X1  g183(.A1(G286), .A2(G868), .ZN(new_n609));
  INV_X1    g184(.A(G299), .ZN(new_n610));
  OAI21_X1  g185(.A(new_n609), .B1(new_n610), .B2(G868), .ZN(G297));
  OAI21_X1  g186(.A(new_n609), .B1(new_n610), .B2(G868), .ZN(G280));
  XNOR2_X1  g187(.A(KEYINPUT78), .B(G559), .ZN(new_n613));
  INV_X1    g188(.A(new_n613), .ZN(new_n614));
  OAI21_X1  g189(.A(new_n606), .B1(G860), .B2(new_n614), .ZN(G148));
  INV_X1    g190(.A(G868), .ZN(new_n616));
  NAND2_X1  g191(.A1(new_n551), .A2(new_n616), .ZN(new_n617));
  NOR2_X1   g192(.A1(new_n605), .A2(new_n613), .ZN(new_n618));
  OAI21_X1  g193(.A(new_n617), .B1(new_n618), .B2(new_n616), .ZN(G323));
  XNOR2_X1  g194(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g195(.A1(new_n484), .A2(G123), .ZN(new_n621));
  NAND2_X1  g196(.A1(new_n478), .A2(G135), .ZN(new_n622));
  OAI221_X1 g197(.A(G2104), .B1(G99), .B2(G2105), .C1(new_n459), .C2(G111), .ZN(new_n623));
  NAND3_X1  g198(.A1(new_n621), .A2(new_n622), .A3(new_n623), .ZN(new_n624));
  XOR2_X1   g199(.A(new_n624), .B(G2096), .Z(new_n625));
  NAND2_X1  g200(.A1(KEYINPUT80), .A2(G2100), .ZN(new_n626));
  NOR2_X1   g201(.A1(new_n477), .A2(new_n474), .ZN(new_n627));
  XOR2_X1   g202(.A(KEYINPUT79), .B(KEYINPUT12), .Z(new_n628));
  XNOR2_X1  g203(.A(new_n627), .B(new_n628), .ZN(new_n629));
  NOR2_X1   g204(.A1(KEYINPUT80), .A2(G2100), .ZN(new_n630));
  XOR2_X1   g205(.A(new_n630), .B(KEYINPUT13), .Z(new_n631));
  XNOR2_X1  g206(.A(new_n629), .B(new_n631), .ZN(new_n632));
  NAND3_X1  g207(.A1(new_n625), .A2(new_n626), .A3(new_n632), .ZN(G156));
  XNOR2_X1  g208(.A(G2443), .B(G2446), .ZN(new_n634));
  INV_X1    g209(.A(new_n634), .ZN(new_n635));
  XNOR2_X1  g210(.A(KEYINPUT15), .B(G2430), .ZN(new_n636));
  XNOR2_X1  g211(.A(new_n636), .B(G2435), .ZN(new_n637));
  XOR2_X1   g212(.A(G2427), .B(G2438), .Z(new_n638));
  XNOR2_X1  g213(.A(new_n637), .B(new_n638), .ZN(new_n639));
  NAND2_X1  g214(.A1(new_n639), .A2(KEYINPUT14), .ZN(new_n640));
  XNOR2_X1  g215(.A(G2451), .B(G2454), .ZN(new_n641));
  XOR2_X1   g216(.A(new_n641), .B(KEYINPUT16), .Z(new_n642));
  NAND2_X1  g217(.A1(new_n640), .A2(new_n642), .ZN(new_n643));
  XNOR2_X1  g218(.A(G1341), .B(G1348), .ZN(new_n644));
  INV_X1    g219(.A(new_n644), .ZN(new_n645));
  INV_X1    g220(.A(new_n642), .ZN(new_n646));
  NAND3_X1  g221(.A1(new_n639), .A2(KEYINPUT14), .A3(new_n646), .ZN(new_n647));
  NAND3_X1  g222(.A1(new_n643), .A2(new_n645), .A3(new_n647), .ZN(new_n648));
  INV_X1    g223(.A(new_n648), .ZN(new_n649));
  AOI21_X1  g224(.A(new_n645), .B1(new_n643), .B2(new_n647), .ZN(new_n650));
  OAI21_X1  g225(.A(new_n635), .B1(new_n649), .B2(new_n650), .ZN(new_n651));
  INV_X1    g226(.A(new_n650), .ZN(new_n652));
  NAND3_X1  g227(.A1(new_n652), .A2(new_n634), .A3(new_n648), .ZN(new_n653));
  NAND3_X1  g228(.A1(new_n651), .A2(new_n653), .A3(G14), .ZN(new_n654));
  INV_X1    g229(.A(KEYINPUT81), .ZN(new_n655));
  XNOR2_X1  g230(.A(new_n654), .B(new_n655), .ZN(new_n656));
  INV_X1    g231(.A(new_n656), .ZN(G401));
  XNOR2_X1  g232(.A(G2072), .B(G2078), .ZN(new_n658));
  XOR2_X1   g233(.A(new_n658), .B(KEYINPUT17), .Z(new_n659));
  XNOR2_X1  g234(.A(G2084), .B(G2090), .ZN(new_n660));
  INV_X1    g235(.A(new_n660), .ZN(new_n661));
  XNOR2_X1  g236(.A(G2067), .B(G2678), .ZN(new_n662));
  INV_X1    g237(.A(new_n662), .ZN(new_n663));
  NAND3_X1  g238(.A1(new_n659), .A2(new_n661), .A3(new_n663), .ZN(new_n664));
  XNOR2_X1  g239(.A(new_n664), .B(KEYINPUT82), .ZN(new_n665));
  NAND3_X1  g240(.A1(new_n661), .A2(new_n658), .A3(new_n662), .ZN(new_n666));
  XOR2_X1   g241(.A(new_n666), .B(KEYINPUT18), .Z(new_n667));
  NOR2_X1   g242(.A1(new_n658), .A2(new_n662), .ZN(new_n668));
  OAI21_X1  g243(.A(new_n660), .B1(new_n659), .B2(new_n663), .ZN(new_n669));
  OAI211_X1 g244(.A(new_n665), .B(new_n667), .C1(new_n668), .C2(new_n669), .ZN(new_n670));
  XNOR2_X1  g245(.A(new_n670), .B(G2096), .ZN(new_n671));
  XNOR2_X1  g246(.A(new_n671), .B(G2100), .ZN(new_n672));
  INV_X1    g247(.A(new_n672), .ZN(G227));
  XNOR2_X1  g248(.A(G1971), .B(G1976), .ZN(new_n674));
  XNOR2_X1  g249(.A(new_n674), .B(KEYINPUT19), .ZN(new_n675));
  INV_X1    g250(.A(new_n675), .ZN(new_n676));
  XOR2_X1   g251(.A(G1956), .B(G2474), .Z(new_n677));
  XNOR2_X1  g252(.A(new_n677), .B(KEYINPUT83), .ZN(new_n678));
  XNOR2_X1  g253(.A(G1961), .B(G1966), .ZN(new_n679));
  XNOR2_X1  g254(.A(new_n679), .B(KEYINPUT84), .ZN(new_n680));
  NAND3_X1  g255(.A1(new_n676), .A2(new_n678), .A3(new_n680), .ZN(new_n681));
  INV_X1    g256(.A(KEYINPUT20), .ZN(new_n682));
  NOR2_X1   g257(.A1(new_n678), .A2(new_n680), .ZN(new_n683));
  AOI22_X1  g258(.A1(new_n681), .A2(new_n682), .B1(new_n683), .B2(new_n676), .ZN(new_n684));
  INV_X1    g259(.A(new_n683), .ZN(new_n685));
  NAND2_X1  g260(.A1(new_n678), .A2(new_n680), .ZN(new_n686));
  NAND3_X1  g261(.A1(new_n685), .A2(new_n675), .A3(new_n686), .ZN(new_n687));
  OAI211_X1 g262(.A(new_n684), .B(new_n687), .C1(new_n682), .C2(new_n681), .ZN(new_n688));
  XNOR2_X1  g263(.A(G1991), .B(G1996), .ZN(new_n689));
  XNOR2_X1  g264(.A(new_n689), .B(G1981), .ZN(new_n690));
  XNOR2_X1  g265(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n691));
  XNOR2_X1  g266(.A(new_n690), .B(new_n691), .ZN(new_n692));
  XNOR2_X1  g267(.A(new_n688), .B(new_n692), .ZN(new_n693));
  XNOR2_X1  g268(.A(KEYINPUT85), .B(G1986), .ZN(new_n694));
  XNOR2_X1  g269(.A(new_n693), .B(new_n694), .ZN(new_n695));
  INV_X1    g270(.A(new_n695), .ZN(G229));
  NAND2_X1  g271(.A1(new_n484), .A2(G128), .ZN(new_n697));
  NAND2_X1  g272(.A1(new_n478), .A2(G140), .ZN(new_n698));
  OAI221_X1 g273(.A(G2104), .B1(G104), .B2(G2105), .C1(new_n459), .C2(G116), .ZN(new_n699));
  NAND3_X1  g274(.A1(new_n697), .A2(new_n698), .A3(new_n699), .ZN(new_n700));
  INV_X1    g275(.A(KEYINPUT89), .ZN(new_n701));
  NAND2_X1  g276(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  NAND4_X1  g277(.A1(new_n697), .A2(new_n698), .A3(new_n699), .A4(KEYINPUT89), .ZN(new_n703));
  AND2_X1   g278(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  INV_X1    g279(.A(G29), .ZN(new_n705));
  NOR2_X1   g280(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  AND2_X1   g281(.A1(new_n705), .A2(G26), .ZN(new_n707));
  OAI21_X1  g282(.A(KEYINPUT28), .B1(new_n706), .B2(new_n707), .ZN(new_n708));
  INV_X1    g283(.A(G2067), .ZN(new_n709));
  OR2_X1    g284(.A1(new_n707), .A2(KEYINPUT28), .ZN(new_n710));
  AND3_X1   g285(.A1(new_n708), .A2(new_n709), .A3(new_n710), .ZN(new_n711));
  NAND2_X1  g286(.A1(new_n606), .A2(G16), .ZN(new_n712));
  OAI21_X1  g287(.A(new_n712), .B1(G4), .B2(G16), .ZN(new_n713));
  INV_X1    g288(.A(G1348), .ZN(new_n714));
  NOR2_X1   g289(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  AOI21_X1  g290(.A(new_n709), .B1(new_n708), .B2(new_n710), .ZN(new_n716));
  NOR3_X1   g291(.A1(new_n711), .A2(new_n715), .A3(new_n716), .ZN(new_n717));
  INV_X1    g292(.A(G16), .ZN(new_n718));
  NAND3_X1  g293(.A1(new_n718), .A2(KEYINPUT23), .A3(G20), .ZN(new_n719));
  INV_X1    g294(.A(KEYINPUT23), .ZN(new_n720));
  INV_X1    g295(.A(G20), .ZN(new_n721));
  OAI21_X1  g296(.A(new_n720), .B1(new_n721), .B2(G16), .ZN(new_n722));
  OAI211_X1 g297(.A(new_n719), .B(new_n722), .C1(new_n610), .C2(new_n718), .ZN(new_n723));
  XNOR2_X1  g298(.A(new_n723), .B(G1956), .ZN(new_n724));
  NAND2_X1  g299(.A1(G171), .A2(G16), .ZN(new_n725));
  OAI21_X1  g300(.A(new_n725), .B1(G5), .B2(G16), .ZN(new_n726));
  INV_X1    g301(.A(G1961), .ZN(new_n727));
  OR2_X1    g302(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  NAND2_X1  g303(.A1(new_n726), .A2(new_n727), .ZN(new_n729));
  INV_X1    g304(.A(G2072), .ZN(new_n730));
  NAND3_X1  g305(.A1(new_n459), .A2(G103), .A3(G2104), .ZN(new_n731));
  XNOR2_X1  g306(.A(new_n731), .B(KEYINPUT25), .ZN(new_n732));
  AOI22_X1  g307(.A1(new_n460), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n733));
  NOR2_X1   g308(.A1(new_n733), .A2(new_n459), .ZN(new_n734));
  AND2_X1   g309(.A1(new_n478), .A2(G139), .ZN(new_n735));
  NOR3_X1   g310(.A1(new_n732), .A2(new_n734), .A3(new_n735), .ZN(new_n736));
  NAND2_X1  g311(.A1(new_n736), .A2(G29), .ZN(new_n737));
  OAI21_X1  g312(.A(new_n737), .B1(G29), .B2(G33), .ZN(new_n738));
  OAI211_X1 g313(.A(new_n728), .B(new_n729), .C1(new_n730), .C2(new_n738), .ZN(new_n739));
  NOR2_X1   g314(.A1(new_n724), .A2(new_n739), .ZN(new_n740));
  NAND2_X1  g315(.A1(new_n705), .A2(G35), .ZN(new_n741));
  OAI21_X1  g316(.A(new_n741), .B1(G162), .B2(new_n705), .ZN(new_n742));
  INV_X1    g317(.A(KEYINPUT93), .ZN(new_n743));
  XNOR2_X1  g318(.A(new_n742), .B(new_n743), .ZN(new_n744));
  AND2_X1   g319(.A1(new_n744), .A2(KEYINPUT29), .ZN(new_n745));
  NOR2_X1   g320(.A1(new_n744), .A2(KEYINPUT29), .ZN(new_n746));
  OR3_X1    g321(.A1(new_n745), .A2(new_n746), .A3(G2090), .ZN(new_n747));
  OAI21_X1  g322(.A(G2090), .B1(new_n745), .B2(new_n746), .ZN(new_n748));
  NAND4_X1  g323(.A1(new_n717), .A2(new_n740), .A3(new_n747), .A4(new_n748), .ZN(new_n749));
  AOI22_X1  g324(.A1(G129), .A2(new_n484), .B1(new_n478), .B2(G141), .ZN(new_n750));
  NAND3_X1  g325(.A1(new_n473), .A2(G105), .A3(G2104), .ZN(new_n751));
  NAND3_X1  g326(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n752));
  XOR2_X1   g327(.A(new_n752), .B(KEYINPUT26), .Z(new_n753));
  NAND3_X1  g328(.A1(new_n750), .A2(new_n751), .A3(new_n753), .ZN(new_n754));
  XOR2_X1   g329(.A(new_n754), .B(KEYINPUT90), .Z(new_n755));
  NAND2_X1  g330(.A1(new_n755), .A2(G29), .ZN(new_n756));
  XNOR2_X1  g331(.A(KEYINPUT27), .B(G1996), .ZN(new_n757));
  NAND2_X1  g332(.A1(new_n705), .A2(G32), .ZN(new_n758));
  AND3_X1   g333(.A1(new_n756), .A2(new_n757), .A3(new_n758), .ZN(new_n759));
  AOI21_X1  g334(.A(new_n757), .B1(new_n756), .B2(new_n758), .ZN(new_n760));
  XNOR2_X1  g335(.A(KEYINPUT92), .B(G28), .ZN(new_n761));
  XNOR2_X1  g336(.A(new_n761), .B(KEYINPUT30), .ZN(new_n762));
  NOR2_X1   g337(.A1(new_n762), .A2(G29), .ZN(new_n763));
  NOR3_X1   g338(.A1(new_n759), .A2(new_n760), .A3(new_n763), .ZN(new_n764));
  INV_X1    g339(.A(G34), .ZN(new_n765));
  AND2_X1   g340(.A1(new_n765), .A2(KEYINPUT24), .ZN(new_n766));
  NOR2_X1   g341(.A1(new_n765), .A2(KEYINPUT24), .ZN(new_n767));
  OAI21_X1  g342(.A(new_n705), .B1(new_n766), .B2(new_n767), .ZN(new_n768));
  OAI21_X1  g343(.A(new_n768), .B1(G160), .B2(new_n705), .ZN(new_n769));
  INV_X1    g344(.A(G2084), .ZN(new_n770));
  XNOR2_X1  g345(.A(new_n769), .B(new_n770), .ZN(new_n771));
  NAND2_X1  g346(.A1(new_n552), .A2(G16), .ZN(new_n772));
  OAI21_X1  g347(.A(new_n772), .B1(G16), .B2(G19), .ZN(new_n773));
  INV_X1    g348(.A(G1341), .ZN(new_n774));
  NAND2_X1  g349(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  OR2_X1    g350(.A1(new_n624), .A2(new_n705), .ZN(new_n776));
  NAND4_X1  g351(.A1(new_n764), .A2(new_n771), .A3(new_n775), .A4(new_n776), .ZN(new_n777));
  NAND2_X1  g352(.A1(new_n713), .A2(new_n714), .ZN(new_n778));
  INV_X1    g353(.A(new_n778), .ZN(new_n779));
  NOR2_X1   g354(.A1(new_n773), .A2(new_n774), .ZN(new_n780));
  NOR4_X1   g355(.A1(new_n749), .A2(new_n777), .A3(new_n779), .A4(new_n780), .ZN(new_n781));
  XNOR2_X1  g356(.A(KEYINPUT31), .B(G11), .ZN(new_n782));
  XNOR2_X1  g357(.A(new_n782), .B(KEYINPUT91), .ZN(new_n783));
  NAND2_X1  g358(.A1(new_n718), .A2(G22), .ZN(new_n784));
  OAI21_X1  g359(.A(new_n784), .B1(G166), .B2(new_n718), .ZN(new_n785));
  INV_X1    g360(.A(G1971), .ZN(new_n786));
  XNOR2_X1  g361(.A(new_n785), .B(new_n786), .ZN(new_n787));
  MUX2_X1   g362(.A(G23), .B(G288), .S(G16), .Z(new_n788));
  XNOR2_X1  g363(.A(KEYINPUT33), .B(G1976), .ZN(new_n789));
  XNOR2_X1  g364(.A(new_n788), .B(new_n789), .ZN(new_n790));
  NAND2_X1  g365(.A1(new_n787), .A2(new_n790), .ZN(new_n791));
  NAND2_X1  g366(.A1(new_n718), .A2(G6), .ZN(new_n792));
  INV_X1    g367(.A(G305), .ZN(new_n793));
  OAI21_X1  g368(.A(new_n792), .B1(new_n793), .B2(new_n718), .ZN(new_n794));
  XOR2_X1   g369(.A(KEYINPUT32), .B(G1981), .Z(new_n795));
  XOR2_X1   g370(.A(new_n794), .B(new_n795), .Z(new_n796));
  NOR2_X1   g371(.A1(new_n791), .A2(new_n796), .ZN(new_n797));
  INV_X1    g372(.A(KEYINPUT88), .ZN(new_n798));
  NAND3_X1  g373(.A1(new_n797), .A2(new_n798), .A3(KEYINPUT34), .ZN(new_n799));
  OR2_X1    g374(.A1(new_n798), .A2(KEYINPUT34), .ZN(new_n800));
  NAND2_X1  g375(.A1(new_n798), .A2(KEYINPUT34), .ZN(new_n801));
  OAI211_X1 g376(.A(new_n800), .B(new_n801), .C1(new_n791), .C2(new_n796), .ZN(new_n802));
  NAND2_X1  g377(.A1(new_n799), .A2(new_n802), .ZN(new_n803));
  NAND2_X1  g378(.A1(new_n484), .A2(G119), .ZN(new_n804));
  NAND2_X1  g379(.A1(new_n478), .A2(G131), .ZN(new_n805));
  OAI221_X1 g380(.A(G2104), .B1(G95), .B2(G2105), .C1(new_n459), .C2(G107), .ZN(new_n806));
  NAND3_X1  g381(.A1(new_n804), .A2(new_n805), .A3(new_n806), .ZN(new_n807));
  MUX2_X1   g382(.A(G25), .B(new_n807), .S(G29), .Z(new_n808));
  XNOR2_X1  g383(.A(KEYINPUT35), .B(G1991), .ZN(new_n809));
  XNOR2_X1  g384(.A(new_n808), .B(new_n809), .ZN(new_n810));
  NOR2_X1   g385(.A1(G16), .A2(G24), .ZN(new_n811));
  INV_X1    g386(.A(new_n811), .ZN(new_n812));
  XNOR2_X1  g387(.A(G290), .B(KEYINPUT86), .ZN(new_n813));
  OAI21_X1  g388(.A(new_n812), .B1(new_n813), .B2(new_n718), .ZN(new_n814));
  XOR2_X1   g389(.A(KEYINPUT87), .B(G1986), .Z(new_n815));
  NAND2_X1  g390(.A1(new_n814), .A2(new_n815), .ZN(new_n816));
  INV_X1    g391(.A(new_n815), .ZN(new_n817));
  OAI211_X1 g392(.A(new_n817), .B(new_n812), .C1(new_n813), .C2(new_n718), .ZN(new_n818));
  AOI21_X1  g393(.A(new_n810), .B1(new_n816), .B2(new_n818), .ZN(new_n819));
  INV_X1    g394(.A(KEYINPUT36), .ZN(new_n820));
  AND3_X1   g395(.A1(new_n803), .A2(new_n819), .A3(new_n820), .ZN(new_n821));
  AOI21_X1  g396(.A(new_n820), .B1(new_n803), .B2(new_n819), .ZN(new_n822));
  OAI211_X1 g397(.A(new_n781), .B(new_n783), .C1(new_n821), .C2(new_n822), .ZN(new_n823));
  NAND2_X1  g398(.A1(new_n718), .A2(G21), .ZN(new_n824));
  OAI21_X1  g399(.A(new_n824), .B1(G168), .B2(new_n718), .ZN(new_n825));
  XNOR2_X1  g400(.A(new_n825), .B(G1966), .ZN(new_n826));
  NAND2_X1  g401(.A1(new_n705), .A2(G27), .ZN(new_n827));
  OAI21_X1  g402(.A(new_n827), .B1(G164), .B2(new_n705), .ZN(new_n828));
  INV_X1    g403(.A(G2078), .ZN(new_n829));
  XNOR2_X1  g404(.A(new_n828), .B(new_n829), .ZN(new_n830));
  INV_X1    g405(.A(new_n830), .ZN(new_n831));
  NAND2_X1  g406(.A1(new_n738), .A2(new_n730), .ZN(new_n832));
  INV_X1    g407(.A(new_n832), .ZN(new_n833));
  NOR4_X1   g408(.A1(new_n823), .A2(new_n826), .A3(new_n831), .A4(new_n833), .ZN(G311));
  NOR3_X1   g409(.A1(new_n749), .A2(new_n780), .A3(new_n777), .ZN(new_n835));
  NAND3_X1  g410(.A1(new_n835), .A2(new_n783), .A3(new_n778), .ZN(new_n836));
  NOR2_X1   g411(.A1(new_n821), .A2(new_n822), .ZN(new_n837));
  NOR2_X1   g412(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  INV_X1    g413(.A(new_n826), .ZN(new_n839));
  NAND4_X1  g414(.A1(new_n838), .A2(new_n839), .A3(new_n830), .A4(new_n832), .ZN(G150));
  NAND2_X1  g415(.A1(new_n543), .A2(G93), .ZN(new_n841));
  NAND2_X1  g416(.A1(G80), .A2(G543), .ZN(new_n842));
  INV_X1    g417(.A(G67), .ZN(new_n843));
  OAI21_X1  g418(.A(new_n842), .B1(new_n510), .B2(new_n843), .ZN(new_n844));
  AOI22_X1  g419(.A1(new_n844), .A2(G651), .B1(new_n516), .B2(G55), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n841), .A2(new_n845), .ZN(new_n846));
  NAND2_X1  g421(.A1(new_n846), .A2(G860), .ZN(new_n847));
  XOR2_X1   g422(.A(KEYINPUT94), .B(KEYINPUT37), .Z(new_n848));
  XNOR2_X1  g423(.A(new_n847), .B(new_n848), .ZN(new_n849));
  NAND3_X1  g424(.A1(new_n551), .A2(new_n841), .A3(new_n845), .ZN(new_n850));
  OAI211_X1 g425(.A(new_n846), .B(new_n546), .C1(new_n549), .C2(new_n550), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  XNOR2_X1  g427(.A(KEYINPUT38), .B(KEYINPUT39), .ZN(new_n853));
  XNOR2_X1  g428(.A(new_n852), .B(new_n853), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n606), .A2(G559), .ZN(new_n855));
  XNOR2_X1  g430(.A(new_n854), .B(new_n855), .ZN(new_n856));
  OAI21_X1  g431(.A(new_n849), .B1(new_n856), .B2(G860), .ZN(G145));
  INV_X1    g432(.A(G37), .ZN(new_n858));
  INV_X1    g433(.A(new_n755), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n702), .A2(new_n703), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n860), .A2(new_n503), .ZN(new_n861));
  INV_X1    g436(.A(KEYINPUT95), .ZN(new_n862));
  NAND3_X1  g437(.A1(new_n702), .A2(G164), .A3(new_n703), .ZN(new_n863));
  AND3_X1   g438(.A1(new_n861), .A2(new_n862), .A3(new_n863), .ZN(new_n864));
  AOI21_X1  g439(.A(new_n862), .B1(new_n861), .B2(new_n863), .ZN(new_n865));
  OAI21_X1  g440(.A(new_n859), .B1(new_n864), .B2(new_n865), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n861), .A2(new_n863), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n867), .A2(KEYINPUT95), .ZN(new_n868));
  NAND3_X1  g443(.A1(new_n861), .A2(new_n862), .A3(new_n863), .ZN(new_n869));
  NAND3_X1  g444(.A1(new_n868), .A2(new_n755), .A3(new_n869), .ZN(new_n870));
  NAND3_X1  g445(.A1(new_n866), .A2(new_n870), .A3(new_n736), .ZN(new_n871));
  INV_X1    g446(.A(new_n736), .ZN(new_n872));
  INV_X1    g447(.A(new_n754), .ZN(new_n873));
  AND3_X1   g448(.A1(new_n861), .A2(new_n873), .A3(new_n863), .ZN(new_n874));
  AOI21_X1  g449(.A(new_n873), .B1(new_n861), .B2(new_n863), .ZN(new_n875));
  OAI21_X1  g450(.A(new_n872), .B1(new_n874), .B2(new_n875), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n876), .A2(KEYINPUT96), .ZN(new_n877));
  INV_X1    g452(.A(KEYINPUT96), .ZN(new_n878));
  OAI211_X1 g453(.A(new_n878), .B(new_n872), .C1(new_n874), .C2(new_n875), .ZN(new_n879));
  NAND3_X1  g454(.A1(new_n871), .A2(new_n877), .A3(new_n879), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n484), .A2(G130), .ZN(new_n881));
  XNOR2_X1  g456(.A(new_n881), .B(KEYINPUT97), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n478), .A2(G142), .ZN(new_n883));
  OAI21_X1  g458(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n884));
  NOR2_X1   g459(.A1(new_n459), .A2(G118), .ZN(new_n885));
  XOR2_X1   g460(.A(new_n885), .B(KEYINPUT98), .Z(new_n886));
  OAI211_X1 g461(.A(new_n882), .B(new_n883), .C1(new_n884), .C2(new_n886), .ZN(new_n887));
  XNOR2_X1  g462(.A(new_n887), .B(new_n807), .ZN(new_n888));
  XNOR2_X1  g463(.A(new_n888), .B(new_n629), .ZN(new_n889));
  NOR2_X1   g464(.A1(new_n880), .A2(new_n889), .ZN(new_n890));
  INV_X1    g465(.A(new_n890), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n880), .A2(new_n889), .ZN(new_n892));
  XNOR2_X1  g467(.A(new_n487), .B(G160), .ZN(new_n893));
  XOR2_X1   g468(.A(new_n893), .B(new_n624), .Z(new_n894));
  NAND2_X1  g469(.A1(new_n894), .A2(KEYINPUT100), .ZN(new_n895));
  OR2_X1    g470(.A1(new_n894), .A2(KEYINPUT100), .ZN(new_n896));
  NAND4_X1  g471(.A1(new_n891), .A2(new_n892), .A3(new_n895), .A4(new_n896), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n892), .A2(KEYINPUT99), .ZN(new_n898));
  INV_X1    g473(.A(KEYINPUT99), .ZN(new_n899));
  NAND3_X1  g474(.A1(new_n880), .A2(new_n889), .A3(new_n899), .ZN(new_n900));
  AOI21_X1  g475(.A(new_n890), .B1(new_n898), .B2(new_n900), .ZN(new_n901));
  INV_X1    g476(.A(new_n894), .ZN(new_n902));
  OAI211_X1 g477(.A(new_n858), .B(new_n897), .C1(new_n901), .C2(new_n902), .ZN(new_n903));
  XNOR2_X1  g478(.A(new_n903), .B(KEYINPUT40), .ZN(G395));
  INV_X1    g479(.A(new_n852), .ZN(new_n905));
  INV_X1    g480(.A(new_n618), .ZN(new_n906));
  NAND2_X1  g481(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n852), .A2(new_n618), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n610), .A2(new_n605), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n606), .A2(G299), .ZN(new_n910));
  NAND3_X1  g485(.A1(new_n909), .A2(new_n910), .A3(KEYINPUT41), .ZN(new_n911));
  INV_X1    g486(.A(new_n911), .ZN(new_n912));
  AOI21_X1  g487(.A(KEYINPUT41), .B1(new_n909), .B2(new_n910), .ZN(new_n913));
  OAI211_X1 g488(.A(new_n907), .B(new_n908), .C1(new_n912), .C2(new_n913), .ZN(new_n914));
  INV_X1    g489(.A(KEYINPUT102), .ZN(new_n915));
  NOR2_X1   g490(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  INV_X1    g491(.A(new_n913), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n917), .A2(new_n911), .ZN(new_n918));
  INV_X1    g493(.A(new_n908), .ZN(new_n919));
  NOR2_X1   g494(.A1(new_n852), .A2(new_n618), .ZN(new_n920));
  NOR2_X1   g495(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  AOI21_X1  g496(.A(KEYINPUT102), .B1(new_n918), .B2(new_n921), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n909), .A2(new_n910), .ZN(new_n923));
  OAI21_X1  g498(.A(new_n923), .B1(new_n919), .B2(new_n920), .ZN(new_n924));
  NOR2_X1   g499(.A1(new_n924), .A2(KEYINPUT101), .ZN(new_n925));
  INV_X1    g500(.A(KEYINPUT101), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n907), .A2(new_n908), .ZN(new_n927));
  AOI21_X1  g502(.A(new_n926), .B1(new_n927), .B2(new_n923), .ZN(new_n928));
  OAI22_X1  g503(.A1(new_n916), .A2(new_n922), .B1(new_n925), .B2(new_n928), .ZN(new_n929));
  XNOR2_X1  g504(.A(KEYINPUT103), .B(KEYINPUT42), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  INV_X1    g506(.A(new_n930), .ZN(new_n932));
  OAI221_X1 g507(.A(new_n932), .B1(new_n925), .B2(new_n928), .C1(new_n916), .C2(new_n922), .ZN(new_n933));
  INV_X1    g508(.A(G290), .ZN(new_n934));
  XNOR2_X1  g509(.A(G303), .B(G288), .ZN(new_n935));
  XNOR2_X1  g510(.A(new_n934), .B(new_n935), .ZN(new_n936));
  XNOR2_X1  g511(.A(new_n936), .B(new_n793), .ZN(new_n937));
  AND3_X1   g512(.A1(new_n931), .A2(new_n933), .A3(new_n937), .ZN(new_n938));
  AOI21_X1  g513(.A(new_n937), .B1(new_n931), .B2(new_n933), .ZN(new_n939));
  OAI21_X1  g514(.A(G868), .B1(new_n938), .B2(new_n939), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n846), .A2(new_n616), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n940), .A2(new_n941), .ZN(G295));
  NAND2_X1  g517(.A1(new_n940), .A2(new_n941), .ZN(G331));
  INV_X1    g518(.A(KEYINPUT106), .ZN(new_n944));
  OAI21_X1  g519(.A(G168), .B1(G301), .B2(KEYINPUT104), .ZN(new_n945));
  INV_X1    g520(.A(KEYINPUT104), .ZN(new_n946));
  NOR3_X1   g521(.A1(G171), .A2(new_n946), .A3(KEYINPUT105), .ZN(new_n947));
  INV_X1    g522(.A(KEYINPUT105), .ZN(new_n948));
  AOI21_X1  g523(.A(new_n948), .B1(G301), .B2(KEYINPUT104), .ZN(new_n949));
  OAI21_X1  g524(.A(new_n945), .B1(new_n947), .B2(new_n949), .ZN(new_n950));
  OAI21_X1  g525(.A(KEYINPUT105), .B1(G171), .B2(new_n946), .ZN(new_n951));
  AOI21_X1  g526(.A(G286), .B1(G171), .B2(new_n946), .ZN(new_n952));
  NAND3_X1  g527(.A1(G301), .A2(KEYINPUT104), .A3(new_n948), .ZN(new_n953));
  NAND3_X1  g528(.A1(new_n951), .A2(new_n952), .A3(new_n953), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n950), .A2(new_n954), .ZN(new_n955));
  AOI21_X1  g530(.A(new_n944), .B1(new_n905), .B2(new_n955), .ZN(new_n956));
  INV_X1    g531(.A(new_n956), .ZN(new_n957));
  XNOR2_X1  g532(.A(new_n955), .B(new_n852), .ZN(new_n958));
  OAI211_X1 g533(.A(new_n923), .B(new_n957), .C1(new_n958), .C2(KEYINPUT106), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n905), .A2(new_n955), .ZN(new_n960));
  NAND3_X1  g535(.A1(new_n852), .A2(new_n954), .A3(new_n950), .ZN(new_n961));
  AOI22_X1  g536(.A1(new_n917), .A2(new_n911), .B1(new_n960), .B2(new_n961), .ZN(new_n962));
  INV_X1    g537(.A(new_n962), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n959), .A2(new_n963), .ZN(new_n964));
  XNOR2_X1  g539(.A(new_n936), .B(G305), .ZN(new_n965));
  OAI21_X1  g540(.A(new_n858), .B1(new_n964), .B2(new_n965), .ZN(new_n966));
  INV_X1    g541(.A(KEYINPUT43), .ZN(new_n967));
  AOI21_X1  g542(.A(KEYINPUT106), .B1(new_n960), .B2(new_n961), .ZN(new_n968));
  OAI21_X1  g543(.A(new_n918), .B1(new_n968), .B2(new_n956), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n958), .A2(new_n923), .ZN(new_n970));
  AOI21_X1  g545(.A(new_n937), .B1(new_n969), .B2(new_n970), .ZN(new_n971));
  NOR3_X1   g546(.A1(new_n966), .A2(new_n967), .A3(new_n971), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n960), .A2(new_n961), .ZN(new_n973));
  AOI21_X1  g548(.A(new_n956), .B1(new_n973), .B2(new_n944), .ZN(new_n974));
  AOI21_X1  g549(.A(new_n962), .B1(new_n974), .B2(new_n923), .ZN(new_n975));
  AOI21_X1  g550(.A(G37), .B1(new_n975), .B2(new_n937), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n964), .A2(new_n965), .ZN(new_n977));
  AOI21_X1  g552(.A(KEYINPUT43), .B1(new_n976), .B2(new_n977), .ZN(new_n978));
  OAI21_X1  g553(.A(KEYINPUT44), .B1(new_n972), .B2(new_n978), .ZN(new_n979));
  NOR3_X1   g554(.A1(new_n966), .A2(KEYINPUT43), .A3(new_n971), .ZN(new_n980));
  AOI21_X1  g555(.A(new_n967), .B1(new_n976), .B2(new_n977), .ZN(new_n981));
  NOR2_X1   g556(.A1(new_n980), .A2(new_n981), .ZN(new_n982));
  OAI21_X1  g557(.A(new_n979), .B1(new_n982), .B2(KEYINPUT44), .ZN(G397));
  XOR2_X1   g558(.A(KEYINPUT107), .B(G1384), .Z(new_n984));
  NAND2_X1  g559(.A1(new_n503), .A2(new_n984), .ZN(new_n985));
  INV_X1    g560(.A(G40), .ZN(new_n986));
  NOR3_X1   g561(.A1(new_n463), .A2(new_n475), .A3(new_n986), .ZN(new_n987));
  INV_X1    g562(.A(KEYINPUT45), .ZN(new_n988));
  NAND3_X1  g563(.A1(new_n985), .A2(new_n987), .A3(new_n988), .ZN(new_n989));
  OR2_X1    g564(.A1(new_n989), .A2(KEYINPUT108), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n989), .A2(KEYINPUT108), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n990), .A2(new_n991), .ZN(new_n992));
  NOR3_X1   g567(.A1(new_n992), .A2(G1996), .A3(new_n755), .ZN(new_n993));
  OR2_X1    g568(.A1(new_n993), .A2(KEYINPUT110), .ZN(new_n994));
  INV_X1    g569(.A(new_n992), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n704), .A2(new_n709), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n860), .A2(G2067), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n996), .A2(new_n997), .ZN(new_n998));
  AND2_X1   g573(.A1(new_n754), .A2(G1996), .ZN(new_n999));
  OAI21_X1  g574(.A(new_n995), .B1(new_n998), .B2(new_n999), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n993), .A2(KEYINPUT110), .ZN(new_n1001));
  NOR2_X1   g576(.A1(new_n807), .A2(new_n809), .ZN(new_n1002));
  AND2_X1   g577(.A1(new_n807), .A2(new_n809), .ZN(new_n1003));
  OAI21_X1  g578(.A(new_n995), .B1(new_n1002), .B2(new_n1003), .ZN(new_n1004));
  NAND4_X1  g579(.A1(new_n994), .A2(new_n1000), .A3(new_n1001), .A4(new_n1004), .ZN(new_n1005));
  OR2_X1    g580(.A1(G290), .A2(G1986), .ZN(new_n1006));
  XNOR2_X1  g581(.A(new_n1006), .B(KEYINPUT109), .ZN(new_n1007));
  NAND2_X1  g582(.A1(G290), .A2(G1986), .ZN(new_n1008));
  AOI21_X1  g583(.A(new_n992), .B1(new_n1007), .B2(new_n1008), .ZN(new_n1009));
  NOR2_X1   g584(.A1(new_n1005), .A2(new_n1009), .ZN(new_n1010));
  INV_X1    g585(.A(G8), .ZN(new_n1011));
  INV_X1    g586(.A(G1384), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n503), .A2(new_n1012), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n1013), .A2(new_n988), .ZN(new_n1014));
  INV_X1    g589(.A(KEYINPUT112), .ZN(new_n1015));
  NAND3_X1  g590(.A1(new_n1014), .A2(new_n1015), .A3(new_n987), .ZN(new_n1016));
  NAND3_X1  g591(.A1(new_n503), .A2(KEYINPUT45), .A3(new_n1012), .ZN(new_n1017));
  AOI21_X1  g592(.A(KEYINPUT45), .B1(new_n503), .B2(new_n1012), .ZN(new_n1018));
  NAND2_X1  g593(.A1(G160), .A2(G40), .ZN(new_n1019));
  OAI21_X1  g594(.A(KEYINPUT112), .B1(new_n1018), .B2(new_n1019), .ZN(new_n1020));
  NAND3_X1  g595(.A1(new_n1016), .A2(new_n1017), .A3(new_n1020), .ZN(new_n1021));
  INV_X1    g596(.A(G1966), .ZN(new_n1022));
  INV_X1    g597(.A(KEYINPUT50), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n1013), .A2(new_n1023), .ZN(new_n1024));
  NAND3_X1  g599(.A1(new_n503), .A2(KEYINPUT50), .A3(new_n1012), .ZN(new_n1025));
  AOI21_X1  g600(.A(new_n1019), .B1(new_n1024), .B2(new_n1025), .ZN(new_n1026));
  AOI22_X1  g601(.A1(new_n1021), .A2(new_n1022), .B1(new_n770), .B2(new_n1026), .ZN(new_n1027));
  AOI21_X1  g602(.A(new_n1011), .B1(new_n1027), .B2(G168), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n1021), .A2(new_n1022), .ZN(new_n1029));
  NAND2_X1  g604(.A1(new_n1026), .A2(new_n770), .ZN(new_n1030));
  NAND2_X1  g605(.A1(new_n1029), .A2(new_n1030), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n1031), .A2(G286), .ZN(new_n1032));
  NAND3_X1  g607(.A1(new_n1028), .A2(new_n1032), .A3(KEYINPUT51), .ZN(new_n1033));
  INV_X1    g608(.A(KEYINPUT51), .ZN(new_n1034));
  AOI221_X4 g609(.A(G286), .B1(new_n1026), .B2(new_n770), .C1(new_n1021), .C2(new_n1022), .ZN(new_n1035));
  OAI21_X1  g610(.A(new_n1034), .B1(new_n1035), .B2(new_n1011), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n1033), .A2(new_n1036), .ZN(new_n1037));
  INV_X1    g612(.A(KEYINPUT62), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n1037), .A2(new_n1038), .ZN(new_n1039));
  INV_X1    g614(.A(KEYINPUT49), .ZN(new_n1040));
  INV_X1    g615(.A(G1981), .ZN(new_n1041));
  AND2_X1   g616(.A1(new_n582), .A2(new_n583), .ZN(new_n1042));
  AOI21_X1  g617(.A(KEYINPUT75), .B1(new_n586), .B2(G651), .ZN(new_n1043));
  AOI211_X1 g618(.A(new_n579), .B(new_n539), .C1(new_n584), .C2(new_n585), .ZN(new_n1044));
  NOR2_X1   g619(.A1(new_n1043), .A2(new_n1044), .ZN(new_n1045));
  AOI21_X1  g620(.A(new_n1041), .B1(new_n1042), .B2(new_n1045), .ZN(new_n1046));
  NOR2_X1   g621(.A1(G305), .A2(G1981), .ZN(new_n1047));
  OAI21_X1  g622(.A(new_n1040), .B1(new_n1046), .B2(new_n1047), .ZN(new_n1048));
  NOR2_X1   g623(.A1(new_n1019), .A2(new_n1013), .ZN(new_n1049));
  NOR2_X1   g624(.A1(new_n1049), .A2(new_n1011), .ZN(new_n1050));
  NAND3_X1  g625(.A1(new_n1042), .A2(new_n1041), .A3(new_n1045), .ZN(new_n1051));
  NAND2_X1  g626(.A1(G305), .A2(G1981), .ZN(new_n1052));
  NAND3_X1  g627(.A1(new_n1051), .A2(new_n1052), .A3(KEYINPUT49), .ZN(new_n1053));
  NAND3_X1  g628(.A1(new_n1048), .A2(new_n1050), .A3(new_n1053), .ZN(new_n1054));
  INV_X1    g629(.A(G1976), .ZN(new_n1055));
  OR2_X1    g630(.A1(G288), .A2(new_n1055), .ZN(new_n1056));
  AOI21_X1  g631(.A(KEYINPUT52), .B1(G288), .B2(new_n1055), .ZN(new_n1057));
  NAND3_X1  g632(.A1(new_n1050), .A2(new_n1056), .A3(new_n1057), .ZN(new_n1058));
  NAND3_X1  g633(.A1(new_n987), .A2(new_n1012), .A3(new_n503), .ZN(new_n1059));
  NAND3_X1  g634(.A1(new_n1056), .A2(G8), .A3(new_n1059), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n1060), .A2(KEYINPUT52), .ZN(new_n1061));
  NAND3_X1  g636(.A1(new_n1054), .A2(new_n1058), .A3(new_n1061), .ZN(new_n1062));
  NAND3_X1  g637(.A1(new_n503), .A2(KEYINPUT45), .A3(new_n984), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n1063), .A2(new_n987), .ZN(new_n1064));
  OAI21_X1  g639(.A(new_n786), .B1(new_n1064), .B2(new_n1018), .ZN(new_n1065));
  INV_X1    g640(.A(G2090), .ZN(new_n1066));
  AND3_X1   g641(.A1(new_n503), .A2(KEYINPUT50), .A3(new_n1012), .ZN(new_n1067));
  AOI21_X1  g642(.A(KEYINPUT50), .B1(new_n503), .B2(new_n1012), .ZN(new_n1068));
  OAI211_X1 g643(.A(new_n1066), .B(new_n987), .C1(new_n1067), .C2(new_n1068), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n1065), .A2(new_n1069), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n1070), .A2(G8), .ZN(new_n1071));
  INV_X1    g646(.A(KEYINPUT55), .ZN(new_n1072));
  AND3_X1   g647(.A1(G303), .A2(new_n1072), .A3(G8), .ZN(new_n1073));
  AOI21_X1  g648(.A(new_n1072), .B1(G303), .B2(G8), .ZN(new_n1074));
  NOR2_X1   g649(.A1(new_n1073), .A2(new_n1074), .ZN(new_n1075));
  INV_X1    g650(.A(new_n1075), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n1071), .A2(new_n1076), .ZN(new_n1077));
  INV_X1    g652(.A(KEYINPUT111), .ZN(new_n1078));
  AOI21_X1  g653(.A(new_n1062), .B1(new_n1077), .B2(new_n1078), .ZN(new_n1079));
  AND3_X1   g654(.A1(new_n1070), .A2(G8), .A3(new_n1075), .ZN(new_n1080));
  AOI21_X1  g655(.A(new_n1075), .B1(new_n1070), .B2(G8), .ZN(new_n1081));
  OAI21_X1  g656(.A(KEYINPUT111), .B1(new_n1080), .B2(new_n1081), .ZN(new_n1082));
  AND2_X1   g657(.A1(new_n1079), .A2(new_n1082), .ZN(new_n1083));
  NAND4_X1  g658(.A1(new_n1014), .A2(new_n829), .A3(new_n987), .A4(new_n1063), .ZN(new_n1084));
  INV_X1    g659(.A(KEYINPUT53), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n1084), .A2(new_n1085), .ZN(new_n1086));
  OAI21_X1  g661(.A(new_n987), .B1(new_n1067), .B2(new_n1068), .ZN(new_n1087));
  XOR2_X1   g662(.A(KEYINPUT123), .B(G1961), .Z(new_n1088));
  NAND2_X1  g663(.A1(new_n1087), .A2(new_n1088), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n829), .A2(KEYINPUT53), .ZN(new_n1090));
  OAI211_X1 g665(.A(new_n1086), .B(new_n1089), .C1(new_n1021), .C2(new_n1090), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n1091), .A2(G171), .ZN(new_n1092));
  INV_X1    g667(.A(new_n1092), .ZN(new_n1093));
  NAND3_X1  g668(.A1(new_n1033), .A2(KEYINPUT62), .A3(new_n1036), .ZN(new_n1094));
  NAND4_X1  g669(.A1(new_n1039), .A2(new_n1083), .A3(new_n1093), .A4(new_n1094), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n1095), .A2(KEYINPUT125), .ZN(new_n1096));
  AND2_X1   g671(.A1(new_n1094), .A2(new_n1093), .ZN(new_n1097));
  INV_X1    g672(.A(KEYINPUT125), .ZN(new_n1098));
  NAND4_X1  g673(.A1(new_n1097), .A2(new_n1098), .A3(new_n1083), .A4(new_n1039), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n1096), .A2(new_n1099), .ZN(new_n1100));
  XNOR2_X1  g675(.A(KEYINPUT56), .B(G2072), .ZN(new_n1101));
  NAND4_X1  g676(.A1(new_n1014), .A2(new_n987), .A3(new_n1063), .A4(new_n1101), .ZN(new_n1102));
  INV_X1    g677(.A(KEYINPUT118), .ZN(new_n1103));
  NAND2_X1  g678(.A1(new_n1102), .A2(new_n1103), .ZN(new_n1104));
  AND2_X1   g679(.A1(new_n1063), .A2(new_n987), .ZN(new_n1105));
  NAND4_X1  g680(.A1(new_n1105), .A2(KEYINPUT118), .A3(new_n1014), .A4(new_n1101), .ZN(new_n1106));
  NAND2_X1  g681(.A1(new_n1104), .A2(new_n1106), .ZN(new_n1107));
  XOR2_X1   g682(.A(KEYINPUT114), .B(G1956), .Z(new_n1108));
  INV_X1    g683(.A(new_n1108), .ZN(new_n1109));
  NAND3_X1  g684(.A1(new_n1087), .A2(KEYINPUT115), .A3(new_n1109), .ZN(new_n1110));
  INV_X1    g685(.A(new_n1110), .ZN(new_n1111));
  AOI21_X1  g686(.A(KEYINPUT115), .B1(new_n1087), .B2(new_n1109), .ZN(new_n1112));
  OAI21_X1  g687(.A(new_n1107), .B1(new_n1111), .B2(new_n1112), .ZN(new_n1113));
  INV_X1    g688(.A(KEYINPUT117), .ZN(new_n1114));
  OR2_X1    g689(.A1(new_n1114), .A2(KEYINPUT57), .ZN(new_n1115));
  NAND3_X1  g690(.A1(new_n564), .A2(new_n570), .A3(new_n1115), .ZN(new_n1116));
  AOI22_X1  g691(.A1(new_n561), .A2(new_n563), .B1(G651), .B2(new_n569), .ZN(new_n1117));
  OAI211_X1 g692(.A(new_n1116), .B(new_n566), .C1(new_n1114), .C2(new_n1117), .ZN(new_n1118));
  OR2_X1    g693(.A1(KEYINPUT116), .A2(KEYINPUT57), .ZN(new_n1119));
  NAND3_X1  g694(.A1(G299), .A2(KEYINPUT116), .A3(KEYINPUT57), .ZN(new_n1120));
  NAND3_X1  g695(.A1(new_n1118), .A2(new_n1119), .A3(new_n1120), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n1113), .A2(new_n1121), .ZN(new_n1122));
  AND3_X1   g697(.A1(new_n1118), .A2(new_n1119), .A3(new_n1120), .ZN(new_n1123));
  INV_X1    g698(.A(KEYINPUT115), .ZN(new_n1124));
  OAI21_X1  g699(.A(new_n1124), .B1(new_n1026), .B2(new_n1108), .ZN(new_n1125));
  NAND2_X1  g700(.A1(new_n1125), .A2(new_n1110), .ZN(new_n1126));
  INV_X1    g701(.A(KEYINPUT121), .ZN(new_n1127));
  NAND4_X1  g702(.A1(new_n1123), .A2(new_n1126), .A3(new_n1127), .A4(new_n1107), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n1122), .A2(new_n1128), .ZN(new_n1129));
  AOI22_X1  g704(.A1(new_n1125), .A2(new_n1110), .B1(new_n1104), .B2(new_n1106), .ZN(new_n1130));
  OAI22_X1  g705(.A1(new_n1026), .A2(G1348), .B1(G2067), .B2(new_n1059), .ZN(new_n1131));
  AOI21_X1  g706(.A(KEYINPUT121), .B1(new_n1131), .B2(new_n606), .ZN(new_n1132));
  AOI22_X1  g707(.A1(new_n1123), .A2(new_n1130), .B1(new_n1132), .B2(KEYINPUT61), .ZN(new_n1133));
  OAI211_X1 g708(.A(new_n1036), .B(new_n1033), .C1(new_n1129), .C2(new_n1133), .ZN(new_n1134));
  INV_X1    g709(.A(new_n1134), .ZN(new_n1135));
  INV_X1    g710(.A(KEYINPUT54), .ZN(new_n1136));
  NAND2_X1  g711(.A1(new_n985), .A2(new_n988), .ZN(new_n1137));
  NAND4_X1  g712(.A1(new_n1105), .A2(KEYINPUT53), .A3(new_n829), .A4(new_n1137), .ZN(new_n1138));
  NAND3_X1  g713(.A1(new_n1086), .A2(new_n1138), .A3(new_n1089), .ZN(new_n1139));
  AOI21_X1  g714(.A(new_n1136), .B1(new_n1139), .B2(G171), .ZN(new_n1140));
  OAI21_X1  g715(.A(new_n1140), .B1(G171), .B2(new_n1091), .ZN(new_n1141));
  INV_X1    g716(.A(KEYINPUT61), .ZN(new_n1142));
  NAND3_X1  g717(.A1(new_n1130), .A2(new_n1142), .A3(new_n1123), .ZN(new_n1143));
  AND4_X1   g718(.A1(new_n1082), .A2(new_n1141), .A3(new_n1079), .A4(new_n1143), .ZN(new_n1144));
  NAND4_X1  g719(.A1(new_n1086), .A2(new_n1138), .A3(new_n1089), .A4(G301), .ZN(new_n1145));
  NAND2_X1  g720(.A1(new_n1092), .A2(new_n1145), .ZN(new_n1146));
  AOI21_X1  g721(.A(KEYINPUT124), .B1(new_n1146), .B2(new_n1136), .ZN(new_n1147));
  INV_X1    g722(.A(KEYINPUT124), .ZN(new_n1148));
  AOI211_X1 g723(.A(new_n1148), .B(KEYINPUT54), .C1(new_n1092), .C2(new_n1145), .ZN(new_n1149));
  NOR2_X1   g724(.A1(new_n1147), .A2(new_n1149), .ZN(new_n1150));
  OAI211_X1 g725(.A(new_n606), .B(new_n1131), .C1(new_n1113), .C2(new_n1121), .ZN(new_n1151));
  XOR2_X1   g726(.A(new_n605), .B(KEYINPUT122), .Z(new_n1152));
  AOI22_X1  g727(.A1(new_n1087), .A2(new_n714), .B1(new_n709), .B2(new_n1049), .ZN(new_n1153));
  NAND2_X1  g728(.A1(new_n1153), .A2(KEYINPUT60), .ZN(new_n1154));
  NOR2_X1   g729(.A1(new_n1152), .A2(new_n1154), .ZN(new_n1155));
  OAI22_X1  g730(.A1(new_n1153), .A2(KEYINPUT60), .B1(KEYINPUT122), .B2(new_n606), .ZN(new_n1156));
  AOI21_X1  g731(.A(new_n1155), .B1(new_n1154), .B2(new_n1156), .ZN(new_n1157));
  INV_X1    g732(.A(G1996), .ZN(new_n1158));
  NAND3_X1  g733(.A1(new_n1105), .A2(new_n1158), .A3(new_n1014), .ZN(new_n1159));
  XOR2_X1   g734(.A(KEYINPUT58), .B(G1341), .Z(new_n1160));
  NAND2_X1  g735(.A1(new_n1059), .A2(new_n1160), .ZN(new_n1161));
  AOI21_X1  g736(.A(new_n551), .B1(new_n1159), .B2(new_n1161), .ZN(new_n1162));
  NAND2_X1  g737(.A1(KEYINPUT119), .A2(KEYINPUT59), .ZN(new_n1163));
  XOR2_X1   g738(.A(new_n1163), .B(KEYINPUT120), .Z(new_n1164));
  XNOR2_X1  g739(.A(new_n1162), .B(new_n1164), .ZN(new_n1165));
  OAI211_X1 g740(.A(new_n1122), .B(new_n1151), .C1(new_n1157), .C2(new_n1165), .ZN(new_n1166));
  NAND4_X1  g741(.A1(new_n1135), .A2(new_n1144), .A3(new_n1150), .A4(new_n1166), .ZN(new_n1167));
  NOR3_X1   g742(.A1(new_n1027), .A2(new_n1011), .A3(G286), .ZN(new_n1168));
  NAND3_X1  g743(.A1(new_n1079), .A2(new_n1082), .A3(new_n1168), .ZN(new_n1169));
  INV_X1    g744(.A(KEYINPUT63), .ZN(new_n1170));
  NAND2_X1  g745(.A1(new_n1169), .A2(new_n1170), .ZN(new_n1171));
  NAND2_X1  g746(.A1(new_n1171), .A2(KEYINPUT113), .ZN(new_n1172));
  INV_X1    g747(.A(KEYINPUT113), .ZN(new_n1173));
  NAND3_X1  g748(.A1(new_n1169), .A2(new_n1173), .A3(new_n1170), .ZN(new_n1174));
  NOR2_X1   g749(.A1(new_n1080), .A2(new_n1081), .ZN(new_n1175));
  INV_X1    g750(.A(new_n1062), .ZN(new_n1176));
  NAND4_X1  g751(.A1(new_n1168), .A2(new_n1175), .A3(KEYINPUT63), .A4(new_n1176), .ZN(new_n1177));
  NAND3_X1  g752(.A1(new_n1172), .A2(new_n1174), .A3(new_n1177), .ZN(new_n1178));
  NAND2_X1  g753(.A1(new_n1054), .A2(new_n1055), .ZN(new_n1179));
  OAI21_X1  g754(.A(new_n1051), .B1(new_n1179), .B2(G288), .ZN(new_n1180));
  AOI22_X1  g755(.A1(new_n1180), .A2(new_n1050), .B1(new_n1176), .B2(new_n1080), .ZN(new_n1181));
  NAND3_X1  g756(.A1(new_n1167), .A2(new_n1178), .A3(new_n1181), .ZN(new_n1182));
  OAI21_X1  g757(.A(new_n1010), .B1(new_n1100), .B2(new_n1182), .ZN(new_n1183));
  NOR2_X1   g758(.A1(new_n1007), .A2(new_n992), .ZN(new_n1184));
  XNOR2_X1  g759(.A(new_n1184), .B(KEYINPUT48), .ZN(new_n1185));
  NOR2_X1   g760(.A1(new_n1185), .A2(new_n1005), .ZN(new_n1186));
  XOR2_X1   g761(.A(new_n1002), .B(KEYINPUT126), .Z(new_n1187));
  NAND4_X1  g762(.A1(new_n994), .A2(new_n1000), .A3(new_n1001), .A4(new_n1187), .ZN(new_n1188));
  AOI21_X1  g763(.A(new_n992), .B1(new_n1188), .B2(new_n996), .ZN(new_n1189));
  NOR2_X1   g764(.A1(new_n992), .A2(G1996), .ZN(new_n1190));
  OR2_X1    g765(.A1(new_n1190), .A2(KEYINPUT46), .ZN(new_n1191));
  OAI21_X1  g766(.A(new_n995), .B1(new_n754), .B2(new_n998), .ZN(new_n1192));
  NAND2_X1  g767(.A1(new_n1190), .A2(KEYINPUT46), .ZN(new_n1193));
  NAND3_X1  g768(.A1(new_n1191), .A2(new_n1192), .A3(new_n1193), .ZN(new_n1194));
  XOR2_X1   g769(.A(new_n1194), .B(KEYINPUT47), .Z(new_n1195));
  NOR3_X1   g770(.A1(new_n1186), .A2(new_n1189), .A3(new_n1195), .ZN(new_n1196));
  NAND2_X1  g771(.A1(new_n1183), .A2(new_n1196), .ZN(G329));
  assign    G231 = 1'b0;
  OAI21_X1  g772(.A(new_n695), .B1(new_n980), .B2(new_n981), .ZN(new_n1199));
  NAND3_X1  g773(.A1(new_n656), .A2(G319), .A3(new_n672), .ZN(new_n1200));
  INV_X1    g774(.A(KEYINPUT127), .ZN(new_n1201));
  NAND2_X1  g775(.A1(new_n1200), .A2(new_n1201), .ZN(new_n1202));
  NAND4_X1  g776(.A1(new_n656), .A2(KEYINPUT127), .A3(G319), .A4(new_n672), .ZN(new_n1203));
  NAND2_X1  g777(.A1(new_n1202), .A2(new_n1203), .ZN(new_n1204));
  NAND2_X1  g778(.A1(new_n903), .A2(new_n1204), .ZN(new_n1205));
  NOR2_X1   g779(.A1(new_n1199), .A2(new_n1205), .ZN(G308));
  AND2_X1   g780(.A1(new_n969), .A2(new_n970), .ZN(new_n1207));
  OAI211_X1 g781(.A(new_n976), .B(new_n967), .C1(new_n937), .C2(new_n1207), .ZN(new_n1208));
  AND2_X1   g782(.A1(new_n976), .A2(new_n977), .ZN(new_n1209));
  OAI21_X1  g783(.A(new_n1208), .B1(new_n1209), .B2(new_n967), .ZN(new_n1210));
  NAND4_X1  g784(.A1(new_n1210), .A2(new_n695), .A3(new_n903), .A4(new_n1204), .ZN(G225));
endmodule


