//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 0 0 0 1 1 0 1 0 0 1 1 0 0 1 0 0 1 0 0 0 1 1 0 1 0 0 0 0 0 1 0 1 1 1 1 0 1 0 1 0 1 0 0 0 1 0 1 0 0 1 0 0 1 0 1 1 1 1 0 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:17:36 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n630,
    new_n631, new_n632, new_n633, new_n635, new_n636, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n709, new_n710, new_n711, new_n712, new_n714, new_n715,
    new_n716, new_n717, new_n718, new_n720, new_n721, new_n722, new_n724,
    new_n725, new_n726, new_n727, new_n728, new_n729, new_n730, new_n731,
    new_n732, new_n733, new_n734, new_n735, new_n736, new_n737, new_n738,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n758, new_n759, new_n760, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n812, new_n813,
    new_n814, new_n815, new_n816, new_n817, new_n819, new_n820, new_n822,
    new_n823, new_n824, new_n825, new_n826, new_n827, new_n828, new_n829,
    new_n830, new_n831, new_n832, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n882, new_n883, new_n885, new_n886, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n897, new_n898,
    new_n899, new_n901, new_n902, new_n903, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n928, new_n929, new_n930, new_n931,
    new_n932, new_n933, new_n934, new_n935, new_n937, new_n938, new_n939,
    new_n940;
  XNOR2_X1  g000(.A(G15gat), .B(G22gat), .ZN(new_n202));
  NAND2_X1  g001(.A1(new_n202), .A2(KEYINPUT89), .ZN(new_n203));
  INV_X1    g002(.A(G1gat), .ZN(new_n204));
  NAND2_X1  g003(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  NAND3_X1  g004(.A1(new_n202), .A2(KEYINPUT89), .A3(G1gat), .ZN(new_n206));
  INV_X1    g005(.A(KEYINPUT16), .ZN(new_n207));
  NAND2_X1  g006(.A1(new_n202), .A2(new_n207), .ZN(new_n208));
  NAND3_X1  g007(.A1(new_n205), .A2(new_n206), .A3(new_n208), .ZN(new_n209));
  OR2_X1    g008(.A1(new_n209), .A2(G8gat), .ZN(new_n210));
  NAND2_X1  g009(.A1(new_n209), .A2(G8gat), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  INV_X1    g011(.A(KEYINPUT90), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  NAND3_X1  g013(.A1(new_n210), .A2(KEYINPUT90), .A3(new_n211), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n214), .A2(new_n215), .ZN(new_n216));
  NOR2_X1   g015(.A1(G29gat), .A2(G36gat), .ZN(new_n217));
  INV_X1    g016(.A(KEYINPUT14), .ZN(new_n218));
  XNOR2_X1  g017(.A(new_n217), .B(new_n218), .ZN(new_n219));
  INV_X1    g018(.A(G29gat), .ZN(new_n220));
  INV_X1    g019(.A(G36gat), .ZN(new_n221));
  OAI21_X1  g020(.A(new_n219), .B1(new_n220), .B2(new_n221), .ZN(new_n222));
  XNOR2_X1  g021(.A(G43gat), .B(G50gat), .ZN(new_n223));
  NAND3_X1  g022(.A1(new_n222), .A2(KEYINPUT15), .A3(new_n223), .ZN(new_n224));
  OAI21_X1  g023(.A(KEYINPUT88), .B1(new_n220), .B2(new_n221), .ZN(new_n225));
  OR3_X1    g024(.A1(new_n220), .A2(new_n221), .A3(KEYINPUT88), .ZN(new_n226));
  NAND3_X1  g025(.A1(new_n219), .A2(new_n225), .A3(new_n226), .ZN(new_n227));
  XNOR2_X1  g026(.A(new_n223), .B(KEYINPUT15), .ZN(new_n228));
  OAI21_X1  g027(.A(new_n224), .B1(new_n227), .B2(new_n228), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n216), .A2(new_n229), .ZN(new_n230));
  NAND2_X1  g029(.A1(G229gat), .A2(G233gat), .ZN(new_n231));
  XNOR2_X1  g030(.A(new_n229), .B(KEYINPUT17), .ZN(new_n232));
  INV_X1    g031(.A(new_n212), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n232), .A2(new_n233), .ZN(new_n234));
  NAND3_X1  g033(.A1(new_n230), .A2(new_n231), .A3(new_n234), .ZN(new_n235));
  NOR2_X1   g034(.A1(KEYINPUT91), .A2(KEYINPUT18), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n235), .A2(new_n236), .ZN(new_n237));
  XNOR2_X1  g036(.A(KEYINPUT92), .B(KEYINPUT13), .ZN(new_n238));
  XNOR2_X1  g037(.A(new_n238), .B(new_n231), .ZN(new_n239));
  NOR2_X1   g038(.A1(new_n216), .A2(new_n229), .ZN(new_n240));
  INV_X1    g039(.A(new_n229), .ZN(new_n241));
  AOI21_X1  g040(.A(new_n241), .B1(new_n214), .B2(new_n215), .ZN(new_n242));
  OAI21_X1  g041(.A(new_n239), .B1(new_n240), .B2(new_n242), .ZN(new_n243));
  INV_X1    g042(.A(new_n236), .ZN(new_n244));
  NAND4_X1  g043(.A1(new_n230), .A2(new_n234), .A3(new_n231), .A4(new_n244), .ZN(new_n245));
  NAND3_X1  g044(.A1(new_n237), .A2(new_n243), .A3(new_n245), .ZN(new_n246));
  XNOR2_X1  g045(.A(G113gat), .B(G141gat), .ZN(new_n247));
  XNOR2_X1  g046(.A(new_n247), .B(G197gat), .ZN(new_n248));
  XOR2_X1   g047(.A(KEYINPUT11), .B(G169gat), .Z(new_n249));
  XNOR2_X1  g048(.A(new_n248), .B(new_n249), .ZN(new_n250));
  XOR2_X1   g049(.A(new_n250), .B(KEYINPUT12), .Z(new_n251));
  NAND2_X1  g050(.A1(new_n246), .A2(new_n251), .ZN(new_n252));
  INV_X1    g051(.A(new_n251), .ZN(new_n253));
  NAND4_X1  g052(.A1(new_n237), .A2(new_n253), .A3(new_n243), .A4(new_n245), .ZN(new_n254));
  AND2_X1   g053(.A1(new_n252), .A2(new_n254), .ZN(new_n255));
  XNOR2_X1  g054(.A(G1gat), .B(G29gat), .ZN(new_n256));
  XNOR2_X1  g055(.A(new_n256), .B(KEYINPUT0), .ZN(new_n257));
  XNOR2_X1  g056(.A(G57gat), .B(G85gat), .ZN(new_n258));
  XOR2_X1   g057(.A(new_n257), .B(new_n258), .Z(new_n259));
  INV_X1    g058(.A(new_n259), .ZN(new_n260));
  INV_X1    g059(.A(KEYINPUT5), .ZN(new_n261));
  XOR2_X1   g060(.A(G155gat), .B(G162gat), .Z(new_n262));
  XOR2_X1   g061(.A(G141gat), .B(G148gat), .Z(new_n263));
  AOI21_X1  g062(.A(new_n262), .B1(KEYINPUT77), .B2(new_n263), .ZN(new_n264));
  INV_X1    g063(.A(G155gat), .ZN(new_n265));
  INV_X1    g064(.A(G162gat), .ZN(new_n266));
  OAI21_X1  g065(.A(KEYINPUT2), .B1(new_n265), .B2(new_n266), .ZN(new_n267));
  NAND2_X1  g066(.A1(new_n263), .A2(new_n267), .ZN(new_n268));
  XNOR2_X1  g067(.A(new_n264), .B(new_n268), .ZN(new_n269));
  XNOR2_X1  g068(.A(G113gat), .B(G120gat), .ZN(new_n270));
  INV_X1    g069(.A(KEYINPUT67), .ZN(new_n271));
  OR2_X1    g070(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  INV_X1    g071(.A(KEYINPUT1), .ZN(new_n273));
  XNOR2_X1  g072(.A(G127gat), .B(G134gat), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n270), .A2(new_n271), .ZN(new_n275));
  NAND4_X1  g074(.A1(new_n272), .A2(new_n273), .A3(new_n274), .A4(new_n275), .ZN(new_n276));
  INV_X1    g075(.A(KEYINPUT66), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n274), .A2(new_n277), .ZN(new_n278));
  INV_X1    g077(.A(G127gat), .ZN(new_n279));
  NAND3_X1  g078(.A1(new_n279), .A2(KEYINPUT66), .A3(G134gat), .ZN(new_n280));
  OAI211_X1 g079(.A(new_n278), .B(new_n280), .C1(KEYINPUT1), .C2(new_n270), .ZN(new_n281));
  AND2_X1   g080(.A1(new_n276), .A2(new_n281), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n269), .A2(new_n282), .ZN(new_n283));
  INV_X1    g082(.A(KEYINPUT79), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  NAND3_X1  g084(.A1(new_n269), .A2(new_n282), .A3(KEYINPUT79), .ZN(new_n286));
  NAND3_X1  g085(.A1(new_n285), .A2(KEYINPUT4), .A3(new_n286), .ZN(new_n287));
  INV_X1    g086(.A(KEYINPUT81), .ZN(new_n288));
  OR2_X1    g087(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  OAI211_X1 g088(.A(new_n287), .B(new_n288), .C1(KEYINPUT4), .C2(new_n283), .ZN(new_n290));
  XOR2_X1   g089(.A(new_n264), .B(new_n268), .Z(new_n291));
  NOR2_X1   g090(.A1(new_n291), .A2(KEYINPUT3), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n276), .A2(new_n281), .ZN(new_n293));
  INV_X1    g092(.A(KEYINPUT3), .ZN(new_n294));
  OAI21_X1  g093(.A(new_n293), .B1(new_n269), .B2(new_n294), .ZN(new_n295));
  NOR2_X1   g094(.A1(new_n292), .A2(new_n295), .ZN(new_n296));
  NAND2_X1  g095(.A1(G225gat), .A2(G233gat), .ZN(new_n297));
  XNOR2_X1  g096(.A(new_n297), .B(KEYINPUT78), .ZN(new_n298));
  NOR2_X1   g097(.A1(new_n296), .A2(new_n298), .ZN(new_n299));
  AND4_X1   g098(.A1(new_n261), .A2(new_n289), .A3(new_n290), .A4(new_n299), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n291), .A2(new_n293), .ZN(new_n301));
  NAND3_X1  g100(.A1(new_n285), .A2(new_n286), .A3(new_n301), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n302), .A2(new_n298), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n303), .A2(KEYINPUT5), .ZN(new_n304));
  INV_X1    g103(.A(new_n298), .ZN(new_n305));
  NAND3_X1  g104(.A1(new_n269), .A2(new_n282), .A3(KEYINPUT4), .ZN(new_n306));
  OAI211_X1 g105(.A(new_n305), .B(new_n306), .C1(new_n292), .C2(new_n295), .ZN(new_n307));
  INV_X1    g106(.A(new_n307), .ZN(new_n308));
  INV_X1    g107(.A(KEYINPUT4), .ZN(new_n309));
  NAND3_X1  g108(.A1(new_n285), .A2(new_n309), .A3(new_n286), .ZN(new_n310));
  NAND3_X1  g109(.A1(new_n308), .A2(KEYINPUT80), .A3(new_n310), .ZN(new_n311));
  INV_X1    g110(.A(KEYINPUT80), .ZN(new_n312));
  AND3_X1   g111(.A1(new_n285), .A2(new_n309), .A3(new_n286), .ZN(new_n313));
  OAI21_X1  g112(.A(new_n312), .B1(new_n313), .B2(new_n307), .ZN(new_n314));
  AOI21_X1  g113(.A(new_n304), .B1(new_n311), .B2(new_n314), .ZN(new_n315));
  OAI21_X1  g114(.A(new_n260), .B1(new_n300), .B2(new_n315), .ZN(new_n316));
  INV_X1    g115(.A(KEYINPUT6), .ZN(new_n317));
  AOI21_X1  g116(.A(new_n261), .B1(new_n302), .B2(new_n298), .ZN(new_n318));
  AOI21_X1  g117(.A(KEYINPUT80), .B1(new_n308), .B2(new_n310), .ZN(new_n319));
  NOR3_X1   g118(.A1(new_n313), .A2(new_n307), .A3(new_n312), .ZN(new_n320));
  OAI21_X1  g119(.A(new_n318), .B1(new_n319), .B2(new_n320), .ZN(new_n321));
  NAND4_X1  g120(.A1(new_n289), .A2(new_n290), .A3(new_n261), .A4(new_n299), .ZN(new_n322));
  NAND3_X1  g121(.A1(new_n321), .A2(new_n259), .A3(new_n322), .ZN(new_n323));
  NAND3_X1  g122(.A1(new_n316), .A2(new_n317), .A3(new_n323), .ZN(new_n324));
  INV_X1    g123(.A(KEYINPUT82), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n324), .A2(new_n325), .ZN(new_n326));
  NAND4_X1  g125(.A1(new_n316), .A2(new_n323), .A3(KEYINPUT82), .A4(new_n317), .ZN(new_n327));
  AOI211_X1 g126(.A(new_n317), .B(new_n259), .C1(new_n321), .C2(new_n322), .ZN(new_n328));
  INV_X1    g127(.A(new_n328), .ZN(new_n329));
  NAND3_X1  g128(.A1(new_n326), .A2(new_n327), .A3(new_n329), .ZN(new_n330));
  NAND2_X1  g129(.A1(G169gat), .A2(G176gat), .ZN(new_n331));
  INV_X1    g130(.A(new_n331), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n332), .A2(KEYINPUT64), .ZN(new_n333));
  INV_X1    g132(.A(KEYINPUT64), .ZN(new_n334));
  NAND2_X1  g133(.A1(new_n331), .A2(new_n334), .ZN(new_n335));
  NOR2_X1   g134(.A1(G169gat), .A2(G176gat), .ZN(new_n336));
  OAI211_X1 g135(.A(new_n333), .B(new_n335), .C1(KEYINPUT23), .C2(new_n336), .ZN(new_n337));
  INV_X1    g136(.A(KEYINPUT24), .ZN(new_n338));
  NAND3_X1  g137(.A1(new_n338), .A2(G183gat), .A3(G190gat), .ZN(new_n339));
  XNOR2_X1  g138(.A(G183gat), .B(G190gat), .ZN(new_n340));
  OAI21_X1  g139(.A(new_n339), .B1(new_n340), .B2(new_n338), .ZN(new_n341));
  INV_X1    g140(.A(KEYINPUT25), .ZN(new_n342));
  AND2_X1   g141(.A1(new_n336), .A2(KEYINPUT23), .ZN(new_n343));
  NOR4_X1   g142(.A1(new_n337), .A2(new_n341), .A3(new_n342), .A4(new_n343), .ZN(new_n344));
  INV_X1    g143(.A(new_n341), .ZN(new_n345));
  NOR2_X1   g144(.A1(new_n336), .A2(KEYINPUT23), .ZN(new_n346));
  NOR3_X1   g145(.A1(new_n343), .A2(new_n346), .A3(new_n332), .ZN(new_n347));
  AOI21_X1  g146(.A(KEYINPUT25), .B1(new_n345), .B2(new_n347), .ZN(new_n348));
  NOR2_X1   g147(.A1(new_n344), .A2(new_n348), .ZN(new_n349));
  INV_X1    g148(.A(new_n349), .ZN(new_n350));
  XNOR2_X1  g149(.A(KEYINPUT27), .B(G183gat), .ZN(new_n351));
  INV_X1    g150(.A(G190gat), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n351), .A2(new_n352), .ZN(new_n353));
  AND2_X1   g152(.A1(KEYINPUT65), .A2(KEYINPUT28), .ZN(new_n354));
  NOR2_X1   g153(.A1(KEYINPUT65), .A2(KEYINPUT28), .ZN(new_n355));
  OR3_X1    g154(.A1(new_n353), .A2(new_n354), .A3(new_n355), .ZN(new_n356));
  AOI22_X1  g155(.A1(new_n353), .A2(new_n354), .B1(G183gat), .B2(G190gat), .ZN(new_n357));
  XNOR2_X1  g156(.A(new_n336), .B(KEYINPUT26), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n358), .A2(new_n331), .ZN(new_n359));
  NAND3_X1  g158(.A1(new_n356), .A2(new_n357), .A3(new_n359), .ZN(new_n360));
  AOI21_X1  g159(.A(KEYINPUT29), .B1(new_n350), .B2(new_n360), .ZN(new_n361));
  NAND2_X1  g160(.A1(G226gat), .A2(G233gat), .ZN(new_n362));
  XOR2_X1   g161(.A(new_n362), .B(KEYINPUT72), .Z(new_n363));
  OAI21_X1  g162(.A(KEYINPUT74), .B1(new_n361), .B2(new_n363), .ZN(new_n364));
  INV_X1    g163(.A(KEYINPUT22), .ZN(new_n365));
  INV_X1    g164(.A(G211gat), .ZN(new_n366));
  INV_X1    g165(.A(G218gat), .ZN(new_n367));
  OAI21_X1  g166(.A(new_n365), .B1(new_n366), .B2(new_n367), .ZN(new_n368));
  OR2_X1    g167(.A1(new_n368), .A2(KEYINPUT71), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n368), .A2(KEYINPUT71), .ZN(new_n370));
  XNOR2_X1  g169(.A(G197gat), .B(G204gat), .ZN(new_n371));
  NAND3_X1  g170(.A1(new_n369), .A2(new_n370), .A3(new_n371), .ZN(new_n372));
  XOR2_X1   g171(.A(G211gat), .B(G218gat), .Z(new_n373));
  XOR2_X1   g172(.A(new_n372), .B(new_n373), .Z(new_n374));
  INV_X1    g173(.A(new_n374), .ZN(new_n375));
  XOR2_X1   g174(.A(new_n363), .B(KEYINPUT73), .Z(new_n376));
  INV_X1    g175(.A(new_n360), .ZN(new_n377));
  OAI21_X1  g176(.A(new_n376), .B1(new_n349), .B2(new_n377), .ZN(new_n378));
  INV_X1    g177(.A(KEYINPUT74), .ZN(new_n379));
  INV_X1    g178(.A(new_n363), .ZN(new_n380));
  NOR2_X1   g179(.A1(new_n349), .A2(new_n377), .ZN(new_n381));
  OAI211_X1 g180(.A(new_n379), .B(new_n380), .C1(new_n381), .C2(KEYINPUT29), .ZN(new_n382));
  NAND4_X1  g181(.A1(new_n364), .A2(new_n375), .A3(new_n378), .A4(new_n382), .ZN(new_n383));
  XNOR2_X1  g182(.A(G8gat), .B(G36gat), .ZN(new_n384));
  XNOR2_X1  g183(.A(G64gat), .B(G92gat), .ZN(new_n385));
  XOR2_X1   g184(.A(new_n384), .B(new_n385), .Z(new_n386));
  OAI22_X1  g185(.A1(new_n361), .A2(new_n376), .B1(new_n381), .B2(new_n380), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n387), .A2(new_n374), .ZN(new_n388));
  NAND3_X1  g187(.A1(new_n383), .A2(new_n386), .A3(new_n388), .ZN(new_n389));
  INV_X1    g188(.A(KEYINPUT30), .ZN(new_n390));
  AND3_X1   g189(.A1(new_n389), .A2(KEYINPUT76), .A3(new_n390), .ZN(new_n391));
  AOI21_X1  g190(.A(new_n390), .B1(new_n389), .B2(KEYINPUT76), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n383), .A2(new_n388), .ZN(new_n393));
  XOR2_X1   g192(.A(new_n386), .B(KEYINPUT75), .Z(new_n394));
  AND2_X1   g193(.A1(new_n393), .A2(new_n394), .ZN(new_n395));
  NOR3_X1   g194(.A1(new_n391), .A2(new_n392), .A3(new_n395), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n330), .A2(new_n396), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n381), .A2(new_n293), .ZN(new_n398));
  OAI21_X1  g197(.A(new_n282), .B1(new_n349), .B2(new_n377), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n398), .A2(new_n399), .ZN(new_n400));
  INV_X1    g199(.A(G227gat), .ZN(new_n401));
  INV_X1    g200(.A(G233gat), .ZN(new_n402));
  NOR2_X1   g201(.A1(new_n401), .A2(new_n402), .ZN(new_n403));
  INV_X1    g202(.A(new_n403), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n400), .A2(new_n404), .ZN(new_n405));
  AND2_X1   g204(.A1(new_n405), .A2(KEYINPUT34), .ZN(new_n406));
  NOR2_X1   g205(.A1(new_n405), .A2(KEYINPUT34), .ZN(new_n407));
  NOR2_X1   g206(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  INV_X1    g207(.A(new_n408), .ZN(new_n409));
  INV_X1    g208(.A(KEYINPUT32), .ZN(new_n410));
  NAND3_X1  g209(.A1(new_n398), .A2(new_n403), .A3(new_n399), .ZN(new_n411));
  INV_X1    g210(.A(KEYINPUT68), .ZN(new_n412));
  NAND2_X1  g211(.A1(new_n411), .A2(new_n412), .ZN(new_n413));
  NAND4_X1  g212(.A1(new_n398), .A2(new_n399), .A3(KEYINPUT68), .A4(new_n403), .ZN(new_n414));
  AOI21_X1  g213(.A(new_n410), .B1(new_n413), .B2(new_n414), .ZN(new_n415));
  AOI21_X1  g214(.A(KEYINPUT33), .B1(new_n413), .B2(new_n414), .ZN(new_n416));
  XOR2_X1   g215(.A(G15gat), .B(G43gat), .Z(new_n417));
  XNOR2_X1  g216(.A(G71gat), .B(G99gat), .ZN(new_n418));
  XNOR2_X1  g217(.A(new_n417), .B(new_n418), .ZN(new_n419));
  INV_X1    g218(.A(new_n419), .ZN(new_n420));
  NOR3_X1   g219(.A1(new_n415), .A2(new_n416), .A3(new_n420), .ZN(new_n421));
  AOI221_X4 g220(.A(new_n410), .B1(KEYINPUT33), .B2(new_n419), .C1(new_n413), .C2(new_n414), .ZN(new_n422));
  OAI21_X1  g221(.A(new_n409), .B1(new_n421), .B2(new_n422), .ZN(new_n423));
  INV_X1    g222(.A(KEYINPUT69), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n423), .A2(new_n424), .ZN(new_n425));
  OAI21_X1  g224(.A(new_n374), .B1(new_n292), .B2(KEYINPUT29), .ZN(new_n426));
  INV_X1    g225(.A(KEYINPUT29), .ZN(new_n427));
  AOI21_X1  g226(.A(KEYINPUT3), .B1(new_n375), .B2(new_n427), .ZN(new_n428));
  OAI21_X1  g227(.A(new_n426), .B1(new_n428), .B2(new_n269), .ZN(new_n429));
  XOR2_X1   g228(.A(G78gat), .B(G106gat), .Z(new_n430));
  XNOR2_X1  g229(.A(new_n429), .B(new_n430), .ZN(new_n431));
  NAND2_X1  g230(.A1(G228gat), .A2(G233gat), .ZN(new_n432));
  XNOR2_X1  g231(.A(new_n432), .B(G22gat), .ZN(new_n433));
  XOR2_X1   g232(.A(KEYINPUT31), .B(G50gat), .Z(new_n434));
  XNOR2_X1  g233(.A(new_n433), .B(new_n434), .ZN(new_n435));
  XOR2_X1   g234(.A(new_n431), .B(new_n435), .Z(new_n436));
  OAI211_X1 g235(.A(KEYINPUT69), .B(new_n409), .C1(new_n421), .C2(new_n422), .ZN(new_n437));
  NOR2_X1   g236(.A1(new_n416), .A2(new_n420), .ZN(new_n438));
  INV_X1    g237(.A(new_n415), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n438), .A2(new_n439), .ZN(new_n440));
  INV_X1    g239(.A(new_n422), .ZN(new_n441));
  NAND3_X1  g240(.A1(new_n440), .A2(new_n408), .A3(new_n441), .ZN(new_n442));
  NAND4_X1  g241(.A1(new_n425), .A2(new_n436), .A3(new_n437), .A4(new_n442), .ZN(new_n443));
  OAI21_X1  g242(.A(KEYINPUT35), .B1(new_n397), .B2(new_n443), .ZN(new_n444));
  INV_X1    g243(.A(new_n396), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n423), .A2(new_n442), .ZN(new_n446));
  NOR2_X1   g245(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  INV_X1    g246(.A(new_n436), .ZN(new_n448));
  NOR2_X1   g247(.A1(new_n448), .A2(KEYINPUT35), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n329), .A2(new_n324), .ZN(new_n450));
  NAND3_X1  g249(.A1(new_n447), .A2(new_n449), .A3(new_n450), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n444), .A2(new_n451), .ZN(new_n452));
  INV_X1    g251(.A(new_n296), .ZN(new_n453));
  NAND3_X1  g252(.A1(new_n289), .A2(new_n290), .A3(new_n453), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n454), .A2(new_n298), .ZN(new_n455));
  OR2_X1    g254(.A1(new_n455), .A2(KEYINPUT39), .ZN(new_n456));
  OR2_X1    g255(.A1(new_n302), .A2(new_n298), .ZN(new_n457));
  NAND3_X1  g256(.A1(new_n455), .A2(KEYINPUT39), .A3(new_n457), .ZN(new_n458));
  NAND3_X1  g257(.A1(new_n456), .A2(new_n259), .A3(new_n458), .ZN(new_n459));
  INV_X1    g258(.A(KEYINPUT40), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  NAND4_X1  g260(.A1(new_n456), .A2(KEYINPUT40), .A3(new_n259), .A4(new_n458), .ZN(new_n462));
  NAND3_X1  g261(.A1(new_n461), .A2(new_n316), .A3(new_n462), .ZN(new_n463));
  OAI21_X1  g262(.A(new_n436), .B1(new_n463), .B2(new_n396), .ZN(new_n464));
  XNOR2_X1  g263(.A(KEYINPUT84), .B(KEYINPUT38), .ZN(new_n465));
  AOI21_X1  g264(.A(new_n386), .B1(new_n393), .B2(KEYINPUT37), .ZN(new_n466));
  INV_X1    g265(.A(KEYINPUT37), .ZN(new_n467));
  NAND3_X1  g266(.A1(new_n383), .A2(new_n467), .A3(new_n388), .ZN(new_n468));
  AOI21_X1  g267(.A(new_n465), .B1(new_n466), .B2(new_n468), .ZN(new_n469));
  INV_X1    g268(.A(new_n389), .ZN(new_n470));
  AOI21_X1  g269(.A(new_n467), .B1(new_n387), .B2(new_n375), .ZN(new_n471));
  NAND4_X1  g270(.A1(new_n364), .A2(new_n374), .A3(new_n378), .A4(new_n382), .ZN(new_n472));
  AND3_X1   g271(.A1(new_n471), .A2(new_n472), .A3(KEYINPUT83), .ZN(new_n473));
  AOI21_X1  g272(.A(KEYINPUT83), .B1(new_n471), .B2(new_n472), .ZN(new_n474));
  NOR2_X1   g273(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  NAND3_X1  g274(.A1(new_n468), .A2(new_n394), .A3(new_n465), .ZN(new_n476));
  NOR2_X1   g275(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  INV_X1    g276(.A(KEYINPUT85), .ZN(new_n478));
  AOI21_X1  g277(.A(new_n470), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n321), .A2(new_n322), .ZN(new_n480));
  AOI21_X1  g279(.A(KEYINPUT6), .B1(new_n480), .B2(new_n260), .ZN(new_n481));
  AOI21_X1  g280(.A(new_n328), .B1(new_n481), .B2(new_n323), .ZN(new_n482));
  OAI21_X1  g281(.A(KEYINPUT85), .B1(new_n475), .B2(new_n476), .ZN(new_n483));
  NAND3_X1  g282(.A1(new_n479), .A2(new_n482), .A3(new_n483), .ZN(new_n484));
  AOI21_X1  g283(.A(new_n469), .B1(new_n484), .B2(KEYINPUT86), .ZN(new_n485));
  INV_X1    g284(.A(KEYINPUT86), .ZN(new_n486));
  NAND4_X1  g285(.A1(new_n479), .A2(new_n482), .A3(new_n486), .A4(new_n483), .ZN(new_n487));
  AOI21_X1  g286(.A(new_n464), .B1(new_n485), .B2(new_n487), .ZN(new_n488));
  NAND2_X1  g287(.A1(new_n397), .A2(new_n448), .ZN(new_n489));
  INV_X1    g288(.A(KEYINPUT36), .ZN(new_n490));
  AOI21_X1  g289(.A(KEYINPUT70), .B1(new_n423), .B2(new_n442), .ZN(new_n491));
  INV_X1    g290(.A(new_n491), .ZN(new_n492));
  NAND3_X1  g291(.A1(new_n425), .A2(new_n437), .A3(new_n442), .ZN(new_n493));
  AOI21_X1  g292(.A(new_n490), .B1(new_n492), .B2(new_n493), .ZN(new_n494));
  NAND3_X1  g293(.A1(new_n446), .A2(KEYINPUT70), .A3(new_n490), .ZN(new_n495));
  INV_X1    g294(.A(new_n495), .ZN(new_n496));
  OAI21_X1  g295(.A(new_n489), .B1(new_n494), .B2(new_n496), .ZN(new_n497));
  OAI21_X1  g296(.A(new_n452), .B1(new_n488), .B2(new_n497), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n498), .A2(KEYINPUT87), .ZN(new_n499));
  INV_X1    g298(.A(KEYINPUT87), .ZN(new_n500));
  OAI211_X1 g299(.A(new_n500), .B(new_n452), .C1(new_n488), .C2(new_n497), .ZN(new_n501));
  AOI21_X1  g300(.A(new_n255), .B1(new_n499), .B2(new_n501), .ZN(new_n502));
  INV_X1    g301(.A(KEYINPUT95), .ZN(new_n503));
  INV_X1    g302(.A(G71gat), .ZN(new_n504));
  INV_X1    g303(.A(G78gat), .ZN(new_n505));
  NOR2_X1   g304(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  NOR2_X1   g305(.A1(G71gat), .A2(G78gat), .ZN(new_n507));
  AOI21_X1  g306(.A(new_n506), .B1(KEYINPUT9), .B2(new_n507), .ZN(new_n508));
  INV_X1    g307(.A(G57gat), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n509), .A2(KEYINPUT93), .ZN(new_n510));
  INV_X1    g309(.A(KEYINPUT93), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n511), .A2(G57gat), .ZN(new_n512));
  NAND3_X1  g311(.A1(new_n510), .A2(new_n512), .A3(G64gat), .ZN(new_n513));
  OR2_X1    g312(.A1(new_n509), .A2(G64gat), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  INV_X1    g314(.A(KEYINPUT94), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  NAND3_X1  g316(.A1(new_n513), .A2(KEYINPUT94), .A3(new_n514), .ZN(new_n518));
  AOI21_X1  g317(.A(new_n508), .B1(new_n517), .B2(new_n518), .ZN(new_n519));
  XOR2_X1   g318(.A(G57gat), .B(G64gat), .Z(new_n520));
  NAND2_X1  g319(.A1(new_n520), .A2(KEYINPUT9), .ZN(new_n521));
  NOR2_X1   g320(.A1(new_n506), .A2(new_n507), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  INV_X1    g322(.A(new_n523), .ZN(new_n524));
  OAI21_X1  g323(.A(new_n503), .B1(new_n519), .B2(new_n524), .ZN(new_n525));
  INV_X1    g324(.A(new_n508), .ZN(new_n526));
  AND3_X1   g325(.A1(new_n513), .A2(KEYINPUT94), .A3(new_n514), .ZN(new_n527));
  AOI21_X1  g326(.A(KEYINPUT94), .B1(new_n513), .B2(new_n514), .ZN(new_n528));
  OAI21_X1  g327(.A(new_n526), .B1(new_n527), .B2(new_n528), .ZN(new_n529));
  NAND3_X1  g328(.A1(new_n529), .A2(KEYINPUT95), .A3(new_n523), .ZN(new_n530));
  NAND2_X1  g329(.A1(new_n525), .A2(new_n530), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n531), .A2(KEYINPUT21), .ZN(new_n532));
  NAND3_X1  g331(.A1(new_n532), .A2(new_n215), .A3(new_n214), .ZN(new_n533));
  XNOR2_X1  g332(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n534));
  XOR2_X1   g333(.A(new_n533), .B(new_n534), .Z(new_n535));
  INV_X1    g334(.A(new_n535), .ZN(new_n536));
  NOR2_X1   g335(.A1(new_n531), .A2(KEYINPUT21), .ZN(new_n537));
  NAND2_X1  g336(.A1(G231gat), .A2(G233gat), .ZN(new_n538));
  XNOR2_X1  g337(.A(new_n537), .B(new_n538), .ZN(new_n539));
  XNOR2_X1  g338(.A(G127gat), .B(G155gat), .ZN(new_n540));
  XNOR2_X1  g339(.A(new_n540), .B(KEYINPUT96), .ZN(new_n541));
  XNOR2_X1  g340(.A(new_n539), .B(new_n541), .ZN(new_n542));
  XOR2_X1   g341(.A(G183gat), .B(G211gat), .Z(new_n543));
  INV_X1    g342(.A(new_n543), .ZN(new_n544));
  NAND2_X1  g343(.A1(new_n542), .A2(new_n544), .ZN(new_n545));
  INV_X1    g344(.A(new_n545), .ZN(new_n546));
  NOR2_X1   g345(.A1(new_n542), .A2(new_n544), .ZN(new_n547));
  OAI21_X1  g346(.A(new_n536), .B1(new_n546), .B2(new_n547), .ZN(new_n548));
  INV_X1    g347(.A(new_n547), .ZN(new_n549));
  NAND3_X1  g348(.A1(new_n549), .A2(new_n535), .A3(new_n545), .ZN(new_n550));
  XNOR2_X1  g349(.A(G190gat), .B(G218gat), .ZN(new_n551));
  INV_X1    g350(.A(new_n551), .ZN(new_n552));
  NAND2_X1  g351(.A1(G85gat), .A2(G92gat), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n553), .A2(KEYINPUT7), .ZN(new_n554));
  INV_X1    g353(.A(KEYINPUT7), .ZN(new_n555));
  NAND3_X1  g354(.A1(new_n555), .A2(G85gat), .A3(G92gat), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n554), .A2(new_n556), .ZN(new_n557));
  NAND2_X1  g356(.A1(G99gat), .A2(G106gat), .ZN(new_n558));
  INV_X1    g357(.A(G85gat), .ZN(new_n559));
  INV_X1    g358(.A(G92gat), .ZN(new_n560));
  AOI22_X1  g359(.A1(KEYINPUT8), .A2(new_n558), .B1(new_n559), .B2(new_n560), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n557), .A2(new_n561), .ZN(new_n562));
  OR2_X1    g361(.A1(G99gat), .A2(G106gat), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n563), .A2(new_n558), .ZN(new_n564));
  XOR2_X1   g363(.A(new_n562), .B(new_n564), .Z(new_n565));
  INV_X1    g364(.A(new_n565), .ZN(new_n566));
  AND2_X1   g365(.A1(G232gat), .A2(G233gat), .ZN(new_n567));
  AOI22_X1  g366(.A1(new_n566), .A2(new_n229), .B1(KEYINPUT41), .B2(new_n567), .ZN(new_n568));
  INV_X1    g367(.A(new_n232), .ZN(new_n569));
  OAI211_X1 g368(.A(new_n552), .B(new_n568), .C1(new_n569), .C2(new_n566), .ZN(new_n570));
  INV_X1    g369(.A(KEYINPUT98), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  NOR2_X1   g371(.A1(new_n567), .A2(KEYINPUT41), .ZN(new_n573));
  XOR2_X1   g372(.A(new_n573), .B(KEYINPUT97), .Z(new_n574));
  XNOR2_X1  g373(.A(new_n574), .B(G134gat), .ZN(new_n575));
  XNOR2_X1  g374(.A(new_n575), .B(new_n266), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n572), .A2(new_n576), .ZN(new_n577));
  OAI21_X1  g376(.A(new_n568), .B1(new_n569), .B2(new_n566), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n578), .A2(new_n551), .ZN(new_n579));
  NAND2_X1  g378(.A1(new_n579), .A2(new_n570), .ZN(new_n580));
  NAND2_X1  g379(.A1(new_n577), .A2(new_n580), .ZN(new_n581));
  NAND4_X1  g380(.A1(new_n579), .A2(KEYINPUT98), .A3(new_n570), .A4(new_n576), .ZN(new_n582));
  NAND2_X1  g381(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  INV_X1    g382(.A(new_n583), .ZN(new_n584));
  NAND3_X1  g383(.A1(new_n548), .A2(new_n550), .A3(new_n584), .ZN(new_n585));
  NAND3_X1  g384(.A1(new_n563), .A2(KEYINPUT99), .A3(new_n558), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n562), .A2(new_n586), .ZN(new_n587));
  AND3_X1   g386(.A1(new_n563), .A2(KEYINPUT99), .A3(new_n558), .ZN(new_n588));
  NAND3_X1  g387(.A1(new_n588), .A2(new_n557), .A3(new_n561), .ZN(new_n589));
  NAND2_X1  g388(.A1(new_n587), .A2(new_n589), .ZN(new_n590));
  NAND3_X1  g389(.A1(new_n529), .A2(new_n523), .A3(new_n590), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n591), .A2(KEYINPUT100), .ZN(new_n592));
  INV_X1    g391(.A(KEYINPUT100), .ZN(new_n593));
  NAND4_X1  g392(.A1(new_n529), .A2(new_n593), .A3(new_n590), .A4(new_n523), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n592), .A2(new_n594), .ZN(new_n595));
  INV_X1    g394(.A(KEYINPUT10), .ZN(new_n596));
  NAND3_X1  g395(.A1(new_n525), .A2(new_n565), .A3(new_n530), .ZN(new_n597));
  NAND3_X1  g396(.A1(new_n595), .A2(new_n596), .A3(new_n597), .ZN(new_n598));
  NAND3_X1  g397(.A1(new_n531), .A2(KEYINPUT10), .A3(new_n566), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  NAND2_X1  g399(.A1(new_n600), .A2(KEYINPUT101), .ZN(new_n601));
  NAND2_X1  g400(.A1(G230gat), .A2(G233gat), .ZN(new_n602));
  INV_X1    g401(.A(KEYINPUT101), .ZN(new_n603));
  NAND3_X1  g402(.A1(new_n598), .A2(new_n599), .A3(new_n603), .ZN(new_n604));
  NAND3_X1  g403(.A1(new_n601), .A2(new_n602), .A3(new_n604), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n595), .A2(new_n597), .ZN(new_n606));
  INV_X1    g405(.A(new_n602), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  XNOR2_X1  g407(.A(G120gat), .B(G148gat), .ZN(new_n609));
  XNOR2_X1  g408(.A(G176gat), .B(G204gat), .ZN(new_n610));
  XOR2_X1   g409(.A(new_n609), .B(new_n610), .Z(new_n611));
  NAND3_X1  g410(.A1(new_n605), .A2(new_n608), .A3(new_n611), .ZN(new_n612));
  NAND2_X1  g411(.A1(new_n600), .A2(new_n602), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n613), .A2(new_n608), .ZN(new_n614));
  INV_X1    g413(.A(new_n611), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n612), .A2(new_n616), .ZN(new_n617));
  NOR2_X1   g416(.A1(new_n585), .A2(new_n617), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n502), .A2(new_n618), .ZN(new_n619));
  NOR2_X1   g418(.A1(new_n619), .A2(new_n330), .ZN(new_n620));
  XNOR2_X1  g419(.A(new_n620), .B(new_n204), .ZN(G1324gat));
  INV_X1    g420(.A(G8gat), .ZN(new_n622));
  INV_X1    g421(.A(new_n619), .ZN(new_n623));
  AOI21_X1  g422(.A(new_n622), .B1(new_n623), .B2(new_n445), .ZN(new_n624));
  NOR2_X1   g423(.A1(new_n207), .A2(new_n622), .ZN(new_n625));
  NOR2_X1   g424(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n626));
  NOR4_X1   g425(.A1(new_n619), .A2(new_n396), .A3(new_n625), .A4(new_n626), .ZN(new_n627));
  OAI21_X1  g426(.A(KEYINPUT42), .B1(new_n624), .B2(new_n627), .ZN(new_n628));
  OAI21_X1  g427(.A(new_n628), .B1(KEYINPUT42), .B2(new_n627), .ZN(G1325gat));
  NOR2_X1   g428(.A1(new_n494), .A2(new_n496), .ZN(new_n630));
  INV_X1    g429(.A(new_n630), .ZN(new_n631));
  OAI21_X1  g430(.A(G15gat), .B1(new_n619), .B2(new_n631), .ZN(new_n632));
  OR2_X1    g431(.A1(new_n446), .A2(G15gat), .ZN(new_n633));
  OAI21_X1  g432(.A(new_n632), .B1(new_n619), .B2(new_n633), .ZN(G1326gat));
  NOR2_X1   g433(.A1(new_n619), .A2(new_n436), .ZN(new_n635));
  XOR2_X1   g434(.A(KEYINPUT43), .B(G22gat), .Z(new_n636));
  XNOR2_X1  g435(.A(new_n635), .B(new_n636), .ZN(G1327gat));
  INV_X1    g436(.A(KEYINPUT44), .ZN(new_n638));
  NOR2_X1   g437(.A1(new_n584), .A2(new_n638), .ZN(new_n639));
  INV_X1    g438(.A(new_n501), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n437), .A2(new_n442), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n440), .A2(new_n441), .ZN(new_n642));
  AOI21_X1  g441(.A(KEYINPUT69), .B1(new_n642), .B2(new_n409), .ZN(new_n643));
  NOR2_X1   g442(.A1(new_n641), .A2(new_n643), .ZN(new_n644));
  OAI21_X1  g443(.A(KEYINPUT36), .B1(new_n644), .B2(new_n491), .ZN(new_n645));
  AOI22_X1  g444(.A1(new_n645), .A2(new_n495), .B1(new_n397), .B2(new_n448), .ZN(new_n646));
  AND3_X1   g445(.A1(new_n461), .A2(new_n316), .A3(new_n462), .ZN(new_n647));
  AOI21_X1  g446(.A(new_n448), .B1(new_n647), .B2(new_n445), .ZN(new_n648));
  AND3_X1   g447(.A1(new_n468), .A2(new_n394), .A3(new_n465), .ZN(new_n649));
  OAI211_X1 g448(.A(new_n649), .B(new_n478), .C1(new_n474), .C2(new_n473), .ZN(new_n650));
  NAND3_X1  g449(.A1(new_n650), .A2(new_n483), .A3(new_n389), .ZN(new_n651));
  OAI21_X1  g450(.A(KEYINPUT86), .B1(new_n651), .B2(new_n450), .ZN(new_n652));
  INV_X1    g451(.A(new_n469), .ZN(new_n653));
  NAND3_X1  g452(.A1(new_n652), .A2(new_n487), .A3(new_n653), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n648), .A2(new_n654), .ZN(new_n655));
  NAND2_X1  g454(.A1(new_n646), .A2(new_n655), .ZN(new_n656));
  AOI21_X1  g455(.A(new_n500), .B1(new_n656), .B2(new_n452), .ZN(new_n657));
  OAI21_X1  g456(.A(new_n639), .B1(new_n640), .B2(new_n657), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n498), .A2(new_n583), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n659), .A2(new_n638), .ZN(new_n660));
  AND2_X1   g459(.A1(new_n658), .A2(new_n660), .ZN(new_n661));
  NAND2_X1  g460(.A1(new_n548), .A2(new_n550), .ZN(new_n662));
  INV_X1    g461(.A(new_n662), .ZN(new_n663));
  NOR2_X1   g462(.A1(new_n663), .A2(new_n617), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n252), .A2(new_n254), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  XOR2_X1   g465(.A(new_n666), .B(KEYINPUT102), .Z(new_n667));
  NAND2_X1  g466(.A1(new_n661), .A2(new_n667), .ZN(new_n668));
  OAI21_X1  g467(.A(G29gat), .B1(new_n668), .B2(new_n330), .ZN(new_n669));
  INV_X1    g468(.A(KEYINPUT45), .ZN(new_n670));
  NAND2_X1  g469(.A1(new_n664), .A2(new_n583), .ZN(new_n671));
  INV_X1    g470(.A(new_n671), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n502), .A2(new_n672), .ZN(new_n673));
  INV_X1    g472(.A(new_n330), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n674), .A2(new_n220), .ZN(new_n675));
  OAI21_X1  g474(.A(new_n670), .B1(new_n673), .B2(new_n675), .ZN(new_n676));
  OR3_X1    g475(.A1(new_n673), .A2(new_n670), .A3(new_n675), .ZN(new_n677));
  NAND3_X1  g476(.A1(new_n669), .A2(new_n676), .A3(new_n677), .ZN(G1328gat));
  INV_X1    g477(.A(new_n673), .ZN(new_n679));
  NAND3_X1  g478(.A1(new_n679), .A2(new_n221), .A3(new_n445), .ZN(new_n680));
  INV_X1    g479(.A(KEYINPUT46), .ZN(new_n681));
  NOR2_X1   g480(.A1(new_n681), .A2(KEYINPUT103), .ZN(new_n682));
  AND2_X1   g481(.A1(new_n681), .A2(KEYINPUT103), .ZN(new_n683));
  OAI21_X1  g482(.A(new_n680), .B1(new_n682), .B2(new_n683), .ZN(new_n684));
  OAI21_X1  g483(.A(G36gat), .B1(new_n668), .B2(new_n396), .ZN(new_n685));
  OAI211_X1 g484(.A(new_n684), .B(new_n685), .C1(new_n682), .C2(new_n680), .ZN(G1329gat));
  NAND4_X1  g485(.A1(new_n661), .A2(G43gat), .A3(new_n630), .A4(new_n667), .ZN(new_n687));
  INV_X1    g486(.A(G43gat), .ZN(new_n688));
  OAI21_X1  g487(.A(new_n688), .B1(new_n673), .B2(new_n446), .ZN(new_n689));
  XNOR2_X1  g488(.A(KEYINPUT104), .B(KEYINPUT47), .ZN(new_n690));
  AND3_X1   g489(.A1(new_n687), .A2(new_n689), .A3(new_n690), .ZN(new_n691));
  AOI21_X1  g490(.A(new_n690), .B1(new_n687), .B2(new_n689), .ZN(new_n692));
  NOR2_X1   g491(.A1(new_n691), .A2(new_n692), .ZN(G1330gat));
  INV_X1    g492(.A(G50gat), .ZN(new_n694));
  NAND3_X1  g493(.A1(new_n679), .A2(new_n694), .A3(new_n448), .ZN(new_n695));
  AOI21_X1  g494(.A(KEYINPUT48), .B1(new_n695), .B2(KEYINPUT105), .ZN(new_n696));
  NAND4_X1  g495(.A1(new_n658), .A2(new_n448), .A3(new_n660), .A4(new_n667), .ZN(new_n697));
  NAND2_X1  g496(.A1(new_n697), .A2(G50gat), .ZN(new_n698));
  NAND2_X1  g497(.A1(new_n695), .A2(new_n698), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n696), .A2(new_n699), .ZN(new_n700));
  OAI211_X1 g499(.A(new_n695), .B(new_n698), .C1(KEYINPUT105), .C2(KEYINPUT48), .ZN(new_n701));
  NAND2_X1  g500(.A1(new_n700), .A2(new_n701), .ZN(G1331gat));
  INV_X1    g501(.A(new_n617), .ZN(new_n703));
  NOR3_X1   g502(.A1(new_n585), .A2(new_n665), .A3(new_n703), .ZN(new_n704));
  AND2_X1   g503(.A1(new_n498), .A2(new_n704), .ZN(new_n705));
  NAND2_X1  g504(.A1(new_n705), .A2(new_n674), .ZN(new_n706));
  NAND2_X1  g505(.A1(new_n510), .A2(new_n512), .ZN(new_n707));
  XNOR2_X1  g506(.A(new_n706), .B(new_n707), .ZN(G1332gat));
  AOI21_X1  g507(.A(new_n396), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n705), .A2(new_n709), .ZN(new_n710));
  XOR2_X1   g509(.A(new_n710), .B(KEYINPUT106), .Z(new_n711));
  NOR2_X1   g510(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n712));
  XNOR2_X1  g511(.A(new_n711), .B(new_n712), .ZN(G1333gat));
  NAND2_X1  g512(.A1(new_n498), .A2(new_n704), .ZN(new_n714));
  NOR3_X1   g513(.A1(new_n714), .A2(new_n504), .A3(new_n631), .ZN(new_n715));
  XNOR2_X1  g514(.A(new_n715), .B(KEYINPUT107), .ZN(new_n716));
  OAI21_X1  g515(.A(new_n504), .B1(new_n714), .B2(new_n446), .ZN(new_n717));
  NAND2_X1  g516(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  XNOR2_X1  g517(.A(new_n718), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g518(.A1(new_n705), .A2(new_n448), .ZN(new_n720));
  XNOR2_X1  g519(.A(new_n720), .B(KEYINPUT109), .ZN(new_n721));
  XNOR2_X1  g520(.A(KEYINPUT108), .B(G78gat), .ZN(new_n722));
  XNOR2_X1  g521(.A(new_n721), .B(new_n722), .ZN(G1335gat));
  NAND3_X1  g522(.A1(new_n498), .A2(KEYINPUT111), .A3(new_n583), .ZN(new_n724));
  NOR2_X1   g523(.A1(new_n663), .A2(new_n665), .ZN(new_n725));
  NAND2_X1  g524(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  INV_X1    g525(.A(new_n726), .ZN(new_n727));
  AOI21_X1  g526(.A(KEYINPUT111), .B1(new_n498), .B2(new_n583), .ZN(new_n728));
  INV_X1    g527(.A(new_n728), .ZN(new_n729));
  AOI21_X1  g528(.A(KEYINPUT51), .B1(new_n727), .B2(new_n729), .ZN(new_n730));
  INV_X1    g529(.A(KEYINPUT51), .ZN(new_n731));
  NOR3_X1   g530(.A1(new_n726), .A2(new_n731), .A3(new_n728), .ZN(new_n732));
  OR2_X1    g531(.A1(new_n730), .A2(new_n732), .ZN(new_n733));
  NAND4_X1  g532(.A1(new_n733), .A2(new_n559), .A3(new_n674), .A4(new_n617), .ZN(new_n734));
  NAND3_X1  g533(.A1(new_n662), .A2(new_n255), .A3(new_n617), .ZN(new_n735));
  XOR2_X1   g534(.A(new_n735), .B(KEYINPUT110), .Z(new_n736));
  NAND2_X1  g535(.A1(new_n661), .A2(new_n736), .ZN(new_n737));
  OAI21_X1  g536(.A(G85gat), .B1(new_n737), .B2(new_n330), .ZN(new_n738));
  NAND2_X1  g537(.A1(new_n734), .A2(new_n738), .ZN(G1336gat));
  NOR2_X1   g538(.A1(new_n396), .A2(G92gat), .ZN(new_n740));
  OAI211_X1 g539(.A(new_n617), .B(new_n740), .C1(new_n730), .C2(new_n732), .ZN(new_n741));
  XOR2_X1   g540(.A(KEYINPUT114), .B(KEYINPUT52), .Z(new_n742));
  NAND4_X1  g541(.A1(new_n658), .A2(new_n445), .A3(new_n660), .A4(new_n736), .ZN(new_n743));
  AOI21_X1  g542(.A(new_n742), .B1(new_n743), .B2(G92gat), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n741), .A2(new_n744), .ZN(new_n745));
  AND2_X1   g544(.A1(new_n743), .A2(G92gat), .ZN(new_n746));
  XOR2_X1   g545(.A(KEYINPUT112), .B(KEYINPUT51), .Z(new_n747));
  OAI21_X1  g546(.A(new_n747), .B1(new_n726), .B2(new_n728), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n748), .A2(KEYINPUT113), .ZN(new_n749));
  NAND3_X1  g548(.A1(new_n727), .A2(KEYINPUT51), .A3(new_n729), .ZN(new_n750));
  INV_X1    g549(.A(KEYINPUT113), .ZN(new_n751));
  OAI211_X1 g550(.A(new_n751), .B(new_n747), .C1(new_n726), .C2(new_n728), .ZN(new_n752));
  NAND3_X1  g551(.A1(new_n749), .A2(new_n750), .A3(new_n752), .ZN(new_n753));
  NOR3_X1   g552(.A1(new_n396), .A2(G92gat), .A3(new_n703), .ZN(new_n754));
  AOI21_X1  g553(.A(new_n746), .B1(new_n753), .B2(new_n754), .ZN(new_n755));
  INV_X1    g554(.A(KEYINPUT52), .ZN(new_n756));
  OAI21_X1  g555(.A(new_n745), .B1(new_n755), .B2(new_n756), .ZN(G1337gat));
  NOR2_X1   g556(.A1(new_n446), .A2(G99gat), .ZN(new_n758));
  NAND3_X1  g557(.A1(new_n733), .A2(new_n617), .A3(new_n758), .ZN(new_n759));
  OAI21_X1  g558(.A(G99gat), .B1(new_n737), .B2(new_n631), .ZN(new_n760));
  NAND2_X1  g559(.A1(new_n759), .A2(new_n760), .ZN(G1338gat));
  NOR2_X1   g560(.A1(new_n436), .A2(G106gat), .ZN(new_n762));
  OAI211_X1 g561(.A(new_n617), .B(new_n762), .C1(new_n730), .C2(new_n732), .ZN(new_n763));
  NAND4_X1  g562(.A1(new_n658), .A2(new_n448), .A3(new_n660), .A4(new_n736), .ZN(new_n764));
  AOI21_X1  g563(.A(KEYINPUT53), .B1(new_n764), .B2(G106gat), .ZN(new_n765));
  NAND2_X1  g564(.A1(new_n763), .A2(new_n765), .ZN(new_n766));
  AND2_X1   g565(.A1(new_n764), .A2(G106gat), .ZN(new_n767));
  NOR3_X1   g566(.A1(new_n436), .A2(G106gat), .A3(new_n703), .ZN(new_n768));
  AOI21_X1  g567(.A(new_n767), .B1(new_n753), .B2(new_n768), .ZN(new_n769));
  INV_X1    g568(.A(KEYINPUT53), .ZN(new_n770));
  OAI21_X1  g569(.A(new_n766), .B1(new_n769), .B2(new_n770), .ZN(G1339gat));
  NOR2_X1   g570(.A1(new_n613), .A2(KEYINPUT54), .ZN(new_n772));
  NOR2_X1   g571(.A1(new_n772), .A2(new_n611), .ZN(new_n773));
  INV_X1    g572(.A(KEYINPUT115), .ZN(new_n774));
  NAND3_X1  g573(.A1(new_n598), .A2(new_n599), .A3(new_n607), .ZN(new_n775));
  AND2_X1   g574(.A1(new_n775), .A2(KEYINPUT54), .ZN(new_n776));
  AND3_X1   g575(.A1(new_n605), .A2(new_n774), .A3(new_n776), .ZN(new_n777));
  AOI21_X1  g576(.A(new_n774), .B1(new_n605), .B2(new_n776), .ZN(new_n778));
  OAI21_X1  g577(.A(new_n773), .B1(new_n777), .B2(new_n778), .ZN(new_n779));
  INV_X1    g578(.A(KEYINPUT55), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  OAI211_X1 g580(.A(KEYINPUT55), .B(new_n773), .C1(new_n777), .C2(new_n778), .ZN(new_n782));
  NAND4_X1  g581(.A1(new_n781), .A2(new_n665), .A3(new_n612), .A4(new_n782), .ZN(new_n783));
  NOR3_X1   g582(.A1(new_n240), .A2(new_n242), .A3(new_n239), .ZN(new_n784));
  AOI21_X1  g583(.A(new_n231), .B1(new_n230), .B2(new_n234), .ZN(new_n785));
  OAI21_X1  g584(.A(new_n250), .B1(new_n784), .B2(new_n785), .ZN(new_n786));
  AND2_X1   g585(.A1(new_n254), .A2(new_n786), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n787), .A2(new_n617), .ZN(new_n788));
  AOI21_X1  g587(.A(new_n583), .B1(new_n783), .B2(new_n788), .ZN(new_n789));
  AND2_X1   g588(.A1(new_n782), .A2(new_n612), .ZN(new_n790));
  AND2_X1   g589(.A1(new_n787), .A2(new_n583), .ZN(new_n791));
  AND3_X1   g590(.A1(new_n790), .A2(new_n781), .A3(new_n791), .ZN(new_n792));
  OAI21_X1  g591(.A(KEYINPUT116), .B1(new_n789), .B2(new_n792), .ZN(new_n793));
  INV_X1    g592(.A(KEYINPUT116), .ZN(new_n794));
  NAND3_X1  g593(.A1(new_n790), .A2(new_n781), .A3(new_n791), .ZN(new_n795));
  INV_X1    g594(.A(new_n788), .ZN(new_n796));
  AOI21_X1  g595(.A(new_n255), .B1(new_n780), .B2(new_n779), .ZN(new_n797));
  AOI21_X1  g596(.A(new_n796), .B1(new_n797), .B2(new_n790), .ZN(new_n798));
  OAI211_X1 g597(.A(new_n794), .B(new_n795), .C1(new_n798), .C2(new_n583), .ZN(new_n799));
  NAND3_X1  g598(.A1(new_n793), .A2(new_n799), .A3(new_n662), .ZN(new_n800));
  NOR3_X1   g599(.A1(new_n585), .A2(new_n665), .A3(new_n617), .ZN(new_n801));
  INV_X1    g600(.A(new_n801), .ZN(new_n802));
  AOI21_X1  g601(.A(new_n448), .B1(new_n800), .B2(new_n802), .ZN(new_n803));
  AND2_X1   g602(.A1(new_n803), .A2(new_n674), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n804), .A2(new_n447), .ZN(new_n805));
  INV_X1    g604(.A(G113gat), .ZN(new_n806));
  NOR3_X1   g605(.A1(new_n805), .A2(new_n806), .A3(new_n255), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n804), .A2(new_n644), .ZN(new_n808));
  NOR2_X1   g607(.A1(new_n808), .A2(new_n445), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n809), .A2(new_n665), .ZN(new_n810));
  AOI21_X1  g609(.A(new_n807), .B1(new_n810), .B2(new_n806), .ZN(G1340gat));
  INV_X1    g610(.A(G120gat), .ZN(new_n812));
  NAND3_X1  g611(.A1(new_n809), .A2(new_n812), .A3(new_n617), .ZN(new_n813));
  INV_X1    g612(.A(KEYINPUT117), .ZN(new_n814));
  OAI21_X1  g613(.A(G120gat), .B1(new_n805), .B2(new_n703), .ZN(new_n815));
  AND3_X1   g614(.A1(new_n813), .A2(new_n814), .A3(new_n815), .ZN(new_n816));
  AOI21_X1  g615(.A(new_n814), .B1(new_n813), .B2(new_n815), .ZN(new_n817));
  NOR2_X1   g616(.A1(new_n816), .A2(new_n817), .ZN(G1341gat));
  NAND3_X1  g617(.A1(new_n809), .A2(new_n279), .A3(new_n663), .ZN(new_n819));
  OAI21_X1  g618(.A(G127gat), .B1(new_n805), .B2(new_n662), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n819), .A2(new_n820), .ZN(G1342gat));
  NOR2_X1   g620(.A1(new_n445), .A2(new_n584), .ZN(new_n822));
  INV_X1    g621(.A(new_n822), .ZN(new_n823));
  NOR3_X1   g622(.A1(new_n808), .A2(G134gat), .A3(new_n823), .ZN(new_n824));
  INV_X1    g623(.A(KEYINPUT56), .ZN(new_n825));
  OR2_X1    g624(.A1(new_n824), .A2(new_n825), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n824), .A2(new_n825), .ZN(new_n827));
  INV_X1    g626(.A(KEYINPUT118), .ZN(new_n828));
  NAND3_X1  g627(.A1(new_n804), .A2(new_n447), .A3(new_n583), .ZN(new_n829));
  AOI21_X1  g628(.A(new_n828), .B1(new_n829), .B2(G134gat), .ZN(new_n830));
  NAND3_X1  g629(.A1(new_n829), .A2(new_n828), .A3(G134gat), .ZN(new_n831));
  INV_X1    g630(.A(new_n831), .ZN(new_n832));
  OAI211_X1 g631(.A(new_n826), .B(new_n827), .C1(new_n830), .C2(new_n832), .ZN(G1343gat));
  INV_X1    g632(.A(G141gat), .ZN(new_n834));
  NAND2_X1  g633(.A1(new_n631), .A2(new_n674), .ZN(new_n835));
  NOR2_X1   g634(.A1(new_n835), .A2(new_n445), .ZN(new_n836));
  INV_X1    g635(.A(new_n836), .ZN(new_n837));
  OAI21_X1  g636(.A(new_n662), .B1(new_n789), .B2(new_n792), .ZN(new_n838));
  AOI21_X1  g637(.A(new_n436), .B1(new_n838), .B2(new_n802), .ZN(new_n839));
  INV_X1    g638(.A(new_n839), .ZN(new_n840));
  INV_X1    g639(.A(KEYINPUT57), .ZN(new_n841));
  NOR2_X1   g640(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  AOI21_X1  g641(.A(new_n436), .B1(new_n800), .B2(new_n802), .ZN(new_n843));
  XNOR2_X1  g642(.A(KEYINPUT119), .B(KEYINPUT57), .ZN(new_n844));
  INV_X1    g643(.A(new_n844), .ZN(new_n845));
  NOR2_X1   g644(.A1(new_n843), .A2(new_n845), .ZN(new_n846));
  AOI21_X1  g645(.A(new_n842), .B1(new_n846), .B2(KEYINPUT120), .ZN(new_n847));
  INV_X1    g646(.A(KEYINPUT120), .ZN(new_n848));
  OAI21_X1  g647(.A(new_n848), .B1(new_n843), .B2(new_n845), .ZN(new_n849));
  AOI21_X1  g648(.A(new_n837), .B1(new_n847), .B2(new_n849), .ZN(new_n850));
  AOI21_X1  g649(.A(new_n834), .B1(new_n850), .B2(new_n665), .ZN(new_n851));
  NAND2_X1  g650(.A1(new_n800), .A2(new_n802), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n852), .A2(new_n448), .ZN(new_n853));
  NOR3_X1   g652(.A1(new_n853), .A2(new_n445), .A3(new_n835), .ZN(new_n854));
  NAND3_X1  g653(.A1(new_n854), .A2(new_n834), .A3(new_n665), .ZN(new_n855));
  NAND2_X1  g654(.A1(new_n855), .A2(KEYINPUT121), .ZN(new_n856));
  OAI21_X1  g655(.A(KEYINPUT58), .B1(new_n851), .B2(new_n856), .ZN(new_n857));
  NAND3_X1  g656(.A1(new_n853), .A2(KEYINPUT120), .A3(new_n844), .ZN(new_n858));
  OAI21_X1  g657(.A(new_n858), .B1(new_n841), .B2(new_n840), .ZN(new_n859));
  INV_X1    g658(.A(new_n849), .ZN(new_n860));
  OAI211_X1 g659(.A(new_n665), .B(new_n836), .C1(new_n859), .C2(new_n860), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n861), .A2(G141gat), .ZN(new_n862));
  INV_X1    g661(.A(KEYINPUT58), .ZN(new_n863));
  INV_X1    g662(.A(new_n856), .ZN(new_n864));
  NAND3_X1  g663(.A1(new_n862), .A2(new_n863), .A3(new_n864), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n857), .A2(new_n865), .ZN(G1344gat));
  INV_X1    g665(.A(G148gat), .ZN(new_n867));
  NAND3_X1  g666(.A1(new_n854), .A2(new_n867), .A3(new_n617), .ZN(new_n868));
  AOI211_X1 g667(.A(KEYINPUT59), .B(new_n867), .C1(new_n850), .C2(new_n617), .ZN(new_n869));
  INV_X1    g668(.A(KEYINPUT59), .ZN(new_n870));
  INV_X1    g669(.A(KEYINPUT122), .ZN(new_n871));
  OAI21_X1  g670(.A(new_n871), .B1(new_n839), .B2(KEYINPUT57), .ZN(new_n872));
  OAI21_X1  g671(.A(new_n795), .B1(new_n798), .B2(new_n583), .ZN(new_n873));
  AOI21_X1  g672(.A(new_n801), .B1(new_n873), .B2(new_n662), .ZN(new_n874));
  OAI211_X1 g673(.A(KEYINPUT122), .B(new_n841), .C1(new_n874), .C2(new_n436), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n872), .A2(new_n875), .ZN(new_n876));
  AOI211_X1 g675(.A(new_n436), .B(new_n844), .C1(new_n800), .C2(new_n802), .ZN(new_n877));
  OR2_X1    g676(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  NAND3_X1  g677(.A1(new_n878), .A2(new_n617), .A3(new_n836), .ZN(new_n879));
  AOI21_X1  g678(.A(new_n870), .B1(new_n879), .B2(G148gat), .ZN(new_n880));
  OAI21_X1  g679(.A(new_n868), .B1(new_n869), .B2(new_n880), .ZN(G1345gat));
  AOI21_X1  g680(.A(new_n265), .B1(new_n850), .B2(new_n663), .ZN(new_n882));
  AND3_X1   g681(.A1(new_n854), .A2(new_n265), .A3(new_n663), .ZN(new_n883));
  OR2_X1    g682(.A1(new_n882), .A2(new_n883), .ZN(G1346gat));
  AOI21_X1  g683(.A(new_n266), .B1(new_n850), .B2(new_n583), .ZN(new_n885));
  NOR4_X1   g684(.A1(new_n853), .A2(G162gat), .A3(new_n823), .A4(new_n835), .ZN(new_n886));
  OR2_X1    g685(.A1(new_n885), .A2(new_n886), .ZN(G1347gat));
  NAND2_X1  g686(.A1(new_n330), .A2(new_n445), .ZN(new_n888));
  NOR2_X1   g687(.A1(new_n888), .A2(new_n446), .ZN(new_n889));
  NAND2_X1  g688(.A1(new_n803), .A2(new_n889), .ZN(new_n890));
  INV_X1    g689(.A(G169gat), .ZN(new_n891));
  NOR3_X1   g690(.A1(new_n890), .A2(new_n891), .A3(new_n255), .ZN(new_n892));
  AOI21_X1  g691(.A(new_n674), .B1(new_n800), .B2(new_n802), .ZN(new_n893));
  AND4_X1   g692(.A1(new_n445), .A2(new_n893), .A3(new_n436), .A4(new_n644), .ZN(new_n894));
  NAND2_X1  g693(.A1(new_n894), .A2(new_n665), .ZN(new_n895));
  AOI21_X1  g694(.A(new_n892), .B1(new_n895), .B2(new_n891), .ZN(G1348gat));
  INV_X1    g695(.A(G176gat), .ZN(new_n897));
  NAND3_X1  g696(.A1(new_n894), .A2(new_n897), .A3(new_n617), .ZN(new_n898));
  OAI21_X1  g697(.A(G176gat), .B1(new_n890), .B2(new_n703), .ZN(new_n899));
  NAND2_X1  g698(.A1(new_n898), .A2(new_n899), .ZN(G1349gat));
  NAND3_X1  g699(.A1(new_n894), .A2(new_n351), .A3(new_n663), .ZN(new_n901));
  OAI21_X1  g700(.A(G183gat), .B1(new_n890), .B2(new_n662), .ZN(new_n902));
  NAND2_X1  g701(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  XNOR2_X1  g702(.A(new_n903), .B(KEYINPUT60), .ZN(G1350gat));
  NAND3_X1  g703(.A1(new_n894), .A2(new_n352), .A3(new_n583), .ZN(new_n905));
  NAND3_X1  g704(.A1(new_n803), .A2(new_n583), .A3(new_n889), .ZN(new_n906));
  INV_X1    g705(.A(KEYINPUT61), .ZN(new_n907));
  AND3_X1   g706(.A1(new_n906), .A2(new_n907), .A3(G190gat), .ZN(new_n908));
  AOI21_X1  g707(.A(new_n907), .B1(new_n906), .B2(G190gat), .ZN(new_n909));
  OAI21_X1  g708(.A(new_n905), .B1(new_n908), .B2(new_n909), .ZN(new_n910));
  XNOR2_X1  g709(.A(new_n910), .B(KEYINPUT123), .ZN(G1351gat));
  NAND3_X1  g710(.A1(new_n631), .A2(new_n445), .A3(new_n448), .ZN(new_n912));
  XNOR2_X1  g711(.A(new_n912), .B(KEYINPUT124), .ZN(new_n913));
  AND2_X1   g712(.A1(new_n913), .A2(new_n893), .ZN(new_n914));
  AOI21_X1  g713(.A(G197gat), .B1(new_n914), .B2(new_n665), .ZN(new_n915));
  NOR2_X1   g714(.A1(new_n630), .A2(new_n888), .ZN(new_n916));
  AND2_X1   g715(.A1(new_n878), .A2(new_n916), .ZN(new_n917));
  AND2_X1   g716(.A1(new_n665), .A2(G197gat), .ZN(new_n918));
  AOI21_X1  g717(.A(new_n915), .B1(new_n917), .B2(new_n918), .ZN(G1352gat));
  NAND2_X1  g718(.A1(new_n917), .A2(new_n617), .ZN(new_n920));
  NAND2_X1  g719(.A1(new_n920), .A2(G204gat), .ZN(new_n921));
  INV_X1    g720(.A(G204gat), .ZN(new_n922));
  NAND3_X1  g721(.A1(new_n914), .A2(new_n922), .A3(new_n617), .ZN(new_n923));
  AND2_X1   g722(.A1(KEYINPUT125), .A2(KEYINPUT62), .ZN(new_n924));
  NOR2_X1   g723(.A1(KEYINPUT125), .A2(KEYINPUT62), .ZN(new_n925));
  OAI21_X1  g724(.A(new_n923), .B1(new_n924), .B2(new_n925), .ZN(new_n926));
  OAI211_X1 g725(.A(new_n921), .B(new_n926), .C1(new_n924), .C2(new_n923), .ZN(G1353gat));
  NAND3_X1  g726(.A1(new_n914), .A2(new_n366), .A3(new_n663), .ZN(new_n928));
  OAI211_X1 g727(.A(new_n663), .B(new_n916), .C1(new_n876), .C2(new_n877), .ZN(new_n929));
  AND3_X1   g728(.A1(new_n929), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n930));
  AOI21_X1  g729(.A(KEYINPUT63), .B1(new_n929), .B2(G211gat), .ZN(new_n931));
  OAI21_X1  g730(.A(new_n928), .B1(new_n930), .B2(new_n931), .ZN(new_n932));
  NAND2_X1  g731(.A1(new_n932), .A2(KEYINPUT126), .ZN(new_n933));
  INV_X1    g732(.A(KEYINPUT126), .ZN(new_n934));
  OAI211_X1 g733(.A(new_n934), .B(new_n928), .C1(new_n930), .C2(new_n931), .ZN(new_n935));
  NAND2_X1  g734(.A1(new_n933), .A2(new_n935), .ZN(G1354gat));
  NAND3_X1  g735(.A1(new_n914), .A2(new_n367), .A3(new_n583), .ZN(new_n937));
  OAI211_X1 g736(.A(new_n583), .B(new_n916), .C1(new_n876), .C2(new_n877), .ZN(new_n938));
  NAND2_X1  g737(.A1(new_n938), .A2(G218gat), .ZN(new_n939));
  NAND2_X1  g738(.A1(new_n937), .A2(new_n939), .ZN(new_n940));
  XNOR2_X1  g739(.A(new_n940), .B(KEYINPUT127), .ZN(G1355gat));
endmodule


