//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 1 1 0 0 1 0 0 1 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 0 0 0 0 0 0 0 1 0 0 0 1 1 1 0 0 0 1 1 0 0 0 0 1 1 1 0 1 0 0 1 0 0 0 0 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:17:44 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n768, new_n769, new_n770,
    new_n772, new_n773, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n799, new_n800, new_n801,
    new_n802, new_n803, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n814, new_n815, new_n816, new_n817,
    new_n818, new_n819, new_n820, new_n821, new_n823, new_n824, new_n825,
    new_n826, new_n828, new_n829, new_n830, new_n831, new_n832, new_n834,
    new_n835, new_n836, new_n837, new_n839, new_n841, new_n842, new_n843,
    new_n844, new_n845, new_n846, new_n847, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n867, new_n868, new_n869, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n912, new_n913, new_n914, new_n915, new_n916, new_n917,
    new_n918, new_n919, new_n920, new_n921, new_n922, new_n923, new_n924,
    new_n926, new_n927, new_n929, new_n930, new_n932, new_n933, new_n934,
    new_n935, new_n937, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n951, new_n952, new_n953, new_n954, new_n955, new_n956,
    new_n957, new_n958, new_n959, new_n960, new_n961, new_n962, new_n963,
    new_n964, new_n965, new_n966, new_n967, new_n968, new_n969, new_n971,
    new_n972, new_n973, new_n974, new_n975, new_n976, new_n977, new_n978,
    new_n979, new_n980, new_n981, new_n982, new_n983, new_n984, new_n985,
    new_n986, new_n987, new_n988, new_n989, new_n990, new_n992, new_n993,
    new_n994, new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1012, new_n1013, new_n1015, new_n1016,
    new_n1017, new_n1018, new_n1020, new_n1021, new_n1022, new_n1023,
    new_n1025, new_n1026, new_n1027, new_n1028, new_n1029, new_n1030,
    new_n1031, new_n1032, new_n1034, new_n1035, new_n1036, new_n1037,
    new_n1038, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1050, new_n1051,
    new_n1052;
  NAND2_X1  g000(.A1(KEYINPUT97), .A2(G57gat), .ZN(new_n202));
  XNOR2_X1  g001(.A(new_n202), .B(G64gat), .ZN(new_n203));
  NAND2_X1  g002(.A1(G71gat), .A2(G78gat), .ZN(new_n204));
  OR2_X1    g003(.A1(G71gat), .A2(G78gat), .ZN(new_n205));
  INV_X1    g004(.A(KEYINPUT9), .ZN(new_n206));
  OAI21_X1  g005(.A(new_n204), .B1(new_n205), .B2(new_n206), .ZN(new_n207));
  AND2_X1   g006(.A1(new_n203), .A2(new_n207), .ZN(new_n208));
  OAI21_X1  g007(.A(KEYINPUT9), .B1(G57gat), .B2(G64gat), .ZN(new_n209));
  AND2_X1   g008(.A1(G57gat), .A2(G64gat), .ZN(new_n210));
  OR2_X1    g009(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  AND2_X1   g010(.A1(new_n205), .A2(new_n204), .ZN(new_n212));
  AND2_X1   g011(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  OAI21_X1  g012(.A(KEYINPUT98), .B1(new_n208), .B2(new_n213), .ZN(new_n214));
  AOI22_X1  g013(.A1(new_n207), .A2(new_n203), .B1(new_n211), .B2(new_n212), .ZN(new_n215));
  INV_X1    g014(.A(KEYINPUT98), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  NAND2_X1  g016(.A1(new_n214), .A2(new_n217), .ZN(new_n218));
  NOR2_X1   g017(.A1(new_n218), .A2(KEYINPUT21), .ZN(new_n219));
  NAND2_X1  g018(.A1(G231gat), .A2(G233gat), .ZN(new_n220));
  XNOR2_X1  g019(.A(new_n219), .B(new_n220), .ZN(new_n221));
  XNOR2_X1  g020(.A(G127gat), .B(G155gat), .ZN(new_n222));
  XNOR2_X1  g021(.A(new_n222), .B(KEYINPUT99), .ZN(new_n223));
  XNOR2_X1  g022(.A(new_n221), .B(new_n223), .ZN(new_n224));
  XOR2_X1   g023(.A(G183gat), .B(G211gat), .Z(new_n225));
  XNOR2_X1  g024(.A(new_n224), .B(new_n225), .ZN(new_n226));
  INV_X1    g025(.A(G1gat), .ZN(new_n227));
  INV_X1    g026(.A(G15gat), .ZN(new_n228));
  NOR2_X1   g027(.A1(new_n228), .A2(G22gat), .ZN(new_n229));
  INV_X1    g028(.A(G22gat), .ZN(new_n230));
  NOR2_X1   g029(.A1(new_n230), .A2(G15gat), .ZN(new_n231));
  OAI21_X1  g030(.A(new_n227), .B1(new_n229), .B2(new_n231), .ZN(new_n232));
  XNOR2_X1  g031(.A(KEYINPUT93), .B(G8gat), .ZN(new_n233));
  AND2_X1   g032(.A1(new_n232), .A2(new_n233), .ZN(new_n234));
  XNOR2_X1  g033(.A(G15gat), .B(G22gat), .ZN(new_n235));
  INV_X1    g034(.A(KEYINPUT16), .ZN(new_n236));
  OAI21_X1  g035(.A(new_n235), .B1(new_n236), .B2(G1gat), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n237), .A2(KEYINPUT92), .ZN(new_n238));
  INV_X1    g037(.A(KEYINPUT92), .ZN(new_n239));
  OAI211_X1 g038(.A(new_n235), .B(new_n239), .C1(new_n236), .C2(G1gat), .ZN(new_n240));
  NAND3_X1  g039(.A1(new_n234), .A2(new_n238), .A3(new_n240), .ZN(new_n241));
  INV_X1    g040(.A(KEYINPUT94), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n241), .A2(new_n242), .ZN(new_n243));
  NAND4_X1  g042(.A1(new_n234), .A2(new_n238), .A3(KEYINPUT94), .A4(new_n240), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n243), .A2(new_n244), .ZN(new_n245));
  INV_X1    g044(.A(G8gat), .ZN(new_n246));
  AOI21_X1  g045(.A(new_n246), .B1(new_n237), .B2(new_n232), .ZN(new_n247));
  INV_X1    g046(.A(new_n247), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n245), .A2(new_n248), .ZN(new_n249));
  AOI21_X1  g048(.A(new_n249), .B1(KEYINPUT21), .B2(new_n218), .ZN(new_n250));
  XNOR2_X1  g049(.A(new_n250), .B(KEYINPUT100), .ZN(new_n251));
  XOR2_X1   g050(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n252));
  XNOR2_X1  g051(.A(new_n251), .B(new_n252), .ZN(new_n253));
  XNOR2_X1  g052(.A(new_n226), .B(new_n253), .ZN(new_n254));
  NAND2_X1  g053(.A1(G230gat), .A2(G233gat), .ZN(new_n255));
  XNOR2_X1  g054(.A(new_n255), .B(KEYINPUT105), .ZN(new_n256));
  INV_X1    g055(.A(KEYINPUT10), .ZN(new_n257));
  NAND2_X1  g056(.A1(G85gat), .A2(G92gat), .ZN(new_n258));
  XNOR2_X1  g057(.A(new_n258), .B(KEYINPUT7), .ZN(new_n259));
  NAND2_X1  g058(.A1(G99gat), .A2(G106gat), .ZN(new_n260));
  INV_X1    g059(.A(G85gat), .ZN(new_n261));
  INV_X1    g060(.A(G92gat), .ZN(new_n262));
  AOI22_X1  g061(.A1(KEYINPUT8), .A2(new_n260), .B1(new_n261), .B2(new_n262), .ZN(new_n263));
  NAND2_X1  g062(.A1(new_n259), .A2(new_n263), .ZN(new_n264));
  XOR2_X1   g063(.A(G99gat), .B(G106gat), .Z(new_n265));
  NAND2_X1  g064(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  INV_X1    g065(.A(new_n265), .ZN(new_n267));
  NAND3_X1  g066(.A1(new_n267), .A2(new_n259), .A3(new_n263), .ZN(new_n268));
  NAND3_X1  g067(.A1(new_n266), .A2(new_n215), .A3(new_n268), .ZN(new_n269));
  INV_X1    g068(.A(KEYINPUT104), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  NAND4_X1  g070(.A1(new_n266), .A2(new_n215), .A3(KEYINPUT104), .A4(new_n268), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n266), .A2(new_n268), .ZN(new_n274));
  NAND3_X1  g073(.A1(new_n214), .A2(new_n274), .A3(new_n217), .ZN(new_n275));
  AND2_X1   g074(.A1(new_n275), .A2(KEYINPUT103), .ZN(new_n276));
  INV_X1    g075(.A(KEYINPUT103), .ZN(new_n277));
  NAND4_X1  g076(.A1(new_n214), .A2(new_n274), .A3(new_n217), .A4(new_n277), .ZN(new_n278));
  INV_X1    g077(.A(new_n278), .ZN(new_n279));
  OAI211_X1 g078(.A(new_n257), .B(new_n273), .C1(new_n276), .C2(new_n279), .ZN(new_n280));
  INV_X1    g079(.A(new_n274), .ZN(new_n281));
  NAND3_X1  g080(.A1(new_n218), .A2(KEYINPUT10), .A3(new_n281), .ZN(new_n282));
  AOI21_X1  g081(.A(new_n256), .B1(new_n280), .B2(new_n282), .ZN(new_n283));
  INV_X1    g082(.A(new_n256), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n275), .A2(KEYINPUT103), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n285), .A2(new_n278), .ZN(new_n286));
  AOI21_X1  g085(.A(new_n284), .B1(new_n286), .B2(new_n273), .ZN(new_n287));
  XOR2_X1   g086(.A(G120gat), .B(G148gat), .Z(new_n288));
  XNOR2_X1  g087(.A(new_n288), .B(KEYINPUT106), .ZN(new_n289));
  XNOR2_X1  g088(.A(G176gat), .B(G204gat), .ZN(new_n290));
  XOR2_X1   g089(.A(new_n289), .B(new_n290), .Z(new_n291));
  INV_X1    g090(.A(new_n291), .ZN(new_n292));
  NOR3_X1   g091(.A1(new_n283), .A2(new_n287), .A3(new_n292), .ZN(new_n293));
  INV_X1    g092(.A(new_n293), .ZN(new_n294));
  OAI21_X1  g093(.A(new_n292), .B1(new_n283), .B2(new_n287), .ZN(new_n295));
  NAND2_X1  g094(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  XOR2_X1   g095(.A(G43gat), .B(G50gat), .Z(new_n297));
  INV_X1    g096(.A(G36gat), .ZN(new_n298));
  AND2_X1   g097(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n299));
  NOR2_X1   g098(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n300));
  OAI21_X1  g099(.A(new_n298), .B1(new_n299), .B2(new_n300), .ZN(new_n301));
  INV_X1    g100(.A(G29gat), .ZN(new_n302));
  NAND3_X1  g101(.A1(new_n302), .A2(KEYINPUT14), .A3(G36gat), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n301), .A2(new_n303), .ZN(new_n304));
  AOI21_X1  g103(.A(new_n297), .B1(new_n304), .B2(KEYINPUT15), .ZN(new_n305));
  OAI21_X1  g104(.A(new_n305), .B1(KEYINPUT15), .B2(new_n304), .ZN(new_n306));
  NAND3_X1  g105(.A1(new_n304), .A2(KEYINPUT15), .A3(new_n297), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n306), .A2(new_n307), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n308), .A2(KEYINPUT17), .ZN(new_n309));
  INV_X1    g108(.A(KEYINPUT17), .ZN(new_n310));
  NAND3_X1  g109(.A1(new_n306), .A2(new_n310), .A3(new_n307), .ZN(new_n311));
  AOI21_X1  g110(.A(new_n281), .B1(new_n309), .B2(new_n311), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n308), .A2(new_n281), .ZN(new_n313));
  INV_X1    g112(.A(KEYINPUT41), .ZN(new_n314));
  NAND2_X1  g113(.A1(G232gat), .A2(G233gat), .ZN(new_n315));
  OAI21_X1  g114(.A(new_n313), .B1(new_n314), .B2(new_n315), .ZN(new_n316));
  NOR2_X1   g115(.A1(new_n312), .A2(new_n316), .ZN(new_n317));
  XNOR2_X1  g116(.A(G190gat), .B(G218gat), .ZN(new_n318));
  INV_X1    g117(.A(new_n318), .ZN(new_n319));
  INV_X1    g118(.A(KEYINPUT102), .ZN(new_n320));
  XNOR2_X1  g119(.A(G134gat), .B(G162gat), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n315), .A2(new_n314), .ZN(new_n322));
  XNOR2_X1  g121(.A(new_n321), .B(new_n322), .ZN(new_n323));
  AOI22_X1  g122(.A1(new_n317), .A2(new_n319), .B1(new_n320), .B2(new_n323), .ZN(new_n324));
  INV_X1    g123(.A(KEYINPUT101), .ZN(new_n325));
  OAI21_X1  g124(.A(new_n325), .B1(new_n317), .B2(new_n319), .ZN(new_n326));
  OAI211_X1 g125(.A(KEYINPUT101), .B(new_n318), .C1(new_n312), .C2(new_n316), .ZN(new_n327));
  NAND3_X1  g126(.A1(new_n324), .A2(new_n326), .A3(new_n327), .ZN(new_n328));
  NOR2_X1   g127(.A1(new_n323), .A2(new_n320), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n328), .A2(new_n329), .ZN(new_n330));
  INV_X1    g129(.A(new_n329), .ZN(new_n331));
  NAND4_X1  g130(.A1(new_n324), .A2(new_n326), .A3(new_n331), .A4(new_n327), .ZN(new_n332));
  AND2_X1   g131(.A1(new_n330), .A2(new_n332), .ZN(new_n333));
  NOR3_X1   g132(.A1(new_n254), .A2(new_n296), .A3(new_n333), .ZN(new_n334));
  INV_X1    g133(.A(new_n334), .ZN(new_n335));
  INV_X1    g134(.A(G169gat), .ZN(new_n336));
  INV_X1    g135(.A(G176gat), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n336), .A2(new_n337), .ZN(new_n338));
  INV_X1    g137(.A(KEYINPUT26), .ZN(new_n339));
  NAND2_X1  g138(.A1(G169gat), .A2(G176gat), .ZN(new_n340));
  NAND3_X1  g139(.A1(new_n338), .A2(new_n339), .A3(new_n340), .ZN(new_n341));
  NOR2_X1   g140(.A1(G169gat), .A2(G176gat), .ZN(new_n342));
  AOI22_X1  g141(.A1(new_n342), .A2(KEYINPUT26), .B1(G183gat), .B2(G190gat), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n341), .A2(new_n343), .ZN(new_n344));
  XOR2_X1   g143(.A(KEYINPUT27), .B(G183gat), .Z(new_n345));
  INV_X1    g144(.A(G190gat), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n346), .A2(KEYINPUT28), .ZN(new_n347));
  OR2_X1    g146(.A1(new_n345), .A2(new_n347), .ZN(new_n348));
  INV_X1    g147(.A(KEYINPUT27), .ZN(new_n349));
  NAND3_X1  g148(.A1(new_n349), .A2(KEYINPUT67), .A3(G183gat), .ZN(new_n350));
  AND2_X1   g149(.A1(KEYINPUT67), .A2(G183gat), .ZN(new_n351));
  OAI211_X1 g150(.A(new_n346), .B(new_n350), .C1(new_n351), .C2(new_n349), .ZN(new_n352));
  INV_X1    g151(.A(KEYINPUT28), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n352), .A2(new_n353), .ZN(new_n354));
  AOI21_X1  g153(.A(new_n344), .B1(new_n348), .B2(new_n354), .ZN(new_n355));
  INV_X1    g154(.A(new_n355), .ZN(new_n356));
  INV_X1    g155(.A(KEYINPUT23), .ZN(new_n357));
  NOR2_X1   g156(.A1(new_n357), .A2(G176gat), .ZN(new_n358));
  INV_X1    g157(.A(KEYINPUT65), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n359), .A2(new_n336), .ZN(new_n360));
  NAND2_X1  g159(.A1(KEYINPUT65), .A2(G169gat), .ZN(new_n361));
  NAND3_X1  g160(.A1(new_n358), .A2(new_n360), .A3(new_n361), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n340), .A2(KEYINPUT23), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n363), .A2(new_n338), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n362), .A2(new_n364), .ZN(new_n365));
  INV_X1    g164(.A(KEYINPUT24), .ZN(new_n366));
  NAND3_X1  g165(.A1(new_n366), .A2(G183gat), .A3(G190gat), .ZN(new_n367));
  XNOR2_X1  g166(.A(G183gat), .B(G190gat), .ZN(new_n368));
  OAI21_X1  g167(.A(new_n367), .B1(new_n368), .B2(new_n366), .ZN(new_n369));
  AOI21_X1  g168(.A(new_n365), .B1(KEYINPUT64), .B2(new_n369), .ZN(new_n370));
  INV_X1    g169(.A(KEYINPUT64), .ZN(new_n371));
  OAI211_X1 g170(.A(new_n371), .B(new_n367), .C1(new_n368), .C2(new_n366), .ZN(new_n372));
  AOI21_X1  g171(.A(KEYINPUT25), .B1(new_n370), .B2(new_n372), .ZN(new_n373));
  INV_X1    g172(.A(KEYINPUT66), .ZN(new_n374));
  NAND3_X1  g173(.A1(new_n336), .A2(new_n337), .A3(KEYINPUT23), .ZN(new_n375));
  AOI21_X1  g174(.A(new_n357), .B1(G169gat), .B2(G176gat), .ZN(new_n376));
  OAI211_X1 g175(.A(KEYINPUT25), .B(new_n375), .C1(new_n376), .C2(new_n342), .ZN(new_n377));
  OAI21_X1  g176(.A(new_n374), .B1(new_n369), .B2(new_n377), .ZN(new_n378));
  AOI21_X1  g177(.A(new_n342), .B1(KEYINPUT23), .B2(new_n340), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n375), .A2(KEYINPUT25), .ZN(new_n380));
  NOR2_X1   g179(.A1(new_n379), .A2(new_n380), .ZN(new_n381));
  AND3_X1   g180(.A1(new_n366), .A2(G183gat), .A3(G190gat), .ZN(new_n382));
  INV_X1    g181(.A(G183gat), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n383), .A2(G190gat), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n346), .A2(G183gat), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n384), .A2(new_n385), .ZN(new_n386));
  AOI21_X1  g185(.A(new_n382), .B1(new_n386), .B2(KEYINPUT24), .ZN(new_n387));
  NAND3_X1  g186(.A1(new_n381), .A2(KEYINPUT66), .A3(new_n387), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n378), .A2(new_n388), .ZN(new_n389));
  OAI21_X1  g188(.A(new_n356), .B1(new_n373), .B2(new_n389), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n390), .A2(KEYINPUT73), .ZN(new_n391));
  NAND2_X1  g190(.A1(G226gat), .A2(G233gat), .ZN(new_n392));
  INV_X1    g191(.A(new_n392), .ZN(new_n393));
  NOR3_X1   g192(.A1(new_n369), .A2(new_n377), .A3(new_n374), .ZN(new_n394));
  AOI21_X1  g193(.A(KEYINPUT66), .B1(new_n381), .B2(new_n387), .ZN(new_n395));
  NOR2_X1   g194(.A1(new_n394), .A2(new_n395), .ZN(new_n396));
  AOI21_X1  g195(.A(new_n366), .B1(new_n384), .B2(new_n385), .ZN(new_n397));
  OAI21_X1  g196(.A(KEYINPUT64), .B1(new_n397), .B2(new_n382), .ZN(new_n398));
  INV_X1    g197(.A(new_n361), .ZN(new_n399));
  NOR2_X1   g198(.A1(KEYINPUT65), .A2(G169gat), .ZN(new_n400));
  NOR2_X1   g199(.A1(new_n399), .A2(new_n400), .ZN(new_n401));
  AOI22_X1  g200(.A1(new_n401), .A2(new_n358), .B1(new_n338), .B2(new_n363), .ZN(new_n402));
  NAND3_X1  g201(.A1(new_n398), .A2(new_n402), .A3(new_n372), .ZN(new_n403));
  INV_X1    g202(.A(KEYINPUT25), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n403), .A2(new_n404), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n396), .A2(new_n405), .ZN(new_n406));
  INV_X1    g205(.A(KEYINPUT73), .ZN(new_n407));
  NAND3_X1  g206(.A1(new_n406), .A2(new_n407), .A3(new_n356), .ZN(new_n408));
  NAND3_X1  g207(.A1(new_n391), .A2(new_n393), .A3(new_n408), .ZN(new_n409));
  INV_X1    g208(.A(KEYINPUT29), .ZN(new_n410));
  NAND3_X1  g209(.A1(new_n390), .A2(new_n410), .A3(new_n392), .ZN(new_n411));
  AND2_X1   g210(.A1(G211gat), .A2(G218gat), .ZN(new_n412));
  NOR2_X1   g211(.A1(G211gat), .A2(G218gat), .ZN(new_n413));
  NOR2_X1   g212(.A1(new_n412), .A2(new_n413), .ZN(new_n414));
  AND2_X1   g213(.A1(G197gat), .A2(G204gat), .ZN(new_n415));
  NOR2_X1   g214(.A1(G197gat), .A2(G204gat), .ZN(new_n416));
  NOR2_X1   g215(.A1(new_n415), .A2(new_n416), .ZN(new_n417));
  AOI21_X1  g216(.A(KEYINPUT22), .B1(G211gat), .B2(G218gat), .ZN(new_n418));
  OAI21_X1  g217(.A(new_n414), .B1(new_n417), .B2(new_n418), .ZN(new_n419));
  XNOR2_X1  g218(.A(G211gat), .B(G218gat), .ZN(new_n420));
  XNOR2_X1  g219(.A(G197gat), .B(G204gat), .ZN(new_n421));
  INV_X1    g220(.A(new_n418), .ZN(new_n422));
  NAND3_X1  g221(.A1(new_n420), .A2(new_n421), .A3(new_n422), .ZN(new_n423));
  INV_X1    g222(.A(KEYINPUT71), .ZN(new_n424));
  NAND3_X1  g223(.A1(new_n419), .A2(new_n423), .A3(new_n424), .ZN(new_n425));
  OAI211_X1 g224(.A(KEYINPUT71), .B(new_n414), .C1(new_n417), .C2(new_n418), .ZN(new_n426));
  AND3_X1   g225(.A1(new_n425), .A2(KEYINPUT72), .A3(new_n426), .ZN(new_n427));
  AOI21_X1  g226(.A(KEYINPUT72), .B1(new_n425), .B2(new_n426), .ZN(new_n428));
  NOR2_X1   g227(.A1(new_n427), .A2(new_n428), .ZN(new_n429));
  INV_X1    g228(.A(new_n429), .ZN(new_n430));
  NAND3_X1  g229(.A1(new_n409), .A2(new_n411), .A3(new_n430), .ZN(new_n431));
  XNOR2_X1  g230(.A(G8gat), .B(G36gat), .ZN(new_n432));
  XNOR2_X1  g231(.A(G64gat), .B(G92gat), .ZN(new_n433));
  XOR2_X1   g232(.A(new_n432), .B(new_n433), .Z(new_n434));
  NAND2_X1  g233(.A1(new_n391), .A2(new_n408), .ZN(new_n435));
  AOI21_X1  g234(.A(new_n393), .B1(new_n435), .B2(new_n410), .ZN(new_n436));
  AOI21_X1  g235(.A(new_n355), .B1(new_n396), .B2(new_n405), .ZN(new_n437));
  INV_X1    g236(.A(KEYINPUT74), .ZN(new_n438));
  NOR3_X1   g237(.A1(new_n437), .A2(new_n438), .A3(new_n392), .ZN(new_n439));
  AOI21_X1  g238(.A(KEYINPUT74), .B1(new_n390), .B2(new_n393), .ZN(new_n440));
  OAI21_X1  g239(.A(new_n429), .B1(new_n439), .B2(new_n440), .ZN(new_n441));
  OAI211_X1 g240(.A(new_n431), .B(new_n434), .C1(new_n436), .C2(new_n441), .ZN(new_n442));
  INV_X1    g241(.A(KEYINPUT30), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  OAI21_X1  g243(.A(new_n431), .B1(new_n436), .B2(new_n441), .ZN(new_n445));
  INV_X1    g244(.A(new_n434), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  OAI21_X1  g246(.A(new_n438), .B1(new_n437), .B2(new_n392), .ZN(new_n448));
  NAND3_X1  g247(.A1(new_n390), .A2(KEYINPUT74), .A3(new_n393), .ZN(new_n449));
  AOI21_X1  g248(.A(new_n430), .B1(new_n448), .B2(new_n449), .ZN(new_n450));
  AOI21_X1  g249(.A(KEYINPUT29), .B1(new_n391), .B2(new_n408), .ZN(new_n451));
  OAI21_X1  g250(.A(new_n450), .B1(new_n393), .B2(new_n451), .ZN(new_n452));
  NAND4_X1  g251(.A1(new_n452), .A2(KEYINPUT30), .A3(new_n431), .A4(new_n434), .ZN(new_n453));
  NAND3_X1  g252(.A1(new_n444), .A2(new_n447), .A3(new_n453), .ZN(new_n454));
  INV_X1    g253(.A(KEYINPUT82), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  NAND4_X1  g255(.A1(new_n444), .A2(new_n447), .A3(KEYINPUT82), .A4(new_n453), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  XOR2_X1   g257(.A(G15gat), .B(G43gat), .Z(new_n459));
  XNOR2_X1  g258(.A(G71gat), .B(G99gat), .ZN(new_n460));
  XNOR2_X1  g259(.A(new_n459), .B(new_n460), .ZN(new_n461));
  INV_X1    g260(.A(new_n461), .ZN(new_n462));
  INV_X1    g261(.A(G227gat), .ZN(new_n463));
  INV_X1    g262(.A(G233gat), .ZN(new_n464));
  NOR2_X1   g263(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  INV_X1    g264(.A(G134gat), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n466), .A2(G127gat), .ZN(new_n467));
  INV_X1    g266(.A(G127gat), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n468), .A2(G134gat), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n467), .A2(new_n469), .ZN(new_n470));
  XNOR2_X1  g269(.A(G113gat), .B(G120gat), .ZN(new_n471));
  OAI21_X1  g270(.A(new_n470), .B1(new_n471), .B2(KEYINPUT1), .ZN(new_n472));
  INV_X1    g271(.A(G113gat), .ZN(new_n473));
  NAND3_X1  g272(.A1(new_n473), .A2(KEYINPUT68), .A3(G120gat), .ZN(new_n474));
  INV_X1    g273(.A(KEYINPUT1), .ZN(new_n475));
  NAND4_X1  g274(.A1(new_n474), .A2(new_n467), .A3(new_n469), .A4(new_n475), .ZN(new_n476));
  INV_X1    g275(.A(new_n476), .ZN(new_n477));
  INV_X1    g276(.A(KEYINPUT68), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n471), .A2(new_n478), .ZN(new_n479));
  AOI21_X1  g278(.A(KEYINPUT69), .B1(new_n477), .B2(new_n479), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n473), .A2(G120gat), .ZN(new_n481));
  INV_X1    g280(.A(G120gat), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n482), .A2(G113gat), .ZN(new_n483));
  AND3_X1   g282(.A1(new_n481), .A2(new_n483), .A3(new_n478), .ZN(new_n484));
  INV_X1    g283(.A(KEYINPUT69), .ZN(new_n485));
  NOR3_X1   g284(.A1(new_n484), .A2(new_n476), .A3(new_n485), .ZN(new_n486));
  OAI21_X1  g285(.A(new_n472), .B1(new_n480), .B2(new_n486), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n487), .A2(KEYINPUT70), .ZN(new_n488));
  NAND3_X1  g287(.A1(new_n477), .A2(KEYINPUT69), .A3(new_n479), .ZN(new_n489));
  OAI21_X1  g288(.A(new_n485), .B1(new_n484), .B2(new_n476), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  INV_X1    g290(.A(KEYINPUT70), .ZN(new_n492));
  NAND3_X1  g291(.A1(new_n491), .A2(new_n492), .A3(new_n472), .ZN(new_n493));
  NAND4_X1  g292(.A1(new_n406), .A2(new_n488), .A3(new_n493), .A4(new_n356), .ZN(new_n494));
  INV_X1    g293(.A(new_n494), .ZN(new_n495));
  AOI22_X1  g294(.A1(new_n356), .A2(new_n406), .B1(new_n488), .B2(new_n493), .ZN(new_n496));
  OAI21_X1  g295(.A(new_n465), .B1(new_n495), .B2(new_n496), .ZN(new_n497));
  INV_X1    g296(.A(KEYINPUT33), .ZN(new_n498));
  AOI21_X1  g297(.A(new_n462), .B1(new_n497), .B2(new_n498), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n488), .A2(new_n493), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n500), .A2(new_n390), .ZN(new_n501));
  INV_X1    g300(.A(new_n465), .ZN(new_n502));
  NAND3_X1  g301(.A1(new_n501), .A2(new_n502), .A3(new_n494), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n503), .A2(KEYINPUT34), .ZN(new_n504));
  INV_X1    g303(.A(KEYINPUT34), .ZN(new_n505));
  NAND4_X1  g304(.A1(new_n501), .A2(new_n494), .A3(new_n505), .A4(new_n502), .ZN(new_n506));
  NAND2_X1  g305(.A1(new_n504), .A2(new_n506), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n499), .A2(new_n507), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n501), .A2(new_n494), .ZN(new_n509));
  AOI21_X1  g308(.A(KEYINPUT33), .B1(new_n509), .B2(new_n465), .ZN(new_n510));
  OAI211_X1 g309(.A(new_n504), .B(new_n506), .C1(new_n510), .C2(new_n462), .ZN(new_n511));
  AND2_X1   g310(.A1(new_n497), .A2(KEYINPUT32), .ZN(new_n512));
  AND3_X1   g311(.A1(new_n508), .A2(new_n511), .A3(new_n512), .ZN(new_n513));
  NAND2_X1  g312(.A1(G155gat), .A2(G162gat), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n514), .A2(KEYINPUT2), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n515), .A2(KEYINPUT75), .ZN(new_n516));
  XNOR2_X1  g315(.A(G155gat), .B(G162gat), .ZN(new_n517));
  XNOR2_X1  g316(.A(G141gat), .B(G148gat), .ZN(new_n518));
  AND2_X1   g317(.A1(new_n514), .A2(KEYINPUT2), .ZN(new_n519));
  OAI211_X1 g318(.A(new_n516), .B(new_n517), .C1(new_n518), .C2(new_n519), .ZN(new_n520));
  INV_X1    g319(.A(G141gat), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n521), .A2(G148gat), .ZN(new_n522));
  INV_X1    g321(.A(G148gat), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n523), .A2(G141gat), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n522), .A2(new_n524), .ZN(new_n525));
  AND2_X1   g324(.A1(G155gat), .A2(G162gat), .ZN(new_n526));
  NOR2_X1   g325(.A1(G155gat), .A2(G162gat), .ZN(new_n527));
  NOR2_X1   g326(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  OAI211_X1 g327(.A(new_n515), .B(new_n525), .C1(new_n528), .C2(KEYINPUT75), .ZN(new_n529));
  NAND2_X1  g328(.A1(new_n520), .A2(new_n529), .ZN(new_n530));
  XOR2_X1   g329(.A(KEYINPUT76), .B(KEYINPUT3), .Z(new_n531));
  NAND2_X1  g330(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  NAND3_X1  g331(.A1(new_n532), .A2(KEYINPUT80), .A3(new_n410), .ZN(new_n533));
  INV_X1    g332(.A(KEYINPUT80), .ZN(new_n534));
  INV_X1    g333(.A(new_n531), .ZN(new_n535));
  AOI21_X1  g334(.A(new_n535), .B1(new_n520), .B2(new_n529), .ZN(new_n536));
  OAI21_X1  g335(.A(new_n534), .B1(new_n536), .B2(KEYINPUT29), .ZN(new_n537));
  OAI211_X1 g336(.A(new_n533), .B(new_n537), .C1(new_n427), .C2(new_n428), .ZN(new_n538));
  NAND2_X1  g337(.A1(G228gat), .A2(G233gat), .ZN(new_n539));
  INV_X1    g338(.A(KEYINPUT3), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n425), .A2(new_n426), .ZN(new_n541));
  OAI21_X1  g340(.A(new_n540), .B1(new_n541), .B2(KEYINPUT29), .ZN(new_n542));
  INV_X1    g341(.A(new_n530), .ZN(new_n543));
  AOI21_X1  g342(.A(new_n539), .B1(new_n542), .B2(new_n543), .ZN(new_n544));
  NAND2_X1  g343(.A1(new_n538), .A2(new_n544), .ZN(new_n545));
  AOI21_X1  g344(.A(KEYINPUT29), .B1(new_n530), .B2(new_n531), .ZN(new_n546));
  INV_X1    g345(.A(KEYINPUT72), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n541), .A2(new_n547), .ZN(new_n548));
  NAND3_X1  g347(.A1(new_n425), .A2(KEYINPUT72), .A3(new_n426), .ZN(new_n549));
  AOI21_X1  g348(.A(new_n546), .B1(new_n548), .B2(new_n549), .ZN(new_n550));
  NAND3_X1  g349(.A1(new_n419), .A2(new_n423), .A3(KEYINPUT79), .ZN(new_n551));
  INV_X1    g350(.A(KEYINPUT79), .ZN(new_n552));
  NAND4_X1  g351(.A1(new_n420), .A2(new_n421), .A3(new_n552), .A4(new_n422), .ZN(new_n553));
  NAND3_X1  g352(.A1(new_n551), .A2(new_n410), .A3(new_n553), .ZN(new_n554));
  AOI21_X1  g353(.A(new_n530), .B1(new_n554), .B2(new_n531), .ZN(new_n555));
  OAI21_X1  g354(.A(new_n539), .B1(new_n550), .B2(new_n555), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n545), .A2(new_n556), .ZN(new_n557));
  XNOR2_X1  g356(.A(G78gat), .B(G106gat), .ZN(new_n558));
  XNOR2_X1  g357(.A(KEYINPUT31), .B(G50gat), .ZN(new_n559));
  XOR2_X1   g358(.A(new_n558), .B(new_n559), .Z(new_n560));
  INV_X1    g359(.A(new_n560), .ZN(new_n561));
  AOI21_X1  g360(.A(KEYINPUT81), .B1(new_n557), .B2(new_n561), .ZN(new_n562));
  OAI22_X1  g361(.A1(new_n427), .A2(new_n428), .B1(KEYINPUT29), .B2(new_n536), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n554), .A2(new_n531), .ZN(new_n564));
  NAND2_X1  g363(.A1(new_n564), .A2(new_n543), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n563), .A2(new_n565), .ZN(new_n566));
  AOI22_X1  g365(.A1(new_n566), .A2(new_n539), .B1(new_n538), .B2(new_n544), .ZN(new_n567));
  AOI21_X1  g366(.A(new_n230), .B1(new_n567), .B2(new_n560), .ZN(new_n568));
  AND4_X1   g367(.A1(new_n230), .A2(new_n545), .A3(new_n556), .A4(new_n560), .ZN(new_n569));
  OAI21_X1  g368(.A(new_n562), .B1(new_n568), .B2(new_n569), .ZN(new_n570));
  INV_X1    g369(.A(KEYINPUT81), .ZN(new_n571));
  OAI21_X1  g370(.A(new_n571), .B1(new_n567), .B2(new_n560), .ZN(new_n572));
  OAI21_X1  g371(.A(G22gat), .B1(new_n557), .B2(new_n561), .ZN(new_n573));
  NAND3_X1  g372(.A1(new_n567), .A2(new_n230), .A3(new_n560), .ZN(new_n574));
  NAND3_X1  g373(.A1(new_n572), .A2(new_n573), .A3(new_n574), .ZN(new_n575));
  AND2_X1   g374(.A1(new_n570), .A2(new_n575), .ZN(new_n576));
  AOI21_X1  g375(.A(new_n512), .B1(new_n508), .B2(new_n511), .ZN(new_n577));
  NOR3_X1   g376(.A1(new_n513), .A2(new_n576), .A3(new_n577), .ZN(new_n578));
  INV_X1    g377(.A(KEYINPUT35), .ZN(new_n579));
  XOR2_X1   g378(.A(G1gat), .B(G29gat), .Z(new_n580));
  XNOR2_X1  g379(.A(KEYINPUT77), .B(KEYINPUT0), .ZN(new_n581));
  XNOR2_X1  g380(.A(new_n580), .B(new_n581), .ZN(new_n582));
  XNOR2_X1  g381(.A(G57gat), .B(G85gat), .ZN(new_n583));
  XNOR2_X1  g382(.A(new_n582), .B(new_n583), .ZN(new_n584));
  NAND3_X1  g383(.A1(new_n491), .A2(new_n530), .A3(new_n472), .ZN(new_n585));
  INV_X1    g384(.A(new_n585), .ZN(new_n586));
  NOR2_X1   g385(.A1(new_n586), .A2(KEYINPUT4), .ZN(new_n587));
  OAI21_X1  g386(.A(new_n532), .B1(new_n540), .B2(new_n530), .ZN(new_n588));
  INV_X1    g387(.A(new_n487), .ZN(new_n589));
  NOR2_X1   g388(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  NAND2_X1  g389(.A1(G225gat), .A2(G233gat), .ZN(new_n591));
  INV_X1    g390(.A(new_n591), .ZN(new_n592));
  NOR3_X1   g391(.A1(new_n587), .A2(new_n590), .A3(new_n592), .ZN(new_n593));
  NAND4_X1  g392(.A1(new_n488), .A2(KEYINPUT4), .A3(new_n530), .A4(new_n493), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  AOI21_X1  g394(.A(new_n530), .B1(new_n491), .B2(new_n472), .ZN(new_n596));
  OAI21_X1  g395(.A(new_n592), .B1(new_n586), .B2(new_n596), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n597), .A2(KEYINPUT5), .ZN(new_n598));
  INV_X1    g397(.A(new_n598), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n595), .A2(new_n599), .ZN(new_n600));
  INV_X1    g399(.A(KEYINPUT4), .ZN(new_n601));
  NAND4_X1  g400(.A1(new_n488), .A2(new_n601), .A3(new_n530), .A4(new_n493), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n585), .A2(KEYINPUT4), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  NAND2_X1  g403(.A1(new_n604), .A2(KEYINPUT78), .ZN(new_n605));
  INV_X1    g404(.A(KEYINPUT78), .ZN(new_n606));
  NAND3_X1  g405(.A1(new_n602), .A2(new_n606), .A3(new_n603), .ZN(new_n607));
  NOR3_X1   g406(.A1(new_n590), .A2(KEYINPUT5), .A3(new_n592), .ZN(new_n608));
  NAND3_X1  g407(.A1(new_n605), .A2(new_n607), .A3(new_n608), .ZN(new_n609));
  AOI21_X1  g408(.A(new_n584), .B1(new_n600), .B2(new_n609), .ZN(new_n610));
  NAND2_X1  g409(.A1(new_n610), .A2(KEYINPUT6), .ZN(new_n611));
  XOR2_X1   g410(.A(new_n584), .B(KEYINPUT83), .Z(new_n612));
  INV_X1    g411(.A(new_n612), .ZN(new_n613));
  INV_X1    g412(.A(KEYINPUT85), .ZN(new_n614));
  AND3_X1   g413(.A1(new_n602), .A2(new_n606), .A3(new_n603), .ZN(new_n615));
  AOI21_X1  g414(.A(new_n606), .B1(new_n602), .B2(new_n603), .ZN(new_n616));
  OR2_X1    g415(.A1(new_n588), .A2(new_n589), .ZN(new_n617));
  INV_X1    g416(.A(KEYINPUT5), .ZN(new_n618));
  NAND3_X1  g417(.A1(new_n617), .A2(new_n618), .A3(new_n591), .ZN(new_n619));
  NOR3_X1   g418(.A1(new_n615), .A2(new_n616), .A3(new_n619), .ZN(new_n620));
  AOI21_X1  g419(.A(new_n598), .B1(new_n593), .B2(new_n594), .ZN(new_n621));
  OAI21_X1  g420(.A(new_n614), .B1(new_n620), .B2(new_n621), .ZN(new_n622));
  NAND3_X1  g421(.A1(new_n600), .A2(KEYINPUT85), .A3(new_n609), .ZN(new_n623));
  AOI21_X1  g422(.A(new_n613), .B1(new_n622), .B2(new_n623), .ZN(new_n624));
  INV_X1    g423(.A(KEYINPUT6), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n600), .A2(new_n609), .ZN(new_n626));
  INV_X1    g425(.A(new_n584), .ZN(new_n627));
  OAI21_X1  g426(.A(new_n625), .B1(new_n626), .B2(new_n627), .ZN(new_n628));
  OAI21_X1  g427(.A(new_n611), .B1(new_n624), .B2(new_n628), .ZN(new_n629));
  NAND4_X1  g428(.A1(new_n458), .A2(new_n578), .A3(new_n579), .A4(new_n629), .ZN(new_n630));
  INV_X1    g429(.A(KEYINPUT89), .ZN(new_n631));
  NOR2_X1   g430(.A1(new_n513), .A2(new_n577), .ZN(new_n632));
  OAI21_X1  g431(.A(new_n611), .B1(new_n628), .B2(new_n610), .ZN(new_n633));
  INV_X1    g432(.A(new_n576), .ZN(new_n634));
  INV_X1    g433(.A(new_n454), .ZN(new_n635));
  NAND4_X1  g434(.A1(new_n632), .A2(new_n633), .A3(new_n634), .A4(new_n635), .ZN(new_n636));
  AOI22_X1  g435(.A1(new_n630), .A2(new_n631), .B1(KEYINPUT35), .B2(new_n636), .ZN(new_n637));
  NOR4_X1   g436(.A1(new_n513), .A2(new_n576), .A3(new_n577), .A4(KEYINPUT35), .ZN(new_n638));
  NAND4_X1  g437(.A1(new_n638), .A2(KEYINPUT89), .A3(new_n458), .A4(new_n629), .ZN(new_n639));
  INV_X1    g438(.A(KEYINPUT40), .ZN(new_n640));
  NOR2_X1   g439(.A1(new_n615), .A2(new_n616), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n641), .A2(new_n617), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n642), .A2(new_n592), .ZN(new_n643));
  OR2_X1    g442(.A1(new_n586), .A2(new_n596), .ZN(new_n644));
  OAI21_X1  g443(.A(KEYINPUT39), .B1(new_n644), .B2(new_n592), .ZN(new_n645));
  INV_X1    g444(.A(new_n645), .ZN(new_n646));
  AOI21_X1  g445(.A(new_n640), .B1(new_n643), .B2(new_n646), .ZN(new_n647));
  AOI21_X1  g446(.A(new_n591), .B1(new_n641), .B2(new_n617), .ZN(new_n648));
  INV_X1    g447(.A(KEYINPUT39), .ZN(new_n649));
  AOI21_X1  g448(.A(new_n612), .B1(new_n648), .B2(new_n649), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n622), .A2(new_n623), .ZN(new_n651));
  AOI22_X1  g450(.A1(new_n647), .A2(new_n650), .B1(new_n651), .B2(new_n612), .ZN(new_n652));
  XNOR2_X1  g451(.A(KEYINPUT84), .B(KEYINPUT40), .ZN(new_n653));
  OAI21_X1  g452(.A(new_n613), .B1(new_n643), .B2(KEYINPUT39), .ZN(new_n654));
  NOR2_X1   g453(.A1(new_n648), .A2(new_n645), .ZN(new_n655));
  OAI21_X1  g454(.A(new_n653), .B1(new_n654), .B2(new_n655), .ZN(new_n656));
  NAND4_X1  g455(.A1(new_n652), .A2(new_n656), .A3(new_n456), .A4(new_n457), .ZN(new_n657));
  INV_X1    g456(.A(KEYINPUT37), .ZN(new_n658));
  NOR2_X1   g457(.A1(new_n434), .A2(new_n658), .ZN(new_n659));
  AOI21_X1  g458(.A(new_n659), .B1(new_n445), .B2(new_n446), .ZN(new_n660));
  NOR2_X1   g459(.A1(new_n660), .A2(KEYINPUT38), .ZN(new_n661));
  NAND2_X1  g460(.A1(new_n409), .A2(new_n411), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n662), .A2(new_n429), .ZN(new_n663));
  AOI21_X1  g462(.A(new_n407), .B1(new_n406), .B2(new_n356), .ZN(new_n664));
  AOI211_X1 g463(.A(KEYINPUT73), .B(new_n355), .C1(new_n396), .C2(new_n405), .ZN(new_n665));
  OAI21_X1  g464(.A(new_n410), .B1(new_n664), .B2(new_n665), .ZN(new_n666));
  AOI22_X1  g465(.A1(new_n666), .A2(new_n392), .B1(new_n448), .B2(new_n449), .ZN(new_n667));
  OAI211_X1 g466(.A(new_n663), .B(KEYINPUT86), .C1(new_n667), .C2(new_n429), .ZN(new_n668));
  INV_X1    g467(.A(KEYINPUT87), .ZN(new_n669));
  AOI21_X1  g468(.A(new_n430), .B1(new_n409), .B2(new_n411), .ZN(new_n670));
  INV_X1    g469(.A(KEYINPUT86), .ZN(new_n671));
  AOI21_X1  g470(.A(new_n658), .B1(new_n670), .B2(new_n671), .ZN(new_n672));
  AND3_X1   g471(.A1(new_n668), .A2(new_n669), .A3(new_n672), .ZN(new_n673));
  AOI21_X1  g472(.A(new_n669), .B1(new_n668), .B2(new_n672), .ZN(new_n674));
  OAI21_X1  g473(.A(new_n661), .B1(new_n673), .B2(new_n674), .ZN(new_n675));
  NAND2_X1  g474(.A1(new_n651), .A2(new_n612), .ZN(new_n676));
  INV_X1    g475(.A(new_n628), .ZN(new_n677));
  NAND2_X1  g476(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  AND2_X1   g477(.A1(new_n611), .A2(new_n442), .ZN(new_n679));
  NAND3_X1  g478(.A1(new_n675), .A2(new_n678), .A3(new_n679), .ZN(new_n680));
  AOI21_X1  g479(.A(new_n658), .B1(new_n452), .B2(new_n431), .ZN(new_n681));
  OAI211_X1 g480(.A(KEYINPUT88), .B(KEYINPUT38), .C1(new_n660), .C2(new_n681), .ZN(new_n682));
  INV_X1    g481(.A(new_n682), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n445), .A2(KEYINPUT37), .ZN(new_n684));
  AOI21_X1  g483(.A(new_n434), .B1(new_n452), .B2(new_n431), .ZN(new_n685));
  OAI21_X1  g484(.A(new_n684), .B1(new_n685), .B2(new_n659), .ZN(new_n686));
  AOI21_X1  g485(.A(KEYINPUT88), .B1(new_n686), .B2(KEYINPUT38), .ZN(new_n687));
  NOR2_X1   g486(.A1(new_n683), .A2(new_n687), .ZN(new_n688));
  OAI211_X1 g487(.A(new_n634), .B(new_n657), .C1(new_n680), .C2(new_n688), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n632), .A2(KEYINPUT36), .ZN(new_n690));
  INV_X1    g489(.A(KEYINPUT36), .ZN(new_n691));
  OAI21_X1  g490(.A(new_n691), .B1(new_n513), .B2(new_n577), .ZN(new_n692));
  NAND2_X1  g491(.A1(new_n633), .A2(new_n635), .ZN(new_n693));
  AOI22_X1  g492(.A1(new_n690), .A2(new_n692), .B1(new_n693), .B2(new_n576), .ZN(new_n694));
  AOI22_X1  g493(.A1(new_n637), .A2(new_n639), .B1(new_n689), .B2(new_n694), .ZN(new_n695));
  NAND2_X1  g494(.A1(new_n249), .A2(new_n308), .ZN(new_n696));
  AOI21_X1  g495(.A(new_n247), .B1(new_n243), .B2(new_n244), .ZN(new_n697));
  INV_X1    g496(.A(new_n311), .ZN(new_n698));
  AOI21_X1  g497(.A(new_n310), .B1(new_n306), .B2(new_n307), .ZN(new_n699));
  OAI21_X1  g498(.A(new_n697), .B1(new_n698), .B2(new_n699), .ZN(new_n700));
  NAND2_X1  g499(.A1(G229gat), .A2(G233gat), .ZN(new_n701));
  NAND3_X1  g500(.A1(new_n696), .A2(new_n700), .A3(new_n701), .ZN(new_n702));
  INV_X1    g501(.A(KEYINPUT95), .ZN(new_n703));
  NAND2_X1  g502(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n704), .A2(KEYINPUT18), .ZN(new_n705));
  INV_X1    g504(.A(KEYINPUT18), .ZN(new_n706));
  NAND3_X1  g505(.A1(new_n702), .A2(new_n703), .A3(new_n706), .ZN(new_n707));
  XOR2_X1   g506(.A(new_n701), .B(KEYINPUT13), .Z(new_n708));
  INV_X1    g507(.A(new_n696), .ZN(new_n709));
  NOR2_X1   g508(.A1(new_n249), .A2(new_n308), .ZN(new_n710));
  OAI21_X1  g509(.A(new_n708), .B1(new_n709), .B2(new_n710), .ZN(new_n711));
  NAND3_X1  g510(.A1(new_n705), .A2(new_n707), .A3(new_n711), .ZN(new_n712));
  XNOR2_X1  g511(.A(G113gat), .B(G141gat), .ZN(new_n713));
  XNOR2_X1  g512(.A(new_n713), .B(KEYINPUT91), .ZN(new_n714));
  XOR2_X1   g513(.A(G169gat), .B(G197gat), .Z(new_n715));
  XNOR2_X1  g514(.A(new_n714), .B(new_n715), .ZN(new_n716));
  XNOR2_X1  g515(.A(KEYINPUT90), .B(KEYINPUT11), .ZN(new_n717));
  XNOR2_X1  g516(.A(new_n716), .B(new_n717), .ZN(new_n718));
  XNOR2_X1  g517(.A(new_n718), .B(KEYINPUT12), .ZN(new_n719));
  INV_X1    g518(.A(new_n719), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n712), .A2(new_n720), .ZN(new_n721));
  NAND4_X1  g520(.A1(new_n705), .A2(new_n719), .A3(new_n707), .A4(new_n711), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  INV_X1    g522(.A(new_n723), .ZN(new_n724));
  OAI21_X1  g523(.A(KEYINPUT96), .B1(new_n695), .B2(new_n724), .ZN(new_n725));
  INV_X1    g524(.A(KEYINPUT96), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n630), .A2(new_n631), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n636), .A2(KEYINPUT35), .ZN(new_n728));
  AND3_X1   g527(.A1(new_n727), .A2(new_n639), .A3(new_n728), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n690), .A2(new_n692), .ZN(new_n730));
  NAND2_X1  g529(.A1(new_n693), .A2(new_n576), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  AND2_X1   g531(.A1(new_n657), .A2(new_n634), .ZN(new_n733));
  NAND2_X1  g532(.A1(new_n686), .A2(KEYINPUT38), .ZN(new_n734));
  INV_X1    g533(.A(KEYINPUT88), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n736), .A2(new_n682), .ZN(new_n737));
  NAND4_X1  g536(.A1(new_n737), .A2(new_n678), .A3(new_n675), .A4(new_n679), .ZN(new_n738));
  AOI21_X1  g537(.A(new_n732), .B1(new_n733), .B2(new_n738), .ZN(new_n739));
  OAI211_X1 g538(.A(new_n726), .B(new_n723), .C1(new_n729), .C2(new_n739), .ZN(new_n740));
  AOI21_X1  g539(.A(new_n335), .B1(new_n725), .B2(new_n740), .ZN(new_n741));
  INV_X1    g540(.A(new_n633), .ZN(new_n742));
  NAND2_X1  g541(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  XNOR2_X1  g542(.A(new_n743), .B(G1gat), .ZN(G1324gat));
  INV_X1    g543(.A(KEYINPUT42), .ZN(new_n745));
  INV_X1    g544(.A(new_n458), .ZN(new_n746));
  NAND3_X1  g545(.A1(new_n727), .A2(new_n639), .A3(new_n728), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n689), .A2(new_n694), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  AOI21_X1  g548(.A(new_n726), .B1(new_n749), .B2(new_n723), .ZN(new_n750));
  AOI211_X1 g549(.A(KEYINPUT96), .B(new_n724), .C1(new_n747), .C2(new_n748), .ZN(new_n751));
  OAI211_X1 g550(.A(new_n746), .B(new_n334), .C1(new_n750), .C2(new_n751), .ZN(new_n752));
  NAND2_X1  g551(.A1(new_n752), .A2(G8gat), .ZN(new_n753));
  XNOR2_X1  g552(.A(KEYINPUT107), .B(KEYINPUT16), .ZN(new_n754));
  XNOR2_X1  g553(.A(new_n754), .B(new_n246), .ZN(new_n755));
  NAND3_X1  g554(.A1(new_n741), .A2(new_n746), .A3(new_n755), .ZN(new_n756));
  AOI21_X1  g555(.A(new_n745), .B1(new_n753), .B2(new_n756), .ZN(new_n757));
  AND2_X1   g556(.A1(new_n756), .A2(new_n745), .ZN(new_n758));
  OAI21_X1  g557(.A(KEYINPUT108), .B1(new_n757), .B2(new_n758), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n725), .A2(new_n740), .ZN(new_n760));
  AND4_X1   g559(.A1(new_n746), .A2(new_n760), .A3(new_n334), .A4(new_n755), .ZN(new_n761));
  AOI21_X1  g560(.A(new_n246), .B1(new_n741), .B2(new_n746), .ZN(new_n762));
  OAI21_X1  g561(.A(KEYINPUT42), .B1(new_n761), .B2(new_n762), .ZN(new_n763));
  INV_X1    g562(.A(KEYINPUT108), .ZN(new_n764));
  NAND2_X1  g563(.A1(new_n756), .A2(new_n745), .ZN(new_n765));
  NAND3_X1  g564(.A1(new_n763), .A2(new_n764), .A3(new_n765), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n759), .A2(new_n766), .ZN(G1325gat));
  INV_X1    g566(.A(new_n741), .ZN(new_n768));
  OAI21_X1  g567(.A(G15gat), .B1(new_n768), .B2(new_n730), .ZN(new_n769));
  NAND3_X1  g568(.A1(new_n741), .A2(new_n228), .A3(new_n632), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n769), .A2(new_n770), .ZN(G1326gat));
  NAND2_X1  g570(.A1(new_n741), .A2(new_n576), .ZN(new_n772));
  XNOR2_X1  g571(.A(KEYINPUT43), .B(G22gat), .ZN(new_n773));
  XNOR2_X1  g572(.A(new_n772), .B(new_n773), .ZN(G1327gat));
  INV_X1    g573(.A(new_n254), .ZN(new_n775));
  INV_X1    g574(.A(new_n333), .ZN(new_n776));
  NOR3_X1   g575(.A1(new_n775), .A2(new_n296), .A3(new_n776), .ZN(new_n777));
  AND2_X1   g576(.A1(new_n760), .A2(new_n777), .ZN(new_n778));
  XOR2_X1   g577(.A(KEYINPUT109), .B(KEYINPUT45), .Z(new_n779));
  NAND2_X1  g578(.A1(new_n742), .A2(new_n302), .ZN(new_n780));
  INV_X1    g579(.A(new_n780), .ZN(new_n781));
  AND3_X1   g580(.A1(new_n778), .A2(new_n779), .A3(new_n781), .ZN(new_n782));
  AOI21_X1  g581(.A(new_n779), .B1(new_n778), .B2(new_n781), .ZN(new_n783));
  NOR2_X1   g582(.A1(new_n782), .A2(new_n783), .ZN(new_n784));
  INV_X1    g583(.A(KEYINPUT110), .ZN(new_n785));
  NOR2_X1   g584(.A1(new_n785), .A2(KEYINPUT44), .ZN(new_n786));
  NAND2_X1  g585(.A1(new_n785), .A2(KEYINPUT44), .ZN(new_n787));
  INV_X1    g586(.A(new_n787), .ZN(new_n788));
  OAI22_X1  g587(.A1(new_n695), .A2(new_n776), .B1(new_n786), .B2(new_n788), .ZN(new_n789));
  NAND3_X1  g588(.A1(new_n749), .A2(new_n333), .A3(new_n787), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  NOR2_X1   g590(.A1(new_n775), .A2(new_n296), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n792), .A2(new_n723), .ZN(new_n793));
  INV_X1    g592(.A(new_n793), .ZN(new_n794));
  NAND3_X1  g593(.A1(new_n791), .A2(new_n742), .A3(new_n794), .ZN(new_n795));
  AOI21_X1  g594(.A(new_n302), .B1(new_n795), .B2(KEYINPUT111), .ZN(new_n796));
  OAI21_X1  g595(.A(new_n796), .B1(KEYINPUT111), .B2(new_n795), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n784), .A2(new_n797), .ZN(G1328gat));
  NAND3_X1  g597(.A1(new_n778), .A2(new_n298), .A3(new_n746), .ZN(new_n799));
  OR2_X1    g598(.A1(new_n799), .A2(KEYINPUT46), .ZN(new_n800));
  NAND3_X1  g599(.A1(new_n791), .A2(new_n746), .A3(new_n794), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n801), .A2(G36gat), .ZN(new_n802));
  NAND2_X1  g601(.A1(new_n799), .A2(KEYINPUT46), .ZN(new_n803));
  NAND3_X1  g602(.A1(new_n800), .A2(new_n802), .A3(new_n803), .ZN(G1329gat));
  INV_X1    g603(.A(new_n730), .ZN(new_n805));
  NAND4_X1  g604(.A1(new_n791), .A2(G43gat), .A3(new_n805), .A4(new_n794), .ZN(new_n806));
  INV_X1    g605(.A(KEYINPUT47), .ZN(new_n807));
  AND2_X1   g606(.A1(new_n778), .A2(new_n632), .ZN(new_n808));
  OAI211_X1 g607(.A(new_n806), .B(new_n807), .C1(new_n808), .C2(G43gat), .ZN(new_n809));
  AOI21_X1  g608(.A(G43gat), .B1(new_n778), .B2(new_n632), .ZN(new_n810));
  INV_X1    g609(.A(new_n806), .ZN(new_n811));
  OAI21_X1  g610(.A(KEYINPUT47), .B1(new_n810), .B2(new_n811), .ZN(new_n812));
  NAND2_X1  g611(.A1(new_n809), .A2(new_n812), .ZN(G1330gat));
  AOI211_X1 g612(.A(new_n634), .B(new_n793), .C1(new_n789), .C2(new_n790), .ZN(new_n814));
  INV_X1    g613(.A(G50gat), .ZN(new_n815));
  OAI21_X1  g614(.A(KEYINPUT112), .B1(new_n814), .B2(new_n815), .ZN(new_n816));
  NAND4_X1  g615(.A1(new_n760), .A2(new_n815), .A3(new_n576), .A4(new_n777), .ZN(new_n817));
  OAI21_X1  g616(.A(new_n817), .B1(new_n814), .B2(new_n815), .ZN(new_n818));
  INV_X1    g617(.A(KEYINPUT48), .ZN(new_n819));
  NAND3_X1  g618(.A1(new_n816), .A2(new_n818), .A3(new_n819), .ZN(new_n820));
  OAI221_X1 g619(.A(new_n817), .B1(KEYINPUT112), .B2(KEYINPUT48), .C1(new_n814), .C2(new_n815), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n820), .A2(new_n821), .ZN(G1331gat));
  NAND4_X1  g621(.A1(new_n775), .A2(new_n724), .A3(new_n296), .A4(new_n776), .ZN(new_n823));
  XNOR2_X1  g622(.A(new_n823), .B(KEYINPUT113), .ZN(new_n824));
  NOR2_X1   g623(.A1(new_n824), .A2(new_n695), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n825), .A2(new_n742), .ZN(new_n826));
  XNOR2_X1  g625(.A(new_n826), .B(G57gat), .ZN(G1332gat));
  AOI21_X1  g626(.A(new_n458), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n825), .A2(new_n828), .ZN(new_n829));
  XNOR2_X1  g628(.A(new_n829), .B(KEYINPUT114), .ZN(new_n830));
  NOR2_X1   g629(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n831));
  INV_X1    g630(.A(new_n831), .ZN(new_n832));
  XNOR2_X1  g631(.A(new_n830), .B(new_n832), .ZN(G1333gat));
  NAND2_X1  g632(.A1(new_n825), .A2(new_n805), .ZN(new_n834));
  INV_X1    g633(.A(new_n632), .ZN(new_n835));
  NOR2_X1   g634(.A1(new_n835), .A2(G71gat), .ZN(new_n836));
  AOI22_X1  g635(.A1(new_n834), .A2(G71gat), .B1(new_n825), .B2(new_n836), .ZN(new_n837));
  XNOR2_X1  g636(.A(new_n837), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g637(.A1(new_n825), .A2(new_n576), .ZN(new_n839));
  XNOR2_X1  g638(.A(new_n839), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g639(.A1(new_n775), .A2(new_n723), .ZN(new_n841));
  NAND2_X1  g640(.A1(new_n841), .A2(new_n296), .ZN(new_n842));
  AOI21_X1  g641(.A(new_n842), .B1(new_n789), .B2(new_n790), .ZN(new_n843));
  AND2_X1   g642(.A1(new_n843), .A2(new_n742), .ZN(new_n844));
  NAND3_X1  g643(.A1(new_n749), .A2(new_n333), .A3(new_n841), .ZN(new_n845));
  XNOR2_X1  g644(.A(new_n845), .B(KEYINPUT51), .ZN(new_n846));
  NAND3_X1  g645(.A1(new_n742), .A2(new_n261), .A3(new_n296), .ZN(new_n847));
  OAI22_X1  g646(.A1(new_n844), .A2(new_n261), .B1(new_n846), .B2(new_n847), .ZN(G1336gat));
  INV_X1    g647(.A(KEYINPUT116), .ZN(new_n849));
  NAND2_X1  g648(.A1(new_n845), .A2(new_n849), .ZN(new_n850));
  INV_X1    g649(.A(KEYINPUT51), .ZN(new_n851));
  NAND2_X1  g650(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  NAND3_X1  g651(.A1(new_n845), .A2(new_n849), .A3(KEYINPUT51), .ZN(new_n853));
  INV_X1    g652(.A(new_n296), .ZN(new_n854));
  NOR3_X1   g653(.A1(new_n458), .A2(G92gat), .A3(new_n854), .ZN(new_n855));
  NAND3_X1  g654(.A1(new_n852), .A2(new_n853), .A3(new_n855), .ZN(new_n856));
  AOI21_X1  g655(.A(new_n262), .B1(new_n843), .B2(new_n746), .ZN(new_n857));
  OAI21_X1  g656(.A(new_n856), .B1(new_n857), .B2(KEYINPUT115), .ZN(new_n858));
  INV_X1    g657(.A(KEYINPUT115), .ZN(new_n859));
  AOI211_X1 g658(.A(new_n859), .B(new_n262), .C1(new_n843), .C2(new_n746), .ZN(new_n860));
  OAI21_X1  g659(.A(KEYINPUT52), .B1(new_n858), .B2(new_n860), .ZN(new_n861));
  XOR2_X1   g660(.A(KEYINPUT117), .B(KEYINPUT52), .Z(new_n862));
  INV_X1    g661(.A(new_n855), .ZN(new_n863));
  OAI21_X1  g662(.A(new_n862), .B1(new_n846), .B2(new_n863), .ZN(new_n864));
  OR2_X1    g663(.A1(new_n864), .A2(new_n857), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n861), .A2(new_n865), .ZN(G1337gat));
  AND2_X1   g665(.A1(new_n843), .A2(new_n805), .ZN(new_n867));
  INV_X1    g666(.A(G99gat), .ZN(new_n868));
  NAND3_X1  g667(.A1(new_n632), .A2(new_n868), .A3(new_n296), .ZN(new_n869));
  OAI22_X1  g668(.A1(new_n867), .A2(new_n868), .B1(new_n846), .B2(new_n869), .ZN(G1338gat));
  NAND2_X1  g669(.A1(new_n852), .A2(new_n853), .ZN(new_n871));
  INV_X1    g670(.A(G106gat), .ZN(new_n872));
  NAND3_X1  g671(.A1(new_n296), .A2(new_n576), .A3(new_n872), .ZN(new_n873));
  NOR2_X1   g672(.A1(new_n871), .A2(new_n873), .ZN(new_n874));
  AOI21_X1  g673(.A(new_n872), .B1(new_n843), .B2(new_n576), .ZN(new_n875));
  OAI21_X1  g674(.A(KEYINPUT53), .B1(new_n874), .B2(new_n875), .ZN(new_n876));
  INV_X1    g675(.A(KEYINPUT53), .ZN(new_n877));
  OAI21_X1  g676(.A(new_n877), .B1(new_n846), .B2(new_n873), .ZN(new_n878));
  OAI21_X1  g677(.A(new_n876), .B1(new_n875), .B2(new_n878), .ZN(G1339gat));
  NOR4_X1   g678(.A1(new_n254), .A2(new_n723), .A3(new_n296), .A4(new_n333), .ZN(new_n880));
  INV_X1    g679(.A(KEYINPUT54), .ZN(new_n881));
  NOR2_X1   g680(.A1(new_n283), .A2(new_n881), .ZN(new_n882));
  NAND3_X1  g681(.A1(new_n280), .A2(new_n256), .A3(new_n282), .ZN(new_n883));
  NAND2_X1  g682(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  AOI221_X4 g683(.A(KEYINPUT10), .B1(new_n271), .B2(new_n272), .C1(new_n285), .C2(new_n278), .ZN(new_n885));
  INV_X1    g684(.A(new_n282), .ZN(new_n886));
  OAI211_X1 g685(.A(new_n881), .B(new_n284), .C1(new_n885), .C2(new_n886), .ZN(new_n887));
  INV_X1    g686(.A(KEYINPUT118), .ZN(new_n888));
  AND3_X1   g687(.A1(new_n887), .A2(new_n888), .A3(new_n292), .ZN(new_n889));
  AOI21_X1  g688(.A(new_n888), .B1(new_n887), .B2(new_n292), .ZN(new_n890));
  OAI21_X1  g689(.A(new_n884), .B1(new_n889), .B2(new_n890), .ZN(new_n891));
  INV_X1    g690(.A(KEYINPUT55), .ZN(new_n892));
  NAND2_X1  g691(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  NOR3_X1   g692(.A1(new_n709), .A2(new_n710), .A3(new_n708), .ZN(new_n894));
  AOI21_X1  g693(.A(new_n701), .B1(new_n696), .B2(new_n700), .ZN(new_n895));
  OAI21_X1  g694(.A(new_n718), .B1(new_n894), .B2(new_n895), .ZN(new_n896));
  AND2_X1   g695(.A1(new_n722), .A2(new_n896), .ZN(new_n897));
  NAND3_X1  g696(.A1(new_n893), .A2(new_n333), .A3(new_n897), .ZN(new_n898));
  OAI211_X1 g697(.A(KEYINPUT55), .B(new_n884), .C1(new_n889), .C2(new_n890), .ZN(new_n899));
  NAND2_X1  g698(.A1(new_n899), .A2(new_n294), .ZN(new_n900));
  OAI21_X1  g699(.A(KEYINPUT119), .B1(new_n898), .B2(new_n900), .ZN(new_n901));
  NAND4_X1  g700(.A1(new_n330), .A2(new_n722), .A3(new_n896), .A4(new_n332), .ZN(new_n902));
  AOI21_X1  g701(.A(new_n902), .B1(new_n892), .B2(new_n891), .ZN(new_n903));
  INV_X1    g702(.A(KEYINPUT119), .ZN(new_n904));
  NAND2_X1  g703(.A1(new_n887), .A2(new_n292), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n905), .A2(KEYINPUT118), .ZN(new_n906));
  NAND3_X1  g705(.A1(new_n887), .A2(new_n888), .A3(new_n292), .ZN(new_n907));
  AOI22_X1  g706(.A1(new_n906), .A2(new_n907), .B1(new_n883), .B2(new_n882), .ZN(new_n908));
  AOI21_X1  g707(.A(new_n293), .B1(new_n908), .B2(KEYINPUT55), .ZN(new_n909));
  NAND3_X1  g708(.A1(new_n903), .A2(new_n904), .A3(new_n909), .ZN(new_n910));
  NAND2_X1  g709(.A1(new_n897), .A2(new_n296), .ZN(new_n911));
  INV_X1    g710(.A(new_n911), .ZN(new_n912));
  AND3_X1   g711(.A1(new_n723), .A2(new_n899), .A3(new_n294), .ZN(new_n913));
  AOI21_X1  g712(.A(new_n912), .B1(new_n913), .B2(new_n893), .ZN(new_n914));
  OAI211_X1 g713(.A(new_n901), .B(new_n910), .C1(new_n914), .C2(new_n333), .ZN(new_n915));
  AOI21_X1  g714(.A(new_n880), .B1(new_n915), .B2(new_n254), .ZN(new_n916));
  NOR2_X1   g715(.A1(new_n746), .A2(new_n633), .ZN(new_n917));
  INV_X1    g716(.A(new_n917), .ZN(new_n918));
  NOR4_X1   g717(.A1(new_n916), .A2(new_n576), .A3(new_n835), .A4(new_n918), .ZN(new_n919));
  AOI21_X1  g718(.A(G113gat), .B1(new_n919), .B2(new_n723), .ZN(new_n920));
  NOR2_X1   g719(.A1(new_n916), .A2(new_n576), .ZN(new_n921));
  NAND3_X1  g720(.A1(new_n921), .A2(new_n632), .A3(new_n917), .ZN(new_n922));
  INV_X1    g721(.A(new_n922), .ZN(new_n923));
  NOR2_X1   g722(.A1(new_n724), .A2(new_n473), .ZN(new_n924));
  AOI21_X1  g723(.A(new_n920), .B1(new_n923), .B2(new_n924), .ZN(G1340gat));
  AOI21_X1  g724(.A(G120gat), .B1(new_n919), .B2(new_n296), .ZN(new_n926));
  NOR2_X1   g725(.A1(new_n854), .A2(new_n482), .ZN(new_n927));
  AOI21_X1  g726(.A(new_n926), .B1(new_n923), .B2(new_n927), .ZN(G1341gat));
  OAI21_X1  g727(.A(G127gat), .B1(new_n922), .B2(new_n254), .ZN(new_n929));
  NAND3_X1  g728(.A1(new_n919), .A2(new_n468), .A3(new_n775), .ZN(new_n930));
  NAND2_X1  g729(.A1(new_n929), .A2(new_n930), .ZN(G1342gat));
  NAND3_X1  g730(.A1(new_n919), .A2(new_n466), .A3(new_n333), .ZN(new_n932));
  OR2_X1    g731(.A1(new_n932), .A2(KEYINPUT56), .ZN(new_n933));
  OAI21_X1  g732(.A(G134gat), .B1(new_n922), .B2(new_n776), .ZN(new_n934));
  NAND2_X1  g733(.A1(new_n932), .A2(KEYINPUT56), .ZN(new_n935));
  NAND3_X1  g734(.A1(new_n933), .A2(new_n934), .A3(new_n935), .ZN(G1343gat));
  NAND2_X1  g735(.A1(new_n891), .A2(KEYINPUT121), .ZN(new_n937));
  INV_X1    g736(.A(KEYINPUT121), .ZN(new_n938));
  OAI211_X1 g737(.A(new_n938), .B(new_n884), .C1(new_n889), .C2(new_n890), .ZN(new_n939));
  NAND3_X1  g738(.A1(new_n937), .A2(new_n892), .A3(new_n939), .ZN(new_n940));
  AOI21_X1  g739(.A(new_n912), .B1(new_n940), .B2(new_n913), .ZN(new_n941));
  OAI211_X1 g740(.A(new_n901), .B(new_n910), .C1(new_n941), .C2(new_n333), .ZN(new_n942));
  AOI21_X1  g741(.A(new_n880), .B1(new_n942), .B2(new_n254), .ZN(new_n943));
  INV_X1    g742(.A(KEYINPUT57), .ZN(new_n944));
  NOR2_X1   g743(.A1(new_n634), .A2(new_n944), .ZN(new_n945));
  INV_X1    g744(.A(new_n945), .ZN(new_n946));
  OAI21_X1  g745(.A(KEYINPUT122), .B1(new_n943), .B2(new_n946), .ZN(new_n947));
  XOR2_X1   g746(.A(KEYINPUT120), .B(KEYINPUT57), .Z(new_n948));
  OAI21_X1  g747(.A(new_n948), .B1(new_n916), .B2(new_n634), .ZN(new_n949));
  INV_X1    g748(.A(KEYINPUT122), .ZN(new_n950));
  NOR3_X1   g749(.A1(new_n898), .A2(new_n900), .A3(KEYINPUT119), .ZN(new_n951));
  AOI21_X1  g750(.A(new_n904), .B1(new_n903), .B2(new_n909), .ZN(new_n952));
  NOR2_X1   g751(.A1(new_n951), .A2(new_n952), .ZN(new_n953));
  NAND3_X1  g752(.A1(new_n723), .A2(new_n899), .A3(new_n294), .ZN(new_n954));
  AOI21_X1  g753(.A(KEYINPUT55), .B1(new_n891), .B2(KEYINPUT121), .ZN(new_n955));
  AOI21_X1  g754(.A(new_n954), .B1(new_n939), .B2(new_n955), .ZN(new_n956));
  OAI21_X1  g755(.A(new_n776), .B1(new_n956), .B2(new_n912), .ZN(new_n957));
  AOI21_X1  g756(.A(new_n775), .B1(new_n953), .B2(new_n957), .ZN(new_n958));
  OAI211_X1 g757(.A(new_n950), .B(new_n945), .C1(new_n958), .C2(new_n880), .ZN(new_n959));
  NAND3_X1  g758(.A1(new_n947), .A2(new_n949), .A3(new_n959), .ZN(new_n960));
  NOR2_X1   g759(.A1(new_n918), .A2(new_n805), .ZN(new_n961));
  NAND3_X1  g760(.A1(new_n960), .A2(new_n723), .A3(new_n961), .ZN(new_n962));
  NAND2_X1  g761(.A1(new_n962), .A2(G141gat), .ZN(new_n963));
  NOR4_X1   g762(.A1(new_n916), .A2(new_n634), .A3(new_n805), .A4(new_n918), .ZN(new_n964));
  NAND3_X1  g763(.A1(new_n964), .A2(new_n521), .A3(new_n723), .ZN(new_n965));
  NAND2_X1  g764(.A1(new_n963), .A2(new_n965), .ZN(new_n966));
  NAND2_X1  g765(.A1(new_n966), .A2(KEYINPUT58), .ZN(new_n967));
  INV_X1    g766(.A(KEYINPUT58), .ZN(new_n968));
  NAND3_X1  g767(.A1(new_n963), .A2(new_n968), .A3(new_n965), .ZN(new_n969));
  NAND2_X1  g768(.A1(new_n967), .A2(new_n969), .ZN(G1344gat));
  NAND2_X1  g769(.A1(new_n901), .A2(new_n910), .ZN(new_n971));
  NAND3_X1  g770(.A1(new_n909), .A2(new_n723), .A3(new_n893), .ZN(new_n972));
  AOI21_X1  g771(.A(new_n333), .B1(new_n972), .B2(new_n911), .ZN(new_n973));
  OAI21_X1  g772(.A(new_n254), .B1(new_n971), .B2(new_n973), .ZN(new_n974));
  INV_X1    g773(.A(new_n880), .ZN(new_n975));
  NAND2_X1  g774(.A1(new_n974), .A2(new_n975), .ZN(new_n976));
  INV_X1    g775(.A(new_n948), .ZN(new_n977));
  NAND3_X1  g776(.A1(new_n976), .A2(new_n576), .A3(new_n977), .ZN(new_n978));
  OAI22_X1  g777(.A1(new_n941), .A2(new_n333), .B1(new_n900), .B2(new_n898), .ZN(new_n979));
  AOI21_X1  g778(.A(new_n880), .B1(new_n979), .B2(new_n254), .ZN(new_n980));
  OAI21_X1  g779(.A(new_n944), .B1(new_n980), .B2(new_n634), .ZN(new_n981));
  AND2_X1   g780(.A1(new_n978), .A2(new_n981), .ZN(new_n982));
  NAND2_X1  g781(.A1(new_n961), .A2(new_n296), .ZN(new_n983));
  OAI21_X1  g782(.A(G148gat), .B1(new_n982), .B2(new_n983), .ZN(new_n984));
  NAND2_X1  g783(.A1(new_n984), .A2(KEYINPUT59), .ZN(new_n985));
  NOR2_X1   g784(.A1(new_n523), .A2(KEYINPUT59), .ZN(new_n986));
  NAND2_X1  g785(.A1(new_n960), .A2(new_n961), .ZN(new_n987));
  OAI21_X1  g786(.A(new_n986), .B1(new_n987), .B2(new_n854), .ZN(new_n988));
  NAND2_X1  g787(.A1(new_n985), .A2(new_n988), .ZN(new_n989));
  NAND3_X1  g788(.A1(new_n964), .A2(new_n523), .A3(new_n296), .ZN(new_n990));
  NAND2_X1  g789(.A1(new_n989), .A2(new_n990), .ZN(G1345gat));
  OAI21_X1  g790(.A(G155gat), .B1(new_n987), .B2(new_n254), .ZN(new_n992));
  INV_X1    g791(.A(G155gat), .ZN(new_n993));
  NAND3_X1  g792(.A1(new_n964), .A2(new_n993), .A3(new_n775), .ZN(new_n994));
  NAND2_X1  g793(.A1(new_n992), .A2(new_n994), .ZN(G1346gat));
  INV_X1    g794(.A(G162gat), .ZN(new_n996));
  NAND3_X1  g795(.A1(new_n964), .A2(new_n996), .A3(new_n333), .ZN(new_n997));
  OAI21_X1  g796(.A(KEYINPUT123), .B1(new_n987), .B2(new_n776), .ZN(new_n998));
  NAND2_X1  g797(.A1(new_n998), .A2(G162gat), .ZN(new_n999));
  NOR3_X1   g798(.A1(new_n987), .A2(KEYINPUT123), .A3(new_n776), .ZN(new_n1000));
  OAI21_X1  g799(.A(new_n997), .B1(new_n999), .B2(new_n1000), .ZN(G1347gat));
  NOR2_X1   g800(.A1(new_n916), .A2(new_n742), .ZN(new_n1002));
  NAND3_X1  g801(.A1(new_n1002), .A2(new_n746), .A3(new_n578), .ZN(new_n1003));
  XNOR2_X1  g802(.A(new_n1003), .B(KEYINPUT124), .ZN(new_n1004));
  NAND3_X1  g803(.A1(new_n1004), .A2(new_n723), .A3(new_n401), .ZN(new_n1005));
  NAND2_X1  g804(.A1(new_n746), .A2(new_n633), .ZN(new_n1006));
  NOR2_X1   g805(.A1(new_n1006), .A2(new_n835), .ZN(new_n1007));
  AND2_X1   g806(.A1(new_n921), .A2(new_n1007), .ZN(new_n1008));
  INV_X1    g807(.A(new_n1008), .ZN(new_n1009));
  OAI21_X1  g808(.A(G169gat), .B1(new_n1009), .B2(new_n724), .ZN(new_n1010));
  NAND2_X1  g809(.A1(new_n1005), .A2(new_n1010), .ZN(G1348gat));
  NAND3_X1  g810(.A1(new_n1004), .A2(new_n337), .A3(new_n296), .ZN(new_n1012));
  OAI21_X1  g811(.A(G176gat), .B1(new_n1009), .B2(new_n854), .ZN(new_n1013));
  NAND2_X1  g812(.A1(new_n1012), .A2(new_n1013), .ZN(G1349gat));
  AOI21_X1  g813(.A(new_n383), .B1(new_n1008), .B2(new_n775), .ZN(new_n1015));
  NOR3_X1   g814(.A1(new_n1003), .A2(new_n345), .A3(new_n254), .ZN(new_n1016));
  NOR2_X1   g815(.A1(new_n1015), .A2(new_n1016), .ZN(new_n1017));
  INV_X1    g816(.A(KEYINPUT60), .ZN(new_n1018));
  XNOR2_X1  g817(.A(new_n1017), .B(new_n1018), .ZN(G1350gat));
  NAND3_X1  g818(.A1(new_n1004), .A2(new_n346), .A3(new_n333), .ZN(new_n1020));
  OAI21_X1  g819(.A(G190gat), .B1(new_n1009), .B2(new_n776), .ZN(new_n1021));
  AND2_X1   g820(.A1(new_n1021), .A2(KEYINPUT61), .ZN(new_n1022));
  NOR2_X1   g821(.A1(new_n1021), .A2(KEYINPUT61), .ZN(new_n1023));
  OAI21_X1  g822(.A(new_n1020), .B1(new_n1022), .B2(new_n1023), .ZN(G1351gat));
  NAND3_X1  g823(.A1(new_n730), .A2(new_n576), .A3(new_n746), .ZN(new_n1025));
  XNOR2_X1  g824(.A(new_n1025), .B(KEYINPUT125), .ZN(new_n1026));
  AND2_X1   g825(.A1(new_n1002), .A2(new_n1026), .ZN(new_n1027));
  AOI21_X1  g826(.A(G197gat), .B1(new_n1027), .B2(new_n723), .ZN(new_n1028));
  NOR2_X1   g827(.A1(new_n805), .A2(new_n1006), .ZN(new_n1029));
  XOR2_X1   g828(.A(new_n1029), .B(KEYINPUT126), .Z(new_n1030));
  NOR2_X1   g829(.A1(new_n982), .A2(new_n1030), .ZN(new_n1031));
  AND2_X1   g830(.A1(new_n723), .A2(G197gat), .ZN(new_n1032));
  AOI21_X1  g831(.A(new_n1028), .B1(new_n1031), .B2(new_n1032), .ZN(G1352gat));
  INV_X1    g832(.A(G204gat), .ZN(new_n1034));
  NAND3_X1  g833(.A1(new_n1027), .A2(new_n1034), .A3(new_n296), .ZN(new_n1035));
  OR2_X1    g834(.A1(new_n1035), .A2(KEYINPUT62), .ZN(new_n1036));
  NAND2_X1  g835(.A1(new_n1035), .A2(KEYINPUT62), .ZN(new_n1037));
  NOR3_X1   g836(.A1(new_n982), .A2(new_n854), .A3(new_n1030), .ZN(new_n1038));
  OAI211_X1 g837(.A(new_n1036), .B(new_n1037), .C1(new_n1034), .C2(new_n1038), .ZN(G1353gat));
  INV_X1    g838(.A(G211gat), .ZN(new_n1040));
  NAND3_X1  g839(.A1(new_n1027), .A2(new_n1040), .A3(new_n775), .ZN(new_n1041));
  NAND2_X1  g840(.A1(new_n1029), .A2(new_n775), .ZN(new_n1042));
  OAI21_X1  g841(.A(KEYINPUT127), .B1(new_n982), .B2(new_n1042), .ZN(new_n1043));
  AOI21_X1  g842(.A(new_n1042), .B1(new_n978), .B2(new_n981), .ZN(new_n1044));
  INV_X1    g843(.A(KEYINPUT127), .ZN(new_n1045));
  AOI21_X1  g844(.A(new_n1040), .B1(new_n1044), .B2(new_n1045), .ZN(new_n1046));
  AND3_X1   g845(.A1(new_n1043), .A2(new_n1046), .A3(KEYINPUT63), .ZN(new_n1047));
  AOI21_X1  g846(.A(KEYINPUT63), .B1(new_n1043), .B2(new_n1046), .ZN(new_n1048));
  OAI21_X1  g847(.A(new_n1041), .B1(new_n1047), .B2(new_n1048), .ZN(G1354gat));
  INV_X1    g848(.A(G218gat), .ZN(new_n1050));
  NAND3_X1  g849(.A1(new_n1027), .A2(new_n1050), .A3(new_n333), .ZN(new_n1051));
  NOR3_X1   g850(.A1(new_n982), .A2(new_n776), .A3(new_n1030), .ZN(new_n1052));
  OAI21_X1  g851(.A(new_n1051), .B1(new_n1052), .B2(new_n1050), .ZN(G1355gat));
endmodule


