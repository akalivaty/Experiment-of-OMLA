

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601,
         n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612,
         n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623,
         n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634,
         n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645,
         n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656,
         n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667,
         n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678,
         n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689,
         n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700,
         n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711,
         n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722,
         n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733,
         n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744,
         n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, n755,
         n756, n757, n758, n759, n760, n761, n762, n763, n764, n765, n766,
         n767, n768, n769, n770, n771, n772, n773, n774, n775, n776, n777,
         n778, n779, n780, n781, n782, n783, n784, n785, n786, n787, n788,
         n789, n790, n791, n792, n793, n794, n795, n796, n797, n798, n799,
         n800, n801, n802, n803, n804, n805, n806, n807, n808, n809, n810,
         n811, n812, n813, n814, n815, n816, n817, n818, n819, n820, n821,
         n822, n823, n824, n825, n826, n827, n828, n829, n830, n831, n832,
         n833, n834, n835, n836, n837, n838, n839, n840, n841, n842, n843,
         n844, n845, n846, n847, n848, n849, n850, n851, n852, n853, n854,
         n855, n856, n857, n858, n859, n860, n861, n862, n863, n864, n865,
         n866, n867, n868, n869, n870, n871, n872, n873, n874, n875, n876,
         n877, n878, n879, n880, n881, n882, n883, n884, n885, n886, n887,
         n888, n889, n890, n891, n892, n893, n894, n895, n896, n897, n898,
         n899, n900, n901, n902, n903, n904, n905, n906, n907, n908, n909,
         n910, n911, n912, n913, n914, n915, n916, n917, n918, n919, n920,
         n921, n922, n923, n924, n925, n926, n927, n928, n929, n930, n931,
         n932, n933, n934, n935, n936, n937, n938, n939, n940, n941, n942,
         n943, n944, n945, n946, n947, n948, n949, n950, n951, n952, n953,
         n954, n955, n956, n957, n958, n959, n960, n961, n962, n963, n964,
         n965, n966, n967, n968, n969, n970, n971, n972, n973, n974, n975,
         n976, n977, n978, n979, n980, n981, n982, n983, n984, n985, n986,
         n987, n988, n989, n990, n991, n992, n993, n994, n995, n996, n997,
         n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007,
         n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017,
         n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  OR2_X1 U553 ( .A1(n736), .A2(n735), .ZN(n752) );
  NOR2_X1 U554 ( .A1(n707), .A2(n898), .ZN(n701) );
  XNOR2_X1 U555 ( .A(KEYINPUT29), .B(KEYINPUT101), .ZN(n721) );
  XNOR2_X1 U556 ( .A(n722), .B(n721), .ZN(n723) );
  NOR2_X2 U557 ( .A1(n691), .A2(n690), .ZN(n711) );
  NOR2_X1 U558 ( .A1(G164), .A2(G1384), .ZN(n689) );
  AND2_X1 U559 ( .A1(G2104), .A2(G2105), .ZN(n873) );
  NAND2_X1 U560 ( .A1(G114), .A2(n873), .ZN(n522) );
  INV_X1 U561 ( .A(G2105), .ZN(n524) );
  NOR2_X1 U562 ( .A1(G2104), .A2(n524), .ZN(n874) );
  NAND2_X1 U563 ( .A1(G126), .A2(n874), .ZN(n521) );
  NAND2_X1 U564 ( .A1(n522), .A2(n521), .ZN(n530) );
  NOR2_X1 U565 ( .A1(G2104), .A2(G2105), .ZN(n523) );
  XOR2_X2 U566 ( .A(KEYINPUT17), .B(n523), .Z(n869) );
  NAND2_X1 U567 ( .A1(G138), .A2(n869), .ZN(n526) );
  AND2_X1 U568 ( .A1(n524), .A2(G2104), .ZN(n870) );
  NAND2_X1 U569 ( .A1(G102), .A2(n870), .ZN(n525) );
  NAND2_X1 U570 ( .A1(n526), .A2(n525), .ZN(n528) );
  INV_X1 U571 ( .A(KEYINPUT93), .ZN(n527) );
  XNOR2_X1 U572 ( .A(n528), .B(n527), .ZN(n529) );
  NOR2_X1 U573 ( .A1(n530), .A2(n529), .ZN(G164) );
  INV_X1 U574 ( .A(KEYINPUT23), .ZN(n532) );
  NAND2_X1 U575 ( .A1(n870), .A2(G101), .ZN(n531) );
  XNOR2_X1 U576 ( .A(n532), .B(n531), .ZN(n534) );
  NAND2_X1 U577 ( .A1(n874), .A2(G125), .ZN(n533) );
  NAND2_X1 U578 ( .A1(n534), .A2(n533), .ZN(n535) );
  XNOR2_X1 U579 ( .A(n535), .B(KEYINPUT65), .ZN(n537) );
  NAND2_X1 U580 ( .A1(G113), .A2(n873), .ZN(n536) );
  AND2_X1 U581 ( .A1(n537), .A2(n536), .ZN(n540) );
  NAND2_X1 U582 ( .A1(n869), .A2(G137), .ZN(n538) );
  XNOR2_X1 U583 ( .A(KEYINPUT66), .B(n538), .ZN(n539) );
  AND2_X1 U584 ( .A1(n540), .A2(n539), .ZN(G160) );
  INV_X1 U585 ( .A(G57), .ZN(G237) );
  INV_X1 U586 ( .A(G120), .ZN(G236) );
  INV_X1 U587 ( .A(G132), .ZN(G219) );
  INV_X1 U588 ( .A(G82), .ZN(G220) );
  XNOR2_X1 U589 ( .A(G651), .B(KEYINPUT67), .ZN(n546) );
  NOR2_X1 U590 ( .A1(G543), .A2(n546), .ZN(n541) );
  XOR2_X1 U591 ( .A(KEYINPUT1), .B(n541), .Z(n654) );
  NAND2_X1 U592 ( .A1(G64), .A2(n654), .ZN(n544) );
  XOR2_X1 U593 ( .A(KEYINPUT0), .B(G543), .Z(n626) );
  NOR2_X1 U594 ( .A1(G651), .A2(n626), .ZN(n542) );
  XNOR2_X1 U595 ( .A(KEYINPUT64), .B(n542), .ZN(n653) );
  NAND2_X1 U596 ( .A1(G52), .A2(n653), .ZN(n543) );
  NAND2_X1 U597 ( .A1(n544), .A2(n543), .ZN(n551) );
  NOR2_X1 U598 ( .A1(G651), .A2(G543), .ZN(n649) );
  NAND2_X1 U599 ( .A1(n649), .A2(G90), .ZN(n545) );
  XNOR2_X1 U600 ( .A(n545), .B(KEYINPUT70), .ZN(n548) );
  NOR2_X1 U601 ( .A1(n626), .A2(n546), .ZN(n647) );
  NAND2_X1 U602 ( .A1(G77), .A2(n647), .ZN(n547) );
  NAND2_X1 U603 ( .A1(n548), .A2(n547), .ZN(n549) );
  XOR2_X1 U604 ( .A(KEYINPUT9), .B(n549), .Z(n550) );
  NOR2_X1 U605 ( .A1(n551), .A2(n550), .ZN(G171) );
  NAND2_X1 U606 ( .A1(G89), .A2(n649), .ZN(n552) );
  XOR2_X1 U607 ( .A(KEYINPUT77), .B(n552), .Z(n553) );
  XNOR2_X1 U608 ( .A(n553), .B(KEYINPUT4), .ZN(n555) );
  NAND2_X1 U609 ( .A1(G76), .A2(n647), .ZN(n554) );
  NAND2_X1 U610 ( .A1(n555), .A2(n554), .ZN(n556) );
  XNOR2_X1 U611 ( .A(KEYINPUT5), .B(n556), .ZN(n563) );
  XNOR2_X1 U612 ( .A(KEYINPUT78), .B(KEYINPUT79), .ZN(n561) );
  NAND2_X1 U613 ( .A1(G63), .A2(n654), .ZN(n558) );
  NAND2_X1 U614 ( .A1(G51), .A2(n653), .ZN(n557) );
  NAND2_X1 U615 ( .A1(n558), .A2(n557), .ZN(n559) );
  XNOR2_X1 U616 ( .A(n559), .B(KEYINPUT6), .ZN(n560) );
  XNOR2_X1 U617 ( .A(n561), .B(n560), .ZN(n562) );
  NAND2_X1 U618 ( .A1(n563), .A2(n562), .ZN(n564) );
  XNOR2_X1 U619 ( .A(KEYINPUT7), .B(n564), .ZN(G168) );
  XOR2_X1 U620 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U621 ( .A1(G94), .A2(G452), .ZN(n565) );
  XNOR2_X1 U622 ( .A(n565), .B(KEYINPUT71), .ZN(G173) );
  NAND2_X1 U623 ( .A1(G7), .A2(G661), .ZN(n566) );
  XNOR2_X1 U624 ( .A(n566), .B(KEYINPUT10), .ZN(G223) );
  XOR2_X1 U625 ( .A(G223), .B(KEYINPUT74), .Z(n824) );
  NAND2_X1 U626 ( .A1(n824), .A2(G567), .ZN(n567) );
  XOR2_X1 U627 ( .A(KEYINPUT11), .B(n567), .Z(G234) );
  NAND2_X1 U628 ( .A1(n654), .A2(G56), .ZN(n568) );
  XNOR2_X1 U629 ( .A(KEYINPUT14), .B(n568), .ZN(n578) );
  XNOR2_X1 U630 ( .A(KEYINPUT13), .B(KEYINPUT75), .ZN(n573) );
  NAND2_X1 U631 ( .A1(n649), .A2(G81), .ZN(n569) );
  XNOR2_X1 U632 ( .A(n569), .B(KEYINPUT12), .ZN(n571) );
  NAND2_X1 U633 ( .A1(G68), .A2(n647), .ZN(n570) );
  NAND2_X1 U634 ( .A1(n571), .A2(n570), .ZN(n572) );
  XNOR2_X1 U635 ( .A(n573), .B(n572), .ZN(n576) );
  NAND2_X1 U636 ( .A1(n653), .A2(G43), .ZN(n574) );
  XOR2_X1 U637 ( .A(KEYINPUT76), .B(n574), .Z(n575) );
  NOR2_X1 U638 ( .A1(n576), .A2(n575), .ZN(n577) );
  NAND2_X1 U639 ( .A1(n578), .A2(n577), .ZN(n1000) );
  INV_X1 U640 ( .A(G860), .ZN(n599) );
  OR2_X1 U641 ( .A1(n1000), .A2(n599), .ZN(G153) );
  INV_X1 U642 ( .A(G171), .ZN(G301) );
  NAND2_X1 U643 ( .A1(G868), .A2(G301), .ZN(n587) );
  NAND2_X1 U644 ( .A1(G79), .A2(n647), .ZN(n580) );
  NAND2_X1 U645 ( .A1(G54), .A2(n653), .ZN(n579) );
  NAND2_X1 U646 ( .A1(n580), .A2(n579), .ZN(n584) );
  NAND2_X1 U647 ( .A1(G92), .A2(n649), .ZN(n582) );
  NAND2_X1 U648 ( .A1(G66), .A2(n654), .ZN(n581) );
  NAND2_X1 U649 ( .A1(n582), .A2(n581), .ZN(n583) );
  NOR2_X1 U650 ( .A1(n584), .A2(n583), .ZN(n585) );
  XOR2_X1 U651 ( .A(n585), .B(KEYINPUT15), .Z(n1005) );
  INV_X1 U652 ( .A(n1005), .ZN(n898) );
  INV_X1 U653 ( .A(G868), .ZN(n669) );
  NAND2_X1 U654 ( .A1(n898), .A2(n669), .ZN(n586) );
  NAND2_X1 U655 ( .A1(n587), .A2(n586), .ZN(G284) );
  NAND2_X1 U656 ( .A1(n647), .A2(G78), .ZN(n588) );
  XNOR2_X1 U657 ( .A(n588), .B(KEYINPUT72), .ZN(n590) );
  NAND2_X1 U658 ( .A1(G91), .A2(n649), .ZN(n589) );
  NAND2_X1 U659 ( .A1(n590), .A2(n589), .ZN(n591) );
  XNOR2_X1 U660 ( .A(KEYINPUT73), .B(n591), .ZN(n595) );
  NAND2_X1 U661 ( .A1(n653), .A2(G53), .ZN(n593) );
  NAND2_X1 U662 ( .A1(G65), .A2(n654), .ZN(n592) );
  AND2_X1 U663 ( .A1(n593), .A2(n592), .ZN(n594) );
  NAND2_X1 U664 ( .A1(n595), .A2(n594), .ZN(G299) );
  NOR2_X1 U665 ( .A1(G286), .A2(n669), .ZN(n596) );
  XNOR2_X1 U666 ( .A(n596), .B(KEYINPUT80), .ZN(n598) );
  NOR2_X1 U667 ( .A1(G299), .A2(G868), .ZN(n597) );
  NOR2_X1 U668 ( .A1(n598), .A2(n597), .ZN(G297) );
  NAND2_X1 U669 ( .A1(n599), .A2(G559), .ZN(n600) );
  NAND2_X1 U670 ( .A1(n600), .A2(n1005), .ZN(n601) );
  XNOR2_X1 U671 ( .A(n601), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U672 ( .A1(n898), .A2(n669), .ZN(n602) );
  XNOR2_X1 U673 ( .A(n602), .B(KEYINPUT81), .ZN(n603) );
  NOR2_X1 U674 ( .A1(G559), .A2(n603), .ZN(n605) );
  NOR2_X1 U675 ( .A1(G868), .A2(n1000), .ZN(n604) );
  NOR2_X1 U676 ( .A1(n605), .A2(n604), .ZN(G282) );
  NAND2_X1 U677 ( .A1(G123), .A2(n874), .ZN(n606) );
  XNOR2_X1 U678 ( .A(n606), .B(KEYINPUT18), .ZN(n608) );
  NAND2_X1 U679 ( .A1(n869), .A2(G135), .ZN(n607) );
  NAND2_X1 U680 ( .A1(n608), .A2(n607), .ZN(n612) );
  NAND2_X1 U681 ( .A1(G99), .A2(n870), .ZN(n610) );
  NAND2_X1 U682 ( .A1(G111), .A2(n873), .ZN(n609) );
  NAND2_X1 U683 ( .A1(n610), .A2(n609), .ZN(n611) );
  NOR2_X1 U684 ( .A1(n612), .A2(n611), .ZN(n920) );
  XOR2_X1 U685 ( .A(n920), .B(G2096), .Z(n613) );
  XNOR2_X1 U686 ( .A(KEYINPUT82), .B(n613), .ZN(n614) );
  NOR2_X1 U687 ( .A1(G2100), .A2(n614), .ZN(n615) );
  XNOR2_X1 U688 ( .A(KEYINPUT83), .B(n615), .ZN(G156) );
  NAND2_X1 U689 ( .A1(n1005), .A2(G559), .ZN(n666) );
  XNOR2_X1 U690 ( .A(n1000), .B(n666), .ZN(n616) );
  NOR2_X1 U691 ( .A1(n616), .A2(G860), .ZN(n625) );
  NAND2_X1 U692 ( .A1(G80), .A2(n647), .ZN(n618) );
  NAND2_X1 U693 ( .A1(G67), .A2(n654), .ZN(n617) );
  NAND2_X1 U694 ( .A1(n618), .A2(n617), .ZN(n621) );
  NAND2_X1 U695 ( .A1(G93), .A2(n649), .ZN(n619) );
  XNOR2_X1 U696 ( .A(KEYINPUT85), .B(n619), .ZN(n620) );
  NOR2_X1 U697 ( .A1(n621), .A2(n620), .ZN(n623) );
  NAND2_X1 U698 ( .A1(G55), .A2(n653), .ZN(n622) );
  NAND2_X1 U699 ( .A1(n623), .A2(n622), .ZN(n668) );
  XOR2_X1 U700 ( .A(n668), .B(KEYINPUT84), .Z(n624) );
  XNOR2_X1 U701 ( .A(n625), .B(n624), .ZN(G145) );
  NAND2_X1 U702 ( .A1(G87), .A2(n626), .ZN(n628) );
  NAND2_X1 U703 ( .A1(G74), .A2(G651), .ZN(n627) );
  NAND2_X1 U704 ( .A1(n628), .A2(n627), .ZN(n629) );
  NOR2_X1 U705 ( .A1(n654), .A2(n629), .ZN(n631) );
  NAND2_X1 U706 ( .A1(G49), .A2(n653), .ZN(n630) );
  NAND2_X1 U707 ( .A1(n631), .A2(n630), .ZN(G288) );
  NAND2_X1 U708 ( .A1(n653), .A2(G48), .ZN(n638) );
  NAND2_X1 U709 ( .A1(G86), .A2(n649), .ZN(n633) );
  NAND2_X1 U710 ( .A1(G61), .A2(n654), .ZN(n632) );
  NAND2_X1 U711 ( .A1(n633), .A2(n632), .ZN(n636) );
  NAND2_X1 U712 ( .A1(n647), .A2(G73), .ZN(n634) );
  XOR2_X1 U713 ( .A(KEYINPUT2), .B(n634), .Z(n635) );
  NOR2_X1 U714 ( .A1(n636), .A2(n635), .ZN(n637) );
  NAND2_X1 U715 ( .A1(n638), .A2(n637), .ZN(n639) );
  XNOR2_X1 U716 ( .A(n639), .B(KEYINPUT86), .ZN(G305) );
  NAND2_X1 U717 ( .A1(G88), .A2(n649), .ZN(n641) );
  NAND2_X1 U718 ( .A1(G62), .A2(n654), .ZN(n640) );
  NAND2_X1 U719 ( .A1(n641), .A2(n640), .ZN(n644) );
  NAND2_X1 U720 ( .A1(G75), .A2(n647), .ZN(n642) );
  XNOR2_X1 U721 ( .A(KEYINPUT87), .B(n642), .ZN(n643) );
  NOR2_X1 U722 ( .A1(n644), .A2(n643), .ZN(n646) );
  NAND2_X1 U723 ( .A1(G50), .A2(n653), .ZN(n645) );
  NAND2_X1 U724 ( .A1(n646), .A2(n645), .ZN(G303) );
  NAND2_X1 U725 ( .A1(n647), .A2(G72), .ZN(n648) );
  XNOR2_X1 U726 ( .A(n648), .B(KEYINPUT68), .ZN(n651) );
  NAND2_X1 U727 ( .A1(G85), .A2(n649), .ZN(n650) );
  NAND2_X1 U728 ( .A1(n651), .A2(n650), .ZN(n652) );
  XNOR2_X1 U729 ( .A(KEYINPUT69), .B(n652), .ZN(n658) );
  NAND2_X1 U730 ( .A1(n653), .A2(G47), .ZN(n656) );
  NAND2_X1 U731 ( .A1(G60), .A2(n654), .ZN(n655) );
  AND2_X1 U732 ( .A1(n656), .A2(n655), .ZN(n657) );
  NAND2_X1 U733 ( .A1(n658), .A2(n657), .ZN(G290) );
  XOR2_X1 U734 ( .A(KEYINPUT19), .B(KEYINPUT88), .Z(n659) );
  XNOR2_X1 U735 ( .A(n1000), .B(n659), .ZN(n660) );
  XNOR2_X1 U736 ( .A(n660), .B(G288), .ZN(n663) );
  XOR2_X1 U737 ( .A(G305), .B(G303), .Z(n661) );
  XNOR2_X1 U738 ( .A(n661), .B(n668), .ZN(n662) );
  XNOR2_X1 U739 ( .A(n663), .B(n662), .ZN(n664) );
  XOR2_X1 U740 ( .A(G299), .B(n664), .Z(n665) );
  XNOR2_X1 U741 ( .A(n665), .B(G290), .ZN(n896) );
  XNOR2_X1 U742 ( .A(n666), .B(n896), .ZN(n667) );
  NAND2_X1 U743 ( .A1(n667), .A2(G868), .ZN(n671) );
  NAND2_X1 U744 ( .A1(n669), .A2(n668), .ZN(n670) );
  NAND2_X1 U745 ( .A1(n671), .A2(n670), .ZN(G295) );
  NAND2_X1 U746 ( .A1(G2084), .A2(G2078), .ZN(n672) );
  XNOR2_X1 U747 ( .A(n672), .B(KEYINPUT20), .ZN(n673) );
  XNOR2_X1 U748 ( .A(KEYINPUT89), .B(n673), .ZN(n674) );
  NAND2_X1 U749 ( .A1(n674), .A2(G2090), .ZN(n675) );
  XNOR2_X1 U750 ( .A(KEYINPUT21), .B(n675), .ZN(n676) );
  NAND2_X1 U751 ( .A1(n676), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U752 ( .A(KEYINPUT90), .B(G44), .ZN(n677) );
  XNOR2_X1 U753 ( .A(n677), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U754 ( .A1(G220), .A2(G219), .ZN(n678) );
  XOR2_X1 U755 ( .A(KEYINPUT22), .B(n678), .Z(n679) );
  NOR2_X1 U756 ( .A1(G218), .A2(n679), .ZN(n680) );
  NAND2_X1 U757 ( .A1(G96), .A2(n680), .ZN(n831) );
  AND2_X1 U758 ( .A1(G2106), .A2(n831), .ZN(n686) );
  NOR2_X1 U759 ( .A1(G236), .A2(G237), .ZN(n681) );
  NAND2_X1 U760 ( .A1(G69), .A2(n681), .ZN(n682) );
  XNOR2_X1 U761 ( .A(KEYINPUT91), .B(n682), .ZN(n683) );
  NAND2_X1 U762 ( .A1(n683), .A2(G108), .ZN(n830) );
  NAND2_X1 U763 ( .A1(G567), .A2(n830), .ZN(n684) );
  XOR2_X1 U764 ( .A(KEYINPUT92), .B(n684), .Z(n685) );
  NOR2_X1 U765 ( .A1(n686), .A2(n685), .ZN(G319) );
  INV_X1 U766 ( .A(G319), .ZN(n688) );
  NAND2_X1 U767 ( .A1(G483), .A2(G661), .ZN(n687) );
  NOR2_X1 U768 ( .A1(n688), .A2(n687), .ZN(n828) );
  NAND2_X1 U769 ( .A1(n828), .A2(G36), .ZN(G176) );
  XNOR2_X1 U770 ( .A(G1986), .B(G290), .ZN(n1015) );
  NAND2_X1 U771 ( .A1(G160), .A2(G40), .ZN(n690) );
  NOR2_X1 U772 ( .A1(n689), .A2(n690), .ZN(n819) );
  NAND2_X1 U773 ( .A1(n1015), .A2(n819), .ZN(n807) );
  INV_X1 U774 ( .A(n689), .ZN(n691) );
  INV_X1 U775 ( .A(n711), .ZN(n737) );
  NAND2_X1 U776 ( .A1(G8), .A2(n737), .ZN(n761) );
  NOR2_X1 U777 ( .A1(G1981), .A2(G305), .ZN(n692) );
  XOR2_X1 U778 ( .A(n692), .B(KEYINPUT24), .Z(n693) );
  NOR2_X1 U779 ( .A1(n761), .A2(n693), .ZN(n777) );
  INV_X1 U780 ( .A(G1961), .ZN(n837) );
  NAND2_X1 U781 ( .A1(n737), .A2(n837), .ZN(n695) );
  XNOR2_X1 U782 ( .A(G2078), .B(KEYINPUT25), .ZN(n972) );
  NAND2_X1 U783 ( .A1(n711), .A2(n972), .ZN(n694) );
  NAND2_X1 U784 ( .A1(n695), .A2(n694), .ZN(n728) );
  AND2_X1 U785 ( .A1(n728), .A2(G171), .ZN(n696) );
  XOR2_X1 U786 ( .A(KEYINPUT98), .B(n696), .Z(n724) );
  NAND2_X1 U787 ( .A1(G1996), .A2(n711), .ZN(n697) );
  XOR2_X1 U788 ( .A(KEYINPUT26), .B(n697), .Z(n698) );
  NOR2_X1 U789 ( .A1(n1000), .A2(n698), .ZN(n700) );
  NAND2_X1 U790 ( .A1(G1341), .A2(n737), .ZN(n699) );
  NAND2_X1 U791 ( .A1(n700), .A2(n699), .ZN(n707) );
  XNOR2_X1 U792 ( .A(n701), .B(KEYINPUT99), .ZN(n706) );
  NAND2_X1 U793 ( .A1(n737), .A2(G1348), .ZN(n702) );
  XNOR2_X1 U794 ( .A(n702), .B(KEYINPUT100), .ZN(n704) );
  NAND2_X1 U795 ( .A1(n711), .A2(G2067), .ZN(n703) );
  NAND2_X1 U796 ( .A1(n704), .A2(n703), .ZN(n705) );
  NAND2_X1 U797 ( .A1(n706), .A2(n705), .ZN(n709) );
  NAND2_X1 U798 ( .A1(n707), .A2(n898), .ZN(n708) );
  NAND2_X1 U799 ( .A1(n709), .A2(n708), .ZN(n715) );
  INV_X1 U800 ( .A(G299), .ZN(n717) );
  NAND2_X1 U801 ( .A1(n711), .A2(G2072), .ZN(n710) );
  XNOR2_X1 U802 ( .A(n710), .B(KEYINPUT27), .ZN(n713) );
  INV_X1 U803 ( .A(G1956), .ZN(n1009) );
  NOR2_X1 U804 ( .A1(n1009), .A2(n711), .ZN(n712) );
  NOR2_X1 U805 ( .A1(n713), .A2(n712), .ZN(n716) );
  NAND2_X1 U806 ( .A1(n717), .A2(n716), .ZN(n714) );
  NAND2_X1 U807 ( .A1(n715), .A2(n714), .ZN(n720) );
  NOR2_X1 U808 ( .A1(n717), .A2(n716), .ZN(n718) );
  XOR2_X1 U809 ( .A(n718), .B(KEYINPUT28), .Z(n719) );
  NAND2_X1 U810 ( .A1(n720), .A2(n719), .ZN(n722) );
  NAND2_X1 U811 ( .A1(n724), .A2(n723), .ZN(n745) );
  NOR2_X1 U812 ( .A1(G1966), .A2(n761), .ZN(n733) );
  NOR2_X1 U813 ( .A1(G2084), .A2(n737), .ZN(n732) );
  NOR2_X1 U814 ( .A1(n733), .A2(n732), .ZN(n725) );
  NAND2_X1 U815 ( .A1(G8), .A2(n725), .ZN(n726) );
  XNOR2_X1 U816 ( .A(KEYINPUT30), .B(n726), .ZN(n727) );
  NOR2_X1 U817 ( .A1(G168), .A2(n727), .ZN(n730) );
  NOR2_X1 U818 ( .A1(G171), .A2(n728), .ZN(n729) );
  NOR2_X1 U819 ( .A1(n730), .A2(n729), .ZN(n731) );
  XOR2_X1 U820 ( .A(KEYINPUT31), .B(n731), .Z(n743) );
  AND2_X1 U821 ( .A1(n745), .A2(n743), .ZN(n736) );
  AND2_X1 U822 ( .A1(G8), .A2(n732), .ZN(n734) );
  OR2_X1 U823 ( .A1(n734), .A2(n733), .ZN(n735) );
  INV_X1 U824 ( .A(G8), .ZN(n742) );
  NOR2_X1 U825 ( .A1(G1971), .A2(n761), .ZN(n739) );
  NOR2_X1 U826 ( .A1(G2090), .A2(n737), .ZN(n738) );
  NOR2_X1 U827 ( .A1(n739), .A2(n738), .ZN(n740) );
  NAND2_X1 U828 ( .A1(n740), .A2(G303), .ZN(n741) );
  OR2_X1 U829 ( .A1(n742), .A2(n741), .ZN(n746) );
  AND2_X1 U830 ( .A1(n743), .A2(n746), .ZN(n744) );
  NAND2_X1 U831 ( .A1(n745), .A2(n744), .ZN(n749) );
  INV_X1 U832 ( .A(n746), .ZN(n747) );
  OR2_X1 U833 ( .A1(n747), .A2(G286), .ZN(n748) );
  NAND2_X1 U834 ( .A1(n749), .A2(n748), .ZN(n750) );
  XNOR2_X1 U835 ( .A(n750), .B(KEYINPUT32), .ZN(n751) );
  NAND2_X1 U836 ( .A1(n752), .A2(n751), .ZN(n770) );
  NOR2_X1 U837 ( .A1(G2090), .A2(G303), .ZN(n753) );
  NAND2_X1 U838 ( .A1(G8), .A2(n753), .ZN(n754) );
  NAND2_X1 U839 ( .A1(n770), .A2(n754), .ZN(n755) );
  NAND2_X1 U840 ( .A1(n755), .A2(n761), .ZN(n774) );
  XOR2_X1 U841 ( .A(G1981), .B(G305), .Z(n756) );
  XNOR2_X1 U842 ( .A(KEYINPUT104), .B(n756), .ZN(n996) );
  NAND2_X1 U843 ( .A1(G1976), .A2(G288), .ZN(n1008) );
  INV_X1 U844 ( .A(n1008), .ZN(n757) );
  NOR2_X1 U845 ( .A1(n761), .A2(n757), .ZN(n758) );
  NOR2_X1 U846 ( .A1(KEYINPUT33), .A2(n758), .ZN(n763) );
  NOR2_X1 U847 ( .A1(G1976), .A2(G288), .ZN(n766) );
  NAND2_X1 U848 ( .A1(KEYINPUT33), .A2(n766), .ZN(n759) );
  XOR2_X1 U849 ( .A(KEYINPUT103), .B(n759), .Z(n760) );
  NOR2_X1 U850 ( .A1(n761), .A2(n760), .ZN(n762) );
  NOR2_X1 U851 ( .A1(n763), .A2(n762), .ZN(n764) );
  AND2_X1 U852 ( .A1(n996), .A2(n764), .ZN(n772) );
  NOR2_X1 U853 ( .A1(G1971), .A2(G303), .ZN(n765) );
  NOR2_X1 U854 ( .A1(n766), .A2(n765), .ZN(n1013) );
  XNOR2_X1 U855 ( .A(KEYINPUT102), .B(n1013), .ZN(n768) );
  INV_X1 U856 ( .A(KEYINPUT33), .ZN(n767) );
  AND2_X1 U857 ( .A1(n768), .A2(n767), .ZN(n769) );
  NAND2_X1 U858 ( .A1(n770), .A2(n769), .ZN(n771) );
  NAND2_X1 U859 ( .A1(n772), .A2(n771), .ZN(n773) );
  NAND2_X1 U860 ( .A1(n774), .A2(n773), .ZN(n775) );
  XOR2_X1 U861 ( .A(KEYINPUT105), .B(n775), .Z(n776) );
  NOR2_X1 U862 ( .A1(n777), .A2(n776), .ZN(n805) );
  NAND2_X1 U863 ( .A1(G140), .A2(n869), .ZN(n779) );
  NAND2_X1 U864 ( .A1(G104), .A2(n870), .ZN(n778) );
  NAND2_X1 U865 ( .A1(n779), .A2(n778), .ZN(n780) );
  XNOR2_X1 U866 ( .A(KEYINPUT34), .B(n780), .ZN(n787) );
  NAND2_X1 U867 ( .A1(n873), .A2(G116), .ZN(n781) );
  XNOR2_X1 U868 ( .A(KEYINPUT95), .B(n781), .ZN(n784) );
  NAND2_X1 U869 ( .A1(n874), .A2(G128), .ZN(n782) );
  XOR2_X1 U870 ( .A(KEYINPUT94), .B(n782), .Z(n783) );
  NOR2_X1 U871 ( .A1(n784), .A2(n783), .ZN(n785) );
  XNOR2_X1 U872 ( .A(n785), .B(KEYINPUT35), .ZN(n786) );
  NOR2_X1 U873 ( .A1(n787), .A2(n786), .ZN(n788) );
  XNOR2_X1 U874 ( .A(KEYINPUT36), .B(n788), .ZN(n885) );
  XNOR2_X1 U875 ( .A(G2067), .B(KEYINPUT37), .ZN(n816) );
  NOR2_X1 U876 ( .A1(n885), .A2(n816), .ZN(n931) );
  NAND2_X1 U877 ( .A1(n819), .A2(n931), .ZN(n814) );
  NAND2_X1 U878 ( .A1(G141), .A2(n869), .ZN(n790) );
  NAND2_X1 U879 ( .A1(G117), .A2(n873), .ZN(n789) );
  NAND2_X1 U880 ( .A1(n790), .A2(n789), .ZN(n793) );
  NAND2_X1 U881 ( .A1(n870), .A2(G105), .ZN(n791) );
  XOR2_X1 U882 ( .A(KEYINPUT38), .B(n791), .Z(n792) );
  NOR2_X1 U883 ( .A1(n793), .A2(n792), .ZN(n795) );
  NAND2_X1 U884 ( .A1(n874), .A2(G129), .ZN(n794) );
  NAND2_X1 U885 ( .A1(n795), .A2(n794), .ZN(n884) );
  AND2_X1 U886 ( .A1(n884), .A2(G1996), .ZN(n921) );
  NAND2_X1 U887 ( .A1(G131), .A2(n869), .ZN(n797) );
  NAND2_X1 U888 ( .A1(G107), .A2(n873), .ZN(n796) );
  NAND2_X1 U889 ( .A1(n797), .A2(n796), .ZN(n800) );
  NAND2_X1 U890 ( .A1(n874), .A2(G119), .ZN(n798) );
  XOR2_X1 U891 ( .A(KEYINPUT96), .B(n798), .Z(n799) );
  NOR2_X1 U892 ( .A1(n800), .A2(n799), .ZN(n802) );
  NAND2_X1 U893 ( .A1(n870), .A2(G95), .ZN(n801) );
  AND2_X1 U894 ( .A1(n802), .A2(n801), .ZN(n889) );
  XNOR2_X1 U895 ( .A(KEYINPUT97), .B(G1991), .ZN(n973) );
  NOR2_X1 U896 ( .A1(n889), .A2(n973), .ZN(n927) );
  OR2_X1 U897 ( .A1(n921), .A2(n927), .ZN(n803) );
  NAND2_X1 U898 ( .A1(n803), .A2(n819), .ZN(n808) );
  NAND2_X1 U899 ( .A1(n814), .A2(n808), .ZN(n804) );
  NOR2_X1 U900 ( .A1(n805), .A2(n804), .ZN(n806) );
  NAND2_X1 U901 ( .A1(n807), .A2(n806), .ZN(n822) );
  NOR2_X1 U902 ( .A1(G1996), .A2(n884), .ZN(n917) );
  INV_X1 U903 ( .A(n808), .ZN(n811) );
  NOR2_X1 U904 ( .A1(G1986), .A2(G290), .ZN(n809) );
  AND2_X1 U905 ( .A1(n973), .A2(n889), .ZN(n923) );
  NOR2_X1 U906 ( .A1(n809), .A2(n923), .ZN(n810) );
  NOR2_X1 U907 ( .A1(n811), .A2(n810), .ZN(n812) );
  NOR2_X1 U908 ( .A1(n917), .A2(n812), .ZN(n813) );
  XNOR2_X1 U909 ( .A(n813), .B(KEYINPUT39), .ZN(n815) );
  NAND2_X1 U910 ( .A1(n815), .A2(n814), .ZN(n817) );
  NAND2_X1 U911 ( .A1(n885), .A2(n816), .ZN(n932) );
  NAND2_X1 U912 ( .A1(n817), .A2(n932), .ZN(n818) );
  XNOR2_X1 U913 ( .A(KEYINPUT106), .B(n818), .ZN(n820) );
  NAND2_X1 U914 ( .A1(n820), .A2(n819), .ZN(n821) );
  NAND2_X1 U915 ( .A1(n822), .A2(n821), .ZN(n823) );
  XNOR2_X1 U916 ( .A(KEYINPUT40), .B(n823), .ZN(G329) );
  NAND2_X1 U917 ( .A1(G2106), .A2(n824), .ZN(G217) );
  NAND2_X1 U918 ( .A1(G15), .A2(G2), .ZN(n825) );
  XNOR2_X1 U919 ( .A(KEYINPUT107), .B(n825), .ZN(n826) );
  NAND2_X1 U920 ( .A1(n826), .A2(G661), .ZN(G259) );
  NAND2_X1 U921 ( .A1(G3), .A2(G1), .ZN(n827) );
  XNOR2_X1 U922 ( .A(KEYINPUT108), .B(n827), .ZN(n829) );
  NAND2_X1 U923 ( .A1(n829), .A2(n828), .ZN(G188) );
  INV_X1 U925 ( .A(G108), .ZN(G238) );
  INV_X1 U926 ( .A(G96), .ZN(G221) );
  NOR2_X1 U927 ( .A1(n831), .A2(n830), .ZN(G325) );
  INV_X1 U928 ( .A(G325), .ZN(G261) );
  XOR2_X1 U929 ( .A(KEYINPUT110), .B(G1981), .Z(n833) );
  XNOR2_X1 U930 ( .A(G1996), .B(G1991), .ZN(n832) );
  XNOR2_X1 U931 ( .A(n833), .B(n832), .ZN(n834) );
  XOR2_X1 U932 ( .A(n834), .B(KEYINPUT41), .Z(n836) );
  XNOR2_X1 U933 ( .A(G1986), .B(G1976), .ZN(n835) );
  XNOR2_X1 U934 ( .A(n836), .B(n835), .ZN(n841) );
  XNOR2_X1 U935 ( .A(G1971), .B(n837), .ZN(n839) );
  XOR2_X1 U936 ( .A(G1966), .B(n1009), .Z(n838) );
  XNOR2_X1 U937 ( .A(n839), .B(n838), .ZN(n840) );
  XOR2_X1 U938 ( .A(n841), .B(n840), .Z(n843) );
  XNOR2_X1 U939 ( .A(G2474), .B(KEYINPUT111), .ZN(n842) );
  XNOR2_X1 U940 ( .A(n843), .B(n842), .ZN(G229) );
  XOR2_X1 U941 ( .A(KEYINPUT42), .B(G2090), .Z(n845) );
  XNOR2_X1 U942 ( .A(G2067), .B(G2084), .ZN(n844) );
  XNOR2_X1 U943 ( .A(n845), .B(n844), .ZN(n846) );
  XOR2_X1 U944 ( .A(n846), .B(G2100), .Z(n848) );
  XNOR2_X1 U945 ( .A(G2072), .B(G2078), .ZN(n847) );
  XNOR2_X1 U946 ( .A(n848), .B(n847), .ZN(n852) );
  XOR2_X1 U947 ( .A(G2096), .B(KEYINPUT43), .Z(n850) );
  XNOR2_X1 U948 ( .A(G2678), .B(KEYINPUT109), .ZN(n849) );
  XNOR2_X1 U949 ( .A(n850), .B(n849), .ZN(n851) );
  XOR2_X1 U950 ( .A(n852), .B(n851), .Z(G227) );
  NAND2_X1 U951 ( .A1(G124), .A2(n874), .ZN(n853) );
  XNOR2_X1 U952 ( .A(n853), .B(KEYINPUT44), .ZN(n855) );
  NAND2_X1 U953 ( .A1(n873), .A2(G112), .ZN(n854) );
  NAND2_X1 U954 ( .A1(n855), .A2(n854), .ZN(n859) );
  NAND2_X1 U955 ( .A1(G136), .A2(n869), .ZN(n857) );
  NAND2_X1 U956 ( .A1(G100), .A2(n870), .ZN(n856) );
  NAND2_X1 U957 ( .A1(n857), .A2(n856), .ZN(n858) );
  NOR2_X1 U958 ( .A1(n859), .A2(n858), .ZN(G162) );
  NAND2_X1 U959 ( .A1(G142), .A2(n869), .ZN(n861) );
  NAND2_X1 U960 ( .A1(G106), .A2(n870), .ZN(n860) );
  NAND2_X1 U961 ( .A1(n861), .A2(n860), .ZN(n862) );
  XNOR2_X1 U962 ( .A(n862), .B(KEYINPUT45), .ZN(n867) );
  NAND2_X1 U963 ( .A1(G118), .A2(n873), .ZN(n864) );
  NAND2_X1 U964 ( .A1(G130), .A2(n874), .ZN(n863) );
  NAND2_X1 U965 ( .A1(n864), .A2(n863), .ZN(n865) );
  XOR2_X1 U966 ( .A(KEYINPUT112), .B(n865), .Z(n866) );
  NAND2_X1 U967 ( .A1(n867), .A2(n866), .ZN(n868) );
  XNOR2_X1 U968 ( .A(n868), .B(G160), .ZN(n893) );
  NAND2_X1 U969 ( .A1(G139), .A2(n869), .ZN(n872) );
  NAND2_X1 U970 ( .A1(G103), .A2(n870), .ZN(n871) );
  NAND2_X1 U971 ( .A1(n872), .A2(n871), .ZN(n880) );
  NAND2_X1 U972 ( .A1(G115), .A2(n873), .ZN(n876) );
  NAND2_X1 U973 ( .A1(G127), .A2(n874), .ZN(n875) );
  NAND2_X1 U974 ( .A1(n876), .A2(n875), .ZN(n877) );
  XNOR2_X1 U975 ( .A(KEYINPUT47), .B(n877), .ZN(n878) );
  XNOR2_X1 U976 ( .A(KEYINPUT113), .B(n878), .ZN(n879) );
  NOR2_X1 U977 ( .A1(n880), .A2(n879), .ZN(n935) );
  XOR2_X1 U978 ( .A(KEYINPUT114), .B(KEYINPUT48), .Z(n882) );
  XNOR2_X1 U979 ( .A(n920), .B(KEYINPUT46), .ZN(n881) );
  XNOR2_X1 U980 ( .A(n882), .B(n881), .ZN(n883) );
  XNOR2_X1 U981 ( .A(n935), .B(n883), .ZN(n887) );
  XOR2_X1 U982 ( .A(n885), .B(n884), .Z(n886) );
  XNOR2_X1 U983 ( .A(n887), .B(n886), .ZN(n888) );
  XOR2_X1 U984 ( .A(n888), .B(G162), .Z(n891) );
  XNOR2_X1 U985 ( .A(G164), .B(n889), .ZN(n890) );
  XNOR2_X1 U986 ( .A(n891), .B(n890), .ZN(n892) );
  XOR2_X1 U987 ( .A(n893), .B(n892), .Z(n894) );
  NOR2_X1 U988 ( .A1(G37), .A2(n894), .ZN(n895) );
  XOR2_X1 U989 ( .A(KEYINPUT115), .B(n895), .Z(G395) );
  XOR2_X1 U990 ( .A(G286), .B(G171), .Z(n897) );
  XNOR2_X1 U991 ( .A(n897), .B(n896), .ZN(n899) );
  XOR2_X1 U992 ( .A(n899), .B(n898), .Z(n900) );
  NOR2_X1 U993 ( .A1(G37), .A2(n900), .ZN(G397) );
  XOR2_X1 U994 ( .A(G2451), .B(G2430), .Z(n902) );
  XNOR2_X1 U995 ( .A(G2438), .B(G2443), .ZN(n901) );
  XNOR2_X1 U996 ( .A(n902), .B(n901), .ZN(n908) );
  XOR2_X1 U997 ( .A(G2435), .B(G2454), .Z(n904) );
  XNOR2_X1 U998 ( .A(G1341), .B(G1348), .ZN(n903) );
  XNOR2_X1 U999 ( .A(n904), .B(n903), .ZN(n906) );
  XOR2_X1 U1000 ( .A(G2446), .B(G2427), .Z(n905) );
  XNOR2_X1 U1001 ( .A(n906), .B(n905), .ZN(n907) );
  XOR2_X1 U1002 ( .A(n908), .B(n907), .Z(n909) );
  NAND2_X1 U1003 ( .A1(G14), .A2(n909), .ZN(n915) );
  NAND2_X1 U1004 ( .A1(G319), .A2(n915), .ZN(n912) );
  NOR2_X1 U1005 ( .A1(G229), .A2(G227), .ZN(n910) );
  XNOR2_X1 U1006 ( .A(KEYINPUT49), .B(n910), .ZN(n911) );
  NOR2_X1 U1007 ( .A1(n912), .A2(n911), .ZN(n914) );
  NOR2_X1 U1008 ( .A1(G395), .A2(G397), .ZN(n913) );
  NAND2_X1 U1009 ( .A1(n914), .A2(n913), .ZN(G225) );
  INV_X1 U1010 ( .A(G225), .ZN(G308) );
  INV_X1 U1011 ( .A(G69), .ZN(G235) );
  INV_X1 U1012 ( .A(n915), .ZN(G401) );
  XNOR2_X1 U1013 ( .A(KEYINPUT55), .B(KEYINPUT118), .ZN(n988) );
  XOR2_X1 U1014 ( .A(G2090), .B(G162), .Z(n916) );
  NOR2_X1 U1015 ( .A1(n917), .A2(n916), .ZN(n918) );
  XOR2_X1 U1016 ( .A(KEYINPUT116), .B(n918), .Z(n919) );
  XNOR2_X1 U1017 ( .A(KEYINPUT51), .B(n919), .ZN(n929) );
  NOR2_X1 U1018 ( .A1(n921), .A2(n920), .ZN(n925) );
  XOR2_X1 U1019 ( .A(G160), .B(G2084), .Z(n922) );
  NOR2_X1 U1020 ( .A1(n923), .A2(n922), .ZN(n924) );
  NAND2_X1 U1021 ( .A1(n925), .A2(n924), .ZN(n926) );
  NOR2_X1 U1022 ( .A1(n927), .A2(n926), .ZN(n928) );
  NAND2_X1 U1023 ( .A1(n929), .A2(n928), .ZN(n930) );
  NOR2_X1 U1024 ( .A1(n931), .A2(n930), .ZN(n933) );
  NAND2_X1 U1025 ( .A1(n933), .A2(n932), .ZN(n934) );
  XOR2_X1 U1026 ( .A(KEYINPUT117), .B(n934), .Z(n940) );
  XOR2_X1 U1027 ( .A(G2072), .B(n935), .Z(n937) );
  XOR2_X1 U1028 ( .A(G164), .B(G2078), .Z(n936) );
  NOR2_X1 U1029 ( .A1(n937), .A2(n936), .ZN(n938) );
  XOR2_X1 U1030 ( .A(KEYINPUT50), .B(n938), .Z(n939) );
  NOR2_X1 U1031 ( .A1(n940), .A2(n939), .ZN(n941) );
  XOR2_X1 U1032 ( .A(KEYINPUT52), .B(n941), .Z(n942) );
  NOR2_X1 U1033 ( .A1(n988), .A2(n942), .ZN(n943) );
  XNOR2_X1 U1034 ( .A(KEYINPUT119), .B(n943), .ZN(n944) );
  NAND2_X1 U1035 ( .A1(n944), .A2(G29), .ZN(n995) );
  XOR2_X1 U1036 ( .A(G5), .B(G1961), .Z(n957) );
  XOR2_X1 U1037 ( .A(G1348), .B(KEYINPUT59), .Z(n945) );
  XNOR2_X1 U1038 ( .A(G4), .B(n945), .ZN(n952) );
  XOR2_X1 U1039 ( .A(G1981), .B(G6), .Z(n947) );
  XOR2_X1 U1040 ( .A(G1956), .B(G20), .Z(n946) );
  NAND2_X1 U1041 ( .A1(n947), .A2(n946), .ZN(n949) );
  XNOR2_X1 U1042 ( .A(G19), .B(G1341), .ZN(n948) );
  NOR2_X1 U1043 ( .A1(n949), .A2(n948), .ZN(n950) );
  XNOR2_X1 U1044 ( .A(n950), .B(KEYINPUT125), .ZN(n951) );
  NOR2_X1 U1045 ( .A1(n952), .A2(n951), .ZN(n953) );
  XOR2_X1 U1046 ( .A(KEYINPUT60), .B(n953), .Z(n955) );
  XNOR2_X1 U1047 ( .A(G1966), .B(G21), .ZN(n954) );
  NOR2_X1 U1048 ( .A1(n955), .A2(n954), .ZN(n956) );
  NAND2_X1 U1049 ( .A1(n957), .A2(n956), .ZN(n965) );
  XNOR2_X1 U1050 ( .A(G1986), .B(G24), .ZN(n959) );
  XNOR2_X1 U1051 ( .A(G23), .B(G1976), .ZN(n958) );
  NOR2_X1 U1052 ( .A1(n959), .A2(n958), .ZN(n962) );
  XOR2_X1 U1053 ( .A(G1971), .B(KEYINPUT126), .Z(n960) );
  XNOR2_X1 U1054 ( .A(G22), .B(n960), .ZN(n961) );
  NAND2_X1 U1055 ( .A1(n962), .A2(n961), .ZN(n963) );
  XNOR2_X1 U1056 ( .A(KEYINPUT58), .B(n963), .ZN(n964) );
  NOR2_X1 U1057 ( .A1(n965), .A2(n964), .ZN(n966) );
  XOR2_X1 U1058 ( .A(KEYINPUT61), .B(n966), .Z(n967) );
  NOR2_X1 U1059 ( .A1(G16), .A2(n967), .ZN(n968) );
  XOR2_X1 U1060 ( .A(KEYINPUT127), .B(n968), .Z(n993) );
  XOR2_X1 U1061 ( .A(G2090), .B(G35), .Z(n983) );
  XOR2_X1 U1062 ( .A(G32), .B(G1996), .Z(n969) );
  NAND2_X1 U1063 ( .A1(n969), .A2(G28), .ZN(n979) );
  XNOR2_X1 U1064 ( .A(G2067), .B(G26), .ZN(n971) );
  XNOR2_X1 U1065 ( .A(G33), .B(G2072), .ZN(n970) );
  NOR2_X1 U1066 ( .A1(n971), .A2(n970), .ZN(n977) );
  XOR2_X1 U1067 ( .A(n972), .B(G27), .Z(n975) );
  XOR2_X1 U1068 ( .A(n973), .B(G25), .Z(n974) );
  NOR2_X1 U1069 ( .A1(n975), .A2(n974), .ZN(n976) );
  NAND2_X1 U1070 ( .A1(n977), .A2(n976), .ZN(n978) );
  NOR2_X1 U1071 ( .A1(n979), .A2(n978), .ZN(n980) );
  XOR2_X1 U1072 ( .A(KEYINPUT120), .B(n980), .Z(n981) );
  XNOR2_X1 U1073 ( .A(n981), .B(KEYINPUT53), .ZN(n982) );
  NAND2_X1 U1074 ( .A1(n983), .A2(n982), .ZN(n986) );
  XNOR2_X1 U1075 ( .A(G34), .B(G2084), .ZN(n984) );
  XNOR2_X1 U1076 ( .A(KEYINPUT54), .B(n984), .ZN(n985) );
  NOR2_X1 U1077 ( .A1(n986), .A2(n985), .ZN(n987) );
  XNOR2_X1 U1078 ( .A(n988), .B(n987), .ZN(n990) );
  INV_X1 U1079 ( .A(G29), .ZN(n989) );
  NAND2_X1 U1080 ( .A1(n990), .A2(n989), .ZN(n991) );
  NAND2_X1 U1081 ( .A1(n991), .A2(G11), .ZN(n992) );
  NOR2_X1 U1082 ( .A1(n993), .A2(n992), .ZN(n994) );
  NAND2_X1 U1083 ( .A1(n995), .A2(n994), .ZN(n1025) );
  XOR2_X1 U1084 ( .A(KEYINPUT56), .B(G16), .Z(n1023) );
  XNOR2_X1 U1085 ( .A(G1966), .B(G168), .ZN(n997) );
  NAND2_X1 U1086 ( .A1(n997), .A2(n996), .ZN(n998) );
  XNOR2_X1 U1087 ( .A(n998), .B(KEYINPUT57), .ZN(n1004) );
  XOR2_X1 U1088 ( .A(G301), .B(KEYINPUT122), .Z(n999) );
  XOR2_X1 U1089 ( .A(n999), .B(G1961), .Z(n1002) );
  XNOR2_X1 U1090 ( .A(G1341), .B(n1000), .ZN(n1001) );
  NOR2_X1 U1091 ( .A1(n1002), .A2(n1001), .ZN(n1003) );
  NAND2_X1 U1092 ( .A1(n1004), .A2(n1003), .ZN(n1020) );
  XNOR2_X1 U1093 ( .A(G1348), .B(KEYINPUT121), .ZN(n1006) );
  XOR2_X1 U1094 ( .A(n1006), .B(n1005), .Z(n1018) );
  NAND2_X1 U1095 ( .A1(G1971), .A2(G303), .ZN(n1007) );
  NAND2_X1 U1096 ( .A1(n1008), .A2(n1007), .ZN(n1011) );
  XOR2_X1 U1097 ( .A(n1009), .B(G299), .Z(n1010) );
  NOR2_X1 U1098 ( .A1(n1011), .A2(n1010), .ZN(n1012) );
  NAND2_X1 U1099 ( .A1(n1013), .A2(n1012), .ZN(n1014) );
  NOR2_X1 U1100 ( .A1(n1015), .A2(n1014), .ZN(n1016) );
  XOR2_X1 U1101 ( .A(KEYINPUT123), .B(n1016), .Z(n1017) );
  NAND2_X1 U1102 ( .A1(n1018), .A2(n1017), .ZN(n1019) );
  NOR2_X1 U1103 ( .A1(n1020), .A2(n1019), .ZN(n1021) );
  XNOR2_X1 U1104 ( .A(KEYINPUT124), .B(n1021), .ZN(n1022) );
  NOR2_X1 U1105 ( .A1(n1023), .A2(n1022), .ZN(n1024) );
  NOR2_X1 U1106 ( .A1(n1025), .A2(n1024), .ZN(n1026) );
  XOR2_X1 U1107 ( .A(n1026), .B(KEYINPUT62), .Z(G150) );
  INV_X1 U1108 ( .A(G150), .ZN(G311) );
  INV_X1 U1109 ( .A(G303), .ZN(G166) );
endmodule

