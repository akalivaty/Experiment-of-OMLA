

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360,
         n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371,
         n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382,
         n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393,
         n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404,
         n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415,
         n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426,
         n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437,
         n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448,
         n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459,
         n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470,
         n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481,
         n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492,
         n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503,
         n504, n505, n506, n507, n508, n509, n510, n511, n512, n513, n514,
         n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525,
         n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536,
         n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547,
         n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558,
         n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569,
         n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580,
         n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591,
         n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602,
         n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613,
         n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624,
         n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635,
         n636, n637, n638, n639, n640, n641, n643, n644, n645, n646, n647,
         n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659,
         n660, n661, n663, n664, n665, n666, n667, n668, n669, n670, n671,
         n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682,
         n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693,
         n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704,
         n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715,
         n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726,
         n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737,
         n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748,
         n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759,
         n760, n761, n762, n763, n764, n765, n766;

  AND2_X1 U372 ( .A1(n351), .A2(n350), .ZN(n650) );
  AND2_X1 U373 ( .A1(n354), .A2(n353), .ZN(n663) );
  AND2_X1 U374 ( .A1(n357), .A2(n356), .ZN(n644) );
  INV_X1 U375 ( .A(n738), .ZN(n350) );
  INV_X1 U376 ( .A(n738), .ZN(n353) );
  INV_X1 U377 ( .A(n738), .ZN(n356) );
  AND2_X1 U378 ( .A1(n626), .A2(n625), .ZN(n627) );
  NOR2_X1 U379 ( .A1(n696), .A2(n594), .ZN(n666) );
  XNOR2_X1 U380 ( .A(n647), .B(n352), .ZN(n351) );
  INV_X1 U381 ( .A(n646), .ZN(n352) );
  XNOR2_X1 U382 ( .A(n661), .B(n355), .ZN(n354) );
  INV_X1 U383 ( .A(n660), .ZN(n355) );
  XNOR2_X1 U384 ( .A(n641), .B(n358), .ZN(n357) );
  INV_X1 U385 ( .A(n640), .ZN(n358) );
  AND2_X2 U386 ( .A1(n743), .A2(n421), .ZN(n420) );
  INV_X1 U387 ( .A(G953), .ZN(n757) );
  NAND2_X1 U388 ( .A1(n743), .A2(n423), .ZN(n729) );
  XNOR2_X2 U389 ( .A(n384), .B(n500), .ZN(n652) );
  XNOR2_X2 U390 ( .A(n750), .B(G146), .ZN(n384) );
  NAND2_X1 U391 ( .A1(n627), .A2(n628), .ZN(n365) );
  XNOR2_X1 U392 ( .A(n607), .B(KEYINPUT89), .ZN(n628) );
  XNOR2_X1 U393 ( .A(n429), .B(n427), .ZN(n762) );
  XNOR2_X1 U394 ( .A(n527), .B(KEYINPUT1), .ZN(n571) );
  NAND2_X1 U395 ( .A1(n405), .A2(n403), .ZN(n527) );
  AND2_X1 U396 ( .A1(n407), .A2(n406), .ZN(n405) );
  XNOR2_X1 U397 ( .A(n410), .B(n409), .ZN(n408) );
  XNOR2_X1 U398 ( .A(n494), .B(n493), .ZN(n750) );
  AND2_X1 U399 ( .A1(n630), .A2(n629), .ZN(n421) );
  XNOR2_X1 U400 ( .A(n464), .B(n438), .ZN(n751) );
  XNOR2_X1 U401 ( .A(n418), .B(n447), .ZN(n492) );
  XNOR2_X1 U402 ( .A(n415), .B(G146), .ZN(n464) );
  INV_X1 U403 ( .A(G125), .ZN(n415) );
  XNOR2_X1 U404 ( .A(KEYINPUT66), .B(KEYINPUT67), .ZN(n418) );
  XNOR2_X2 U405 ( .A(n370), .B(G143), .ZN(n391) );
  XNOR2_X2 U406 ( .A(G128), .B(KEYINPUT82), .ZN(n370) );
  NAND2_X2 U407 ( .A1(n568), .A2(n707), .ZN(n416) );
  XNOR2_X2 U408 ( .A(n474), .B(n473), .ZN(n568) );
  INV_X1 U409 ( .A(KEYINPUT68), .ZN(n389) );
  XNOR2_X1 U410 ( .A(n751), .B(n437), .ZN(n436) );
  INV_X1 U411 ( .A(KEYINPUT24), .ZN(n437) );
  NAND2_X1 U412 ( .A1(n396), .A2(n395), .ZN(n394) );
  INV_X1 U413 ( .A(n583), .ZN(n395) );
  AND2_X1 U414 ( .A1(n762), .A2(n766), .ZN(n558) );
  NOR2_X1 U415 ( .A1(n373), .A2(n372), .ZN(n371) );
  AND2_X1 U416 ( .A1(n710), .A2(n376), .ZN(n372) );
  OR2_X1 U417 ( .A1(n652), .A2(n404), .ZN(n403) );
  NAND2_X1 U418 ( .A1(G469), .A2(n513), .ZN(n404) );
  OR2_X1 U419 ( .A1(G902), .A2(G237), .ZN(n515) );
  AND2_X1 U420 ( .A1(n677), .A2(n530), .ZN(n390) );
  NAND2_X1 U421 ( .A1(n488), .A2(G217), .ZN(n410) );
  XNOR2_X1 U422 ( .A(n384), .B(n512), .ZN(n639) );
  XNOR2_X1 U423 ( .A(n387), .B(n386), .ZN(n385) );
  XNOR2_X1 U424 ( .A(n479), .B(n436), .ZN(n484) );
  XNOR2_X1 U425 ( .A(G137), .B(G119), .ZN(n481) );
  XNOR2_X1 U426 ( .A(n756), .B(KEYINPUT79), .ZN(n419) );
  XNOR2_X1 U427 ( .A(n739), .B(KEYINPUT72), .ZN(n499) );
  XNOR2_X1 U428 ( .A(n463), .B(G478), .ZN(n547) );
  NOR2_X1 U429 ( .A1(n710), .A2(n376), .ZN(n375) );
  INV_X1 U430 ( .A(KEYINPUT105), .ZN(n376) );
  AND2_X1 U431 ( .A1(n679), .A2(n375), .ZN(n373) );
  NAND2_X1 U432 ( .A1(n501), .A2(G902), .ZN(n406) );
  XNOR2_X1 U433 ( .A(n556), .B(KEYINPUT46), .ZN(n557) );
  OR2_X1 U434 ( .A1(n592), .A2(KEYINPUT34), .ZN(n398) );
  NOR2_X1 U435 ( .A1(G953), .A2(G237), .ZN(n508) );
  INV_X1 U436 ( .A(KEYINPUT48), .ZN(n386) );
  AND2_X1 U437 ( .A1(n381), .A2(n380), .ZN(n605) );
  XOR2_X1 U438 ( .A(KEYINPUT71), .B(KEYINPUT23), .Z(n477) );
  XNOR2_X1 U439 ( .A(G110), .B(G128), .ZN(n475) );
  XNOR2_X1 U440 ( .A(G113), .B(G143), .ZN(n442) );
  XOR2_X1 U441 ( .A(KEYINPUT101), .B(KEYINPUT11), .Z(n443) );
  INV_X1 U442 ( .A(G131), .ZN(n447) );
  XNOR2_X1 U443 ( .A(KEYINPUT10), .B(G140), .ZN(n438) );
  NOR2_X1 U444 ( .A1(n413), .A2(G953), .ZN(n412) );
  INV_X1 U445 ( .A(G224), .ZN(n413) );
  XNOR2_X1 U446 ( .A(n452), .B(n451), .ZN(n548) );
  BUF_X1 U447 ( .A(n527), .Z(n533) );
  XNOR2_X1 U448 ( .A(n470), .B(n469), .ZN(n511) );
  INV_X1 U449 ( .A(G113), .ZN(n467) );
  XOR2_X1 U450 ( .A(KEYINPUT103), .B(KEYINPUT102), .Z(n455) );
  XNOR2_X1 U451 ( .A(n391), .B(G134), .ZN(n494) );
  XNOR2_X1 U452 ( .A(n391), .B(n368), .ZN(n367) );
  XNOR2_X1 U453 ( .A(n369), .B(KEYINPUT80), .ZN(n368) );
  XNOR2_X1 U454 ( .A(KEYINPUT4), .B(KEYINPUT17), .ZN(n369) );
  XNOR2_X1 U455 ( .A(n411), .B(n400), .ZN(n399) );
  XNOR2_X1 U456 ( .A(n414), .B(n412), .ZN(n411) );
  INV_X1 U457 ( .A(n464), .ZN(n400) );
  XNOR2_X1 U458 ( .A(KEYINPUT93), .B(KEYINPUT18), .ZN(n414) );
  BUF_X1 U459 ( .A(n588), .Z(n697) );
  XNOR2_X1 U460 ( .A(KEYINPUT25), .B(KEYINPUT99), .ZN(n409) );
  NOR2_X1 U461 ( .A1(n533), .A2(n686), .ZN(n417) );
  XOR2_X1 U462 ( .A(KEYINPUT62), .B(n639), .Z(n640) );
  XNOR2_X1 U463 ( .A(n511), .B(n431), .ZN(n740) );
  XNOR2_X1 U464 ( .A(n472), .B(KEYINPUT16), .ZN(n431) );
  INV_X1 U465 ( .A(n471), .ZN(n472) );
  NAND2_X2 U466 ( .A1(n422), .A2(n402), .ZN(n734) );
  NAND2_X1 U467 ( .A1(n729), .A2(n434), .ZN(n422) );
  NOR2_X1 U468 ( .A1(n485), .A2(n629), .ZN(n434) );
  XNOR2_X1 U469 ( .A(n645), .B(KEYINPUT59), .ZN(n646) );
  XNOR2_X1 U470 ( .A(n366), .B(n740), .ZN(n659) );
  XNOR2_X1 U471 ( .A(n433), .B(n432), .ZN(n366) );
  INV_X1 U472 ( .A(n499), .ZN(n432) );
  XNOR2_X1 U473 ( .A(n367), .B(n399), .ZN(n433) );
  AND2_X1 U474 ( .A1(n634), .A2(G953), .ZN(n738) );
  NAND2_X1 U475 ( .A1(n729), .A2(KEYINPUT2), .ZN(n726) );
  XNOR2_X1 U476 ( .A(n426), .B(n424), .ZN(n766) );
  XNOR2_X1 U477 ( .A(n425), .B(KEYINPUT42), .ZN(n424) );
  OR2_X1 U478 ( .A1(n703), .A2(n551), .ZN(n426) );
  INV_X1 U479 ( .A(KEYINPUT113), .ZN(n425) );
  XNOR2_X1 U480 ( .A(n428), .B(KEYINPUT40), .ZN(n427) );
  AND2_X1 U481 ( .A1(n559), .A2(n677), .ZN(n429) );
  INV_X1 U482 ( .A(KEYINPUT112), .ZN(n428) );
  INV_X1 U483 ( .A(KEYINPUT36), .ZN(n401) );
  XOR2_X1 U484 ( .A(KEYINPUT70), .B(G101), .Z(n359) );
  AND2_X1 U485 ( .A1(n382), .A2(n543), .ZN(n360) );
  XOR2_X1 U486 ( .A(n558), .B(n557), .Z(n361) );
  AND2_X1 U487 ( .A1(n417), .A2(n440), .ZN(n362) );
  AND2_X1 U488 ( .A1(n377), .A2(n374), .ZN(n363) );
  XNOR2_X1 U489 ( .A(n574), .B(KEYINPUT33), .ZN(n364) );
  INV_X1 U490 ( .A(n485), .ZN(n630) );
  XNOR2_X1 U491 ( .A(G902), .B(KEYINPUT15), .ZN(n485) );
  XNOR2_X2 U492 ( .A(n365), .B(KEYINPUT45), .ZN(n743) );
  XNOR2_X1 U493 ( .A(n710), .B(KEYINPUT76), .ZN(n539) );
  XNOR2_X1 U494 ( .A(n519), .B(KEYINPUT104), .ZN(n680) );
  NOR2_X1 U495 ( .A1(n683), .A2(n398), .ZN(n397) );
  NAND2_X2 U496 ( .A1(n385), .A2(n570), .ZN(n756) );
  XNOR2_X1 U497 ( .A(n545), .B(n389), .ZN(n388) );
  NOR2_X1 U498 ( .A1(n679), .A2(KEYINPUT105), .ZN(n379) );
  NAND2_X1 U499 ( .A1(n363), .A2(n371), .ZN(n381) );
  NAND2_X1 U500 ( .A1(n666), .A2(n375), .ZN(n374) );
  NAND2_X1 U501 ( .A1(n379), .A2(n378), .ZN(n377) );
  INV_X1 U502 ( .A(n666), .ZN(n378) );
  INV_X1 U503 ( .A(n764), .ZN(n380) );
  INV_X1 U504 ( .A(n383), .ZN(n382) );
  XNOR2_X1 U505 ( .A(n383), .B(G125), .ZN(n765) );
  XNOR2_X1 U506 ( .A(n529), .B(KEYINPUT114), .ZN(n383) );
  NAND2_X1 U507 ( .A1(n361), .A2(n388), .ZN(n387) );
  NAND2_X1 U508 ( .A1(n608), .A2(n390), .ZN(n562) );
  XNOR2_X1 U509 ( .A(n587), .B(n525), .ZN(n608) );
  XNOR2_X2 U510 ( .A(n514), .B(G472), .ZN(n587) );
  NAND2_X1 U511 ( .A1(n393), .A2(n392), .ZN(n585) );
  NAND2_X1 U512 ( .A1(n683), .A2(KEYINPUT34), .ZN(n392) );
  NOR2_X1 U513 ( .A1(n397), .A2(n394), .ZN(n393) );
  NAND2_X1 U514 ( .A1(n592), .A2(KEYINPUT34), .ZN(n396) );
  XNOR2_X2 U515 ( .A(n435), .B(n364), .ZN(n683) );
  XNOR2_X1 U516 ( .A(n526), .B(n401), .ZN(n528) );
  NAND2_X1 U517 ( .A1(n420), .A2(n419), .ZN(n402) );
  NAND2_X1 U518 ( .A1(n652), .A2(n501), .ZN(n407) );
  XNOR2_X2 U519 ( .A(n487), .B(n408), .ZN(n600) );
  XNOR2_X2 U520 ( .A(n416), .B(KEYINPUT19), .ZN(n581) );
  NOR2_X1 U521 ( .A1(n562), .A2(n416), .ZN(n526) );
  NAND2_X1 U522 ( .A1(n593), .A2(n417), .ZN(n594) );
  INV_X1 U523 ( .A(n756), .ZN(n423) );
  OR2_X2 U524 ( .A1(n624), .A2(n439), .ZN(n621) );
  XNOR2_X2 U525 ( .A(n430), .B(KEYINPUT91), .ZN(n624) );
  NOR2_X2 U526 ( .A1(n763), .A2(n670), .ZN(n430) );
  XNOR2_X2 U527 ( .A(n614), .B(n613), .ZN(n763) );
  NAND2_X1 U528 ( .A1(n573), .A2(n608), .ZN(n435) );
  XNOR2_X2 U529 ( .A(n599), .B(n598), .ZN(n617) );
  XNOR2_X2 U530 ( .A(n465), .B(KEYINPUT78), .ZN(n739) );
  XOR2_X2 U531 ( .A(G110), .B(G107), .Z(n465) );
  NAND2_X1 U532 ( .A1(n618), .A2(KEYINPUT90), .ZN(n439) );
  XNOR2_X1 U533 ( .A(KEYINPUT83), .B(n507), .ZN(n440) );
  XOR2_X1 U534 ( .A(KEYINPUT30), .B(n516), .Z(n441) );
  XNOR2_X1 U535 ( .A(n478), .B(n477), .ZN(n479) );
  BUF_X1 U536 ( .A(n683), .Z(n715) );
  BUF_X1 U537 ( .A(n581), .Z(n536) );
  XNOR2_X1 U538 ( .A(n555), .B(n554), .ZN(n559) );
  INV_X1 U539 ( .A(n536), .ZN(n537) );
  INV_X1 U540 ( .A(KEYINPUT125), .ZN(n636) );
  BUF_X1 U541 ( .A(n622), .Z(n638) );
  XOR2_X1 U542 ( .A(G122), .B(G104), .Z(n471) );
  XNOR2_X1 U543 ( .A(n751), .B(n471), .ZN(n450) );
  XNOR2_X1 U544 ( .A(n443), .B(n442), .ZN(n446) );
  NAND2_X1 U545 ( .A1(n508), .A2(G214), .ZN(n444) );
  XNOR2_X1 U546 ( .A(n444), .B(KEYINPUT12), .ZN(n445) );
  XNOR2_X1 U547 ( .A(n446), .B(n445), .ZN(n448) );
  XNOR2_X1 U548 ( .A(n448), .B(n492), .ZN(n449) );
  XNOR2_X1 U549 ( .A(n449), .B(n450), .ZN(n645) );
  INV_X1 U550 ( .A(G902), .ZN(n513) );
  NAND2_X1 U551 ( .A1(n645), .A2(n513), .ZN(n452) );
  XOR2_X1 U552 ( .A(KEYINPUT13), .B(G475), .Z(n451) );
  XNOR2_X1 U553 ( .A(G116), .B(G122), .ZN(n453) );
  XNOR2_X1 U554 ( .A(n453), .B(KEYINPUT7), .ZN(n457) );
  XNOR2_X1 U555 ( .A(G107), .B(KEYINPUT9), .ZN(n454) );
  XNOR2_X1 U556 ( .A(n455), .B(n454), .ZN(n456) );
  XOR2_X1 U557 ( .A(n457), .B(n456), .Z(n461) );
  NAND2_X1 U558 ( .A1(n757), .A2(G234), .ZN(n459) );
  XNOR2_X1 U559 ( .A(KEYINPUT8), .B(KEYINPUT65), .ZN(n458) );
  XNOR2_X1 U560 ( .A(n459), .B(n458), .ZN(n480) );
  NAND2_X1 U561 ( .A1(G217), .A2(n480), .ZN(n460) );
  XNOR2_X1 U562 ( .A(n461), .B(n460), .ZN(n462) );
  XNOR2_X1 U563 ( .A(n494), .B(n462), .ZN(n736) );
  NAND2_X1 U564 ( .A1(n736), .A2(n513), .ZN(n463) );
  NAND2_X1 U565 ( .A1(n548), .A2(n547), .ZN(n583) );
  XNOR2_X1 U566 ( .A(KEYINPUT3), .B(KEYINPUT69), .ZN(n466) );
  XNOR2_X1 U567 ( .A(n359), .B(n466), .ZN(n470) );
  XNOR2_X1 U568 ( .A(G119), .B(G116), .ZN(n468) );
  XNOR2_X1 U569 ( .A(n468), .B(n467), .ZN(n469) );
  NAND2_X1 U570 ( .A1(n659), .A2(n485), .ZN(n474) );
  AND2_X1 U571 ( .A1(G210), .A2(n515), .ZN(n473) );
  INV_X1 U572 ( .A(n568), .ZN(n546) );
  XOR2_X1 U573 ( .A(KEYINPUT98), .B(KEYINPUT97), .Z(n476) );
  XNOR2_X1 U574 ( .A(n476), .B(n475), .ZN(n478) );
  AND2_X1 U575 ( .A1(n480), .A2(G221), .ZN(n482) );
  XNOR2_X1 U576 ( .A(n482), .B(n481), .ZN(n483) );
  XNOR2_X1 U577 ( .A(n484), .B(n483), .ZN(n631) );
  NAND2_X1 U578 ( .A1(n631), .A2(n513), .ZN(n487) );
  NAND2_X1 U579 ( .A1(G234), .A2(n485), .ZN(n486) );
  XNOR2_X1 U580 ( .A(KEYINPUT20), .B(n486), .ZN(n488) );
  NAND2_X1 U581 ( .A1(n488), .A2(G221), .ZN(n490) );
  XOR2_X1 U582 ( .A(KEYINPUT21), .B(KEYINPUT100), .Z(n489) );
  XNOR2_X1 U583 ( .A(n490), .B(n489), .ZN(n689) );
  NAND2_X1 U584 ( .A1(n600), .A2(n689), .ZN(n686) );
  XNOR2_X1 U585 ( .A(KEYINPUT4), .B(G137), .ZN(n491) );
  XNOR2_X1 U586 ( .A(n492), .B(n491), .ZN(n493) );
  NAND2_X1 U587 ( .A1(n757), .A2(G227), .ZN(n495) );
  XNOR2_X1 U588 ( .A(n495), .B(G101), .ZN(n497) );
  XNOR2_X1 U589 ( .A(G140), .B(G104), .ZN(n496) );
  XNOR2_X1 U590 ( .A(n497), .B(n496), .ZN(n498) );
  XNOR2_X1 U591 ( .A(n499), .B(n498), .ZN(n500) );
  INV_X1 U592 ( .A(G469), .ZN(n501) );
  NAND2_X1 U593 ( .A1(G237), .A2(G234), .ZN(n502) );
  XNOR2_X1 U594 ( .A(n502), .B(KEYINPUT14), .ZN(n503) );
  NAND2_X1 U595 ( .A1(G952), .A2(n503), .ZN(n721) );
  NOR2_X1 U596 ( .A1(G953), .A2(n721), .ZN(n575) );
  NAND2_X1 U597 ( .A1(n503), .A2(G902), .ZN(n504) );
  XOR2_X1 U598 ( .A(KEYINPUT94), .B(n504), .Z(n576) );
  NAND2_X1 U599 ( .A1(n576), .A2(G953), .ZN(n505) );
  NOR2_X1 U600 ( .A1(G900), .A2(n505), .ZN(n506) );
  NOR2_X1 U601 ( .A1(n575), .A2(n506), .ZN(n507) );
  NAND2_X1 U602 ( .A1(n508), .A2(G210), .ZN(n509) );
  XNOR2_X1 U603 ( .A(n509), .B(KEYINPUT5), .ZN(n510) );
  XNOR2_X1 U604 ( .A(n511), .B(n510), .ZN(n512) );
  NAND2_X1 U605 ( .A1(n639), .A2(n513), .ZN(n514) );
  NAND2_X1 U606 ( .A1(G214), .A2(n515), .ZN(n707) );
  NAND2_X1 U607 ( .A1(n587), .A2(n707), .ZN(n516) );
  NAND2_X1 U608 ( .A1(n362), .A2(n441), .ZN(n552) );
  NOR2_X1 U609 ( .A1(n546), .A2(n552), .ZN(n517) );
  XNOR2_X1 U610 ( .A(n517), .B(KEYINPUT109), .ZN(n518) );
  NOR2_X2 U611 ( .A1(n583), .A2(n518), .ZN(n673) );
  XNOR2_X1 U612 ( .A(n673), .B(KEYINPUT87), .ZN(n522) );
  INV_X1 U613 ( .A(n548), .ZN(n520) );
  AND2_X1 U614 ( .A1(n520), .A2(n547), .ZN(n519) );
  NOR2_X1 U615 ( .A1(n520), .A2(n547), .ZN(n677) );
  NOR2_X1 U616 ( .A1(n680), .A2(n677), .ZN(n710) );
  NAND2_X1 U617 ( .A1(n710), .A2(KEYINPUT47), .ZN(n521) );
  NAND2_X1 U618 ( .A1(n522), .A2(n521), .ZN(n523) );
  XNOR2_X1 U619 ( .A(n523), .B(KEYINPUT85), .ZN(n544) );
  NAND2_X1 U620 ( .A1(n689), .A2(n440), .ZN(n524) );
  NOR2_X1 U621 ( .A1(n600), .A2(n524), .ZN(n530) );
  INV_X1 U622 ( .A(KEYINPUT6), .ZN(n525) );
  BUF_X2 U623 ( .A(n571), .Z(n687) );
  NOR2_X1 U624 ( .A1(n528), .A2(n687), .ZN(n529) );
  NAND2_X1 U625 ( .A1(n530), .A2(n587), .ZN(n531) );
  XNOR2_X1 U626 ( .A(n531), .B(KEYINPUT111), .ZN(n532) );
  XNOR2_X1 U627 ( .A(KEYINPUT28), .B(n532), .ZN(n535) );
  XOR2_X1 U628 ( .A(KEYINPUT110), .B(n533), .Z(n534) );
  NAND2_X1 U629 ( .A1(n535), .A2(n534), .ZN(n551) );
  NOR2_X1 U630 ( .A1(n551), .A2(n537), .ZN(n675) );
  NAND2_X1 U631 ( .A1(KEYINPUT76), .A2(n675), .ZN(n538) );
  NAND2_X1 U632 ( .A1(n538), .A2(KEYINPUT47), .ZN(n542) );
  NOR2_X1 U633 ( .A1(KEYINPUT47), .A2(n539), .ZN(n540) );
  NAND2_X1 U634 ( .A1(n540), .A2(n675), .ZN(n541) );
  AND2_X1 U635 ( .A1(n541), .A2(n542), .ZN(n543) );
  NAND2_X1 U636 ( .A1(n544), .A2(n360), .ZN(n545) );
  XNOR2_X1 U637 ( .A(KEYINPUT38), .B(n546), .ZN(n708) );
  NOR2_X1 U638 ( .A1(n548), .A2(n547), .ZN(n704) );
  AND2_X1 U639 ( .A1(n707), .A2(n704), .ZN(n549) );
  AND2_X1 U640 ( .A1(n708), .A2(n549), .ZN(n550) );
  XNOR2_X1 U641 ( .A(KEYINPUT41), .B(n550), .ZN(n703) );
  XOR2_X1 U642 ( .A(KEYINPUT73), .B(KEYINPUT39), .Z(n555) );
  INV_X1 U643 ( .A(n552), .ZN(n553) );
  NAND2_X1 U644 ( .A1(n553), .A2(n708), .ZN(n554) );
  INV_X1 U645 ( .A(KEYINPUT88), .ZN(n556) );
  NAND2_X1 U646 ( .A1(n680), .A2(n559), .ZN(n561) );
  INV_X1 U647 ( .A(KEYINPUT115), .ZN(n560) );
  XNOR2_X1 U648 ( .A(n561), .B(n560), .ZN(n761) );
  INV_X1 U649 ( .A(n761), .ZN(n569) );
  INV_X1 U650 ( .A(n562), .ZN(n563) );
  NAND2_X1 U651 ( .A1(n563), .A2(n707), .ZN(n565) );
  INV_X1 U652 ( .A(n687), .ZN(n564) );
  NOR2_X1 U653 ( .A1(n565), .A2(n564), .ZN(n566) );
  XNOR2_X1 U654 ( .A(n566), .B(KEYINPUT43), .ZN(n567) );
  NOR2_X1 U655 ( .A1(n568), .A2(n567), .ZN(n682) );
  NOR2_X1 U656 ( .A1(n569), .A2(n682), .ZN(n570) );
  NOR2_X2 U657 ( .A1(n571), .A2(n686), .ZN(n572) );
  XNOR2_X2 U658 ( .A(n572), .B(KEYINPUT77), .ZN(n588) );
  XNOR2_X1 U659 ( .A(n588), .B(KEYINPUT107), .ZN(n573) );
  INV_X1 U660 ( .A(KEYINPUT108), .ZN(n574) );
  INV_X1 U661 ( .A(n575), .ZN(n578) );
  NOR2_X1 U662 ( .A1(G898), .A2(n757), .ZN(n741) );
  NAND2_X1 U663 ( .A1(n741), .A2(n576), .ZN(n577) );
  NAND2_X1 U664 ( .A1(n578), .A2(n577), .ZN(n579) );
  XOR2_X1 U665 ( .A(KEYINPUT95), .B(n579), .Z(n580) );
  NAND2_X1 U666 ( .A1(n581), .A2(n580), .ZN(n582) );
  XNOR2_X2 U667 ( .A(n582), .B(KEYINPUT0), .ZN(n596) );
  XNOR2_X1 U668 ( .A(n596), .B(KEYINPUT96), .ZN(n592) );
  INV_X1 U669 ( .A(KEYINPUT35), .ZN(n584) );
  XNOR2_X1 U670 ( .A(n585), .B(n584), .ZN(n622) );
  INV_X1 U671 ( .A(n622), .ZN(n586) );
  NAND2_X1 U672 ( .A1(n586), .A2(KEYINPUT44), .ZN(n606) );
  INV_X1 U673 ( .A(n587), .ZN(n694) );
  NOR2_X1 U674 ( .A1(n596), .A2(n694), .ZN(n590) );
  INV_X1 U675 ( .A(n697), .ZN(n589) );
  NAND2_X1 U676 ( .A1(n590), .A2(n589), .ZN(n591) );
  XNOR2_X1 U677 ( .A(n591), .B(KEYINPUT31), .ZN(n679) );
  INV_X1 U678 ( .A(n694), .ZN(n696) );
  INV_X1 U679 ( .A(n592), .ZN(n593) );
  NAND2_X1 U680 ( .A1(n704), .A2(n689), .ZN(n595) );
  NOR2_X2 U681 ( .A1(n596), .A2(n595), .ZN(n599) );
  XOR2_X1 U682 ( .A(KEYINPUT22), .B(KEYINPUT74), .Z(n597) );
  XNOR2_X1 U683 ( .A(KEYINPUT75), .B(n597), .ZN(n598) );
  NAND2_X1 U684 ( .A1(n687), .A2(n600), .ZN(n601) );
  NOR2_X1 U685 ( .A1(n608), .A2(n601), .ZN(n602) );
  NAND2_X1 U686 ( .A1(n617), .A2(n602), .ZN(n604) );
  INV_X1 U687 ( .A(KEYINPUT106), .ZN(n603) );
  XNOR2_X1 U688 ( .A(n604), .B(n603), .ZN(n764) );
  NAND2_X1 U689 ( .A1(n606), .A2(n605), .ZN(n607) );
  INV_X1 U690 ( .A(n608), .ZN(n610) );
  NOR2_X1 U691 ( .A1(n687), .A2(n600), .ZN(n609) );
  NAND2_X1 U692 ( .A1(n610), .A2(n609), .ZN(n611) );
  XNOR2_X1 U693 ( .A(KEYINPUT81), .B(n611), .ZN(n612) );
  NAND2_X1 U694 ( .A1(n617), .A2(n612), .ZN(n614) );
  XOR2_X1 U695 ( .A(KEYINPUT64), .B(KEYINPUT32), .Z(n613) );
  NOR2_X1 U696 ( .A1(n600), .A2(n696), .ZN(n615) );
  AND2_X1 U697 ( .A1(n615), .A2(n687), .ZN(n616) );
  AND2_X1 U698 ( .A1(n617), .A2(n616), .ZN(n670) );
  INV_X1 U699 ( .A(KEYINPUT44), .ZN(n618) );
  INV_X1 U700 ( .A(KEYINPUT90), .ZN(n619) );
  NAND2_X1 U701 ( .A1(n624), .A2(n619), .ZN(n620) );
  NAND2_X1 U702 ( .A1(n621), .A2(n620), .ZN(n623) );
  NAND2_X1 U703 ( .A1(n623), .A2(n638), .ZN(n626) );
  NAND2_X1 U704 ( .A1(n624), .A2(KEYINPUT44), .ZN(n625) );
  INV_X1 U705 ( .A(KEYINPUT2), .ZN(n629) );
  NAND2_X1 U706 ( .A1(n734), .A2(G217), .ZN(n633) );
  INV_X1 U707 ( .A(n631), .ZN(n632) );
  XNOR2_X1 U708 ( .A(n633), .B(n632), .ZN(n635) );
  INV_X1 U709 ( .A(G952), .ZN(n634) );
  NOR2_X2 U710 ( .A1(n635), .A2(n738), .ZN(n637) );
  XNOR2_X1 U711 ( .A(n637), .B(n636), .ZN(G66) );
  XNOR2_X1 U712 ( .A(n638), .B(G122), .ZN(G24) );
  NAND2_X1 U713 ( .A1(n734), .A2(G472), .ZN(n641) );
  XOR2_X1 U714 ( .A(KEYINPUT92), .B(KEYINPUT63), .Z(n643) );
  XNOR2_X1 U715 ( .A(n644), .B(n643), .ZN(G57) );
  NAND2_X1 U716 ( .A1(n734), .A2(G475), .ZN(n647) );
  XNOR2_X1 U717 ( .A(KEYINPUT124), .B(KEYINPUT60), .ZN(n649) );
  XNOR2_X1 U718 ( .A(n650), .B(n649), .ZN(G60) );
  NAND2_X1 U719 ( .A1(n734), .A2(G469), .ZN(n654) );
  XNOR2_X1 U720 ( .A(KEYINPUT57), .B(KEYINPUT58), .ZN(n651) );
  XNOR2_X1 U721 ( .A(n652), .B(n651), .ZN(n653) );
  XNOR2_X1 U722 ( .A(n654), .B(n653), .ZN(n656) );
  INV_X1 U723 ( .A(n738), .ZN(n655) );
  AND2_X1 U724 ( .A1(n656), .A2(n655), .ZN(G54) );
  NAND2_X1 U725 ( .A1(n734), .A2(G210), .ZN(n661) );
  XNOR2_X1 U726 ( .A(KEYINPUT86), .B(KEYINPUT54), .ZN(n657) );
  XNOR2_X1 U727 ( .A(n657), .B(KEYINPUT55), .ZN(n658) );
  XNOR2_X1 U728 ( .A(n659), .B(n658), .ZN(n660) );
  XNOR2_X1 U729 ( .A(n663), .B(KEYINPUT56), .ZN(G51) );
  NAND2_X1 U730 ( .A1(n666), .A2(n677), .ZN(n664) );
  XNOR2_X1 U731 ( .A(n664), .B(KEYINPUT116), .ZN(n665) );
  XNOR2_X1 U732 ( .A(G104), .B(n665), .ZN(G6) );
  XOR2_X1 U733 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n668) );
  NAND2_X1 U734 ( .A1(n666), .A2(n680), .ZN(n667) );
  XNOR2_X1 U735 ( .A(n668), .B(n667), .ZN(n669) );
  XNOR2_X1 U736 ( .A(G107), .B(n669), .ZN(G9) );
  XOR2_X1 U737 ( .A(n670), .B(G110), .Z(G12) );
  XOR2_X1 U738 ( .A(G128), .B(KEYINPUT29), .Z(n672) );
  NAND2_X1 U739 ( .A1(n675), .A2(n680), .ZN(n671) );
  XNOR2_X1 U740 ( .A(n672), .B(n671), .ZN(G30) );
  XNOR2_X1 U741 ( .A(n673), .B(G143), .ZN(n674) );
  XNOR2_X1 U742 ( .A(n674), .B(KEYINPUT117), .ZN(G45) );
  NAND2_X1 U743 ( .A1(n675), .A2(n677), .ZN(n676) );
  XNOR2_X1 U744 ( .A(n676), .B(G146), .ZN(G48) );
  NAND2_X1 U745 ( .A1(n679), .A2(n677), .ZN(n678) );
  XNOR2_X1 U746 ( .A(n678), .B(G113), .ZN(G15) );
  NAND2_X1 U747 ( .A1(n680), .A2(n679), .ZN(n681) );
  XNOR2_X1 U748 ( .A(n681), .B(G116), .ZN(G18) );
  XOR2_X1 U749 ( .A(G140), .B(n682), .Z(G42) );
  NOR2_X1 U750 ( .A1(n715), .A2(n703), .ZN(n684) );
  XNOR2_X1 U751 ( .A(n684), .B(KEYINPUT123), .ZN(n685) );
  NAND2_X1 U752 ( .A1(n757), .A2(n685), .ZN(n724) );
  XOR2_X1 U753 ( .A(KEYINPUT122), .B(KEYINPUT121), .Z(n720) );
  NAND2_X1 U754 ( .A1(n687), .A2(n686), .ZN(n688) );
  XNOR2_X1 U755 ( .A(n688), .B(KEYINPUT50), .ZN(n693) );
  NOR2_X1 U756 ( .A1(n689), .A2(n600), .ZN(n691) );
  XNOR2_X1 U757 ( .A(KEYINPUT49), .B(KEYINPUT118), .ZN(n690) );
  XNOR2_X1 U758 ( .A(n691), .B(n690), .ZN(n692) );
  NAND2_X1 U759 ( .A1(n693), .A2(n692), .ZN(n695) );
  NAND2_X1 U760 ( .A1(n695), .A2(n694), .ZN(n699) );
  NAND2_X1 U761 ( .A1(n697), .A2(n696), .ZN(n698) );
  NAND2_X1 U762 ( .A1(n699), .A2(n698), .ZN(n700) );
  XNOR2_X1 U763 ( .A(n700), .B(KEYINPUT119), .ZN(n701) );
  XNOR2_X1 U764 ( .A(n701), .B(KEYINPUT51), .ZN(n702) );
  NOR2_X1 U765 ( .A1(n703), .A2(n702), .ZN(n717) );
  INV_X1 U766 ( .A(n704), .ZN(n706) );
  NOR2_X1 U767 ( .A1(n708), .A2(n707), .ZN(n705) );
  NOR2_X1 U768 ( .A1(n706), .A2(n705), .ZN(n712) );
  NAND2_X1 U769 ( .A1(n708), .A2(n707), .ZN(n709) );
  NOR2_X1 U770 ( .A1(n710), .A2(n709), .ZN(n711) );
  NOR2_X1 U771 ( .A1(n712), .A2(n711), .ZN(n713) );
  XNOR2_X1 U772 ( .A(n713), .B(KEYINPUT120), .ZN(n714) );
  NOR2_X1 U773 ( .A1(n715), .A2(n714), .ZN(n716) );
  NOR2_X1 U774 ( .A1(n717), .A2(n716), .ZN(n718) );
  XNOR2_X1 U775 ( .A(n718), .B(KEYINPUT52), .ZN(n719) );
  XNOR2_X1 U776 ( .A(n720), .B(n719), .ZN(n722) );
  NOR2_X1 U777 ( .A1(n722), .A2(n721), .ZN(n723) );
  NOR2_X1 U778 ( .A1(n724), .A2(n723), .ZN(n728) );
  INV_X1 U779 ( .A(KEYINPUT84), .ZN(n725) );
  OR2_X1 U780 ( .A1(n726), .A2(n725), .ZN(n727) );
  NAND2_X1 U781 ( .A1(n728), .A2(n727), .ZN(n732) );
  XNOR2_X1 U782 ( .A(n729), .B(KEYINPUT84), .ZN(n730) );
  NOR2_X1 U783 ( .A1(n730), .A2(KEYINPUT2), .ZN(n731) );
  NOR2_X1 U784 ( .A1(n732), .A2(n731), .ZN(n733) );
  XNOR2_X1 U785 ( .A(n733), .B(KEYINPUT53), .ZN(G75) );
  NAND2_X1 U786 ( .A1(n734), .A2(G478), .ZN(n735) );
  XOR2_X1 U787 ( .A(n736), .B(n735), .Z(n737) );
  NOR2_X1 U788 ( .A1(n738), .A2(n737), .ZN(G63) );
  XNOR2_X1 U789 ( .A(n740), .B(n739), .ZN(n742) );
  NOR2_X1 U790 ( .A1(n742), .A2(n741), .ZN(n749) );
  NAND2_X1 U791 ( .A1(n743), .A2(n757), .ZN(n747) );
  NAND2_X1 U792 ( .A1(G953), .A2(G224), .ZN(n744) );
  XNOR2_X1 U793 ( .A(KEYINPUT61), .B(n744), .ZN(n745) );
  NAND2_X1 U794 ( .A1(n745), .A2(G898), .ZN(n746) );
  NAND2_X1 U795 ( .A1(n747), .A2(n746), .ZN(n748) );
  XNOR2_X1 U796 ( .A(n749), .B(n748), .ZN(G69) );
  XNOR2_X1 U797 ( .A(n750), .B(n751), .ZN(n755) );
  XNOR2_X1 U798 ( .A(n755), .B(G227), .ZN(n752) );
  NAND2_X1 U799 ( .A1(n752), .A2(G900), .ZN(n753) );
  NAND2_X1 U800 ( .A1(n753), .A2(G953), .ZN(n754) );
  XNOR2_X1 U801 ( .A(n754), .B(KEYINPUT126), .ZN(n760) );
  XNOR2_X1 U802 ( .A(n756), .B(n755), .ZN(n758) );
  NAND2_X1 U803 ( .A1(n758), .A2(n757), .ZN(n759) );
  NAND2_X1 U804 ( .A1(n760), .A2(n759), .ZN(G72) );
  XNOR2_X1 U805 ( .A(G134), .B(n761), .ZN(G36) );
  XNOR2_X1 U806 ( .A(G131), .B(n762), .ZN(G33) );
  XOR2_X1 U807 ( .A(n763), .B(G119), .Z(G21) );
  XOR2_X1 U808 ( .A(G101), .B(n764), .Z(G3) );
  XNOR2_X1 U809 ( .A(KEYINPUT37), .B(n765), .ZN(G27) );
  XNOR2_X1 U810 ( .A(G137), .B(n766), .ZN(G39) );
endmodule

