

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
         n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597,
         n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608,
         n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619,
         n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630,
         n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641,
         n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652,
         n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663,
         n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674,
         n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685,
         n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696,
         n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707,
         n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718,
         n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729,
         n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740,
         n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751,
         n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762,
         n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773,
         n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784,
         n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, n795,
         n796, n797, n798, n799, n800, n801, n802, n803, n804, n805, n806,
         n807, n808, n809, n810, n811, n812, n813, n814, n815, n816, n817,
         n818, n819, n820, n821, n822, n823, n824, n825, n826, n827, n828,
         n829, n830, n831, n832, n833, n834, n835, n836, n837, n838, n839,
         n840, n841, n842, n843, n844, n845, n846, n847, n848, n849, n850,
         n851, n852, n853, n854, n855, n856, n857, n858, n859, n860, n861,
         n862, n863, n864, n865, n866, n867, n868, n869, n870, n871, n872,
         n873, n874, n875, n876, n877, n878, n879, n880, n881, n882, n883,
         n884, n885, n886, n887, n888, n889, n890, n891, n892, n893, n894,
         n895, n896, n897, n898, n899, n900, n901, n902, n903, n904, n905,
         n906, n907, n908, n909, n910, n911, n912, n913, n914, n915, n916,
         n917, n918, n919, n920, n921, n922, n923, n924, n925, n926, n927,
         n928, n929, n930, n931, n932, n933, n934, n935, n936, n937, n938,
         n939, n940, n941, n942, n943, n944, n945, n946, n947, n948, n949,
         n950, n951, n952, n953, n954, n955, n956, n957, n958, n959, n960,
         n961, n962, n963, n964, n965, n966, n967, n968, n969, n970, n971,
         n972, n973, n974, n975, n976, n977, n978, n979, n980, n981, n982,
         n983, n984, n985, n986, n987, n988, n989, n990, n991, n992, n993,
         n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
         n1025, n1026, n1027, n1028, n1029;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  AND2_X1 U552 ( .A1(G2105), .A2(G2104), .ZN(n881) );
  AND2_X1 U553 ( .A1(n740), .A2(n739), .ZN(n742) );
  XNOR2_X2 U554 ( .A(n742), .B(n741), .ZN(n766) );
  XNOR2_X1 U555 ( .A(n532), .B(KEYINPUT65), .ZN(n648) );
  INV_X1 U556 ( .A(G2105), .ZN(n525) );
  XNOR2_X1 U557 ( .A(G543), .B(KEYINPUT0), .ZN(n532) );
  XNOR2_X1 U558 ( .A(n715), .B(n517), .ZN(n719) );
  NOR2_X1 U559 ( .A1(n727), .A2(n726), .ZN(n729) );
  NOR2_X1 U560 ( .A1(n820), .A2(n811), .ZN(n812) );
  NOR2_X1 U561 ( .A1(G543), .A2(n538), .ZN(n539) );
  NOR2_X1 U562 ( .A1(n546), .A2(n545), .ZN(n547) );
  XOR2_X1 U563 ( .A(KEYINPUT29), .B(KEYINPUT100), .Z(n517) );
  OR2_X1 U564 ( .A1(G301), .A2(n720), .ZN(n518) );
  AND2_X1 U565 ( .A1(n744), .A2(G8), .ZN(n519) );
  XOR2_X1 U566 ( .A(n729), .B(n728), .Z(n520) );
  XNOR2_X1 U567 ( .A(KEYINPUT102), .B(KEYINPUT31), .ZN(n728) );
  OR2_X2 U568 ( .A1(n795), .A2(n797), .ZN(n722) );
  OR2_X1 U569 ( .A1(G1384), .A2(G164), .ZN(n690) );
  NOR2_X1 U570 ( .A1(n777), .A2(n776), .ZN(n778) );
  INV_X1 U571 ( .A(KEYINPUT77), .ZN(n592) );
  XNOR2_X1 U572 ( .A(n690), .B(KEYINPUT64), .ZN(n795) );
  NAND2_X1 U573 ( .A1(n813), .A2(n812), .ZN(n814) );
  INV_X1 U574 ( .A(KEYINPUT15), .ZN(n598) );
  NOR2_X1 U575 ( .A1(G2105), .A2(G2104), .ZN(n528) );
  NOR2_X2 U576 ( .A1(n648), .A2(n538), .ZN(n655) );
  NOR2_X2 U577 ( .A1(G2104), .A2(n525), .ZN(n882) );
  NOR2_X2 U578 ( .A1(G651), .A2(n648), .ZN(n654) );
  AND2_X4 U579 ( .A1(n525), .A2(G2104), .ZN(n877) );
  NAND2_X1 U580 ( .A1(G102), .A2(n877), .ZN(n521) );
  XOR2_X1 U581 ( .A(KEYINPUT92), .B(n521), .Z(n524) );
  NAND2_X1 U582 ( .A1(G114), .A2(n881), .ZN(n522) );
  XNOR2_X1 U583 ( .A(KEYINPUT91), .B(n522), .ZN(n523) );
  NOR2_X1 U584 ( .A1(n524), .A2(n523), .ZN(n527) );
  NAND2_X1 U585 ( .A1(n882), .A2(G126), .ZN(n526) );
  NAND2_X1 U586 ( .A1(n527), .A2(n526), .ZN(n531) );
  XOR2_X1 U587 ( .A(KEYINPUT17), .B(n528), .Z(n558) );
  NAND2_X1 U588 ( .A1(G138), .A2(n558), .ZN(n529) );
  XNOR2_X1 U589 ( .A(n529), .B(KEYINPUT93), .ZN(n530) );
  NOR2_X2 U590 ( .A1(n531), .A2(n530), .ZN(G164) );
  AND2_X1 U591 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U592 ( .A(G860), .ZN(n613) );
  INV_X1 U593 ( .A(G651), .ZN(n538) );
  NAND2_X1 U594 ( .A1(n655), .A2(G68), .ZN(n533) );
  XNOR2_X1 U595 ( .A(KEYINPUT72), .B(n533), .ZN(n536) );
  NOR2_X1 U596 ( .A1(G543), .A2(G651), .ZN(n656) );
  NAND2_X1 U597 ( .A1(n656), .A2(G81), .ZN(n534) );
  XNOR2_X1 U598 ( .A(KEYINPUT12), .B(n534), .ZN(n535) );
  NAND2_X1 U599 ( .A1(n536), .A2(n535), .ZN(n537) );
  XNOR2_X1 U600 ( .A(n537), .B(KEYINPUT13), .ZN(n543) );
  XOR2_X1 U601 ( .A(KEYINPUT1), .B(n539), .Z(n659) );
  NAND2_X1 U602 ( .A1(n659), .A2(G56), .ZN(n541) );
  XOR2_X1 U603 ( .A(KEYINPUT14), .B(KEYINPUT71), .Z(n540) );
  XNOR2_X1 U604 ( .A(n541), .B(n540), .ZN(n542) );
  NAND2_X1 U605 ( .A1(n543), .A2(n542), .ZN(n546) );
  NAND2_X1 U606 ( .A1(G43), .A2(n654), .ZN(n544) );
  XNOR2_X1 U607 ( .A(KEYINPUT73), .B(n544), .ZN(n545) );
  XOR2_X2 U608 ( .A(KEYINPUT74), .B(n547), .Z(n973) );
  OR2_X1 U609 ( .A1(n613), .A2(n973), .ZN(G153) );
  INV_X1 U610 ( .A(G132), .ZN(G219) );
  INV_X1 U611 ( .A(G82), .ZN(G220) );
  INV_X1 U612 ( .A(G57), .ZN(G237) );
  NAND2_X1 U613 ( .A1(n656), .A2(G88), .ZN(n550) );
  NAND2_X1 U614 ( .A1(G62), .A2(n659), .ZN(n548) );
  XOR2_X1 U615 ( .A(KEYINPUT89), .B(n548), .Z(n549) );
  NAND2_X1 U616 ( .A1(n550), .A2(n549), .ZN(n554) );
  NAND2_X1 U617 ( .A1(G75), .A2(n655), .ZN(n552) );
  NAND2_X1 U618 ( .A1(G50), .A2(n654), .ZN(n551) );
  NAND2_X1 U619 ( .A1(n552), .A2(n551), .ZN(n553) );
  NOR2_X1 U620 ( .A1(n554), .A2(n553), .ZN(G166) );
  NAND2_X1 U621 ( .A1(n881), .A2(G113), .ZN(n557) );
  NAND2_X1 U622 ( .A1(G101), .A2(n877), .ZN(n555) );
  XOR2_X1 U623 ( .A(KEYINPUT23), .B(n555), .Z(n556) );
  NAND2_X1 U624 ( .A1(n557), .A2(n556), .ZN(n563) );
  INV_X1 U625 ( .A(n558), .ZN(n559) );
  INV_X1 U626 ( .A(n559), .ZN(n878) );
  NAND2_X1 U627 ( .A1(G137), .A2(n878), .ZN(n561) );
  NAND2_X1 U628 ( .A1(G125), .A2(n882), .ZN(n560) );
  NAND2_X1 U629 ( .A1(n561), .A2(n560), .ZN(n562) );
  NOR2_X1 U630 ( .A1(n563), .A2(n562), .ZN(G160) );
  NAND2_X1 U631 ( .A1(G51), .A2(n654), .ZN(n565) );
  NAND2_X1 U632 ( .A1(G63), .A2(n659), .ZN(n564) );
  NAND2_X1 U633 ( .A1(n565), .A2(n564), .ZN(n566) );
  XNOR2_X1 U634 ( .A(KEYINPUT6), .B(n566), .ZN(n573) );
  NAND2_X1 U635 ( .A1(n656), .A2(G89), .ZN(n567) );
  XNOR2_X1 U636 ( .A(n567), .B(KEYINPUT4), .ZN(n569) );
  NAND2_X1 U637 ( .A1(G76), .A2(n655), .ZN(n568) );
  NAND2_X1 U638 ( .A1(n569), .A2(n568), .ZN(n570) );
  XOR2_X1 U639 ( .A(KEYINPUT5), .B(n570), .Z(n571) );
  XNOR2_X1 U640 ( .A(KEYINPUT80), .B(n571), .ZN(n572) );
  NOR2_X1 U641 ( .A1(n573), .A2(n572), .ZN(n574) );
  XOR2_X1 U642 ( .A(KEYINPUT7), .B(n574), .Z(G168) );
  XNOR2_X1 U643 ( .A(G168), .B(KEYINPUT8), .ZN(n575) );
  XNOR2_X1 U644 ( .A(n575), .B(KEYINPUT81), .ZN(G286) );
  XOR2_X1 U645 ( .A(KEYINPUT10), .B(KEYINPUT69), .Z(n577) );
  NAND2_X1 U646 ( .A1(G7), .A2(G661), .ZN(n576) );
  XNOR2_X1 U647 ( .A(n577), .B(n576), .ZN(G223) );
  XOR2_X1 U648 ( .A(KEYINPUT11), .B(KEYINPUT70), .Z(n579) );
  INV_X1 U649 ( .A(G223), .ZN(n833) );
  NAND2_X1 U650 ( .A1(G567), .A2(n833), .ZN(n578) );
  XNOR2_X1 U651 ( .A(n579), .B(n578), .ZN(G234) );
  NAND2_X1 U652 ( .A1(n656), .A2(G90), .ZN(n580) );
  XNOR2_X1 U653 ( .A(n580), .B(KEYINPUT68), .ZN(n582) );
  NAND2_X1 U654 ( .A1(G77), .A2(n655), .ZN(n581) );
  NAND2_X1 U655 ( .A1(n582), .A2(n581), .ZN(n583) );
  XNOR2_X1 U656 ( .A(KEYINPUT9), .B(n583), .ZN(n587) );
  NAND2_X1 U657 ( .A1(n654), .A2(G52), .ZN(n585) );
  NAND2_X1 U658 ( .A1(G64), .A2(n659), .ZN(n584) );
  AND2_X1 U659 ( .A1(n585), .A2(n584), .ZN(n586) );
  NAND2_X1 U660 ( .A1(n587), .A2(n586), .ZN(G301) );
  NAND2_X1 U661 ( .A1(G868), .A2(G301), .ZN(n588) );
  XNOR2_X1 U662 ( .A(n588), .B(KEYINPUT75), .ZN(n602) );
  NAND2_X1 U663 ( .A1(n654), .A2(G54), .ZN(n589) );
  XNOR2_X1 U664 ( .A(n589), .B(KEYINPUT76), .ZN(n591) );
  NAND2_X1 U665 ( .A1(G79), .A2(n655), .ZN(n590) );
  NAND2_X1 U666 ( .A1(n591), .A2(n590), .ZN(n593) );
  XNOR2_X1 U667 ( .A(n593), .B(n592), .ZN(n597) );
  NAND2_X1 U668 ( .A1(G92), .A2(n656), .ZN(n595) );
  NAND2_X1 U669 ( .A1(G66), .A2(n659), .ZN(n594) );
  NAND2_X1 U670 ( .A1(n595), .A2(n594), .ZN(n596) );
  NOR2_X1 U671 ( .A1(n597), .A2(n596), .ZN(n599) );
  XNOR2_X1 U672 ( .A(n599), .B(n598), .ZN(n600) );
  XNOR2_X2 U673 ( .A(KEYINPUT78), .B(n600), .ZN(n972) );
  NOR2_X1 U674 ( .A1(n972), .A2(G868), .ZN(n601) );
  NOR2_X1 U675 ( .A1(n602), .A2(n601), .ZN(n603) );
  XNOR2_X1 U676 ( .A(KEYINPUT79), .B(n603), .ZN(G284) );
  INV_X1 U677 ( .A(G301), .ZN(G171) );
  NAND2_X1 U678 ( .A1(G53), .A2(n654), .ZN(n605) );
  NAND2_X1 U679 ( .A1(G65), .A2(n659), .ZN(n604) );
  NAND2_X1 U680 ( .A1(n605), .A2(n604), .ZN(n609) );
  NAND2_X1 U681 ( .A1(G78), .A2(n655), .ZN(n607) );
  NAND2_X1 U682 ( .A1(G91), .A2(n656), .ZN(n606) );
  NAND2_X1 U683 ( .A1(n607), .A2(n606), .ZN(n608) );
  NOR2_X1 U684 ( .A1(n609), .A2(n608), .ZN(n978) );
  INV_X1 U685 ( .A(n978), .ZN(G299) );
  NOR2_X1 U686 ( .A1(G868), .A2(G299), .ZN(n610) );
  XNOR2_X1 U687 ( .A(n610), .B(KEYINPUT82), .ZN(n612) );
  INV_X1 U688 ( .A(G868), .ZN(n674) );
  NOR2_X1 U689 ( .A1(n674), .A2(G286), .ZN(n611) );
  NOR2_X1 U690 ( .A1(n612), .A2(n611), .ZN(G297) );
  NAND2_X1 U691 ( .A1(n613), .A2(G559), .ZN(n614) );
  NAND2_X1 U692 ( .A1(n614), .A2(n972), .ZN(n615) );
  XNOR2_X1 U693 ( .A(n615), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U694 ( .A1(n973), .A2(G868), .ZN(n618) );
  NAND2_X1 U695 ( .A1(n972), .A2(G868), .ZN(n616) );
  NOR2_X1 U696 ( .A1(G559), .A2(n616), .ZN(n617) );
  NOR2_X1 U697 ( .A1(n618), .A2(n617), .ZN(G282) );
  NAND2_X1 U698 ( .A1(n881), .A2(G111), .ZN(n619) );
  XOR2_X1 U699 ( .A(KEYINPUT83), .B(n619), .Z(n621) );
  NAND2_X1 U700 ( .A1(n877), .A2(G99), .ZN(n620) );
  NAND2_X1 U701 ( .A1(n621), .A2(n620), .ZN(n622) );
  XNOR2_X1 U702 ( .A(KEYINPUT84), .B(n622), .ZN(n625) );
  NAND2_X1 U703 ( .A1(n882), .A2(G123), .ZN(n623) );
  XOR2_X1 U704 ( .A(KEYINPUT18), .B(n623), .Z(n624) );
  NOR2_X1 U705 ( .A1(n625), .A2(n624), .ZN(n627) );
  NAND2_X1 U706 ( .A1(n878), .A2(G135), .ZN(n626) );
  NAND2_X1 U707 ( .A1(n627), .A2(n626), .ZN(n925) );
  XOR2_X1 U708 ( .A(n925), .B(G2096), .Z(n629) );
  XNOR2_X1 U709 ( .A(G2100), .B(KEYINPUT85), .ZN(n628) );
  NAND2_X1 U710 ( .A1(n629), .A2(n628), .ZN(G156) );
  NAND2_X1 U711 ( .A1(n972), .A2(G559), .ZN(n630) );
  XNOR2_X1 U712 ( .A(n630), .B(n973), .ZN(n671) );
  NOR2_X1 U713 ( .A1(n671), .A2(G860), .ZN(n640) );
  NAND2_X1 U714 ( .A1(G80), .A2(n655), .ZN(n632) );
  NAND2_X1 U715 ( .A1(G93), .A2(n656), .ZN(n631) );
  NAND2_X1 U716 ( .A1(n632), .A2(n631), .ZN(n633) );
  XNOR2_X1 U717 ( .A(n633), .B(KEYINPUT87), .ZN(n635) );
  NAND2_X1 U718 ( .A1(G55), .A2(n654), .ZN(n634) );
  NAND2_X1 U719 ( .A1(n635), .A2(n634), .ZN(n638) );
  NAND2_X1 U720 ( .A1(n659), .A2(G67), .ZN(n636) );
  XOR2_X1 U721 ( .A(KEYINPUT88), .B(n636), .Z(n637) );
  NOR2_X1 U722 ( .A1(n638), .A2(n637), .ZN(n673) );
  XNOR2_X1 U723 ( .A(n673), .B(KEYINPUT86), .ZN(n639) );
  XNOR2_X1 U724 ( .A(n640), .B(n639), .ZN(G145) );
  NAND2_X1 U725 ( .A1(G86), .A2(n656), .ZN(n642) );
  NAND2_X1 U726 ( .A1(G61), .A2(n659), .ZN(n641) );
  NAND2_X1 U727 ( .A1(n642), .A2(n641), .ZN(n645) );
  NAND2_X1 U728 ( .A1(n655), .A2(G73), .ZN(n643) );
  XOR2_X1 U729 ( .A(KEYINPUT2), .B(n643), .Z(n644) );
  NOR2_X1 U730 ( .A1(n645), .A2(n644), .ZN(n647) );
  NAND2_X1 U731 ( .A1(n654), .A2(G48), .ZN(n646) );
  NAND2_X1 U732 ( .A1(n647), .A2(n646), .ZN(G305) );
  NAND2_X1 U733 ( .A1(G49), .A2(n654), .ZN(n650) );
  NAND2_X1 U734 ( .A1(G87), .A2(n648), .ZN(n649) );
  NAND2_X1 U735 ( .A1(n650), .A2(n649), .ZN(n651) );
  NOR2_X1 U736 ( .A1(n659), .A2(n651), .ZN(n653) );
  NAND2_X1 U737 ( .A1(G651), .A2(G74), .ZN(n652) );
  NAND2_X1 U738 ( .A1(n653), .A2(n652), .ZN(G288) );
  NAND2_X1 U739 ( .A1(n654), .A2(G47), .ZN(n664) );
  NAND2_X1 U740 ( .A1(G72), .A2(n655), .ZN(n658) );
  NAND2_X1 U741 ( .A1(G85), .A2(n656), .ZN(n657) );
  NAND2_X1 U742 ( .A1(n658), .A2(n657), .ZN(n662) );
  NAND2_X1 U743 ( .A1(G60), .A2(n659), .ZN(n660) );
  XOR2_X1 U744 ( .A(KEYINPUT66), .B(n660), .Z(n661) );
  NOR2_X1 U745 ( .A1(n662), .A2(n661), .ZN(n663) );
  NAND2_X1 U746 ( .A1(n664), .A2(n663), .ZN(n665) );
  XOR2_X1 U747 ( .A(KEYINPUT67), .B(n665), .Z(G290) );
  XNOR2_X1 U748 ( .A(KEYINPUT19), .B(G305), .ZN(n666) );
  XNOR2_X1 U749 ( .A(n666), .B(G288), .ZN(n667) );
  XOR2_X1 U750 ( .A(n667), .B(n673), .Z(n669) );
  XNOR2_X1 U751 ( .A(G166), .B(n978), .ZN(n668) );
  XNOR2_X1 U752 ( .A(n669), .B(n668), .ZN(n670) );
  XNOR2_X1 U753 ( .A(n670), .B(G290), .ZN(n903) );
  XOR2_X1 U754 ( .A(n903), .B(n671), .Z(n672) );
  NOR2_X1 U755 ( .A1(n674), .A2(n672), .ZN(n676) );
  AND2_X1 U756 ( .A1(n674), .A2(n673), .ZN(n675) );
  NOR2_X1 U757 ( .A1(n676), .A2(n675), .ZN(G295) );
  NAND2_X1 U758 ( .A1(G2084), .A2(G2078), .ZN(n677) );
  XOR2_X1 U759 ( .A(KEYINPUT20), .B(n677), .Z(n678) );
  NAND2_X1 U760 ( .A1(G2090), .A2(n678), .ZN(n679) );
  XNOR2_X1 U761 ( .A(KEYINPUT21), .B(n679), .ZN(n680) );
  NAND2_X1 U762 ( .A1(n680), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U763 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NAND2_X1 U764 ( .A1(G120), .A2(G69), .ZN(n681) );
  NOR2_X1 U765 ( .A1(G237), .A2(n681), .ZN(n682) );
  XNOR2_X1 U766 ( .A(KEYINPUT90), .B(n682), .ZN(n683) );
  NAND2_X1 U767 ( .A1(n683), .A2(G108), .ZN(n837) );
  NAND2_X1 U768 ( .A1(G567), .A2(n837), .ZN(n688) );
  NOR2_X1 U769 ( .A1(G220), .A2(G219), .ZN(n684) );
  XOR2_X1 U770 ( .A(KEYINPUT22), .B(n684), .Z(n685) );
  NOR2_X1 U771 ( .A1(G218), .A2(n685), .ZN(n686) );
  NAND2_X1 U772 ( .A1(G96), .A2(n686), .ZN(n838) );
  NAND2_X1 U773 ( .A1(G2106), .A2(n838), .ZN(n687) );
  NAND2_X1 U774 ( .A1(n688), .A2(n687), .ZN(n857) );
  NAND2_X1 U775 ( .A1(G661), .A2(G483), .ZN(n689) );
  NOR2_X1 U776 ( .A1(n857), .A2(n689), .ZN(n836) );
  NAND2_X1 U777 ( .A1(n836), .A2(G36), .ZN(G176) );
  INV_X1 U778 ( .A(G166), .ZN(G303) );
  NAND2_X1 U779 ( .A1(G160), .A2(G40), .ZN(n797) );
  AND2_X1 U780 ( .A1(n722), .A2(G1341), .ZN(n691) );
  NOR2_X1 U781 ( .A1(n973), .A2(n691), .ZN(n694) );
  INV_X2 U782 ( .A(n722), .ZN(n716) );
  AND2_X1 U783 ( .A1(n716), .A2(G1996), .ZN(n692) );
  XOR2_X1 U784 ( .A(KEYINPUT26), .B(n692), .Z(n693) );
  AND2_X1 U785 ( .A1(n694), .A2(n693), .ZN(n700) );
  NAND2_X1 U786 ( .A1(n972), .A2(n700), .ZN(n699) );
  INV_X1 U787 ( .A(G1348), .ZN(n971) );
  NOR2_X1 U788 ( .A1(n716), .A2(n971), .ZN(n695) );
  XNOR2_X1 U789 ( .A(n695), .B(KEYINPUT99), .ZN(n697) );
  NAND2_X1 U790 ( .A1(n716), .A2(G2067), .ZN(n696) );
  NAND2_X1 U791 ( .A1(n697), .A2(n696), .ZN(n698) );
  NAND2_X1 U792 ( .A1(n699), .A2(n698), .ZN(n704) );
  INV_X1 U793 ( .A(n972), .ZN(n702) );
  INV_X1 U794 ( .A(n700), .ZN(n701) );
  NAND2_X1 U795 ( .A1(n702), .A2(n701), .ZN(n703) );
  NAND2_X1 U796 ( .A1(n704), .A2(n703), .ZN(n709) );
  NAND2_X1 U797 ( .A1(n716), .A2(G2072), .ZN(n705) );
  XNOR2_X1 U798 ( .A(n705), .B(KEYINPUT27), .ZN(n707) );
  INV_X1 U799 ( .A(G1956), .ZN(n1008) );
  NOR2_X1 U800 ( .A1(n1008), .A2(n716), .ZN(n706) );
  NOR2_X1 U801 ( .A1(n707), .A2(n706), .ZN(n710) );
  NAND2_X1 U802 ( .A1(n710), .A2(n978), .ZN(n708) );
  NAND2_X1 U803 ( .A1(n709), .A2(n708), .ZN(n714) );
  NOR2_X1 U804 ( .A1(n710), .A2(n978), .ZN(n712) );
  XOR2_X1 U805 ( .A(KEYINPUT28), .B(KEYINPUT98), .Z(n711) );
  XNOR2_X1 U806 ( .A(n712), .B(n711), .ZN(n713) );
  NAND2_X1 U807 ( .A1(n714), .A2(n713), .ZN(n715) );
  BUF_X1 U808 ( .A(n722), .Z(n732) );
  NAND2_X1 U809 ( .A1(G1961), .A2(n732), .ZN(n718) );
  XOR2_X1 U810 ( .A(G2078), .B(KEYINPUT25), .Z(n955) );
  NAND2_X1 U811 ( .A1(n716), .A2(n955), .ZN(n717) );
  NAND2_X1 U812 ( .A1(n718), .A2(n717), .ZN(n720) );
  NAND2_X1 U813 ( .A1(n719), .A2(n518), .ZN(n730) );
  NAND2_X1 U814 ( .A1(G301), .A2(n720), .ZN(n721) );
  XNOR2_X1 U815 ( .A(n721), .B(KEYINPUT101), .ZN(n727) );
  NAND2_X1 U816 ( .A1(n722), .A2(G8), .ZN(n731) );
  NOR2_X1 U817 ( .A1(n731), .A2(G1966), .ZN(n745) );
  NOR2_X1 U818 ( .A1(G2084), .A2(n722), .ZN(n744) );
  NOR2_X1 U819 ( .A1(n745), .A2(n744), .ZN(n723) );
  NAND2_X1 U820 ( .A1(n723), .A2(G8), .ZN(n724) );
  XNOR2_X1 U821 ( .A(n724), .B(KEYINPUT30), .ZN(n725) );
  NOR2_X1 U822 ( .A1(n725), .A2(G168), .ZN(n726) );
  NAND2_X1 U823 ( .A1(n730), .A2(n520), .ZN(n743) );
  NAND2_X1 U824 ( .A1(n743), .A2(G286), .ZN(n740) );
  INV_X1 U825 ( .A(G8), .ZN(n738) );
  NOR2_X1 U826 ( .A1(G1971), .A2(n731), .ZN(n734) );
  NOR2_X1 U827 ( .A1(G2090), .A2(n732), .ZN(n733) );
  NOR2_X1 U828 ( .A1(n734), .A2(n733), .ZN(n735) );
  NAND2_X1 U829 ( .A1(n735), .A2(G303), .ZN(n736) );
  XOR2_X1 U830 ( .A(KEYINPUT103), .B(n736), .Z(n737) );
  OR2_X1 U831 ( .A1(n738), .A2(n737), .ZN(n739) );
  XNOR2_X1 U832 ( .A(KEYINPUT104), .B(KEYINPUT32), .ZN(n741) );
  NOR2_X1 U833 ( .A1(n745), .A2(n519), .ZN(n746) );
  NAND2_X1 U834 ( .A1(n743), .A2(n746), .ZN(n767) );
  NAND2_X1 U835 ( .A1(G1976), .A2(G288), .ZN(n977) );
  INV_X1 U836 ( .A(KEYINPUT33), .ZN(n747) );
  NAND2_X1 U837 ( .A1(n977), .A2(n747), .ZN(n748) );
  NOR2_X1 U838 ( .A1(n748), .A2(n731), .ZN(n750) );
  AND2_X1 U839 ( .A1(n767), .A2(n750), .ZN(n749) );
  NAND2_X1 U840 ( .A1(n766), .A2(n749), .ZN(n759) );
  INV_X1 U841 ( .A(n750), .ZN(n752) );
  NOR2_X1 U842 ( .A1(G1976), .A2(G288), .ZN(n754) );
  NOR2_X1 U843 ( .A1(G1971), .A2(G303), .ZN(n751) );
  NOR2_X1 U844 ( .A1(n754), .A2(n751), .ZN(n979) );
  OR2_X1 U845 ( .A1(n752), .A2(n979), .ZN(n757) );
  INV_X1 U846 ( .A(n731), .ZN(n753) );
  NAND2_X1 U847 ( .A1(n754), .A2(n753), .ZN(n755) );
  NAND2_X1 U848 ( .A1(n755), .A2(KEYINPUT33), .ZN(n756) );
  AND2_X1 U849 ( .A1(n757), .A2(n756), .ZN(n758) );
  NAND2_X1 U850 ( .A1(n759), .A2(n758), .ZN(n760) );
  XNOR2_X1 U851 ( .A(n760), .B(KEYINPUT105), .ZN(n763) );
  XOR2_X1 U852 ( .A(G1981), .B(KEYINPUT106), .Z(n761) );
  XNOR2_X1 U853 ( .A(G305), .B(n761), .ZN(n987) );
  INV_X1 U854 ( .A(n987), .ZN(n762) );
  OR2_X1 U855 ( .A1(n763), .A2(n762), .ZN(n772) );
  NAND2_X1 U856 ( .A1(G8), .A2(G166), .ZN(n764) );
  NOR2_X1 U857 ( .A1(G2090), .A2(n764), .ZN(n765) );
  XNOR2_X1 U858 ( .A(n765), .B(KEYINPUT107), .ZN(n769) );
  NAND2_X1 U859 ( .A1(n767), .A2(n766), .ZN(n768) );
  NAND2_X1 U860 ( .A1(n769), .A2(n768), .ZN(n770) );
  NAND2_X1 U861 ( .A1(n770), .A2(n731), .ZN(n771) );
  NAND2_X1 U862 ( .A1(n772), .A2(n771), .ZN(n773) );
  XNOR2_X1 U863 ( .A(n773), .B(KEYINPUT108), .ZN(n777) );
  NOR2_X1 U864 ( .A1(G1981), .A2(G305), .ZN(n774) );
  XOR2_X1 U865 ( .A(n774), .B(KEYINPUT24), .Z(n775) );
  NOR2_X1 U866 ( .A1(n731), .A2(n775), .ZN(n776) );
  INV_X1 U867 ( .A(n778), .ZN(n813) );
  NAND2_X1 U868 ( .A1(n881), .A2(G107), .ZN(n781) );
  NAND2_X1 U869 ( .A1(G119), .A2(n882), .ZN(n779) );
  XOR2_X1 U870 ( .A(KEYINPUT97), .B(n779), .Z(n780) );
  NAND2_X1 U871 ( .A1(n781), .A2(n780), .ZN(n785) );
  NAND2_X1 U872 ( .A1(G95), .A2(n877), .ZN(n783) );
  NAND2_X1 U873 ( .A1(G131), .A2(n878), .ZN(n782) );
  NAND2_X1 U874 ( .A1(n783), .A2(n782), .ZN(n784) );
  NOR2_X1 U875 ( .A1(n785), .A2(n784), .ZN(n896) );
  INV_X1 U876 ( .A(G1991), .ZN(n951) );
  NOR2_X1 U877 ( .A1(n896), .A2(n951), .ZN(n794) );
  NAND2_X1 U878 ( .A1(G117), .A2(n881), .ZN(n787) );
  NAND2_X1 U879 ( .A1(G129), .A2(n882), .ZN(n786) );
  NAND2_X1 U880 ( .A1(n787), .A2(n786), .ZN(n790) );
  NAND2_X1 U881 ( .A1(n877), .A2(G105), .ZN(n788) );
  XOR2_X1 U882 ( .A(KEYINPUT38), .B(n788), .Z(n789) );
  NOR2_X1 U883 ( .A1(n790), .A2(n789), .ZN(n792) );
  NAND2_X1 U884 ( .A1(n878), .A2(G141), .ZN(n791) );
  NAND2_X1 U885 ( .A1(n792), .A2(n791), .ZN(n888) );
  AND2_X1 U886 ( .A1(n888), .A2(G1996), .ZN(n793) );
  NOR2_X1 U887 ( .A1(n794), .A2(n793), .ZN(n928) );
  INV_X1 U888 ( .A(n795), .ZN(n796) );
  NOR2_X1 U889 ( .A1(n797), .A2(n796), .ZN(n827) );
  INV_X1 U890 ( .A(n827), .ZN(n798) );
  NOR2_X1 U891 ( .A1(n928), .A2(n798), .ZN(n820) );
  XNOR2_X1 U892 ( .A(G2067), .B(KEYINPUT37), .ZN(n825) );
  XNOR2_X1 U893 ( .A(KEYINPUT34), .B(KEYINPUT94), .ZN(n802) );
  NAND2_X1 U894 ( .A1(G104), .A2(n877), .ZN(n800) );
  NAND2_X1 U895 ( .A1(G140), .A2(n878), .ZN(n799) );
  NAND2_X1 U896 ( .A1(n800), .A2(n799), .ZN(n801) );
  XNOR2_X1 U897 ( .A(n802), .B(n801), .ZN(n808) );
  XNOR2_X1 U898 ( .A(KEYINPUT95), .B(KEYINPUT35), .ZN(n806) );
  NAND2_X1 U899 ( .A1(G116), .A2(n881), .ZN(n804) );
  NAND2_X1 U900 ( .A1(G128), .A2(n882), .ZN(n803) );
  NAND2_X1 U901 ( .A1(n804), .A2(n803), .ZN(n805) );
  XNOR2_X1 U902 ( .A(n806), .B(n805), .ZN(n807) );
  NOR2_X1 U903 ( .A1(n808), .A2(n807), .ZN(n809) );
  XNOR2_X1 U904 ( .A(n809), .B(KEYINPUT36), .ZN(n897) );
  NOR2_X1 U905 ( .A1(n825), .A2(n897), .ZN(n810) );
  XNOR2_X1 U906 ( .A(n810), .B(KEYINPUT96), .ZN(n944) );
  NAND2_X1 U907 ( .A1(n827), .A2(n944), .ZN(n823) );
  INV_X1 U908 ( .A(n823), .ZN(n811) );
  XNOR2_X1 U909 ( .A(n814), .B(KEYINPUT109), .ZN(n816) );
  XNOR2_X1 U910 ( .A(G1986), .B(G290), .ZN(n984) );
  NAND2_X1 U911 ( .A1(n984), .A2(n827), .ZN(n815) );
  NAND2_X1 U912 ( .A1(n816), .A2(n815), .ZN(n830) );
  NOR2_X1 U913 ( .A1(G1996), .A2(n888), .ZN(n936) );
  AND2_X1 U914 ( .A1(n951), .A2(n896), .ZN(n924) );
  NOR2_X1 U915 ( .A1(G1986), .A2(G290), .ZN(n817) );
  XNOR2_X1 U916 ( .A(KEYINPUT110), .B(n817), .ZN(n818) );
  NOR2_X1 U917 ( .A1(n924), .A2(n818), .ZN(n819) );
  NOR2_X1 U918 ( .A1(n820), .A2(n819), .ZN(n821) );
  NOR2_X1 U919 ( .A1(n936), .A2(n821), .ZN(n822) );
  XNOR2_X1 U920 ( .A(KEYINPUT39), .B(n822), .ZN(n824) );
  NAND2_X1 U921 ( .A1(n824), .A2(n823), .ZN(n826) );
  NAND2_X1 U922 ( .A1(n897), .A2(n825), .ZN(n927) );
  NAND2_X1 U923 ( .A1(n826), .A2(n927), .ZN(n828) );
  NAND2_X1 U924 ( .A1(n828), .A2(n827), .ZN(n829) );
  NAND2_X1 U925 ( .A1(n830), .A2(n829), .ZN(n832) );
  XOR2_X1 U926 ( .A(KEYINPUT40), .B(KEYINPUT111), .Z(n831) );
  XNOR2_X1 U927 ( .A(n832), .B(n831), .ZN(G329) );
  NAND2_X1 U928 ( .A1(G2106), .A2(n833), .ZN(G217) );
  AND2_X1 U929 ( .A1(G15), .A2(G2), .ZN(n834) );
  NAND2_X1 U930 ( .A1(G661), .A2(n834), .ZN(G259) );
  NAND2_X1 U931 ( .A1(G3), .A2(G1), .ZN(n835) );
  NAND2_X1 U932 ( .A1(n836), .A2(n835), .ZN(G188) );
  XOR2_X1 U933 ( .A(G96), .B(KEYINPUT112), .Z(G221) );
  INV_X1 U935 ( .A(G120), .ZN(G236) );
  INV_X1 U936 ( .A(G108), .ZN(G238) );
  INV_X1 U937 ( .A(G69), .ZN(G235) );
  NOR2_X1 U938 ( .A1(n838), .A2(n837), .ZN(G325) );
  INV_X1 U939 ( .A(G325), .ZN(G261) );
  XOR2_X1 U940 ( .A(G2100), .B(G2096), .Z(n840) );
  XNOR2_X1 U941 ( .A(KEYINPUT42), .B(G2678), .ZN(n839) );
  XNOR2_X1 U942 ( .A(n840), .B(n839), .ZN(n844) );
  XOR2_X1 U943 ( .A(KEYINPUT43), .B(G2090), .Z(n842) );
  XNOR2_X1 U944 ( .A(G2067), .B(G2072), .ZN(n841) );
  XNOR2_X1 U945 ( .A(n842), .B(n841), .ZN(n843) );
  XOR2_X1 U946 ( .A(n844), .B(n843), .Z(n846) );
  XNOR2_X1 U947 ( .A(G2084), .B(G2078), .ZN(n845) );
  XNOR2_X1 U948 ( .A(n846), .B(n845), .ZN(G227) );
  XNOR2_X1 U949 ( .A(G1956), .B(G2474), .ZN(n856) );
  XOR2_X1 U950 ( .A(G1961), .B(G1971), .Z(n848) );
  XNOR2_X1 U951 ( .A(G1986), .B(G1976), .ZN(n847) );
  XNOR2_X1 U952 ( .A(n848), .B(n847), .ZN(n852) );
  XOR2_X1 U953 ( .A(G1966), .B(G1981), .Z(n850) );
  XNOR2_X1 U954 ( .A(G1996), .B(G1991), .ZN(n849) );
  XNOR2_X1 U955 ( .A(n850), .B(n849), .ZN(n851) );
  XOR2_X1 U956 ( .A(n852), .B(n851), .Z(n854) );
  XNOR2_X1 U957 ( .A(KEYINPUT114), .B(KEYINPUT41), .ZN(n853) );
  XNOR2_X1 U958 ( .A(n854), .B(n853), .ZN(n855) );
  XNOR2_X1 U959 ( .A(n856), .B(n855), .ZN(G229) );
  XNOR2_X1 U960 ( .A(KEYINPUT113), .B(n857), .ZN(G319) );
  NAND2_X1 U961 ( .A1(G124), .A2(n882), .ZN(n858) );
  XOR2_X1 U962 ( .A(KEYINPUT44), .B(n858), .Z(n859) );
  XNOR2_X1 U963 ( .A(n859), .B(KEYINPUT115), .ZN(n861) );
  NAND2_X1 U964 ( .A1(G112), .A2(n881), .ZN(n860) );
  NAND2_X1 U965 ( .A1(n861), .A2(n860), .ZN(n865) );
  NAND2_X1 U966 ( .A1(G100), .A2(n877), .ZN(n863) );
  NAND2_X1 U967 ( .A1(G136), .A2(n878), .ZN(n862) );
  NAND2_X1 U968 ( .A1(n863), .A2(n862), .ZN(n864) );
  NOR2_X1 U969 ( .A1(n865), .A2(n864), .ZN(G162) );
  XOR2_X1 U970 ( .A(KEYINPUT118), .B(KEYINPUT46), .Z(n867) );
  XNOR2_X1 U971 ( .A(G164), .B(KEYINPUT48), .ZN(n866) );
  XNOR2_X1 U972 ( .A(n867), .B(n866), .ZN(n895) );
  NAND2_X1 U973 ( .A1(n877), .A2(G106), .ZN(n868) );
  XOR2_X1 U974 ( .A(KEYINPUT117), .B(n868), .Z(n870) );
  NAND2_X1 U975 ( .A1(n878), .A2(G142), .ZN(n869) );
  NAND2_X1 U976 ( .A1(n870), .A2(n869), .ZN(n871) );
  XNOR2_X1 U977 ( .A(n871), .B(KEYINPUT45), .ZN(n873) );
  NAND2_X1 U978 ( .A1(G130), .A2(n882), .ZN(n872) );
  NAND2_X1 U979 ( .A1(n873), .A2(n872), .ZN(n876) );
  NAND2_X1 U980 ( .A1(n881), .A2(G118), .ZN(n874) );
  XOR2_X1 U981 ( .A(KEYINPUT116), .B(n874), .Z(n875) );
  NOR2_X1 U982 ( .A1(n876), .A2(n875), .ZN(n892) );
  NAND2_X1 U983 ( .A1(G103), .A2(n877), .ZN(n880) );
  NAND2_X1 U984 ( .A1(G139), .A2(n878), .ZN(n879) );
  NAND2_X1 U985 ( .A1(n880), .A2(n879), .ZN(n887) );
  NAND2_X1 U986 ( .A1(G115), .A2(n881), .ZN(n884) );
  NAND2_X1 U987 ( .A1(G127), .A2(n882), .ZN(n883) );
  NAND2_X1 U988 ( .A1(n884), .A2(n883), .ZN(n885) );
  XOR2_X1 U989 ( .A(KEYINPUT47), .B(n885), .Z(n886) );
  NOR2_X1 U990 ( .A1(n887), .A2(n886), .ZN(n931) );
  XOR2_X1 U991 ( .A(G162), .B(n931), .Z(n890) );
  XOR2_X1 U992 ( .A(G160), .B(n888), .Z(n889) );
  XNOR2_X1 U993 ( .A(n890), .B(n889), .ZN(n891) );
  XOR2_X1 U994 ( .A(n892), .B(n891), .Z(n893) );
  XNOR2_X1 U995 ( .A(n925), .B(n893), .ZN(n894) );
  XNOR2_X1 U996 ( .A(n895), .B(n894), .ZN(n899) );
  XNOR2_X1 U997 ( .A(n897), .B(n896), .ZN(n898) );
  XNOR2_X1 U998 ( .A(n899), .B(n898), .ZN(n900) );
  NOR2_X1 U999 ( .A1(G37), .A2(n900), .ZN(G395) );
  XOR2_X1 U1000 ( .A(KEYINPUT119), .B(n973), .Z(n902) );
  XNOR2_X1 U1001 ( .A(G286), .B(G171), .ZN(n901) );
  XNOR2_X1 U1002 ( .A(n902), .B(n901), .ZN(n905) );
  XNOR2_X1 U1003 ( .A(n972), .B(n903), .ZN(n904) );
  XNOR2_X1 U1004 ( .A(n905), .B(n904), .ZN(n906) );
  NOR2_X1 U1005 ( .A1(G37), .A2(n906), .ZN(G397) );
  XNOR2_X1 U1006 ( .A(KEYINPUT49), .B(KEYINPUT120), .ZN(n908) );
  NOR2_X1 U1007 ( .A1(G227), .A2(G229), .ZN(n907) );
  XNOR2_X1 U1008 ( .A(n908), .B(n907), .ZN(n919) );
  XOR2_X1 U1009 ( .A(G2451), .B(G2430), .Z(n910) );
  XNOR2_X1 U1010 ( .A(G2438), .B(G2443), .ZN(n909) );
  XNOR2_X1 U1011 ( .A(n910), .B(n909), .ZN(n916) );
  XOR2_X1 U1012 ( .A(G2435), .B(G2454), .Z(n912) );
  XNOR2_X1 U1013 ( .A(G1341), .B(G1348), .ZN(n911) );
  XNOR2_X1 U1014 ( .A(n912), .B(n911), .ZN(n914) );
  XOR2_X1 U1015 ( .A(G2446), .B(G2427), .Z(n913) );
  XNOR2_X1 U1016 ( .A(n914), .B(n913), .ZN(n915) );
  XOR2_X1 U1017 ( .A(n916), .B(n915), .Z(n917) );
  NAND2_X1 U1018 ( .A1(G14), .A2(n917), .ZN(n922) );
  NAND2_X1 U1019 ( .A1(G319), .A2(n922), .ZN(n918) );
  NOR2_X1 U1020 ( .A1(n919), .A2(n918), .ZN(n921) );
  NOR2_X1 U1021 ( .A1(G395), .A2(G397), .ZN(n920) );
  NAND2_X1 U1022 ( .A1(n921), .A2(n920), .ZN(G225) );
  INV_X1 U1023 ( .A(G225), .ZN(G308) );
  INV_X1 U1024 ( .A(n922), .ZN(G401) );
  XOR2_X1 U1025 ( .A(G160), .B(G2084), .Z(n923) );
  NOR2_X1 U1026 ( .A1(n924), .A2(n923), .ZN(n926) );
  NAND2_X1 U1027 ( .A1(n926), .A2(n925), .ZN(n930) );
  NAND2_X1 U1028 ( .A1(n928), .A2(n927), .ZN(n929) );
  NOR2_X1 U1029 ( .A1(n930), .A2(n929), .ZN(n942) );
  XOR2_X1 U1030 ( .A(G2072), .B(n931), .Z(n933) );
  XOR2_X1 U1031 ( .A(G164), .B(G2078), .Z(n932) );
  NOR2_X1 U1032 ( .A1(n933), .A2(n932), .ZN(n934) );
  XOR2_X1 U1033 ( .A(KEYINPUT50), .B(n934), .Z(n940) );
  XOR2_X1 U1034 ( .A(G2090), .B(G162), .Z(n935) );
  NOR2_X1 U1035 ( .A1(n936), .A2(n935), .ZN(n937) );
  XOR2_X1 U1036 ( .A(KEYINPUT121), .B(n937), .Z(n938) );
  XNOR2_X1 U1037 ( .A(KEYINPUT51), .B(n938), .ZN(n939) );
  NOR2_X1 U1038 ( .A1(n940), .A2(n939), .ZN(n941) );
  NAND2_X1 U1039 ( .A1(n942), .A2(n941), .ZN(n943) );
  NOR2_X1 U1040 ( .A1(n944), .A2(n943), .ZN(n945) );
  XNOR2_X1 U1041 ( .A(KEYINPUT52), .B(n945), .ZN(n946) );
  INV_X1 U1042 ( .A(KEYINPUT55), .ZN(n967) );
  NAND2_X1 U1043 ( .A1(n946), .A2(n967), .ZN(n947) );
  NAND2_X1 U1044 ( .A1(n947), .A2(G29), .ZN(n1028) );
  XNOR2_X1 U1045 ( .A(G2084), .B(G34), .ZN(n948) );
  XNOR2_X1 U1046 ( .A(n948), .B(KEYINPUT54), .ZN(n950) );
  XNOR2_X1 U1047 ( .A(G35), .B(G2090), .ZN(n949) );
  NOR2_X1 U1048 ( .A1(n950), .A2(n949), .ZN(n965) );
  XNOR2_X1 U1049 ( .A(G25), .B(n951), .ZN(n952) );
  NAND2_X1 U1050 ( .A1(n952), .A2(G28), .ZN(n961) );
  XNOR2_X1 U1051 ( .A(G2067), .B(G26), .ZN(n954) );
  XNOR2_X1 U1052 ( .A(G33), .B(G2072), .ZN(n953) );
  NOR2_X1 U1053 ( .A1(n954), .A2(n953), .ZN(n959) );
  XNOR2_X1 U1054 ( .A(G1996), .B(G32), .ZN(n957) );
  XNOR2_X1 U1055 ( .A(G27), .B(n955), .ZN(n956) );
  NOR2_X1 U1056 ( .A1(n957), .A2(n956), .ZN(n958) );
  NAND2_X1 U1057 ( .A1(n959), .A2(n958), .ZN(n960) );
  NOR2_X1 U1058 ( .A1(n961), .A2(n960), .ZN(n962) );
  XOR2_X1 U1059 ( .A(n962), .B(KEYINPUT122), .Z(n963) );
  XNOR2_X1 U1060 ( .A(KEYINPUT53), .B(n963), .ZN(n964) );
  NAND2_X1 U1061 ( .A1(n965), .A2(n964), .ZN(n966) );
  XNOR2_X1 U1062 ( .A(n967), .B(n966), .ZN(n969) );
  INV_X1 U1063 ( .A(G29), .ZN(n968) );
  NAND2_X1 U1064 ( .A1(n969), .A2(n968), .ZN(n970) );
  NAND2_X1 U1065 ( .A1(G11), .A2(n970), .ZN(n1026) );
  XNOR2_X1 U1066 ( .A(G16), .B(KEYINPUT56), .ZN(n996) );
  XNOR2_X1 U1067 ( .A(n972), .B(n971), .ZN(n975) );
  XNOR2_X1 U1068 ( .A(G1341), .B(n973), .ZN(n974) );
  NOR2_X1 U1069 ( .A1(n975), .A2(n974), .ZN(n994) );
  NAND2_X1 U1070 ( .A1(G1971), .A2(G303), .ZN(n976) );
  NAND2_X1 U1071 ( .A1(n977), .A2(n976), .ZN(n982) );
  XNOR2_X1 U1072 ( .A(n978), .B(G1956), .ZN(n980) );
  NAND2_X1 U1073 ( .A1(n980), .A2(n979), .ZN(n981) );
  NOR2_X1 U1074 ( .A1(n982), .A2(n981), .ZN(n986) );
  XNOR2_X1 U1075 ( .A(G1961), .B(G301), .ZN(n983) );
  NOR2_X1 U1076 ( .A1(n984), .A2(n983), .ZN(n985) );
  NAND2_X1 U1077 ( .A1(n986), .A2(n985), .ZN(n992) );
  XNOR2_X1 U1078 ( .A(G168), .B(G1966), .ZN(n988) );
  NAND2_X1 U1079 ( .A1(n988), .A2(n987), .ZN(n989) );
  XNOR2_X1 U1080 ( .A(n989), .B(KEYINPUT57), .ZN(n990) );
  XNOR2_X1 U1081 ( .A(n990), .B(KEYINPUT123), .ZN(n991) );
  NOR2_X1 U1082 ( .A1(n992), .A2(n991), .ZN(n993) );
  NAND2_X1 U1083 ( .A1(n994), .A2(n993), .ZN(n995) );
  NAND2_X1 U1084 ( .A1(n996), .A2(n995), .ZN(n1024) );
  INV_X1 U1085 ( .A(G16), .ZN(n1022) );
  XOR2_X1 U1086 ( .A(G1971), .B(KEYINPUT126), .Z(n997) );
  XNOR2_X1 U1087 ( .A(G22), .B(n997), .ZN(n1001) );
  XNOR2_X1 U1088 ( .A(G1986), .B(G24), .ZN(n999) );
  XNOR2_X1 U1089 ( .A(G23), .B(G1976), .ZN(n998) );
  NOR2_X1 U1090 ( .A1(n999), .A2(n998), .ZN(n1000) );
  NAND2_X1 U1091 ( .A1(n1001), .A2(n1000), .ZN(n1002) );
  XNOR2_X1 U1092 ( .A(n1002), .B(KEYINPUT58), .ZN(n1005) );
  XOR2_X1 U1093 ( .A(G1966), .B(KEYINPUT125), .Z(n1003) );
  XNOR2_X1 U1094 ( .A(G21), .B(n1003), .ZN(n1004) );
  NOR2_X1 U1095 ( .A1(n1005), .A2(n1004), .ZN(n1017) );
  XOR2_X1 U1096 ( .A(KEYINPUT124), .B(G4), .Z(n1007) );
  XNOR2_X1 U1097 ( .A(G1348), .B(KEYINPUT59), .ZN(n1006) );
  XNOR2_X1 U1098 ( .A(n1007), .B(n1006), .ZN(n1014) );
  XNOR2_X1 U1099 ( .A(G20), .B(n1008), .ZN(n1012) );
  XNOR2_X1 U1100 ( .A(G1981), .B(G6), .ZN(n1010) );
  XNOR2_X1 U1101 ( .A(G1341), .B(G19), .ZN(n1009) );
  NOR2_X1 U1102 ( .A1(n1010), .A2(n1009), .ZN(n1011) );
  NAND2_X1 U1103 ( .A1(n1012), .A2(n1011), .ZN(n1013) );
  NOR2_X1 U1104 ( .A1(n1014), .A2(n1013), .ZN(n1015) );
  XNOR2_X1 U1105 ( .A(n1015), .B(KEYINPUT60), .ZN(n1016) );
  NAND2_X1 U1106 ( .A1(n1017), .A2(n1016), .ZN(n1019) );
  XNOR2_X1 U1107 ( .A(G5), .B(G1961), .ZN(n1018) );
  NOR2_X1 U1108 ( .A1(n1019), .A2(n1018), .ZN(n1020) );
  XNOR2_X1 U1109 ( .A(KEYINPUT61), .B(n1020), .ZN(n1021) );
  NAND2_X1 U1110 ( .A1(n1022), .A2(n1021), .ZN(n1023) );
  NAND2_X1 U1111 ( .A1(n1024), .A2(n1023), .ZN(n1025) );
  NOR2_X1 U1112 ( .A1(n1026), .A2(n1025), .ZN(n1027) );
  NAND2_X1 U1113 ( .A1(n1028), .A2(n1027), .ZN(n1029) );
  XOR2_X1 U1114 ( .A(KEYINPUT62), .B(n1029), .Z(G311) );
  INV_X1 U1115 ( .A(G311), .ZN(G150) );
endmodule

