

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300,
         n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311,
         n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322,
         n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333,
         n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344,
         n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583;

  XOR2_X1 U322 ( .A(n384), .B(n383), .Z(n290) );
  XOR2_X1 U323 ( .A(n380), .B(G204GAT), .Z(n291) );
  XOR2_X1 U324 ( .A(n378), .B(KEYINPUT89), .Z(n292) );
  NOR2_X1 U325 ( .A1(n467), .A2(n453), .ZN(n454) );
  XNOR2_X1 U326 ( .A(n298), .B(n297), .ZN(n299) );
  XNOR2_X1 U327 ( .A(KEYINPUT48), .B(KEYINPUT110), .ZN(n372) );
  XNOR2_X1 U328 ( .A(n300), .B(n299), .ZN(n305) );
  XNOR2_X1 U329 ( .A(n373), .B(n372), .ZN(n525) );
  XOR2_X1 U330 ( .A(n307), .B(n306), .Z(n573) );
  XOR2_X1 U331 ( .A(n444), .B(n443), .Z(n529) );
  XNOR2_X1 U332 ( .A(KEYINPUT38), .B(n488), .ZN(n497) );
  XNOR2_X1 U333 ( .A(G190GAT), .B(KEYINPUT58), .ZN(n448) );
  XNOR2_X1 U334 ( .A(n449), .B(n448), .ZN(G1351GAT) );
  XOR2_X1 U335 ( .A(G99GAT), .B(G85GAT), .Z(n326) );
  XOR2_X1 U336 ( .A(G71GAT), .B(KEYINPUT13), .Z(n345) );
  XNOR2_X1 U337 ( .A(n326), .B(n345), .ZN(n307) );
  XOR2_X1 U338 ( .A(G64GAT), .B(KEYINPUT74), .Z(n294) );
  XNOR2_X1 U339 ( .A(G176GAT), .B(G92GAT), .ZN(n293) );
  XNOR2_X1 U340 ( .A(n294), .B(n293), .ZN(n378) );
  XNOR2_X1 U341 ( .A(KEYINPUT33), .B(n378), .ZN(n300) );
  XOR2_X1 U342 ( .A(KEYINPUT31), .B(KEYINPUT32), .Z(n296) );
  XNOR2_X1 U343 ( .A(KEYINPUT71), .B(KEYINPUT73), .ZN(n295) );
  XNOR2_X1 U344 ( .A(n296), .B(n295), .ZN(n298) );
  AND2_X1 U345 ( .A1(G230GAT), .A2(G233GAT), .ZN(n297) );
  XNOR2_X1 U346 ( .A(G120GAT), .B(G57GAT), .ZN(n301) );
  XNOR2_X1 U347 ( .A(n301), .B(G148GAT), .ZN(n396) );
  XOR2_X1 U348 ( .A(G78GAT), .B(G204GAT), .Z(n303) );
  XNOR2_X1 U349 ( .A(G106GAT), .B(KEYINPUT72), .ZN(n302) );
  XNOR2_X1 U350 ( .A(n303), .B(n302), .ZN(n420) );
  XOR2_X1 U351 ( .A(n396), .B(n420), .Z(n304) );
  XNOR2_X1 U352 ( .A(n305), .B(n304), .ZN(n306) );
  XOR2_X1 U353 ( .A(KEYINPUT41), .B(n573), .Z(n500) );
  XOR2_X1 U354 ( .A(G197GAT), .B(G36GAT), .Z(n309) );
  XNOR2_X1 U355 ( .A(G50GAT), .B(G29GAT), .ZN(n308) );
  XNOR2_X1 U356 ( .A(n309), .B(n308), .ZN(n313) );
  XOR2_X1 U357 ( .A(KEYINPUT29), .B(KEYINPUT70), .Z(n311) );
  XNOR2_X1 U358 ( .A(G169GAT), .B(G141GAT), .ZN(n310) );
  XNOR2_X1 U359 ( .A(n311), .B(n310), .ZN(n312) );
  XNOR2_X1 U360 ( .A(n313), .B(n312), .ZN(n323) );
  XOR2_X1 U361 ( .A(G113GAT), .B(G1GAT), .Z(n399) );
  XOR2_X1 U362 ( .A(G8GAT), .B(G15GAT), .Z(n315) );
  XNOR2_X1 U363 ( .A(KEYINPUT69), .B(G22GAT), .ZN(n314) );
  XNOR2_X1 U364 ( .A(n315), .B(n314), .ZN(n346) );
  XOR2_X1 U365 ( .A(n399), .B(n346), .Z(n317) );
  NAND2_X1 U366 ( .A1(G229GAT), .A2(G233GAT), .ZN(n316) );
  XNOR2_X1 U367 ( .A(n317), .B(n316), .ZN(n318) );
  XOR2_X1 U368 ( .A(n318), .B(KEYINPUT30), .Z(n321) );
  XNOR2_X1 U369 ( .A(G43GAT), .B(KEYINPUT8), .ZN(n319) );
  XNOR2_X1 U370 ( .A(n319), .B(KEYINPUT7), .ZN(n329) );
  XNOR2_X1 U371 ( .A(n329), .B(KEYINPUT68), .ZN(n320) );
  XNOR2_X1 U372 ( .A(n321), .B(n320), .ZN(n322) );
  XOR2_X1 U373 ( .A(n323), .B(n322), .Z(n501) );
  INV_X1 U374 ( .A(n501), .ZN(n570) );
  NAND2_X1 U375 ( .A1(n500), .A2(n570), .ZN(n324) );
  XNOR2_X1 U376 ( .A(n324), .B(KEYINPUT108), .ZN(n325) );
  XNOR2_X1 U377 ( .A(KEYINPUT46), .B(n325), .ZN(n361) );
  XOR2_X1 U378 ( .A(G36GAT), .B(G190GAT), .Z(n381) );
  XOR2_X1 U379 ( .A(n381), .B(n326), .Z(n328) );
  XOR2_X1 U380 ( .A(G29GAT), .B(G134GAT), .Z(n398) );
  XOR2_X1 U381 ( .A(G50GAT), .B(KEYINPUT75), .Z(n419) );
  XNOR2_X1 U382 ( .A(n398), .B(n419), .ZN(n327) );
  XNOR2_X1 U383 ( .A(n328), .B(n327), .ZN(n333) );
  XOR2_X1 U384 ( .A(n329), .B(KEYINPUT67), .Z(n331) );
  NAND2_X1 U385 ( .A1(G232GAT), .A2(G233GAT), .ZN(n330) );
  XNOR2_X1 U386 ( .A(n331), .B(n330), .ZN(n332) );
  XOR2_X1 U387 ( .A(n333), .B(n332), .Z(n341) );
  XOR2_X1 U388 ( .A(G106GAT), .B(KEYINPUT9), .Z(n335) );
  XNOR2_X1 U389 ( .A(G162GAT), .B(G218GAT), .ZN(n334) );
  XNOR2_X1 U390 ( .A(n335), .B(n334), .ZN(n339) );
  XOR2_X1 U391 ( .A(KEYINPUT10), .B(KEYINPUT11), .Z(n337) );
  XNOR2_X1 U392 ( .A(G92GAT), .B(KEYINPUT65), .ZN(n336) );
  XNOR2_X1 U393 ( .A(n337), .B(n336), .ZN(n338) );
  XNOR2_X1 U394 ( .A(n339), .B(n338), .ZN(n340) );
  XNOR2_X1 U395 ( .A(n341), .B(n340), .ZN(n363) );
  INV_X1 U396 ( .A(n363), .ZN(n342) );
  INV_X1 U397 ( .A(n342), .ZN(n551) );
  XOR2_X1 U398 ( .A(KEYINPUT12), .B(G57GAT), .Z(n344) );
  XNOR2_X1 U399 ( .A(G1GAT), .B(G183GAT), .ZN(n343) );
  XNOR2_X1 U400 ( .A(n344), .B(n343), .ZN(n359) );
  XOR2_X1 U401 ( .A(G64GAT), .B(G78GAT), .Z(n348) );
  XNOR2_X1 U402 ( .A(n346), .B(n345), .ZN(n347) );
  XNOR2_X1 U403 ( .A(n348), .B(n347), .ZN(n352) );
  XOR2_X1 U404 ( .A(G155GAT), .B(KEYINPUT14), .Z(n350) );
  NAND2_X1 U405 ( .A1(G231GAT), .A2(G233GAT), .ZN(n349) );
  XNOR2_X1 U406 ( .A(n350), .B(n349), .ZN(n351) );
  XOR2_X1 U407 ( .A(n352), .B(n351), .Z(n357) );
  XOR2_X1 U408 ( .A(KEYINPUT15), .B(KEYINPUT77), .Z(n354) );
  XNOR2_X1 U409 ( .A(G211GAT), .B(KEYINPUT76), .ZN(n353) );
  XNOR2_X1 U410 ( .A(n354), .B(n353), .ZN(n355) );
  XNOR2_X1 U411 ( .A(G127GAT), .B(n355), .ZN(n356) );
  XNOR2_X1 U412 ( .A(n357), .B(n356), .ZN(n358) );
  XOR2_X1 U413 ( .A(n359), .B(n358), .Z(n451) );
  INV_X1 U414 ( .A(n451), .ZN(n577) );
  NOR2_X1 U415 ( .A1(n551), .A2(n577), .ZN(n360) );
  AND2_X1 U416 ( .A1(n361), .A2(n360), .ZN(n362) );
  XNOR2_X1 U417 ( .A(n362), .B(KEYINPUT47), .ZN(n371) );
  INV_X1 U418 ( .A(n573), .ZN(n450) );
  XOR2_X1 U419 ( .A(KEYINPUT66), .B(KEYINPUT45), .Z(n366) );
  XOR2_X1 U420 ( .A(n363), .B(KEYINPUT99), .Z(n364) );
  XNOR2_X1 U421 ( .A(KEYINPUT36), .B(n364), .ZN(n580) );
  NAND2_X1 U422 ( .A1(n580), .A2(n577), .ZN(n365) );
  XNOR2_X1 U423 ( .A(n366), .B(n365), .ZN(n367) );
  NAND2_X1 U424 ( .A1(n450), .A2(n367), .ZN(n368) );
  NOR2_X1 U425 ( .A1(n570), .A2(n368), .ZN(n369) );
  XNOR2_X1 U426 ( .A(KEYINPUT109), .B(n369), .ZN(n370) );
  AND2_X1 U427 ( .A1(n371), .A2(n370), .ZN(n373) );
  XOR2_X1 U428 ( .A(KEYINPUT19), .B(KEYINPUT78), .Z(n375) );
  XNOR2_X1 U429 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n374) );
  XNOR2_X1 U430 ( .A(n375), .B(n374), .ZN(n377) );
  XOR2_X1 U431 ( .A(G169GAT), .B(G183GAT), .Z(n376) );
  XOR2_X1 U432 ( .A(n377), .B(n376), .Z(n443) );
  INV_X1 U433 ( .A(n443), .ZN(n384) );
  NAND2_X1 U434 ( .A1(G226GAT), .A2(G233GAT), .ZN(n379) );
  XNOR2_X1 U435 ( .A(n292), .B(n379), .ZN(n380) );
  XNOR2_X1 U436 ( .A(G8GAT), .B(n381), .ZN(n382) );
  XNOR2_X1 U437 ( .A(n291), .B(n382), .ZN(n383) );
  XOR2_X1 U438 ( .A(KEYINPUT82), .B(KEYINPUT81), .Z(n386) );
  XNOR2_X1 U439 ( .A(G211GAT), .B(KEYINPUT21), .ZN(n385) );
  XNOR2_X1 U440 ( .A(n386), .B(n385), .ZN(n388) );
  XOR2_X1 U441 ( .A(G197GAT), .B(G218GAT), .Z(n387) );
  XOR2_X1 U442 ( .A(n388), .B(n387), .Z(n424) );
  XOR2_X1 U443 ( .A(n290), .B(n424), .Z(n456) );
  NOR2_X1 U444 ( .A1(n525), .A2(n456), .ZN(n390) );
  INV_X1 U445 ( .A(KEYINPUT54), .ZN(n389) );
  XNOR2_X1 U446 ( .A(n390), .B(n389), .ZN(n411) );
  XOR2_X1 U447 ( .A(KEYINPUT87), .B(KEYINPUT4), .Z(n392) );
  XNOR2_X1 U448 ( .A(KEYINPUT85), .B(KEYINPUT84), .ZN(n391) );
  XNOR2_X1 U449 ( .A(n392), .B(n391), .ZN(n393) );
  XOR2_X1 U450 ( .A(n393), .B(KEYINPUT6), .Z(n395) );
  XOR2_X1 U451 ( .A(G127GAT), .B(KEYINPUT0), .Z(n431) );
  XNOR2_X1 U452 ( .A(n431), .B(G85GAT), .ZN(n394) );
  XNOR2_X1 U453 ( .A(n395), .B(n394), .ZN(n397) );
  XOR2_X1 U454 ( .A(n397), .B(n396), .Z(n401) );
  XNOR2_X1 U455 ( .A(n399), .B(n398), .ZN(n400) );
  XNOR2_X1 U456 ( .A(n401), .B(n400), .ZN(n405) );
  XOR2_X1 U457 ( .A(KEYINPUT86), .B(KEYINPUT1), .Z(n403) );
  NAND2_X1 U458 ( .A1(G225GAT), .A2(G233GAT), .ZN(n402) );
  XNOR2_X1 U459 ( .A(n403), .B(n402), .ZN(n404) );
  XOR2_X1 U460 ( .A(n405), .B(n404), .Z(n410) );
  XOR2_X1 U461 ( .A(G162GAT), .B(KEYINPUT2), .Z(n407) );
  XNOR2_X1 U462 ( .A(G141GAT), .B(KEYINPUT3), .ZN(n406) );
  XNOR2_X1 U463 ( .A(n407), .B(n406), .ZN(n408) );
  XNOR2_X1 U464 ( .A(G155GAT), .B(n408), .ZN(n427) );
  XOR2_X1 U465 ( .A(n427), .B(KEYINPUT5), .Z(n409) );
  XNOR2_X1 U466 ( .A(n410), .B(n409), .ZN(n462) );
  XNOR2_X1 U467 ( .A(KEYINPUT88), .B(n462), .ZN(n515) );
  NOR2_X1 U468 ( .A1(n411), .A2(n515), .ZN(n412) );
  XOR2_X1 U469 ( .A(KEYINPUT64), .B(n412), .Z(n568) );
  XOR2_X1 U470 ( .A(KEYINPUT79), .B(KEYINPUT22), .Z(n414) );
  XNOR2_X1 U471 ( .A(G22GAT), .B(G148GAT), .ZN(n413) );
  XNOR2_X1 U472 ( .A(n414), .B(n413), .ZN(n418) );
  XOR2_X1 U473 ( .A(KEYINPUT80), .B(KEYINPUT24), .Z(n416) );
  XNOR2_X1 U474 ( .A(KEYINPUT23), .B(KEYINPUT83), .ZN(n415) );
  XNOR2_X1 U475 ( .A(n416), .B(n415), .ZN(n417) );
  XOR2_X1 U476 ( .A(n418), .B(n417), .Z(n426) );
  XOR2_X1 U477 ( .A(n420), .B(n419), .Z(n422) );
  NAND2_X1 U478 ( .A1(G228GAT), .A2(G233GAT), .ZN(n421) );
  XNOR2_X1 U479 ( .A(n422), .B(n421), .ZN(n423) );
  XNOR2_X1 U480 ( .A(n424), .B(n423), .ZN(n425) );
  XNOR2_X1 U481 ( .A(n426), .B(n425), .ZN(n428) );
  XNOR2_X1 U482 ( .A(n428), .B(n427), .ZN(n467) );
  NOR2_X1 U483 ( .A1(n568), .A2(n467), .ZN(n430) );
  XNOR2_X1 U484 ( .A(KEYINPUT119), .B(KEYINPUT55), .ZN(n429) );
  XNOR2_X1 U485 ( .A(n430), .B(n429), .ZN(n445) );
  XOR2_X1 U486 ( .A(n431), .B(KEYINPUT20), .Z(n433) );
  NAND2_X1 U487 ( .A1(G227GAT), .A2(G233GAT), .ZN(n432) );
  XNOR2_X1 U488 ( .A(n433), .B(n432), .ZN(n437) );
  XOR2_X1 U489 ( .A(G120GAT), .B(G71GAT), .Z(n435) );
  XNOR2_X1 U490 ( .A(G113GAT), .B(G176GAT), .ZN(n434) );
  XNOR2_X1 U491 ( .A(n435), .B(n434), .ZN(n436) );
  XOR2_X1 U492 ( .A(n437), .B(n436), .Z(n442) );
  XOR2_X1 U493 ( .A(G190GAT), .B(G99GAT), .Z(n439) );
  XNOR2_X1 U494 ( .A(G43GAT), .B(G134GAT), .ZN(n438) );
  XNOR2_X1 U495 ( .A(n439), .B(n438), .ZN(n440) );
  XNOR2_X1 U496 ( .A(G15GAT), .B(n440), .ZN(n441) );
  XNOR2_X1 U497 ( .A(n442), .B(n441), .ZN(n444) );
  NAND2_X1 U498 ( .A1(n445), .A2(n529), .ZN(n447) );
  INV_X1 U499 ( .A(KEYINPUT120), .ZN(n446) );
  XNOR2_X1 U500 ( .A(n447), .B(n446), .ZN(n563) );
  NAND2_X1 U501 ( .A1(n563), .A2(n551), .ZN(n449) );
  NAND2_X1 U502 ( .A1(n570), .A2(n450), .ZN(n487) );
  NOR2_X1 U503 ( .A1(n551), .A2(n451), .ZN(n452) );
  XNOR2_X1 U504 ( .A(n452), .B(KEYINPUT16), .ZN(n472) );
  INV_X1 U505 ( .A(n529), .ZN(n468) );
  NOR2_X1 U506 ( .A1(n456), .A2(n468), .ZN(n453) );
  XNOR2_X1 U507 ( .A(n454), .B(KEYINPUT91), .ZN(n455) );
  XNOR2_X1 U508 ( .A(n455), .B(KEYINPUT25), .ZN(n460) );
  INV_X1 U509 ( .A(n456), .ZN(n517) );
  XOR2_X1 U510 ( .A(KEYINPUT27), .B(n517), .Z(n465) );
  NAND2_X1 U511 ( .A1(n468), .A2(n467), .ZN(n457) );
  XNOR2_X1 U512 ( .A(n457), .B(KEYINPUT90), .ZN(n458) );
  XNOR2_X1 U513 ( .A(KEYINPUT26), .B(n458), .ZN(n567) );
  NOR2_X1 U514 ( .A1(n465), .A2(n567), .ZN(n459) );
  NOR2_X1 U515 ( .A1(n460), .A2(n459), .ZN(n461) );
  XNOR2_X1 U516 ( .A(n461), .B(KEYINPUT92), .ZN(n463) );
  NOR2_X1 U517 ( .A1(n463), .A2(n462), .ZN(n464) );
  XNOR2_X1 U518 ( .A(n464), .B(KEYINPUT93), .ZN(n471) );
  INV_X1 U519 ( .A(n465), .ZN(n466) );
  NAND2_X1 U520 ( .A1(n515), .A2(n466), .ZN(n526) );
  XNOR2_X1 U521 ( .A(n467), .B(KEYINPUT28), .ZN(n528) );
  NOR2_X1 U522 ( .A1(n526), .A2(n528), .ZN(n469) );
  NAND2_X1 U523 ( .A1(n469), .A2(n468), .ZN(n470) );
  NAND2_X1 U524 ( .A1(n471), .A2(n470), .ZN(n484) );
  NAND2_X1 U525 ( .A1(n472), .A2(n484), .ZN(n503) );
  NOR2_X1 U526 ( .A1(n487), .A2(n503), .ZN(n473) );
  XNOR2_X1 U527 ( .A(KEYINPUT94), .B(n473), .ZN(n482) );
  NAND2_X1 U528 ( .A1(n482), .A2(n515), .ZN(n477) );
  XOR2_X1 U529 ( .A(KEYINPUT96), .B(KEYINPUT95), .Z(n475) );
  XNOR2_X1 U530 ( .A(G1GAT), .B(KEYINPUT34), .ZN(n474) );
  XNOR2_X1 U531 ( .A(n475), .B(n474), .ZN(n476) );
  XNOR2_X1 U532 ( .A(n477), .B(n476), .ZN(G1324GAT) );
  NAND2_X1 U533 ( .A1(n482), .A2(n517), .ZN(n478) );
  XNOR2_X1 U534 ( .A(n478), .B(G8GAT), .ZN(G1325GAT) );
  XOR2_X1 U535 ( .A(KEYINPUT97), .B(KEYINPUT35), .Z(n480) );
  NAND2_X1 U536 ( .A1(n529), .A2(n482), .ZN(n479) );
  XNOR2_X1 U537 ( .A(n480), .B(n479), .ZN(n481) );
  XOR2_X1 U538 ( .A(G15GAT), .B(n481), .Z(G1326GAT) );
  NAND2_X1 U539 ( .A1(n482), .A2(n528), .ZN(n483) );
  XNOR2_X1 U540 ( .A(n483), .B(G22GAT), .ZN(G1327GAT) );
  NAND2_X1 U541 ( .A1(n484), .A2(n580), .ZN(n485) );
  NOR2_X1 U542 ( .A1(n577), .A2(n485), .ZN(n486) );
  XNOR2_X1 U543 ( .A(KEYINPUT37), .B(n486), .ZN(n514) );
  NOR2_X1 U544 ( .A1(n514), .A2(n487), .ZN(n488) );
  NAND2_X1 U545 ( .A1(n497), .A2(n515), .ZN(n492) );
  XOR2_X1 U546 ( .A(KEYINPUT100), .B(KEYINPUT39), .Z(n490) );
  XNOR2_X1 U547 ( .A(G29GAT), .B(KEYINPUT98), .ZN(n489) );
  XNOR2_X1 U548 ( .A(n490), .B(n489), .ZN(n491) );
  XNOR2_X1 U549 ( .A(n492), .B(n491), .ZN(G1328GAT) );
  NAND2_X1 U550 ( .A1(n517), .A2(n497), .ZN(n493) );
  XNOR2_X1 U551 ( .A(G36GAT), .B(n493), .ZN(G1329GAT) );
  XOR2_X1 U552 ( .A(KEYINPUT40), .B(KEYINPUT101), .Z(n495) );
  NAND2_X1 U553 ( .A1(n529), .A2(n497), .ZN(n494) );
  XNOR2_X1 U554 ( .A(n495), .B(n494), .ZN(n496) );
  XNOR2_X1 U555 ( .A(n496), .B(G43GAT), .ZN(G1330GAT) );
  NAND2_X1 U556 ( .A1(n497), .A2(n528), .ZN(n498) );
  XNOR2_X1 U557 ( .A(n498), .B(KEYINPUT102), .ZN(n499) );
  XNOR2_X1 U558 ( .A(G50GAT), .B(n499), .ZN(G1331GAT) );
  XOR2_X1 U559 ( .A(KEYINPUT42), .B(KEYINPUT104), .Z(n505) );
  BUF_X1 U560 ( .A(n500), .Z(n560) );
  NAND2_X1 U561 ( .A1(n560), .A2(n501), .ZN(n502) );
  XOR2_X1 U562 ( .A(KEYINPUT103), .B(n502), .Z(n513) );
  NOR2_X1 U563 ( .A1(n503), .A2(n513), .ZN(n510) );
  NAND2_X1 U564 ( .A1(n510), .A2(n515), .ZN(n504) );
  XNOR2_X1 U565 ( .A(n505), .B(n504), .ZN(n506) );
  XOR2_X1 U566 ( .A(G57GAT), .B(n506), .Z(G1332GAT) );
  NAND2_X1 U567 ( .A1(n510), .A2(n517), .ZN(n507) );
  XNOR2_X1 U568 ( .A(n507), .B(G64GAT), .ZN(G1333GAT) );
  XOR2_X1 U569 ( .A(G71GAT), .B(KEYINPUT105), .Z(n509) );
  NAND2_X1 U570 ( .A1(n510), .A2(n529), .ZN(n508) );
  XNOR2_X1 U571 ( .A(n509), .B(n508), .ZN(G1334GAT) );
  XOR2_X1 U572 ( .A(G78GAT), .B(KEYINPUT43), .Z(n512) );
  NAND2_X1 U573 ( .A1(n510), .A2(n528), .ZN(n511) );
  XNOR2_X1 U574 ( .A(n512), .B(n511), .ZN(G1335GAT) );
  NOR2_X1 U575 ( .A1(n514), .A2(n513), .ZN(n521) );
  NAND2_X1 U576 ( .A1(n515), .A2(n521), .ZN(n516) );
  XNOR2_X1 U577 ( .A(n516), .B(G85GAT), .ZN(G1336GAT) );
  NAND2_X1 U578 ( .A1(n521), .A2(n517), .ZN(n518) );
  XNOR2_X1 U579 ( .A(n518), .B(KEYINPUT106), .ZN(n519) );
  XNOR2_X1 U580 ( .A(G92GAT), .B(n519), .ZN(G1337GAT) );
  NAND2_X1 U581 ( .A1(n521), .A2(n529), .ZN(n520) );
  XNOR2_X1 U582 ( .A(n520), .B(G99GAT), .ZN(G1338GAT) );
  XOR2_X1 U583 ( .A(KEYINPUT44), .B(KEYINPUT107), .Z(n523) );
  NAND2_X1 U584 ( .A1(n521), .A2(n528), .ZN(n522) );
  XNOR2_X1 U585 ( .A(n523), .B(n522), .ZN(n524) );
  XNOR2_X1 U586 ( .A(G106GAT), .B(n524), .ZN(G1339GAT) );
  XOR2_X1 U587 ( .A(G113GAT), .B(KEYINPUT113), .Z(n533) );
  NOR2_X1 U588 ( .A1(n526), .A2(n525), .ZN(n527) );
  XNOR2_X1 U589 ( .A(n527), .B(KEYINPUT111), .ZN(n543) );
  NOR2_X1 U590 ( .A1(n528), .A2(n543), .ZN(n530) );
  NAND2_X1 U591 ( .A1(n530), .A2(n529), .ZN(n531) );
  XOR2_X1 U592 ( .A(KEYINPUT112), .B(n531), .Z(n540) );
  NAND2_X1 U593 ( .A1(n570), .A2(n540), .ZN(n532) );
  XNOR2_X1 U594 ( .A(n533), .B(n532), .ZN(G1340GAT) );
  XOR2_X1 U595 ( .A(KEYINPUT114), .B(KEYINPUT49), .Z(n535) );
  NAND2_X1 U596 ( .A1(n540), .A2(n560), .ZN(n534) );
  XNOR2_X1 U597 ( .A(n535), .B(n534), .ZN(n536) );
  XNOR2_X1 U598 ( .A(G120GAT), .B(n536), .ZN(G1341GAT) );
  XOR2_X1 U599 ( .A(KEYINPUT115), .B(KEYINPUT50), .Z(n538) );
  NAND2_X1 U600 ( .A1(n540), .A2(n577), .ZN(n537) );
  XNOR2_X1 U601 ( .A(n538), .B(n537), .ZN(n539) );
  XNOR2_X1 U602 ( .A(G127GAT), .B(n539), .ZN(G1342GAT) );
  XOR2_X1 U603 ( .A(G134GAT), .B(KEYINPUT51), .Z(n542) );
  NAND2_X1 U604 ( .A1(n551), .A2(n540), .ZN(n541) );
  XNOR2_X1 U605 ( .A(n542), .B(n541), .ZN(G1343GAT) );
  NOR2_X1 U606 ( .A1(n567), .A2(n543), .ZN(n552) );
  NAND2_X1 U607 ( .A1(n570), .A2(n552), .ZN(n544) );
  XNOR2_X1 U608 ( .A(G141GAT), .B(n544), .ZN(G1344GAT) );
  XOR2_X1 U609 ( .A(KEYINPUT53), .B(KEYINPUT52), .Z(n546) );
  NAND2_X1 U610 ( .A1(n552), .A2(n560), .ZN(n545) );
  XNOR2_X1 U611 ( .A(n546), .B(n545), .ZN(n547) );
  XNOR2_X1 U612 ( .A(G148GAT), .B(n547), .ZN(G1345GAT) );
  XOR2_X1 U613 ( .A(KEYINPUT116), .B(KEYINPUT117), .Z(n549) );
  NAND2_X1 U614 ( .A1(n552), .A2(n577), .ZN(n548) );
  XNOR2_X1 U615 ( .A(n549), .B(n548), .ZN(n550) );
  XNOR2_X1 U616 ( .A(G155GAT), .B(n550), .ZN(G1346GAT) );
  NAND2_X1 U617 ( .A1(n552), .A2(n551), .ZN(n553) );
  XNOR2_X1 U618 ( .A(n553), .B(KEYINPUT118), .ZN(n554) );
  XNOR2_X1 U619 ( .A(G162GAT), .B(n554), .ZN(G1347GAT) );
  XOR2_X1 U620 ( .A(G169GAT), .B(KEYINPUT121), .Z(n556) );
  NAND2_X1 U621 ( .A1(n570), .A2(n563), .ZN(n555) );
  XNOR2_X1 U622 ( .A(n556), .B(n555), .ZN(G1348GAT) );
  XOR2_X1 U623 ( .A(KEYINPUT122), .B(KEYINPUT123), .Z(n558) );
  XNOR2_X1 U624 ( .A(G176GAT), .B(KEYINPUT57), .ZN(n557) );
  XNOR2_X1 U625 ( .A(n558), .B(n557), .ZN(n559) );
  XOR2_X1 U626 ( .A(KEYINPUT56), .B(n559), .Z(n562) );
  NAND2_X1 U627 ( .A1(n563), .A2(n560), .ZN(n561) );
  XNOR2_X1 U628 ( .A(n562), .B(n561), .ZN(G1349GAT) );
  NAND2_X1 U629 ( .A1(n563), .A2(n577), .ZN(n564) );
  XNOR2_X1 U630 ( .A(n564), .B(G183GAT), .ZN(G1350GAT) );
  XOR2_X1 U631 ( .A(KEYINPUT60), .B(KEYINPUT125), .Z(n566) );
  XNOR2_X1 U632 ( .A(G197GAT), .B(KEYINPUT59), .ZN(n565) );
  XNOR2_X1 U633 ( .A(n566), .B(n565), .ZN(n572) );
  NOR2_X1 U634 ( .A1(n568), .A2(n567), .ZN(n569) );
  XNOR2_X1 U635 ( .A(KEYINPUT124), .B(n569), .ZN(n581) );
  NAND2_X1 U636 ( .A1(n581), .A2(n570), .ZN(n571) );
  XOR2_X1 U637 ( .A(n572), .B(n571), .Z(G1352GAT) );
  XOR2_X1 U638 ( .A(KEYINPUT126), .B(KEYINPUT61), .Z(n575) );
  NAND2_X1 U639 ( .A1(n581), .A2(n573), .ZN(n574) );
  XNOR2_X1 U640 ( .A(n575), .B(n574), .ZN(n576) );
  XNOR2_X1 U641 ( .A(G204GAT), .B(n576), .ZN(G1353GAT) );
  XOR2_X1 U642 ( .A(G211GAT), .B(KEYINPUT127), .Z(n579) );
  NAND2_X1 U643 ( .A1(n581), .A2(n577), .ZN(n578) );
  XNOR2_X1 U644 ( .A(n579), .B(n578), .ZN(G1354GAT) );
  NAND2_X1 U645 ( .A1(n581), .A2(n580), .ZN(n582) );
  XNOR2_X1 U646 ( .A(n582), .B(KEYINPUT62), .ZN(n583) );
  XNOR2_X1 U647 ( .A(G218GAT), .B(n583), .ZN(G1355GAT) );
endmodule

