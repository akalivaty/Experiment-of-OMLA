//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 0 1 0 0 1 1 0 0 0 1 1 1 0 0 1 1 0 0 1 1 1 0 1 1 1 1 1 1 1 1 1 0 1 1 1 1 0 0 0 0 1 0 1 1 0 0 0 1 0 1 0 1 0 1 0 1 0 0 0 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:28:03 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n636, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n647, new_n648, new_n649, new_n650, new_n651, new_n652,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n683, new_n684, new_n685, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n697, new_n699,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n705, new_n707,
    new_n708, new_n709, new_n710, new_n711, new_n712, new_n713, new_n714,
    new_n715, new_n716, new_n717, new_n719, new_n720, new_n721, new_n722,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n741, new_n742, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n896, new_n897, new_n898,
    new_n899, new_n900, new_n901, new_n902, new_n904, new_n905, new_n906,
    new_n907, new_n908, new_n909, new_n910, new_n911, new_n912, new_n913,
    new_n914, new_n915, new_n916, new_n917, new_n918, new_n919, new_n920,
    new_n921, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n960, new_n961, new_n962, new_n963, new_n964, new_n965, new_n966,
    new_n967, new_n968;
  XNOR2_X1  g000(.A(KEYINPUT9), .B(G234), .ZN(new_n187));
  XNOR2_X1  g001(.A(new_n187), .B(KEYINPUT75), .ZN(new_n188));
  OAI21_X1  g002(.A(G221), .B1(new_n188), .B2(G902), .ZN(new_n189));
  XNOR2_X1  g003(.A(KEYINPUT69), .B(G902), .ZN(new_n190));
  XNOR2_X1  g004(.A(KEYINPUT79), .B(G469), .ZN(new_n191));
  INV_X1    g005(.A(KEYINPUT64), .ZN(new_n192));
  INV_X1    g006(.A(G143), .ZN(new_n193));
  OAI21_X1  g007(.A(new_n192), .B1(new_n193), .B2(G146), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n193), .A2(G146), .ZN(new_n195));
  INV_X1    g009(.A(G146), .ZN(new_n196));
  NAND3_X1  g010(.A1(new_n196), .A2(KEYINPUT64), .A3(G143), .ZN(new_n197));
  NAND3_X1  g011(.A1(new_n194), .A2(new_n195), .A3(new_n197), .ZN(new_n198));
  NOR2_X1   g012(.A1(new_n193), .A2(G146), .ZN(new_n199));
  INV_X1    g013(.A(KEYINPUT1), .ZN(new_n200));
  OAI21_X1  g014(.A(G128), .B1(new_n199), .B2(new_n200), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n198), .A2(new_n201), .ZN(new_n202));
  INV_X1    g016(.A(G128), .ZN(new_n203));
  NOR2_X1   g017(.A1(new_n203), .A2(KEYINPUT1), .ZN(new_n204));
  NAND4_X1  g018(.A1(new_n194), .A2(new_n197), .A3(new_n204), .A4(new_n195), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n202), .A2(new_n205), .ZN(new_n206));
  INV_X1    g020(.A(G104), .ZN(new_n207));
  OAI21_X1  g021(.A(KEYINPUT3), .B1(new_n207), .B2(G107), .ZN(new_n208));
  INV_X1    g022(.A(KEYINPUT3), .ZN(new_n209));
  INV_X1    g023(.A(G107), .ZN(new_n210));
  NAND3_X1  g024(.A1(new_n209), .A2(new_n210), .A3(G104), .ZN(new_n211));
  INV_X1    g025(.A(G101), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n207), .A2(G107), .ZN(new_n213));
  NAND4_X1  g027(.A1(new_n208), .A2(new_n211), .A3(new_n212), .A4(new_n213), .ZN(new_n214));
  NOR2_X1   g028(.A1(new_n210), .A2(G104), .ZN(new_n215));
  NOR2_X1   g029(.A1(new_n207), .A2(G107), .ZN(new_n216));
  OAI21_X1  g030(.A(G101), .B1(new_n215), .B2(new_n216), .ZN(new_n217));
  AND2_X1   g031(.A1(new_n214), .A2(new_n217), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n206), .A2(new_n218), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n196), .A2(G143), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n195), .A2(new_n220), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n201), .A2(new_n221), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n222), .A2(new_n205), .ZN(new_n223));
  OAI21_X1  g037(.A(new_n219), .B1(new_n223), .B2(new_n218), .ZN(new_n224));
  INV_X1    g038(.A(KEYINPUT11), .ZN(new_n225));
  INV_X1    g039(.A(G134), .ZN(new_n226));
  OAI21_X1  g040(.A(new_n225), .B1(new_n226), .B2(G137), .ZN(new_n227));
  INV_X1    g041(.A(G137), .ZN(new_n228));
  NAND3_X1  g042(.A1(new_n228), .A2(KEYINPUT11), .A3(G134), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n226), .A2(G137), .ZN(new_n230));
  NAND3_X1  g044(.A1(new_n227), .A2(new_n229), .A3(new_n230), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n231), .A2(G131), .ZN(new_n232));
  INV_X1    g046(.A(KEYINPUT66), .ZN(new_n233));
  INV_X1    g047(.A(G131), .ZN(new_n234));
  NAND4_X1  g048(.A1(new_n227), .A2(new_n229), .A3(new_n234), .A4(new_n230), .ZN(new_n235));
  NAND3_X1  g049(.A1(new_n232), .A2(new_n233), .A3(new_n235), .ZN(new_n236));
  NAND3_X1  g050(.A1(new_n231), .A2(KEYINPUT66), .A3(G131), .ZN(new_n237));
  AND2_X1   g051(.A1(new_n236), .A2(new_n237), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n224), .A2(new_n238), .ZN(new_n239));
  INV_X1    g053(.A(KEYINPUT12), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n239), .A2(new_n240), .ZN(new_n241));
  NAND3_X1  g055(.A1(new_n224), .A2(KEYINPUT12), .A3(new_n238), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n241), .A2(new_n242), .ZN(new_n243));
  XNOR2_X1  g057(.A(G110), .B(G140), .ZN(new_n244));
  INV_X1    g058(.A(G227), .ZN(new_n245));
  NOR2_X1   g059(.A1(new_n245), .A2(G953), .ZN(new_n246));
  XOR2_X1   g060(.A(new_n244), .B(new_n246), .Z(new_n247));
  NAND3_X1  g061(.A1(new_n208), .A2(new_n211), .A3(new_n213), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n248), .A2(G101), .ZN(new_n249));
  NOR2_X1   g063(.A1(new_n249), .A2(KEYINPUT4), .ZN(new_n250));
  AND2_X1   g064(.A1(new_n248), .A2(G101), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n214), .A2(KEYINPUT4), .ZN(new_n252));
  OAI21_X1  g066(.A(KEYINPUT76), .B1(new_n251), .B2(new_n252), .ZN(new_n253));
  INV_X1    g067(.A(KEYINPUT76), .ZN(new_n254));
  NAND4_X1  g068(.A1(new_n249), .A2(new_n254), .A3(KEYINPUT4), .A4(new_n214), .ZN(new_n255));
  AOI21_X1  g069(.A(new_n250), .B1(new_n253), .B2(new_n255), .ZN(new_n256));
  NAND2_X1  g070(.A1(KEYINPUT0), .A2(G128), .ZN(new_n257));
  OR2_X1    g071(.A1(KEYINPUT0), .A2(G128), .ZN(new_n258));
  NOR2_X1   g072(.A1(new_n196), .A2(G143), .ZN(new_n259));
  OAI211_X1 g073(.A(new_n257), .B(new_n258), .C1(new_n259), .C2(new_n199), .ZN(new_n260));
  INV_X1    g074(.A(new_n257), .ZN(new_n261));
  NAND4_X1  g075(.A1(new_n194), .A2(new_n197), .A3(new_n195), .A4(new_n261), .ZN(new_n262));
  AND2_X1   g076(.A1(new_n260), .A2(new_n262), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n256), .A2(new_n263), .ZN(new_n264));
  INV_X1    g078(.A(new_n238), .ZN(new_n265));
  XOR2_X1   g079(.A(KEYINPUT77), .B(KEYINPUT10), .Z(new_n266));
  INV_X1    g080(.A(KEYINPUT10), .ZN(new_n267));
  AOI21_X1  g081(.A(new_n267), .B1(new_n222), .B2(new_n205), .ZN(new_n268));
  AOI22_X1  g082(.A1(new_n219), .A2(new_n266), .B1(new_n218), .B2(new_n268), .ZN(new_n269));
  NAND3_X1  g083(.A1(new_n264), .A2(new_n265), .A3(new_n269), .ZN(new_n270));
  NAND3_X1  g084(.A1(new_n243), .A2(new_n247), .A3(new_n270), .ZN(new_n271));
  INV_X1    g085(.A(new_n271), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n264), .A2(new_n269), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n273), .A2(new_n238), .ZN(new_n274));
  AOI21_X1  g088(.A(new_n247), .B1(new_n274), .B2(new_n270), .ZN(new_n275));
  OAI211_X1 g089(.A(new_n190), .B(new_n191), .C1(new_n272), .C2(new_n275), .ZN(new_n276));
  INV_X1    g090(.A(G469), .ZN(new_n277));
  INV_X1    g091(.A(G902), .ZN(new_n278));
  NOR2_X1   g092(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  INV_X1    g093(.A(new_n279), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n276), .A2(new_n280), .ZN(new_n281));
  AOI21_X1  g095(.A(new_n247), .B1(new_n243), .B2(new_n270), .ZN(new_n282));
  AOI21_X1  g096(.A(new_n265), .B1(new_n264), .B2(new_n269), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n270), .A2(new_n247), .ZN(new_n284));
  INV_X1    g098(.A(KEYINPUT78), .ZN(new_n285));
  AOI21_X1  g099(.A(new_n283), .B1(new_n284), .B2(new_n285), .ZN(new_n286));
  NAND3_X1  g100(.A1(new_n270), .A2(KEYINPUT78), .A3(new_n247), .ZN(new_n287));
  AOI211_X1 g101(.A(new_n277), .B(new_n282), .C1(new_n286), .C2(new_n287), .ZN(new_n288));
  OAI21_X1  g102(.A(new_n189), .B1(new_n281), .B2(new_n288), .ZN(new_n289));
  XNOR2_X1  g103(.A(G113), .B(G122), .ZN(new_n290));
  XNOR2_X1  g104(.A(new_n290), .B(new_n207), .ZN(new_n291));
  NOR2_X1   g105(.A1(G237), .A2(G953), .ZN(new_n292));
  AOI21_X1  g106(.A(G143), .B1(new_n292), .B2(G214), .ZN(new_n293));
  INV_X1    g107(.A(G237), .ZN(new_n294));
  INV_X1    g108(.A(G953), .ZN(new_n295));
  NAND4_X1  g109(.A1(new_n294), .A2(new_n295), .A3(G143), .A4(G214), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n296), .A2(KEYINPUT84), .ZN(new_n297));
  INV_X1    g111(.A(KEYINPUT84), .ZN(new_n298));
  NAND4_X1  g112(.A1(new_n292), .A2(new_n298), .A3(G143), .A4(G214), .ZN(new_n299));
  AOI21_X1  g113(.A(new_n293), .B1(new_n297), .B2(new_n299), .ZN(new_n300));
  NOR2_X1   g114(.A1(new_n300), .A2(new_n234), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n301), .A2(KEYINPUT18), .ZN(new_n302));
  NAND2_X1  g116(.A1(KEYINPUT18), .A2(G131), .ZN(new_n303));
  XNOR2_X1  g117(.A(G125), .B(G140), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n304), .A2(new_n196), .ZN(new_n305));
  XOR2_X1   g119(.A(G125), .B(G140), .Z(new_n306));
  NAND2_X1  g120(.A1(new_n306), .A2(G146), .ZN(new_n307));
  AOI22_X1  g121(.A1(new_n300), .A2(new_n303), .B1(new_n305), .B2(new_n307), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n302), .A2(new_n308), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n301), .A2(KEYINPUT17), .ZN(new_n310));
  INV_X1    g124(.A(G125), .ZN(new_n311));
  NOR3_X1   g125(.A1(new_n311), .A2(KEYINPUT16), .A3(G140), .ZN(new_n312));
  AOI211_X1 g126(.A(new_n196), .B(new_n312), .C1(KEYINPUT16), .C2(new_n304), .ZN(new_n313));
  INV_X1    g127(.A(new_n313), .ZN(new_n314));
  AOI21_X1  g128(.A(new_n312), .B1(new_n304), .B2(KEYINPUT16), .ZN(new_n315));
  OAI21_X1  g129(.A(KEYINPUT72), .B1(new_n315), .B2(G146), .ZN(new_n316));
  INV_X1    g130(.A(KEYINPUT72), .ZN(new_n317));
  AND2_X1   g131(.A1(new_n304), .A2(KEYINPUT16), .ZN(new_n318));
  OAI211_X1 g132(.A(new_n317), .B(new_n196), .C1(new_n318), .C2(new_n312), .ZN(new_n319));
  NAND4_X1  g133(.A1(new_n310), .A2(new_n314), .A3(new_n316), .A4(new_n319), .ZN(new_n320));
  AND2_X1   g134(.A1(new_n300), .A2(new_n234), .ZN(new_n321));
  NOR3_X1   g135(.A1(new_n321), .A2(new_n301), .A3(KEYINPUT17), .ZN(new_n322));
  OAI211_X1 g136(.A(new_n291), .B(new_n309), .C1(new_n320), .C2(new_n322), .ZN(new_n323));
  INV_X1    g137(.A(KEYINPUT19), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n306), .A2(new_n324), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n304), .A2(KEYINPUT19), .ZN(new_n326));
  AOI21_X1  g140(.A(G146), .B1(new_n325), .B2(new_n326), .ZN(new_n327));
  NOR2_X1   g141(.A1(new_n327), .A2(new_n313), .ZN(new_n328));
  OAI21_X1  g142(.A(new_n328), .B1(new_n321), .B2(new_n301), .ZN(new_n329));
  NAND3_X1  g143(.A1(new_n329), .A2(new_n309), .A3(KEYINPUT85), .ZN(new_n330));
  INV_X1    g144(.A(new_n291), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n330), .A2(new_n331), .ZN(new_n332));
  AOI21_X1  g146(.A(KEYINPUT85), .B1(new_n329), .B2(new_n309), .ZN(new_n333));
  OAI21_X1  g147(.A(new_n323), .B1(new_n332), .B2(new_n333), .ZN(new_n334));
  NOR2_X1   g148(.A1(G475), .A2(G902), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n336), .A2(KEYINPUT20), .ZN(new_n337));
  INV_X1    g151(.A(KEYINPUT20), .ZN(new_n338));
  NAND3_X1  g152(.A1(new_n334), .A2(new_n338), .A3(new_n335), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n337), .A2(new_n339), .ZN(new_n340));
  INV_X1    g154(.A(G475), .ZN(new_n341));
  OAI21_X1  g155(.A(new_n309), .B1(new_n320), .B2(new_n322), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n342), .A2(new_n331), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n343), .A2(new_n323), .ZN(new_n344));
  AOI21_X1  g158(.A(new_n341), .B1(new_n344), .B2(new_n278), .ZN(new_n345));
  INV_X1    g159(.A(new_n345), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n340), .A2(new_n346), .ZN(new_n347));
  INV_X1    g161(.A(new_n347), .ZN(new_n348));
  INV_X1    g162(.A(G122), .ZN(new_n349));
  OAI21_X1  g163(.A(KEYINPUT86), .B1(new_n349), .B2(G116), .ZN(new_n350));
  INV_X1    g164(.A(KEYINPUT86), .ZN(new_n351));
  INV_X1    g165(.A(G116), .ZN(new_n352));
  NAND3_X1  g166(.A1(new_n351), .A2(new_n352), .A3(G122), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n350), .A2(new_n353), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n349), .A2(G116), .ZN(new_n355));
  NAND3_X1  g169(.A1(new_n354), .A2(new_n210), .A3(new_n355), .ZN(new_n356));
  INV_X1    g170(.A(KEYINPUT89), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n193), .A2(G128), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n203), .A2(G143), .ZN(new_n359));
  NAND3_X1  g173(.A1(new_n358), .A2(new_n359), .A3(new_n226), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n358), .A2(new_n359), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n361), .A2(G134), .ZN(new_n362));
  AOI22_X1  g176(.A1(new_n356), .A2(new_n357), .B1(new_n360), .B2(new_n362), .ZN(new_n363));
  NAND4_X1  g177(.A1(new_n354), .A2(KEYINPUT89), .A3(new_n210), .A4(new_n355), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n363), .A2(new_n364), .ZN(new_n365));
  OR2_X1    g179(.A1(new_n354), .A2(KEYINPUT14), .ZN(new_n366));
  AOI22_X1  g180(.A1(new_n354), .A2(KEYINPUT14), .B1(G116), .B2(new_n349), .ZN(new_n367));
  AOI21_X1  g181(.A(new_n210), .B1(new_n366), .B2(new_n367), .ZN(new_n368));
  OAI21_X1  g182(.A(KEYINPUT90), .B1(new_n365), .B2(new_n368), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n366), .A2(new_n367), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n370), .A2(G107), .ZN(new_n371));
  INV_X1    g185(.A(KEYINPUT90), .ZN(new_n372));
  NAND4_X1  g186(.A1(new_n371), .A2(new_n372), .A3(new_n363), .A4(new_n364), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n369), .A2(new_n373), .ZN(new_n374));
  INV_X1    g188(.A(G217), .ZN(new_n375));
  NOR3_X1   g189(.A1(new_n188), .A2(new_n375), .A3(G953), .ZN(new_n376));
  INV_X1    g190(.A(KEYINPUT87), .ZN(new_n377));
  INV_X1    g191(.A(KEYINPUT13), .ZN(new_n378));
  NAND3_X1  g192(.A1(new_n358), .A2(new_n377), .A3(new_n378), .ZN(new_n379));
  OAI211_X1 g193(.A(new_n379), .B(new_n359), .C1(new_n378), .C2(new_n358), .ZN(new_n380));
  AOI21_X1  g194(.A(new_n377), .B1(new_n358), .B2(new_n378), .ZN(new_n381));
  OAI21_X1  g195(.A(G134), .B1(new_n380), .B2(new_n381), .ZN(new_n382));
  INV_X1    g196(.A(KEYINPUT88), .ZN(new_n383));
  OR2_X1    g197(.A1(new_n382), .A2(new_n383), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n354), .A2(new_n355), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n385), .A2(G107), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n386), .A2(new_n356), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n382), .A2(new_n383), .ZN(new_n388));
  NAND4_X1  g202(.A1(new_n384), .A2(new_n387), .A3(new_n360), .A4(new_n388), .ZN(new_n389));
  AND3_X1   g203(.A1(new_n374), .A2(new_n376), .A3(new_n389), .ZN(new_n390));
  AOI21_X1  g204(.A(new_n376), .B1(new_n374), .B2(new_n389), .ZN(new_n391));
  OAI21_X1  g205(.A(new_n190), .B1(new_n390), .B2(new_n391), .ZN(new_n392));
  INV_X1    g206(.A(G478), .ZN(new_n393));
  INV_X1    g207(.A(KEYINPUT91), .ZN(new_n394));
  NOR2_X1   g208(.A1(new_n394), .A2(KEYINPUT15), .ZN(new_n395));
  INV_X1    g209(.A(new_n395), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n394), .A2(KEYINPUT15), .ZN(new_n397));
  AOI21_X1  g211(.A(new_n393), .B1(new_n396), .B2(new_n397), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n392), .A2(new_n398), .ZN(new_n399));
  INV_X1    g213(.A(new_n398), .ZN(new_n400));
  OAI211_X1 g214(.A(new_n190), .B(new_n400), .C1(new_n390), .C2(new_n391), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n399), .A2(new_n401), .ZN(new_n402));
  NAND2_X1  g216(.A1(G234), .A2(G237), .ZN(new_n403));
  NAND3_X1  g217(.A1(new_n403), .A2(G952), .A3(new_n295), .ZN(new_n404));
  XNOR2_X1  g218(.A(new_n404), .B(KEYINPUT92), .ZN(new_n405));
  INV_X1    g219(.A(new_n405), .ZN(new_n406));
  INV_X1    g220(.A(new_n190), .ZN(new_n407));
  AND3_X1   g221(.A1(new_n407), .A2(G953), .A3(new_n403), .ZN(new_n408));
  XNOR2_X1  g222(.A(KEYINPUT21), .B(G898), .ZN(new_n409));
  AOI21_X1  g223(.A(new_n406), .B1(new_n408), .B2(new_n409), .ZN(new_n410));
  NOR2_X1   g224(.A1(new_n402), .A2(new_n410), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n348), .A2(new_n411), .ZN(new_n412));
  INV_X1    g226(.A(KEYINPUT93), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n412), .A2(new_n413), .ZN(new_n414));
  NAND3_X1  g228(.A1(new_n348), .A2(KEYINPUT93), .A3(new_n411), .ZN(new_n415));
  AOI21_X1  g229(.A(new_n289), .B1(new_n414), .B2(new_n415), .ZN(new_n416));
  INV_X1    g230(.A(G472), .ZN(new_n417));
  INV_X1    g231(.A(KEYINPUT29), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n292), .A2(G210), .ZN(new_n419));
  XNOR2_X1  g233(.A(new_n419), .B(KEYINPUT27), .ZN(new_n420));
  XNOR2_X1  g234(.A(KEYINPUT26), .B(G101), .ZN(new_n421));
  XNOR2_X1  g235(.A(new_n420), .B(new_n421), .ZN(new_n422));
  INV_X1    g236(.A(new_n422), .ZN(new_n423));
  INV_X1    g237(.A(G119), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n424), .A2(G116), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n352), .A2(G119), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n425), .A2(new_n426), .ZN(new_n427));
  XNOR2_X1  g241(.A(KEYINPUT2), .B(G113), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n427), .A2(new_n428), .ZN(new_n429));
  INV_X1    g243(.A(G113), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n430), .A2(KEYINPUT2), .ZN(new_n431));
  INV_X1    g245(.A(KEYINPUT2), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n432), .A2(G113), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n431), .A2(new_n433), .ZN(new_n434));
  XNOR2_X1  g248(.A(G116), .B(G119), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  NAND3_X1  g250(.A1(new_n429), .A2(new_n436), .A3(KEYINPUT67), .ZN(new_n437));
  INV_X1    g251(.A(KEYINPUT67), .ZN(new_n438));
  NAND3_X1  g252(.A1(new_n427), .A2(new_n428), .A3(new_n438), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n437), .A2(new_n439), .ZN(new_n440));
  NAND3_X1  g254(.A1(new_n236), .A2(new_n263), .A3(new_n237), .ZN(new_n441));
  NOR2_X1   g255(.A1(new_n226), .A2(G137), .ZN(new_n442));
  NOR2_X1   g256(.A1(new_n228), .A2(G134), .ZN(new_n443));
  OAI21_X1  g257(.A(G131), .B1(new_n442), .B2(new_n443), .ZN(new_n444));
  NAND3_X1  g258(.A1(new_n223), .A2(new_n235), .A3(new_n444), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n441), .A2(new_n445), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n446), .A2(KEYINPUT30), .ZN(new_n447));
  NAND3_X1  g261(.A1(new_n260), .A2(KEYINPUT65), .A3(new_n262), .ZN(new_n448));
  INV_X1    g262(.A(new_n448), .ZN(new_n449));
  AOI21_X1  g263(.A(KEYINPUT65), .B1(new_n260), .B2(new_n262), .ZN(new_n450));
  OAI211_X1 g264(.A(new_n237), .B(new_n236), .C1(new_n449), .C2(new_n450), .ZN(new_n451));
  INV_X1    g265(.A(KEYINPUT30), .ZN(new_n452));
  NAND3_X1  g266(.A1(new_n451), .A2(new_n452), .A3(new_n445), .ZN(new_n453));
  AOI21_X1  g267(.A(new_n440), .B1(new_n447), .B2(new_n453), .ZN(new_n454));
  NAND3_X1  g268(.A1(new_n441), .A2(new_n440), .A3(new_n445), .ZN(new_n455));
  INV_X1    g269(.A(new_n455), .ZN(new_n456));
  OAI21_X1  g270(.A(new_n423), .B1(new_n454), .B2(new_n456), .ZN(new_n457));
  AOI21_X1  g271(.A(new_n440), .B1(new_n451), .B2(new_n445), .ZN(new_n458));
  OAI21_X1  g272(.A(KEYINPUT28), .B1(new_n458), .B2(new_n456), .ZN(new_n459));
  INV_X1    g273(.A(new_n440), .ZN(new_n460));
  INV_X1    g274(.A(KEYINPUT68), .ZN(new_n461));
  AOI21_X1  g275(.A(new_n461), .B1(new_n441), .B2(new_n445), .ZN(new_n462));
  INV_X1    g276(.A(new_n462), .ZN(new_n463));
  NAND3_X1  g277(.A1(new_n441), .A2(new_n461), .A3(new_n445), .ZN(new_n464));
  AOI21_X1  g278(.A(new_n460), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  OAI21_X1  g279(.A(new_n459), .B1(new_n465), .B2(KEYINPUT28), .ZN(new_n466));
  OAI211_X1 g280(.A(new_n418), .B(new_n457), .C1(new_n466), .C2(new_n423), .ZN(new_n467));
  INV_X1    g281(.A(KEYINPUT28), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n446), .A2(new_n460), .ZN(new_n469));
  AOI21_X1  g283(.A(new_n468), .B1(new_n469), .B2(new_n455), .ZN(new_n470));
  AND3_X1   g284(.A1(new_n441), .A2(new_n461), .A3(new_n445), .ZN(new_n471));
  OAI21_X1  g285(.A(new_n440), .B1(new_n471), .B2(new_n462), .ZN(new_n472));
  AOI21_X1  g286(.A(new_n470), .B1(new_n468), .B2(new_n472), .ZN(new_n473));
  NOR2_X1   g287(.A1(new_n423), .A2(new_n418), .ZN(new_n474));
  AOI21_X1  g288(.A(new_n407), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  AOI21_X1  g289(.A(new_n417), .B1(new_n467), .B2(new_n475), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n472), .A2(new_n468), .ZN(new_n477));
  AOI21_X1  g291(.A(new_n422), .B1(new_n477), .B2(new_n459), .ZN(new_n478));
  AOI21_X1  g292(.A(new_n452), .B1(new_n441), .B2(new_n445), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n235), .A2(new_n444), .ZN(new_n480));
  AOI21_X1  g294(.A(new_n480), .B1(new_n222), .B2(new_n205), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n260), .A2(new_n262), .ZN(new_n482));
  INV_X1    g296(.A(KEYINPUT65), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n484), .A2(new_n448), .ZN(new_n485));
  AOI21_X1  g299(.A(new_n481), .B1(new_n238), .B2(new_n485), .ZN(new_n486));
  AOI21_X1  g300(.A(new_n479), .B1(new_n486), .B2(new_n452), .ZN(new_n487));
  OAI211_X1 g301(.A(new_n455), .B(new_n422), .C1(new_n487), .C2(new_n440), .ZN(new_n488));
  INV_X1    g302(.A(KEYINPUT31), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n447), .A2(new_n453), .ZN(new_n491));
  AOI21_X1  g305(.A(new_n456), .B1(new_n491), .B2(new_n460), .ZN(new_n492));
  NAND3_X1  g306(.A1(new_n492), .A2(KEYINPUT31), .A3(new_n422), .ZN(new_n493));
  AOI21_X1  g307(.A(new_n478), .B1(new_n490), .B2(new_n493), .ZN(new_n494));
  NOR2_X1   g308(.A1(G472), .A2(G902), .ZN(new_n495));
  INV_X1    g309(.A(new_n495), .ZN(new_n496));
  OAI21_X1  g310(.A(KEYINPUT32), .B1(new_n494), .B2(new_n496), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n466), .A2(new_n423), .ZN(new_n498));
  AOI21_X1  g312(.A(KEYINPUT31), .B1(new_n492), .B2(new_n422), .ZN(new_n499));
  NOR4_X1   g313(.A1(new_n454), .A2(new_n489), .A3(new_n456), .A4(new_n423), .ZN(new_n500));
  OAI21_X1  g314(.A(new_n498), .B1(new_n499), .B2(new_n500), .ZN(new_n501));
  INV_X1    g315(.A(KEYINPUT32), .ZN(new_n502));
  NAND3_X1  g316(.A1(new_n501), .A2(new_n502), .A3(new_n495), .ZN(new_n503));
  AOI21_X1  g317(.A(new_n476), .B1(new_n497), .B2(new_n503), .ZN(new_n504));
  AOI21_X1  g318(.A(new_n375), .B1(new_n190), .B2(G234), .ZN(new_n505));
  INV_X1    g319(.A(new_n505), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n203), .A2(G119), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n424), .A2(G128), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  XNOR2_X1  g323(.A(KEYINPUT24), .B(G110), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  INV_X1    g325(.A(KEYINPUT71), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n507), .A2(new_n512), .ZN(new_n513));
  NAND3_X1  g327(.A1(new_n203), .A2(KEYINPUT71), .A3(G119), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  OR2_X1    g329(.A1(KEYINPUT70), .A2(KEYINPUT23), .ZN(new_n516));
  NAND2_X1  g330(.A1(KEYINPUT70), .A2(KEYINPUT23), .ZN(new_n517));
  AOI22_X1  g331(.A1(new_n516), .A2(new_n517), .B1(new_n424), .B2(G128), .ZN(new_n518));
  INV_X1    g332(.A(KEYINPUT23), .ZN(new_n519));
  OAI22_X1  g333(.A1(new_n515), .A2(new_n518), .B1(new_n519), .B2(new_n507), .ZN(new_n520));
  OAI21_X1  g334(.A(new_n511), .B1(new_n520), .B2(G110), .ZN(new_n521));
  INV_X1    g335(.A(new_n305), .ZN(new_n522));
  NOR2_X1   g336(.A1(new_n313), .A2(new_n522), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n521), .A2(new_n523), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n524), .A2(KEYINPUT73), .ZN(new_n525));
  INV_X1    g339(.A(KEYINPUT73), .ZN(new_n526));
  NAND3_X1  g340(.A1(new_n521), .A2(new_n526), .A3(new_n523), .ZN(new_n527));
  NAND3_X1  g341(.A1(new_n314), .A2(new_n319), .A3(new_n316), .ZN(new_n528));
  NOR2_X1   g342(.A1(new_n509), .A2(new_n510), .ZN(new_n529));
  AOI21_X1  g343(.A(new_n529), .B1(new_n520), .B2(G110), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n528), .A2(new_n530), .ZN(new_n531));
  NAND3_X1  g345(.A1(new_n525), .A2(new_n527), .A3(new_n531), .ZN(new_n532));
  INV_X1    g346(.A(KEYINPUT74), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  XNOR2_X1  g348(.A(KEYINPUT22), .B(G137), .ZN(new_n535));
  AND3_X1   g349(.A1(new_n295), .A2(G221), .A3(G234), .ZN(new_n536));
  XNOR2_X1  g350(.A(new_n535), .B(new_n536), .ZN(new_n537));
  NAND4_X1  g351(.A1(new_n525), .A2(KEYINPUT74), .A3(new_n527), .A4(new_n531), .ZN(new_n538));
  NAND3_X1  g352(.A1(new_n534), .A2(new_n537), .A3(new_n538), .ZN(new_n539));
  INV_X1    g353(.A(new_n537), .ZN(new_n540));
  NAND3_X1  g354(.A1(new_n532), .A2(new_n533), .A3(new_n540), .ZN(new_n541));
  AOI21_X1  g355(.A(new_n407), .B1(new_n539), .B2(new_n541), .ZN(new_n542));
  INV_X1    g356(.A(KEYINPUT25), .ZN(new_n543));
  AOI21_X1  g357(.A(new_n506), .B1(new_n542), .B2(new_n543), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n538), .A2(new_n537), .ZN(new_n545));
  AOI22_X1  g359(.A1(new_n524), .A2(KEYINPUT73), .B1(new_n528), .B2(new_n530), .ZN(new_n546));
  AOI21_X1  g360(.A(KEYINPUT74), .B1(new_n546), .B2(new_n527), .ZN(new_n547));
  NOR2_X1   g361(.A1(new_n545), .A2(new_n547), .ZN(new_n548));
  INV_X1    g362(.A(new_n541), .ZN(new_n549));
  OAI21_X1  g363(.A(new_n190), .B1(new_n548), .B2(new_n549), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n550), .A2(KEYINPUT25), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n544), .A2(new_n551), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n539), .A2(new_n541), .ZN(new_n553));
  NOR2_X1   g367(.A1(new_n505), .A2(G902), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n552), .A2(new_n555), .ZN(new_n556));
  NOR2_X1   g370(.A1(new_n504), .A2(new_n556), .ZN(new_n557));
  OAI21_X1  g371(.A(G214), .B1(G237), .B2(G902), .ZN(new_n558));
  OAI21_X1  g372(.A(G210), .B1(G237), .B2(G902), .ZN(new_n559));
  XNOR2_X1  g373(.A(G110), .B(G122), .ZN(new_n560));
  INV_X1    g374(.A(new_n560), .ZN(new_n561));
  AOI211_X1 g375(.A(new_n250), .B(new_n440), .C1(new_n255), .C2(new_n253), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n435), .A2(KEYINPUT5), .ZN(new_n563));
  OAI211_X1 g377(.A(new_n563), .B(G113), .C1(KEYINPUT5), .C2(new_n425), .ZN(new_n564));
  NAND3_X1  g378(.A1(new_n564), .A2(new_n218), .A3(new_n436), .ZN(new_n565));
  INV_X1    g379(.A(new_n565), .ZN(new_n566));
  OAI21_X1  g380(.A(new_n561), .B1(new_n562), .B2(new_n566), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n256), .A2(new_n460), .ZN(new_n568));
  NAND3_X1  g382(.A1(new_n568), .A2(new_n565), .A3(new_n560), .ZN(new_n569));
  INV_X1    g383(.A(KEYINPUT80), .ZN(new_n570));
  INV_X1    g384(.A(KEYINPUT6), .ZN(new_n571));
  NOR2_X1   g385(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  NAND3_X1  g386(.A1(new_n567), .A2(new_n569), .A3(new_n572), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n482), .A2(G125), .ZN(new_n574));
  NAND3_X1  g388(.A1(new_n222), .A2(new_n311), .A3(new_n205), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n295), .A2(G224), .ZN(new_n577));
  XOR2_X1   g391(.A(new_n576), .B(new_n577), .Z(new_n578));
  OAI221_X1 g392(.A(new_n561), .B1(new_n570), .B2(new_n571), .C1(new_n562), .C2(new_n566), .ZN(new_n579));
  NAND3_X1  g393(.A1(new_n573), .A2(new_n578), .A3(new_n579), .ZN(new_n580));
  INV_X1    g394(.A(KEYINPUT81), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  NAND4_X1  g396(.A1(new_n573), .A2(new_n579), .A3(KEYINPUT81), .A4(new_n578), .ZN(new_n583));
  INV_X1    g397(.A(new_n569), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n577), .A2(KEYINPUT7), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n575), .A2(KEYINPUT83), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n586), .A2(new_n574), .ZN(new_n587));
  NOR2_X1   g401(.A1(new_n575), .A2(KEYINPUT83), .ZN(new_n588));
  OAI21_X1  g402(.A(new_n585), .B1(new_n587), .B2(new_n588), .ZN(new_n589));
  XOR2_X1   g403(.A(KEYINPUT82), .B(KEYINPUT8), .Z(new_n590));
  XNOR2_X1  g404(.A(new_n590), .B(new_n560), .ZN(new_n591));
  AOI21_X1  g405(.A(new_n218), .B1(new_n436), .B2(new_n564), .ZN(new_n592));
  OAI21_X1  g406(.A(new_n591), .B1(new_n566), .B2(new_n592), .ZN(new_n593));
  NAND4_X1  g407(.A1(new_n574), .A2(new_n575), .A3(KEYINPUT7), .A4(new_n577), .ZN(new_n594));
  NAND3_X1  g408(.A1(new_n589), .A2(new_n593), .A3(new_n594), .ZN(new_n595));
  OAI21_X1  g409(.A(new_n278), .B1(new_n584), .B2(new_n595), .ZN(new_n596));
  INV_X1    g410(.A(new_n596), .ZN(new_n597));
  AND4_X1   g411(.A1(new_n559), .A2(new_n582), .A3(new_n583), .A4(new_n597), .ZN(new_n598));
  AOI21_X1  g412(.A(new_n596), .B1(new_n580), .B2(new_n581), .ZN(new_n599));
  AOI21_X1  g413(.A(new_n559), .B1(new_n599), .B2(new_n583), .ZN(new_n600));
  OAI21_X1  g414(.A(new_n558), .B1(new_n598), .B2(new_n600), .ZN(new_n601));
  INV_X1    g415(.A(new_n601), .ZN(new_n602));
  NAND3_X1  g416(.A1(new_n416), .A2(new_n557), .A3(new_n602), .ZN(new_n603));
  XNOR2_X1  g417(.A(new_n603), .B(G101), .ZN(G3));
  NOR2_X1   g418(.A1(new_n390), .A2(new_n391), .ZN(new_n605));
  AOI21_X1  g419(.A(KEYINPUT95), .B1(new_n374), .B2(new_n389), .ZN(new_n606));
  INV_X1    g420(.A(KEYINPUT33), .ZN(new_n607));
  NOR2_X1   g421(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n605), .A2(new_n608), .ZN(new_n609));
  OAI22_X1  g423(.A1(new_n390), .A2(new_n391), .B1(new_n606), .B2(new_n607), .ZN(new_n610));
  NAND3_X1  g424(.A1(new_n609), .A2(new_n190), .A3(new_n610), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n611), .A2(G478), .ZN(new_n612));
  OR2_X1    g426(.A1(new_n392), .A2(G478), .ZN(new_n613));
  AND2_X1   g427(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n614), .A2(new_n347), .ZN(new_n615));
  INV_X1    g429(.A(KEYINPUT94), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n601), .A2(new_n616), .ZN(new_n617));
  OAI211_X1 g431(.A(KEYINPUT94), .B(new_n558), .C1(new_n598), .C2(new_n600), .ZN(new_n618));
  AOI211_X1 g432(.A(new_n410), .B(new_n615), .C1(new_n617), .C2(new_n618), .ZN(new_n619));
  OAI21_X1  g433(.A(G472), .B1(new_n494), .B2(new_n407), .ZN(new_n620));
  OAI21_X1  g434(.A(new_n620), .B1(new_n496), .B2(new_n494), .ZN(new_n621));
  NOR3_X1   g435(.A1(new_n621), .A2(new_n556), .A3(new_n289), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n619), .A2(new_n622), .ZN(new_n623));
  XOR2_X1   g437(.A(KEYINPUT34), .B(G104), .Z(new_n624));
  XNOR2_X1  g438(.A(new_n623), .B(new_n624), .ZN(G6));
  INV_X1    g439(.A(new_n410), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n617), .A2(new_n618), .ZN(new_n627));
  AOI21_X1  g441(.A(new_n345), .B1(new_n399), .B2(new_n401), .ZN(new_n628));
  INV_X1    g442(.A(KEYINPUT96), .ZN(new_n629));
  NAND3_X1  g443(.A1(new_n336), .A2(new_n629), .A3(KEYINPUT20), .ZN(new_n630));
  NAND3_X1  g444(.A1(new_n337), .A2(KEYINPUT96), .A3(new_n339), .ZN(new_n631));
  AND3_X1   g445(.A1(new_n628), .A2(new_n630), .A3(new_n631), .ZN(new_n632));
  AND4_X1   g446(.A1(new_n626), .A2(new_n627), .A3(new_n622), .A4(new_n632), .ZN(new_n633));
  XNOR2_X1  g447(.A(KEYINPUT35), .B(G107), .ZN(new_n634));
  XNOR2_X1  g448(.A(new_n633), .B(new_n634), .ZN(G9));
  INV_X1    g449(.A(KEYINPUT97), .ZN(new_n636));
  NOR2_X1   g450(.A1(new_n537), .A2(KEYINPUT36), .ZN(new_n637));
  XNOR2_X1  g451(.A(new_n532), .B(new_n637), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n638), .A2(new_n554), .ZN(new_n639));
  AOI21_X1  g453(.A(new_n636), .B1(new_n552), .B2(new_n639), .ZN(new_n640));
  INV_X1    g454(.A(new_n639), .ZN(new_n641));
  AOI211_X1 g455(.A(KEYINPUT97), .B(new_n641), .C1(new_n544), .C2(new_n551), .ZN(new_n642));
  NOR3_X1   g456(.A1(new_n640), .A2(new_n642), .A3(new_n621), .ZN(new_n643));
  NAND3_X1  g457(.A1(new_n416), .A2(new_n602), .A3(new_n643), .ZN(new_n644));
  XOR2_X1   g458(.A(KEYINPUT37), .B(G110), .Z(new_n645));
  XNOR2_X1  g459(.A(new_n644), .B(new_n645), .ZN(G12));
  INV_X1    g460(.A(new_n408), .ZN(new_n647));
  XNOR2_X1  g461(.A(KEYINPUT98), .B(G900), .ZN(new_n648));
  OAI21_X1  g462(.A(new_n405), .B1(new_n647), .B2(new_n648), .ZN(new_n649));
  NAND4_X1  g463(.A1(new_n628), .A2(new_n631), .A3(new_n630), .A4(new_n649), .ZN(new_n650));
  NOR3_X1   g464(.A1(new_n504), .A2(new_n289), .A3(new_n650), .ZN(new_n651));
  NOR2_X1   g465(.A1(new_n640), .A2(new_n642), .ZN(new_n652));
  NAND3_X1  g466(.A1(new_n582), .A2(new_n583), .A3(new_n597), .ZN(new_n653));
  INV_X1    g467(.A(new_n559), .ZN(new_n654));
  NAND2_X1  g468(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  NAND3_X1  g469(.A1(new_n599), .A2(new_n559), .A3(new_n583), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  AOI21_X1  g471(.A(KEYINPUT94), .B1(new_n657), .B2(new_n558), .ZN(new_n658));
  INV_X1    g472(.A(new_n558), .ZN(new_n659));
  AOI211_X1 g473(.A(new_n616), .B(new_n659), .C1(new_n655), .C2(new_n656), .ZN(new_n660));
  OAI211_X1 g474(.A(new_n651), .B(new_n652), .C1(new_n658), .C2(new_n660), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n661), .A2(KEYINPUT99), .ZN(new_n662));
  INV_X1    g476(.A(KEYINPUT99), .ZN(new_n663));
  NAND4_X1  g477(.A1(new_n627), .A2(new_n663), .A3(new_n652), .A4(new_n651), .ZN(new_n664));
  NAND2_X1  g478(.A1(new_n662), .A2(new_n664), .ZN(new_n665));
  XNOR2_X1  g479(.A(new_n665), .B(G128), .ZN(G30));
  AOI21_X1  g480(.A(new_n641), .B1(new_n544), .B2(new_n551), .ZN(new_n667));
  NAND4_X1  g481(.A1(new_n667), .A2(new_n558), .A3(new_n347), .A4(new_n402), .ZN(new_n668));
  AND2_X1   g482(.A1(new_n497), .A2(new_n503), .ZN(new_n669));
  AND2_X1   g483(.A1(new_n469), .A2(new_n455), .ZN(new_n670));
  OAI21_X1  g484(.A(new_n488), .B1(new_n422), .B2(new_n670), .ZN(new_n671));
  AOI21_X1  g485(.A(new_n417), .B1(new_n671), .B2(new_n278), .ZN(new_n672));
  NOR2_X1   g486(.A1(new_n669), .A2(new_n672), .ZN(new_n673));
  XNOR2_X1  g487(.A(new_n649), .B(KEYINPUT39), .ZN(new_n674));
  OAI211_X1 g488(.A(new_n189), .B(new_n674), .C1(new_n281), .C2(new_n288), .ZN(new_n675));
  AOI211_X1 g489(.A(new_n668), .B(new_n673), .C1(KEYINPUT40), .C2(new_n675), .ZN(new_n676));
  NOR2_X1   g490(.A1(new_n598), .A2(new_n600), .ZN(new_n677));
  XNOR2_X1  g491(.A(new_n677), .B(KEYINPUT38), .ZN(new_n678));
  INV_X1    g492(.A(new_n678), .ZN(new_n679));
  OAI211_X1 g493(.A(new_n676), .B(new_n679), .C1(KEYINPUT40), .C2(new_n675), .ZN(new_n680));
  XNOR2_X1  g494(.A(KEYINPUT100), .B(G143), .ZN(new_n681));
  XNOR2_X1  g495(.A(new_n680), .B(new_n681), .ZN(G45));
  NAND4_X1  g496(.A1(new_n347), .A2(new_n612), .A3(new_n613), .A4(new_n649), .ZN(new_n683));
  NOR3_X1   g497(.A1(new_n683), .A2(new_n504), .A3(new_n289), .ZN(new_n684));
  NAND3_X1  g498(.A1(new_n627), .A2(new_n652), .A3(new_n684), .ZN(new_n685));
  XNOR2_X1  g499(.A(new_n685), .B(G146), .ZN(G48));
  NAND2_X1  g500(.A1(new_n612), .A2(new_n613), .ZN(new_n687));
  NOR2_X1   g501(.A1(new_n687), .A2(new_n348), .ZN(new_n688));
  INV_X1    g502(.A(new_n275), .ZN(new_n689));
  AOI21_X1  g503(.A(new_n407), .B1(new_n689), .B2(new_n271), .ZN(new_n690));
  OR2_X1    g504(.A1(new_n690), .A2(new_n277), .ZN(new_n691));
  NAND3_X1  g505(.A1(new_n691), .A2(new_n189), .A3(new_n276), .ZN(new_n692));
  NOR3_X1   g506(.A1(new_n692), .A2(new_n504), .A3(new_n556), .ZN(new_n693));
  NAND4_X1  g507(.A1(new_n627), .A2(new_n626), .A3(new_n688), .A4(new_n693), .ZN(new_n694));
  XNOR2_X1  g508(.A(KEYINPUT41), .B(G113), .ZN(new_n695));
  XNOR2_X1  g509(.A(new_n694), .B(new_n695), .ZN(G15));
  NAND4_X1  g510(.A1(new_n627), .A2(new_n626), .A3(new_n632), .A4(new_n693), .ZN(new_n697));
  XNOR2_X1  g511(.A(new_n697), .B(G116), .ZN(G18));
  AOI21_X1  g512(.A(new_n504), .B1(new_n414), .B2(new_n415), .ZN(new_n699));
  INV_X1    g513(.A(new_n692), .ZN(new_n700));
  AOI21_X1  g514(.A(KEYINPUT101), .B1(new_n627), .B2(new_n700), .ZN(new_n701));
  INV_X1    g515(.A(KEYINPUT101), .ZN(new_n702));
  AOI211_X1 g516(.A(new_n702), .B(new_n692), .C1(new_n617), .C2(new_n618), .ZN(new_n703));
  OAI211_X1 g517(.A(new_n652), .B(new_n699), .C1(new_n701), .C2(new_n703), .ZN(new_n704));
  XOR2_X1   g518(.A(KEYINPUT102), .B(G119), .Z(new_n705));
  XNOR2_X1  g519(.A(new_n704), .B(new_n705), .ZN(G21));
  NAND4_X1  g520(.A1(new_n691), .A2(new_n626), .A3(new_n189), .A4(new_n276), .ZN(new_n707));
  NAND2_X1  g521(.A1(new_n620), .A2(KEYINPUT103), .ZN(new_n708));
  NOR2_X1   g522(.A1(new_n499), .A2(new_n500), .ZN(new_n709));
  NOR2_X1   g523(.A1(new_n473), .A2(new_n422), .ZN(new_n710));
  OAI21_X1  g524(.A(new_n495), .B1(new_n709), .B2(new_n710), .ZN(new_n711));
  NAND2_X1  g525(.A1(new_n708), .A2(new_n711), .ZN(new_n712));
  NOR2_X1   g526(.A1(new_n620), .A2(KEYINPUT103), .ZN(new_n713));
  NOR4_X1   g527(.A1(new_n707), .A2(new_n712), .A3(new_n556), .A4(new_n713), .ZN(new_n714));
  NAND2_X1  g528(.A1(new_n347), .A2(new_n402), .ZN(new_n715));
  AOI21_X1  g529(.A(new_n715), .B1(new_n617), .B2(new_n618), .ZN(new_n716));
  NAND2_X1  g530(.A1(new_n714), .A2(new_n716), .ZN(new_n717));
  XNOR2_X1  g531(.A(new_n717), .B(G122), .ZN(G24));
  NOR3_X1   g532(.A1(new_n712), .A2(new_n667), .A3(new_n713), .ZN(new_n719));
  INV_X1    g533(.A(new_n683), .ZN(new_n720));
  AND2_X1   g534(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  OAI21_X1  g535(.A(new_n721), .B1(new_n701), .B2(new_n703), .ZN(new_n722));
  XNOR2_X1  g536(.A(new_n722), .B(G125), .ZN(G27));
  INV_X1    g537(.A(new_n189), .ZN(new_n724));
  NOR3_X1   g538(.A1(new_n657), .A2(new_n659), .A3(new_n724), .ZN(new_n725));
  INV_X1    g539(.A(new_n281), .ZN(new_n726));
  NAND2_X1  g540(.A1(new_n286), .A2(new_n287), .ZN(new_n727));
  INV_X1    g541(.A(new_n282), .ZN(new_n728));
  NAND2_X1  g542(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  OAI21_X1  g543(.A(KEYINPUT104), .B1(new_n729), .B2(new_n277), .ZN(new_n730));
  INV_X1    g544(.A(KEYINPUT104), .ZN(new_n731));
  NAND2_X1  g545(.A1(new_n288), .A2(new_n731), .ZN(new_n732));
  NAND3_X1  g546(.A1(new_n726), .A2(new_n730), .A3(new_n732), .ZN(new_n733));
  NAND4_X1  g547(.A1(new_n725), .A2(new_n720), .A3(new_n557), .A4(new_n733), .ZN(new_n734));
  INV_X1    g548(.A(KEYINPUT42), .ZN(new_n735));
  NAND2_X1  g549(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  AND4_X1   g550(.A1(new_n558), .A2(new_n733), .A3(new_n677), .A4(new_n189), .ZN(new_n737));
  NAND4_X1  g551(.A1(new_n737), .A2(KEYINPUT42), .A3(new_n557), .A4(new_n720), .ZN(new_n738));
  NAND2_X1  g552(.A1(new_n736), .A2(new_n738), .ZN(new_n739));
  XNOR2_X1  g553(.A(new_n739), .B(G131), .ZN(G33));
  NAND4_X1  g554(.A1(new_n737), .A2(new_n557), .A3(new_n632), .A4(new_n649), .ZN(new_n741));
  XOR2_X1   g555(.A(KEYINPUT105), .B(G134), .Z(new_n742));
  XNOR2_X1  g556(.A(new_n741), .B(new_n742), .ZN(G36));
  NOR2_X1   g557(.A1(new_n657), .A2(new_n659), .ZN(new_n744));
  INV_X1    g558(.A(new_n744), .ZN(new_n745));
  XNOR2_X1  g559(.A(new_n347), .B(KEYINPUT106), .ZN(new_n746));
  NOR2_X1   g560(.A1(new_n746), .A2(new_n687), .ZN(new_n747));
  NAND2_X1  g561(.A1(new_n747), .A2(KEYINPUT43), .ZN(new_n748));
  NOR2_X1   g562(.A1(new_n687), .A2(new_n347), .ZN(new_n749));
  OAI21_X1  g563(.A(new_n748), .B1(KEYINPUT43), .B2(new_n749), .ZN(new_n750));
  INV_X1    g564(.A(new_n667), .ZN(new_n751));
  NAND3_X1  g565(.A1(new_n750), .A2(new_n621), .A3(new_n751), .ZN(new_n752));
  INV_X1    g566(.A(new_n752), .ZN(new_n753));
  AOI21_X1  g567(.A(new_n745), .B1(new_n753), .B2(KEYINPUT44), .ZN(new_n754));
  XOR2_X1   g568(.A(new_n729), .B(KEYINPUT45), .Z(new_n755));
  NOR2_X1   g569(.A1(new_n755), .A2(new_n277), .ZN(new_n756));
  NOR2_X1   g570(.A1(new_n756), .A2(new_n279), .ZN(new_n757));
  AOI22_X1  g571(.A1(new_n757), .A2(KEYINPUT46), .B1(new_n690), .B2(new_n191), .ZN(new_n758));
  OAI21_X1  g572(.A(new_n758), .B1(KEYINPUT46), .B2(new_n757), .ZN(new_n759));
  NAND3_X1  g573(.A1(new_n759), .A2(new_n189), .A3(new_n674), .ZN(new_n760));
  INV_X1    g574(.A(new_n760), .ZN(new_n761));
  OAI211_X1 g575(.A(new_n754), .B(new_n761), .C1(KEYINPUT44), .C2(new_n753), .ZN(new_n762));
  XNOR2_X1  g576(.A(new_n762), .B(G137), .ZN(G39));
  NAND2_X1  g577(.A1(KEYINPUT107), .A2(KEYINPUT47), .ZN(new_n764));
  NAND3_X1  g578(.A1(new_n759), .A2(new_n189), .A3(new_n764), .ZN(new_n765));
  NOR2_X1   g579(.A1(KEYINPUT107), .A2(KEYINPUT47), .ZN(new_n766));
  XNOR2_X1  g580(.A(new_n765), .B(new_n766), .ZN(new_n767));
  AND4_X1   g581(.A1(new_n556), .A2(new_n744), .A3(new_n504), .A4(new_n720), .ZN(new_n768));
  AND2_X1   g582(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  XOR2_X1   g583(.A(new_n769), .B(G140), .Z(G42));
  AND2_X1   g584(.A1(new_n750), .A2(new_n406), .ZN(new_n771));
  AND2_X1   g585(.A1(new_n691), .A2(new_n276), .ZN(new_n772));
  AND2_X1   g586(.A1(new_n725), .A2(new_n772), .ZN(new_n773));
  NAND2_X1  g587(.A1(new_n771), .A2(new_n773), .ZN(new_n774));
  INV_X1    g588(.A(KEYINPUT117), .ZN(new_n775));
  XNOR2_X1  g589(.A(new_n774), .B(new_n775), .ZN(new_n776));
  NAND2_X1  g590(.A1(new_n776), .A2(new_n557), .ZN(new_n777));
  AND2_X1   g591(.A1(new_n777), .A2(KEYINPUT119), .ZN(new_n778));
  INV_X1    g592(.A(KEYINPUT48), .ZN(new_n779));
  NAND2_X1  g593(.A1(new_n778), .A2(new_n779), .ZN(new_n780));
  OR3_X1    g594(.A1(new_n712), .A2(new_n556), .A3(new_n713), .ZN(new_n781));
  INV_X1    g595(.A(new_n781), .ZN(new_n782));
  NAND2_X1  g596(.A1(new_n771), .A2(new_n782), .ZN(new_n783));
  NOR2_X1   g597(.A1(new_n701), .A2(new_n703), .ZN(new_n784));
  NOR2_X1   g598(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  OR2_X1    g599(.A1(new_n669), .A2(new_n672), .ZN(new_n786));
  NOR3_X1   g600(.A1(new_n786), .A2(new_n556), .A3(new_n405), .ZN(new_n787));
  AND3_X1   g601(.A1(new_n773), .A2(new_n688), .A3(new_n787), .ZN(new_n788));
  NAND2_X1  g602(.A1(new_n295), .A2(G952), .ZN(new_n789));
  XOR2_X1   g603(.A(new_n789), .B(KEYINPUT118), .Z(new_n790));
  NOR3_X1   g604(.A1(new_n785), .A2(new_n788), .A3(new_n790), .ZN(new_n791));
  OAI21_X1  g605(.A(KEYINPUT48), .B1(new_n777), .B2(KEYINPUT119), .ZN(new_n792));
  OAI211_X1 g606(.A(new_n780), .B(new_n791), .C1(new_n778), .C2(new_n792), .ZN(new_n793));
  INV_X1    g607(.A(KEYINPUT51), .ZN(new_n794));
  NOR4_X1   g608(.A1(new_n783), .A2(new_n558), .A3(new_n679), .A4(new_n692), .ZN(new_n795));
  XNOR2_X1  g609(.A(new_n795), .B(KEYINPUT50), .ZN(new_n796));
  INV_X1    g610(.A(new_n783), .ZN(new_n797));
  NAND2_X1  g611(.A1(new_n772), .A2(new_n724), .ZN(new_n798));
  INV_X1    g612(.A(new_n798), .ZN(new_n799));
  OAI211_X1 g613(.A(new_n744), .B(new_n797), .C1(new_n767), .C2(new_n799), .ZN(new_n800));
  NAND2_X1  g614(.A1(new_n776), .A2(new_n719), .ZN(new_n801));
  NAND4_X1  g615(.A1(new_n787), .A2(new_n773), .A3(new_n348), .A4(new_n687), .ZN(new_n802));
  NAND4_X1  g616(.A1(new_n796), .A2(new_n800), .A3(new_n801), .A4(new_n802), .ZN(new_n803));
  AOI21_X1  g617(.A(new_n793), .B1(new_n794), .B2(new_n803), .ZN(new_n804));
  INV_X1    g618(.A(KEYINPUT116), .ZN(new_n805));
  AND2_X1   g619(.A1(new_n649), .A2(new_n189), .ZN(new_n806));
  NAND3_X1  g620(.A1(new_n733), .A2(new_n667), .A3(new_n806), .ZN(new_n807));
  AND2_X1   g621(.A1(new_n807), .A2(KEYINPUT112), .ZN(new_n808));
  NOR2_X1   g622(.A1(new_n807), .A2(KEYINPUT112), .ZN(new_n809));
  OAI211_X1 g623(.A(new_n786), .B(new_n716), .C1(new_n808), .C2(new_n809), .ZN(new_n810));
  NAND4_X1  g624(.A1(new_n722), .A2(new_n665), .A3(new_n685), .A4(new_n810), .ZN(new_n811));
  INV_X1    g625(.A(KEYINPUT52), .ZN(new_n812));
  NAND2_X1  g626(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  INV_X1    g627(.A(new_n685), .ZN(new_n814));
  AOI21_X1  g628(.A(new_n814), .B1(new_n664), .B2(new_n662), .ZN(new_n815));
  NAND4_X1  g629(.A1(new_n815), .A2(KEYINPUT52), .A3(new_n722), .A4(new_n810), .ZN(new_n816));
  NAND2_X1  g630(.A1(new_n813), .A2(new_n816), .ZN(new_n817));
  INV_X1    g631(.A(KEYINPUT113), .ZN(new_n818));
  NAND2_X1  g632(.A1(new_n817), .A2(new_n818), .ZN(new_n819));
  NAND3_X1  g633(.A1(new_n813), .A2(KEYINPUT113), .A3(new_n816), .ZN(new_n820));
  AND3_X1   g634(.A1(new_n717), .A2(new_n694), .A3(new_n697), .ZN(new_n821));
  NAND3_X1  g635(.A1(new_n821), .A2(new_n704), .A3(new_n739), .ZN(new_n822));
  XNOR2_X1  g636(.A(new_n688), .B(KEYINPUT109), .ZN(new_n823));
  NOR2_X1   g637(.A1(new_n601), .A2(new_n410), .ZN(new_n824));
  NAND3_X1  g638(.A1(new_n823), .A2(new_n622), .A3(new_n824), .ZN(new_n825));
  OAI211_X1 g639(.A(new_n416), .B(new_n602), .C1(new_n557), .C2(new_n643), .ZN(new_n826));
  AND2_X1   g640(.A1(new_n628), .A2(new_n340), .ZN(new_n827));
  NAND3_X1  g641(.A1(new_n824), .A2(KEYINPUT110), .A3(new_n827), .ZN(new_n828));
  NAND2_X1  g642(.A1(new_n828), .A2(new_n622), .ZN(new_n829));
  AOI21_X1  g643(.A(KEYINPUT110), .B1(new_n824), .B2(new_n827), .ZN(new_n830));
  OAI211_X1 g644(.A(new_n825), .B(new_n826), .C1(new_n829), .C2(new_n830), .ZN(new_n831));
  AND4_X1   g645(.A1(new_n346), .A2(new_n399), .A3(new_n401), .A4(new_n649), .ZN(new_n832));
  NAND3_X1  g646(.A1(new_n832), .A2(new_n630), .A3(new_n631), .ZN(new_n833));
  XNOR2_X1  g647(.A(new_n833), .B(KEYINPUT111), .ZN(new_n834));
  NOR2_X1   g648(.A1(new_n504), .A2(new_n289), .ZN(new_n835));
  NAND4_X1  g649(.A1(new_n834), .A2(new_n652), .A3(new_n835), .A4(new_n744), .ZN(new_n836));
  NAND3_X1  g650(.A1(new_n737), .A2(new_n720), .A3(new_n719), .ZN(new_n837));
  NAND3_X1  g651(.A1(new_n836), .A2(new_n741), .A3(new_n837), .ZN(new_n838));
  NOR3_X1   g652(.A1(new_n822), .A2(new_n831), .A3(new_n838), .ZN(new_n839));
  NAND4_X1  g653(.A1(new_n819), .A2(KEYINPUT53), .A3(new_n820), .A4(new_n839), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n817), .A2(new_n839), .ZN(new_n841));
  INV_X1    g655(.A(KEYINPUT53), .ZN(new_n842));
  NAND2_X1  g656(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  NAND2_X1  g657(.A1(new_n840), .A2(new_n843), .ZN(new_n844));
  INV_X1    g658(.A(KEYINPUT114), .ZN(new_n845));
  NAND3_X1  g659(.A1(new_n844), .A2(new_n845), .A3(KEYINPUT54), .ZN(new_n846));
  NAND3_X1  g660(.A1(new_n819), .A2(new_n820), .A3(new_n839), .ZN(new_n847));
  NAND2_X1  g661(.A1(new_n847), .A2(new_n842), .ZN(new_n848));
  INV_X1    g662(.A(KEYINPUT54), .ZN(new_n849));
  INV_X1    g663(.A(new_n817), .ZN(new_n850));
  NAND2_X1  g664(.A1(new_n822), .A2(KEYINPUT115), .ZN(new_n851));
  INV_X1    g665(.A(KEYINPUT115), .ZN(new_n852));
  NAND4_X1  g666(.A1(new_n821), .A2(new_n704), .A3(new_n852), .A4(new_n739), .ZN(new_n853));
  NOR3_X1   g667(.A1(new_n831), .A2(new_n838), .A3(new_n842), .ZN(new_n854));
  NAND3_X1  g668(.A1(new_n851), .A2(new_n853), .A3(new_n854), .ZN(new_n855));
  NOR2_X1   g669(.A1(new_n850), .A2(new_n855), .ZN(new_n856));
  INV_X1    g670(.A(new_n856), .ZN(new_n857));
  NAND3_X1  g671(.A1(new_n848), .A2(new_n849), .A3(new_n857), .ZN(new_n858));
  NAND2_X1  g672(.A1(new_n846), .A2(new_n858), .ZN(new_n859));
  AOI21_X1  g673(.A(new_n849), .B1(new_n840), .B2(new_n843), .ZN(new_n860));
  NOR2_X1   g674(.A1(new_n860), .A2(new_n845), .ZN(new_n861));
  OAI21_X1  g675(.A(new_n805), .B1(new_n859), .B2(new_n861), .ZN(new_n862));
  AOI21_X1  g676(.A(new_n856), .B1(new_n847), .B2(new_n842), .ZN(new_n863));
  AOI22_X1  g677(.A1(new_n845), .A2(new_n860), .B1(new_n863), .B2(new_n849), .ZN(new_n864));
  NAND2_X1  g678(.A1(new_n844), .A2(KEYINPUT54), .ZN(new_n865));
  NAND2_X1  g679(.A1(new_n865), .A2(KEYINPUT114), .ZN(new_n866));
  NAND3_X1  g680(.A1(new_n864), .A2(KEYINPUT116), .A3(new_n866), .ZN(new_n867));
  OR2_X1    g681(.A1(new_n803), .A2(new_n794), .ZN(new_n868));
  NAND4_X1  g682(.A1(new_n804), .A2(new_n862), .A3(new_n867), .A4(new_n868), .ZN(new_n869));
  OAI21_X1  g683(.A(new_n869), .B1(G952), .B2(G953), .ZN(new_n870));
  XNOR2_X1  g684(.A(new_n772), .B(KEYINPUT49), .ZN(new_n871));
  AND2_X1   g685(.A1(new_n871), .A2(new_n747), .ZN(new_n872));
  NOR3_X1   g686(.A1(new_n556), .A2(new_n659), .A3(new_n724), .ZN(new_n873));
  XNOR2_X1  g687(.A(new_n873), .B(KEYINPUT108), .ZN(new_n874));
  NAND4_X1  g688(.A1(new_n872), .A2(new_n874), .A3(new_n678), .A4(new_n673), .ZN(new_n875));
  NAND2_X1  g689(.A1(new_n870), .A2(new_n875), .ZN(new_n876));
  INV_X1    g690(.A(KEYINPUT120), .ZN(new_n877));
  NAND2_X1  g691(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  NAND3_X1  g692(.A1(new_n870), .A2(KEYINPUT120), .A3(new_n875), .ZN(new_n879));
  NAND2_X1  g693(.A1(new_n878), .A2(new_n879), .ZN(G75));
  NOR2_X1   g694(.A1(new_n295), .A2(G952), .ZN(new_n881));
  INV_X1    g695(.A(new_n881), .ZN(new_n882));
  NOR2_X1   g696(.A1(new_n863), .A2(new_n190), .ZN(new_n883));
  AOI21_X1  g697(.A(KEYINPUT56), .B1(new_n883), .B2(new_n654), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n573), .A2(new_n579), .ZN(new_n885));
  XNOR2_X1  g699(.A(new_n885), .B(new_n578), .ZN(new_n886));
  XNOR2_X1  g700(.A(new_n886), .B(KEYINPUT55), .ZN(new_n887));
  OAI21_X1  g701(.A(new_n882), .B1(new_n884), .B2(new_n887), .ZN(new_n888));
  AOI21_X1  g702(.A(new_n888), .B1(new_n884), .B2(new_n887), .ZN(G51));
  XNOR2_X1  g703(.A(new_n863), .B(new_n849), .ZN(new_n890));
  XNOR2_X1  g704(.A(new_n279), .B(KEYINPUT57), .ZN(new_n891));
  NAND2_X1  g705(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  OAI21_X1  g706(.A(new_n892), .B1(new_n275), .B2(new_n272), .ZN(new_n893));
  NAND2_X1  g707(.A1(new_n883), .A2(new_n756), .ZN(new_n894));
  AOI21_X1  g708(.A(new_n881), .B1(new_n893), .B2(new_n894), .ZN(G54));
  NAND3_X1  g709(.A1(new_n883), .A2(KEYINPUT58), .A3(G475), .ZN(new_n896));
  INV_X1    g710(.A(new_n334), .ZN(new_n897));
  NAND2_X1  g711(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  INV_X1    g712(.A(new_n898), .ZN(new_n899));
  AND2_X1   g713(.A1(new_n899), .A2(KEYINPUT121), .ZN(new_n900));
  NOR2_X1   g714(.A1(new_n899), .A2(KEYINPUT121), .ZN(new_n901));
  OAI21_X1  g715(.A(new_n882), .B1(new_n896), .B2(new_n897), .ZN(new_n902));
  NOR3_X1   g716(.A1(new_n900), .A2(new_n901), .A3(new_n902), .ZN(G60));
  NAND2_X1  g717(.A1(G478), .A2(G902), .ZN(new_n904));
  XOR2_X1   g718(.A(new_n904), .B(KEYINPUT59), .Z(new_n905));
  INV_X1    g719(.A(new_n905), .ZN(new_n906));
  NOR3_X1   g720(.A1(new_n859), .A2(new_n805), .A3(new_n861), .ZN(new_n907));
  AOI21_X1  g721(.A(KEYINPUT116), .B1(new_n864), .B2(new_n866), .ZN(new_n908));
  OAI21_X1  g722(.A(new_n906), .B1(new_n907), .B2(new_n908), .ZN(new_n909));
  INV_X1    g723(.A(KEYINPUT122), .ZN(new_n910));
  NAND2_X1  g724(.A1(new_n609), .A2(new_n610), .ZN(new_n911));
  NAND3_X1  g725(.A1(new_n909), .A2(new_n910), .A3(new_n911), .ZN(new_n912));
  AOI21_X1  g726(.A(new_n905), .B1(new_n862), .B2(new_n867), .ZN(new_n913));
  INV_X1    g727(.A(new_n911), .ZN(new_n914));
  OAI21_X1  g728(.A(KEYINPUT122), .B1(new_n913), .B2(new_n914), .ZN(new_n915));
  NOR2_X1   g729(.A1(new_n911), .A2(new_n905), .ZN(new_n916));
  AOI21_X1  g730(.A(new_n881), .B1(new_n890), .B2(new_n916), .ZN(new_n917));
  NAND3_X1  g731(.A1(new_n912), .A2(new_n915), .A3(new_n917), .ZN(new_n918));
  NAND2_X1  g732(.A1(new_n918), .A2(KEYINPUT123), .ZN(new_n919));
  INV_X1    g733(.A(KEYINPUT123), .ZN(new_n920));
  NAND4_X1  g734(.A1(new_n912), .A2(new_n915), .A3(new_n920), .A4(new_n917), .ZN(new_n921));
  NAND2_X1  g735(.A1(new_n919), .A2(new_n921), .ZN(G63));
  NAND2_X1  g736(.A1(G217), .A2(G902), .ZN(new_n923));
  XNOR2_X1  g737(.A(new_n923), .B(KEYINPUT60), .ZN(new_n924));
  OR2_X1    g738(.A1(new_n863), .A2(new_n924), .ZN(new_n925));
  XNOR2_X1  g739(.A(new_n925), .B(KEYINPUT124), .ZN(new_n926));
  AND2_X1   g740(.A1(new_n926), .A2(new_n638), .ZN(new_n927));
  XNOR2_X1  g741(.A(new_n553), .B(KEYINPUT125), .ZN(new_n928));
  OAI21_X1  g742(.A(new_n882), .B1(new_n926), .B2(new_n928), .ZN(new_n929));
  NOR2_X1   g743(.A1(new_n927), .A2(new_n929), .ZN(new_n930));
  XNOR2_X1  g744(.A(new_n930), .B(KEYINPUT61), .ZN(G66));
  NAND2_X1  g745(.A1(new_n821), .A2(new_n704), .ZN(new_n932));
  NOR2_X1   g746(.A1(new_n932), .A2(new_n831), .ZN(new_n933));
  INV_X1    g747(.A(new_n933), .ZN(new_n934));
  NAND2_X1  g748(.A1(G224), .A2(G953), .ZN(new_n935));
  OAI22_X1  g749(.A1(new_n934), .A2(G953), .B1(new_n409), .B2(new_n935), .ZN(new_n936));
  OAI21_X1  g750(.A(new_n885), .B1(G898), .B2(new_n295), .ZN(new_n937));
  XOR2_X1   g751(.A(new_n936), .B(new_n937), .Z(G69));
  AND2_X1   g752(.A1(new_n325), .A2(new_n326), .ZN(new_n939));
  XNOR2_X1  g753(.A(new_n487), .B(new_n939), .ZN(new_n940));
  NAND3_X1  g754(.A1(new_n245), .A2(G900), .A3(G953), .ZN(new_n941));
  NAND3_X1  g755(.A1(new_n761), .A2(new_n557), .A3(new_n716), .ZN(new_n942));
  NAND4_X1  g756(.A1(new_n762), .A2(new_n739), .A3(new_n741), .A4(new_n942), .ZN(new_n943));
  NAND2_X1  g757(.A1(new_n815), .A2(new_n722), .ZN(new_n944));
  NOR3_X1   g758(.A1(new_n943), .A2(new_n769), .A3(new_n944), .ZN(new_n945));
  OAI211_X1 g759(.A(new_n940), .B(new_n941), .C1(new_n945), .C2(G953), .ZN(new_n946));
  NOR3_X1   g760(.A1(new_n504), .A2(new_n675), .A3(new_n556), .ZN(new_n947));
  OAI211_X1 g761(.A(new_n744), .B(new_n947), .C1(new_n823), .C2(new_n827), .ZN(new_n948));
  NAND2_X1  g762(.A1(new_n762), .A2(new_n948), .ZN(new_n949));
  NAND3_X1  g763(.A1(new_n815), .A2(new_n680), .A3(new_n722), .ZN(new_n950));
  OAI21_X1  g764(.A(new_n950), .B1(KEYINPUT126), .B2(KEYINPUT62), .ZN(new_n951));
  NAND2_X1  g765(.A1(KEYINPUT126), .A2(KEYINPUT62), .ZN(new_n952));
  AND2_X1   g766(.A1(new_n951), .A2(new_n952), .ZN(new_n953));
  NOR2_X1   g767(.A1(new_n951), .A2(new_n952), .ZN(new_n954));
  OR4_X1    g768(.A1(new_n769), .A2(new_n949), .A3(new_n953), .A4(new_n954), .ZN(new_n955));
  NOR2_X1   g769(.A1(new_n955), .A2(G953), .ZN(new_n956));
  AND3_X1   g770(.A1(G227), .A2(G900), .A3(G953), .ZN(new_n957));
  OR2_X1    g771(.A1(new_n940), .A2(new_n957), .ZN(new_n958));
  OAI21_X1  g772(.A(new_n946), .B1(new_n956), .B2(new_n958), .ZN(G72));
  NAND2_X1  g773(.A1(G472), .A2(G902), .ZN(new_n960));
  XOR2_X1   g774(.A(new_n960), .B(KEYINPUT63), .Z(new_n961));
  INV_X1    g775(.A(new_n961), .ZN(new_n962));
  AOI21_X1  g776(.A(new_n962), .B1(new_n945), .B2(new_n933), .ZN(new_n963));
  NAND2_X1  g777(.A1(new_n492), .A2(new_n423), .ZN(new_n964));
  OAI21_X1  g778(.A(new_n882), .B1(new_n963), .B2(new_n964), .ZN(new_n965));
  OR2_X1    g779(.A1(new_n955), .A2(new_n934), .ZN(new_n966));
  AOI211_X1 g780(.A(new_n423), .B(new_n492), .C1(new_n966), .C2(new_n961), .ZN(new_n967));
  AOI21_X1  g781(.A(new_n962), .B1(new_n457), .B2(new_n488), .ZN(new_n968));
  AOI211_X1 g782(.A(new_n965), .B(new_n967), .C1(new_n844), .C2(new_n968), .ZN(G57));
endmodule


