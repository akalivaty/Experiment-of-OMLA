//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 1 1 0 1 1 1 0 1 0 0 1 0 1 1 1 0 1 1 0 1 1 0 0 0 0 0 1 0 0 0 1 0 0 1 1 0 0 0 0 1 0 0 0 0 0 1 1 0 0 0 0 0 1 1 1 0 0 0 1 1 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:40:10 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n204, new_n205, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n237, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n244, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1231, new_n1232, new_n1233, new_n1234, new_n1235, new_n1236,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1295, new_n1296, new_n1297, new_n1298, new_n1299,
    new_n1300;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(new_n201), .ZN(new_n202));
  NOR3_X1   g0002(.A1(new_n202), .A2(G50), .A3(G77), .ZN(G353));
  NOR2_X1   g0003(.A1(G97), .A2(G107), .ZN(new_n204));
  INV_X1    g0004(.A(new_n204), .ZN(new_n205));
  NAND2_X1  g0005(.A1(new_n205), .A2(G87), .ZN(G355));
  NAND2_X1  g0006(.A1(G1), .A2(G20), .ZN(new_n207));
  XNOR2_X1  g0007(.A(new_n207), .B(KEYINPUT64), .ZN(new_n208));
  AOI22_X1  g0008(.A1(G68), .A2(G238), .B1(G107), .B2(G264), .ZN(new_n209));
  INV_X1    g0009(.A(G50), .ZN(new_n210));
  INV_X1    g0010(.A(G226), .ZN(new_n211));
  INV_X1    g0011(.A(G87), .ZN(new_n212));
  INV_X1    g0012(.A(G250), .ZN(new_n213));
  OAI221_X1 g0013(.A(new_n209), .B1(new_n210), .B2(new_n211), .C1(new_n212), .C2(new_n213), .ZN(new_n214));
  AOI22_X1  g0014(.A1(G77), .A2(G244), .B1(G116), .B2(G270), .ZN(new_n215));
  AOI22_X1  g0015(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n216));
  NAND2_X1  g0016(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  OAI21_X1  g0017(.A(new_n208), .B1(new_n214), .B2(new_n217), .ZN(new_n218));
  XNOR2_X1  g0018(.A(new_n218), .B(KEYINPUT1), .ZN(new_n219));
  NOR2_X1   g0019(.A1(new_n208), .A2(G13), .ZN(new_n220));
  OAI211_X1 g0020(.A(new_n220), .B(G250), .C1(G257), .C2(G264), .ZN(new_n221));
  XOR2_X1   g0021(.A(new_n221), .B(KEYINPUT0), .Z(new_n222));
  NAND2_X1  g0022(.A1(G1), .A2(G13), .ZN(new_n223));
  INV_X1    g0023(.A(G20), .ZN(new_n224));
  NOR2_X1   g0024(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  NAND2_X1  g0025(.A1(new_n202), .A2(G50), .ZN(new_n226));
  INV_X1    g0026(.A(new_n226), .ZN(new_n227));
  AOI211_X1 g0027(.A(new_n219), .B(new_n222), .C1(new_n225), .C2(new_n227), .ZN(G361));
  XNOR2_X1  g0028(.A(G238), .B(G244), .ZN(new_n229));
  XNOR2_X1  g0029(.A(new_n229), .B(G232), .ZN(new_n230));
  XNOR2_X1  g0030(.A(KEYINPUT2), .B(G226), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n230), .B(new_n231), .ZN(new_n232));
  XNOR2_X1  g0032(.A(G250), .B(G257), .ZN(new_n233));
  XNOR2_X1  g0033(.A(G264), .B(G270), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XOR2_X1   g0035(.A(new_n232), .B(new_n235), .Z(G358));
  XNOR2_X1  g0036(.A(G87), .B(G97), .ZN(new_n237));
  XNOR2_X1  g0037(.A(G107), .B(G116), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XNOR2_X1  g0039(.A(G50), .B(G68), .ZN(new_n240));
  XNOR2_X1  g0040(.A(G58), .B(G77), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n239), .B(new_n242), .ZN(G351));
  INV_X1    g0043(.A(KEYINPUT3), .ZN(new_n244));
  NOR2_X1   g0044(.A1(new_n244), .A2(G33), .ZN(new_n245));
  INV_X1    g0045(.A(G33), .ZN(new_n246));
  NOR2_X1   g0046(.A1(new_n246), .A2(KEYINPUT3), .ZN(new_n247));
  OAI21_X1  g0047(.A(KEYINPUT67), .B1(new_n245), .B2(new_n247), .ZN(new_n248));
  NAND2_X1  g0048(.A1(new_n246), .A2(KEYINPUT3), .ZN(new_n249));
  NAND2_X1  g0049(.A1(new_n244), .A2(G33), .ZN(new_n250));
  INV_X1    g0050(.A(KEYINPUT67), .ZN(new_n251));
  NAND3_X1  g0051(.A1(new_n249), .A2(new_n250), .A3(new_n251), .ZN(new_n252));
  NAND4_X1  g0052(.A1(new_n248), .A2(G232), .A3(G1698), .A4(new_n252), .ZN(new_n253));
  INV_X1    g0053(.A(G1698), .ZN(new_n254));
  NAND4_X1  g0054(.A1(new_n248), .A2(G226), .A3(new_n254), .A4(new_n252), .ZN(new_n255));
  NAND2_X1  g0055(.A1(G33), .A2(G97), .ZN(new_n256));
  NAND3_X1  g0056(.A1(new_n253), .A2(new_n255), .A3(new_n256), .ZN(new_n257));
  AND2_X1   g0057(.A1(G1), .A2(G13), .ZN(new_n258));
  INV_X1    g0058(.A(G41), .ZN(new_n259));
  OAI21_X1  g0059(.A(new_n258), .B1(new_n246), .B2(new_n259), .ZN(new_n260));
  INV_X1    g0060(.A(new_n260), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n257), .A2(new_n261), .ZN(new_n262));
  INV_X1    g0062(.A(KEYINPUT13), .ZN(new_n263));
  XNOR2_X1  g0063(.A(KEYINPUT65), .B(G41), .ZN(new_n264));
  INV_X1    g0064(.A(G45), .ZN(new_n265));
  AOI21_X1  g0065(.A(G1), .B1(new_n264), .B2(new_n265), .ZN(new_n266));
  INV_X1    g0066(.A(KEYINPUT66), .ZN(new_n267));
  NAND4_X1  g0067(.A1(new_n266), .A2(new_n267), .A3(G274), .A4(new_n260), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n259), .A2(KEYINPUT65), .ZN(new_n269));
  INV_X1    g0069(.A(KEYINPUT65), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n270), .A2(G41), .ZN(new_n271));
  NAND3_X1  g0071(.A1(new_n269), .A2(new_n271), .A3(new_n265), .ZN(new_n272));
  INV_X1    g0072(.A(G1), .ZN(new_n273));
  NAND4_X1  g0073(.A1(new_n272), .A2(new_n260), .A3(new_n273), .A4(G274), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n274), .A2(KEYINPUT66), .ZN(new_n275));
  OAI21_X1  g0075(.A(new_n273), .B1(G41), .B2(G45), .ZN(new_n276));
  AND2_X1   g0076(.A1(new_n260), .A2(new_n276), .ZN(new_n277));
  AOI22_X1  g0077(.A1(new_n268), .A2(new_n275), .B1(G238), .B2(new_n277), .ZN(new_n278));
  AND3_X1   g0078(.A1(new_n262), .A2(new_n263), .A3(new_n278), .ZN(new_n279));
  AOI21_X1  g0079(.A(new_n263), .B1(new_n262), .B2(new_n278), .ZN(new_n280));
  NOR2_X1   g0080(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  INV_X1    g0081(.A(G169), .ZN(new_n282));
  OAI21_X1  g0082(.A(KEYINPUT14), .B1(new_n281), .B2(new_n282), .ZN(new_n283));
  INV_X1    g0083(.A(KEYINPUT14), .ZN(new_n284));
  OAI211_X1 g0084(.A(new_n284), .B(G169), .C1(new_n279), .C2(new_n280), .ZN(new_n285));
  AOI21_X1  g0085(.A(KEYINPUT72), .B1(new_n281), .B2(G179), .ZN(new_n286));
  INV_X1    g0086(.A(KEYINPUT72), .ZN(new_n287));
  INV_X1    g0087(.A(G179), .ZN(new_n288));
  NOR4_X1   g0088(.A1(new_n279), .A2(new_n280), .A3(new_n287), .A4(new_n288), .ZN(new_n289));
  OAI211_X1 g0089(.A(new_n283), .B(new_n285), .C1(new_n286), .C2(new_n289), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n224), .A2(G33), .ZN(new_n291));
  XOR2_X1   g0091(.A(new_n291), .B(KEYINPUT70), .Z(new_n292));
  NAND2_X1  g0092(.A1(new_n292), .A2(G77), .ZN(new_n293));
  NOR2_X1   g0093(.A1(G20), .A2(G33), .ZN(new_n294));
  INV_X1    g0094(.A(new_n294), .ZN(new_n295));
  OAI221_X1 g0095(.A(new_n293), .B1(new_n224), .B2(G68), .C1(new_n210), .C2(new_n295), .ZN(new_n296));
  NAND3_X1  g0096(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n297), .A2(new_n223), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n296), .A2(new_n298), .ZN(new_n299));
  INV_X1    g0099(.A(KEYINPUT11), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n299), .A2(new_n300), .ZN(new_n301));
  NAND3_X1  g0101(.A1(new_n273), .A2(G13), .A3(G20), .ZN(new_n302));
  INV_X1    g0102(.A(new_n302), .ZN(new_n303));
  INV_X1    g0103(.A(G68), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  OAI21_X1  g0105(.A(KEYINPUT12), .B1(new_n305), .B2(KEYINPUT71), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n305), .A2(KEYINPUT71), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n306), .A2(new_n307), .ZN(new_n308));
  NAND3_X1  g0108(.A1(new_n305), .A2(KEYINPUT71), .A3(KEYINPUT12), .ZN(new_n309));
  AOI21_X1  g0109(.A(new_n298), .B1(new_n273), .B2(G20), .ZN(new_n310));
  AOI22_X1  g0110(.A1(new_n308), .A2(new_n309), .B1(G68), .B2(new_n310), .ZN(new_n311));
  NAND3_X1  g0111(.A1(new_n296), .A2(KEYINPUT11), .A3(new_n298), .ZN(new_n312));
  NAND3_X1  g0112(.A1(new_n301), .A2(new_n311), .A3(new_n312), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n290), .A2(new_n313), .ZN(new_n314));
  INV_X1    g0114(.A(G238), .ZN(new_n315));
  AND3_X1   g0115(.A1(new_n249), .A2(new_n250), .A3(new_n251), .ZN(new_n316));
  AOI21_X1  g0116(.A(new_n251), .B1(new_n249), .B2(new_n250), .ZN(new_n317));
  NOR2_X1   g0117(.A1(new_n316), .A2(new_n317), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n318), .A2(G1698), .ZN(new_n319));
  OR2_X1    g0119(.A1(new_n319), .A2(KEYINPUT68), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n319), .A2(KEYINPUT68), .ZN(new_n321));
  AOI21_X1  g0121(.A(new_n315), .B1(new_n320), .B2(new_n321), .ZN(new_n322));
  NAND3_X1  g0122(.A1(new_n318), .A2(G232), .A3(new_n254), .ZN(new_n323));
  INV_X1    g0123(.A(G107), .ZN(new_n324));
  OAI21_X1  g0124(.A(new_n323), .B1(new_n324), .B2(new_n318), .ZN(new_n325));
  OAI21_X1  g0125(.A(new_n261), .B1(new_n322), .B2(new_n325), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n268), .A2(new_n275), .ZN(new_n327));
  INV_X1    g0127(.A(new_n327), .ZN(new_n328));
  AOI21_X1  g0128(.A(new_n328), .B1(G244), .B2(new_n277), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n326), .A2(new_n329), .ZN(new_n330));
  NOR2_X1   g0130(.A1(new_n330), .A2(G179), .ZN(new_n331));
  NAND2_X1  g0131(.A1(G20), .A2(G77), .ZN(new_n332));
  XNOR2_X1  g0132(.A(KEYINPUT8), .B(G58), .ZN(new_n333));
  XNOR2_X1  g0133(.A(KEYINPUT15), .B(G87), .ZN(new_n334));
  OAI221_X1 g0134(.A(new_n332), .B1(new_n333), .B2(new_n295), .C1(new_n291), .C2(new_n334), .ZN(new_n335));
  AND2_X1   g0135(.A1(new_n335), .A2(new_n298), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n310), .A2(G77), .ZN(new_n337));
  OAI21_X1  g0137(.A(new_n337), .B1(G77), .B2(new_n302), .ZN(new_n338));
  NOR2_X1   g0138(.A1(new_n336), .A2(new_n338), .ZN(new_n339));
  AOI21_X1  g0139(.A(G169), .B1(new_n326), .B2(new_n329), .ZN(new_n340));
  OR3_X1    g0140(.A1(new_n331), .A2(new_n339), .A3(new_n340), .ZN(new_n341));
  AOI21_X1  g0141(.A(new_n313), .B1(G190), .B2(new_n281), .ZN(new_n342));
  OAI21_X1  g0142(.A(G200), .B1(new_n279), .B2(new_n280), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n342), .A2(new_n343), .ZN(new_n344));
  INV_X1    g0144(.A(G200), .ZN(new_n345));
  AOI21_X1  g0145(.A(new_n345), .B1(new_n326), .B2(new_n329), .ZN(new_n346));
  INV_X1    g0146(.A(new_n346), .ZN(new_n347));
  INV_X1    g0147(.A(G190), .ZN(new_n348));
  OAI211_X1 g0148(.A(new_n347), .B(new_n339), .C1(new_n348), .C2(new_n330), .ZN(new_n349));
  AND4_X1   g0149(.A1(new_n314), .A2(new_n341), .A3(new_n344), .A4(new_n349), .ZN(new_n350));
  AND2_X1   g0150(.A1(new_n297), .A2(new_n223), .ZN(new_n351));
  INV_X1    g0151(.A(KEYINPUT7), .ZN(new_n352));
  XNOR2_X1  g0152(.A(KEYINPUT3), .B(G33), .ZN(new_n353));
  OAI21_X1  g0153(.A(new_n352), .B1(new_n353), .B2(G20), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n249), .A2(new_n250), .ZN(new_n355));
  NAND3_X1  g0155(.A1(new_n355), .A2(KEYINPUT7), .A3(new_n224), .ZN(new_n356));
  AOI21_X1  g0156(.A(new_n304), .B1(new_n354), .B2(new_n356), .ZN(new_n357));
  INV_X1    g0157(.A(G58), .ZN(new_n358));
  NOR2_X1   g0158(.A1(new_n358), .A2(new_n304), .ZN(new_n359));
  OAI21_X1  g0159(.A(G20), .B1(new_n359), .B2(new_n201), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n294), .A2(G159), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  OR2_X1    g0162(.A1(new_n357), .A2(new_n362), .ZN(new_n363));
  INV_X1    g0163(.A(KEYINPUT16), .ZN(new_n364));
  OAI21_X1  g0164(.A(KEYINPUT73), .B1(new_n363), .B2(new_n364), .ZN(new_n365));
  NOR4_X1   g0165(.A1(new_n357), .A2(new_n362), .A3(KEYINPUT73), .A4(new_n364), .ZN(new_n366));
  INV_X1    g0166(.A(new_n366), .ZN(new_n367));
  AOI21_X1  g0167(.A(new_n351), .B1(new_n365), .B2(new_n367), .ZN(new_n368));
  INV_X1    g0168(.A(new_n356), .ZN(new_n369));
  OAI21_X1  g0169(.A(new_n224), .B1(new_n316), .B2(new_n317), .ZN(new_n370));
  AOI21_X1  g0170(.A(new_n369), .B1(new_n370), .B2(new_n352), .ZN(new_n371));
  OAI21_X1  g0171(.A(KEYINPUT74), .B1(new_n371), .B2(new_n304), .ZN(new_n372));
  INV_X1    g0172(.A(KEYINPUT74), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n248), .A2(new_n252), .ZN(new_n374));
  AOI21_X1  g0174(.A(KEYINPUT7), .B1(new_n374), .B2(new_n224), .ZN(new_n375));
  OAI211_X1 g0175(.A(new_n373), .B(G68), .C1(new_n375), .C2(new_n369), .ZN(new_n376));
  INV_X1    g0176(.A(new_n362), .ZN(new_n377));
  NAND3_X1  g0177(.A1(new_n372), .A2(new_n376), .A3(new_n377), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n378), .A2(new_n364), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n368), .A2(new_n379), .ZN(new_n380));
  INV_X1    g0180(.A(KEYINPUT69), .ZN(new_n381));
  XNOR2_X1  g0181(.A(new_n333), .B(new_n381), .ZN(new_n382));
  INV_X1    g0182(.A(new_n382), .ZN(new_n383));
  NOR2_X1   g0183(.A1(new_n383), .A2(new_n310), .ZN(new_n384));
  AOI21_X1  g0184(.A(new_n384), .B1(new_n383), .B2(new_n302), .ZN(new_n385));
  INV_X1    g0185(.A(new_n385), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n211), .A2(G1698), .ZN(new_n387));
  OAI21_X1  g0187(.A(new_n387), .B1(G223), .B2(G1698), .ZN(new_n388));
  OAI22_X1  g0188(.A1(new_n388), .A2(new_n355), .B1(new_n246), .B2(new_n212), .ZN(new_n389));
  AOI22_X1  g0189(.A1(new_n261), .A2(new_n389), .B1(new_n277), .B2(G232), .ZN(new_n390));
  AOI21_X1  g0190(.A(G200), .B1(new_n327), .B2(new_n390), .ZN(new_n391));
  AND2_X1   g0191(.A1(new_n327), .A2(new_n390), .ZN(new_n392));
  AOI21_X1  g0192(.A(new_n391), .B1(new_n348), .B2(new_n392), .ZN(new_n393));
  INV_X1    g0193(.A(new_n393), .ZN(new_n394));
  NAND3_X1  g0194(.A1(new_n380), .A2(new_n386), .A3(new_n394), .ZN(new_n395));
  INV_X1    g0195(.A(KEYINPUT17), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n395), .A2(new_n396), .ZN(new_n397));
  AOI21_X1  g0197(.A(new_n385), .B1(new_n368), .B2(new_n379), .ZN(new_n398));
  AND3_X1   g0198(.A1(new_n327), .A2(G179), .A3(new_n390), .ZN(new_n399));
  AOI21_X1  g0199(.A(new_n282), .B1(new_n327), .B2(new_n390), .ZN(new_n400));
  NOR2_X1   g0200(.A1(new_n399), .A2(new_n400), .ZN(new_n401));
  OAI21_X1  g0201(.A(KEYINPUT18), .B1(new_n398), .B2(new_n401), .ZN(new_n402));
  INV_X1    g0202(.A(KEYINPUT18), .ZN(new_n403));
  INV_X1    g0203(.A(new_n401), .ZN(new_n404));
  INV_X1    g0204(.A(KEYINPUT73), .ZN(new_n405));
  NOR2_X1   g0205(.A1(new_n357), .A2(new_n362), .ZN(new_n406));
  AOI21_X1  g0206(.A(new_n405), .B1(new_n406), .B2(KEYINPUT16), .ZN(new_n407));
  OAI21_X1  g0207(.A(new_n298), .B1(new_n407), .B2(new_n366), .ZN(new_n408));
  AOI21_X1  g0208(.A(new_n408), .B1(new_n364), .B2(new_n378), .ZN(new_n409));
  OAI211_X1 g0209(.A(new_n403), .B(new_n404), .C1(new_n409), .C2(new_n385), .ZN(new_n410));
  NAND3_X1  g0210(.A1(new_n398), .A2(KEYINPUT17), .A3(new_n394), .ZN(new_n411));
  NAND4_X1  g0211(.A1(new_n397), .A2(new_n402), .A3(new_n410), .A4(new_n411), .ZN(new_n412));
  INV_X1    g0212(.A(new_n412), .ZN(new_n413));
  INV_X1    g0213(.A(G223), .ZN(new_n414));
  AOI21_X1  g0214(.A(new_n414), .B1(new_n320), .B2(new_n321), .ZN(new_n415));
  NAND3_X1  g0215(.A1(new_n318), .A2(G222), .A3(new_n254), .ZN(new_n416));
  INV_X1    g0216(.A(G77), .ZN(new_n417));
  OAI21_X1  g0217(.A(new_n416), .B1(new_n417), .B2(new_n318), .ZN(new_n418));
  OAI21_X1  g0218(.A(new_n261), .B1(new_n415), .B2(new_n418), .ZN(new_n419));
  AOI21_X1  g0219(.A(new_n328), .B1(G226), .B2(new_n277), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  NOR2_X1   g0221(.A1(new_n421), .A2(G179), .ZN(new_n422));
  OAI21_X1  g0222(.A(G20), .B1(new_n202), .B2(G50), .ZN(new_n423));
  INV_X1    g0223(.A(G150), .ZN(new_n424));
  OAI21_X1  g0224(.A(new_n423), .B1(new_n424), .B2(new_n295), .ZN(new_n425));
  AOI21_X1  g0225(.A(new_n425), .B1(new_n382), .B2(new_n292), .ZN(new_n426));
  NOR2_X1   g0226(.A1(new_n426), .A2(new_n351), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n310), .A2(G50), .ZN(new_n428));
  OAI21_X1  g0228(.A(new_n428), .B1(G50), .B2(new_n302), .ZN(new_n429));
  NOR2_X1   g0229(.A1(new_n427), .A2(new_n429), .ZN(new_n430));
  AOI21_X1  g0230(.A(G169), .B1(new_n419), .B2(new_n420), .ZN(new_n431));
  NOR3_X1   g0231(.A1(new_n422), .A2(new_n430), .A3(new_n431), .ZN(new_n432));
  XNOR2_X1  g0232(.A(new_n430), .B(KEYINPUT9), .ZN(new_n433));
  INV_X1    g0233(.A(new_n433), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n421), .A2(G200), .ZN(new_n435));
  NAND3_X1  g0235(.A1(new_n419), .A2(G190), .A3(new_n420), .ZN(new_n436));
  NAND3_X1  g0236(.A1(new_n434), .A2(new_n435), .A3(new_n436), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n437), .A2(KEYINPUT10), .ZN(new_n438));
  INV_X1    g0238(.A(KEYINPUT10), .ZN(new_n439));
  NAND4_X1  g0239(.A1(new_n435), .A2(new_n434), .A3(new_n439), .A4(new_n436), .ZN(new_n440));
  AOI21_X1  g0240(.A(new_n432), .B1(new_n438), .B2(new_n440), .ZN(new_n441));
  NAND3_X1  g0241(.A1(new_n350), .A2(new_n413), .A3(new_n441), .ZN(new_n442));
  XNOR2_X1  g0242(.A(G97), .B(G107), .ZN(new_n443));
  INV_X1    g0243(.A(KEYINPUT6), .ZN(new_n444));
  AND2_X1   g0244(.A1(new_n443), .A2(new_n444), .ZN(new_n445));
  INV_X1    g0245(.A(G97), .ZN(new_n446));
  NOR3_X1   g0246(.A1(new_n444), .A2(new_n446), .A3(G107), .ZN(new_n447));
  NOR2_X1   g0247(.A1(new_n445), .A2(new_n447), .ZN(new_n448));
  OAI22_X1  g0248(.A1(new_n448), .A2(new_n224), .B1(new_n417), .B2(new_n295), .ZN(new_n449));
  OAI21_X1  g0249(.A(G107), .B1(new_n375), .B2(new_n369), .ZN(new_n450));
  AOI21_X1  g0250(.A(new_n449), .B1(new_n450), .B2(KEYINPUT75), .ZN(new_n451));
  INV_X1    g0251(.A(KEYINPUT75), .ZN(new_n452));
  OAI211_X1 g0252(.A(new_n452), .B(G107), .C1(new_n375), .C2(new_n369), .ZN(new_n453));
  AOI21_X1  g0253(.A(new_n351), .B1(new_n451), .B2(new_n453), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n303), .A2(new_n446), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n273), .A2(G33), .ZN(new_n456));
  NAND3_X1  g0256(.A1(new_n351), .A2(new_n302), .A3(new_n456), .ZN(new_n457));
  OAI21_X1  g0257(.A(new_n455), .B1(new_n457), .B2(new_n446), .ZN(new_n458));
  OAI21_X1  g0258(.A(KEYINPUT76), .B1(new_n454), .B2(new_n458), .ZN(new_n459));
  OAI21_X1  g0259(.A(KEYINPUT75), .B1(new_n371), .B2(new_n324), .ZN(new_n460));
  INV_X1    g0260(.A(new_n449), .ZN(new_n461));
  NAND3_X1  g0261(.A1(new_n460), .A2(new_n461), .A3(new_n453), .ZN(new_n462));
  AOI21_X1  g0262(.A(new_n458), .B1(new_n462), .B2(new_n298), .ZN(new_n463));
  INV_X1    g0263(.A(KEYINPUT76), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n273), .A2(G45), .ZN(new_n466));
  INV_X1    g0266(.A(new_n466), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n259), .A2(KEYINPUT5), .ZN(new_n468));
  OAI211_X1 g0268(.A(new_n467), .B(new_n468), .C1(new_n264), .C2(KEYINPUT5), .ZN(new_n469));
  NAND3_X1  g0269(.A1(new_n469), .A2(G257), .A3(new_n260), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n470), .A2(KEYINPUT80), .ZN(new_n471));
  INV_X1    g0271(.A(KEYINPUT80), .ZN(new_n472));
  NAND4_X1  g0272(.A1(new_n469), .A2(new_n472), .A3(G257), .A4(new_n260), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n471), .A2(new_n473), .ZN(new_n474));
  NAND4_X1  g0274(.A1(new_n248), .A2(G250), .A3(G1698), .A4(new_n252), .ZN(new_n475));
  AND2_X1   g0275(.A1(new_n254), .A2(G244), .ZN(new_n476));
  NAND4_X1  g0276(.A1(new_n248), .A2(KEYINPUT4), .A3(new_n252), .A4(new_n476), .ZN(new_n477));
  NAND4_X1  g0277(.A1(new_n249), .A2(new_n250), .A3(G244), .A4(new_n254), .ZN(new_n478));
  INV_X1    g0278(.A(KEYINPUT4), .ZN(new_n479));
  AOI21_X1  g0279(.A(KEYINPUT77), .B1(G33), .B2(G283), .ZN(new_n480));
  INV_X1    g0280(.A(new_n480), .ZN(new_n481));
  NAND3_X1  g0281(.A1(KEYINPUT77), .A2(G33), .A3(G283), .ZN(new_n482));
  AOI22_X1  g0282(.A1(new_n478), .A2(new_n479), .B1(new_n481), .B2(new_n482), .ZN(new_n483));
  NAND3_X1  g0283(.A1(new_n475), .A2(new_n477), .A3(new_n483), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n484), .A2(new_n261), .ZN(new_n485));
  INV_X1    g0285(.A(KEYINPUT5), .ZN(new_n486));
  OAI21_X1  g0286(.A(KEYINPUT79), .B1(new_n486), .B2(G41), .ZN(new_n487));
  INV_X1    g0287(.A(KEYINPUT79), .ZN(new_n488));
  NAND3_X1  g0288(.A1(new_n488), .A2(new_n259), .A3(KEYINPUT5), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n487), .A2(new_n489), .ZN(new_n490));
  NAND3_X1  g0290(.A1(new_n490), .A2(G274), .A3(new_n260), .ZN(new_n491));
  INV_X1    g0291(.A(new_n491), .ZN(new_n492));
  NOR2_X1   g0292(.A1(new_n270), .A2(G41), .ZN(new_n493));
  NOR2_X1   g0293(.A1(new_n259), .A2(KEYINPUT65), .ZN(new_n494));
  OAI21_X1  g0294(.A(new_n486), .B1(new_n493), .B2(new_n494), .ZN(new_n495));
  AOI21_X1  g0295(.A(KEYINPUT78), .B1(new_n495), .B2(new_n467), .ZN(new_n496));
  AOI21_X1  g0296(.A(KEYINPUT5), .B1(new_n269), .B2(new_n271), .ZN(new_n497));
  INV_X1    g0297(.A(KEYINPUT78), .ZN(new_n498));
  NOR3_X1   g0298(.A1(new_n497), .A2(new_n498), .A3(new_n466), .ZN(new_n499));
  OAI21_X1  g0299(.A(new_n492), .B1(new_n496), .B2(new_n499), .ZN(new_n500));
  NAND3_X1  g0300(.A1(new_n474), .A2(new_n485), .A3(new_n500), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n501), .A2(new_n345), .ZN(new_n502));
  OAI21_X1  g0302(.A(new_n502), .B1(G190), .B2(new_n501), .ZN(new_n503));
  NAND3_X1  g0303(.A1(new_n459), .A2(new_n465), .A3(new_n503), .ZN(new_n504));
  INV_X1    g0304(.A(new_n463), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n501), .A2(G169), .ZN(new_n506));
  OAI21_X1  g0306(.A(new_n498), .B1(new_n497), .B2(new_n466), .ZN(new_n507));
  OAI211_X1 g0307(.A(KEYINPUT78), .B(new_n467), .C1(new_n264), .C2(KEYINPUT5), .ZN(new_n508));
  AOI21_X1  g0308(.A(new_n491), .B1(new_n507), .B2(new_n508), .ZN(new_n509));
  AOI21_X1  g0309(.A(new_n509), .B1(new_n484), .B2(new_n261), .ZN(new_n510));
  NAND3_X1  g0310(.A1(new_n510), .A2(G179), .A3(new_n474), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n506), .A2(new_n511), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n505), .A2(new_n512), .ZN(new_n513));
  NAND3_X1  g0313(.A1(new_n353), .A2(G244), .A3(G1698), .ZN(new_n514));
  NAND3_X1  g0314(.A1(new_n353), .A2(G238), .A3(new_n254), .ZN(new_n515));
  NAND2_X1  g0315(.A1(G33), .A2(G116), .ZN(new_n516));
  NAND3_X1  g0316(.A1(new_n514), .A2(new_n515), .A3(new_n516), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n517), .A2(new_n261), .ZN(new_n518));
  OR2_X1    g0318(.A1(new_n466), .A2(G274), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n466), .A2(new_n213), .ZN(new_n520));
  NAND3_X1  g0320(.A1(new_n519), .A2(new_n260), .A3(new_n520), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n518), .A2(new_n521), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n522), .A2(G200), .ZN(new_n523));
  INV_X1    g0323(.A(KEYINPUT19), .ZN(new_n524));
  OAI21_X1  g0324(.A(new_n224), .B1(new_n256), .B2(new_n524), .ZN(new_n525));
  OAI21_X1  g0325(.A(new_n525), .B1(G87), .B2(new_n205), .ZN(new_n526));
  OAI21_X1  g0326(.A(new_n524), .B1(new_n291), .B2(new_n446), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n353), .A2(new_n224), .ZN(new_n528));
  OAI211_X1 g0328(.A(new_n526), .B(new_n527), .C1(new_n528), .C2(new_n304), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n529), .A2(new_n298), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n334), .A2(new_n303), .ZN(new_n531));
  AND3_X1   g0331(.A1(new_n351), .A2(new_n302), .A3(new_n456), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n532), .A2(G87), .ZN(new_n533));
  AND3_X1   g0333(.A1(new_n530), .A2(new_n531), .A3(new_n533), .ZN(new_n534));
  INV_X1    g0334(.A(new_n521), .ZN(new_n535));
  AOI21_X1  g0335(.A(new_n535), .B1(new_n517), .B2(new_n261), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n536), .A2(G190), .ZN(new_n537));
  NAND3_X1  g0337(.A1(new_n523), .A2(new_n534), .A3(new_n537), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n522), .A2(new_n282), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n536), .A2(new_n288), .ZN(new_n540));
  OR3_X1    g0340(.A1(new_n457), .A2(KEYINPUT81), .A3(new_n334), .ZN(new_n541));
  OAI21_X1  g0341(.A(KEYINPUT81), .B1(new_n457), .B2(new_n334), .ZN(new_n542));
  NAND4_X1  g0342(.A1(new_n530), .A2(new_n541), .A3(new_n531), .A4(new_n542), .ZN(new_n543));
  NAND3_X1  g0343(.A1(new_n539), .A2(new_n540), .A3(new_n543), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n538), .A2(new_n544), .ZN(new_n545));
  INV_X1    g0345(.A(KEYINPUT23), .ZN(new_n546));
  NOR3_X1   g0346(.A1(new_n546), .A2(new_n224), .A3(G107), .ZN(new_n547));
  AOI21_X1  g0347(.A(KEYINPUT23), .B1(new_n324), .B2(G20), .ZN(new_n548));
  OAI22_X1  g0348(.A1(new_n547), .A2(new_n548), .B1(G20), .B2(new_n516), .ZN(new_n549));
  OAI21_X1  g0349(.A(KEYINPUT22), .B1(new_n528), .B2(new_n212), .ZN(new_n550));
  NOR3_X1   g0350(.A1(new_n212), .A2(KEYINPUT22), .A3(G20), .ZN(new_n551));
  NAND3_X1  g0351(.A1(new_n248), .A2(new_n252), .A3(new_n551), .ZN(new_n552));
  AOI21_X1  g0352(.A(new_n549), .B1(new_n550), .B2(new_n552), .ZN(new_n553));
  INV_X1    g0353(.A(KEYINPUT24), .ZN(new_n554));
  NOR2_X1   g0354(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  AOI211_X1 g0355(.A(KEYINPUT24), .B(new_n549), .C1(new_n550), .C2(new_n552), .ZN(new_n556));
  OAI21_X1  g0356(.A(new_n298), .B1(new_n555), .B2(new_n556), .ZN(new_n557));
  NOR2_X1   g0357(.A1(new_n302), .A2(G107), .ZN(new_n558));
  XNOR2_X1  g0358(.A(KEYINPUT84), .B(KEYINPUT25), .ZN(new_n559));
  XNOR2_X1  g0359(.A(new_n558), .B(new_n559), .ZN(new_n560));
  AOI21_X1  g0360(.A(new_n560), .B1(G107), .B2(new_n532), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n557), .A2(new_n561), .ZN(new_n562));
  INV_X1    g0362(.A(new_n562), .ZN(new_n563));
  NAND3_X1  g0363(.A1(new_n469), .A2(G264), .A3(new_n260), .ZN(new_n564));
  NAND3_X1  g0364(.A1(new_n353), .A2(G257), .A3(G1698), .ZN(new_n565));
  NAND3_X1  g0365(.A1(new_n353), .A2(G250), .A3(new_n254), .ZN(new_n566));
  NAND2_X1  g0366(.A1(G33), .A2(G294), .ZN(new_n567));
  NAND3_X1  g0367(.A1(new_n565), .A2(new_n566), .A3(new_n567), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n568), .A2(new_n261), .ZN(new_n569));
  NAND3_X1  g0369(.A1(new_n500), .A2(new_n564), .A3(new_n569), .ZN(new_n570));
  NOR2_X1   g0370(.A1(new_n570), .A2(new_n348), .ZN(new_n571));
  AOI21_X1  g0371(.A(new_n571), .B1(G200), .B2(new_n570), .ZN(new_n572));
  AOI21_X1  g0372(.A(new_n545), .B1(new_n563), .B2(new_n572), .ZN(new_n573));
  NAND3_X1  g0373(.A1(new_n504), .A2(new_n513), .A3(new_n573), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n570), .A2(new_n282), .ZN(new_n575));
  NAND4_X1  g0375(.A1(new_n500), .A2(new_n288), .A3(new_n569), .A4(new_n564), .ZN(new_n576));
  AND2_X1   g0376(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n577), .A2(new_n562), .ZN(new_n578));
  INV_X1    g0378(.A(G303), .ZN(new_n579));
  AOI21_X1  g0379(.A(new_n579), .B1(new_n248), .B2(new_n252), .ZN(new_n580));
  NAND4_X1  g0380(.A1(new_n249), .A2(new_n250), .A3(G264), .A4(G1698), .ZN(new_n581));
  NAND4_X1  g0381(.A1(new_n249), .A2(new_n250), .A3(G257), .A4(new_n254), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  OAI21_X1  g0383(.A(new_n261), .B1(new_n580), .B2(new_n583), .ZN(new_n584));
  NAND3_X1  g0384(.A1(new_n469), .A2(G270), .A3(new_n260), .ZN(new_n585));
  NAND3_X1  g0385(.A1(new_n500), .A2(new_n584), .A3(new_n585), .ZN(new_n586));
  INV_X1    g0386(.A(KEYINPUT20), .ZN(new_n587));
  OAI21_X1  g0387(.A(new_n224), .B1(new_n446), .B2(G33), .ZN(new_n588));
  AOI21_X1  g0388(.A(new_n588), .B1(new_n481), .B2(new_n482), .ZN(new_n589));
  INV_X1    g0389(.A(G116), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n590), .A2(G20), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n298), .A2(new_n591), .ZN(new_n592));
  OAI21_X1  g0392(.A(new_n587), .B1(new_n589), .B2(new_n592), .ZN(new_n593));
  AOI21_X1  g0393(.A(G20), .B1(new_n246), .B2(G97), .ZN(new_n594));
  INV_X1    g0394(.A(new_n482), .ZN(new_n595));
  OAI21_X1  g0395(.A(new_n594), .B1(new_n595), .B2(new_n480), .ZN(new_n596));
  NAND4_X1  g0396(.A1(new_n596), .A2(KEYINPUT20), .A3(new_n298), .A4(new_n591), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n593), .A2(new_n597), .ZN(new_n598));
  NOR2_X1   g0398(.A1(new_n302), .A2(G116), .ZN(new_n599));
  AOI21_X1  g0399(.A(new_n599), .B1(new_n532), .B2(G116), .ZN(new_n600));
  AOI21_X1  g0400(.A(new_n282), .B1(new_n598), .B2(new_n600), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n586), .A2(new_n601), .ZN(new_n602));
  INV_X1    g0402(.A(KEYINPUT21), .ZN(new_n603));
  AND3_X1   g0403(.A1(new_n500), .A2(new_n584), .A3(new_n585), .ZN(new_n604));
  AOI21_X1  g0404(.A(new_n288), .B1(new_n598), .B2(new_n600), .ZN(new_n605));
  AOI22_X1  g0405(.A1(new_n602), .A2(new_n603), .B1(new_n604), .B2(new_n605), .ZN(new_n606));
  NAND4_X1  g0406(.A1(new_n586), .A2(new_n601), .A3(KEYINPUT82), .A4(KEYINPUT21), .ZN(new_n607));
  NAND3_X1  g0407(.A1(new_n586), .A2(new_n601), .A3(KEYINPUT21), .ZN(new_n608));
  INV_X1    g0408(.A(KEYINPUT82), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  AND2_X1   g0410(.A1(new_n598), .A2(new_n600), .ZN(new_n611));
  NAND4_X1  g0411(.A1(new_n500), .A2(new_n584), .A3(G190), .A4(new_n585), .ZN(new_n612));
  OAI211_X1 g0412(.A(new_n611), .B(new_n612), .C1(new_n604), .C2(new_n345), .ZN(new_n613));
  NAND4_X1  g0413(.A1(new_n606), .A2(new_n607), .A3(new_n610), .A4(new_n613), .ZN(new_n614));
  INV_X1    g0414(.A(KEYINPUT83), .ZN(new_n615));
  AND2_X1   g0415(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  NOR2_X1   g0416(.A1(new_n614), .A2(new_n615), .ZN(new_n617));
  OAI21_X1  g0417(.A(new_n578), .B1(new_n616), .B2(new_n617), .ZN(new_n618));
  NOR3_X1   g0418(.A1(new_n442), .A2(new_n574), .A3(new_n618), .ZN(G372));
  NAND2_X1  g0419(.A1(new_n402), .A2(new_n410), .ZN(new_n620));
  INV_X1    g0420(.A(new_n620), .ZN(new_n621));
  NOR3_X1   g0421(.A1(new_n331), .A2(new_n340), .A3(new_n339), .ZN(new_n622));
  AOI22_X1  g0422(.A1(new_n622), .A2(new_n344), .B1(new_n313), .B2(new_n290), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n397), .A2(new_n411), .ZN(new_n624));
  OAI21_X1  g0424(.A(new_n621), .B1(new_n623), .B2(new_n624), .ZN(new_n625));
  OR2_X1    g0425(.A1(new_n625), .A2(KEYINPUT88), .ZN(new_n626));
  AOI22_X1  g0426(.A1(new_n625), .A2(KEYINPUT88), .B1(new_n438), .B2(new_n440), .ZN(new_n627));
  AOI21_X1  g0427(.A(new_n432), .B1(new_n626), .B2(new_n627), .ZN(new_n628));
  AND3_X1   g0428(.A1(new_n504), .A2(new_n513), .A3(new_n573), .ZN(new_n629));
  NAND3_X1  g0429(.A1(new_n606), .A2(new_n607), .A3(new_n610), .ZN(new_n630));
  INV_X1    g0430(.A(KEYINPUT85), .ZN(new_n631));
  XNOR2_X1  g0431(.A(new_n578), .B(new_n631), .ZN(new_n632));
  OAI21_X1  g0432(.A(new_n629), .B1(new_n630), .B2(new_n632), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n459), .A2(new_n465), .ZN(new_n634));
  AND3_X1   g0434(.A1(new_n510), .A2(G179), .A3(new_n474), .ZN(new_n635));
  AOI21_X1  g0435(.A(new_n282), .B1(new_n510), .B2(new_n474), .ZN(new_n636));
  INV_X1    g0436(.A(KEYINPUT86), .ZN(new_n637));
  NOR3_X1   g0437(.A1(new_n635), .A2(new_n636), .A3(new_n637), .ZN(new_n638));
  AOI21_X1  g0438(.A(KEYINPUT86), .B1(new_n506), .B2(new_n511), .ZN(new_n639));
  NOR2_X1   g0439(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  INV_X1    g0440(.A(KEYINPUT26), .ZN(new_n641));
  AND2_X1   g0441(.A1(new_n538), .A2(new_n544), .ZN(new_n642));
  NAND4_X1  g0442(.A1(new_n634), .A2(new_n640), .A3(new_n641), .A4(new_n642), .ZN(new_n643));
  INV_X1    g0443(.A(KEYINPUT87), .ZN(new_n644));
  INV_X1    g0444(.A(new_n544), .ZN(new_n645));
  NAND3_X1  g0445(.A1(new_n505), .A2(new_n642), .A3(new_n512), .ZN(new_n646));
  AOI21_X1  g0446(.A(new_n645), .B1(new_n646), .B2(KEYINPUT26), .ZN(new_n647));
  AND3_X1   g0447(.A1(new_n643), .A2(new_n644), .A3(new_n647), .ZN(new_n648));
  AOI21_X1  g0448(.A(new_n644), .B1(new_n643), .B2(new_n647), .ZN(new_n649));
  OAI21_X1  g0449(.A(new_n633), .B1(new_n648), .B2(new_n649), .ZN(new_n650));
  INV_X1    g0450(.A(new_n650), .ZN(new_n651));
  OAI21_X1  g0451(.A(new_n628), .B1(new_n442), .B2(new_n651), .ZN(G369));
  NAND3_X1  g0452(.A1(new_n273), .A2(new_n224), .A3(G13), .ZN(new_n653));
  OR2_X1    g0453(.A1(new_n653), .A2(KEYINPUT27), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n653), .A2(KEYINPUT27), .ZN(new_n655));
  NAND3_X1  g0455(.A1(new_n654), .A2(G213), .A3(new_n655), .ZN(new_n656));
  INV_X1    g0456(.A(G343), .ZN(new_n657));
  NOR2_X1   g0457(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  INV_X1    g0458(.A(new_n658), .ZN(new_n659));
  NOR2_X1   g0459(.A1(new_n611), .A2(new_n659), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n630), .A2(new_n660), .ZN(new_n661));
  XOR2_X1   g0461(.A(new_n661), .B(KEYINPUT89), .Z(new_n662));
  NOR2_X1   g0462(.A1(new_n616), .A2(new_n617), .ZN(new_n663));
  OAI21_X1  g0463(.A(new_n662), .B1(new_n663), .B2(new_n660), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n563), .A2(new_n572), .ZN(new_n665));
  OAI211_X1 g0465(.A(new_n665), .B(new_n578), .C1(new_n563), .C2(new_n659), .ZN(new_n666));
  INV_X1    g0466(.A(new_n578), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n667), .A2(new_n658), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n666), .A2(new_n668), .ZN(new_n669));
  NAND3_X1  g0469(.A1(new_n664), .A2(G330), .A3(new_n669), .ZN(new_n670));
  XNOR2_X1  g0470(.A(new_n670), .B(KEYINPUT90), .ZN(new_n671));
  INV_X1    g0471(.A(new_n671), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n630), .A2(new_n659), .ZN(new_n673));
  NOR2_X1   g0473(.A1(new_n666), .A2(new_n673), .ZN(new_n674));
  AOI21_X1  g0474(.A(new_n674), .B1(new_n632), .B2(new_n659), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n672), .A2(new_n675), .ZN(G399));
  NAND2_X1  g0476(.A1(new_n220), .A2(new_n264), .ZN(new_n677));
  NOR3_X1   g0477(.A1(new_n205), .A2(G87), .A3(G116), .ZN(new_n678));
  AND3_X1   g0478(.A1(new_n677), .A2(G1), .A3(new_n678), .ZN(new_n679));
  INV_X1    g0479(.A(new_n677), .ZN(new_n680));
  AOI21_X1  g0480(.A(new_n679), .B1(new_n227), .B2(new_n680), .ZN(new_n681));
  XOR2_X1   g0481(.A(new_n681), .B(KEYINPUT28), .Z(new_n682));
  INV_X1    g0482(.A(KEYINPUT29), .ZN(new_n683));
  AND3_X1   g0483(.A1(new_n650), .A2(new_n683), .A3(new_n659), .ZN(new_n684));
  OAI21_X1  g0484(.A(new_n637), .B1(new_n635), .B2(new_n636), .ZN(new_n685));
  NAND3_X1  g0485(.A1(new_n506), .A2(KEYINPUT86), .A3(new_n511), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  AOI21_X1  g0487(.A(new_n687), .B1(new_n459), .B2(new_n465), .ZN(new_n688));
  NAND4_X1  g0488(.A1(new_n688), .A2(KEYINPUT92), .A3(KEYINPUT26), .A4(new_n642), .ZN(new_n689));
  NAND4_X1  g0489(.A1(new_n634), .A2(new_n640), .A3(KEYINPUT26), .A4(new_n642), .ZN(new_n690));
  NOR2_X1   g0490(.A1(new_n635), .A2(new_n636), .ZN(new_n691));
  NOR3_X1   g0491(.A1(new_n691), .A2(new_n463), .A3(new_n545), .ZN(new_n692));
  OAI21_X1  g0492(.A(KEYINPUT92), .B1(new_n692), .B2(KEYINPUT26), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n690), .A2(new_n693), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n689), .A2(new_n694), .ZN(new_n695));
  NAND4_X1  g0495(.A1(new_n578), .A2(new_n607), .A3(new_n610), .A4(new_n606), .ZN(new_n696));
  NAND4_X1  g0496(.A1(new_n504), .A2(new_n573), .A3(new_n696), .A4(new_n513), .ZN(new_n697));
  AND2_X1   g0497(.A1(new_n697), .A2(new_n544), .ZN(new_n698));
  AOI21_X1  g0498(.A(new_n658), .B1(new_n695), .B2(new_n698), .ZN(new_n699));
  NOR2_X1   g0499(.A1(new_n699), .A2(new_n683), .ZN(new_n700));
  NOR2_X1   g0500(.A1(new_n684), .A2(new_n700), .ZN(new_n701));
  INV_X1    g0501(.A(G330), .ZN(new_n702));
  OR2_X1    g0502(.A1(new_n614), .A2(new_n615), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n614), .A2(new_n615), .ZN(new_n704));
  AOI21_X1  g0504(.A(new_n667), .B1(new_n703), .B2(new_n704), .ZN(new_n705));
  NAND3_X1  g0505(.A1(new_n705), .A2(new_n629), .A3(new_n659), .ZN(new_n706));
  INV_X1    g0506(.A(KEYINPUT30), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n569), .A2(new_n564), .ZN(new_n708));
  OAI21_X1  g0508(.A(KEYINPUT91), .B1(new_n522), .B2(new_n708), .ZN(new_n709));
  INV_X1    g0509(.A(KEYINPUT91), .ZN(new_n710));
  NAND4_X1  g0510(.A1(new_n536), .A2(new_n710), .A3(new_n564), .A4(new_n569), .ZN(new_n711));
  AND2_X1   g0511(.A1(new_n709), .A2(new_n711), .ZN(new_n712));
  NAND4_X1  g0512(.A1(new_n604), .A2(G179), .A3(new_n474), .A4(new_n510), .ZN(new_n713));
  OAI21_X1  g0513(.A(new_n707), .B1(new_n712), .B2(new_n713), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n709), .A2(new_n711), .ZN(new_n715));
  NAND4_X1  g0515(.A1(new_n715), .A2(new_n635), .A3(KEYINPUT30), .A4(new_n604), .ZN(new_n716));
  NOR2_X1   g0516(.A1(new_n536), .A2(G179), .ZN(new_n717));
  NAND4_X1  g0517(.A1(new_n501), .A2(new_n570), .A3(new_n586), .A4(new_n717), .ZN(new_n718));
  NAND3_X1  g0518(.A1(new_n714), .A2(new_n716), .A3(new_n718), .ZN(new_n719));
  AND3_X1   g0519(.A1(new_n719), .A2(KEYINPUT31), .A3(new_n658), .ZN(new_n720));
  AOI21_X1  g0520(.A(KEYINPUT31), .B1(new_n719), .B2(new_n658), .ZN(new_n721));
  NOR2_X1   g0521(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  AOI21_X1  g0522(.A(new_n702), .B1(new_n706), .B2(new_n722), .ZN(new_n723));
  INV_X1    g0523(.A(new_n723), .ZN(new_n724));
  NAND2_X1  g0524(.A1(new_n701), .A2(new_n724), .ZN(new_n725));
  INV_X1    g0525(.A(new_n725), .ZN(new_n726));
  OAI21_X1  g0526(.A(new_n682), .B1(new_n726), .B2(G1), .ZN(G364));
  AND2_X1   g0527(.A1(new_n224), .A2(G13), .ZN(new_n728));
  AOI21_X1  g0528(.A(new_n273), .B1(new_n728), .B2(G45), .ZN(new_n729));
  INV_X1    g0529(.A(new_n729), .ZN(new_n730));
  NOR2_X1   g0530(.A1(new_n680), .A2(new_n730), .ZN(new_n731));
  AOI21_X1  g0531(.A(new_n731), .B1(new_n664), .B2(G330), .ZN(new_n732));
  OAI21_X1  g0532(.A(new_n732), .B1(G330), .B2(new_n664), .ZN(new_n733));
  INV_X1    g0533(.A(new_n731), .ZN(new_n734));
  OAI21_X1  g0534(.A(new_n258), .B1(new_n224), .B2(G169), .ZN(new_n735));
  XOR2_X1   g0535(.A(new_n735), .B(KEYINPUT94), .Z(new_n736));
  NOR2_X1   g0536(.A1(new_n224), .A2(new_n288), .ZN(new_n737));
  INV_X1    g0537(.A(new_n737), .ZN(new_n738));
  NOR3_X1   g0538(.A1(new_n738), .A2(new_n345), .A3(G190), .ZN(new_n739));
  INV_X1    g0539(.A(new_n739), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n740), .A2(KEYINPUT95), .ZN(new_n741));
  INV_X1    g0541(.A(new_n741), .ZN(new_n742));
  NOR2_X1   g0542(.A1(new_n740), .A2(KEYINPUT95), .ZN(new_n743));
  NOR2_X1   g0543(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  INV_X1    g0544(.A(new_n744), .ZN(new_n745));
  XNOR2_X1  g0545(.A(KEYINPUT33), .B(G317), .ZN(new_n746));
  NAND2_X1  g0546(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  NOR3_X1   g0547(.A1(new_n738), .A2(new_n348), .A3(G200), .ZN(new_n748));
  INV_X1    g0548(.A(new_n748), .ZN(new_n749));
  INV_X1    g0549(.A(G322), .ZN(new_n750));
  NOR2_X1   g0550(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  NOR3_X1   g0551(.A1(new_n738), .A2(new_n348), .A3(new_n345), .ZN(new_n752));
  INV_X1    g0552(.A(new_n752), .ZN(new_n753));
  INV_X1    g0553(.A(G326), .ZN(new_n754));
  NOR2_X1   g0554(.A1(G190), .A2(G200), .ZN(new_n755));
  NAND2_X1  g0555(.A1(new_n737), .A2(new_n755), .ZN(new_n756));
  INV_X1    g0556(.A(G311), .ZN(new_n757));
  OAI22_X1  g0557(.A1(new_n753), .A2(new_n754), .B1(new_n756), .B2(new_n757), .ZN(new_n758));
  NOR2_X1   g0558(.A1(new_n224), .A2(G179), .ZN(new_n759));
  NAND2_X1  g0559(.A1(new_n759), .A2(new_n755), .ZN(new_n760));
  INV_X1    g0560(.A(new_n760), .ZN(new_n761));
  AOI211_X1 g0561(.A(new_n751), .B(new_n758), .C1(G329), .C2(new_n761), .ZN(new_n762));
  NAND3_X1  g0562(.A1(new_n759), .A2(G190), .A3(G200), .ZN(new_n763));
  INV_X1    g0563(.A(new_n763), .ZN(new_n764));
  AOI21_X1  g0564(.A(new_n318), .B1(G303), .B2(new_n764), .ZN(new_n765));
  NOR3_X1   g0565(.A1(new_n348), .A2(G179), .A3(G200), .ZN(new_n766));
  NOR2_X1   g0566(.A1(new_n766), .A2(new_n224), .ZN(new_n767));
  INV_X1    g0567(.A(new_n767), .ZN(new_n768));
  NAND3_X1  g0568(.A1(new_n759), .A2(new_n348), .A3(G200), .ZN(new_n769));
  INV_X1    g0569(.A(new_n769), .ZN(new_n770));
  AOI22_X1  g0570(.A1(new_n768), .A2(G294), .B1(new_n770), .B2(G283), .ZN(new_n771));
  NAND4_X1  g0571(.A1(new_n747), .A2(new_n762), .A3(new_n765), .A4(new_n771), .ZN(new_n772));
  AOI22_X1  g0572(.A1(new_n748), .A2(G58), .B1(new_n752), .B2(G50), .ZN(new_n773));
  OAI21_X1  g0573(.A(new_n773), .B1(new_n417), .B2(new_n756), .ZN(new_n774));
  INV_X1    g0574(.A(KEYINPUT32), .ZN(new_n775));
  INV_X1    g0575(.A(G159), .ZN(new_n776));
  OAI21_X1  g0576(.A(new_n775), .B1(new_n760), .B2(new_n776), .ZN(new_n777));
  NAND3_X1  g0577(.A1(new_n761), .A2(KEYINPUT32), .A3(G159), .ZN(new_n778));
  AOI21_X1  g0578(.A(new_n774), .B1(new_n777), .B2(new_n778), .ZN(new_n779));
  NAND2_X1  g0579(.A1(new_n764), .A2(G87), .ZN(new_n780));
  OAI21_X1  g0580(.A(new_n780), .B1(new_n324), .B2(new_n769), .ZN(new_n781));
  AOI211_X1 g0581(.A(new_n374), .B(new_n781), .C1(G97), .C2(new_n768), .ZN(new_n782));
  OAI211_X1 g0582(.A(new_n779), .B(new_n782), .C1(new_n304), .C2(new_n744), .ZN(new_n783));
  AOI21_X1  g0583(.A(new_n736), .B1(new_n772), .B2(new_n783), .ZN(new_n784));
  INV_X1    g0584(.A(new_n736), .ZN(new_n785));
  NOR2_X1   g0585(.A1(G13), .A2(G33), .ZN(new_n786));
  INV_X1    g0586(.A(new_n786), .ZN(new_n787));
  NOR2_X1   g0587(.A1(new_n787), .A2(G20), .ZN(new_n788));
  NOR2_X1   g0588(.A1(new_n785), .A2(new_n788), .ZN(new_n789));
  INV_X1    g0589(.A(new_n220), .ZN(new_n790));
  NOR2_X1   g0590(.A1(new_n790), .A2(new_n353), .ZN(new_n791));
  OAI21_X1  g0591(.A(new_n791), .B1(G45), .B2(new_n226), .ZN(new_n792));
  AOI21_X1  g0592(.A(new_n792), .B1(G45), .B2(new_n242), .ZN(new_n793));
  NAND2_X1  g0593(.A1(new_n220), .A2(new_n318), .ZN(new_n794));
  XNOR2_X1  g0594(.A(G355), .B(KEYINPUT93), .ZN(new_n795));
  OAI22_X1  g0595(.A1(new_n794), .A2(new_n795), .B1(G116), .B2(new_n220), .ZN(new_n796));
  OR2_X1    g0596(.A1(new_n793), .A2(new_n796), .ZN(new_n797));
  AOI211_X1 g0597(.A(new_n734), .B(new_n784), .C1(new_n789), .C2(new_n797), .ZN(new_n798));
  INV_X1    g0598(.A(new_n788), .ZN(new_n799));
  OAI21_X1  g0599(.A(new_n798), .B1(new_n664), .B2(new_n799), .ZN(new_n800));
  AND2_X1   g0600(.A1(new_n733), .A2(new_n800), .ZN(new_n801));
  INV_X1    g0601(.A(new_n801), .ZN(G396));
  OAI21_X1  g0602(.A(new_n658), .B1(new_n336), .B2(new_n338), .ZN(new_n803));
  OAI21_X1  g0603(.A(new_n339), .B1(new_n330), .B2(new_n348), .ZN(new_n804));
  OAI21_X1  g0604(.A(new_n803), .B1(new_n804), .B2(new_n346), .ZN(new_n805));
  NAND2_X1  g0605(.A1(new_n341), .A2(new_n805), .ZN(new_n806));
  NAND2_X1  g0606(.A1(new_n622), .A2(new_n659), .ZN(new_n807));
  NAND2_X1  g0607(.A1(new_n806), .A2(new_n807), .ZN(new_n808));
  OAI21_X1  g0608(.A(new_n808), .B1(new_n651), .B2(new_n658), .ZN(new_n809));
  INV_X1    g0609(.A(new_n808), .ZN(new_n810));
  NAND3_X1  g0610(.A1(new_n650), .A2(new_n810), .A3(new_n659), .ZN(new_n811));
  NAND2_X1  g0611(.A1(new_n809), .A2(new_n811), .ZN(new_n812));
  AOI21_X1  g0612(.A(new_n731), .B1(new_n812), .B2(new_n724), .ZN(new_n813));
  OAI21_X1  g0613(.A(new_n813), .B1(new_n724), .B2(new_n812), .ZN(new_n814));
  NAND2_X1  g0614(.A1(new_n808), .A2(new_n786), .ZN(new_n815));
  INV_X1    g0615(.A(new_n756), .ZN(new_n816));
  AOI22_X1  g0616(.A1(new_n752), .A2(G137), .B1(G159), .B2(new_n816), .ZN(new_n817));
  INV_X1    g0617(.A(G143), .ZN(new_n818));
  OAI221_X1 g0618(.A(new_n817), .B1(new_n818), .B2(new_n749), .C1(new_n744), .C2(new_n424), .ZN(new_n819));
  XOR2_X1   g0619(.A(new_n819), .B(KEYINPUT34), .Z(new_n820));
  INV_X1    g0620(.A(G132), .ZN(new_n821));
  OAI221_X1 g0621(.A(new_n353), .B1(new_n760), .B2(new_n821), .C1(new_n767), .C2(new_n358), .ZN(new_n822));
  NOR2_X1   g0622(.A1(new_n763), .A2(new_n210), .ZN(new_n823));
  NOR2_X1   g0623(.A1(new_n769), .A2(new_n304), .ZN(new_n824));
  NOR4_X1   g0624(.A1(new_n820), .A2(new_n822), .A3(new_n823), .A4(new_n824), .ZN(new_n825));
  INV_X1    g0625(.A(G283), .ZN(new_n826));
  NOR2_X1   g0626(.A1(new_n744), .A2(new_n826), .ZN(new_n827));
  NOR2_X1   g0627(.A1(new_n769), .A2(new_n212), .ZN(new_n828));
  AOI21_X1  g0628(.A(new_n828), .B1(G107), .B2(new_n764), .ZN(new_n829));
  OAI211_X1 g0629(.A(new_n829), .B(new_n374), .C1(new_n446), .C2(new_n767), .ZN(new_n830));
  OAI22_X1  g0630(.A1(new_n753), .A2(new_n579), .B1(new_n760), .B2(new_n757), .ZN(new_n831));
  INV_X1    g0631(.A(G294), .ZN(new_n832));
  OAI22_X1  g0632(.A1(new_n749), .A2(new_n832), .B1(new_n756), .B2(new_n590), .ZN(new_n833));
  NOR4_X1   g0633(.A1(new_n827), .A2(new_n830), .A3(new_n831), .A4(new_n833), .ZN(new_n834));
  OAI21_X1  g0634(.A(new_n785), .B1(new_n825), .B2(new_n834), .ZN(new_n835));
  NAND2_X1  g0635(.A1(new_n736), .A2(new_n787), .ZN(new_n836));
  XOR2_X1   g0636(.A(new_n836), .B(KEYINPUT96), .Z(new_n837));
  XNOR2_X1  g0637(.A(new_n837), .B(KEYINPUT97), .ZN(new_n838));
  OR2_X1    g0638(.A1(new_n838), .A2(G77), .ZN(new_n839));
  NAND4_X1  g0639(.A1(new_n815), .A2(new_n731), .A3(new_n835), .A4(new_n839), .ZN(new_n840));
  NAND2_X1  g0640(.A1(new_n814), .A2(new_n840), .ZN(G384));
  INV_X1    g0641(.A(new_n448), .ZN(new_n842));
  OR2_X1    g0642(.A1(new_n842), .A2(KEYINPUT35), .ZN(new_n843));
  NAND2_X1  g0643(.A1(new_n842), .A2(KEYINPUT35), .ZN(new_n844));
  NAND4_X1  g0644(.A1(new_n843), .A2(G116), .A3(new_n225), .A4(new_n844), .ZN(new_n845));
  XOR2_X1   g0645(.A(new_n845), .B(KEYINPUT36), .Z(new_n846));
  OR3_X1    g0646(.A1(new_n226), .A2(new_n417), .A3(new_n359), .ZN(new_n847));
  NAND2_X1  g0647(.A1(new_n210), .A2(G68), .ZN(new_n848));
  AOI211_X1 g0648(.A(new_n273), .B(G13), .C1(new_n847), .C2(new_n848), .ZN(new_n849));
  NOR2_X1   g0649(.A1(new_n846), .A2(new_n849), .ZN(new_n850));
  NAND2_X1  g0650(.A1(new_n314), .A2(KEYINPUT98), .ZN(new_n851));
  INV_X1    g0651(.A(KEYINPUT98), .ZN(new_n852));
  NAND3_X1  g0652(.A1(new_n290), .A2(new_n852), .A3(new_n313), .ZN(new_n853));
  NAND2_X1  g0653(.A1(new_n851), .A2(new_n853), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n854), .A2(new_n659), .ZN(new_n855));
  INV_X1    g0655(.A(new_n855), .ZN(new_n856));
  INV_X1    g0656(.A(KEYINPUT99), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n363), .A2(new_n364), .ZN(new_n858));
  OAI211_X1 g0658(.A(new_n298), .B(new_n858), .C1(new_n407), .C2(new_n366), .ZN(new_n859));
  AOI22_X1  g0659(.A1(new_n859), .A2(new_n386), .B1(new_n401), .B2(new_n656), .ZN(new_n860));
  AOI21_X1  g0660(.A(new_n860), .B1(new_n398), .B2(new_n394), .ZN(new_n861));
  INV_X1    g0661(.A(KEYINPUT37), .ZN(new_n862));
  OAI21_X1  g0662(.A(new_n857), .B1(new_n861), .B2(new_n862), .ZN(new_n863));
  OAI21_X1  g0663(.A(new_n404), .B1(new_n409), .B2(new_n385), .ZN(new_n864));
  INV_X1    g0664(.A(new_n656), .ZN(new_n865));
  OAI21_X1  g0665(.A(new_n865), .B1(new_n409), .B2(new_n385), .ZN(new_n866));
  NAND4_X1  g0666(.A1(new_n864), .A2(new_n866), .A3(new_n862), .A4(new_n395), .ZN(new_n867));
  AOI211_X1 g0667(.A(new_n385), .B(new_n393), .C1(new_n368), .C2(new_n379), .ZN(new_n868));
  OAI211_X1 g0668(.A(KEYINPUT99), .B(KEYINPUT37), .C1(new_n868), .C2(new_n860), .ZN(new_n869));
  NAND3_X1  g0669(.A1(new_n863), .A2(new_n867), .A3(new_n869), .ZN(new_n870));
  AOI21_X1  g0670(.A(new_n656), .B1(new_n859), .B2(new_n386), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n412), .A2(new_n871), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n870), .A2(new_n872), .ZN(new_n873));
  INV_X1    g0673(.A(KEYINPUT38), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  NAND3_X1  g0675(.A1(new_n870), .A2(new_n872), .A3(KEYINPUT38), .ZN(new_n876));
  NAND3_X1  g0676(.A1(new_n875), .A2(KEYINPUT39), .A3(new_n876), .ZN(new_n877));
  INV_X1    g0677(.A(KEYINPUT101), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n876), .A2(new_n878), .ZN(new_n879));
  NAND4_X1  g0679(.A1(new_n870), .A2(new_n872), .A3(KEYINPUT101), .A4(KEYINPUT38), .ZN(new_n880));
  NOR2_X1   g0680(.A1(new_n398), .A2(new_n401), .ZN(new_n881));
  NOR2_X1   g0681(.A1(new_n881), .A2(new_n868), .ZN(new_n882));
  NAND4_X1  g0682(.A1(new_n882), .A2(KEYINPUT100), .A3(new_n862), .A4(new_n866), .ZN(new_n883));
  INV_X1    g0683(.A(KEYINPUT100), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n867), .A2(new_n884), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n864), .A2(new_n395), .ZN(new_n886));
  INV_X1    g0686(.A(new_n866), .ZN(new_n887));
  OAI21_X1  g0687(.A(KEYINPUT37), .B1(new_n886), .B2(new_n887), .ZN(new_n888));
  NAND3_X1  g0688(.A1(new_n883), .A2(new_n885), .A3(new_n888), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n412), .A2(new_n887), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  AOI22_X1  g0691(.A1(new_n879), .A2(new_n880), .B1(new_n891), .B2(new_n874), .ZN(new_n892));
  OAI211_X1 g0692(.A(new_n856), .B(new_n877), .C1(new_n892), .C2(KEYINPUT39), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n313), .A2(new_n658), .ZN(new_n894));
  NAND4_X1  g0694(.A1(new_n851), .A2(new_n344), .A3(new_n853), .A4(new_n894), .ZN(new_n895));
  INV_X1    g0695(.A(new_n344), .ZN(new_n896));
  OAI211_X1 g0696(.A(new_n313), .B(new_n658), .C1(new_n896), .C2(new_n290), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n895), .A2(new_n897), .ZN(new_n898));
  INV_X1    g0698(.A(new_n898), .ZN(new_n899));
  AOI21_X1  g0699(.A(new_n899), .B1(new_n811), .B2(new_n807), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n875), .A2(new_n876), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n620), .A2(new_n656), .ZN(new_n903));
  NAND3_X1  g0703(.A1(new_n893), .A2(new_n902), .A3(new_n903), .ZN(new_n904));
  INV_X1    g0704(.A(new_n442), .ZN(new_n905));
  OAI21_X1  g0705(.A(new_n905), .B1(new_n684), .B2(new_n700), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n906), .A2(new_n628), .ZN(new_n907));
  XOR2_X1   g0707(.A(new_n904), .B(new_n907), .Z(new_n908));
  AOI21_X1  g0708(.A(new_n808), .B1(new_n895), .B2(new_n897), .ZN(new_n909));
  NOR3_X1   g0709(.A1(new_n618), .A2(new_n574), .A3(new_n658), .ZN(new_n910));
  INV_X1    g0710(.A(new_n721), .ZN(new_n911));
  NAND3_X1  g0711(.A1(new_n719), .A2(KEYINPUT31), .A3(new_n658), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  OAI21_X1  g0713(.A(KEYINPUT102), .B1(new_n910), .B2(new_n913), .ZN(new_n914));
  INV_X1    g0714(.A(KEYINPUT102), .ZN(new_n915));
  NAND3_X1  g0715(.A1(new_n706), .A2(new_n722), .A3(new_n915), .ZN(new_n916));
  NAND3_X1  g0716(.A1(new_n909), .A2(new_n914), .A3(new_n916), .ZN(new_n917));
  OAI21_X1  g0717(.A(KEYINPUT40), .B1(new_n892), .B2(new_n917), .ZN(new_n918));
  AND2_X1   g0718(.A1(new_n914), .A2(new_n916), .ZN(new_n919));
  INV_X1    g0719(.A(KEYINPUT40), .ZN(new_n920));
  NAND4_X1  g0720(.A1(new_n919), .A2(new_n901), .A3(new_n920), .A4(new_n909), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n918), .A2(new_n921), .ZN(new_n922));
  AND2_X1   g0722(.A1(new_n919), .A2(new_n905), .ZN(new_n923));
  AND2_X1   g0723(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  NOR2_X1   g0724(.A1(new_n922), .A2(new_n923), .ZN(new_n925));
  NOR3_X1   g0725(.A1(new_n924), .A2(new_n925), .A3(new_n702), .ZN(new_n926));
  OAI22_X1  g0726(.A1(new_n908), .A2(new_n926), .B1(new_n273), .B2(new_n728), .ZN(new_n927));
  AND2_X1   g0727(.A1(new_n908), .A2(new_n926), .ZN(new_n928));
  OAI21_X1  g0728(.A(new_n850), .B1(new_n927), .B2(new_n928), .ZN(G367));
  NAND2_X1  g0729(.A1(new_n634), .A2(new_n658), .ZN(new_n930));
  NAND3_X1  g0730(.A1(new_n930), .A2(new_n513), .A3(new_n504), .ZN(new_n931));
  INV_X1    g0731(.A(KEYINPUT103), .ZN(new_n932));
  XNOR2_X1  g0732(.A(new_n931), .B(new_n932), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n688), .A2(new_n658), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n933), .A2(new_n934), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n935), .A2(new_n674), .ZN(new_n936));
  INV_X1    g0736(.A(KEYINPUT42), .ZN(new_n937));
  XNOR2_X1  g0737(.A(new_n936), .B(new_n937), .ZN(new_n938));
  INV_X1    g0738(.A(new_n935), .ZN(new_n939));
  OAI21_X1  g0739(.A(new_n513), .B1(new_n939), .B2(new_n578), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n940), .A2(new_n659), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n938), .A2(new_n941), .ZN(new_n942));
  OR2_X1    g0742(.A1(new_n534), .A2(new_n659), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n642), .A2(new_n943), .ZN(new_n944));
  OR2_X1    g0744(.A1(new_n943), .A2(new_n544), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n944), .A2(new_n945), .ZN(new_n946));
  OR3_X1    g0746(.A1(new_n942), .A2(KEYINPUT43), .A3(new_n946), .ZN(new_n947));
  AOI22_X1  g0747(.A1(new_n938), .A2(new_n941), .B1(KEYINPUT43), .B2(new_n946), .ZN(new_n948));
  OAI21_X1  g0748(.A(new_n948), .B1(KEYINPUT43), .B2(new_n946), .ZN(new_n949));
  NAND4_X1  g0749(.A1(new_n947), .A2(new_n949), .A3(new_n671), .A4(new_n935), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n947), .A2(new_n949), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n671), .A2(new_n935), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n951), .A2(new_n952), .ZN(new_n953));
  XNOR2_X1  g0753(.A(new_n677), .B(KEYINPUT41), .ZN(new_n954));
  NOR2_X1   g0754(.A1(new_n935), .A2(new_n675), .ZN(new_n955));
  XNOR2_X1  g0755(.A(new_n955), .B(KEYINPUT44), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n935), .A2(new_n675), .ZN(new_n957));
  INV_X1    g0757(.A(KEYINPUT45), .ZN(new_n958));
  XNOR2_X1  g0758(.A(new_n957), .B(new_n958), .ZN(new_n959));
  AOI21_X1  g0759(.A(new_n672), .B1(new_n956), .B2(new_n959), .ZN(new_n960));
  INV_X1    g0760(.A(new_n960), .ZN(new_n961));
  INV_X1    g0761(.A(new_n669), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n962), .A2(new_n673), .ZN(new_n963));
  INV_X1    g0763(.A(new_n674), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n963), .A2(new_n964), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n664), .A2(G330), .ZN(new_n966));
  AOI21_X1  g0766(.A(new_n965), .B1(new_n966), .B2(KEYINPUT104), .ZN(new_n967));
  INV_X1    g0767(.A(KEYINPUT104), .ZN(new_n968));
  NAND3_X1  g0768(.A1(new_n664), .A2(new_n968), .A3(G330), .ZN(new_n969));
  OR2_X1    g0769(.A1(new_n967), .A2(new_n969), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n967), .A2(new_n969), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n970), .A2(new_n971), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n726), .A2(new_n972), .ZN(new_n973));
  INV_X1    g0773(.A(new_n973), .ZN(new_n974));
  NAND3_X1  g0774(.A1(new_n956), .A2(new_n672), .A3(new_n959), .ZN(new_n975));
  NAND3_X1  g0775(.A1(new_n961), .A2(new_n974), .A3(new_n975), .ZN(new_n976));
  AOI21_X1  g0776(.A(new_n954), .B1(new_n976), .B2(new_n726), .ZN(new_n977));
  OAI211_X1 g0777(.A(new_n950), .B(new_n953), .C1(new_n977), .C2(new_n730), .ZN(new_n978));
  INV_X1    g0778(.A(new_n789), .ZN(new_n979));
  INV_X1    g0779(.A(new_n334), .ZN(new_n980));
  AOI21_X1  g0780(.A(new_n979), .B1(new_n790), .B2(new_n980), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n791), .A2(new_n235), .ZN(new_n982));
  AOI21_X1  g0782(.A(new_n734), .B1(new_n981), .B2(new_n982), .ZN(new_n983));
  NOR2_X1   g0783(.A1(new_n744), .A2(new_n776), .ZN(new_n984));
  AOI21_X1  g0784(.A(new_n374), .B1(G77), .B2(new_n770), .ZN(new_n985));
  XNOR2_X1  g0785(.A(new_n985), .B(KEYINPUT106), .ZN(new_n986));
  AOI22_X1  g0786(.A1(G50), .A2(new_n816), .B1(new_n761), .B2(G137), .ZN(new_n987));
  OAI221_X1 g0787(.A(new_n987), .B1(new_n749), .B2(new_n424), .C1(new_n818), .C2(new_n753), .ZN(new_n988));
  OAI22_X1  g0788(.A1(new_n767), .A2(new_n304), .B1(new_n763), .B2(new_n358), .ZN(new_n989));
  NOR4_X1   g0789(.A1(new_n984), .A2(new_n986), .A3(new_n988), .A4(new_n989), .ZN(new_n990));
  XNOR2_X1  g0790(.A(new_n990), .B(KEYINPUT107), .ZN(new_n991));
  AND3_X1   g0791(.A1(new_n764), .A2(KEYINPUT46), .A3(G116), .ZN(new_n992));
  AOI21_X1  g0792(.A(KEYINPUT46), .B1(new_n764), .B2(G116), .ZN(new_n993));
  AOI211_X1 g0793(.A(new_n992), .B(new_n993), .C1(new_n745), .C2(G294), .ZN(new_n994));
  AOI21_X1  g0794(.A(new_n353), .B1(new_n761), .B2(G317), .ZN(new_n995));
  OAI21_X1  g0795(.A(new_n995), .B1(new_n446), .B2(new_n769), .ZN(new_n996));
  OR2_X1    g0796(.A1(new_n996), .A2(KEYINPUT105), .ZN(new_n997));
  NAND2_X1  g0797(.A1(new_n996), .A2(KEYINPUT105), .ZN(new_n998));
  NOR2_X1   g0798(.A1(new_n756), .A2(new_n826), .ZN(new_n999));
  OAI22_X1  g0799(.A1(new_n749), .A2(new_n579), .B1(new_n753), .B2(new_n757), .ZN(new_n1000));
  AOI211_X1 g0800(.A(new_n999), .B(new_n1000), .C1(G107), .C2(new_n768), .ZN(new_n1001));
  NAND4_X1  g0801(.A1(new_n994), .A2(new_n997), .A3(new_n998), .A4(new_n1001), .ZN(new_n1002));
  NAND3_X1  g0802(.A1(new_n991), .A2(KEYINPUT47), .A3(new_n1002), .ZN(new_n1003));
  NAND2_X1  g0803(.A1(new_n1003), .A2(new_n785), .ZN(new_n1004));
  AOI21_X1  g0804(.A(KEYINPUT47), .B1(new_n991), .B2(new_n1002), .ZN(new_n1005));
  OAI221_X1 g0805(.A(new_n983), .B1(new_n799), .B2(new_n946), .C1(new_n1004), .C2(new_n1005), .ZN(new_n1006));
  NAND2_X1  g0806(.A1(new_n978), .A2(new_n1006), .ZN(G387));
  OAI21_X1  g0807(.A(new_n791), .B1(new_n232), .B2(new_n265), .ZN(new_n1008));
  OAI21_X1  g0808(.A(new_n1008), .B1(new_n678), .B2(new_n794), .ZN(new_n1009));
  OR3_X1    g0809(.A1(new_n333), .A2(KEYINPUT50), .A3(G50), .ZN(new_n1010));
  OAI21_X1  g0810(.A(KEYINPUT50), .B1(new_n333), .B2(G50), .ZN(new_n1011));
  AOI21_X1  g0811(.A(G45), .B1(G68), .B2(G77), .ZN(new_n1012));
  NAND4_X1  g0812(.A1(new_n1010), .A2(new_n678), .A3(new_n1011), .A4(new_n1012), .ZN(new_n1013));
  AOI22_X1  g0813(.A1(new_n1009), .A2(new_n1013), .B1(new_n324), .B2(new_n790), .ZN(new_n1014));
  OAI21_X1  g0814(.A(new_n731), .B1(new_n1014), .B2(new_n979), .ZN(new_n1015));
  AOI22_X1  g0815(.A1(new_n748), .A2(G317), .B1(new_n752), .B2(G322), .ZN(new_n1016));
  OAI221_X1 g0816(.A(new_n1016), .B1(new_n579), .B2(new_n756), .C1(new_n744), .C2(new_n757), .ZN(new_n1017));
  INV_X1    g0817(.A(KEYINPUT48), .ZN(new_n1018));
  OR2_X1    g0818(.A1(new_n1017), .A2(new_n1018), .ZN(new_n1019));
  NAND2_X1  g0819(.A1(new_n1017), .A2(new_n1018), .ZN(new_n1020));
  AOI22_X1  g0820(.A1(new_n768), .A2(G283), .B1(new_n764), .B2(G294), .ZN(new_n1021));
  NAND3_X1  g0821(.A1(new_n1019), .A2(new_n1020), .A3(new_n1021), .ZN(new_n1022));
  INV_X1    g0822(.A(KEYINPUT49), .ZN(new_n1023));
  AND2_X1   g0823(.A1(new_n1022), .A2(new_n1023), .ZN(new_n1024));
  NOR2_X1   g0824(.A1(new_n1022), .A2(new_n1023), .ZN(new_n1025));
  OAI221_X1 g0825(.A(new_n355), .B1(new_n760), .B2(new_n754), .C1(new_n590), .C2(new_n769), .ZN(new_n1026));
  OR3_X1    g0826(.A1(new_n1024), .A2(new_n1025), .A3(new_n1026), .ZN(new_n1027));
  NAND2_X1  g0827(.A1(new_n745), .A2(new_n382), .ZN(new_n1028));
  XOR2_X1   g0828(.A(KEYINPUT108), .B(G150), .Z(new_n1029));
  AOI21_X1  g0829(.A(new_n355), .B1(new_n761), .B2(new_n1029), .ZN(new_n1030));
  OAI221_X1 g0830(.A(new_n1030), .B1(new_n417), .B2(new_n763), .C1(new_n446), .C2(new_n769), .ZN(new_n1031));
  XNOR2_X1  g0831(.A(new_n1031), .B(KEYINPUT109), .ZN(new_n1032));
  NAND2_X1  g0832(.A1(new_n768), .A2(new_n980), .ZN(new_n1033));
  OAI22_X1  g0833(.A1(new_n749), .A2(new_n210), .B1(new_n756), .B2(new_n304), .ZN(new_n1034));
  AOI21_X1  g0834(.A(new_n1034), .B1(G159), .B2(new_n752), .ZN(new_n1035));
  NAND4_X1  g0835(.A1(new_n1028), .A2(new_n1032), .A3(new_n1033), .A4(new_n1035), .ZN(new_n1036));
  AOI21_X1  g0836(.A(new_n736), .B1(new_n1027), .B2(new_n1036), .ZN(new_n1037));
  AOI211_X1 g0837(.A(new_n1015), .B(new_n1037), .C1(new_n962), .C2(new_n788), .ZN(new_n1038));
  AOI21_X1  g0838(.A(new_n1038), .B1(new_n972), .B2(new_n730), .ZN(new_n1039));
  NAND2_X1  g0839(.A1(new_n973), .A2(new_n680), .ZN(new_n1040));
  NOR2_X1   g0840(.A1(new_n726), .A2(new_n972), .ZN(new_n1041));
  OAI21_X1  g0841(.A(new_n1039), .B1(new_n1040), .B2(new_n1041), .ZN(G393));
  INV_X1    g0842(.A(new_n975), .ZN(new_n1043));
  NOR3_X1   g0843(.A1(new_n1043), .A2(new_n960), .A3(new_n729), .ZN(new_n1044));
  NAND2_X1  g0844(.A1(new_n939), .A2(new_n788), .ZN(new_n1045));
  AOI21_X1  g0845(.A(new_n979), .B1(G97), .B2(new_n790), .ZN(new_n1046));
  NAND2_X1  g0846(.A1(new_n791), .A2(new_n239), .ZN(new_n1047));
  AOI21_X1  g0847(.A(new_n734), .B1(new_n1046), .B2(new_n1047), .ZN(new_n1048));
  XNOR2_X1  g0848(.A(new_n1048), .B(KEYINPUT110), .ZN(new_n1049));
  OAI221_X1 g0849(.A(new_n353), .B1(new_n760), .B2(new_n818), .C1(new_n333), .C2(new_n756), .ZN(new_n1050));
  AOI21_X1  g0850(.A(new_n1050), .B1(new_n745), .B2(G50), .ZN(new_n1051));
  AOI22_X1  g0851(.A1(new_n748), .A2(G159), .B1(new_n752), .B2(G150), .ZN(new_n1052));
  XOR2_X1   g0852(.A(new_n1052), .B(KEYINPUT51), .Z(new_n1053));
  NOR2_X1   g0853(.A1(new_n763), .A2(new_n304), .ZN(new_n1054));
  AOI211_X1 g0854(.A(new_n828), .B(new_n1054), .C1(G77), .C2(new_n768), .ZN(new_n1055));
  NAND3_X1  g0855(.A1(new_n1051), .A2(new_n1053), .A3(new_n1055), .ZN(new_n1056));
  AOI22_X1  g0856(.A1(new_n748), .A2(G311), .B1(new_n752), .B2(G317), .ZN(new_n1057));
  XNOR2_X1  g0857(.A(new_n1057), .B(KEYINPUT52), .ZN(new_n1058));
  OAI22_X1  g0858(.A1(new_n324), .A2(new_n769), .B1(new_n763), .B2(new_n826), .ZN(new_n1059));
  AOI21_X1  g0859(.A(new_n1059), .B1(G116), .B2(new_n768), .ZN(new_n1060));
  OAI22_X1  g0860(.A1(new_n756), .A2(new_n832), .B1(new_n760), .B2(new_n750), .ZN(new_n1061));
  NOR2_X1   g0861(.A1(new_n318), .A2(new_n1061), .ZN(new_n1062));
  OAI211_X1 g0862(.A(new_n1060), .B(new_n1062), .C1(new_n744), .C2(new_n579), .ZN(new_n1063));
  OAI21_X1  g0863(.A(new_n1056), .B1(new_n1058), .B2(new_n1063), .ZN(new_n1064));
  AOI21_X1  g0864(.A(new_n1049), .B1(new_n785), .B2(new_n1064), .ZN(new_n1065));
  AOI21_X1  g0865(.A(new_n1044), .B1(new_n1045), .B2(new_n1065), .ZN(new_n1066));
  OAI21_X1  g0866(.A(new_n973), .B1(new_n1043), .B2(new_n960), .ZN(new_n1067));
  NAND3_X1  g0867(.A1(new_n1067), .A2(new_n976), .A3(new_n680), .ZN(new_n1068));
  NAND2_X1  g0868(.A1(new_n1066), .A2(new_n1068), .ZN(G390));
  NAND4_X1  g0869(.A1(new_n905), .A2(G330), .A3(new_n914), .A4(new_n916), .ZN(new_n1070));
  NAND3_X1  g0870(.A1(new_n906), .A2(new_n628), .A3(new_n1070), .ZN(new_n1071));
  NAND2_X1  g0871(.A1(new_n811), .A2(new_n807), .ZN(new_n1072));
  NAND4_X1  g0872(.A1(new_n909), .A2(G330), .A3(new_n914), .A4(new_n916), .ZN(new_n1073));
  INV_X1    g0873(.A(new_n1073), .ZN(new_n1074));
  AOI21_X1  g0874(.A(new_n898), .B1(new_n723), .B2(new_n810), .ZN(new_n1075));
  OAI21_X1  g0875(.A(new_n1072), .B1(new_n1074), .B2(new_n1075), .ZN(new_n1076));
  NAND4_X1  g0876(.A1(new_n914), .A2(G330), .A3(new_n810), .A4(new_n916), .ZN(new_n1077));
  NAND2_X1  g0877(.A1(new_n1077), .A2(new_n899), .ZN(new_n1078));
  NAND3_X1  g0878(.A1(new_n898), .A2(new_n723), .A3(new_n810), .ZN(new_n1079));
  INV_X1    g0879(.A(KEYINPUT112), .ZN(new_n1080));
  INV_X1    g0880(.A(new_n807), .ZN(new_n1081));
  AOI211_X1 g0881(.A(new_n1080), .B(new_n1081), .C1(new_n699), .C2(new_n806), .ZN(new_n1082));
  NAND2_X1  g0882(.A1(new_n695), .A2(new_n698), .ZN(new_n1083));
  NAND3_X1  g0883(.A1(new_n1083), .A2(new_n659), .A3(new_n806), .ZN(new_n1084));
  AOI21_X1  g0884(.A(KEYINPUT112), .B1(new_n1084), .B2(new_n807), .ZN(new_n1085));
  OAI211_X1 g0885(.A(new_n1078), .B(new_n1079), .C1(new_n1082), .C2(new_n1085), .ZN(new_n1086));
  AOI21_X1  g0886(.A(new_n1071), .B1(new_n1076), .B2(new_n1086), .ZN(new_n1087));
  AOI21_X1  g0887(.A(new_n622), .B1(new_n349), .B2(new_n803), .ZN(new_n1088));
  AOI211_X1 g0888(.A(new_n658), .B(new_n1088), .C1(new_n695), .C2(new_n698), .ZN(new_n1089));
  OAI21_X1  g0889(.A(new_n1080), .B1(new_n1089), .B2(new_n1081), .ZN(new_n1090));
  NAND3_X1  g0890(.A1(new_n1084), .A2(KEYINPUT112), .A3(new_n807), .ZN(new_n1091));
  NAND3_X1  g0891(.A1(new_n1090), .A2(new_n898), .A3(new_n1091), .ZN(new_n1092));
  NAND2_X1  g0892(.A1(new_n891), .A2(new_n874), .ZN(new_n1093));
  NAND2_X1  g0893(.A1(new_n879), .A2(new_n880), .ZN(new_n1094));
  OR2_X1    g0894(.A1(new_n855), .A2(KEYINPUT111), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n855), .A2(KEYINPUT111), .ZN(new_n1096));
  AOI22_X1  g0896(.A1(new_n1093), .A2(new_n1094), .B1(new_n1095), .B2(new_n1096), .ZN(new_n1097));
  NAND2_X1  g0897(.A1(new_n1092), .A2(new_n1097), .ZN(new_n1098));
  AOI21_X1  g0898(.A(KEYINPUT39), .B1(new_n1094), .B2(new_n1093), .ZN(new_n1099));
  INV_X1    g0899(.A(new_n877), .ZN(new_n1100));
  OAI22_X1  g0900(.A1(new_n1099), .A2(new_n1100), .B1(new_n900), .B2(new_n856), .ZN(new_n1101));
  NAND3_X1  g0901(.A1(new_n1098), .A2(new_n1101), .A3(new_n1079), .ZN(new_n1102));
  OAI21_X1  g0902(.A(new_n877), .B1(new_n892), .B2(KEYINPUT39), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n1072), .A2(new_n898), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n1104), .A2(new_n855), .ZN(new_n1105));
  AOI22_X1  g0905(.A1(new_n1103), .A2(new_n1105), .B1(new_n1092), .B2(new_n1097), .ZN(new_n1106));
  OAI211_X1 g0906(.A(new_n1087), .B(new_n1102), .C1(new_n1106), .C2(new_n1073), .ZN(new_n1107));
  INV_X1    g0907(.A(KEYINPUT113), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n1107), .A2(new_n1108), .ZN(new_n1109));
  NAND2_X1  g0909(.A1(new_n1098), .A2(new_n1101), .ZN(new_n1110));
  NAND2_X1  g0910(.A1(new_n1110), .A2(new_n1074), .ZN(new_n1111));
  NAND4_X1  g0911(.A1(new_n1111), .A2(KEYINPUT113), .A3(new_n1102), .A4(new_n1087), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n1109), .A2(new_n1112), .ZN(new_n1113));
  AND2_X1   g0913(.A1(new_n1111), .A2(new_n1102), .ZN(new_n1114));
  OAI211_X1 g0914(.A(new_n1113), .B(new_n680), .C1(new_n1114), .C2(new_n1087), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n1103), .A2(new_n786), .ZN(new_n1116));
  OAI21_X1  g0916(.A(new_n731), .B1(new_n838), .B2(new_n382), .ZN(new_n1117));
  AOI22_X1  g0917(.A1(new_n748), .A2(G116), .B1(G97), .B2(new_n816), .ZN(new_n1118));
  OAI221_X1 g0918(.A(new_n1118), .B1(new_n826), .B2(new_n753), .C1(new_n832), .C2(new_n760), .ZN(new_n1119));
  AOI21_X1  g0919(.A(new_n1119), .B1(new_n745), .B2(G107), .ZN(new_n1120));
  AOI21_X1  g0920(.A(new_n824), .B1(G77), .B2(new_n768), .ZN(new_n1121));
  NAND4_X1  g0921(.A1(new_n1120), .A2(new_n374), .A3(new_n780), .A4(new_n1121), .ZN(new_n1122));
  XNOR2_X1  g0922(.A(new_n1122), .B(KEYINPUT115), .ZN(new_n1123));
  INV_X1    g0923(.A(KEYINPUT53), .ZN(new_n1124));
  AND3_X1   g0924(.A1(new_n764), .A2(new_n1124), .A3(new_n1029), .ZN(new_n1125));
  AOI21_X1  g0925(.A(new_n1124), .B1(new_n764), .B2(new_n1029), .ZN(new_n1126));
  AOI211_X1 g0926(.A(new_n1125), .B(new_n1126), .C1(new_n745), .C2(G137), .ZN(new_n1127));
  OAI21_X1  g0927(.A(new_n318), .B1(new_n210), .B2(new_n769), .ZN(new_n1128));
  INV_X1    g0928(.A(KEYINPUT114), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n1128), .A2(new_n1129), .ZN(new_n1130));
  OR2_X1    g0930(.A1(new_n1128), .A2(new_n1129), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n761), .A2(G125), .ZN(new_n1132));
  OAI21_X1  g0932(.A(new_n1132), .B1(new_n749), .B2(new_n821), .ZN(new_n1133));
  INV_X1    g0933(.A(G128), .ZN(new_n1134));
  XNOR2_X1  g0934(.A(KEYINPUT54), .B(G143), .ZN(new_n1135));
  OAI22_X1  g0935(.A1(new_n753), .A2(new_n1134), .B1(new_n756), .B2(new_n1135), .ZN(new_n1136));
  AOI211_X1 g0936(.A(new_n1133), .B(new_n1136), .C1(G159), .C2(new_n768), .ZN(new_n1137));
  AND4_X1   g0937(.A1(new_n1127), .A2(new_n1130), .A3(new_n1131), .A4(new_n1137), .ZN(new_n1138));
  NOR2_X1   g0938(.A1(new_n1123), .A2(new_n1138), .ZN(new_n1139));
  INV_X1    g0939(.A(KEYINPUT116), .ZN(new_n1140));
  AOI21_X1  g0940(.A(new_n736), .B1(new_n1139), .B2(new_n1140), .ZN(new_n1141));
  OAI21_X1  g0941(.A(KEYINPUT116), .B1(new_n1123), .B2(new_n1138), .ZN(new_n1142));
  AOI21_X1  g0942(.A(new_n1117), .B1(new_n1141), .B2(new_n1142), .ZN(new_n1143));
  AOI22_X1  g0943(.A1(new_n1114), .A2(new_n730), .B1(new_n1116), .B2(new_n1143), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n1115), .A2(new_n1144), .ZN(G378));
  INV_X1    g0945(.A(KEYINPUT119), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n922), .A2(G330), .ZN(new_n1147));
  NOR2_X1   g0947(.A1(new_n430), .A2(new_n656), .ZN(new_n1148));
  AND2_X1   g0948(.A1(new_n438), .A2(new_n440), .ZN(new_n1149));
  OAI21_X1  g0949(.A(new_n1148), .B1(new_n1149), .B2(new_n432), .ZN(new_n1150));
  OAI21_X1  g0950(.A(new_n441), .B1(new_n430), .B2(new_n656), .ZN(new_n1151));
  XNOR2_X1  g0951(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1152));
  AND3_X1   g0952(.A1(new_n1150), .A2(new_n1151), .A3(new_n1152), .ZN(new_n1153));
  AOI21_X1  g0953(.A(new_n1152), .B1(new_n1150), .B2(new_n1151), .ZN(new_n1154));
  NOR2_X1   g0954(.A1(new_n1153), .A2(new_n1154), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n1147), .A2(new_n1155), .ZN(new_n1156));
  INV_X1    g0956(.A(new_n904), .ZN(new_n1157));
  INV_X1    g0957(.A(new_n1155), .ZN(new_n1158));
  NAND3_X1  g0958(.A1(new_n922), .A2(G330), .A3(new_n1158), .ZN(new_n1159));
  NAND3_X1  g0959(.A1(new_n1156), .A2(new_n1157), .A3(new_n1159), .ZN(new_n1160));
  AOI21_X1  g0960(.A(new_n1158), .B1(new_n922), .B2(G330), .ZN(new_n1161));
  AOI211_X1 g0961(.A(new_n702), .B(new_n1155), .C1(new_n918), .C2(new_n921), .ZN(new_n1162));
  OAI21_X1  g0962(.A(new_n904), .B1(new_n1161), .B2(new_n1162), .ZN(new_n1163));
  AND2_X1   g0963(.A1(new_n1160), .A2(new_n1163), .ZN(new_n1164));
  INV_X1    g0964(.A(new_n1071), .ZN(new_n1165));
  AOI21_X1  g0965(.A(new_n1164), .B1(new_n1113), .B2(new_n1165), .ZN(new_n1166));
  OAI21_X1  g0966(.A(new_n1146), .B1(new_n1166), .B2(KEYINPUT57), .ZN(new_n1167));
  AOI21_X1  g0967(.A(new_n677), .B1(new_n1166), .B2(KEYINPUT57), .ZN(new_n1168));
  INV_X1    g0968(.A(KEYINPUT57), .ZN(new_n1169));
  AOI21_X1  g0969(.A(new_n1071), .B1(new_n1109), .B2(new_n1112), .ZN(new_n1170));
  OAI211_X1 g0970(.A(KEYINPUT119), .B(new_n1169), .C1(new_n1170), .C2(new_n1164), .ZN(new_n1171));
  NAND3_X1  g0971(.A1(new_n1167), .A2(new_n1168), .A3(new_n1171), .ZN(new_n1172));
  NAND2_X1  g0972(.A1(new_n1160), .A2(new_n1163), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n1155), .A2(new_n786), .ZN(new_n1174));
  AOI22_X1  g0974(.A1(new_n748), .A2(G107), .B1(G283), .B2(new_n761), .ZN(new_n1175));
  OAI221_X1 g0975(.A(new_n1175), .B1(new_n334), .B2(new_n756), .C1(new_n744), .C2(new_n446), .ZN(new_n1176));
  NOR2_X1   g0976(.A1(new_n767), .A2(new_n304), .ZN(new_n1177));
  OAI211_X1 g0977(.A(new_n355), .B(new_n264), .C1(new_n753), .C2(new_n590), .ZN(new_n1178));
  OAI22_X1  g0978(.A1(new_n358), .A2(new_n769), .B1(new_n763), .B2(new_n417), .ZN(new_n1179));
  NOR4_X1   g0979(.A1(new_n1176), .A2(new_n1177), .A3(new_n1178), .A4(new_n1179), .ZN(new_n1180));
  OR2_X1    g0980(.A1(new_n1180), .A2(KEYINPUT58), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n1180), .A2(KEYINPUT58), .ZN(new_n1182));
  NOR2_X1   g0982(.A1(G33), .A2(G41), .ZN(new_n1183));
  XNOR2_X1  g0983(.A(new_n1183), .B(KEYINPUT117), .ZN(new_n1184));
  NAND2_X1  g0984(.A1(new_n355), .A2(new_n264), .ZN(new_n1185));
  NAND3_X1  g0985(.A1(new_n1184), .A2(new_n1185), .A3(new_n210), .ZN(new_n1186));
  NAND3_X1  g0986(.A1(new_n1181), .A2(new_n1182), .A3(new_n1186), .ZN(new_n1187));
  AOI22_X1  g0987(.A1(new_n748), .A2(G128), .B1(new_n752), .B2(G125), .ZN(new_n1188));
  INV_X1    g0988(.A(new_n1135), .ZN(new_n1189));
  AOI22_X1  g0989(.A1(new_n768), .A2(G150), .B1(new_n764), .B2(new_n1189), .ZN(new_n1190));
  INV_X1    g0990(.A(G137), .ZN(new_n1191));
  OAI211_X1 g0991(.A(new_n1188), .B(new_n1190), .C1(new_n1191), .C2(new_n756), .ZN(new_n1192));
  AOI21_X1  g0992(.A(new_n1192), .B1(new_n745), .B2(G132), .ZN(new_n1193));
  INV_X1    g0993(.A(new_n1193), .ZN(new_n1194));
  AND2_X1   g0994(.A1(new_n1194), .A2(KEYINPUT59), .ZN(new_n1195));
  NOR2_X1   g0995(.A1(new_n1194), .A2(KEYINPUT59), .ZN(new_n1196));
  AOI21_X1  g0996(.A(new_n1184), .B1(G124), .B2(new_n761), .ZN(new_n1197));
  OAI21_X1  g0997(.A(new_n1197), .B1(new_n776), .B2(new_n769), .ZN(new_n1198));
  NOR3_X1   g0998(.A1(new_n1195), .A2(new_n1196), .A3(new_n1198), .ZN(new_n1199));
  OAI21_X1  g0999(.A(new_n785), .B1(new_n1187), .B2(new_n1199), .ZN(new_n1200));
  XOR2_X1   g1000(.A(new_n1200), .B(KEYINPUT118), .Z(new_n1201));
  AOI211_X1 g1001(.A(new_n734), .B(new_n1201), .C1(new_n210), .C2(new_n837), .ZN(new_n1202));
  AOI22_X1  g1002(.A1(new_n1173), .A2(new_n730), .B1(new_n1174), .B2(new_n1202), .ZN(new_n1203));
  NAND2_X1  g1003(.A1(new_n1172), .A2(new_n1203), .ZN(G375));
  NAND3_X1  g1004(.A1(new_n1086), .A2(new_n1076), .A3(new_n1071), .ZN(new_n1205));
  INV_X1    g1005(.A(new_n1205), .ZN(new_n1206));
  OR3_X1    g1006(.A1(new_n1206), .A2(new_n954), .A3(new_n1087), .ZN(new_n1207));
  OAI22_X1  g1007(.A1(new_n744), .A2(new_n590), .B1(new_n324), .B2(new_n756), .ZN(new_n1208));
  AOI22_X1  g1008(.A1(new_n1208), .A2(KEYINPUT120), .B1(G294), .B2(new_n752), .ZN(new_n1209));
  OAI21_X1  g1009(.A(new_n1209), .B1(KEYINPUT120), .B2(new_n1208), .ZN(new_n1210));
  XOR2_X1   g1010(.A(new_n1210), .B(KEYINPUT121), .Z(new_n1211));
  OAI221_X1 g1011(.A(new_n374), .B1(new_n579), .B2(new_n760), .C1(new_n749), .C2(new_n826), .ZN(new_n1212));
  NOR2_X1   g1012(.A1(new_n763), .A2(new_n446), .ZN(new_n1213));
  OAI21_X1  g1013(.A(new_n1033), .B1(new_n417), .B2(new_n769), .ZN(new_n1214));
  NOR4_X1   g1014(.A1(new_n1211), .A2(new_n1212), .A3(new_n1213), .A4(new_n1214), .ZN(new_n1215));
  OAI22_X1  g1015(.A1(new_n749), .A2(new_n1191), .B1(new_n753), .B2(new_n821), .ZN(new_n1216));
  AOI21_X1  g1016(.A(new_n1216), .B1(new_n745), .B2(new_n1189), .ZN(new_n1217));
  OR2_X1    g1017(.A1(new_n1217), .A2(KEYINPUT122), .ZN(new_n1218));
  NAND2_X1  g1018(.A1(new_n1217), .A2(KEYINPUT122), .ZN(new_n1219));
  OAI22_X1  g1019(.A1(new_n358), .A2(new_n769), .B1(new_n763), .B2(new_n776), .ZN(new_n1220));
  OAI221_X1 g1020(.A(new_n353), .B1(new_n760), .B2(new_n1134), .C1(new_n424), .C2(new_n756), .ZN(new_n1221));
  AOI211_X1 g1021(.A(new_n1220), .B(new_n1221), .C1(G50), .C2(new_n768), .ZN(new_n1222));
  AND3_X1   g1022(.A1(new_n1218), .A2(new_n1219), .A3(new_n1222), .ZN(new_n1223));
  OAI21_X1  g1023(.A(new_n785), .B1(new_n1215), .B2(new_n1223), .ZN(new_n1224));
  OAI211_X1 g1024(.A(new_n1224), .B(new_n731), .C1(G68), .C2(new_n838), .ZN(new_n1225));
  AOI21_X1  g1025(.A(new_n1225), .B1(new_n899), .B2(new_n786), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n1086), .A2(new_n1076), .ZN(new_n1227));
  AOI21_X1  g1027(.A(new_n1226), .B1(new_n1227), .B2(new_n730), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(new_n1207), .A2(new_n1228), .ZN(new_n1229));
  XOR2_X1   g1029(.A(new_n1229), .B(KEYINPUT123), .Z(G381));
  INV_X1    g1030(.A(G390), .ZN(new_n1231));
  INV_X1    g1031(.A(G384), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(new_n1231), .A2(new_n1232), .ZN(new_n1233));
  OR4_X1    g1033(.A1(G396), .A2(new_n1233), .A3(G387), .A4(G393), .ZN(new_n1234));
  INV_X1    g1034(.A(G378), .ZN(new_n1235));
  NAND3_X1  g1035(.A1(new_n1172), .A2(new_n1235), .A3(new_n1203), .ZN(new_n1236));
  OR3_X1    g1036(.A1(new_n1234), .A2(new_n1236), .A3(G381), .ZN(G407));
  OAI211_X1 g1037(.A(G407), .B(G213), .C1(G343), .C2(new_n1236), .ZN(G409));
  XNOR2_X1  g1038(.A(G393), .B(new_n801), .ZN(new_n1239));
  INV_X1    g1039(.A(new_n1239), .ZN(new_n1240));
  NAND3_X1  g1040(.A1(new_n978), .A2(new_n1006), .A3(G390), .ZN(new_n1241));
  INV_X1    g1041(.A(new_n1241), .ZN(new_n1242));
  AOI21_X1  g1042(.A(G390), .B1(new_n978), .B2(new_n1006), .ZN(new_n1243));
  OAI21_X1  g1043(.A(new_n1240), .B1(new_n1242), .B2(new_n1243), .ZN(new_n1244));
  NAND2_X1  g1044(.A1(G387), .A2(new_n1231), .ZN(new_n1245));
  NAND3_X1  g1045(.A1(new_n1245), .A2(new_n1239), .A3(new_n1241), .ZN(new_n1246));
  AND3_X1   g1046(.A1(new_n1244), .A2(KEYINPUT127), .A3(new_n1246), .ZN(new_n1247));
  AOI21_X1  g1047(.A(KEYINPUT127), .B1(new_n1244), .B2(new_n1246), .ZN(new_n1248));
  NOR2_X1   g1048(.A1(new_n1247), .A2(new_n1248), .ZN(new_n1249));
  INV_X1    g1049(.A(new_n1249), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(G375), .A2(G378), .ZN(new_n1251));
  INV_X1    g1051(.A(KEYINPUT62), .ZN(new_n1252));
  AND3_X1   g1052(.A1(new_n1115), .A2(new_n1144), .A3(new_n1203), .ZN(new_n1253));
  INV_X1    g1053(.A(new_n954), .ZN(new_n1254));
  NAND2_X1  g1054(.A1(new_n1166), .A2(new_n1254), .ZN(new_n1255));
  AOI22_X1  g1055(.A1(new_n1253), .A2(new_n1255), .B1(G213), .B2(new_n657), .ZN(new_n1256));
  NOR2_X1   g1056(.A1(new_n1232), .A2(KEYINPUT125), .ZN(new_n1257));
  INV_X1    g1057(.A(KEYINPUT60), .ZN(new_n1258));
  OAI21_X1  g1058(.A(new_n1205), .B1(new_n1087), .B2(new_n1258), .ZN(new_n1259));
  INV_X1    g1059(.A(KEYINPUT124), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(new_n1259), .A2(new_n1260), .ZN(new_n1261));
  OAI211_X1 g1061(.A(KEYINPUT124), .B(new_n1205), .C1(new_n1087), .C2(new_n1258), .ZN(new_n1262));
  AOI21_X1  g1062(.A(new_n677), .B1(new_n1206), .B2(KEYINPUT60), .ZN(new_n1263));
  NAND3_X1  g1063(.A1(new_n1261), .A2(new_n1262), .A3(new_n1263), .ZN(new_n1264));
  AOI21_X1  g1064(.A(new_n1257), .B1(new_n1264), .B2(new_n1228), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(new_n1232), .A2(KEYINPUT125), .ZN(new_n1266));
  NOR2_X1   g1066(.A1(new_n1265), .A2(new_n1266), .ZN(new_n1267));
  INV_X1    g1067(.A(new_n1267), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1265), .A2(new_n1266), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n1268), .A2(new_n1269), .ZN(new_n1270));
  NAND4_X1  g1070(.A1(new_n1251), .A2(new_n1252), .A3(new_n1256), .A4(new_n1270), .ZN(new_n1271));
  INV_X1    g1071(.A(KEYINPUT61), .ZN(new_n1272));
  NAND3_X1  g1072(.A1(new_n657), .A2(G213), .A3(G2897), .ZN(new_n1273));
  INV_X1    g1073(.A(new_n1273), .ZN(new_n1274));
  INV_X1    g1074(.A(new_n1269), .ZN(new_n1275));
  OAI21_X1  g1075(.A(new_n1274), .B1(new_n1275), .B2(new_n1267), .ZN(new_n1276));
  NAND3_X1  g1076(.A1(new_n1268), .A2(new_n1269), .A3(new_n1273), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(new_n1276), .A2(new_n1277), .ZN(new_n1278));
  AOI21_X1  g1078(.A(new_n1235), .B1(new_n1172), .B2(new_n1203), .ZN(new_n1279));
  INV_X1    g1079(.A(new_n1256), .ZN(new_n1280));
  OAI21_X1  g1080(.A(new_n1278), .B1(new_n1279), .B2(new_n1280), .ZN(new_n1281));
  NAND3_X1  g1081(.A1(new_n1271), .A2(new_n1272), .A3(new_n1281), .ZN(new_n1282));
  NOR2_X1   g1082(.A1(new_n1279), .A2(new_n1280), .ZN(new_n1283));
  AOI21_X1  g1083(.A(new_n1252), .B1(new_n1283), .B2(new_n1270), .ZN(new_n1284));
  OAI21_X1  g1084(.A(new_n1250), .B1(new_n1282), .B2(new_n1284), .ZN(new_n1285));
  NAND3_X1  g1085(.A1(new_n1244), .A2(new_n1246), .A3(new_n1272), .ZN(new_n1286));
  INV_X1    g1086(.A(KEYINPUT126), .ZN(new_n1287));
  XNOR2_X1  g1087(.A(new_n1286), .B(new_n1287), .ZN(new_n1288));
  NAND3_X1  g1088(.A1(new_n1251), .A2(new_n1256), .A3(new_n1270), .ZN(new_n1289));
  INV_X1    g1089(.A(KEYINPUT63), .ZN(new_n1290));
  NAND2_X1  g1090(.A1(new_n1289), .A2(new_n1290), .ZN(new_n1291));
  NAND3_X1  g1091(.A1(new_n1283), .A2(KEYINPUT63), .A3(new_n1270), .ZN(new_n1292));
  NAND4_X1  g1092(.A1(new_n1288), .A2(new_n1291), .A3(new_n1292), .A4(new_n1281), .ZN(new_n1293));
  NAND2_X1  g1093(.A1(new_n1285), .A2(new_n1293), .ZN(G405));
  NOR2_X1   g1094(.A1(G375), .A2(G378), .ZN(new_n1295));
  OAI211_X1 g1095(.A(new_n1268), .B(new_n1269), .C1(new_n1295), .C2(new_n1279), .ZN(new_n1296));
  NAND3_X1  g1096(.A1(new_n1251), .A2(new_n1236), .A3(new_n1270), .ZN(new_n1297));
  NAND2_X1  g1097(.A1(new_n1296), .A2(new_n1297), .ZN(new_n1298));
  NAND2_X1  g1098(.A1(new_n1298), .A2(new_n1250), .ZN(new_n1299));
  NAND3_X1  g1099(.A1(new_n1296), .A2(new_n1249), .A3(new_n1297), .ZN(new_n1300));
  NAND2_X1  g1100(.A1(new_n1299), .A2(new_n1300), .ZN(G402));
endmodule


