//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 0 1 1 1 1 1 1 1 1 1 1 1 0 0 1 0 1 1 0 0 1 1 0 1 1 0 0 0 0 1 0 0 0 0 0 0 0 0 0 1 0 1 0 1 0 1 1 0 1 1 1 1 1 1 1 1 0 1 0 0 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:26:44 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n694, new_n695, new_n696,
    new_n697, new_n698, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n712,
    new_n713, new_n715, new_n716, new_n717, new_n719, new_n720, new_n721,
    new_n722, new_n723, new_n724, new_n725, new_n726, new_n727, new_n728,
    new_n729, new_n730, new_n731, new_n733, new_n734, new_n735, new_n736,
    new_n737, new_n738, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n755, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n783, new_n784, new_n785, new_n786, new_n787, new_n788, new_n789,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n926, new_n927, new_n928, new_n929, new_n930, new_n931,
    new_n932, new_n933, new_n934, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n944, new_n945, new_n946, new_n947,
    new_n949, new_n950, new_n951, new_n952, new_n953, new_n954, new_n955,
    new_n956, new_n957, new_n958, new_n959, new_n960, new_n962, new_n963,
    new_n964, new_n965, new_n966, new_n967, new_n968, new_n969, new_n970,
    new_n971, new_n972, new_n973, new_n974, new_n975, new_n976, new_n977,
    new_n978, new_n980, new_n981, new_n982, new_n983, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1021, new_n1022, new_n1023, new_n1024, new_n1025,
    new_n1026;
  INV_X1    g000(.A(G119), .ZN(new_n187));
  NAND2_X1  g001(.A1(new_n187), .A2(G116), .ZN(new_n188));
  INV_X1    g002(.A(G116), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n189), .A2(G119), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n188), .A2(new_n190), .ZN(new_n191));
  XNOR2_X1  g005(.A(KEYINPUT2), .B(G113), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n191), .A2(new_n192), .ZN(new_n193));
  INV_X1    g007(.A(KEYINPUT2), .ZN(new_n194));
  INV_X1    g008(.A(G113), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n194), .A2(new_n195), .ZN(new_n196));
  NAND2_X1  g010(.A1(KEYINPUT2), .A2(G113), .ZN(new_n197));
  NAND4_X1  g011(.A1(new_n196), .A2(new_n188), .A3(new_n190), .A4(new_n197), .ZN(new_n198));
  AND3_X1   g012(.A1(new_n193), .A2(KEYINPUT69), .A3(new_n198), .ZN(new_n199));
  AOI21_X1  g013(.A(KEYINPUT69), .B1(new_n193), .B2(new_n198), .ZN(new_n200));
  NOR2_X1   g014(.A1(new_n199), .A2(new_n200), .ZN(new_n201));
  INV_X1    g015(.A(KEYINPUT1), .ZN(new_n202));
  INV_X1    g016(.A(G146), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n203), .A2(G143), .ZN(new_n204));
  INV_X1    g018(.A(G143), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n205), .A2(G146), .ZN(new_n206));
  AND4_X1   g020(.A1(new_n202), .A2(new_n204), .A3(new_n206), .A4(G128), .ZN(new_n207));
  OAI21_X1  g021(.A(KEYINPUT1), .B1(new_n205), .B2(G146), .ZN(new_n208));
  INV_X1    g022(.A(KEYINPUT68), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  NAND3_X1  g024(.A1(new_n204), .A2(KEYINPUT68), .A3(KEYINPUT1), .ZN(new_n211));
  NAND3_X1  g025(.A1(new_n210), .A2(G128), .A3(new_n211), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n204), .A2(new_n206), .ZN(new_n213));
  AOI21_X1  g027(.A(new_n207), .B1(new_n212), .B2(new_n213), .ZN(new_n214));
  INV_X1    g028(.A(KEYINPUT67), .ZN(new_n215));
  INV_X1    g029(.A(G137), .ZN(new_n216));
  OAI21_X1  g030(.A(new_n215), .B1(new_n216), .B2(G134), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n216), .A2(G134), .ZN(new_n218));
  INV_X1    g032(.A(G134), .ZN(new_n219));
  NAND3_X1  g033(.A1(new_n219), .A2(KEYINPUT67), .A3(G137), .ZN(new_n220));
  NAND3_X1  g034(.A1(new_n217), .A2(new_n218), .A3(new_n220), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n221), .A2(G131), .ZN(new_n222));
  INV_X1    g036(.A(KEYINPUT11), .ZN(new_n223));
  OAI22_X1  g037(.A1(KEYINPUT65), .A2(new_n223), .B1(new_n219), .B2(G137), .ZN(new_n224));
  INV_X1    g038(.A(KEYINPUT65), .ZN(new_n225));
  NAND4_X1  g039(.A1(new_n225), .A2(new_n216), .A3(KEYINPUT11), .A4(G134), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n223), .A2(KEYINPUT65), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n219), .A2(G137), .ZN(new_n228));
  NAND4_X1  g042(.A1(new_n224), .A2(new_n226), .A3(new_n227), .A4(new_n228), .ZN(new_n229));
  AND2_X1   g043(.A1(KEYINPUT66), .A2(G131), .ZN(new_n230));
  NOR2_X1   g044(.A1(KEYINPUT66), .A2(G131), .ZN(new_n231));
  NOR2_X1   g045(.A1(new_n230), .A2(new_n231), .ZN(new_n232));
  OAI21_X1  g046(.A(new_n222), .B1(new_n229), .B2(new_n232), .ZN(new_n233));
  NOR2_X1   g047(.A1(new_n214), .A2(new_n233), .ZN(new_n234));
  NOR2_X1   g048(.A1(new_n216), .A2(G134), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n225), .A2(KEYINPUT11), .ZN(new_n236));
  AOI21_X1  g050(.A(new_n235), .B1(new_n218), .B2(new_n236), .ZN(new_n237));
  INV_X1    g051(.A(new_n232), .ZN(new_n238));
  NAND4_X1  g052(.A1(new_n237), .A2(new_n238), .A3(new_n227), .A4(new_n226), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n229), .A2(G131), .ZN(new_n240));
  OAI21_X1  g054(.A(KEYINPUT64), .B1(KEYINPUT0), .B2(G128), .ZN(new_n241));
  INV_X1    g055(.A(KEYINPUT64), .ZN(new_n242));
  INV_X1    g056(.A(KEYINPUT0), .ZN(new_n243));
  INV_X1    g057(.A(G128), .ZN(new_n244));
  NAND3_X1  g058(.A1(new_n242), .A2(new_n243), .A3(new_n244), .ZN(new_n245));
  NOR2_X1   g059(.A1(new_n205), .A2(G146), .ZN(new_n246));
  NOR2_X1   g060(.A1(new_n203), .A2(G143), .ZN(new_n247));
  OAI211_X1 g061(.A(new_n241), .B(new_n245), .C1(new_n246), .C2(new_n247), .ZN(new_n248));
  NAND2_X1  g062(.A1(KEYINPUT0), .A2(G128), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n248), .A2(new_n249), .ZN(new_n250));
  NAND3_X1  g064(.A1(new_n213), .A2(KEYINPUT0), .A3(G128), .ZN(new_n251));
  AOI22_X1  g065(.A1(new_n239), .A2(new_n240), .B1(new_n250), .B2(new_n251), .ZN(new_n252));
  OAI21_X1  g066(.A(new_n201), .B1(new_n234), .B2(new_n252), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n239), .A2(new_n240), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n250), .A2(new_n251), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n254), .A2(new_n255), .ZN(new_n256));
  INV_X1    g070(.A(KEYINPUT69), .ZN(new_n257));
  AND4_X1   g071(.A1(new_n188), .A2(new_n196), .A3(new_n190), .A4(new_n197), .ZN(new_n258));
  AOI22_X1  g072(.A1(new_n188), .A2(new_n190), .B1(new_n196), .B2(new_n197), .ZN(new_n259));
  OAI21_X1  g073(.A(new_n257), .B1(new_n258), .B2(new_n259), .ZN(new_n260));
  NAND3_X1  g074(.A1(new_n193), .A2(KEYINPUT69), .A3(new_n198), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  XNOR2_X1  g076(.A(G143), .B(G146), .ZN(new_n263));
  AOI21_X1  g077(.A(new_n244), .B1(new_n208), .B2(new_n209), .ZN(new_n264));
  AOI21_X1  g078(.A(new_n263), .B1(new_n264), .B2(new_n211), .ZN(new_n265));
  OAI211_X1 g079(.A(new_n239), .B(new_n222), .C1(new_n265), .C2(new_n207), .ZN(new_n266));
  NAND3_X1  g080(.A1(new_n256), .A2(new_n262), .A3(new_n266), .ZN(new_n267));
  NAND3_X1  g081(.A1(new_n253), .A2(KEYINPUT71), .A3(new_n267), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n256), .A2(new_n266), .ZN(new_n269));
  INV_X1    g083(.A(KEYINPUT71), .ZN(new_n270));
  NAND3_X1  g084(.A1(new_n269), .A2(new_n270), .A3(new_n201), .ZN(new_n271));
  NAND3_X1  g085(.A1(new_n268), .A2(KEYINPUT28), .A3(new_n271), .ZN(new_n272));
  INV_X1    g086(.A(KEYINPUT28), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n267), .A2(new_n273), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n272), .A2(new_n274), .ZN(new_n275));
  INV_X1    g089(.A(G237), .ZN(new_n276));
  INV_X1    g090(.A(G953), .ZN(new_n277));
  NAND3_X1  g091(.A1(new_n276), .A2(new_n277), .A3(G210), .ZN(new_n278));
  INV_X1    g092(.A(KEYINPUT27), .ZN(new_n279));
  XNOR2_X1  g093(.A(new_n278), .B(new_n279), .ZN(new_n280));
  XNOR2_X1  g094(.A(new_n280), .B(KEYINPUT26), .ZN(new_n281));
  XNOR2_X1  g095(.A(new_n281), .B(G101), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n275), .A2(new_n282), .ZN(new_n283));
  INV_X1    g097(.A(KEYINPUT30), .ZN(new_n284));
  OAI21_X1  g098(.A(new_n284), .B1(new_n234), .B2(new_n252), .ZN(new_n285));
  NAND3_X1  g099(.A1(new_n256), .A2(KEYINPUT30), .A3(new_n266), .ZN(new_n286));
  NAND3_X1  g100(.A1(new_n285), .A2(new_n201), .A3(new_n286), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n267), .A2(KEYINPUT70), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  INV_X1    g103(.A(new_n282), .ZN(new_n290));
  NAND4_X1  g104(.A1(new_n285), .A2(new_n286), .A3(KEYINPUT70), .A4(new_n201), .ZN(new_n291));
  NAND3_X1  g105(.A1(new_n289), .A2(new_n290), .A3(new_n291), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n292), .A2(KEYINPUT31), .ZN(new_n293));
  INV_X1    g107(.A(KEYINPUT31), .ZN(new_n294));
  NAND4_X1  g108(.A1(new_n289), .A2(new_n294), .A3(new_n290), .A4(new_n291), .ZN(new_n295));
  NAND3_X1  g109(.A1(new_n283), .A2(new_n293), .A3(new_n295), .ZN(new_n296));
  NOR2_X1   g110(.A1(G472), .A2(G902), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n296), .A2(new_n297), .ZN(new_n298));
  INV_X1    g112(.A(KEYINPUT32), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n298), .A2(new_n299), .ZN(new_n300));
  NAND3_X1  g114(.A1(new_n296), .A2(KEYINPUT32), .A3(new_n297), .ZN(new_n301));
  NAND3_X1  g115(.A1(new_n253), .A2(KEYINPUT72), .A3(new_n267), .ZN(new_n302));
  INV_X1    g116(.A(KEYINPUT72), .ZN(new_n303));
  NAND3_X1  g117(.A1(new_n269), .A2(new_n303), .A3(new_n201), .ZN(new_n304));
  NAND3_X1  g118(.A1(new_n302), .A2(KEYINPUT28), .A3(new_n304), .ZN(new_n305));
  AND2_X1   g119(.A1(new_n305), .A2(new_n274), .ZN(new_n306));
  INV_X1    g120(.A(KEYINPUT29), .ZN(new_n307));
  NOR2_X1   g121(.A1(new_n282), .A2(new_n307), .ZN(new_n308));
  AOI21_X1  g122(.A(G902), .B1(new_n306), .B2(new_n308), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n289), .A2(new_n291), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n310), .A2(new_n282), .ZN(new_n311));
  NAND3_X1  g125(.A1(new_n272), .A2(new_n274), .A3(new_n290), .ZN(new_n312));
  NAND3_X1  g126(.A1(new_n311), .A2(new_n307), .A3(new_n312), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n309), .A2(new_n313), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n314), .A2(G472), .ZN(new_n315));
  NAND3_X1  g129(.A1(new_n300), .A2(new_n301), .A3(new_n315), .ZN(new_n316));
  INV_X1    g130(.A(G140), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n317), .A2(G125), .ZN(new_n318));
  INV_X1    g132(.A(G125), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n319), .A2(G140), .ZN(new_n320));
  NAND3_X1  g134(.A1(new_n318), .A2(new_n320), .A3(KEYINPUT16), .ZN(new_n321));
  OAI21_X1  g135(.A(new_n321), .B1(KEYINPUT16), .B2(new_n318), .ZN(new_n322));
  XNOR2_X1  g136(.A(new_n322), .B(G146), .ZN(new_n323));
  INV_X1    g137(.A(new_n323), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n187), .A2(G128), .ZN(new_n325));
  XNOR2_X1  g139(.A(new_n325), .B(KEYINPUT74), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n244), .A2(G119), .ZN(new_n327));
  AND2_X1   g141(.A1(new_n326), .A2(new_n327), .ZN(new_n328));
  XOR2_X1   g142(.A(KEYINPUT24), .B(G110), .Z(new_n329));
  NAND2_X1  g143(.A1(new_n328), .A2(new_n329), .ZN(new_n330));
  INV_X1    g144(.A(KEYINPUT75), .ZN(new_n331));
  AOI21_X1  g145(.A(new_n331), .B1(new_n325), .B2(KEYINPUT23), .ZN(new_n332));
  XNOR2_X1  g146(.A(new_n332), .B(new_n327), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n333), .A2(G110), .ZN(new_n334));
  NAND3_X1  g148(.A1(new_n324), .A2(new_n330), .A3(new_n334), .ZN(new_n335));
  NAND3_X1  g149(.A1(new_n318), .A2(new_n320), .A3(new_n203), .ZN(new_n336));
  OR2_X1    g150(.A1(new_n322), .A2(new_n203), .ZN(new_n337));
  NOR2_X1   g151(.A1(new_n328), .A2(new_n329), .ZN(new_n338));
  NOR2_X1   g152(.A1(new_n333), .A2(G110), .ZN(new_n339));
  OAI211_X1 g153(.A(new_n336), .B(new_n337), .C1(new_n338), .C2(new_n339), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n335), .A2(new_n340), .ZN(new_n341));
  NAND3_X1  g155(.A1(new_n277), .A2(G221), .A3(G234), .ZN(new_n342));
  XNOR2_X1  g156(.A(new_n342), .B(KEYINPUT22), .ZN(new_n343));
  XNOR2_X1  g157(.A(new_n343), .B(G137), .ZN(new_n344));
  INV_X1    g158(.A(new_n344), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n341), .A2(new_n345), .ZN(new_n346));
  INV_X1    g160(.A(G902), .ZN(new_n347));
  NAND3_X1  g161(.A1(new_n335), .A2(new_n340), .A3(new_n344), .ZN(new_n348));
  NAND3_X1  g162(.A1(new_n346), .A2(new_n347), .A3(new_n348), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n349), .A2(KEYINPUT25), .ZN(new_n350));
  INV_X1    g164(.A(G234), .ZN(new_n351));
  OAI21_X1  g165(.A(G217), .B1(new_n351), .B2(G902), .ZN(new_n352));
  OR2_X1    g166(.A1(new_n352), .A2(KEYINPUT73), .ZN(new_n353));
  INV_X1    g167(.A(KEYINPUT25), .ZN(new_n354));
  NAND4_X1  g168(.A1(new_n346), .A2(new_n354), .A3(new_n347), .A4(new_n348), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n352), .A2(KEYINPUT73), .ZN(new_n356));
  NAND4_X1  g170(.A1(new_n350), .A2(new_n353), .A3(new_n355), .A4(new_n356), .ZN(new_n357));
  AND2_X1   g171(.A1(new_n346), .A2(new_n348), .ZN(new_n358));
  AOI21_X1  g172(.A(G902), .B1(new_n351), .B2(G217), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n358), .A2(new_n359), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n357), .A2(new_n360), .ZN(new_n361));
  INV_X1    g175(.A(new_n361), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n316), .A2(new_n362), .ZN(new_n363));
  INV_X1    g177(.A(KEYINPUT79), .ZN(new_n364));
  INV_X1    g178(.A(G104), .ZN(new_n365));
  OAI21_X1  g179(.A(KEYINPUT3), .B1(new_n365), .B2(G107), .ZN(new_n366));
  INV_X1    g180(.A(KEYINPUT3), .ZN(new_n367));
  INV_X1    g181(.A(G107), .ZN(new_n368));
  NAND3_X1  g182(.A1(new_n367), .A2(new_n368), .A3(G104), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n365), .A2(G107), .ZN(new_n370));
  NAND3_X1  g184(.A1(new_n366), .A2(new_n369), .A3(new_n370), .ZN(new_n371));
  INV_X1    g185(.A(KEYINPUT4), .ZN(new_n372));
  NAND3_X1  g186(.A1(new_n371), .A2(new_n372), .A3(G101), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n371), .A2(G101), .ZN(new_n374));
  INV_X1    g188(.A(G101), .ZN(new_n375));
  NAND4_X1  g189(.A1(new_n366), .A2(new_n369), .A3(new_n375), .A4(new_n370), .ZN(new_n376));
  NAND3_X1  g190(.A1(new_n374), .A2(KEYINPUT4), .A3(new_n376), .ZN(new_n377));
  NAND4_X1  g191(.A1(new_n201), .A2(new_n364), .A3(new_n373), .A4(new_n377), .ZN(new_n378));
  NAND4_X1  g192(.A1(new_n377), .A2(new_n260), .A3(new_n261), .A4(new_n373), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n379), .A2(KEYINPUT79), .ZN(new_n380));
  XNOR2_X1  g194(.A(KEYINPUT80), .B(KEYINPUT5), .ZN(new_n381));
  OAI21_X1  g195(.A(G113), .B1(new_n381), .B2(new_n188), .ZN(new_n382));
  INV_X1    g196(.A(new_n382), .ZN(new_n383));
  INV_X1    g197(.A(new_n191), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n384), .A2(new_n381), .ZN(new_n385));
  AOI21_X1  g199(.A(new_n258), .B1(new_n383), .B2(new_n385), .ZN(new_n386));
  NOR2_X1   g200(.A1(new_n368), .A2(G104), .ZN(new_n387));
  NOR2_X1   g201(.A1(new_n365), .A2(G107), .ZN(new_n388));
  OAI21_X1  g202(.A(G101), .B1(new_n387), .B2(new_n388), .ZN(new_n389));
  AND2_X1   g203(.A1(new_n376), .A2(new_n389), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n386), .A2(new_n390), .ZN(new_n391));
  NAND3_X1  g205(.A1(new_n378), .A2(new_n380), .A3(new_n391), .ZN(new_n392));
  XOR2_X1   g206(.A(G110), .B(G122), .Z(new_n393));
  NAND2_X1  g207(.A1(new_n392), .A2(new_n393), .ZN(new_n394));
  INV_X1    g208(.A(new_n393), .ZN(new_n395));
  NAND4_X1  g209(.A1(new_n378), .A2(new_n380), .A3(new_n395), .A4(new_n391), .ZN(new_n396));
  NAND3_X1  g210(.A1(new_n394), .A2(KEYINPUT6), .A3(new_n396), .ZN(new_n397));
  NAND3_X1  g211(.A1(new_n250), .A2(G125), .A3(new_n251), .ZN(new_n398));
  AOI22_X1  g212(.A1(new_n398), .A2(KEYINPUT81), .B1(new_n214), .B2(new_n319), .ZN(new_n399));
  OR2_X1    g213(.A1(new_n398), .A2(KEYINPUT81), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n399), .A2(new_n400), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n277), .A2(G224), .ZN(new_n402));
  XNOR2_X1  g216(.A(new_n402), .B(KEYINPUT82), .ZN(new_n403));
  INV_X1    g217(.A(new_n403), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n401), .A2(new_n404), .ZN(new_n405));
  NAND3_X1  g219(.A1(new_n399), .A2(new_n400), .A3(new_n403), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n405), .A2(new_n406), .ZN(new_n407));
  INV_X1    g221(.A(KEYINPUT6), .ZN(new_n408));
  NAND3_X1  g222(.A1(new_n392), .A2(new_n408), .A3(new_n393), .ZN(new_n409));
  NAND3_X1  g223(.A1(new_n397), .A2(new_n407), .A3(new_n409), .ZN(new_n410));
  INV_X1    g224(.A(KEYINPUT83), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n410), .A2(new_n411), .ZN(new_n412));
  INV_X1    g226(.A(new_n396), .ZN(new_n413));
  INV_X1    g227(.A(new_n406), .ZN(new_n414));
  AOI21_X1  g228(.A(new_n413), .B1(new_n414), .B2(KEYINPUT7), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n214), .A2(new_n319), .ZN(new_n416));
  INV_X1    g230(.A(KEYINPUT85), .ZN(new_n417));
  XNOR2_X1  g231(.A(new_n416), .B(new_n417), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n418), .A2(new_n398), .ZN(new_n419));
  INV_X1    g233(.A(KEYINPUT86), .ZN(new_n420));
  OR2_X1    g234(.A1(new_n420), .A2(KEYINPUT7), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n420), .A2(KEYINPUT7), .ZN(new_n422));
  NAND3_X1  g236(.A1(new_n403), .A2(new_n421), .A3(new_n422), .ZN(new_n423));
  OR3_X1    g237(.A1(new_n386), .A2(KEYINPUT84), .A3(new_n390), .ZN(new_n424));
  AND2_X1   g238(.A1(new_n384), .A2(KEYINPUT5), .ZN(new_n425));
  OAI211_X1 g239(.A(new_n390), .B(new_n198), .C1(new_n425), .C2(new_n382), .ZN(new_n426));
  OAI21_X1  g240(.A(KEYINPUT84), .B1(new_n386), .B2(new_n390), .ZN(new_n427));
  NAND3_X1  g241(.A1(new_n424), .A2(new_n426), .A3(new_n427), .ZN(new_n428));
  XOR2_X1   g242(.A(new_n393), .B(KEYINPUT8), .Z(new_n429));
  AOI22_X1  g243(.A1(new_n419), .A2(new_n423), .B1(new_n428), .B2(new_n429), .ZN(new_n430));
  AOI21_X1  g244(.A(G902), .B1(new_n415), .B2(new_n430), .ZN(new_n431));
  NAND4_X1  g245(.A1(new_n397), .A2(new_n407), .A3(KEYINPUT83), .A4(new_n409), .ZN(new_n432));
  NAND3_X1  g246(.A1(new_n412), .A2(new_n431), .A3(new_n432), .ZN(new_n433));
  OAI21_X1  g247(.A(G210), .B1(G237), .B2(G902), .ZN(new_n434));
  INV_X1    g248(.A(new_n434), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n433), .A2(new_n435), .ZN(new_n436));
  NAND4_X1  g250(.A1(new_n412), .A2(new_n431), .A3(new_n434), .A4(new_n432), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n436), .A2(new_n437), .ZN(new_n438));
  OAI21_X1  g252(.A(G214), .B1(G237), .B2(G902), .ZN(new_n439));
  XNOR2_X1  g253(.A(new_n439), .B(KEYINPUT78), .ZN(new_n440));
  INV_X1    g254(.A(new_n440), .ZN(new_n441));
  XOR2_X1   g255(.A(KEYINPUT9), .B(G234), .Z(new_n442));
  XNOR2_X1  g256(.A(new_n442), .B(KEYINPUT76), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n443), .A2(new_n347), .ZN(new_n444));
  AND2_X1   g258(.A1(new_n444), .A2(G221), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n212), .A2(new_n213), .ZN(new_n446));
  INV_X1    g260(.A(new_n207), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n376), .A2(new_n389), .ZN(new_n448));
  NAND3_X1  g262(.A1(new_n446), .A2(new_n447), .A3(new_n448), .ZN(new_n449));
  AOI21_X1  g263(.A(new_n263), .B1(G128), .B2(new_n208), .ZN(new_n450));
  OAI211_X1 g264(.A(new_n376), .B(new_n389), .C1(new_n450), .C2(new_n207), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n449), .A2(new_n451), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n452), .A2(new_n254), .ZN(new_n453));
  INV_X1    g267(.A(KEYINPUT12), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  NAND3_X1  g269(.A1(new_n452), .A2(KEYINPUT12), .A3(new_n254), .ZN(new_n456));
  NAND3_X1  g270(.A1(new_n455), .A2(KEYINPUT77), .A3(new_n456), .ZN(new_n457));
  INV_X1    g271(.A(KEYINPUT77), .ZN(new_n458));
  AOI221_X4 g272(.A(new_n454), .B1(new_n240), .B2(new_n239), .C1(new_n449), .C2(new_n451), .ZN(new_n459));
  AOI21_X1  g273(.A(KEYINPUT12), .B1(new_n452), .B2(new_n254), .ZN(new_n460));
  OAI21_X1  g274(.A(new_n458), .B1(new_n459), .B2(new_n460), .ZN(new_n461));
  INV_X1    g275(.A(KEYINPUT10), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n451), .A2(new_n462), .ZN(new_n463));
  NAND3_X1  g277(.A1(new_n255), .A2(new_n377), .A3(new_n373), .ZN(new_n464));
  INV_X1    g278(.A(new_n254), .ZN(new_n465));
  OAI211_X1 g279(.A(new_n390), .B(KEYINPUT10), .C1(new_n265), .C2(new_n207), .ZN(new_n466));
  NAND4_X1  g280(.A1(new_n463), .A2(new_n464), .A3(new_n465), .A4(new_n466), .ZN(new_n467));
  XNOR2_X1  g281(.A(G110), .B(G140), .ZN(new_n468));
  AND2_X1   g282(.A1(new_n277), .A2(G227), .ZN(new_n469));
  XOR2_X1   g283(.A(new_n468), .B(new_n469), .Z(new_n470));
  AND2_X1   g284(.A1(new_n467), .A2(new_n470), .ZN(new_n471));
  NAND3_X1  g285(.A1(new_n457), .A2(new_n461), .A3(new_n471), .ZN(new_n472));
  NAND3_X1  g286(.A1(new_n463), .A2(new_n464), .A3(new_n466), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n473), .A2(new_n254), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n474), .A2(new_n467), .ZN(new_n475));
  INV_X1    g289(.A(new_n470), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n472), .A2(new_n477), .ZN(new_n478));
  INV_X1    g292(.A(G469), .ZN(new_n479));
  NAND3_X1  g293(.A1(new_n478), .A2(new_n479), .A3(new_n347), .ZN(new_n480));
  OAI21_X1  g294(.A(new_n467), .B1(new_n459), .B2(new_n460), .ZN(new_n481));
  AOI22_X1  g295(.A1(new_n481), .A2(new_n476), .B1(new_n471), .B2(new_n474), .ZN(new_n482));
  OAI21_X1  g296(.A(G469), .B1(new_n482), .B2(G902), .ZN(new_n483));
  AOI21_X1  g297(.A(new_n445), .B1(new_n480), .B2(new_n483), .ZN(new_n484));
  NAND3_X1  g298(.A1(new_n438), .A2(new_n441), .A3(new_n484), .ZN(new_n485));
  NOR2_X1   g299(.A1(new_n363), .A2(new_n485), .ZN(new_n486));
  INV_X1    g300(.A(KEYINPUT87), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n487), .A2(new_n205), .ZN(new_n488));
  NOR2_X1   g302(.A1(G237), .A2(G953), .ZN(new_n489));
  NAND2_X1  g303(.A1(KEYINPUT87), .A2(G143), .ZN(new_n490));
  NAND4_X1  g304(.A1(new_n488), .A2(G214), .A3(new_n489), .A4(new_n490), .ZN(new_n491));
  NAND3_X1  g305(.A1(new_n276), .A2(new_n277), .A3(G214), .ZN(new_n492));
  INV_X1    g306(.A(new_n490), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n491), .A2(new_n494), .ZN(new_n495));
  INV_X1    g309(.A(KEYINPUT17), .ZN(new_n496));
  NOR3_X1   g310(.A1(new_n495), .A2(new_n496), .A3(new_n238), .ZN(new_n497));
  AND3_X1   g311(.A1(new_n491), .A2(new_n494), .A3(new_n232), .ZN(new_n498));
  AOI21_X1  g312(.A(new_n232), .B1(new_n491), .B2(new_n494), .ZN(new_n499));
  NOR2_X1   g313(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  AOI21_X1  g314(.A(new_n497), .B1(new_n500), .B2(new_n496), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n501), .A2(new_n323), .ZN(new_n502));
  XNOR2_X1  g316(.A(G113), .B(G122), .ZN(new_n503));
  XNOR2_X1  g317(.A(new_n503), .B(new_n365), .ZN(new_n504));
  XNOR2_X1  g318(.A(new_n504), .B(KEYINPUT90), .ZN(new_n505));
  INV_X1    g319(.A(KEYINPUT89), .ZN(new_n506));
  INV_X1    g320(.A(KEYINPUT88), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n495), .A2(new_n507), .ZN(new_n508));
  NAND2_X1  g322(.A1(KEYINPUT18), .A2(G131), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  NAND4_X1  g324(.A1(new_n495), .A2(new_n507), .A3(KEYINPUT18), .A4(G131), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n318), .A2(new_n320), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n513), .A2(G146), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n514), .A2(new_n336), .ZN(new_n515));
  AOI21_X1  g329(.A(new_n506), .B1(new_n512), .B2(new_n515), .ZN(new_n516));
  AOI22_X1  g330(.A1(new_n495), .A2(new_n507), .B1(KEYINPUT18), .B2(G131), .ZN(new_n517));
  AOI211_X1 g331(.A(KEYINPUT88), .B(new_n509), .C1(new_n491), .C2(new_n494), .ZN(new_n518));
  OAI211_X1 g332(.A(new_n506), .B(new_n515), .C1(new_n517), .C2(new_n518), .ZN(new_n519));
  INV_X1    g333(.A(new_n519), .ZN(new_n520));
  OAI211_X1 g334(.A(new_n502), .B(new_n505), .C1(new_n516), .C2(new_n520), .ZN(new_n521));
  INV_X1    g335(.A(new_n521), .ZN(new_n522));
  OAI21_X1  g336(.A(new_n515), .B1(new_n517), .B2(new_n518), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n523), .A2(KEYINPUT89), .ZN(new_n524));
  AOI22_X1  g338(.A1(new_n524), .A2(new_n519), .B1(new_n323), .B2(new_n501), .ZN(new_n525));
  INV_X1    g339(.A(KEYINPUT92), .ZN(new_n526));
  AOI21_X1  g340(.A(new_n504), .B1(new_n525), .B2(new_n526), .ZN(new_n527));
  OAI21_X1  g341(.A(new_n502), .B1(new_n516), .B2(new_n520), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n528), .A2(KEYINPUT92), .ZN(new_n529));
  AOI21_X1  g343(.A(new_n522), .B1(new_n527), .B2(new_n529), .ZN(new_n530));
  OAI21_X1  g344(.A(KEYINPUT93), .B1(new_n530), .B2(G902), .ZN(new_n531));
  XOR2_X1   g345(.A(KEYINPUT91), .B(G475), .Z(new_n532));
  OAI211_X1 g346(.A(new_n526), .B(new_n502), .C1(new_n516), .C2(new_n520), .ZN(new_n533));
  INV_X1    g347(.A(new_n504), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  NOR2_X1   g349(.A1(new_n525), .A2(new_n526), .ZN(new_n536));
  OAI21_X1  g350(.A(new_n521), .B1(new_n535), .B2(new_n536), .ZN(new_n537));
  INV_X1    g351(.A(KEYINPUT93), .ZN(new_n538));
  NAND3_X1  g352(.A1(new_n537), .A2(new_n538), .A3(new_n347), .ZN(new_n539));
  NAND3_X1  g353(.A1(new_n531), .A2(new_n532), .A3(new_n539), .ZN(new_n540));
  INV_X1    g354(.A(G475), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n524), .A2(new_n519), .ZN(new_n542));
  XNOR2_X1  g356(.A(new_n513), .B(KEYINPUT19), .ZN(new_n543));
  OAI221_X1 g357(.A(new_n337), .B1(new_n498), .B2(new_n499), .C1(G146), .C2(new_n543), .ZN(new_n544));
  AOI21_X1  g358(.A(new_n504), .B1(new_n542), .B2(new_n544), .ZN(new_n545));
  OAI211_X1 g359(.A(new_n541), .B(new_n347), .C1(new_n522), .C2(new_n545), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n546), .A2(KEYINPUT20), .ZN(new_n547));
  AND2_X1   g361(.A1(new_n542), .A2(new_n544), .ZN(new_n548));
  OAI21_X1  g362(.A(new_n521), .B1(new_n548), .B2(new_n504), .ZN(new_n549));
  INV_X1    g363(.A(KEYINPUT20), .ZN(new_n550));
  NAND4_X1  g364(.A1(new_n549), .A2(new_n550), .A3(new_n541), .A4(new_n347), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n547), .A2(new_n551), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n205), .A2(G128), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n244), .A2(G143), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n555), .A2(G134), .ZN(new_n556));
  NAND3_X1  g370(.A1(new_n553), .A2(new_n554), .A3(new_n219), .ZN(new_n557));
  INV_X1    g371(.A(G122), .ZN(new_n558));
  OAI21_X1  g372(.A(KEYINPUT14), .B1(new_n558), .B2(G116), .ZN(new_n559));
  INV_X1    g373(.A(KEYINPUT14), .ZN(new_n560));
  NAND3_X1  g374(.A1(new_n560), .A2(new_n189), .A3(G122), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n558), .A2(G116), .ZN(new_n562));
  NAND3_X1  g376(.A1(new_n559), .A2(new_n561), .A3(new_n562), .ZN(new_n563));
  AOI22_X1  g377(.A1(new_n556), .A2(new_n557), .B1(new_n563), .B2(G107), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n189), .A2(G122), .ZN(new_n565));
  NAND3_X1  g379(.A1(new_n562), .A2(new_n565), .A3(new_n368), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n566), .A2(KEYINPUT94), .ZN(new_n567));
  OR2_X1    g381(.A1(new_n566), .A2(KEYINPUT94), .ZN(new_n568));
  NAND3_X1  g382(.A1(new_n564), .A2(new_n567), .A3(new_n568), .ZN(new_n569));
  INV_X1    g383(.A(KEYINPUT13), .ZN(new_n570));
  OAI21_X1  g384(.A(new_n554), .B1(new_n553), .B2(new_n570), .ZN(new_n571));
  NOR2_X1   g385(.A1(new_n244), .A2(G143), .ZN(new_n572));
  NOR2_X1   g386(.A1(new_n572), .A2(KEYINPUT13), .ZN(new_n573));
  OAI21_X1  g387(.A(G134), .B1(new_n571), .B2(new_n573), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n562), .A2(new_n565), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n575), .A2(G107), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n576), .A2(new_n566), .ZN(new_n577));
  NAND3_X1  g391(.A1(new_n574), .A2(new_n577), .A3(new_n557), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n569), .A2(new_n578), .ZN(new_n579));
  NAND3_X1  g393(.A1(new_n443), .A2(G217), .A3(new_n277), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  INV_X1    g395(.A(new_n581), .ZN(new_n582));
  NOR2_X1   g396(.A1(new_n579), .A2(new_n580), .ZN(new_n583));
  OAI21_X1  g397(.A(new_n347), .B1(new_n582), .B2(new_n583), .ZN(new_n584));
  INV_X1    g398(.A(G478), .ZN(new_n585));
  NOR2_X1   g399(.A1(new_n585), .A2(KEYINPUT15), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n584), .A2(new_n586), .ZN(new_n587));
  XNOR2_X1  g401(.A(new_n579), .B(new_n580), .ZN(new_n588));
  INV_X1    g402(.A(new_n586), .ZN(new_n589));
  NAND3_X1  g403(.A1(new_n588), .A2(new_n347), .A3(new_n589), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n587), .A2(new_n590), .ZN(new_n591));
  INV_X1    g405(.A(KEYINPUT95), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  NAND3_X1  g407(.A1(new_n587), .A2(new_n590), .A3(KEYINPUT95), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  INV_X1    g409(.A(G952), .ZN(new_n596));
  NOR2_X1   g410(.A1(new_n596), .A2(G953), .ZN(new_n597));
  NAND2_X1  g411(.A1(G234), .A2(G237), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  XOR2_X1   g413(.A(KEYINPUT21), .B(G898), .Z(new_n600));
  NAND3_X1  g414(.A1(new_n598), .A2(G902), .A3(G953), .ZN(new_n601));
  OAI21_X1  g415(.A(new_n599), .B1(new_n600), .B2(new_n601), .ZN(new_n602));
  NAND4_X1  g416(.A1(new_n540), .A2(new_n552), .A3(new_n595), .A4(new_n602), .ZN(new_n603));
  OR2_X1    g417(.A1(new_n603), .A2(KEYINPUT96), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n603), .A2(KEYINPUT96), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n486), .A2(new_n606), .ZN(new_n607));
  XNOR2_X1  g421(.A(new_n607), .B(G101), .ZN(G3));
  NAND2_X1  g422(.A1(new_n296), .A2(new_n347), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n609), .A2(G472), .ZN(new_n610));
  INV_X1    g424(.A(KEYINPUT97), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n298), .A2(new_n611), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n610), .A2(new_n612), .ZN(new_n613));
  NAND3_X1  g427(.A1(new_n609), .A2(new_n611), .A3(G472), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  INV_X1    g429(.A(new_n445), .ZN(new_n616));
  AOI211_X1 g430(.A(G469), .B(G902), .C1(new_n472), .C2(new_n477), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n481), .A2(new_n476), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n471), .A2(new_n474), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  AOI21_X1  g434(.A(new_n479), .B1(new_n620), .B2(new_n347), .ZN(new_n621));
  OAI21_X1  g435(.A(new_n616), .B1(new_n617), .B2(new_n621), .ZN(new_n622));
  NOR2_X1   g436(.A1(new_n615), .A2(new_n622), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n623), .A2(new_n362), .ZN(new_n624));
  XNOR2_X1  g438(.A(new_n624), .B(KEYINPUT98), .ZN(new_n625));
  AOI21_X1  g439(.A(new_n440), .B1(new_n436), .B2(new_n437), .ZN(new_n626));
  NOR2_X1   g440(.A1(new_n585), .A2(new_n347), .ZN(new_n627));
  INV_X1    g441(.A(new_n627), .ZN(new_n628));
  NAND3_X1  g442(.A1(new_n588), .A2(new_n585), .A3(new_n347), .ZN(new_n629));
  XNOR2_X1  g443(.A(KEYINPUT99), .B(KEYINPUT33), .ZN(new_n630));
  AND2_X1   g444(.A1(new_n588), .A2(new_n630), .ZN(new_n631));
  INV_X1    g445(.A(KEYINPUT33), .ZN(new_n632));
  INV_X1    g446(.A(KEYINPUT100), .ZN(new_n633));
  AOI21_X1  g447(.A(new_n632), .B1(new_n588), .B2(new_n633), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n581), .A2(KEYINPUT100), .ZN(new_n635));
  AOI21_X1  g449(.A(new_n631), .B1(new_n634), .B2(new_n635), .ZN(new_n636));
  OAI211_X1 g450(.A(new_n628), .B(new_n629), .C1(new_n636), .C2(new_n585), .ZN(new_n637));
  AOI21_X1  g451(.A(new_n637), .B1(new_n540), .B2(new_n552), .ZN(new_n638));
  NAND3_X1  g452(.A1(new_n626), .A2(new_n602), .A3(new_n638), .ZN(new_n639));
  INV_X1    g453(.A(new_n639), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n625), .A2(new_n640), .ZN(new_n641));
  XOR2_X1   g455(.A(KEYINPUT34), .B(G104), .Z(new_n642));
  XNOR2_X1  g456(.A(new_n641), .B(new_n642), .ZN(G6));
  AND2_X1   g457(.A1(new_n593), .A2(new_n594), .ZN(new_n644));
  NAND3_X1  g458(.A1(new_n546), .A2(KEYINPUT101), .A3(KEYINPUT20), .ZN(new_n645));
  INV_X1    g459(.A(KEYINPUT101), .ZN(new_n646));
  NAND3_X1  g460(.A1(new_n547), .A2(new_n551), .A3(new_n646), .ZN(new_n647));
  AND4_X1   g461(.A1(new_n540), .A2(new_n644), .A3(new_n645), .A4(new_n647), .ZN(new_n648));
  AND3_X1   g462(.A1(new_n626), .A2(new_n648), .A3(new_n602), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n625), .A2(new_n649), .ZN(new_n650));
  XOR2_X1   g464(.A(new_n650), .B(KEYINPUT102), .Z(new_n651));
  XNOR2_X1  g465(.A(new_n651), .B(KEYINPUT35), .ZN(new_n652));
  XNOR2_X1  g466(.A(new_n652), .B(new_n368), .ZN(G9));
  NOR2_X1   g467(.A1(new_n345), .A2(KEYINPUT36), .ZN(new_n654));
  XNOR2_X1  g468(.A(new_n341), .B(new_n654), .ZN(new_n655));
  NAND2_X1  g469(.A1(new_n655), .A2(new_n359), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n357), .A2(new_n656), .ZN(new_n657));
  AND2_X1   g471(.A1(new_n603), .A2(KEYINPUT96), .ZN(new_n658));
  NOR2_X1   g472(.A1(new_n603), .A2(KEYINPUT96), .ZN(new_n659));
  OAI21_X1  g473(.A(new_n657), .B1(new_n658), .B2(new_n659), .ZN(new_n660));
  NAND4_X1  g474(.A1(new_n626), .A2(new_n613), .A3(new_n484), .A4(new_n614), .ZN(new_n661));
  NOR2_X1   g475(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  XNOR2_X1  g476(.A(new_n662), .B(KEYINPUT37), .ZN(new_n663));
  XNOR2_X1  g477(.A(new_n663), .B(G110), .ZN(G12));
  INV_X1    g478(.A(new_n657), .ZN(new_n665));
  AND3_X1   g479(.A1(new_n296), .A2(KEYINPUT32), .A3(new_n297), .ZN(new_n666));
  AOI21_X1  g480(.A(KEYINPUT32), .B1(new_n296), .B2(new_n297), .ZN(new_n667));
  NOR2_X1   g481(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  AOI21_X1  g482(.A(new_n665), .B1(new_n668), .B2(new_n315), .ZN(new_n669));
  AOI211_X1 g483(.A(new_n440), .B(new_n622), .C1(new_n436), .C2(new_n437), .ZN(new_n670));
  NAND3_X1  g484(.A1(new_n540), .A2(new_n645), .A3(new_n647), .ZN(new_n671));
  OAI21_X1  g485(.A(new_n599), .B1(new_n601), .B2(G900), .ZN(new_n672));
  INV_X1    g486(.A(new_n672), .ZN(new_n673));
  NOR3_X1   g487(.A1(new_n671), .A2(new_n595), .A3(new_n673), .ZN(new_n674));
  NAND3_X1  g488(.A1(new_n669), .A2(new_n670), .A3(new_n674), .ZN(new_n675));
  XNOR2_X1  g489(.A(new_n675), .B(G128), .ZN(G30));
  AND2_X1   g490(.A1(new_n302), .A2(new_n304), .ZN(new_n677));
  OAI21_X1  g491(.A(new_n347), .B1(new_n677), .B2(new_n290), .ZN(new_n678));
  AOI21_X1  g492(.A(new_n282), .B1(new_n289), .B2(new_n291), .ZN(new_n679));
  OAI21_X1  g493(.A(G472), .B1(new_n678), .B2(new_n679), .ZN(new_n680));
  NAND2_X1  g494(.A1(new_n668), .A2(new_n680), .ZN(new_n681));
  AOI21_X1  g495(.A(new_n595), .B1(new_n540), .B2(new_n552), .ZN(new_n682));
  NAND2_X1  g496(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  INV_X1    g497(.A(KEYINPUT38), .ZN(new_n684));
  NAND2_X1  g498(.A1(new_n438), .A2(new_n684), .ZN(new_n685));
  NAND3_X1  g499(.A1(new_n436), .A2(KEYINPUT38), .A3(new_n437), .ZN(new_n686));
  NAND3_X1  g500(.A1(new_n685), .A2(new_n665), .A3(new_n686), .ZN(new_n687));
  XOR2_X1   g501(.A(new_n672), .B(KEYINPUT39), .Z(new_n688));
  INV_X1    g502(.A(new_n688), .ZN(new_n689));
  NAND2_X1  g503(.A1(new_n484), .A2(new_n689), .ZN(new_n690));
  XNOR2_X1  g504(.A(new_n690), .B(KEYINPUT40), .ZN(new_n691));
  NOR4_X1   g505(.A1(new_n683), .A2(new_n687), .A3(new_n691), .A4(new_n440), .ZN(new_n692));
  XNOR2_X1  g506(.A(new_n692), .B(new_n205), .ZN(G45));
  NAND2_X1  g507(.A1(new_n540), .A2(new_n552), .ZN(new_n694));
  INV_X1    g508(.A(new_n637), .ZN(new_n695));
  NAND3_X1  g509(.A1(new_n694), .A2(new_n695), .A3(new_n672), .ZN(new_n696));
  INV_X1    g510(.A(new_n696), .ZN(new_n697));
  NAND3_X1  g511(.A1(new_n669), .A2(new_n670), .A3(new_n697), .ZN(new_n698));
  XNOR2_X1  g512(.A(new_n698), .B(G146), .ZN(G48));
  NAND2_X1  g513(.A1(new_n478), .A2(new_n347), .ZN(new_n700));
  NAND2_X1  g514(.A1(new_n700), .A2(G469), .ZN(new_n701));
  NAND3_X1  g515(.A1(new_n701), .A2(new_n616), .A3(new_n480), .ZN(new_n702));
  INV_X1    g516(.A(KEYINPUT103), .ZN(new_n703));
  NAND2_X1  g517(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  AOI21_X1  g518(.A(new_n479), .B1(new_n478), .B2(new_n347), .ZN(new_n705));
  NOR2_X1   g519(.A1(new_n705), .A2(new_n617), .ZN(new_n706));
  NAND3_X1  g520(.A1(new_n706), .A2(KEYINPUT103), .A3(new_n616), .ZN(new_n707));
  NAND4_X1  g521(.A1(new_n316), .A2(new_n362), .A3(new_n704), .A4(new_n707), .ZN(new_n708));
  NOR2_X1   g522(.A1(new_n708), .A2(new_n639), .ZN(new_n709));
  XOR2_X1   g523(.A(KEYINPUT41), .B(G113), .Z(new_n710));
  XNOR2_X1  g524(.A(new_n709), .B(new_n710), .ZN(G15));
  NAND3_X1  g525(.A1(new_n626), .A2(new_n648), .A3(new_n602), .ZN(new_n712));
  NOR2_X1   g526(.A1(new_n708), .A2(new_n712), .ZN(new_n713));
  XNOR2_X1  g527(.A(new_n713), .B(new_n189), .ZN(G18));
  NAND3_X1  g528(.A1(new_n626), .A2(new_n704), .A3(new_n707), .ZN(new_n715));
  INV_X1    g529(.A(new_n715), .ZN(new_n716));
  NAND3_X1  g530(.A1(new_n606), .A2(new_n716), .A3(new_n669), .ZN(new_n717));
  XNOR2_X1  g531(.A(new_n717), .B(G119), .ZN(G21));
  NAND3_X1  g532(.A1(new_n438), .A2(new_n602), .A3(new_n441), .ZN(new_n719));
  OAI211_X1 g533(.A(new_n293), .B(new_n295), .C1(new_n290), .C2(new_n306), .ZN(new_n720));
  NAND2_X1  g534(.A1(new_n720), .A2(new_n297), .ZN(new_n721));
  NAND3_X1  g535(.A1(new_n610), .A2(new_n362), .A3(new_n721), .ZN(new_n722));
  NOR2_X1   g536(.A1(new_n719), .A2(new_n722), .ZN(new_n723));
  NAND3_X1  g537(.A1(new_n704), .A2(new_n707), .A3(new_n682), .ZN(new_n724));
  INV_X1    g538(.A(new_n724), .ZN(new_n725));
  NAND3_X1  g539(.A1(new_n723), .A2(KEYINPUT104), .A3(new_n725), .ZN(new_n726));
  INV_X1    g540(.A(KEYINPUT104), .ZN(new_n727));
  AOI22_X1  g541(.A1(new_n609), .A2(G472), .B1(new_n297), .B2(new_n720), .ZN(new_n728));
  NAND4_X1  g542(.A1(new_n626), .A2(new_n602), .A3(new_n362), .A4(new_n728), .ZN(new_n729));
  OAI21_X1  g543(.A(new_n727), .B1(new_n729), .B2(new_n724), .ZN(new_n730));
  NAND2_X1  g544(.A1(new_n726), .A2(new_n730), .ZN(new_n731));
  XNOR2_X1  g545(.A(new_n731), .B(G122), .ZN(G24));
  NAND2_X1  g546(.A1(new_n728), .A2(new_n657), .ZN(new_n733));
  INV_X1    g547(.A(KEYINPUT105), .ZN(new_n734));
  NAND2_X1  g548(.A1(new_n696), .A2(new_n734), .ZN(new_n735));
  NAND3_X1  g549(.A1(new_n638), .A2(KEYINPUT105), .A3(new_n672), .ZN(new_n736));
  AOI21_X1  g550(.A(new_n733), .B1(new_n735), .B2(new_n736), .ZN(new_n737));
  NAND2_X1  g551(.A1(new_n737), .A2(new_n716), .ZN(new_n738));
  XNOR2_X1  g552(.A(new_n738), .B(G125), .ZN(G27));
  NAND2_X1  g553(.A1(new_n735), .A2(new_n736), .ZN(new_n740));
  INV_X1    g554(.A(G472), .ZN(new_n741));
  AOI21_X1  g555(.A(new_n741), .B1(new_n309), .B2(new_n313), .ZN(new_n742));
  NOR3_X1   g556(.A1(new_n666), .A2(new_n667), .A3(new_n742), .ZN(new_n743));
  NAND4_X1  g557(.A1(new_n436), .A2(new_n441), .A3(new_n484), .A4(new_n437), .ZN(new_n744));
  NOR3_X1   g558(.A1(new_n743), .A2(new_n744), .A3(new_n361), .ZN(new_n745));
  NAND2_X1  g559(.A1(new_n740), .A2(new_n745), .ZN(new_n746));
  INV_X1    g560(.A(KEYINPUT42), .ZN(new_n747));
  NOR2_X1   g561(.A1(new_n747), .A2(KEYINPUT106), .ZN(new_n748));
  INV_X1    g562(.A(new_n748), .ZN(new_n749));
  NAND2_X1  g563(.A1(new_n746), .A2(new_n749), .ZN(new_n750));
  XOR2_X1   g564(.A(KEYINPUT106), .B(KEYINPUT42), .Z(new_n751));
  NAND3_X1  g565(.A1(new_n740), .A2(new_n745), .A3(new_n751), .ZN(new_n752));
  NAND2_X1  g566(.A1(new_n750), .A2(new_n752), .ZN(new_n753));
  XNOR2_X1  g567(.A(new_n753), .B(G131), .ZN(G33));
  NAND2_X1  g568(.A1(new_n745), .A2(new_n674), .ZN(new_n755));
  XNOR2_X1  g569(.A(new_n755), .B(G134), .ZN(G36));
  INV_X1    g570(.A(KEYINPUT46), .ZN(new_n757));
  INV_X1    g571(.A(KEYINPUT45), .ZN(new_n758));
  XNOR2_X1  g572(.A(new_n482), .B(new_n758), .ZN(new_n759));
  OAI211_X1 g573(.A(new_n757), .B(G469), .C1(new_n759), .C2(G902), .ZN(new_n760));
  NAND2_X1  g574(.A1(new_n620), .A2(new_n758), .ZN(new_n761));
  NAND2_X1  g575(.A1(new_n482), .A2(KEYINPUT45), .ZN(new_n762));
  NAND3_X1  g576(.A1(new_n761), .A2(new_n762), .A3(G469), .ZN(new_n763));
  NAND2_X1  g577(.A1(G469), .A2(G902), .ZN(new_n764));
  NAND3_X1  g578(.A1(new_n763), .A2(KEYINPUT46), .A3(new_n764), .ZN(new_n765));
  NAND3_X1  g579(.A1(new_n760), .A2(new_n480), .A3(new_n765), .ZN(new_n766));
  NAND2_X1  g580(.A1(new_n766), .A2(new_n616), .ZN(new_n767));
  NOR2_X1   g581(.A1(new_n767), .A2(new_n688), .ZN(new_n768));
  INV_X1    g582(.A(new_n768), .ZN(new_n769));
  INV_X1    g583(.A(KEYINPUT43), .ZN(new_n770));
  OAI21_X1  g584(.A(new_n770), .B1(new_n694), .B2(new_n637), .ZN(new_n771));
  NAND4_X1  g585(.A1(new_n695), .A2(KEYINPUT43), .A3(new_n552), .A4(new_n540), .ZN(new_n772));
  AOI21_X1  g586(.A(new_n665), .B1(new_n771), .B2(new_n772), .ZN(new_n773));
  NAND3_X1  g587(.A1(new_n773), .A2(KEYINPUT44), .A3(new_n615), .ZN(new_n774));
  OR2_X1    g588(.A1(new_n774), .A2(KEYINPUT107), .ZN(new_n775));
  NAND2_X1  g589(.A1(new_n774), .A2(KEYINPUT107), .ZN(new_n776));
  AOI21_X1  g590(.A(new_n769), .B1(new_n775), .B2(new_n776), .ZN(new_n777));
  AOI21_X1  g591(.A(KEYINPUT44), .B1(new_n773), .B2(new_n615), .ZN(new_n778));
  NAND3_X1  g592(.A1(new_n436), .A2(new_n441), .A3(new_n437), .ZN(new_n779));
  NOR2_X1   g593(.A1(new_n778), .A2(new_n779), .ZN(new_n780));
  NAND2_X1  g594(.A1(new_n777), .A2(new_n780), .ZN(new_n781));
  XNOR2_X1  g595(.A(new_n781), .B(G137), .ZN(G39));
  NAND2_X1  g596(.A1(new_n767), .A2(KEYINPUT47), .ZN(new_n783));
  INV_X1    g597(.A(KEYINPUT47), .ZN(new_n784));
  NAND3_X1  g598(.A1(new_n766), .A2(new_n784), .A3(new_n616), .ZN(new_n785));
  NAND2_X1  g599(.A1(new_n783), .A2(new_n785), .ZN(new_n786));
  NAND3_X1  g600(.A1(new_n697), .A2(new_n743), .A3(new_n361), .ZN(new_n787));
  NOR3_X1   g601(.A1(new_n786), .A2(new_n779), .A3(new_n787), .ZN(new_n788));
  XNOR2_X1  g602(.A(new_n788), .B(KEYINPUT108), .ZN(new_n789));
  XNOR2_X1  g603(.A(new_n789), .B(G140), .ZN(G42));
  NAND2_X1  g604(.A1(new_n704), .A2(new_n707), .ZN(new_n791));
  NOR2_X1   g605(.A1(new_n791), .A2(new_n779), .ZN(new_n792));
  INV_X1    g606(.A(new_n792), .ZN(new_n793));
  OR2_X1    g607(.A1(new_n361), .A2(new_n599), .ZN(new_n794));
  NOR3_X1   g608(.A1(new_n793), .A2(new_n681), .A3(new_n794), .ZN(new_n795));
  NAND2_X1  g609(.A1(new_n795), .A2(new_n638), .ZN(new_n796));
  AND3_X1   g610(.A1(new_n436), .A2(KEYINPUT38), .A3(new_n437), .ZN(new_n797));
  AOI21_X1  g611(.A(KEYINPUT38), .B1(new_n436), .B2(new_n437), .ZN(new_n798));
  OAI21_X1  g612(.A(new_n440), .B1(new_n797), .B2(new_n798), .ZN(new_n799));
  OAI21_X1  g613(.A(KEYINPUT116), .B1(new_n799), .B2(new_n791), .ZN(new_n800));
  AOI211_X1 g614(.A(new_n599), .B(new_n722), .C1(new_n771), .C2(new_n772), .ZN(new_n801));
  NAND2_X1  g615(.A1(new_n685), .A2(new_n686), .ZN(new_n802));
  INV_X1    g616(.A(new_n791), .ZN(new_n803));
  INV_X1    g617(.A(KEYINPUT116), .ZN(new_n804));
  NAND4_X1  g618(.A1(new_n802), .A2(new_n803), .A3(new_n804), .A4(new_n440), .ZN(new_n805));
  NAND3_X1  g619(.A1(new_n800), .A2(new_n801), .A3(new_n805), .ZN(new_n806));
  INV_X1    g620(.A(KEYINPUT50), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n806), .A2(new_n807), .ZN(new_n808));
  NAND4_X1  g622(.A1(new_n800), .A2(new_n805), .A3(new_n801), .A4(KEYINPUT50), .ZN(new_n809));
  NAND2_X1  g623(.A1(new_n808), .A2(new_n809), .ZN(new_n810));
  AOI21_X1  g624(.A(new_n599), .B1(new_n771), .B2(new_n772), .ZN(new_n811));
  INV_X1    g625(.A(new_n733), .ZN(new_n812));
  NAND3_X1  g626(.A1(new_n792), .A2(new_n811), .A3(new_n812), .ZN(new_n813));
  NAND2_X1  g627(.A1(new_n706), .A2(new_n445), .ZN(new_n814));
  AOI21_X1  g628(.A(new_n779), .B1(new_n786), .B2(new_n814), .ZN(new_n815));
  NOR2_X1   g629(.A1(new_n694), .A2(new_n695), .ZN(new_n816));
  AOI22_X1  g630(.A1(new_n815), .A2(new_n801), .B1(new_n795), .B2(new_n816), .ZN(new_n817));
  NAND3_X1  g631(.A1(new_n810), .A2(new_n813), .A3(new_n817), .ZN(new_n818));
  INV_X1    g632(.A(KEYINPUT51), .ZN(new_n819));
  NAND2_X1  g633(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  NAND4_X1  g634(.A1(new_n810), .A2(new_n817), .A3(KEYINPUT51), .A4(new_n813), .ZN(new_n821));
  NAND2_X1  g635(.A1(new_n801), .A2(new_n716), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n822), .A2(new_n597), .ZN(new_n823));
  NAND4_X1  g637(.A1(new_n792), .A2(new_n811), .A3(new_n316), .A4(new_n362), .ZN(new_n824));
  INV_X1    g638(.A(KEYINPUT48), .ZN(new_n825));
  AND2_X1   g639(.A1(new_n825), .A2(KEYINPUT117), .ZN(new_n826));
  NOR2_X1   g640(.A1(new_n825), .A2(KEYINPUT117), .ZN(new_n827));
  NOR3_X1   g641(.A1(new_n824), .A2(new_n826), .A3(new_n827), .ZN(new_n828));
  AOI211_X1 g642(.A(new_n823), .B(new_n828), .C1(new_n826), .C2(new_n824), .ZN(new_n829));
  AND4_X1   g643(.A1(new_n796), .A2(new_n820), .A3(new_n821), .A4(new_n829), .ZN(new_n830));
  INV_X1    g644(.A(KEYINPUT113), .ZN(new_n831));
  AND4_X1   g645(.A1(new_n441), .A2(new_n436), .A3(new_n437), .A4(new_n484), .ZN(new_n832));
  NOR2_X1   g646(.A1(new_n591), .A2(new_n673), .ZN(new_n833));
  NAND4_X1  g647(.A1(new_n540), .A2(new_n645), .A3(new_n647), .A4(new_n833), .ZN(new_n834));
  NOR2_X1   g648(.A1(new_n834), .A2(new_n665), .ZN(new_n835));
  NAND3_X1  g649(.A1(new_n832), .A2(new_n835), .A3(new_n316), .ZN(new_n836));
  NAND2_X1  g650(.A1(new_n836), .A2(KEYINPUT112), .ZN(new_n837));
  INV_X1    g651(.A(KEYINPUT112), .ZN(new_n838));
  NAND4_X1  g652(.A1(new_n832), .A2(new_n835), .A3(new_n838), .A4(new_n316), .ZN(new_n839));
  AND2_X1   g653(.A1(new_n837), .A2(new_n839), .ZN(new_n840));
  AND4_X1   g654(.A1(KEYINPUT105), .A2(new_n694), .A3(new_n695), .A4(new_n672), .ZN(new_n841));
  AOI21_X1  g655(.A(KEYINPUT105), .B1(new_n638), .B2(new_n672), .ZN(new_n842));
  OAI211_X1 g656(.A(new_n812), .B(new_n832), .C1(new_n841), .C2(new_n842), .ZN(new_n843));
  NAND2_X1  g657(.A1(new_n755), .A2(new_n843), .ZN(new_n844));
  OAI21_X1  g658(.A(new_n831), .B1(new_n840), .B2(new_n844), .ZN(new_n845));
  AOI22_X1  g659(.A1(new_n737), .A2(new_n832), .B1(new_n674), .B2(new_n745), .ZN(new_n846));
  NAND2_X1  g660(.A1(new_n837), .A2(new_n839), .ZN(new_n847));
  NAND3_X1  g661(.A1(new_n846), .A2(KEYINPUT113), .A3(new_n847), .ZN(new_n848));
  NAND2_X1  g662(.A1(new_n845), .A2(new_n848), .ZN(new_n849));
  OAI22_X1  g663(.A1(new_n660), .A2(new_n661), .B1(new_n639), .B2(new_n708), .ZN(new_n850));
  NOR2_X1   g664(.A1(new_n658), .A2(new_n659), .ZN(new_n851));
  NAND4_X1  g665(.A1(new_n626), .A2(new_n316), .A3(new_n362), .A4(new_n484), .ZN(new_n852));
  OAI22_X1  g666(.A1(new_n851), .A2(new_n852), .B1(new_n708), .B2(new_n712), .ZN(new_n853));
  NOR2_X1   g667(.A1(new_n850), .A2(new_n853), .ZN(new_n854));
  AOI21_X1  g668(.A(new_n715), .B1(new_n604), .B2(new_n605), .ZN(new_n855));
  AOI22_X1  g669(.A1(new_n730), .A2(new_n726), .B1(new_n855), .B2(new_n669), .ZN(new_n856));
  INV_X1    g670(.A(KEYINPUT111), .ZN(new_n857));
  NAND3_X1  g671(.A1(new_n540), .A2(new_n552), .A3(new_n591), .ZN(new_n858));
  AOI21_X1  g672(.A(new_n638), .B1(new_n857), .B2(new_n858), .ZN(new_n859));
  OAI21_X1  g673(.A(new_n859), .B1(new_n857), .B2(new_n858), .ZN(new_n860));
  INV_X1    g674(.A(new_n719), .ZN(new_n861));
  NAND4_X1  g675(.A1(new_n860), .A2(new_n362), .A3(new_n623), .A4(new_n861), .ZN(new_n862));
  NAND4_X1  g676(.A1(new_n854), .A2(new_n753), .A3(new_n856), .A4(new_n862), .ZN(new_n863));
  NOR2_X1   g677(.A1(new_n849), .A2(new_n863), .ZN(new_n864));
  INV_X1    g678(.A(KEYINPUT114), .ZN(new_n865));
  INV_X1    g679(.A(KEYINPUT52), .ZN(new_n866));
  OAI21_X1  g680(.A(new_n812), .B1(new_n841), .B2(new_n842), .ZN(new_n867));
  OAI211_X1 g681(.A(new_n675), .B(new_n698), .C1(new_n867), .C2(new_n715), .ZN(new_n868));
  NOR4_X1   g682(.A1(new_n683), .A2(new_n485), .A3(new_n657), .A4(new_n673), .ZN(new_n869));
  OAI211_X1 g683(.A(new_n865), .B(new_n866), .C1(new_n868), .C2(new_n869), .ZN(new_n870));
  OAI21_X1  g684(.A(new_n866), .B1(new_n868), .B2(new_n869), .ZN(new_n871));
  NAND2_X1  g685(.A1(new_n316), .A2(new_n657), .ZN(new_n872));
  NOR2_X1   g686(.A1(new_n872), .A2(new_n485), .ZN(new_n873));
  AOI22_X1  g687(.A1(new_n737), .A2(new_n716), .B1(new_n873), .B2(new_n674), .ZN(new_n874));
  NOR3_X1   g688(.A1(new_n485), .A2(new_n657), .A3(new_n673), .ZN(new_n875));
  NAND3_X1  g689(.A1(new_n875), .A2(new_n681), .A3(new_n682), .ZN(new_n876));
  NAND4_X1  g690(.A1(new_n874), .A2(KEYINPUT52), .A3(new_n698), .A4(new_n876), .ZN(new_n877));
  NAND3_X1  g691(.A1(new_n871), .A2(new_n877), .A3(KEYINPUT114), .ZN(new_n878));
  NAND4_X1  g692(.A1(new_n864), .A2(KEYINPUT53), .A3(new_n870), .A4(new_n878), .ZN(new_n879));
  AND3_X1   g693(.A1(new_n846), .A2(KEYINPUT113), .A3(new_n847), .ZN(new_n880));
  AOI21_X1  g694(.A(KEYINPUT113), .B1(new_n846), .B2(new_n847), .ZN(new_n881));
  NOR2_X1   g695(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  AOI21_X1  g696(.A(new_n665), .B1(new_n604), .B2(new_n605), .ZN(new_n883));
  INV_X1    g697(.A(new_n661), .ZN(new_n884));
  AND4_X1   g698(.A1(new_n316), .A2(new_n362), .A3(new_n704), .A4(new_n707), .ZN(new_n885));
  AOI22_X1  g699(.A1(new_n883), .A2(new_n884), .B1(new_n885), .B2(new_n640), .ZN(new_n886));
  AOI22_X1  g700(.A1(new_n606), .A2(new_n486), .B1(new_n885), .B2(new_n649), .ZN(new_n887));
  NAND3_X1  g701(.A1(new_n886), .A2(new_n887), .A3(new_n862), .ZN(new_n888));
  AND3_X1   g702(.A1(new_n740), .A2(new_n745), .A3(new_n751), .ZN(new_n889));
  AOI21_X1  g703(.A(new_n748), .B1(new_n740), .B2(new_n745), .ZN(new_n890));
  NOR2_X1   g704(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  AOI21_X1  g705(.A(KEYINPUT104), .B1(new_n723), .B2(new_n725), .ZN(new_n892));
  NOR3_X1   g706(.A1(new_n729), .A2(new_n727), .A3(new_n724), .ZN(new_n893));
  OAI21_X1  g707(.A(new_n717), .B1(new_n892), .B2(new_n893), .ZN(new_n894));
  NOR3_X1   g708(.A1(new_n888), .A2(new_n891), .A3(new_n894), .ZN(new_n895));
  NAND2_X1  g709(.A1(new_n871), .A2(new_n877), .ZN(new_n896));
  NAND3_X1  g710(.A1(new_n882), .A2(new_n895), .A3(new_n896), .ZN(new_n897));
  XNOR2_X1  g711(.A(KEYINPUT115), .B(KEYINPUT53), .ZN(new_n898));
  INV_X1    g712(.A(new_n898), .ZN(new_n899));
  NAND2_X1  g713(.A1(new_n897), .A2(new_n899), .ZN(new_n900));
  INV_X1    g714(.A(KEYINPUT54), .ZN(new_n901));
  NAND3_X1  g715(.A1(new_n879), .A2(new_n900), .A3(new_n901), .ZN(new_n902));
  AND3_X1   g716(.A1(new_n882), .A2(new_n895), .A3(new_n896), .ZN(new_n903));
  NAND4_X1  g717(.A1(new_n882), .A2(new_n895), .A3(new_n878), .A4(new_n870), .ZN(new_n904));
  INV_X1    g718(.A(KEYINPUT53), .ZN(new_n905));
  AOI22_X1  g719(.A1(new_n903), .A2(new_n898), .B1(new_n904), .B2(new_n905), .ZN(new_n906));
  OAI211_X1 g720(.A(new_n830), .B(new_n902), .C1(new_n906), .C2(new_n901), .ZN(new_n907));
  NAND2_X1  g721(.A1(new_n596), .A2(new_n277), .ZN(new_n908));
  NAND2_X1  g722(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  NOR3_X1   g723(.A1(new_n694), .A2(new_n445), .A3(new_n637), .ZN(new_n910));
  NAND3_X1  g724(.A1(new_n910), .A2(new_n362), .A3(new_n441), .ZN(new_n911));
  XOR2_X1   g725(.A(new_n911), .B(KEYINPUT109), .Z(new_n912));
  INV_X1    g726(.A(new_n706), .ZN(new_n913));
  NAND2_X1  g727(.A1(new_n913), .A2(KEYINPUT49), .ZN(new_n914));
  AOI21_X1  g728(.A(KEYINPUT110), .B1(new_n912), .B2(new_n914), .ZN(new_n915));
  NOR2_X1   g729(.A1(new_n913), .A2(KEYINPUT49), .ZN(new_n916));
  NOR3_X1   g730(.A1(new_n915), .A2(new_n681), .A3(new_n916), .ZN(new_n917));
  INV_X1    g731(.A(KEYINPUT110), .ZN(new_n918));
  NAND2_X1  g732(.A1(new_n912), .A2(new_n914), .ZN(new_n919));
  OAI211_X1 g733(.A(new_n917), .B(new_n802), .C1(new_n918), .C2(new_n919), .ZN(new_n920));
  NAND2_X1  g734(.A1(new_n909), .A2(new_n920), .ZN(new_n921));
  NAND2_X1  g735(.A1(new_n921), .A2(KEYINPUT118), .ZN(new_n922));
  INV_X1    g736(.A(KEYINPUT118), .ZN(new_n923));
  NAND3_X1  g737(.A1(new_n909), .A2(new_n923), .A3(new_n920), .ZN(new_n924));
  NAND2_X1  g738(.A1(new_n922), .A2(new_n924), .ZN(G75));
  AOI21_X1  g739(.A(new_n347), .B1(new_n879), .B2(new_n900), .ZN(new_n926));
  AOI21_X1  g740(.A(KEYINPUT56), .B1(new_n926), .B2(G210), .ZN(new_n927));
  NAND2_X1  g741(.A1(new_n397), .A2(new_n409), .ZN(new_n928));
  XOR2_X1   g742(.A(new_n928), .B(new_n407), .Z(new_n929));
  XNOR2_X1  g743(.A(new_n929), .B(KEYINPUT55), .ZN(new_n930));
  INV_X1    g744(.A(new_n930), .ZN(new_n931));
  AND2_X1   g745(.A1(new_n927), .A2(new_n931), .ZN(new_n932));
  NOR2_X1   g746(.A1(new_n927), .A2(new_n931), .ZN(new_n933));
  NOR2_X1   g747(.A1(new_n277), .A2(G952), .ZN(new_n934));
  NOR3_X1   g748(.A1(new_n932), .A2(new_n933), .A3(new_n934), .ZN(G51));
  NAND3_X1  g749(.A1(new_n926), .A2(G469), .A3(new_n759), .ZN(new_n936));
  XNOR2_X1  g750(.A(new_n936), .B(KEYINPUT119), .ZN(new_n937));
  AND3_X1   g751(.A1(new_n879), .A2(new_n900), .A3(new_n901), .ZN(new_n938));
  AOI21_X1  g752(.A(new_n901), .B1(new_n879), .B2(new_n900), .ZN(new_n939));
  NOR2_X1   g753(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  XNOR2_X1  g754(.A(new_n764), .B(KEYINPUT57), .ZN(new_n941));
  OAI21_X1  g755(.A(new_n478), .B1(new_n940), .B2(new_n941), .ZN(new_n942));
  AOI21_X1  g756(.A(new_n934), .B1(new_n937), .B2(new_n942), .ZN(G54));
  NAND3_X1  g757(.A1(new_n926), .A2(KEYINPUT58), .A3(G475), .ZN(new_n944));
  INV_X1    g758(.A(new_n549), .ZN(new_n945));
  AND2_X1   g759(.A1(new_n944), .A2(new_n945), .ZN(new_n946));
  NOR2_X1   g760(.A1(new_n944), .A2(new_n945), .ZN(new_n947));
  NOR3_X1   g761(.A1(new_n946), .A2(new_n947), .A3(new_n934), .ZN(G60));
  INV_X1    g762(.A(new_n636), .ZN(new_n949));
  XNOR2_X1  g763(.A(KEYINPUT120), .B(KEYINPUT59), .ZN(new_n950));
  XNOR2_X1  g764(.A(new_n950), .B(new_n627), .ZN(new_n951));
  NOR2_X1   g765(.A1(new_n949), .A2(new_n951), .ZN(new_n952));
  OAI21_X1  g766(.A(new_n952), .B1(new_n938), .B2(new_n939), .ZN(new_n953));
  INV_X1    g767(.A(KEYINPUT121), .ZN(new_n954));
  INV_X1    g768(.A(new_n934), .ZN(new_n955));
  AND3_X1   g769(.A1(new_n953), .A2(new_n954), .A3(new_n955), .ZN(new_n956));
  AOI21_X1  g770(.A(new_n954), .B1(new_n953), .B2(new_n955), .ZN(new_n957));
  OAI21_X1  g771(.A(new_n902), .B1(new_n906), .B2(new_n901), .ZN(new_n958));
  INV_X1    g772(.A(new_n951), .ZN(new_n959));
  AOI21_X1  g773(.A(new_n636), .B1(new_n958), .B2(new_n959), .ZN(new_n960));
  NOR3_X1   g774(.A1(new_n956), .A2(new_n957), .A3(new_n960), .ZN(G63));
  NAND2_X1  g775(.A1(new_n879), .A2(new_n900), .ZN(new_n962));
  NAND2_X1  g776(.A1(G217), .A2(G902), .ZN(new_n963));
  XOR2_X1   g777(.A(new_n963), .B(KEYINPUT122), .Z(new_n964));
  XOR2_X1   g778(.A(new_n964), .B(KEYINPUT60), .Z(new_n965));
  NAND2_X1  g779(.A1(new_n962), .A2(new_n965), .ZN(new_n966));
  INV_X1    g780(.A(new_n358), .ZN(new_n967));
  NAND2_X1  g781(.A1(new_n966), .A2(new_n967), .ZN(new_n968));
  INV_X1    g782(.A(new_n965), .ZN(new_n969));
  AOI21_X1  g783(.A(new_n969), .B1(new_n879), .B2(new_n900), .ZN(new_n970));
  AOI21_X1  g784(.A(new_n934), .B1(new_n970), .B2(new_n655), .ZN(new_n971));
  NAND2_X1  g785(.A1(new_n968), .A2(new_n971), .ZN(new_n972));
  INV_X1    g786(.A(KEYINPUT123), .ZN(new_n973));
  INV_X1    g787(.A(new_n655), .ZN(new_n974));
  OAI211_X1 g788(.A(new_n973), .B(new_n955), .C1(new_n966), .C2(new_n974), .ZN(new_n975));
  NAND3_X1  g789(.A1(new_n972), .A2(KEYINPUT61), .A3(new_n975), .ZN(new_n976));
  INV_X1    g790(.A(KEYINPUT61), .ZN(new_n977));
  OAI211_X1 g791(.A(new_n968), .B(new_n971), .C1(new_n973), .C2(new_n977), .ZN(new_n978));
  AND2_X1   g792(.A1(new_n976), .A2(new_n978), .ZN(G66));
  AOI21_X1  g793(.A(new_n277), .B1(new_n600), .B2(G224), .ZN(new_n980));
  NAND3_X1  g794(.A1(new_n854), .A2(new_n856), .A3(new_n862), .ZN(new_n981));
  AOI21_X1  g795(.A(new_n980), .B1(new_n981), .B2(new_n277), .ZN(new_n982));
  OAI21_X1  g796(.A(new_n928), .B1(G898), .B2(new_n277), .ZN(new_n983));
  XOR2_X1   g797(.A(new_n982), .B(new_n983), .Z(G69));
  NOR2_X1   g798(.A1(new_n692), .A2(new_n868), .ZN(new_n985));
  XNOR2_X1  g799(.A(new_n985), .B(KEYINPUT62), .ZN(new_n986));
  AOI21_X1  g800(.A(new_n788), .B1(new_n777), .B2(new_n780), .ZN(new_n987));
  OR2_X1    g801(.A1(new_n860), .A2(KEYINPUT124), .ZN(new_n988));
  NAND2_X1  g802(.A1(new_n860), .A2(KEYINPUT124), .ZN(new_n989));
  NAND4_X1  g803(.A1(new_n988), .A2(new_n689), .A3(new_n745), .A4(new_n989), .ZN(new_n990));
  NAND3_X1  g804(.A1(new_n986), .A2(new_n987), .A3(new_n990), .ZN(new_n991));
  NAND2_X1  g805(.A1(new_n991), .A2(new_n277), .ZN(new_n992));
  INV_X1    g806(.A(new_n992), .ZN(new_n993));
  NAND2_X1  g807(.A1(new_n285), .A2(new_n286), .ZN(new_n994));
  XOR2_X1   g808(.A(new_n994), .B(new_n543), .Z(new_n995));
  INV_X1    g809(.A(new_n995), .ZN(new_n996));
  OAI21_X1  g810(.A(KEYINPUT125), .B1(new_n993), .B2(new_n996), .ZN(new_n997));
  NAND2_X1  g811(.A1(G900), .A2(G953), .ZN(new_n998));
  NAND2_X1  g812(.A1(new_n753), .A2(new_n755), .ZN(new_n999));
  XNOR2_X1  g813(.A(new_n999), .B(KEYINPUT126), .ZN(new_n1000));
  INV_X1    g814(.A(new_n626), .ZN(new_n1001));
  NOR3_X1   g815(.A1(new_n769), .A2(new_n363), .A3(new_n1001), .ZN(new_n1002));
  AOI21_X1  g816(.A(new_n868), .B1(new_n1002), .B2(new_n682), .ZN(new_n1003));
  NAND3_X1  g817(.A1(new_n1000), .A2(new_n1003), .A3(new_n987), .ZN(new_n1004));
  OAI211_X1 g818(.A(new_n998), .B(new_n996), .C1(new_n1004), .C2(G953), .ZN(new_n1005));
  INV_X1    g819(.A(KEYINPUT125), .ZN(new_n1006));
  NAND3_X1  g820(.A1(new_n992), .A2(new_n1006), .A3(new_n995), .ZN(new_n1007));
  NAND3_X1  g821(.A1(new_n997), .A2(new_n1005), .A3(new_n1007), .ZN(new_n1008));
  AOI21_X1  g822(.A(new_n277), .B1(G227), .B2(G900), .ZN(new_n1009));
  NAND2_X1  g823(.A1(new_n1008), .A2(new_n1009), .ZN(new_n1010));
  INV_X1    g824(.A(new_n1009), .ZN(new_n1011));
  NAND4_X1  g825(.A1(new_n997), .A2(new_n1005), .A3(new_n1011), .A4(new_n1007), .ZN(new_n1012));
  NAND2_X1  g826(.A1(new_n1010), .A2(new_n1012), .ZN(G72));
  NAND2_X1  g827(.A1(G472), .A2(G902), .ZN(new_n1014));
  XOR2_X1   g828(.A(new_n1014), .B(KEYINPUT63), .Z(new_n1015));
  OAI21_X1  g829(.A(new_n1015), .B1(new_n991), .B2(new_n981), .ZN(new_n1016));
  NAND2_X1  g830(.A1(new_n1016), .A2(KEYINPUT127), .ZN(new_n1017));
  INV_X1    g831(.A(KEYINPUT127), .ZN(new_n1018));
  OAI211_X1 g832(.A(new_n1018), .B(new_n1015), .C1(new_n991), .C2(new_n981), .ZN(new_n1019));
  NAND3_X1  g833(.A1(new_n1017), .A2(new_n679), .A3(new_n1019), .ZN(new_n1020));
  OAI21_X1  g834(.A(new_n1015), .B1(new_n1004), .B2(new_n981), .ZN(new_n1021));
  NOR2_X1   g835(.A1(new_n310), .A2(new_n290), .ZN(new_n1022));
  NAND2_X1  g836(.A1(new_n1021), .A2(new_n1022), .ZN(new_n1023));
  NAND3_X1  g837(.A1(new_n1020), .A2(new_n1023), .A3(new_n955), .ZN(new_n1024));
  OAI21_X1  g838(.A(new_n1015), .B1(new_n310), .B2(new_n290), .ZN(new_n1025));
  NOR3_X1   g839(.A1(new_n906), .A2(new_n679), .A3(new_n1025), .ZN(new_n1026));
  NOR2_X1   g840(.A1(new_n1024), .A2(new_n1026), .ZN(G57));
endmodule


