//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 1 1 1 1 1 1 1 1 1 0 1 0 0 1 0 0 0 0 0 0 1 0 1 0 1 0 1 1 0 1 0 0 1 0 1 1 1 1 1 1 1 1 1 0 0 1 1 0 1 1 0 1 0 1 1 1 1 1 1 0 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:37:26 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n236, new_n237,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n244, new_n245,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n252, new_n253,
    new_n254, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1188, new_n1189, new_n1190, new_n1191, new_n1192, new_n1193,
    new_n1194, new_n1195, new_n1196, new_n1197, new_n1198, new_n1199,
    new_n1200, new_n1201, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1216, new_n1217, new_n1218, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1288, new_n1289, new_n1290, new_n1291;
  INV_X1    g0000(.A(G58), .ZN(new_n201));
  INV_X1    g0001(.A(G68), .ZN(new_n202));
  NAND3_X1  g0002(.A1(new_n201), .A2(new_n202), .A3(KEYINPUT64), .ZN(new_n203));
  INV_X1    g0003(.A(KEYINPUT64), .ZN(new_n204));
  OAI21_X1  g0004(.A(new_n204), .B1(G58), .B2(G68), .ZN(new_n205));
  AND2_X1   g0005(.A1(new_n203), .A2(new_n205), .ZN(new_n206));
  NOR3_X1   g0006(.A1(new_n206), .A2(G50), .A3(G77), .ZN(G353));
  OAI21_X1  g0007(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0008(.A(G1), .ZN(new_n209));
  INV_X1    g0009(.A(G20), .ZN(new_n210));
  NOR2_X1   g0010(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  INV_X1    g0011(.A(new_n211), .ZN(new_n212));
  NOR2_X1   g0012(.A1(new_n212), .A2(G13), .ZN(new_n213));
  OAI211_X1 g0013(.A(new_n213), .B(G250), .C1(G257), .C2(G264), .ZN(new_n214));
  XNOR2_X1  g0014(.A(new_n214), .B(KEYINPUT0), .ZN(new_n215));
  NAND2_X1  g0015(.A1(new_n206), .A2(G50), .ZN(new_n216));
  INV_X1    g0016(.A(new_n216), .ZN(new_n217));
  NAND2_X1  g0017(.A1(G1), .A2(G13), .ZN(new_n218));
  NOR2_X1   g0018(.A1(new_n218), .A2(new_n210), .ZN(new_n219));
  NAND2_X1  g0019(.A1(new_n217), .A2(new_n219), .ZN(new_n220));
  AOI22_X1  g0020(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n221));
  INV_X1    g0021(.A(G232), .ZN(new_n222));
  INV_X1    g0022(.A(G107), .ZN(new_n223));
  INV_X1    g0023(.A(G264), .ZN(new_n224));
  OAI221_X1 g0024(.A(new_n221), .B1(new_n201), .B2(new_n222), .C1(new_n223), .C2(new_n224), .ZN(new_n225));
  NAND2_X1  g0025(.A1(new_n225), .A2(KEYINPUT66), .ZN(new_n226));
  NAND2_X1  g0026(.A1(G116), .A2(G270), .ZN(new_n227));
  INV_X1    g0027(.A(G50), .ZN(new_n228));
  INV_X1    g0028(.A(G226), .ZN(new_n229));
  OAI21_X1  g0029(.A(new_n227), .B1(new_n228), .B2(new_n229), .ZN(new_n230));
  AOI21_X1  g0030(.A(new_n230), .B1(G68), .B2(G238), .ZN(new_n231));
  INV_X1    g0031(.A(G244), .ZN(new_n232));
  XNOR2_X1  g0032(.A(KEYINPUT65), .B(G77), .ZN(new_n233));
  OAI211_X1 g0033(.A(new_n226), .B(new_n231), .C1(new_n232), .C2(new_n233), .ZN(new_n234));
  NOR2_X1   g0034(.A1(new_n225), .A2(KEYINPUT66), .ZN(new_n235));
  OAI21_X1  g0035(.A(new_n212), .B1(new_n234), .B2(new_n235), .ZN(new_n236));
  OAI211_X1 g0036(.A(new_n215), .B(new_n220), .C1(new_n236), .C2(KEYINPUT1), .ZN(new_n237));
  AOI21_X1  g0037(.A(new_n237), .B1(KEYINPUT1), .B2(new_n236), .ZN(G361));
  XNOR2_X1  g0038(.A(G238), .B(G244), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n239), .B(G232), .ZN(new_n240));
  XNOR2_X1  g0040(.A(KEYINPUT2), .B(G226), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XNOR2_X1  g0042(.A(G250), .B(G257), .ZN(new_n243));
  XNOR2_X1  g0043(.A(G264), .B(G270), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XOR2_X1   g0045(.A(new_n242), .B(new_n245), .Z(G358));
  XOR2_X1   g0046(.A(G87), .B(G97), .Z(new_n247));
  XNOR2_X1  g0047(.A(G107), .B(G116), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n247), .B(new_n248), .ZN(new_n249));
  NAND2_X1  g0049(.A1(new_n228), .A2(G68), .ZN(new_n250));
  NAND2_X1  g0050(.A1(new_n202), .A2(G50), .ZN(new_n251));
  NAND2_X1  g0051(.A1(new_n250), .A2(new_n251), .ZN(new_n252));
  XNOR2_X1  g0052(.A(G58), .B(G77), .ZN(new_n253));
  XNOR2_X1  g0053(.A(new_n252), .B(new_n253), .ZN(new_n254));
  XNOR2_X1  g0054(.A(new_n249), .B(new_n254), .ZN(G351));
  NAND3_X1  g0055(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n256), .A2(new_n218), .ZN(new_n257));
  XOR2_X1   g0057(.A(KEYINPUT70), .B(G107), .Z(new_n258));
  INV_X1    g0058(.A(G33), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n259), .A2(KEYINPUT3), .ZN(new_n260));
  INV_X1    g0060(.A(KEYINPUT3), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n261), .A2(G33), .ZN(new_n262));
  INV_X1    g0062(.A(KEYINPUT75), .ZN(new_n263));
  NAND3_X1  g0063(.A1(new_n260), .A2(new_n262), .A3(new_n263), .ZN(new_n264));
  INV_X1    g0064(.A(KEYINPUT7), .ZN(new_n265));
  NOR2_X1   g0065(.A1(new_n265), .A2(G20), .ZN(new_n266));
  NAND3_X1  g0066(.A1(new_n261), .A2(KEYINPUT75), .A3(G33), .ZN(new_n267));
  NAND3_X1  g0067(.A1(new_n264), .A2(new_n266), .A3(new_n267), .ZN(new_n268));
  XNOR2_X1  g0068(.A(KEYINPUT3), .B(G33), .ZN(new_n269));
  OAI21_X1  g0069(.A(new_n265), .B1(new_n269), .B2(G20), .ZN(new_n270));
  AOI21_X1  g0070(.A(new_n258), .B1(new_n268), .B2(new_n270), .ZN(new_n271));
  NOR2_X1   g0071(.A1(G20), .A2(G33), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n272), .A2(G77), .ZN(new_n273));
  NAND2_X1  g0073(.A1(KEYINPUT6), .A2(G97), .ZN(new_n274));
  NOR2_X1   g0074(.A1(new_n274), .A2(G107), .ZN(new_n275));
  XNOR2_X1  g0075(.A(G97), .B(G107), .ZN(new_n276));
  INV_X1    g0076(.A(KEYINPUT6), .ZN(new_n277));
  AOI21_X1  g0077(.A(new_n275), .B1(new_n276), .B2(new_n277), .ZN(new_n278));
  OAI21_X1  g0078(.A(new_n273), .B1(new_n278), .B2(new_n210), .ZN(new_n279));
  OAI21_X1  g0079(.A(new_n257), .B1(new_n271), .B2(new_n279), .ZN(new_n280));
  INV_X1    g0080(.A(G13), .ZN(new_n281));
  NOR3_X1   g0081(.A1(new_n281), .A2(new_n210), .A3(G1), .ZN(new_n282));
  INV_X1    g0082(.A(new_n282), .ZN(new_n283));
  NOR2_X1   g0083(.A1(new_n283), .A2(G97), .ZN(new_n284));
  AOI211_X1 g0084(.A(new_n257), .B(new_n282), .C1(new_n209), .C2(G33), .ZN(new_n285));
  AOI21_X1  g0085(.A(new_n284), .B1(new_n285), .B2(G97), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n280), .A2(new_n286), .ZN(new_n287));
  NOR2_X1   g0087(.A1(new_n232), .A2(G1698), .ZN(new_n288));
  NAND3_X1  g0088(.A1(new_n288), .A2(new_n260), .A3(new_n262), .ZN(new_n289));
  INV_X1    g0089(.A(KEYINPUT4), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  NAND3_X1  g0091(.A1(new_n269), .A2(G250), .A3(G1698), .ZN(new_n292));
  NAND3_X1  g0092(.A1(new_n269), .A2(KEYINPUT4), .A3(new_n288), .ZN(new_n293));
  NAND2_X1  g0093(.A1(G33), .A2(G283), .ZN(new_n294));
  NAND4_X1  g0094(.A1(new_n291), .A2(new_n292), .A3(new_n293), .A4(new_n294), .ZN(new_n295));
  INV_X1    g0095(.A(new_n218), .ZN(new_n296));
  NAND2_X1  g0096(.A1(G33), .A2(G41), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n296), .A2(new_n297), .ZN(new_n298));
  INV_X1    g0098(.A(new_n298), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n295), .A2(new_n299), .ZN(new_n300));
  INV_X1    g0100(.A(G179), .ZN(new_n301));
  INV_X1    g0101(.A(G41), .ZN(new_n302));
  OAI211_X1 g0102(.A(new_n209), .B(G45), .C1(new_n302), .C2(KEYINPUT5), .ZN(new_n303));
  INV_X1    g0103(.A(KEYINPUT5), .ZN(new_n304));
  NOR2_X1   g0104(.A1(new_n304), .A2(G41), .ZN(new_n305));
  OR2_X1    g0105(.A1(new_n303), .A2(new_n305), .ZN(new_n306));
  INV_X1    g0106(.A(KEYINPUT68), .ZN(new_n307));
  INV_X1    g0107(.A(KEYINPUT67), .ZN(new_n308));
  AOI21_X1  g0108(.A(new_n218), .B1(new_n308), .B2(new_n297), .ZN(new_n309));
  NAND3_X1  g0109(.A1(KEYINPUT67), .A2(G33), .A3(G41), .ZN(new_n310));
  AOI21_X1  g0110(.A(new_n307), .B1(new_n309), .B2(new_n310), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n297), .A2(new_n308), .ZN(new_n312));
  AND4_X1   g0112(.A1(new_n307), .A2(new_n312), .A3(new_n296), .A4(new_n310), .ZN(new_n313));
  OAI211_X1 g0113(.A(new_n306), .B(G257), .C1(new_n311), .C2(new_n313), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n304), .A2(G41), .ZN(new_n315));
  NAND4_X1  g0115(.A1(new_n315), .A2(KEYINPUT80), .A3(new_n209), .A4(G45), .ZN(new_n316));
  OAI21_X1  g0116(.A(G274), .B1(new_n304), .B2(G41), .ZN(new_n317));
  INV_X1    g0117(.A(KEYINPUT80), .ZN(new_n318));
  AOI21_X1  g0118(.A(new_n317), .B1(new_n303), .B2(new_n318), .ZN(new_n319));
  OAI211_X1 g0119(.A(new_n316), .B(new_n319), .C1(new_n311), .C2(new_n313), .ZN(new_n320));
  NAND4_X1  g0120(.A1(new_n300), .A2(new_n301), .A3(new_n314), .A4(new_n320), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n287), .A2(new_n321), .ZN(new_n322));
  AND2_X1   g0122(.A1(new_n319), .A2(new_n316), .ZN(new_n323));
  NAND3_X1  g0123(.A1(new_n312), .A2(new_n296), .A3(new_n310), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n324), .A2(KEYINPUT68), .ZN(new_n325));
  NAND3_X1  g0125(.A1(new_n309), .A2(new_n307), .A3(new_n310), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  AOI22_X1  g0127(.A1(new_n295), .A2(new_n299), .B1(new_n323), .B2(new_n327), .ZN(new_n328));
  AOI21_X1  g0128(.A(G169), .B1(new_n328), .B2(new_n314), .ZN(new_n329));
  OAI21_X1  g0129(.A(KEYINPUT81), .B1(new_n322), .B2(new_n329), .ZN(new_n330));
  NAND3_X1  g0130(.A1(new_n300), .A2(new_n314), .A3(new_n320), .ZN(new_n331));
  INV_X1    g0131(.A(G169), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n331), .A2(new_n332), .ZN(new_n333));
  INV_X1    g0133(.A(KEYINPUT81), .ZN(new_n334));
  NAND4_X1  g0134(.A1(new_n333), .A2(new_n334), .A3(new_n287), .A4(new_n321), .ZN(new_n335));
  AND2_X1   g0135(.A1(new_n280), .A2(new_n286), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n331), .A2(G200), .ZN(new_n337));
  INV_X1    g0137(.A(G190), .ZN(new_n338));
  OAI211_X1 g0138(.A(new_n336), .B(new_n337), .C1(new_n338), .C2(new_n331), .ZN(new_n339));
  NAND3_X1  g0139(.A1(new_n330), .A2(new_n335), .A3(new_n339), .ZN(new_n340));
  INV_X1    g0140(.A(KEYINPUT82), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n340), .A2(new_n341), .ZN(new_n342));
  INV_X1    g0142(.A(G97), .ZN(new_n343));
  NOR2_X1   g0143(.A1(new_n259), .A2(new_n343), .ZN(new_n344));
  AOI21_X1  g0144(.A(G20), .B1(new_n344), .B2(KEYINPUT19), .ZN(new_n345));
  INV_X1    g0145(.A(KEYINPUT83), .ZN(new_n346));
  INV_X1    g0146(.A(new_n258), .ZN(new_n347));
  INV_X1    g0147(.A(G87), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n348), .A2(new_n343), .ZN(new_n349));
  OAI21_X1  g0149(.A(new_n346), .B1(new_n347), .B2(new_n349), .ZN(new_n350));
  NAND4_X1  g0150(.A1(new_n258), .A2(KEYINPUT83), .A3(new_n348), .A4(new_n343), .ZN(new_n351));
  AOI21_X1  g0151(.A(new_n345), .B1(new_n350), .B2(new_n351), .ZN(new_n352));
  NAND3_X1  g0152(.A1(new_n269), .A2(new_n210), .A3(G68), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n210), .A2(G33), .ZN(new_n354));
  NOR2_X1   g0154(.A1(new_n354), .A2(new_n343), .ZN(new_n355));
  OAI21_X1  g0155(.A(new_n353), .B1(KEYINPUT19), .B2(new_n355), .ZN(new_n356));
  OAI21_X1  g0156(.A(new_n257), .B1(new_n352), .B2(new_n356), .ZN(new_n357));
  XNOR2_X1  g0157(.A(KEYINPUT15), .B(G87), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n358), .A2(new_n282), .ZN(new_n359));
  INV_X1    g0159(.A(new_n358), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n285), .A2(new_n360), .ZN(new_n361));
  AND3_X1   g0161(.A1(new_n357), .A2(new_n359), .A3(new_n361), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n209), .A2(G45), .ZN(new_n363));
  NOR2_X1   g0163(.A1(new_n363), .A2(G274), .ZN(new_n364));
  INV_X1    g0164(.A(G250), .ZN(new_n365));
  AOI21_X1  g0165(.A(new_n364), .B1(new_n365), .B2(new_n363), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n327), .A2(new_n366), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n232), .A2(G1698), .ZN(new_n368));
  OAI21_X1  g0168(.A(new_n368), .B1(G238), .B2(G1698), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n260), .A2(new_n262), .ZN(new_n370));
  INV_X1    g0170(.A(G116), .ZN(new_n371));
  OAI22_X1  g0171(.A1(new_n369), .A2(new_n370), .B1(new_n259), .B2(new_n371), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n372), .A2(new_n299), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n367), .A2(new_n373), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n374), .A2(new_n332), .ZN(new_n375));
  OAI21_X1  g0175(.A(new_n375), .B1(G179), .B2(new_n374), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n374), .A2(G200), .ZN(new_n377));
  OAI21_X1  g0177(.A(new_n377), .B1(new_n338), .B2(new_n374), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n285), .A2(G87), .ZN(new_n379));
  NAND3_X1  g0179(.A1(new_n357), .A2(new_n359), .A3(new_n379), .ZN(new_n380));
  OAI22_X1  g0180(.A1(new_n362), .A2(new_n376), .B1(new_n378), .B2(new_n380), .ZN(new_n381));
  INV_X1    g0181(.A(new_n381), .ZN(new_n382));
  NAND4_X1  g0182(.A1(new_n330), .A2(new_n339), .A3(KEYINPUT82), .A4(new_n335), .ZN(new_n383));
  NAND3_X1  g0183(.A1(new_n342), .A2(new_n382), .A3(new_n383), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n384), .A2(KEYINPUT84), .ZN(new_n385));
  AOI21_X1  g0185(.A(new_n381), .B1(new_n340), .B2(new_n341), .ZN(new_n386));
  INV_X1    g0186(.A(KEYINPUT84), .ZN(new_n387));
  NAND3_X1  g0187(.A1(new_n386), .A2(new_n387), .A3(new_n383), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n385), .A2(new_n388), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n269), .A2(G1698), .ZN(new_n390));
  XNOR2_X1  g0190(.A(new_n390), .B(KEYINPUT69), .ZN(new_n391));
  INV_X1    g0191(.A(G223), .ZN(new_n392));
  NOR2_X1   g0192(.A1(new_n391), .A2(new_n392), .ZN(new_n393));
  INV_X1    g0193(.A(G1698), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n269), .A2(new_n394), .ZN(new_n395));
  INV_X1    g0195(.A(G222), .ZN(new_n396));
  OAI22_X1  g0196(.A1(new_n395), .A2(new_n396), .B1(new_n233), .B2(new_n269), .ZN(new_n397));
  OAI21_X1  g0197(.A(new_n299), .B1(new_n393), .B2(new_n397), .ZN(new_n398));
  INV_X1    g0198(.A(G45), .ZN(new_n399));
  AOI21_X1  g0199(.A(G1), .B1(new_n302), .B2(new_n399), .ZN(new_n400));
  NAND3_X1  g0200(.A1(new_n327), .A2(G274), .A3(new_n400), .ZN(new_n401));
  OAI21_X1  g0201(.A(new_n209), .B1(G41), .B2(G45), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n327), .A2(new_n402), .ZN(new_n403));
  INV_X1    g0203(.A(new_n403), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n404), .A2(G226), .ZN(new_n405));
  AND3_X1   g0205(.A1(new_n398), .A2(new_n401), .A3(new_n405), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n406), .A2(G190), .ZN(new_n407));
  OAI21_X1  g0207(.A(G20), .B1(new_n206), .B2(G50), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n272), .A2(G150), .ZN(new_n409));
  XNOR2_X1  g0209(.A(KEYINPUT8), .B(G58), .ZN(new_n410));
  OAI211_X1 g0210(.A(new_n408), .B(new_n409), .C1(new_n354), .C2(new_n410), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n411), .A2(new_n257), .ZN(new_n412));
  NOR2_X1   g0212(.A1(new_n282), .A2(new_n257), .ZN(new_n413));
  AOI21_X1  g0213(.A(new_n228), .B1(new_n209), .B2(G20), .ZN(new_n414));
  AOI22_X1  g0214(.A1(new_n413), .A2(new_n414), .B1(new_n228), .B2(new_n282), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n412), .A2(new_n415), .ZN(new_n416));
  XNOR2_X1  g0216(.A(new_n416), .B(KEYINPUT9), .ZN(new_n417));
  NAND3_X1  g0217(.A1(new_n398), .A2(new_n401), .A3(new_n405), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n418), .A2(G200), .ZN(new_n419));
  NAND3_X1  g0219(.A1(new_n407), .A2(new_n417), .A3(new_n419), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n420), .A2(KEYINPUT10), .ZN(new_n421));
  INV_X1    g0221(.A(KEYINPUT10), .ZN(new_n422));
  NAND4_X1  g0222(.A1(new_n407), .A2(new_n417), .A3(new_n422), .A4(new_n419), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n421), .A2(new_n423), .ZN(new_n424));
  INV_X1    g0224(.A(new_n424), .ZN(new_n425));
  INV_X1    g0225(.A(new_n272), .ZN(new_n426));
  AOI21_X1  g0226(.A(new_n410), .B1(KEYINPUT72), .B2(new_n426), .ZN(new_n427));
  OAI21_X1  g0227(.A(new_n427), .B1(KEYINPUT72), .B2(new_n426), .ZN(new_n428));
  OAI221_X1 g0228(.A(new_n428), .B1(new_n210), .B2(new_n233), .C1(new_n354), .C2(new_n358), .ZN(new_n429));
  AND2_X1   g0229(.A1(new_n429), .A2(new_n257), .ZN(new_n430));
  INV_X1    g0230(.A(new_n413), .ZN(new_n431));
  OAI21_X1  g0231(.A(G77), .B1(new_n210), .B2(G1), .ZN(new_n432));
  INV_X1    g0232(.A(new_n233), .ZN(new_n433));
  OAI22_X1  g0233(.A1(new_n431), .A2(new_n432), .B1(new_n433), .B2(new_n283), .ZN(new_n434));
  NOR2_X1   g0234(.A1(new_n430), .A2(new_n434), .ZN(new_n435));
  INV_X1    g0235(.A(KEYINPUT71), .ZN(new_n436));
  INV_X1    g0236(.A(G238), .ZN(new_n437));
  OR2_X1    g0237(.A1(new_n391), .A2(new_n437), .ZN(new_n438));
  OAI22_X1  g0238(.A1(new_n395), .A2(new_n222), .B1(new_n258), .B2(new_n269), .ZN(new_n439));
  INV_X1    g0239(.A(new_n439), .ZN(new_n440));
  AOI21_X1  g0240(.A(new_n298), .B1(new_n438), .B2(new_n440), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n404), .A2(G244), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n442), .A2(new_n401), .ZN(new_n443));
  OAI21_X1  g0243(.A(new_n436), .B1(new_n441), .B2(new_n443), .ZN(new_n444));
  AND2_X1   g0244(.A1(new_n442), .A2(new_n401), .ZN(new_n445));
  NOR2_X1   g0245(.A1(new_n391), .A2(new_n437), .ZN(new_n446));
  OAI21_X1  g0246(.A(new_n299), .B1(new_n446), .B2(new_n439), .ZN(new_n447));
  NAND3_X1  g0247(.A1(new_n445), .A2(KEYINPUT71), .A3(new_n447), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n444), .A2(new_n448), .ZN(new_n449));
  AOI21_X1  g0249(.A(new_n435), .B1(new_n449), .B2(new_n301), .ZN(new_n450));
  NAND3_X1  g0250(.A1(new_n444), .A2(new_n448), .A3(new_n332), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  INV_X1    g0252(.A(new_n452), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n406), .A2(new_n301), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n418), .A2(new_n332), .ZN(new_n455));
  NAND3_X1  g0255(.A1(new_n454), .A2(new_n416), .A3(new_n455), .ZN(new_n456));
  INV_X1    g0256(.A(new_n456), .ZN(new_n457));
  INV_X1    g0257(.A(G200), .ZN(new_n458));
  OAI21_X1  g0258(.A(new_n435), .B1(new_n449), .B2(new_n458), .ZN(new_n459));
  AOI21_X1  g0259(.A(new_n338), .B1(new_n444), .B2(new_n448), .ZN(new_n460));
  NOR2_X1   g0260(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  OR4_X1    g0261(.A1(new_n425), .A2(new_n453), .A3(new_n457), .A4(new_n461), .ZN(new_n462));
  AOI21_X1  g0262(.A(new_n410), .B1(new_n209), .B2(G20), .ZN(new_n463));
  AOI22_X1  g0263(.A1(new_n463), .A2(new_n413), .B1(new_n282), .B2(new_n410), .ZN(new_n464));
  AOI21_X1  g0264(.A(KEYINPUT7), .B1(new_n370), .B2(new_n210), .ZN(new_n465));
  INV_X1    g0265(.A(new_n266), .ZN(new_n466));
  NOR2_X1   g0266(.A1(new_n269), .A2(new_n466), .ZN(new_n467));
  OAI21_X1  g0267(.A(G68), .B1(new_n465), .B2(new_n467), .ZN(new_n468));
  NAND2_X1  g0268(.A1(G58), .A2(G68), .ZN(new_n469));
  NAND3_X1  g0269(.A1(new_n203), .A2(new_n205), .A3(new_n469), .ZN(new_n470));
  AOI22_X1  g0270(.A1(new_n470), .A2(G20), .B1(G159), .B2(new_n272), .ZN(new_n471));
  NAND3_X1  g0271(.A1(new_n468), .A2(KEYINPUT16), .A3(new_n471), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n472), .A2(new_n257), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n268), .A2(new_n270), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n474), .A2(G68), .ZN(new_n475));
  AOI21_X1  g0275(.A(KEYINPUT16), .B1(new_n475), .B2(new_n471), .ZN(new_n476));
  OAI21_X1  g0276(.A(new_n464), .B1(new_n473), .B2(new_n476), .ZN(new_n477));
  INV_X1    g0277(.A(KEYINPUT76), .ZN(new_n478));
  NOR2_X1   g0278(.A1(new_n259), .A2(new_n348), .ZN(new_n479));
  NOR2_X1   g0279(.A1(G223), .A2(G1698), .ZN(new_n480));
  AOI21_X1  g0280(.A(new_n480), .B1(new_n229), .B2(G1698), .ZN(new_n481));
  AOI21_X1  g0281(.A(new_n479), .B1(new_n481), .B2(new_n269), .ZN(new_n482));
  OAI21_X1  g0282(.A(new_n478), .B1(new_n482), .B2(new_n298), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n392), .A2(new_n394), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n229), .A2(G1698), .ZN(new_n485));
  NAND4_X1  g0285(.A1(new_n260), .A2(new_n484), .A3(new_n262), .A4(new_n485), .ZN(new_n486));
  INV_X1    g0286(.A(new_n479), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n486), .A2(new_n487), .ZN(new_n488));
  NAND3_X1  g0288(.A1(new_n488), .A2(KEYINPUT76), .A3(new_n299), .ZN(new_n489));
  AND2_X1   g0289(.A1(new_n483), .A2(new_n489), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n400), .A2(G274), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n402), .A2(G232), .ZN(new_n492));
  AOI22_X1  g0292(.A1(new_n325), .A2(new_n326), .B1(new_n491), .B2(new_n492), .ZN(new_n493));
  NOR2_X1   g0293(.A1(new_n493), .A2(G179), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n491), .A2(new_n492), .ZN(new_n495));
  OAI21_X1  g0295(.A(new_n495), .B1(new_n311), .B2(new_n313), .ZN(new_n496));
  AOI21_X1  g0296(.A(new_n298), .B1(new_n486), .B2(new_n487), .ZN(new_n497));
  INV_X1    g0297(.A(new_n497), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n496), .A2(new_n498), .ZN(new_n499));
  AOI22_X1  g0299(.A1(new_n490), .A2(new_n494), .B1(new_n332), .B2(new_n499), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n477), .A2(new_n500), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n501), .A2(KEYINPUT18), .ZN(new_n502));
  INV_X1    g0302(.A(KEYINPUT18), .ZN(new_n503));
  NAND3_X1  g0303(.A1(new_n477), .A2(new_n500), .A3(new_n503), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n502), .A2(new_n504), .ZN(new_n505));
  NAND4_X1  g0305(.A1(new_n483), .A2(new_n496), .A3(new_n338), .A4(new_n489), .ZN(new_n506));
  OAI21_X1  g0306(.A(new_n458), .B1(new_n493), .B2(new_n497), .ZN(new_n507));
  AND3_X1   g0307(.A1(new_n506), .A2(KEYINPUT77), .A3(new_n507), .ZN(new_n508));
  AOI21_X1  g0308(.A(KEYINPUT77), .B1(new_n506), .B2(new_n507), .ZN(new_n509));
  NOR2_X1   g0309(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  OAI21_X1  g0310(.A(KEYINPUT78), .B1(new_n510), .B2(new_n477), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n506), .A2(new_n507), .ZN(new_n512));
  INV_X1    g0312(.A(KEYINPUT77), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  NAND3_X1  g0314(.A1(new_n506), .A2(KEYINPUT77), .A3(new_n507), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  INV_X1    g0316(.A(KEYINPUT78), .ZN(new_n517));
  INV_X1    g0317(.A(new_n464), .ZN(new_n518));
  INV_X1    g0318(.A(new_n257), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n370), .A2(new_n266), .ZN(new_n520));
  AOI21_X1  g0320(.A(new_n202), .B1(new_n270), .B2(new_n520), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n470), .A2(G20), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n272), .A2(G159), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  NOR2_X1   g0324(.A1(new_n521), .A2(new_n524), .ZN(new_n525));
  AOI21_X1  g0325(.A(new_n519), .B1(new_n525), .B2(KEYINPUT16), .ZN(new_n526));
  INV_X1    g0326(.A(KEYINPUT16), .ZN(new_n527));
  AOI21_X1  g0327(.A(new_n202), .B1(new_n268), .B2(new_n270), .ZN(new_n528));
  OAI21_X1  g0328(.A(new_n527), .B1(new_n528), .B2(new_n524), .ZN(new_n529));
  AOI21_X1  g0329(.A(new_n518), .B1(new_n526), .B2(new_n529), .ZN(new_n530));
  NAND4_X1  g0330(.A1(new_n516), .A2(new_n517), .A3(KEYINPUT79), .A4(new_n530), .ZN(new_n531));
  NAND3_X1  g0331(.A1(new_n511), .A2(new_n531), .A3(KEYINPUT17), .ZN(new_n532));
  INV_X1    g0332(.A(KEYINPUT17), .ZN(new_n533));
  NAND4_X1  g0333(.A1(new_n516), .A2(KEYINPUT79), .A3(new_n533), .A4(new_n530), .ZN(new_n534));
  AOI21_X1  g0334(.A(new_n505), .B1(new_n532), .B2(new_n534), .ZN(new_n535));
  INV_X1    g0335(.A(new_n535), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n222), .A2(G1698), .ZN(new_n537));
  OAI21_X1  g0337(.A(new_n537), .B1(G226), .B2(G1698), .ZN(new_n538));
  NOR2_X1   g0338(.A1(new_n538), .A2(new_n370), .ZN(new_n539));
  OAI21_X1  g0339(.A(new_n299), .B1(new_n539), .B2(new_n344), .ZN(new_n540));
  OAI211_X1 g0340(.A(new_n401), .B(new_n540), .C1(new_n403), .C2(new_n437), .ZN(new_n541));
  XNOR2_X1  g0341(.A(new_n541), .B(KEYINPUT13), .ZN(new_n542));
  INV_X1    g0342(.A(new_n542), .ZN(new_n543));
  OAI211_X1 g0343(.A(KEYINPUT74), .B(KEYINPUT14), .C1(new_n543), .C2(new_n332), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n543), .A2(G179), .ZN(new_n545));
  NAND2_X1  g0345(.A1(KEYINPUT74), .A2(KEYINPUT14), .ZN(new_n546));
  NAND3_X1  g0346(.A1(new_n542), .A2(G169), .A3(new_n546), .ZN(new_n547));
  NAND3_X1  g0347(.A1(new_n544), .A2(new_n545), .A3(new_n547), .ZN(new_n548));
  OAI22_X1  g0348(.A1(new_n426), .A2(new_n228), .B1(new_n210), .B2(G68), .ZN(new_n549));
  INV_X1    g0349(.A(G77), .ZN(new_n550));
  NOR2_X1   g0350(.A1(new_n354), .A2(new_n550), .ZN(new_n551));
  OAI21_X1  g0351(.A(new_n257), .B1(new_n549), .B2(new_n551), .ZN(new_n552));
  XOR2_X1   g0352(.A(new_n552), .B(KEYINPUT11), .Z(new_n553));
  OR2_X1    g0353(.A1(new_n553), .A2(KEYINPUT73), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n553), .A2(KEYINPUT73), .ZN(new_n555));
  OR3_X1    g0355(.A1(new_n283), .A2(KEYINPUT12), .A3(G68), .ZN(new_n556));
  OAI21_X1  g0356(.A(KEYINPUT12), .B1(new_n283), .B2(G68), .ZN(new_n557));
  AOI21_X1  g0357(.A(new_n202), .B1(new_n209), .B2(G20), .ZN(new_n558));
  AOI22_X1  g0358(.A1(new_n556), .A2(new_n557), .B1(new_n413), .B2(new_n558), .ZN(new_n559));
  NAND3_X1  g0359(.A1(new_n554), .A2(new_n555), .A3(new_n559), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n548), .A2(new_n560), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n543), .A2(G190), .ZN(new_n562));
  INV_X1    g0362(.A(new_n560), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n542), .A2(G200), .ZN(new_n564));
  AND3_X1   g0364(.A1(new_n562), .A2(new_n563), .A3(new_n564), .ZN(new_n565));
  INV_X1    g0365(.A(new_n565), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n561), .A2(new_n566), .ZN(new_n567));
  NOR3_X1   g0367(.A1(new_n462), .A2(new_n536), .A3(new_n567), .ZN(new_n568));
  NAND3_X1  g0368(.A1(new_n269), .A2(G257), .A3(G1698), .ZN(new_n569));
  INV_X1    g0369(.A(G294), .ZN(new_n570));
  OAI221_X1 g0370(.A(new_n569), .B1(new_n259), .B2(new_n570), .C1(new_n395), .C2(new_n365), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n571), .A2(new_n299), .ZN(new_n572));
  AND2_X1   g0372(.A1(new_n572), .A2(new_n320), .ZN(new_n573));
  NAND3_X1  g0373(.A1(new_n327), .A2(G264), .A3(new_n306), .ZN(new_n574));
  NAND3_X1  g0374(.A1(new_n573), .A2(new_n301), .A3(new_n574), .ZN(new_n575));
  NAND3_X1  g0375(.A1(new_n572), .A2(new_n320), .A3(new_n574), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n576), .A2(new_n332), .ZN(new_n577));
  NAND3_X1  g0377(.A1(new_n269), .A2(new_n210), .A3(G87), .ZN(new_n578));
  XNOR2_X1  g0378(.A(new_n578), .B(KEYINPUT22), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n223), .A2(G20), .ZN(new_n580));
  OAI22_X1  g0380(.A1(KEYINPUT23), .A2(new_n580), .B1(new_n354), .B2(new_n371), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n258), .A2(G20), .ZN(new_n582));
  AOI21_X1  g0382(.A(new_n581), .B1(new_n582), .B2(KEYINPUT23), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n579), .A2(new_n583), .ZN(new_n584));
  XOR2_X1   g0384(.A(KEYINPUT87), .B(KEYINPUT24), .Z(new_n585));
  NAND2_X1  g0385(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  INV_X1    g0386(.A(new_n585), .ZN(new_n587));
  NAND3_X1  g0387(.A1(new_n579), .A2(new_n587), .A3(new_n583), .ZN(new_n588));
  AOI21_X1  g0388(.A(new_n519), .B1(new_n586), .B2(new_n588), .ZN(new_n589));
  AND2_X1   g0389(.A1(new_n285), .A2(G107), .ZN(new_n590));
  NOR2_X1   g0390(.A1(new_n281), .A2(G1), .ZN(new_n591));
  NAND3_X1  g0391(.A1(new_n591), .A2(G20), .A3(new_n223), .ZN(new_n592));
  XNOR2_X1  g0392(.A(new_n592), .B(KEYINPUT25), .ZN(new_n593));
  NOR2_X1   g0393(.A1(new_n590), .A2(new_n593), .ZN(new_n594));
  INV_X1    g0394(.A(new_n594), .ZN(new_n595));
  OAI211_X1 g0395(.A(new_n575), .B(new_n577), .C1(new_n589), .C2(new_n595), .ZN(new_n596));
  INV_X1    g0396(.A(new_n588), .ZN(new_n597));
  AOI21_X1  g0397(.A(new_n587), .B1(new_n579), .B2(new_n583), .ZN(new_n598));
  OAI21_X1  g0398(.A(new_n257), .B1(new_n597), .B2(new_n598), .ZN(new_n599));
  NAND3_X1  g0399(.A1(new_n573), .A2(G190), .A3(new_n574), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n576), .A2(G200), .ZN(new_n601));
  NAND4_X1  g0401(.A1(new_n599), .A2(new_n600), .A3(new_n594), .A4(new_n601), .ZN(new_n602));
  AND2_X1   g0402(.A1(new_n596), .A2(new_n602), .ZN(new_n603));
  NAND3_X1  g0403(.A1(new_n327), .A2(G270), .A3(new_n306), .ZN(new_n604));
  AND2_X1   g0404(.A1(new_n604), .A2(new_n320), .ZN(new_n605));
  NAND3_X1  g0405(.A1(new_n269), .A2(G257), .A3(new_n394), .ZN(new_n606));
  INV_X1    g0406(.A(G303), .ZN(new_n607));
  OAI221_X1 g0407(.A(new_n606), .B1(new_n607), .B2(new_n269), .C1(new_n390), .C2(new_n224), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n608), .A2(new_n299), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n605), .A2(new_n609), .ZN(new_n610));
  NOR2_X1   g0410(.A1(new_n283), .A2(G116), .ZN(new_n611));
  AOI21_X1  g0411(.A(new_n611), .B1(new_n285), .B2(G116), .ZN(new_n612));
  OAI211_X1 g0412(.A(new_n294), .B(new_n210), .C1(G33), .C2(new_n343), .ZN(new_n613));
  OAI211_X1 g0413(.A(new_n613), .B(new_n257), .C1(new_n210), .C2(G116), .ZN(new_n614));
  INV_X1    g0414(.A(KEYINPUT20), .ZN(new_n615));
  XNOR2_X1  g0415(.A(new_n614), .B(new_n615), .ZN(new_n616));
  AOI21_X1  g0416(.A(new_n332), .B1(new_n612), .B2(new_n616), .ZN(new_n617));
  NAND3_X1  g0417(.A1(new_n610), .A2(KEYINPUT21), .A3(new_n617), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n612), .A2(new_n616), .ZN(new_n619));
  AOI21_X1  g0419(.A(new_n301), .B1(new_n608), .B2(new_n299), .ZN(new_n620));
  NAND3_X1  g0420(.A1(new_n619), .A2(new_n605), .A3(new_n620), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n618), .A2(new_n621), .ZN(new_n622));
  XNOR2_X1  g0422(.A(KEYINPUT86), .B(KEYINPUT21), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n610), .A2(new_n617), .ZN(new_n624));
  AOI21_X1  g0424(.A(new_n623), .B1(new_n624), .B2(KEYINPUT85), .ZN(new_n625));
  INV_X1    g0425(.A(KEYINPUT85), .ZN(new_n626));
  NAND3_X1  g0426(.A1(new_n610), .A2(new_n626), .A3(new_n617), .ZN(new_n627));
  AOI21_X1  g0427(.A(new_n622), .B1(new_n625), .B2(new_n627), .ZN(new_n628));
  AOI21_X1  g0428(.A(new_n619), .B1(new_n610), .B2(G200), .ZN(new_n629));
  OAI21_X1  g0429(.A(new_n629), .B1(new_n338), .B2(new_n610), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n628), .A2(new_n630), .ZN(new_n631));
  INV_X1    g0431(.A(new_n631), .ZN(new_n632));
  AND4_X1   g0432(.A1(new_n389), .A2(new_n568), .A3(new_n603), .A4(new_n632), .ZN(G372));
  NOR2_X1   g0433(.A1(new_n362), .A2(new_n376), .ZN(new_n634));
  OAI21_X1  g0434(.A(new_n602), .B1(new_n380), .B2(new_n378), .ZN(new_n635));
  NOR2_X1   g0435(.A1(new_n635), .A2(new_n340), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n628), .A2(new_n596), .ZN(new_n637));
  AOI21_X1  g0437(.A(new_n634), .B1(new_n636), .B2(new_n637), .ZN(new_n638));
  INV_X1    g0438(.A(new_n638), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n330), .A2(new_n335), .ZN(new_n640));
  INV_X1    g0440(.A(new_n640), .ZN(new_n641));
  NOR2_X1   g0441(.A1(new_n641), .A2(new_n381), .ZN(new_n642));
  XNOR2_X1  g0442(.A(KEYINPUT88), .B(KEYINPUT26), .ZN(new_n643));
  NAND3_X1  g0443(.A1(new_n333), .A2(new_n287), .A3(new_n321), .ZN(new_n644));
  OR2_X1    g0444(.A1(new_n381), .A2(new_n644), .ZN(new_n645));
  INV_X1    g0445(.A(KEYINPUT26), .ZN(new_n646));
  AOI22_X1  g0446(.A1(new_n642), .A2(new_n643), .B1(new_n645), .B2(new_n646), .ZN(new_n647));
  OR2_X1    g0447(.A1(new_n639), .A2(new_n647), .ZN(new_n648));
  AND2_X1   g0448(.A1(new_n568), .A2(new_n648), .ZN(new_n649));
  INV_X1    g0449(.A(new_n504), .ZN(new_n650));
  AOI21_X1  g0450(.A(new_n503), .B1(new_n477), .B2(new_n500), .ZN(new_n651));
  INV_X1    g0451(.A(KEYINPUT89), .ZN(new_n652));
  NOR3_X1   g0452(.A1(new_n650), .A2(new_n651), .A3(new_n652), .ZN(new_n653));
  AOI21_X1  g0453(.A(KEYINPUT89), .B1(new_n502), .B2(new_n504), .ZN(new_n654));
  NOR2_X1   g0454(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  INV_X1    g0455(.A(new_n655), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n561), .A2(new_n452), .ZN(new_n657));
  INV_X1    g0457(.A(new_n534), .ZN(new_n658));
  OAI21_X1  g0458(.A(new_n530), .B1(new_n509), .B2(new_n508), .ZN(new_n659));
  AOI21_X1  g0459(.A(new_n533), .B1(new_n659), .B2(KEYINPUT78), .ZN(new_n660));
  AOI21_X1  g0460(.A(new_n658), .B1(new_n531), .B2(new_n660), .ZN(new_n661));
  NOR2_X1   g0461(.A1(new_n661), .A2(new_n565), .ZN(new_n662));
  AOI21_X1  g0462(.A(new_n656), .B1(new_n657), .B2(new_n662), .ZN(new_n663));
  OAI21_X1  g0463(.A(new_n456), .B1(new_n663), .B2(new_n425), .ZN(new_n664));
  OR2_X1    g0464(.A1(new_n649), .A2(new_n664), .ZN(G369));
  INV_X1    g0465(.A(new_n596), .ZN(new_n666));
  INV_X1    g0466(.A(G213), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n591), .A2(new_n210), .ZN(new_n668));
  NOR2_X1   g0468(.A1(new_n668), .A2(KEYINPUT27), .ZN(new_n669));
  XNOR2_X1  g0469(.A(new_n669), .B(KEYINPUT90), .ZN(new_n670));
  AOI211_X1 g0470(.A(new_n667), .B(new_n670), .C1(KEYINPUT27), .C2(new_n668), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n671), .A2(G343), .ZN(new_n672));
  INV_X1    g0472(.A(new_n672), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n666), .A2(new_n673), .ZN(new_n674));
  XOR2_X1   g0474(.A(new_n674), .B(KEYINPUT92), .Z(new_n675));
  OAI21_X1  g0475(.A(new_n673), .B1(new_n589), .B2(new_n595), .ZN(new_n676));
  NAND3_X1  g0476(.A1(new_n676), .A2(new_n596), .A3(new_n602), .ZN(new_n677));
  XNOR2_X1  g0477(.A(new_n677), .B(KEYINPUT91), .ZN(new_n678));
  NOR2_X1   g0478(.A1(new_n675), .A2(new_n678), .ZN(new_n679));
  NOR2_X1   g0479(.A1(new_n628), .A2(new_n673), .ZN(new_n680));
  INV_X1    g0480(.A(new_n680), .ZN(new_n681));
  NOR2_X1   g0481(.A1(new_n679), .A2(new_n681), .ZN(new_n682));
  AOI21_X1  g0482(.A(new_n682), .B1(new_n666), .B2(new_n672), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n673), .A2(new_n619), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n632), .A2(new_n684), .ZN(new_n685));
  OAI21_X1  g0485(.A(new_n685), .B1(new_n628), .B2(new_n684), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n686), .A2(G330), .ZN(new_n687));
  NOR2_X1   g0487(.A1(new_n687), .A2(new_n679), .ZN(new_n688));
  INV_X1    g0488(.A(new_n688), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n683), .A2(new_n689), .ZN(G399));
  NAND3_X1  g0490(.A1(new_n350), .A2(new_n371), .A3(new_n351), .ZN(new_n691));
  INV_X1    g0491(.A(new_n691), .ZN(new_n692));
  INV_X1    g0492(.A(new_n213), .ZN(new_n693));
  NOR2_X1   g0493(.A1(new_n693), .A2(G41), .ZN(new_n694));
  INV_X1    g0494(.A(new_n694), .ZN(new_n695));
  NAND3_X1  g0495(.A1(new_n692), .A2(G1), .A3(new_n695), .ZN(new_n696));
  OAI21_X1  g0496(.A(new_n696), .B1(new_n216), .B2(new_n695), .ZN(new_n697));
  XNOR2_X1  g0497(.A(new_n697), .B(KEYINPUT28), .ZN(new_n698));
  INV_X1    g0498(.A(G330), .ZN(new_n699));
  AND4_X1   g0499(.A1(new_n603), .A2(new_n628), .A3(new_n630), .A4(new_n672), .ZN(new_n700));
  AND4_X1   g0500(.A1(new_n387), .A2(new_n342), .A3(new_n383), .A4(new_n382), .ZN(new_n701));
  AOI21_X1  g0501(.A(new_n387), .B1(new_n386), .B2(new_n383), .ZN(new_n702));
  OAI21_X1  g0502(.A(new_n700), .B1(new_n701), .B2(new_n702), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n703), .A2(KEYINPUT93), .ZN(new_n704));
  INV_X1    g0504(.A(KEYINPUT93), .ZN(new_n705));
  NAND3_X1  g0505(.A1(new_n389), .A2(new_n705), .A3(new_n700), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n704), .A2(new_n706), .ZN(new_n707));
  NOR2_X1   g0507(.A1(new_n576), .A2(new_n331), .ZN(new_n708));
  INV_X1    g0508(.A(new_n374), .ZN(new_n709));
  NAND4_X1  g0509(.A1(new_n708), .A2(new_n709), .A3(new_n604), .A4(new_n620), .ZN(new_n710));
  INV_X1    g0510(.A(KEYINPUT30), .ZN(new_n711));
  OR2_X1    g0511(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  NOR2_X1   g0512(.A1(new_n709), .A2(G179), .ZN(new_n713));
  NAND4_X1  g0513(.A1(new_n713), .A2(new_n610), .A3(new_n331), .A4(new_n576), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n710), .A2(new_n711), .ZN(new_n715));
  NAND3_X1  g0515(.A1(new_n712), .A2(new_n714), .A3(new_n715), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n716), .A2(new_n673), .ZN(new_n717));
  INV_X1    g0517(.A(KEYINPUT31), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  NAND3_X1  g0519(.A1(new_n716), .A2(KEYINPUT31), .A3(new_n673), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  INV_X1    g0521(.A(new_n721), .ZN(new_n722));
  AOI21_X1  g0522(.A(new_n699), .B1(new_n707), .B2(new_n722), .ZN(new_n723));
  INV_X1    g0523(.A(KEYINPUT29), .ZN(new_n724));
  OAI211_X1 g0524(.A(new_n724), .B(new_n672), .C1(new_n639), .C2(new_n647), .ZN(new_n725));
  OAI22_X1  g0525(.A1(new_n642), .A2(new_n643), .B1(new_n645), .B2(new_n646), .ZN(new_n726));
  AOI21_X1  g0526(.A(new_n673), .B1(new_n638), .B2(new_n726), .ZN(new_n727));
  OAI21_X1  g0527(.A(new_n725), .B1(new_n727), .B2(new_n724), .ZN(new_n728));
  NOR2_X1   g0528(.A1(new_n723), .A2(new_n728), .ZN(new_n729));
  OAI21_X1  g0529(.A(new_n698), .B1(new_n729), .B2(G1), .ZN(new_n730));
  XOR2_X1   g0530(.A(new_n730), .B(KEYINPUT94), .Z(G364));
  NOR2_X1   g0531(.A1(new_n281), .A2(G20), .ZN(new_n732));
  AOI21_X1  g0532(.A(new_n209), .B1(new_n732), .B2(G45), .ZN(new_n733));
  INV_X1    g0533(.A(new_n733), .ZN(new_n734));
  NOR2_X1   g0534(.A1(new_n694), .A2(new_n734), .ZN(new_n735));
  AOI21_X1  g0535(.A(new_n735), .B1(new_n686), .B2(G330), .ZN(new_n736));
  OAI21_X1  g0536(.A(new_n736), .B1(G330), .B2(new_n686), .ZN(new_n737));
  INV_X1    g0537(.A(new_n735), .ZN(new_n738));
  NOR2_X1   g0538(.A1(G13), .A2(G33), .ZN(new_n739));
  INV_X1    g0539(.A(new_n739), .ZN(new_n740));
  NOR2_X1   g0540(.A1(new_n740), .A2(G20), .ZN(new_n741));
  AOI21_X1  g0541(.A(new_n218), .B1(G20), .B2(new_n332), .ZN(new_n742));
  NOR2_X1   g0542(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  XNOR2_X1  g0543(.A(new_n743), .B(KEYINPUT96), .ZN(new_n744));
  NOR2_X1   g0544(.A1(new_n254), .A2(new_n399), .ZN(new_n745));
  NOR2_X1   g0545(.A1(new_n693), .A2(new_n269), .ZN(new_n746));
  INV_X1    g0546(.A(new_n746), .ZN(new_n747));
  AOI21_X1  g0547(.A(new_n747), .B1(new_n217), .B2(new_n399), .ZN(new_n748));
  INV_X1    g0548(.A(KEYINPUT95), .ZN(new_n749));
  AOI21_X1  g0549(.A(new_n745), .B1(new_n748), .B2(new_n749), .ZN(new_n750));
  OAI21_X1  g0550(.A(new_n750), .B1(new_n749), .B2(new_n748), .ZN(new_n751));
  NOR2_X1   g0551(.A1(new_n693), .A2(new_n370), .ZN(new_n752));
  AOI22_X1  g0552(.A1(new_n752), .A2(G355), .B1(new_n371), .B2(new_n693), .ZN(new_n753));
  AOI21_X1  g0553(.A(new_n744), .B1(new_n751), .B2(new_n753), .ZN(new_n754));
  INV_X1    g0554(.A(G283), .ZN(new_n755));
  AOI21_X1  g0555(.A(KEYINPUT97), .B1(new_n301), .B2(G200), .ZN(new_n756));
  NOR2_X1   g0556(.A1(new_n756), .A2(new_n210), .ZN(new_n757));
  NAND3_X1  g0557(.A1(new_n301), .A2(KEYINPUT97), .A3(G200), .ZN(new_n758));
  NAND2_X1  g0558(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n759), .A2(G190), .ZN(new_n760));
  INV_X1    g0560(.A(new_n760), .ZN(new_n761));
  NOR2_X1   g0561(.A1(new_n759), .A2(new_n338), .ZN(new_n762));
  INV_X1    g0562(.A(new_n762), .ZN(new_n763));
  OAI22_X1  g0563(.A1(new_n755), .A2(new_n761), .B1(new_n763), .B2(new_n607), .ZN(new_n764));
  NOR2_X1   g0564(.A1(new_n210), .A2(new_n301), .ZN(new_n765));
  NAND2_X1  g0565(.A1(new_n765), .A2(G200), .ZN(new_n766));
  NOR2_X1   g0566(.A1(new_n766), .A2(G190), .ZN(new_n767));
  NOR2_X1   g0567(.A1(KEYINPUT33), .A2(G317), .ZN(new_n768));
  AND2_X1   g0568(.A1(KEYINPUT33), .A2(G317), .ZN(new_n769));
  OAI21_X1  g0569(.A(new_n767), .B1(new_n768), .B2(new_n769), .ZN(new_n770));
  NOR3_X1   g0570(.A1(new_n338), .A2(G179), .A3(G200), .ZN(new_n771));
  NOR2_X1   g0571(.A1(new_n771), .A2(new_n210), .ZN(new_n772));
  INV_X1    g0572(.A(G326), .ZN(new_n773));
  NOR2_X1   g0573(.A1(new_n766), .A2(new_n338), .ZN(new_n774));
  INV_X1    g0574(.A(new_n774), .ZN(new_n775));
  OAI221_X1 g0575(.A(new_n770), .B1(new_n570), .B2(new_n772), .C1(new_n773), .C2(new_n775), .ZN(new_n776));
  NAND3_X1  g0576(.A1(new_n765), .A2(G190), .A3(new_n458), .ZN(new_n777));
  INV_X1    g0577(.A(new_n777), .ZN(new_n778));
  NOR2_X1   g0578(.A1(G190), .A2(G200), .ZN(new_n779));
  NAND3_X1  g0579(.A1(new_n779), .A2(G20), .A3(new_n301), .ZN(new_n780));
  INV_X1    g0580(.A(new_n780), .ZN(new_n781));
  AOI22_X1  g0581(.A1(new_n778), .A2(G322), .B1(G329), .B2(new_n781), .ZN(new_n782));
  INV_X1    g0582(.A(G311), .ZN(new_n783));
  NAND2_X1  g0583(.A1(new_n765), .A2(new_n779), .ZN(new_n784));
  OAI211_X1 g0584(.A(new_n782), .B(new_n370), .C1(new_n783), .C2(new_n784), .ZN(new_n785));
  NOR3_X1   g0585(.A1(new_n764), .A2(new_n776), .A3(new_n785), .ZN(new_n786));
  OR2_X1    g0586(.A1(new_n786), .A2(KEYINPUT98), .ZN(new_n787));
  NAND2_X1  g0587(.A1(new_n786), .A2(KEYINPUT98), .ZN(new_n788));
  NOR2_X1   g0588(.A1(new_n772), .A2(new_n343), .ZN(new_n789));
  OAI221_X1 g0589(.A(new_n269), .B1(new_n784), .B2(new_n233), .C1(new_n201), .C2(new_n777), .ZN(new_n790));
  AOI211_X1 g0590(.A(new_n789), .B(new_n790), .C1(G68), .C2(new_n767), .ZN(new_n791));
  INV_X1    g0591(.A(KEYINPUT32), .ZN(new_n792));
  INV_X1    g0592(.A(G159), .ZN(new_n793));
  NOR2_X1   g0593(.A1(new_n780), .A2(new_n793), .ZN(new_n794));
  OAI22_X1  g0594(.A1(new_n775), .A2(new_n228), .B1(new_n792), .B2(new_n794), .ZN(new_n795));
  AOI21_X1  g0595(.A(new_n795), .B1(new_n792), .B2(new_n794), .ZN(new_n796));
  NAND2_X1  g0596(.A1(new_n762), .A2(G87), .ZN(new_n797));
  NAND2_X1  g0597(.A1(new_n760), .A2(G107), .ZN(new_n798));
  NAND4_X1  g0598(.A1(new_n791), .A2(new_n796), .A3(new_n797), .A4(new_n798), .ZN(new_n799));
  NAND3_X1  g0599(.A1(new_n787), .A2(new_n788), .A3(new_n799), .ZN(new_n800));
  AOI211_X1 g0600(.A(new_n738), .B(new_n754), .C1(new_n800), .C2(new_n742), .ZN(new_n801));
  INV_X1    g0601(.A(new_n741), .ZN(new_n802));
  OAI21_X1  g0602(.A(new_n801), .B1(new_n686), .B2(new_n802), .ZN(new_n803));
  AND2_X1   g0603(.A1(new_n737), .A2(new_n803), .ZN(new_n804));
  INV_X1    g0604(.A(new_n804), .ZN(G396));
  NOR2_X1   g0605(.A1(new_n742), .A2(new_n739), .ZN(new_n806));
  AOI21_X1  g0606(.A(new_n738), .B1(new_n550), .B2(new_n806), .ZN(new_n807));
  INV_X1    g0607(.A(new_n742), .ZN(new_n808));
  INV_X1    g0608(.A(new_n784), .ZN(new_n809));
  AOI22_X1  g0609(.A1(new_n778), .A2(G143), .B1(new_n809), .B2(G159), .ZN(new_n810));
  NAND2_X1  g0610(.A1(new_n767), .A2(G150), .ZN(new_n811));
  INV_X1    g0611(.A(G137), .ZN(new_n812));
  OAI211_X1 g0612(.A(new_n810), .B(new_n811), .C1(new_n812), .C2(new_n775), .ZN(new_n813));
  XOR2_X1   g0613(.A(KEYINPUT99), .B(KEYINPUT34), .Z(new_n814));
  XNOR2_X1  g0614(.A(new_n813), .B(new_n814), .ZN(new_n815));
  NAND2_X1  g0615(.A1(new_n760), .A2(G68), .ZN(new_n816));
  AOI21_X1  g0616(.A(new_n370), .B1(new_n781), .B2(G132), .ZN(new_n817));
  OAI211_X1 g0617(.A(new_n816), .B(new_n817), .C1(new_n201), .C2(new_n772), .ZN(new_n818));
  AOI21_X1  g0618(.A(new_n818), .B1(G50), .B2(new_n762), .ZN(new_n819));
  AOI21_X1  g0619(.A(new_n789), .B1(G303), .B2(new_n774), .ZN(new_n820));
  INV_X1    g0620(.A(new_n767), .ZN(new_n821));
  OAI21_X1  g0621(.A(new_n820), .B1(new_n755), .B2(new_n821), .ZN(new_n822));
  OAI21_X1  g0622(.A(new_n370), .B1(new_n777), .B2(new_n570), .ZN(new_n823));
  OAI22_X1  g0623(.A1(new_n784), .A2(new_n371), .B1(new_n780), .B2(new_n783), .ZN(new_n824));
  NOR3_X1   g0624(.A1(new_n822), .A2(new_n823), .A3(new_n824), .ZN(new_n825));
  AOI22_X1  g0625(.A1(G87), .A2(new_n760), .B1(new_n762), .B2(G107), .ZN(new_n826));
  AOI22_X1  g0626(.A1(new_n815), .A2(new_n819), .B1(new_n825), .B2(new_n826), .ZN(new_n827));
  INV_X1    g0627(.A(new_n435), .ZN(new_n828));
  NOR3_X1   g0628(.A1(new_n441), .A2(new_n443), .A3(new_n436), .ZN(new_n829));
  AOI21_X1  g0629(.A(KEYINPUT71), .B1(new_n445), .B2(new_n447), .ZN(new_n830));
  OAI21_X1  g0630(.A(new_n301), .B1(new_n829), .B2(new_n830), .ZN(new_n831));
  AND4_X1   g0631(.A1(new_n828), .A2(new_n831), .A3(new_n451), .A4(new_n672), .ZN(new_n832));
  OAI22_X1  g0632(.A1(new_n459), .A2(new_n460), .B1(new_n435), .B2(new_n672), .ZN(new_n833));
  AOI21_X1  g0633(.A(new_n832), .B1(new_n452), .B2(new_n833), .ZN(new_n834));
  OAI221_X1 g0634(.A(new_n807), .B1(new_n808), .B2(new_n827), .C1(new_n834), .C2(new_n740), .ZN(new_n835));
  INV_X1    g0635(.A(KEYINPUT100), .ZN(new_n836));
  XNOR2_X1  g0636(.A(new_n834), .B(new_n836), .ZN(new_n837));
  NAND2_X1  g0637(.A1(new_n648), .A2(new_n672), .ZN(new_n838));
  NAND2_X1  g0638(.A1(new_n837), .A2(new_n838), .ZN(new_n839));
  OAI211_X1 g0639(.A(new_n834), .B(new_n672), .C1(new_n639), .C2(new_n647), .ZN(new_n840));
  NAND2_X1  g0640(.A1(new_n839), .A2(new_n840), .ZN(new_n841));
  INV_X1    g0641(.A(new_n723), .ZN(new_n842));
  NOR2_X1   g0642(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  XNOR2_X1  g0643(.A(new_n843), .B(KEYINPUT101), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n841), .A2(new_n842), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n845), .A2(new_n738), .ZN(new_n846));
  OAI21_X1  g0646(.A(new_n835), .B1(new_n844), .B2(new_n846), .ZN(G384));
  INV_X1    g0647(.A(new_n278), .ZN(new_n848));
  OR2_X1    g0648(.A1(new_n848), .A2(KEYINPUT35), .ZN(new_n849));
  NAND2_X1  g0649(.A1(new_n848), .A2(KEYINPUT35), .ZN(new_n850));
  NAND4_X1  g0650(.A1(new_n849), .A2(G116), .A3(new_n219), .A4(new_n850), .ZN(new_n851));
  XOR2_X1   g0651(.A(new_n851), .B(KEYINPUT36), .Z(new_n852));
  NAND3_X1  g0652(.A1(new_n217), .A2(new_n433), .A3(new_n469), .ZN(new_n853));
  AOI211_X1 g0653(.A(new_n209), .B(G13), .C1(new_n853), .C2(new_n250), .ZN(new_n854));
  NOR2_X1   g0654(.A1(new_n852), .A2(new_n854), .ZN(new_n855));
  NAND3_X1  g0655(.A1(new_n548), .A2(new_n560), .A3(new_n672), .ZN(new_n856));
  NOR2_X1   g0656(.A1(new_n525), .A2(KEYINPUT16), .ZN(new_n857));
  OAI21_X1  g0657(.A(new_n464), .B1(new_n857), .B2(new_n473), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n858), .A2(new_n671), .ZN(new_n859));
  INV_X1    g0659(.A(new_n859), .ZN(new_n860));
  NAND3_X1  g0660(.A1(new_n516), .A2(new_n517), .A3(new_n530), .ZN(new_n861));
  OAI21_X1  g0661(.A(new_n858), .B1(new_n671), .B2(new_n500), .ZN(new_n862));
  NAND3_X1  g0662(.A1(new_n511), .A2(new_n861), .A3(new_n862), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n863), .A2(KEYINPUT37), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n671), .A2(new_n477), .ZN(new_n865));
  INV_X1    g0665(.A(KEYINPUT37), .ZN(new_n866));
  AND3_X1   g0666(.A1(new_n865), .A2(new_n501), .A3(new_n866), .ZN(new_n867));
  NAND3_X1  g0667(.A1(new_n867), .A2(new_n511), .A3(new_n861), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n864), .A2(new_n868), .ZN(new_n869));
  INV_X1    g0669(.A(KEYINPUT102), .ZN(new_n870));
  AOI22_X1  g0670(.A1(new_n536), .A2(new_n860), .B1(new_n869), .B2(new_n870), .ZN(new_n871));
  NAND3_X1  g0671(.A1(new_n864), .A2(KEYINPUT102), .A3(new_n868), .ZN(new_n872));
  AOI21_X1  g0672(.A(KEYINPUT38), .B1(new_n871), .B2(new_n872), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n869), .A2(new_n870), .ZN(new_n874));
  OAI21_X1  g0674(.A(new_n860), .B1(new_n661), .B2(new_n505), .ZN(new_n875));
  NAND4_X1  g0675(.A1(new_n874), .A2(new_n875), .A3(KEYINPUT38), .A4(new_n872), .ZN(new_n876));
  INV_X1    g0676(.A(new_n876), .ZN(new_n877));
  OAI21_X1  g0677(.A(KEYINPUT39), .B1(new_n873), .B2(new_n877), .ZN(new_n878));
  INV_X1    g0678(.A(KEYINPUT104), .ZN(new_n879));
  INV_X1    g0679(.A(KEYINPUT38), .ZN(new_n880));
  INV_X1    g0680(.A(new_n868), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n499), .A2(new_n332), .ZN(new_n882));
  NAND4_X1  g0682(.A1(new_n483), .A2(new_n496), .A3(new_n301), .A4(new_n489), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  OAI21_X1  g0684(.A(KEYINPUT89), .B1(new_n530), .B2(new_n884), .ZN(new_n885));
  NAND3_X1  g0685(.A1(new_n477), .A2(new_n500), .A3(new_n652), .ZN(new_n886));
  NAND3_X1  g0686(.A1(new_n885), .A2(new_n659), .A3(new_n886), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n887), .A2(KEYINPUT103), .ZN(new_n888));
  INV_X1    g0688(.A(KEYINPUT103), .ZN(new_n889));
  NAND4_X1  g0689(.A1(new_n885), .A2(new_n659), .A3(new_n889), .A4(new_n886), .ZN(new_n890));
  NAND3_X1  g0690(.A1(new_n888), .A2(new_n865), .A3(new_n890), .ZN(new_n891));
  AOI21_X1  g0691(.A(new_n881), .B1(new_n891), .B2(KEYINPUT37), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n532), .A2(new_n534), .ZN(new_n893));
  AOI21_X1  g0693(.A(new_n865), .B1(new_n893), .B2(new_n655), .ZN(new_n894));
  OAI21_X1  g0694(.A(new_n880), .B1(new_n892), .B2(new_n894), .ZN(new_n895));
  INV_X1    g0695(.A(KEYINPUT39), .ZN(new_n896));
  NAND3_X1  g0696(.A1(new_n876), .A2(new_n895), .A3(new_n896), .ZN(new_n897));
  NAND3_X1  g0697(.A1(new_n878), .A2(new_n879), .A3(new_n897), .ZN(new_n898));
  AND2_X1   g0698(.A1(new_n511), .A2(new_n861), .ZN(new_n899));
  AOI22_X1  g0699(.A1(new_n899), .A2(new_n867), .B1(new_n863), .B2(KEYINPUT37), .ZN(new_n900));
  OAI22_X1  g0700(.A1(new_n900), .A2(KEYINPUT102), .B1(new_n535), .B2(new_n859), .ZN(new_n901));
  INV_X1    g0701(.A(new_n872), .ZN(new_n902));
  OAI21_X1  g0702(.A(new_n880), .B1(new_n901), .B2(new_n902), .ZN(new_n903));
  AOI21_X1  g0703(.A(new_n896), .B1(new_n903), .B2(new_n876), .ZN(new_n904));
  AND3_X1   g0704(.A1(new_n876), .A2(new_n895), .A3(new_n896), .ZN(new_n905));
  OAI21_X1  g0705(.A(KEYINPUT104), .B1(new_n904), .B2(new_n905), .ZN(new_n906));
  AOI21_X1  g0706(.A(new_n856), .B1(new_n898), .B2(new_n906), .ZN(new_n907));
  INV_X1    g0707(.A(new_n832), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n840), .A2(new_n908), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n673), .A2(new_n560), .ZN(new_n910));
  NAND3_X1  g0710(.A1(new_n561), .A2(new_n566), .A3(new_n910), .ZN(new_n911));
  OAI211_X1 g0711(.A(new_n560), .B(new_n673), .C1(new_n548), .C2(new_n565), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n909), .A2(new_n913), .ZN(new_n914));
  NOR2_X1   g0714(.A1(new_n873), .A2(new_n877), .ZN(new_n915));
  OAI22_X1  g0715(.A1(new_n914), .A2(new_n915), .B1(new_n655), .B2(new_n671), .ZN(new_n916));
  NOR2_X1   g0716(.A1(new_n907), .A2(new_n916), .ZN(new_n917));
  AOI21_X1  g0717(.A(new_n664), .B1(new_n568), .B2(new_n728), .ZN(new_n918));
  XNOR2_X1  g0718(.A(new_n917), .B(new_n918), .ZN(new_n919));
  NOR2_X1   g0719(.A1(new_n703), .A2(KEYINPUT93), .ZN(new_n920));
  AOI21_X1  g0720(.A(new_n705), .B1(new_n389), .B2(new_n700), .ZN(new_n921));
  OAI21_X1  g0721(.A(new_n722), .B1(new_n920), .B2(new_n921), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n876), .A2(new_n895), .ZN(new_n923));
  INV_X1    g0723(.A(new_n834), .ZN(new_n924));
  AOI21_X1  g0724(.A(new_n924), .B1(new_n911), .B2(new_n912), .ZN(new_n925));
  NAND3_X1  g0725(.A1(new_n922), .A2(new_n923), .A3(new_n925), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n926), .A2(KEYINPUT40), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n913), .A2(new_n834), .ZN(new_n928));
  AOI21_X1  g0728(.A(new_n928), .B1(new_n707), .B2(new_n722), .ZN(new_n929));
  AOI21_X1  g0729(.A(KEYINPUT40), .B1(new_n903), .B2(new_n876), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n927), .A2(new_n931), .ZN(new_n932));
  NAND3_X1  g0732(.A1(new_n932), .A2(new_n568), .A3(new_n922), .ZN(new_n933));
  AOI22_X1  g0733(.A1(new_n926), .A2(KEYINPUT40), .B1(new_n929), .B2(new_n930), .ZN(new_n934));
  INV_X1    g0734(.A(new_n568), .ZN(new_n935));
  AOI21_X1  g0735(.A(new_n721), .B1(new_n704), .B2(new_n706), .ZN(new_n936));
  OAI21_X1  g0736(.A(new_n934), .B1(new_n935), .B2(new_n936), .ZN(new_n937));
  NAND3_X1  g0737(.A1(new_n933), .A2(G330), .A3(new_n937), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n919), .A2(new_n938), .ZN(new_n939));
  OAI21_X1  g0739(.A(new_n939), .B1(new_n209), .B2(new_n732), .ZN(new_n940));
  NOR2_X1   g0740(.A1(new_n919), .A2(new_n938), .ZN(new_n941));
  OAI21_X1  g0741(.A(new_n855), .B1(new_n940), .B2(new_n941), .ZN(G367));
  NAND2_X1  g0742(.A1(new_n673), .A2(new_n380), .ZN(new_n943));
  MUX2_X1   g0743(.A(new_n634), .B(new_n382), .S(new_n943), .Z(new_n944));
  NAND2_X1  g0744(.A1(new_n944), .A2(KEYINPUT43), .ZN(new_n945));
  XOR2_X1   g0745(.A(new_n945), .B(KEYINPUT106), .Z(new_n946));
  OAI211_X1 g0746(.A(new_n641), .B(new_n339), .C1(new_n336), .C2(new_n672), .ZN(new_n947));
  OR2_X1    g0747(.A1(new_n672), .A2(new_n644), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n682), .A2(new_n949), .ZN(new_n950));
  NOR2_X1   g0750(.A1(new_n950), .A2(KEYINPUT42), .ZN(new_n951));
  XOR2_X1   g0751(.A(new_n951), .B(KEYINPUT105), .Z(new_n952));
  NAND2_X1  g0752(.A1(new_n949), .A2(new_n666), .ZN(new_n953));
  AOI21_X1  g0753(.A(new_n673), .B1(new_n953), .B2(new_n641), .ZN(new_n954));
  AOI21_X1  g0754(.A(new_n954), .B1(new_n950), .B2(KEYINPUT42), .ZN(new_n955));
  AOI21_X1  g0755(.A(new_n946), .B1(new_n952), .B2(new_n955), .ZN(new_n956));
  INV_X1    g0756(.A(KEYINPUT107), .ZN(new_n957));
  OR2_X1    g0757(.A1(new_n944), .A2(KEYINPUT43), .ZN(new_n958));
  AOI21_X1  g0758(.A(new_n956), .B1(new_n957), .B2(new_n958), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n688), .A2(new_n949), .ZN(new_n960));
  XNOR2_X1  g0760(.A(new_n959), .B(new_n960), .ZN(new_n961));
  NOR2_X1   g0761(.A1(new_n958), .A2(new_n957), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n961), .A2(new_n962), .ZN(new_n963));
  OR2_X1    g0763(.A1(new_n961), .A2(new_n962), .ZN(new_n964));
  XNOR2_X1  g0764(.A(KEYINPUT108), .B(KEYINPUT41), .ZN(new_n965));
  XOR2_X1   g0765(.A(new_n694), .B(new_n965), .Z(new_n966));
  NAND2_X1  g0766(.A1(new_n683), .A2(new_n949), .ZN(new_n967));
  XOR2_X1   g0767(.A(new_n967), .B(KEYINPUT109), .Z(new_n968));
  NAND2_X1  g0768(.A1(new_n968), .A2(KEYINPUT45), .ZN(new_n969));
  XNOR2_X1  g0769(.A(new_n967), .B(KEYINPUT109), .ZN(new_n970));
  INV_X1    g0770(.A(KEYINPUT45), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n970), .A2(new_n971), .ZN(new_n972));
  NOR2_X1   g0772(.A1(new_n683), .A2(new_n949), .ZN(new_n973));
  XNOR2_X1  g0773(.A(new_n973), .B(KEYINPUT44), .ZN(new_n974));
  NAND3_X1  g0774(.A1(new_n969), .A2(new_n972), .A3(new_n974), .ZN(new_n975));
  XNOR2_X1  g0775(.A(new_n975), .B(new_n689), .ZN(new_n976));
  AOI21_X1  g0776(.A(KEYINPUT110), .B1(new_n679), .B2(new_n681), .ZN(new_n977));
  XOR2_X1   g0777(.A(new_n977), .B(new_n687), .Z(new_n978));
  XNOR2_X1  g0778(.A(new_n978), .B(new_n682), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n979), .A2(new_n729), .ZN(new_n980));
  INV_X1    g0780(.A(new_n980), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n976), .A2(new_n981), .ZN(new_n982));
  AOI21_X1  g0782(.A(new_n966), .B1(new_n982), .B2(new_n729), .ZN(new_n983));
  OAI211_X1 g0783(.A(new_n963), .B(new_n964), .C1(new_n983), .C2(new_n734), .ZN(new_n984));
  AOI21_X1  g0784(.A(new_n744), .B1(new_n693), .B2(new_n360), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n746), .A2(new_n245), .ZN(new_n986));
  AOI21_X1  g0786(.A(new_n738), .B1(new_n985), .B2(new_n986), .ZN(new_n987));
  OAI22_X1  g0787(.A1(new_n201), .A2(new_n763), .B1(new_n761), .B2(new_n233), .ZN(new_n988));
  AOI22_X1  g0788(.A1(new_n778), .A2(G150), .B1(G137), .B2(new_n781), .ZN(new_n989));
  OAI211_X1 g0789(.A(new_n989), .B(new_n269), .C1(new_n228), .C2(new_n784), .ZN(new_n990));
  NAND2_X1  g0790(.A1(new_n774), .A2(G143), .ZN(new_n991));
  OAI221_X1 g0791(.A(new_n991), .B1(new_n202), .B2(new_n772), .C1(new_n821), .C2(new_n793), .ZN(new_n992));
  NOR3_X1   g0792(.A1(new_n988), .A2(new_n990), .A3(new_n992), .ZN(new_n993));
  NOR2_X1   g0793(.A1(new_n761), .A2(new_n343), .ZN(new_n994));
  INV_X1    g0794(.A(new_n772), .ZN(new_n995));
  AOI22_X1  g0795(.A1(new_n347), .A2(new_n995), .B1(new_n774), .B2(G311), .ZN(new_n996));
  AOI21_X1  g0796(.A(new_n269), .B1(new_n781), .B2(G317), .ZN(new_n997));
  AOI22_X1  g0797(.A1(new_n778), .A2(G303), .B1(new_n809), .B2(G283), .ZN(new_n998));
  NAND3_X1  g0798(.A1(new_n996), .A2(new_n997), .A3(new_n998), .ZN(new_n999));
  INV_X1    g0799(.A(KEYINPUT46), .ZN(new_n1000));
  OAI21_X1  g0800(.A(new_n1000), .B1(new_n763), .B2(new_n371), .ZN(new_n1001));
  NAND3_X1  g0801(.A1(new_n762), .A2(KEYINPUT46), .A3(G116), .ZN(new_n1002));
  OAI211_X1 g0802(.A(new_n1001), .B(new_n1002), .C1(new_n570), .C2(new_n821), .ZN(new_n1003));
  AOI211_X1 g0803(.A(new_n994), .B(new_n999), .C1(new_n1003), .C2(KEYINPUT111), .ZN(new_n1004));
  OR2_X1    g0804(.A1(new_n1003), .A2(KEYINPUT111), .ZN(new_n1005));
  AOI21_X1  g0805(.A(new_n993), .B1(new_n1004), .B2(new_n1005), .ZN(new_n1006));
  XNOR2_X1  g0806(.A(new_n1006), .B(KEYINPUT47), .ZN(new_n1007));
  OAI221_X1 g0807(.A(new_n987), .B1(new_n944), .B2(new_n802), .C1(new_n1007), .C2(new_n808), .ZN(new_n1008));
  NAND2_X1  g0808(.A1(new_n984), .A2(new_n1008), .ZN(G387));
  OAI21_X1  g0809(.A(new_n746), .B1(new_n242), .B2(new_n399), .ZN(new_n1010));
  INV_X1    g0810(.A(new_n752), .ZN(new_n1011));
  OAI21_X1  g0811(.A(new_n1010), .B1(new_n692), .B2(new_n1011), .ZN(new_n1012));
  OAI21_X1  g0812(.A(new_n399), .B1(new_n202), .B2(new_n550), .ZN(new_n1013));
  INV_X1    g0813(.A(new_n410), .ZN(new_n1014));
  NAND2_X1  g0814(.A1(new_n1014), .A2(new_n228), .ZN(new_n1015));
  AOI21_X1  g0815(.A(new_n1013), .B1(new_n1015), .B2(KEYINPUT50), .ZN(new_n1016));
  OAI211_X1 g0816(.A(new_n692), .B(new_n1016), .C1(KEYINPUT50), .C2(new_n1015), .ZN(new_n1017));
  AOI22_X1  g0817(.A1(new_n1012), .A2(new_n1017), .B1(new_n223), .B2(new_n693), .ZN(new_n1018));
  AOI22_X1  g0818(.A1(G159), .A2(new_n774), .B1(new_n767), .B2(new_n1014), .ZN(new_n1019));
  OAI21_X1  g0819(.A(new_n1019), .B1(new_n358), .B2(new_n772), .ZN(new_n1020));
  NOR2_X1   g0820(.A1(new_n763), .A2(new_n233), .ZN(new_n1021));
  AOI21_X1  g0821(.A(new_n370), .B1(new_n781), .B2(G150), .ZN(new_n1022));
  OAI221_X1 g0822(.A(new_n1022), .B1(new_n228), .B2(new_n777), .C1(new_n202), .C2(new_n784), .ZN(new_n1023));
  NOR4_X1   g0823(.A1(new_n1020), .A2(new_n994), .A3(new_n1021), .A4(new_n1023), .ZN(new_n1024));
  AOI22_X1  g0824(.A1(new_n778), .A2(G317), .B1(new_n809), .B2(G303), .ZN(new_n1025));
  INV_X1    g0825(.A(G322), .ZN(new_n1026));
  OAI221_X1 g0826(.A(new_n1025), .B1(new_n821), .B2(new_n783), .C1(new_n1026), .C2(new_n775), .ZN(new_n1027));
  INV_X1    g0827(.A(KEYINPUT48), .ZN(new_n1028));
  OR2_X1    g0828(.A1(new_n1027), .A2(new_n1028), .ZN(new_n1029));
  NAND2_X1  g0829(.A1(new_n1027), .A2(new_n1028), .ZN(new_n1030));
  AOI22_X1  g0830(.A1(new_n762), .A2(G294), .B1(G283), .B2(new_n995), .ZN(new_n1031));
  NAND3_X1  g0831(.A1(new_n1029), .A2(new_n1030), .A3(new_n1031), .ZN(new_n1032));
  XOR2_X1   g0832(.A(new_n1032), .B(KEYINPUT49), .Z(new_n1033));
  OR2_X1    g0833(.A1(new_n1033), .A2(KEYINPUT112), .ZN(new_n1034));
  OAI221_X1 g0834(.A(new_n370), .B1(new_n773), .B2(new_n780), .C1(new_n761), .C2(new_n371), .ZN(new_n1035));
  AOI21_X1  g0835(.A(new_n1035), .B1(new_n1033), .B2(KEYINPUT112), .ZN(new_n1036));
  AOI21_X1  g0836(.A(new_n1024), .B1(new_n1034), .B2(new_n1036), .ZN(new_n1037));
  OAI221_X1 g0837(.A(new_n735), .B1(new_n744), .B2(new_n1018), .C1(new_n1037), .C2(new_n808), .ZN(new_n1038));
  AOI21_X1  g0838(.A(new_n1038), .B1(new_n679), .B2(new_n741), .ZN(new_n1039));
  AOI21_X1  g0839(.A(new_n1039), .B1(new_n979), .B2(new_n734), .ZN(new_n1040));
  NAND2_X1  g0840(.A1(new_n980), .A2(new_n694), .ZN(new_n1041));
  NOR2_X1   g0841(.A1(new_n979), .A2(new_n729), .ZN(new_n1042));
  OAI21_X1  g0842(.A(new_n1040), .B1(new_n1041), .B2(new_n1042), .ZN(G393));
  AOI21_X1  g0843(.A(new_n695), .B1(new_n976), .B2(new_n981), .ZN(new_n1044));
  OAI21_X1  g0844(.A(new_n1044), .B1(new_n981), .B2(new_n976), .ZN(new_n1045));
  NAND3_X1  g0845(.A1(new_n947), .A2(new_n741), .A3(new_n948), .ZN(new_n1046));
  INV_X1    g0846(.A(new_n744), .ZN(new_n1047));
  OAI21_X1  g0847(.A(new_n1047), .B1(new_n343), .B2(new_n213), .ZN(new_n1048));
  NOR2_X1   g0848(.A1(new_n747), .A2(new_n249), .ZN(new_n1049));
  OAI21_X1  g0849(.A(new_n735), .B1(new_n1048), .B2(new_n1049), .ZN(new_n1050));
  OAI22_X1  g0850(.A1(new_n821), .A2(new_n607), .B1(new_n371), .B2(new_n772), .ZN(new_n1051));
  XNOR2_X1  g0851(.A(new_n1051), .B(KEYINPUT113), .ZN(new_n1052));
  OAI21_X1  g0852(.A(new_n370), .B1(new_n780), .B2(new_n1026), .ZN(new_n1053));
  AOI21_X1  g0853(.A(new_n1053), .B1(G294), .B2(new_n809), .ZN(new_n1054));
  NAND3_X1  g0854(.A1(new_n1052), .A2(new_n798), .A3(new_n1054), .ZN(new_n1055));
  NAND2_X1  g0855(.A1(new_n774), .A2(G317), .ZN(new_n1056));
  OAI21_X1  g0856(.A(new_n1056), .B1(new_n783), .B2(new_n777), .ZN(new_n1057));
  INV_X1    g0857(.A(KEYINPUT52), .ZN(new_n1058));
  AOI22_X1  g0858(.A1(new_n1057), .A2(new_n1058), .B1(G283), .B2(new_n762), .ZN(new_n1059));
  OAI21_X1  g0859(.A(new_n1059), .B1(new_n1058), .B2(new_n1057), .ZN(new_n1060));
  NAND2_X1  g0860(.A1(new_n760), .A2(G87), .ZN(new_n1061));
  NOR2_X1   g0861(.A1(new_n772), .A2(new_n550), .ZN(new_n1062));
  AOI21_X1  g0862(.A(new_n1062), .B1(G50), .B2(new_n767), .ZN(new_n1063));
  NAND2_X1  g0863(.A1(new_n781), .A2(G143), .ZN(new_n1064));
  AOI21_X1  g0864(.A(new_n370), .B1(new_n809), .B2(new_n1014), .ZN(new_n1065));
  NAND4_X1  g0865(.A1(new_n1061), .A2(new_n1063), .A3(new_n1064), .A4(new_n1065), .ZN(new_n1066));
  AOI22_X1  g0866(.A1(G150), .A2(new_n774), .B1(new_n778), .B2(G159), .ZN(new_n1067));
  AOI22_X1  g0867(.A1(new_n1067), .A2(KEYINPUT51), .B1(new_n762), .B2(G68), .ZN(new_n1068));
  OAI21_X1  g0868(.A(new_n1068), .B1(KEYINPUT51), .B2(new_n1067), .ZN(new_n1069));
  OAI22_X1  g0869(.A1(new_n1055), .A2(new_n1060), .B1(new_n1066), .B2(new_n1069), .ZN(new_n1070));
  AOI21_X1  g0870(.A(new_n1050), .B1(new_n1070), .B2(new_n742), .ZN(new_n1071));
  AOI22_X1  g0871(.A1(new_n976), .A2(new_n734), .B1(new_n1046), .B2(new_n1071), .ZN(new_n1072));
  NAND2_X1  g0872(.A1(new_n1045), .A2(new_n1072), .ZN(G390));
  NAND2_X1  g0873(.A1(new_n914), .A2(new_n856), .ZN(new_n1074));
  NAND3_X1  g0874(.A1(new_n898), .A2(new_n906), .A3(new_n1074), .ZN(new_n1075));
  NAND2_X1  g0875(.A1(new_n833), .A2(new_n452), .ZN(new_n1076));
  AOI21_X1  g0876(.A(new_n832), .B1(new_n727), .B2(new_n1076), .ZN(new_n1077));
  INV_X1    g0877(.A(new_n913), .ZN(new_n1078));
  OAI211_X1 g0878(.A(new_n923), .B(new_n856), .C1(new_n1077), .C2(new_n1078), .ZN(new_n1079));
  NAND2_X1  g0879(.A1(new_n1075), .A2(new_n1079), .ZN(new_n1080));
  NOR4_X1   g0880(.A1(new_n936), .A2(new_n1078), .A3(new_n699), .A4(new_n924), .ZN(new_n1081));
  NAND2_X1  g0881(.A1(new_n1080), .A2(new_n1081), .ZN(new_n1082));
  NAND4_X1  g0882(.A1(new_n922), .A2(G330), .A3(new_n834), .A4(new_n913), .ZN(new_n1083));
  NAND3_X1  g0883(.A1(new_n1075), .A2(new_n1083), .A3(new_n1079), .ZN(new_n1084));
  NAND2_X1  g0884(.A1(new_n1082), .A2(new_n1084), .ZN(new_n1085));
  NAND2_X1  g0885(.A1(new_n723), .A2(new_n568), .ZN(new_n1086));
  NAND2_X1  g0886(.A1(new_n918), .A2(new_n1086), .ZN(new_n1087));
  AOI21_X1  g0887(.A(new_n913), .B1(new_n723), .B2(new_n834), .ZN(new_n1088));
  OAI21_X1  g0888(.A(new_n909), .B1(new_n1088), .B2(new_n1081), .ZN(new_n1089));
  NOR3_X1   g0889(.A1(new_n936), .A2(new_n837), .A3(new_n699), .ZN(new_n1090));
  OAI211_X1 g0890(.A(new_n1083), .B(new_n1077), .C1(new_n1090), .C2(new_n913), .ZN(new_n1091));
  AOI21_X1  g0891(.A(new_n1087), .B1(new_n1089), .B2(new_n1091), .ZN(new_n1092));
  INV_X1    g0892(.A(new_n1092), .ZN(new_n1093));
  AOI21_X1  g0893(.A(new_n695), .B1(new_n1085), .B2(new_n1093), .ZN(new_n1094));
  NAND3_X1  g0894(.A1(new_n1082), .A2(new_n1092), .A3(new_n1084), .ZN(new_n1095));
  AND2_X1   g0895(.A1(new_n1094), .A2(new_n1095), .ZN(new_n1096));
  NAND3_X1  g0896(.A1(new_n898), .A2(new_n906), .A3(new_n739), .ZN(new_n1097));
  INV_X1    g0897(.A(new_n806), .ZN(new_n1098));
  OAI21_X1  g0898(.A(new_n735), .B1(new_n1014), .B2(new_n1098), .ZN(new_n1099));
  NOR2_X1   g0899(.A1(new_n821), .A2(new_n258), .ZN(new_n1100));
  AOI211_X1 g0900(.A(new_n1062), .B(new_n1100), .C1(G283), .C2(new_n774), .ZN(new_n1101));
  OAI22_X1  g0901(.A1(new_n784), .A2(new_n343), .B1(new_n780), .B2(new_n570), .ZN(new_n1102));
  AOI211_X1 g0902(.A(new_n269), .B(new_n1102), .C1(G116), .C2(new_n778), .ZN(new_n1103));
  NAND4_X1  g0903(.A1(new_n1101), .A2(new_n1103), .A3(new_n797), .A4(new_n816), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n762), .A2(G150), .ZN(new_n1105));
  XNOR2_X1  g0905(.A(new_n1105), .B(KEYINPUT53), .ZN(new_n1106));
  OAI22_X1  g0906(.A1(new_n821), .A2(new_n812), .B1(new_n793), .B2(new_n772), .ZN(new_n1107));
  AOI21_X1  g0907(.A(new_n1107), .B1(G128), .B2(new_n774), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n760), .A2(G50), .ZN(new_n1109));
  XOR2_X1   g0909(.A(KEYINPUT54), .B(G143), .Z(new_n1110));
  XNOR2_X1  g0910(.A(new_n1110), .B(KEYINPUT114), .ZN(new_n1111));
  NAND2_X1  g0911(.A1(new_n1111), .A2(new_n809), .ZN(new_n1112));
  AND2_X1   g0912(.A1(new_n781), .A2(G125), .ZN(new_n1113));
  AOI211_X1 g0913(.A(new_n370), .B(new_n1113), .C1(G132), .C2(new_n778), .ZN(new_n1114));
  NAND4_X1  g0914(.A1(new_n1108), .A2(new_n1109), .A3(new_n1112), .A4(new_n1114), .ZN(new_n1115));
  OAI21_X1  g0915(.A(new_n1104), .B1(new_n1106), .B2(new_n1115), .ZN(new_n1116));
  AOI21_X1  g0916(.A(new_n1099), .B1(new_n1116), .B2(new_n742), .ZN(new_n1117));
  NAND2_X1  g0917(.A1(new_n1097), .A2(new_n1117), .ZN(new_n1118));
  OAI21_X1  g0918(.A(new_n1118), .B1(new_n1085), .B2(new_n733), .ZN(new_n1119));
  NOR2_X1   g0919(.A1(new_n1096), .A2(new_n1119), .ZN(new_n1120));
  INV_X1    g0920(.A(new_n1120), .ZN(G378));
  OAI22_X1  g0921(.A1(new_n821), .A2(new_n343), .B1(new_n358), .B2(new_n784), .ZN(new_n1122));
  OAI22_X1  g0922(.A1(new_n1122), .A2(KEYINPUT115), .B1(new_n761), .B2(new_n201), .ZN(new_n1123));
  AOI21_X1  g0923(.A(new_n1123), .B1(KEYINPUT115), .B2(new_n1122), .ZN(new_n1124));
  NOR2_X1   g0924(.A1(new_n269), .A2(G41), .ZN(new_n1125));
  OAI221_X1 g0925(.A(new_n1125), .B1(new_n755), .B2(new_n780), .C1(new_n223), .C2(new_n777), .ZN(new_n1126));
  OAI22_X1  g0926(.A1(new_n775), .A2(new_n371), .B1(new_n202), .B2(new_n772), .ZN(new_n1127));
  NOR3_X1   g0927(.A1(new_n1021), .A2(new_n1126), .A3(new_n1127), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n1124), .A2(new_n1128), .ZN(new_n1129));
  XNOR2_X1  g0929(.A(new_n1129), .B(KEYINPUT116), .ZN(new_n1130));
  NAND2_X1  g0930(.A1(new_n1130), .A2(KEYINPUT58), .ZN(new_n1131));
  AOI211_X1 g0931(.A(G50), .B(new_n1125), .C1(new_n259), .C2(new_n302), .ZN(new_n1132));
  NAND2_X1  g0932(.A1(new_n1111), .A2(new_n762), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n767), .A2(G132), .ZN(new_n1134));
  AOI22_X1  g0934(.A1(new_n778), .A2(G128), .B1(new_n809), .B2(G137), .ZN(new_n1135));
  AOI22_X1  g0935(.A1(G150), .A2(new_n995), .B1(new_n774), .B2(G125), .ZN(new_n1136));
  NAND4_X1  g0936(.A1(new_n1133), .A2(new_n1134), .A3(new_n1135), .A4(new_n1136), .ZN(new_n1137));
  OR2_X1    g0937(.A1(new_n1137), .A2(KEYINPUT59), .ZN(new_n1138));
  AOI211_X1 g0938(.A(G33), .B(G41), .C1(new_n781), .C2(G124), .ZN(new_n1139));
  OAI21_X1  g0939(.A(new_n1139), .B1(new_n761), .B2(new_n793), .ZN(new_n1140));
  AOI21_X1  g0940(.A(new_n1140), .B1(new_n1137), .B2(KEYINPUT59), .ZN(new_n1141));
  AOI21_X1  g0941(.A(new_n1132), .B1(new_n1138), .B2(new_n1141), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n1131), .A2(new_n1142), .ZN(new_n1143));
  NOR2_X1   g0943(.A1(new_n1130), .A2(KEYINPUT58), .ZN(new_n1144));
  OAI21_X1  g0944(.A(new_n742), .B1(new_n1143), .B2(new_n1144), .ZN(new_n1145));
  AOI21_X1  g0945(.A(new_n738), .B1(new_n228), .B2(new_n806), .ZN(new_n1146));
  XOR2_X1   g0946(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1147));
  AOI211_X1 g0947(.A(new_n1147), .B(new_n457), .C1(new_n421), .C2(new_n423), .ZN(new_n1148));
  INV_X1    g0948(.A(new_n1147), .ZN(new_n1149));
  AOI21_X1  g0949(.A(new_n1149), .B1(new_n424), .B2(new_n456), .ZN(new_n1150));
  NOR2_X1   g0950(.A1(new_n1148), .A2(new_n1150), .ZN(new_n1151));
  NAND2_X1  g0951(.A1(new_n671), .A2(new_n416), .ZN(new_n1152));
  XOR2_X1   g0952(.A(new_n1152), .B(KEYINPUT117), .Z(new_n1153));
  NAND2_X1  g0953(.A1(new_n1151), .A2(new_n1153), .ZN(new_n1154));
  INV_X1    g0954(.A(new_n1153), .ZN(new_n1155));
  OAI21_X1  g0955(.A(new_n1155), .B1(new_n1148), .B2(new_n1150), .ZN(new_n1156));
  AND3_X1   g0956(.A1(new_n1154), .A2(KEYINPUT118), .A3(new_n1156), .ZN(new_n1157));
  AOI21_X1  g0957(.A(KEYINPUT118), .B1(new_n1154), .B2(new_n1156), .ZN(new_n1158));
  NOR2_X1   g0958(.A1(new_n1157), .A2(new_n1158), .ZN(new_n1159));
  OAI211_X1 g0959(.A(new_n1145), .B(new_n1146), .C1(new_n1159), .C2(new_n740), .ZN(new_n1160));
  INV_X1    g0960(.A(new_n1160), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n1154), .A2(new_n1156), .ZN(new_n1162));
  AOI21_X1  g0962(.A(new_n1162), .B1(new_n932), .B2(G330), .ZN(new_n1163));
  NOR3_X1   g0963(.A1(new_n934), .A2(new_n699), .A3(new_n1159), .ZN(new_n1164));
  OAI21_X1  g0964(.A(new_n917), .B1(new_n1163), .B2(new_n1164), .ZN(new_n1165));
  OR2_X1    g0965(.A1(new_n1157), .A2(new_n1158), .ZN(new_n1166));
  NAND3_X1  g0966(.A1(new_n932), .A2(G330), .A3(new_n1166), .ZN(new_n1167));
  INV_X1    g0967(.A(new_n1162), .ZN(new_n1168));
  OAI21_X1  g0968(.A(new_n1168), .B1(new_n934), .B2(new_n699), .ZN(new_n1169));
  OAI211_X1 g0969(.A(new_n1167), .B(new_n1169), .C1(new_n907), .C2(new_n916), .ZN(new_n1170));
  NAND2_X1  g0970(.A1(new_n1165), .A2(new_n1170), .ZN(new_n1171));
  AOI21_X1  g0971(.A(new_n1161), .B1(new_n1171), .B2(new_n734), .ZN(new_n1172));
  INV_X1    g0972(.A(new_n1172), .ZN(new_n1173));
  INV_X1    g0973(.A(KEYINPUT57), .ZN(new_n1174));
  AOI21_X1  g0974(.A(new_n1174), .B1(new_n1165), .B2(new_n1170), .ZN(new_n1175));
  INV_X1    g0975(.A(KEYINPUT119), .ZN(new_n1176));
  INV_X1    g0976(.A(new_n1087), .ZN(new_n1177));
  AND3_X1   g0977(.A1(new_n1095), .A2(new_n1176), .A3(new_n1177), .ZN(new_n1178));
  AOI21_X1  g0978(.A(new_n1176), .B1(new_n1095), .B2(new_n1177), .ZN(new_n1179));
  OAI21_X1  g0979(.A(new_n1175), .B1(new_n1178), .B2(new_n1179), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n1180), .A2(new_n694), .ZN(new_n1181));
  OAI21_X1  g0981(.A(new_n1171), .B1(new_n1178), .B2(new_n1179), .ZN(new_n1182));
  AOI22_X1  g0982(.A1(new_n1181), .A2(KEYINPUT120), .B1(new_n1174), .B2(new_n1182), .ZN(new_n1183));
  INV_X1    g0983(.A(KEYINPUT120), .ZN(new_n1184));
  NAND3_X1  g0984(.A1(new_n1180), .A2(new_n1184), .A3(new_n694), .ZN(new_n1185));
  AOI21_X1  g0985(.A(new_n1173), .B1(new_n1183), .B2(new_n1185), .ZN(new_n1186));
  INV_X1    g0986(.A(new_n1186), .ZN(G375));
  INV_X1    g0987(.A(new_n966), .ZN(new_n1188));
  NAND3_X1  g0988(.A1(new_n1089), .A2(new_n1091), .A3(new_n1087), .ZN(new_n1189));
  NAND3_X1  g0989(.A1(new_n1093), .A2(new_n1188), .A3(new_n1189), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n1089), .A2(new_n1091), .ZN(new_n1191));
  NAND2_X1  g0991(.A1(new_n1191), .A2(new_n734), .ZN(new_n1192));
  OAI21_X1  g0992(.A(new_n735), .B1(G68), .B2(new_n1098), .ZN(new_n1193));
  NAND2_X1  g0993(.A1(new_n1111), .A2(new_n767), .ZN(new_n1194));
  AOI21_X1  g0994(.A(new_n370), .B1(new_n781), .B2(G128), .ZN(new_n1195));
  AOI22_X1  g0995(.A1(G50), .A2(new_n995), .B1(new_n774), .B2(G132), .ZN(new_n1196));
  AOI22_X1  g0996(.A1(new_n778), .A2(G137), .B1(new_n809), .B2(G150), .ZN(new_n1197));
  NAND4_X1  g0997(.A1(new_n1194), .A2(new_n1195), .A3(new_n1196), .A4(new_n1197), .ZN(new_n1198));
  OAI22_X1  g0998(.A1(new_n201), .A2(new_n761), .B1(new_n763), .B2(new_n793), .ZN(new_n1199));
  OAI22_X1  g0999(.A1(new_n550), .A2(new_n761), .B1(new_n763), .B2(new_n343), .ZN(new_n1200));
  AOI22_X1  g1000(.A1(new_n360), .A2(new_n995), .B1(new_n774), .B2(G294), .ZN(new_n1201));
  AOI22_X1  g1001(.A1(new_n347), .A2(new_n809), .B1(G303), .B2(new_n781), .ZN(new_n1202));
  AOI21_X1  g1002(.A(new_n269), .B1(new_n778), .B2(G283), .ZN(new_n1203));
  NAND2_X1  g1003(.A1(new_n767), .A2(G116), .ZN(new_n1204));
  NAND4_X1  g1004(.A1(new_n1201), .A2(new_n1202), .A3(new_n1203), .A4(new_n1204), .ZN(new_n1205));
  OAI22_X1  g1005(.A1(new_n1198), .A2(new_n1199), .B1(new_n1200), .B2(new_n1205), .ZN(new_n1206));
  AOI21_X1  g1006(.A(new_n1193), .B1(new_n1206), .B2(new_n742), .ZN(new_n1207));
  OAI21_X1  g1007(.A(new_n1207), .B1(new_n913), .B2(new_n740), .ZN(new_n1208));
  NAND3_X1  g1008(.A1(new_n1190), .A2(new_n1192), .A3(new_n1208), .ZN(G381));
  INV_X1    g1009(.A(G390), .ZN(new_n1210));
  NAND3_X1  g1010(.A1(new_n1210), .A2(new_n984), .A3(new_n1008), .ZN(new_n1211));
  NOR2_X1   g1011(.A1(new_n1211), .A2(G381), .ZN(new_n1212));
  NOR3_X1   g1012(.A1(G393), .A2(G396), .A3(G384), .ZN(new_n1213));
  XNOR2_X1  g1013(.A(new_n1213), .B(KEYINPUT121), .ZN(new_n1214));
  NAND4_X1  g1014(.A1(new_n1212), .A2(new_n1120), .A3(new_n1186), .A4(new_n1214), .ZN(G407));
  NOR2_X1   g1015(.A1(new_n667), .A2(G343), .ZN(new_n1216));
  XNOR2_X1  g1016(.A(new_n1216), .B(KEYINPUT122), .ZN(new_n1217));
  NAND3_X1  g1017(.A1(new_n1186), .A2(new_n1120), .A3(new_n1217), .ZN(new_n1218));
  NAND3_X1  g1018(.A1(G407), .A2(G213), .A3(new_n1218), .ZN(G409));
  NAND2_X1  g1019(.A1(new_n1192), .A2(new_n1208), .ZN(new_n1220));
  NAND2_X1  g1020(.A1(new_n1093), .A2(KEYINPUT60), .ZN(new_n1221));
  NOR2_X1   g1021(.A1(new_n1221), .A2(new_n1189), .ZN(new_n1222));
  NOR2_X1   g1022(.A1(new_n1222), .A2(new_n695), .ZN(new_n1223));
  NAND2_X1  g1023(.A1(new_n1221), .A2(new_n1189), .ZN(new_n1224));
  AOI21_X1  g1024(.A(new_n1220), .B1(new_n1223), .B2(new_n1224), .ZN(new_n1225));
  OR2_X1    g1025(.A1(new_n1225), .A2(G384), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n1225), .A2(G384), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(new_n1226), .A2(new_n1227), .ZN(new_n1228));
  INV_X1    g1028(.A(G2897), .ZN(new_n1229));
  INV_X1    g1029(.A(new_n1216), .ZN(new_n1230));
  NOR3_X1   g1030(.A1(new_n1228), .A2(new_n1229), .A3(new_n1230), .ZN(new_n1231));
  AOI22_X1  g1031(.A1(new_n1226), .A2(new_n1227), .B1(G2897), .B2(new_n1217), .ZN(new_n1232));
  NOR2_X1   g1032(.A1(new_n1231), .A2(new_n1232), .ZN(new_n1233));
  INV_X1    g1033(.A(KEYINPUT124), .ZN(new_n1234));
  AOI21_X1  g1034(.A(new_n733), .B1(new_n1171), .B2(new_n1234), .ZN(new_n1235));
  NAND3_X1  g1035(.A1(new_n1165), .A2(new_n1170), .A3(KEYINPUT124), .ZN(new_n1236));
  AOI21_X1  g1036(.A(new_n1161), .B1(new_n1235), .B2(new_n1236), .ZN(new_n1237));
  OAI21_X1  g1037(.A(new_n1237), .B1(new_n1182), .B2(new_n966), .ZN(new_n1238));
  AND3_X1   g1038(.A1(new_n1238), .A2(KEYINPUT125), .A3(new_n1120), .ZN(new_n1239));
  AOI21_X1  g1039(.A(KEYINPUT125), .B1(new_n1238), .B2(new_n1120), .ZN(new_n1240));
  NOR2_X1   g1040(.A1(new_n1239), .A2(new_n1240), .ZN(new_n1241));
  INV_X1    g1041(.A(new_n1241), .ZN(new_n1242));
  INV_X1    g1042(.A(KEYINPUT123), .ZN(new_n1243));
  AOI21_X1  g1043(.A(new_n1243), .B1(new_n1186), .B2(G378), .ZN(new_n1244));
  NAND2_X1  g1044(.A1(new_n1171), .A2(KEYINPUT57), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n1095), .A2(new_n1177), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(new_n1246), .A2(KEYINPUT119), .ZN(new_n1247));
  NAND3_X1  g1047(.A1(new_n1095), .A2(new_n1176), .A3(new_n1177), .ZN(new_n1248));
  AOI21_X1  g1048(.A(new_n1245), .B1(new_n1247), .B2(new_n1248), .ZN(new_n1249));
  OAI21_X1  g1049(.A(KEYINPUT120), .B1(new_n1249), .B2(new_n695), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(new_n1182), .A2(new_n1174), .ZN(new_n1251));
  NAND3_X1  g1051(.A1(new_n1250), .A2(new_n1185), .A3(new_n1251), .ZN(new_n1252));
  NAND4_X1  g1052(.A1(new_n1252), .A2(new_n1243), .A3(G378), .A4(new_n1172), .ZN(new_n1253));
  INV_X1    g1053(.A(new_n1253), .ZN(new_n1254));
  OAI21_X1  g1054(.A(new_n1242), .B1(new_n1244), .B2(new_n1254), .ZN(new_n1255));
  INV_X1    g1055(.A(new_n1217), .ZN(new_n1256));
  AOI21_X1  g1056(.A(new_n1233), .B1(new_n1255), .B2(new_n1256), .ZN(new_n1257));
  XOR2_X1   g1057(.A(KEYINPUT126), .B(KEYINPUT61), .Z(new_n1258));
  OAI21_X1  g1058(.A(KEYINPUT127), .B1(new_n1257), .B2(new_n1258), .ZN(new_n1259));
  INV_X1    g1059(.A(KEYINPUT127), .ZN(new_n1260));
  INV_X1    g1060(.A(new_n1258), .ZN(new_n1261));
  NAND3_X1  g1061(.A1(new_n1252), .A2(G378), .A3(new_n1172), .ZN(new_n1262));
  NAND2_X1  g1062(.A1(new_n1262), .A2(KEYINPUT123), .ZN(new_n1263));
  AOI21_X1  g1063(.A(new_n1241), .B1(new_n1263), .B2(new_n1253), .ZN(new_n1264));
  NOR2_X1   g1064(.A1(new_n1264), .A2(new_n1217), .ZN(new_n1265));
  OAI211_X1 g1065(.A(new_n1260), .B(new_n1261), .C1(new_n1265), .C2(new_n1233), .ZN(new_n1266));
  INV_X1    g1066(.A(new_n1228), .ZN(new_n1267));
  AND2_X1   g1067(.A1(new_n1267), .A2(KEYINPUT62), .ZN(new_n1268));
  NAND3_X1  g1068(.A1(new_n1255), .A2(new_n1256), .A3(new_n1268), .ZN(new_n1269));
  NOR3_X1   g1069(.A1(new_n1264), .A2(new_n1216), .A3(new_n1228), .ZN(new_n1270));
  OAI21_X1  g1070(.A(new_n1269), .B1(new_n1270), .B2(KEYINPUT62), .ZN(new_n1271));
  NAND3_X1  g1071(.A1(new_n1259), .A2(new_n1266), .A3(new_n1271), .ZN(new_n1272));
  NAND2_X1  g1072(.A1(G387), .A2(G390), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(new_n1273), .A2(new_n1211), .ZN(new_n1274));
  XNOR2_X1  g1074(.A(G393), .B(new_n804), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(new_n1274), .A2(new_n1275), .ZN(new_n1276));
  INV_X1    g1076(.A(new_n1275), .ZN(new_n1277));
  NAND3_X1  g1077(.A1(new_n1273), .A2(new_n1211), .A3(new_n1277), .ZN(new_n1278));
  NAND2_X1  g1078(.A1(new_n1276), .A2(new_n1278), .ZN(new_n1279));
  NAND2_X1  g1079(.A1(new_n1272), .A2(new_n1279), .ZN(new_n1280));
  INV_X1    g1080(.A(KEYINPUT61), .ZN(new_n1281));
  AND3_X1   g1081(.A1(new_n1276), .A2(new_n1281), .A3(new_n1278), .ZN(new_n1282));
  OR2_X1    g1082(.A1(new_n1270), .A2(KEYINPUT63), .ZN(new_n1283));
  NAND3_X1  g1083(.A1(new_n1265), .A2(KEYINPUT63), .A3(new_n1267), .ZN(new_n1284));
  OAI22_X1  g1084(.A1(new_n1264), .A2(new_n1216), .B1(new_n1232), .B2(new_n1231), .ZN(new_n1285));
  NAND4_X1  g1085(.A1(new_n1282), .A2(new_n1283), .A3(new_n1284), .A4(new_n1285), .ZN(new_n1286));
  NAND2_X1  g1086(.A1(new_n1280), .A2(new_n1286), .ZN(G405));
  NOR2_X1   g1087(.A1(new_n1244), .A2(new_n1254), .ZN(new_n1288));
  NOR2_X1   g1088(.A1(new_n1186), .A2(G378), .ZN(new_n1289));
  NOR2_X1   g1089(.A1(new_n1288), .A2(new_n1289), .ZN(new_n1290));
  XNOR2_X1  g1090(.A(new_n1290), .B(new_n1228), .ZN(new_n1291));
  XNOR2_X1  g1091(.A(new_n1291), .B(new_n1279), .ZN(G402));
endmodule


