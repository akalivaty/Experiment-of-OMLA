//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 0 1 0 0 0 1 1 0 0 1 1 1 1 0 1 0 1 0 1 0 0 1 1 0 0 0 0 0 0 0 1 1 1 1 0 0 0 1 1 1 0 1 0 0 0 0 1 1 0 1 1 0 0 0 0 0 0 1 0 0 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:30:47 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n447, new_n449, new_n452, new_n453, new_n454, new_n455,
    new_n458, new_n459, new_n460, new_n461, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n533, new_n534, new_n535, new_n537, new_n538, new_n539,
    new_n540, new_n541, new_n542, new_n543, new_n544, new_n546, new_n547,
    new_n548, new_n549, new_n552, new_n553, new_n554, new_n555, new_n556,
    new_n557, new_n560, new_n561, new_n563, new_n564, new_n565, new_n566,
    new_n567, new_n568, new_n569, new_n570, new_n571, new_n573, new_n574,
    new_n575, new_n578, new_n579, new_n580, new_n581, new_n583, new_n584,
    new_n585, new_n586, new_n587, new_n588, new_n589, new_n590, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n614, new_n616, new_n617, new_n618, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1211, new_n1212, new_n1213, new_n1214,
    new_n1215, new_n1216, new_n1217, new_n1218;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  XNOR2_X1  g015(.A(KEYINPUT64), .B(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  XOR2_X1   g018(.A(KEYINPUT65), .B(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  XNOR2_X1  g020(.A(KEYINPUT66), .B(KEYINPUT1), .ZN(new_n446));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XNOR2_X1  g022(.A(new_n446), .B(new_n447), .ZN(G223));
  INV_X1    g023(.A(new_n447), .ZN(new_n449));
  NAND2_X1  g024(.A1(new_n449), .A2(G567), .ZN(G234));
  NAND2_X1  g025(.A1(new_n449), .A2(G2106), .ZN(G217));
  NOR4_X1   g026(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n452));
  XNOR2_X1  g027(.A(new_n452), .B(KEYINPUT2), .ZN(new_n453));
  NOR4_X1   g028(.A1(G238), .A2(G237), .A3(G235), .A4(G236), .ZN(new_n454));
  NAND2_X1  g029(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  INV_X1    g030(.A(new_n455), .ZN(G325));
  XNOR2_X1  g031(.A(new_n455), .B(KEYINPUT67), .ZN(G261));
  INV_X1    g032(.A(new_n453), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n458), .A2(G2106), .ZN(new_n459));
  INV_X1    g034(.A(G567), .ZN(new_n460));
  OAI22_X1  g035(.A1(new_n459), .A2(KEYINPUT68), .B1(new_n460), .B2(new_n454), .ZN(new_n461));
  AOI21_X1  g036(.A(new_n461), .B1(KEYINPUT68), .B2(new_n459), .ZN(G319));
  INV_X1    g037(.A(G2105), .ZN(new_n463));
  OR2_X1    g038(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n464));
  INV_X1    g039(.A(KEYINPUT69), .ZN(new_n465));
  NAND2_X1  g040(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n466));
  NAND3_X1  g041(.A1(new_n464), .A2(new_n465), .A3(new_n466), .ZN(new_n467));
  AND2_X1   g042(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n468));
  NOR2_X1   g043(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n469));
  OAI21_X1  g044(.A(KEYINPUT69), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  NAND3_X1  g045(.A1(new_n467), .A2(new_n470), .A3(G125), .ZN(new_n471));
  NAND2_X1  g046(.A1(G113), .A2(G2104), .ZN(new_n472));
  XOR2_X1   g047(.A(new_n472), .B(KEYINPUT70), .Z(new_n473));
  AOI21_X1  g048(.A(new_n463), .B1(new_n471), .B2(new_n473), .ZN(new_n474));
  INV_X1    g049(.A(G2104), .ZN(new_n475));
  NOR2_X1   g050(.A1(new_n475), .A2(G2105), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n476), .A2(G101), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n464), .A2(new_n466), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n478), .A2(new_n463), .ZN(new_n479));
  INV_X1    g054(.A(G137), .ZN(new_n480));
  OAI21_X1  g055(.A(new_n477), .B1(new_n479), .B2(new_n480), .ZN(new_n481));
  NOR2_X1   g056(.A1(new_n474), .A2(new_n481), .ZN(new_n482));
  XNOR2_X1  g057(.A(new_n482), .B(KEYINPUT71), .ZN(G160));
  INV_X1    g058(.A(new_n479), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n484), .A2(G136), .ZN(new_n485));
  AOI21_X1  g060(.A(new_n463), .B1(new_n464), .B2(new_n466), .ZN(new_n486));
  NAND2_X1  g061(.A1(new_n486), .A2(G124), .ZN(new_n487));
  OR2_X1    g062(.A1(G100), .A2(G2105), .ZN(new_n488));
  OAI211_X1 g063(.A(new_n488), .B(G2104), .C1(G112), .C2(new_n463), .ZN(new_n489));
  NAND3_X1  g064(.A1(new_n485), .A2(new_n487), .A3(new_n489), .ZN(new_n490));
  INV_X1    g065(.A(new_n490), .ZN(G162));
  NOR2_X1   g066(.A1(new_n463), .A2(G114), .ZN(new_n492));
  OAI21_X1  g067(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n493));
  OR3_X1    g068(.A1(new_n492), .A2(new_n493), .A3(KEYINPUT72), .ZN(new_n494));
  OAI21_X1  g069(.A(KEYINPUT72), .B1(new_n492), .B2(new_n493), .ZN(new_n495));
  AOI22_X1  g070(.A1(new_n494), .A2(new_n495), .B1(G126), .B2(new_n486), .ZN(new_n496));
  OAI211_X1 g071(.A(G138), .B(new_n463), .C1(new_n468), .C2(new_n469), .ZN(new_n497));
  NAND2_X1  g072(.A1(new_n497), .A2(KEYINPUT4), .ZN(new_n498));
  NAND2_X1  g073(.A1(new_n467), .A2(new_n470), .ZN(new_n499));
  INV_X1    g074(.A(KEYINPUT4), .ZN(new_n500));
  NAND3_X1  g075(.A1(new_n500), .A2(new_n463), .A3(G138), .ZN(new_n501));
  OAI21_X1  g076(.A(new_n498), .B1(new_n499), .B2(new_n501), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n496), .A2(new_n502), .ZN(new_n503));
  INV_X1    g078(.A(new_n503), .ZN(G164));
  INV_X1    g079(.A(KEYINPUT73), .ZN(new_n505));
  INV_X1    g080(.A(KEYINPUT6), .ZN(new_n506));
  OAI21_X1  g081(.A(new_n505), .B1(new_n506), .B2(G651), .ZN(new_n507));
  INV_X1    g082(.A(G651), .ZN(new_n508));
  NAND3_X1  g083(.A1(new_n508), .A2(KEYINPUT73), .A3(KEYINPUT6), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n507), .A2(new_n509), .ZN(new_n510));
  INV_X1    g085(.A(KEYINPUT74), .ZN(new_n511));
  OAI21_X1  g086(.A(new_n511), .B1(new_n508), .B2(KEYINPUT6), .ZN(new_n512));
  NAND3_X1  g087(.A1(new_n506), .A2(KEYINPUT74), .A3(G651), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n510), .A2(new_n514), .ZN(new_n515));
  INV_X1    g090(.A(KEYINPUT5), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n516), .A2(G543), .ZN(new_n517));
  INV_X1    g092(.A(KEYINPUT75), .ZN(new_n518));
  INV_X1    g093(.A(G543), .ZN(new_n519));
  AOI21_X1  g094(.A(new_n518), .B1(KEYINPUT5), .B2(new_n519), .ZN(new_n520));
  NOR3_X1   g095(.A1(new_n516), .A2(KEYINPUT75), .A3(G543), .ZN(new_n521));
  OAI21_X1  g096(.A(new_n517), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  NOR2_X1   g097(.A1(new_n515), .A2(new_n522), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n523), .A2(G88), .ZN(new_n524));
  INV_X1    g099(.A(G50), .ZN(new_n525));
  NOR2_X1   g100(.A1(new_n515), .A2(new_n519), .ZN(new_n526));
  INV_X1    g101(.A(new_n526), .ZN(new_n527));
  OAI21_X1  g102(.A(new_n524), .B1(new_n525), .B2(new_n527), .ZN(new_n528));
  OAI21_X1  g103(.A(KEYINPUT75), .B1(new_n516), .B2(G543), .ZN(new_n529));
  NAND3_X1  g104(.A1(new_n518), .A2(new_n519), .A3(KEYINPUT5), .ZN(new_n530));
  AOI22_X1  g105(.A1(new_n529), .A2(new_n530), .B1(new_n516), .B2(G543), .ZN(new_n531));
  NAND2_X1  g106(.A1(new_n531), .A2(G62), .ZN(new_n532));
  NAND2_X1  g107(.A1(G75), .A2(G543), .ZN(new_n533));
  XNOR2_X1  g108(.A(new_n533), .B(KEYINPUT76), .ZN(new_n534));
  AOI21_X1  g109(.A(new_n508), .B1(new_n532), .B2(new_n534), .ZN(new_n535));
  NOR2_X1   g110(.A1(new_n528), .A2(new_n535), .ZN(G166));
  NAND2_X1  g111(.A1(new_n523), .A2(G89), .ZN(new_n537));
  NAND4_X1  g112(.A1(new_n510), .A2(new_n514), .A3(G51), .A4(G543), .ZN(new_n538));
  AND2_X1   g113(.A1(G63), .A2(G651), .ZN(new_n539));
  NAND3_X1  g114(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n540));
  NAND2_X1  g115(.A1(new_n540), .A2(KEYINPUT7), .ZN(new_n541));
  OR2_X1    g116(.A1(new_n540), .A2(KEYINPUT7), .ZN(new_n542));
  AOI22_X1  g117(.A1(new_n531), .A2(new_n539), .B1(new_n541), .B2(new_n542), .ZN(new_n543));
  NAND3_X1  g118(.A1(new_n537), .A2(new_n538), .A3(new_n543), .ZN(new_n544));
  INV_X1    g119(.A(new_n544), .ZN(G168));
  AOI22_X1  g120(.A1(new_n531), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n546));
  OR2_X1    g121(.A1(new_n546), .A2(new_n508), .ZN(new_n547));
  NAND2_X1  g122(.A1(new_n526), .A2(G52), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n523), .A2(G90), .ZN(new_n549));
  NAND3_X1  g124(.A1(new_n547), .A2(new_n548), .A3(new_n549), .ZN(G301));
  INV_X1    g125(.A(G301), .ZN(G171));
  AOI22_X1  g126(.A1(new_n531), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n552));
  OR2_X1    g127(.A1(new_n552), .A2(new_n508), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n526), .A2(G43), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n523), .A2(G81), .ZN(new_n555));
  NAND3_X1  g130(.A1(new_n553), .A2(new_n554), .A3(new_n555), .ZN(new_n556));
  INV_X1    g131(.A(new_n556), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n557), .A2(G860), .ZN(G153));
  NAND4_X1  g133(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g134(.A1(G1), .A2(G3), .ZN(new_n560));
  XNOR2_X1  g135(.A(new_n560), .B(KEYINPUT8), .ZN(new_n561));
  NAND4_X1  g136(.A1(G319), .A2(G483), .A3(G661), .A4(new_n561), .ZN(G188));
  NAND4_X1  g137(.A1(new_n510), .A2(new_n514), .A3(G53), .A4(G543), .ZN(new_n563));
  XNOR2_X1  g138(.A(new_n563), .B(KEYINPUT9), .ZN(new_n564));
  XNOR2_X1  g139(.A(KEYINPUT78), .B(G65), .ZN(new_n565));
  AOI22_X1  g140(.A1(new_n531), .A2(new_n565), .B1(G78), .B2(G543), .ZN(new_n566));
  OR2_X1    g141(.A1(new_n566), .A2(new_n508), .ZN(new_n567));
  OAI21_X1  g142(.A(KEYINPUT77), .B1(new_n515), .B2(new_n522), .ZN(new_n568));
  INV_X1    g143(.A(KEYINPUT77), .ZN(new_n569));
  NAND4_X1  g144(.A1(new_n531), .A2(new_n569), .A3(new_n510), .A4(new_n514), .ZN(new_n570));
  NAND3_X1  g145(.A1(new_n568), .A2(G91), .A3(new_n570), .ZN(new_n571));
  NAND3_X1  g146(.A1(new_n564), .A2(new_n567), .A3(new_n571), .ZN(G299));
  NAND2_X1  g147(.A1(new_n544), .A2(KEYINPUT79), .ZN(new_n573));
  INV_X1    g148(.A(KEYINPUT79), .ZN(new_n574));
  NAND4_X1  g149(.A1(new_n537), .A2(new_n574), .A3(new_n538), .A4(new_n543), .ZN(new_n575));
  AND2_X1   g150(.A1(new_n573), .A2(new_n575), .ZN(G286));
  INV_X1    g151(.A(G166), .ZN(G303));
  OAI21_X1  g152(.A(G651), .B1(new_n531), .B2(G74), .ZN(new_n578));
  XNOR2_X1  g153(.A(new_n578), .B(KEYINPUT80), .ZN(new_n579));
  NAND3_X1  g154(.A1(new_n568), .A2(G87), .A3(new_n570), .ZN(new_n580));
  NAND2_X1  g155(.A1(new_n526), .A2(G49), .ZN(new_n581));
  NAND3_X1  g156(.A1(new_n579), .A2(new_n580), .A3(new_n581), .ZN(G288));
  NAND2_X1  g157(.A1(G73), .A2(G543), .ZN(new_n583));
  INV_X1    g158(.A(G61), .ZN(new_n584));
  OAI21_X1  g159(.A(new_n583), .B1(new_n522), .B2(new_n584), .ZN(new_n585));
  AOI22_X1  g160(.A1(G651), .A2(new_n585), .B1(new_n526), .B2(G48), .ZN(new_n586));
  INV_X1    g161(.A(KEYINPUT81), .ZN(new_n587));
  NAND3_X1  g162(.A1(new_n568), .A2(G86), .A3(new_n570), .ZN(new_n588));
  AND3_X1   g163(.A1(new_n586), .A2(new_n587), .A3(new_n588), .ZN(new_n589));
  AOI21_X1  g164(.A(new_n587), .B1(new_n586), .B2(new_n588), .ZN(new_n590));
  NOR2_X1   g165(.A1(new_n589), .A2(new_n590), .ZN(G305));
  AND2_X1   g166(.A1(new_n531), .A2(G60), .ZN(new_n592));
  AND2_X1   g167(.A1(G72), .A2(G543), .ZN(new_n593));
  OAI21_X1  g168(.A(G651), .B1(new_n592), .B2(new_n593), .ZN(new_n594));
  INV_X1    g169(.A(KEYINPUT82), .ZN(new_n595));
  OR2_X1    g170(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  NAND2_X1  g171(.A1(new_n594), .A2(new_n595), .ZN(new_n597));
  AOI22_X1  g172(.A1(G47), .A2(new_n526), .B1(new_n523), .B2(G85), .ZN(new_n598));
  AND3_X1   g173(.A1(new_n596), .A2(new_n597), .A3(new_n598), .ZN(new_n599));
  INV_X1    g174(.A(new_n599), .ZN(G290));
  NAND2_X1  g175(.A1(G301), .A2(G868), .ZN(new_n601));
  NAND2_X1  g176(.A1(new_n526), .A2(G54), .ZN(new_n602));
  AOI22_X1  g177(.A1(new_n531), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n603));
  OAI21_X1  g178(.A(new_n602), .B1(new_n508), .B2(new_n603), .ZN(new_n604));
  NAND3_X1  g179(.A1(new_n568), .A2(G92), .A3(new_n570), .ZN(new_n605));
  INV_X1    g180(.A(KEYINPUT10), .ZN(new_n606));
  NAND2_X1  g181(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  NAND4_X1  g182(.A1(new_n568), .A2(KEYINPUT10), .A3(G92), .A4(new_n570), .ZN(new_n608));
  AOI21_X1  g183(.A(new_n604), .B1(new_n607), .B2(new_n608), .ZN(new_n609));
  OAI21_X1  g184(.A(new_n601), .B1(new_n609), .B2(G868), .ZN(G321));
  XOR2_X1   g185(.A(G321), .B(KEYINPUT83), .Z(G284));
  MUX2_X1   g186(.A(G299), .B(G286), .S(G868), .Z(G297));
  MUX2_X1   g187(.A(G299), .B(G286), .S(G868), .Z(G280));
  XOR2_X1   g188(.A(KEYINPUT84), .B(G559), .Z(new_n614));
  OAI21_X1  g189(.A(new_n609), .B1(G860), .B2(new_n614), .ZN(G148));
  INV_X1    g190(.A(G868), .ZN(new_n616));
  NAND2_X1  g191(.A1(new_n556), .A2(new_n616), .ZN(new_n617));
  AND2_X1   g192(.A1(new_n609), .A2(new_n614), .ZN(new_n618));
  OAI21_X1  g193(.A(new_n617), .B1(new_n618), .B2(new_n616), .ZN(G323));
  XNOR2_X1  g194(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NOR3_X1   g195(.A1(new_n499), .A2(new_n475), .A3(G2105), .ZN(new_n621));
  INV_X1    g196(.A(KEYINPUT12), .ZN(new_n622));
  OR2_X1    g197(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  NAND2_X1  g198(.A1(new_n621), .A2(new_n622), .ZN(new_n624));
  NAND2_X1  g199(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  XNOR2_X1  g200(.A(new_n625), .B(KEYINPUT13), .ZN(new_n626));
  INV_X1    g201(.A(G2100), .ZN(new_n627));
  OR2_X1    g202(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  NAND2_X1  g203(.A1(new_n626), .A2(new_n627), .ZN(new_n629));
  NAND2_X1  g204(.A1(new_n484), .A2(G135), .ZN(new_n630));
  OR3_X1    g205(.A1(new_n463), .A2(KEYINPUT85), .A3(G111), .ZN(new_n631));
  OAI21_X1  g206(.A(KEYINPUT85), .B1(new_n463), .B2(G111), .ZN(new_n632));
  OR2_X1    g207(.A1(G99), .A2(G2105), .ZN(new_n633));
  NAND4_X1  g208(.A1(new_n631), .A2(G2104), .A3(new_n632), .A4(new_n633), .ZN(new_n634));
  NAND2_X1  g209(.A1(new_n486), .A2(G123), .ZN(new_n635));
  NAND3_X1  g210(.A1(new_n630), .A2(new_n634), .A3(new_n635), .ZN(new_n636));
  XOR2_X1   g211(.A(new_n636), .B(G2096), .Z(new_n637));
  NAND3_X1  g212(.A1(new_n628), .A2(new_n629), .A3(new_n637), .ZN(G156));
  XNOR2_X1  g213(.A(G2451), .B(G2454), .ZN(new_n639));
  XNOR2_X1  g214(.A(G2443), .B(G2446), .ZN(new_n640));
  XNOR2_X1  g215(.A(new_n639), .B(new_n640), .ZN(new_n641));
  XNOR2_X1  g216(.A(KEYINPUT86), .B(KEYINPUT16), .ZN(new_n642));
  XNOR2_X1  g217(.A(new_n641), .B(new_n642), .ZN(new_n643));
  XNOR2_X1  g218(.A(G1341), .B(G1348), .ZN(new_n644));
  XNOR2_X1  g219(.A(new_n644), .B(KEYINPUT88), .ZN(new_n645));
  XNOR2_X1  g220(.A(new_n645), .B(KEYINPUT87), .ZN(new_n646));
  XNOR2_X1  g221(.A(new_n643), .B(new_n646), .ZN(new_n647));
  INV_X1    g222(.A(new_n647), .ZN(new_n648));
  XNOR2_X1  g223(.A(G2427), .B(G2438), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n649), .B(G2430), .ZN(new_n650));
  XNOR2_X1  g225(.A(KEYINPUT15), .B(G2435), .ZN(new_n651));
  OR2_X1    g226(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  NAND2_X1  g227(.A1(new_n650), .A2(new_n651), .ZN(new_n653));
  NAND3_X1  g228(.A1(new_n652), .A2(new_n653), .A3(KEYINPUT14), .ZN(new_n654));
  OR2_X1    g229(.A1(new_n648), .A2(new_n654), .ZN(new_n655));
  NAND2_X1  g230(.A1(new_n648), .A2(new_n654), .ZN(new_n656));
  NAND3_X1  g231(.A1(new_n655), .A2(G14), .A3(new_n656), .ZN(new_n657));
  INV_X1    g232(.A(new_n657), .ZN(G401));
  XNOR2_X1  g233(.A(G2072), .B(G2078), .ZN(new_n659));
  XOR2_X1   g234(.A(new_n659), .B(KEYINPUT17), .Z(new_n660));
  XNOR2_X1  g235(.A(G2067), .B(G2678), .ZN(new_n661));
  INV_X1    g236(.A(new_n661), .ZN(new_n662));
  NOR2_X1   g237(.A1(new_n660), .A2(new_n662), .ZN(new_n663));
  XNOR2_X1  g238(.A(G2084), .B(G2090), .ZN(new_n664));
  OAI21_X1  g239(.A(new_n664), .B1(new_n661), .B2(new_n659), .ZN(new_n665));
  NOR2_X1   g240(.A1(new_n663), .A2(new_n665), .ZN(new_n666));
  XNOR2_X1  g241(.A(new_n666), .B(KEYINPUT89), .ZN(new_n667));
  INV_X1    g242(.A(new_n664), .ZN(new_n668));
  NAND3_X1  g243(.A1(new_n668), .A2(new_n661), .A3(new_n659), .ZN(new_n669));
  XNOR2_X1  g244(.A(new_n669), .B(KEYINPUT18), .ZN(new_n670));
  NOR2_X1   g245(.A1(new_n661), .A2(new_n664), .ZN(new_n671));
  AOI21_X1  g246(.A(new_n670), .B1(new_n660), .B2(new_n671), .ZN(new_n672));
  NAND2_X1  g247(.A1(new_n667), .A2(new_n672), .ZN(new_n673));
  XNOR2_X1  g248(.A(G2096), .B(G2100), .ZN(new_n674));
  XNOR2_X1  g249(.A(new_n673), .B(new_n674), .ZN(new_n675));
  INV_X1    g250(.A(new_n675), .ZN(G227));
  XNOR2_X1  g251(.A(G1981), .B(G1986), .ZN(new_n677));
  XNOR2_X1  g252(.A(new_n677), .B(KEYINPUT95), .ZN(new_n678));
  XNOR2_X1  g253(.A(G1971), .B(G1976), .ZN(new_n679));
  XNOR2_X1  g254(.A(KEYINPUT90), .B(KEYINPUT19), .ZN(new_n680));
  XNOR2_X1  g255(.A(new_n679), .B(new_n680), .ZN(new_n681));
  XNOR2_X1  g256(.A(G1961), .B(G1966), .ZN(new_n682));
  INV_X1    g257(.A(KEYINPUT91), .ZN(new_n683));
  XNOR2_X1  g258(.A(new_n682), .B(new_n683), .ZN(new_n684));
  XNOR2_X1  g259(.A(G1956), .B(G2474), .ZN(new_n685));
  NAND3_X1  g260(.A1(new_n681), .A2(new_n684), .A3(new_n685), .ZN(new_n686));
  INV_X1    g261(.A(KEYINPUT92), .ZN(new_n687));
  NAND2_X1  g262(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  NAND4_X1  g263(.A1(new_n681), .A2(new_n684), .A3(KEYINPUT92), .A4(new_n685), .ZN(new_n689));
  AOI21_X1  g264(.A(new_n681), .B1(new_n684), .B2(new_n685), .ZN(new_n690));
  XNOR2_X1  g265(.A(new_n682), .B(KEYINPUT91), .ZN(new_n691));
  INV_X1    g266(.A(new_n685), .ZN(new_n692));
  NAND2_X1  g267(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  AOI22_X1  g268(.A1(new_n688), .A2(new_n689), .B1(new_n690), .B2(new_n693), .ZN(new_n694));
  NAND3_X1  g269(.A1(new_n681), .A2(new_n691), .A3(new_n692), .ZN(new_n695));
  XNOR2_X1  g270(.A(new_n695), .B(KEYINPUT20), .ZN(new_n696));
  NAND3_X1  g271(.A1(new_n694), .A2(new_n696), .A3(KEYINPUT93), .ZN(new_n697));
  INV_X1    g272(.A(new_n697), .ZN(new_n698));
  AOI21_X1  g273(.A(KEYINPUT93), .B1(new_n694), .B2(new_n696), .ZN(new_n699));
  NOR3_X1   g274(.A1(new_n698), .A2(new_n699), .A3(KEYINPUT94), .ZN(new_n700));
  INV_X1    g275(.A(KEYINPUT94), .ZN(new_n701));
  NAND2_X1  g276(.A1(new_n694), .A2(new_n696), .ZN(new_n702));
  INV_X1    g277(.A(KEYINPUT93), .ZN(new_n703));
  NAND2_X1  g278(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  AOI21_X1  g279(.A(new_n701), .B1(new_n704), .B2(new_n697), .ZN(new_n705));
  OAI21_X1  g280(.A(new_n678), .B1(new_n700), .B2(new_n705), .ZN(new_n706));
  XOR2_X1   g281(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n707));
  XNOR2_X1  g282(.A(G1991), .B(G1996), .ZN(new_n708));
  XOR2_X1   g283(.A(new_n707), .B(new_n708), .Z(new_n709));
  OAI21_X1  g284(.A(KEYINPUT94), .B1(new_n698), .B2(new_n699), .ZN(new_n710));
  NAND3_X1  g285(.A1(new_n704), .A2(new_n701), .A3(new_n697), .ZN(new_n711));
  INV_X1    g286(.A(new_n678), .ZN(new_n712));
  NAND3_X1  g287(.A1(new_n710), .A2(new_n711), .A3(new_n712), .ZN(new_n713));
  AND3_X1   g288(.A1(new_n706), .A2(new_n709), .A3(new_n713), .ZN(new_n714));
  AOI21_X1  g289(.A(new_n709), .B1(new_n706), .B2(new_n713), .ZN(new_n715));
  NOR2_X1   g290(.A1(new_n714), .A2(new_n715), .ZN(G229));
  INV_X1    g291(.A(G16), .ZN(new_n717));
  NAND2_X1  g292(.A1(new_n717), .A2(G24), .ZN(new_n718));
  OAI21_X1  g293(.A(new_n718), .B1(new_n599), .B2(new_n717), .ZN(new_n719));
  XOR2_X1   g294(.A(new_n719), .B(KEYINPUT97), .Z(new_n720));
  INV_X1    g295(.A(G1986), .ZN(new_n721));
  AND2_X1   g296(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  NOR2_X1   g297(.A1(new_n720), .A2(new_n721), .ZN(new_n723));
  NOR2_X1   g298(.A1(G25), .A2(G29), .ZN(new_n724));
  NAND2_X1  g299(.A1(new_n484), .A2(G131), .ZN(new_n725));
  NAND2_X1  g300(.A1(new_n486), .A2(G119), .ZN(new_n726));
  OR2_X1    g301(.A1(G95), .A2(G2105), .ZN(new_n727));
  OAI211_X1 g302(.A(new_n727), .B(G2104), .C1(G107), .C2(new_n463), .ZN(new_n728));
  NAND3_X1  g303(.A1(new_n725), .A2(new_n726), .A3(new_n728), .ZN(new_n729));
  INV_X1    g304(.A(new_n729), .ZN(new_n730));
  AOI21_X1  g305(.A(new_n724), .B1(new_n730), .B2(G29), .ZN(new_n731));
  XNOR2_X1  g306(.A(new_n731), .B(KEYINPUT96), .ZN(new_n732));
  XOR2_X1   g307(.A(KEYINPUT35), .B(G1991), .Z(new_n733));
  XOR2_X1   g308(.A(new_n732), .B(new_n733), .Z(new_n734));
  NOR3_X1   g309(.A1(new_n722), .A2(new_n723), .A3(new_n734), .ZN(new_n735));
  NAND2_X1  g310(.A1(new_n717), .A2(G22), .ZN(new_n736));
  OAI21_X1  g311(.A(new_n736), .B1(G166), .B2(new_n717), .ZN(new_n737));
  XNOR2_X1  g312(.A(new_n737), .B(G1971), .ZN(new_n738));
  NAND2_X1  g313(.A1(new_n717), .A2(G23), .ZN(new_n739));
  INV_X1    g314(.A(G288), .ZN(new_n740));
  OAI21_X1  g315(.A(new_n739), .B1(new_n740), .B2(new_n717), .ZN(new_n741));
  XOR2_X1   g316(.A(KEYINPUT33), .B(G1976), .Z(new_n742));
  NOR2_X1   g317(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  NOR2_X1   g318(.A1(new_n738), .A2(new_n743), .ZN(new_n744));
  NAND2_X1  g319(.A1(new_n741), .A2(new_n742), .ZN(new_n745));
  NAND2_X1  g320(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  MUX2_X1   g321(.A(G6), .B(G305), .S(G16), .Z(new_n747));
  XNOR2_X1  g322(.A(KEYINPUT32), .B(G1981), .ZN(new_n748));
  XNOR2_X1  g323(.A(new_n747), .B(new_n748), .ZN(new_n749));
  OR3_X1    g324(.A1(new_n746), .A2(new_n749), .A3(KEYINPUT34), .ZN(new_n750));
  NAND2_X1  g325(.A1(new_n735), .A2(new_n750), .ZN(new_n751));
  OAI21_X1  g326(.A(KEYINPUT34), .B1(new_n746), .B2(new_n749), .ZN(new_n752));
  INV_X1    g327(.A(new_n752), .ZN(new_n753));
  OAI21_X1  g328(.A(KEYINPUT36), .B1(new_n751), .B2(new_n753), .ZN(new_n754));
  INV_X1    g329(.A(KEYINPUT36), .ZN(new_n755));
  NAND4_X1  g330(.A1(new_n735), .A2(new_n750), .A3(new_n755), .A4(new_n752), .ZN(new_n756));
  NAND2_X1  g331(.A1(new_n754), .A2(new_n756), .ZN(new_n757));
  NAND2_X1  g332(.A1(new_n717), .A2(G21), .ZN(new_n758));
  OAI21_X1  g333(.A(new_n758), .B1(G168), .B2(new_n717), .ZN(new_n759));
  NOR2_X1   g334(.A1(new_n759), .A2(G1966), .ZN(new_n760));
  INV_X1    g335(.A(G29), .ZN(new_n761));
  NAND2_X1  g336(.A1(new_n761), .A2(G35), .ZN(new_n762));
  OAI21_X1  g337(.A(new_n762), .B1(G162), .B2(new_n761), .ZN(new_n763));
  XOR2_X1   g338(.A(new_n763), .B(KEYINPUT29), .Z(new_n764));
  INV_X1    g339(.A(G2090), .ZN(new_n765));
  AOI21_X1  g340(.A(new_n760), .B1(new_n764), .B2(new_n765), .ZN(new_n766));
  OAI21_X1  g341(.A(new_n766), .B1(new_n765), .B2(new_n764), .ZN(new_n767));
  XNOR2_X1  g342(.A(KEYINPUT30), .B(G28), .ZN(new_n768));
  OR2_X1    g343(.A1(KEYINPUT31), .A2(G11), .ZN(new_n769));
  NAND2_X1  g344(.A1(KEYINPUT31), .A2(G11), .ZN(new_n770));
  AOI22_X1  g345(.A1(new_n768), .A2(new_n761), .B1(new_n769), .B2(new_n770), .ZN(new_n771));
  OAI21_X1  g346(.A(new_n771), .B1(new_n636), .B2(new_n761), .ZN(new_n772));
  NAND2_X1  g347(.A1(new_n761), .A2(G26), .ZN(new_n773));
  XNOR2_X1  g348(.A(new_n773), .B(KEYINPUT28), .ZN(new_n774));
  NAND2_X1  g349(.A1(new_n484), .A2(G140), .ZN(new_n775));
  NAND2_X1  g350(.A1(new_n486), .A2(G128), .ZN(new_n776));
  OR2_X1    g351(.A1(G104), .A2(G2105), .ZN(new_n777));
  OAI211_X1 g352(.A(new_n777), .B(G2104), .C1(G116), .C2(new_n463), .ZN(new_n778));
  NAND3_X1  g353(.A1(new_n775), .A2(new_n776), .A3(new_n778), .ZN(new_n779));
  INV_X1    g354(.A(new_n779), .ZN(new_n780));
  OAI21_X1  g355(.A(new_n774), .B1(new_n780), .B2(new_n761), .ZN(new_n781));
  XNOR2_X1  g356(.A(new_n781), .B(G2067), .ZN(new_n782));
  AOI211_X1 g357(.A(new_n772), .B(new_n782), .C1(G1966), .C2(new_n759), .ZN(new_n783));
  NAND2_X1  g358(.A1(new_n717), .A2(G5), .ZN(new_n784));
  OAI21_X1  g359(.A(new_n784), .B1(G171), .B2(new_n717), .ZN(new_n785));
  INV_X1    g360(.A(G1961), .ZN(new_n786));
  XNOR2_X1  g361(.A(new_n785), .B(new_n786), .ZN(new_n787));
  NAND2_X1  g362(.A1(G164), .A2(G29), .ZN(new_n788));
  OAI21_X1  g363(.A(new_n788), .B1(G27), .B2(G29), .ZN(new_n789));
  INV_X1    g364(.A(G2078), .ZN(new_n790));
  OR2_X1    g365(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  NAND2_X1  g366(.A1(new_n761), .A2(G32), .ZN(new_n792));
  INV_X1    g367(.A(G141), .ZN(new_n793));
  AOI21_X1  g368(.A(KEYINPUT101), .B1(new_n476), .B2(G105), .ZN(new_n794));
  NAND2_X1  g369(.A1(new_n476), .A2(G105), .ZN(new_n795));
  INV_X1    g370(.A(KEYINPUT101), .ZN(new_n796));
  NOR2_X1   g371(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  OAI22_X1  g372(.A1(new_n479), .A2(new_n793), .B1(new_n794), .B2(new_n797), .ZN(new_n798));
  NAND2_X1  g373(.A1(new_n486), .A2(G129), .ZN(new_n799));
  NAND3_X1  g374(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n800));
  XOR2_X1   g375(.A(new_n800), .B(KEYINPUT26), .Z(new_n801));
  NAND2_X1  g376(.A1(new_n799), .A2(new_n801), .ZN(new_n802));
  NOR2_X1   g377(.A1(new_n798), .A2(new_n802), .ZN(new_n803));
  OAI21_X1  g378(.A(new_n792), .B1(new_n803), .B2(new_n761), .ZN(new_n804));
  XOR2_X1   g379(.A(KEYINPUT27), .B(G1996), .Z(new_n805));
  XNOR2_X1  g380(.A(new_n804), .B(new_n805), .ZN(new_n806));
  AOI21_X1  g381(.A(new_n806), .B1(new_n790), .B2(new_n789), .ZN(new_n807));
  NAND4_X1  g382(.A1(new_n783), .A2(new_n787), .A3(new_n791), .A4(new_n807), .ZN(new_n808));
  AND2_X1   g383(.A1(KEYINPUT24), .A2(G34), .ZN(new_n809));
  NOR2_X1   g384(.A1(KEYINPUT24), .A2(G34), .ZN(new_n810));
  OAI21_X1  g385(.A(new_n761), .B1(new_n809), .B2(new_n810), .ZN(new_n811));
  XNOR2_X1  g386(.A(new_n811), .B(KEYINPUT100), .ZN(new_n812));
  AOI21_X1  g387(.A(new_n812), .B1(G160), .B2(G29), .ZN(new_n813));
  AOI211_X1 g388(.A(new_n767), .B(new_n808), .C1(G2084), .C2(new_n813), .ZN(new_n814));
  AND2_X1   g389(.A1(new_n761), .A2(G33), .ZN(new_n815));
  NAND3_X1  g390(.A1(new_n467), .A2(new_n470), .A3(G127), .ZN(new_n816));
  NAND2_X1  g391(.A1(G115), .A2(G2104), .ZN(new_n817));
  NAND2_X1  g392(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  NAND2_X1  g393(.A1(new_n818), .A2(G2105), .ZN(new_n819));
  INV_X1    g394(.A(KEYINPUT99), .ZN(new_n820));
  NAND3_X1  g395(.A1(new_n463), .A2(G103), .A3(G2104), .ZN(new_n821));
  INV_X1    g396(.A(KEYINPUT25), .ZN(new_n822));
  XNOR2_X1  g397(.A(new_n821), .B(new_n822), .ZN(new_n823));
  NAND3_X1  g398(.A1(new_n478), .A2(G139), .A3(new_n463), .ZN(new_n824));
  NAND2_X1  g399(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  INV_X1    g400(.A(new_n825), .ZN(new_n826));
  NAND3_X1  g401(.A1(new_n819), .A2(new_n820), .A3(new_n826), .ZN(new_n827));
  AOI21_X1  g402(.A(new_n463), .B1(new_n816), .B2(new_n817), .ZN(new_n828));
  OAI21_X1  g403(.A(KEYINPUT99), .B1(new_n828), .B2(new_n825), .ZN(new_n829));
  NAND2_X1  g404(.A1(new_n827), .A2(new_n829), .ZN(new_n830));
  AOI21_X1  g405(.A(new_n815), .B1(new_n830), .B2(G29), .ZN(new_n831));
  INV_X1    g406(.A(G2072), .ZN(new_n832));
  OR2_X1    g407(.A1(new_n831), .A2(new_n832), .ZN(new_n833));
  OR2_X1    g408(.A1(new_n813), .A2(G2084), .ZN(new_n834));
  NAND2_X1  g409(.A1(new_n831), .A2(new_n832), .ZN(new_n835));
  NAND4_X1  g410(.A1(new_n814), .A2(new_n833), .A3(new_n834), .A4(new_n835), .ZN(new_n836));
  NOR2_X1   g411(.A1(G16), .A2(G19), .ZN(new_n837));
  AOI21_X1  g412(.A(new_n837), .B1(new_n557), .B2(G16), .ZN(new_n838));
  XNOR2_X1  g413(.A(new_n838), .B(KEYINPUT98), .ZN(new_n839));
  XOR2_X1   g414(.A(new_n839), .B(G1341), .Z(new_n840));
  NOR2_X1   g415(.A1(G4), .A2(G16), .ZN(new_n841));
  AOI21_X1  g416(.A(new_n841), .B1(new_n609), .B2(G16), .ZN(new_n842));
  OR2_X1    g417(.A1(new_n842), .A2(G1348), .ZN(new_n843));
  NAND2_X1  g418(.A1(new_n717), .A2(G20), .ZN(new_n844));
  XNOR2_X1  g419(.A(new_n844), .B(KEYINPUT23), .ZN(new_n845));
  INV_X1    g420(.A(G299), .ZN(new_n846));
  OAI21_X1  g421(.A(new_n845), .B1(new_n846), .B2(new_n717), .ZN(new_n847));
  INV_X1    g422(.A(G1956), .ZN(new_n848));
  XNOR2_X1  g423(.A(new_n847), .B(new_n848), .ZN(new_n849));
  NAND2_X1  g424(.A1(new_n842), .A2(G1348), .ZN(new_n850));
  NAND4_X1  g425(.A1(new_n840), .A2(new_n843), .A3(new_n849), .A4(new_n850), .ZN(new_n851));
  NOR2_X1   g426(.A1(new_n836), .A2(new_n851), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n757), .A2(new_n852), .ZN(G150));
  INV_X1    g428(.A(G150), .ZN(G311));
  NAND2_X1  g429(.A1(new_n609), .A2(G559), .ZN(new_n855));
  XNOR2_X1  g430(.A(KEYINPUT102), .B(KEYINPUT38), .ZN(new_n856));
  XNOR2_X1  g431(.A(new_n856), .B(KEYINPUT103), .ZN(new_n857));
  XNOR2_X1  g432(.A(new_n855), .B(new_n857), .ZN(new_n858));
  AND2_X1   g433(.A1(new_n554), .A2(new_n555), .ZN(new_n859));
  AOI22_X1  g434(.A1(G55), .A2(new_n526), .B1(new_n523), .B2(G93), .ZN(new_n860));
  AOI22_X1  g435(.A1(new_n531), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n861));
  OR2_X1    g436(.A1(new_n861), .A2(new_n508), .ZN(new_n862));
  NAND4_X1  g437(.A1(new_n859), .A2(new_n860), .A3(new_n553), .A4(new_n862), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n860), .A2(new_n862), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n864), .A2(new_n556), .ZN(new_n865));
  NAND2_X1  g440(.A1(new_n863), .A2(new_n865), .ZN(new_n866));
  XNOR2_X1  g441(.A(new_n858), .B(new_n866), .ZN(new_n867));
  NOR2_X1   g442(.A1(new_n867), .A2(KEYINPUT39), .ZN(new_n868));
  XOR2_X1   g443(.A(new_n868), .B(KEYINPUT104), .Z(new_n869));
  XNOR2_X1  g444(.A(KEYINPUT105), .B(G860), .ZN(new_n870));
  AOI21_X1  g445(.A(new_n870), .B1(new_n867), .B2(KEYINPUT39), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n869), .A2(new_n871), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n864), .A2(new_n870), .ZN(new_n873));
  XOR2_X1   g448(.A(new_n873), .B(KEYINPUT37), .Z(new_n874));
  NAND2_X1  g449(.A1(new_n872), .A2(new_n874), .ZN(G145));
  XNOR2_X1  g450(.A(G160), .B(G162), .ZN(new_n876));
  XNOR2_X1  g451(.A(new_n876), .B(new_n636), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n484), .A2(G142), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n486), .A2(G130), .ZN(new_n879));
  OR2_X1    g454(.A1(G106), .A2(G2105), .ZN(new_n880));
  OAI211_X1 g455(.A(new_n880), .B(G2104), .C1(G118), .C2(new_n463), .ZN(new_n881));
  NAND3_X1  g456(.A1(new_n878), .A2(new_n879), .A3(new_n881), .ZN(new_n882));
  AND3_X1   g457(.A1(new_n623), .A2(new_n624), .A3(new_n882), .ZN(new_n883));
  AOI21_X1  g458(.A(new_n882), .B1(new_n623), .B2(new_n624), .ZN(new_n884));
  OR3_X1    g459(.A1(new_n883), .A2(new_n884), .A3(new_n729), .ZN(new_n885));
  OAI21_X1  g460(.A(new_n729), .B1(new_n883), .B2(new_n884), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  INV_X1    g462(.A(KEYINPUT106), .ZN(new_n888));
  NAND3_X1  g463(.A1(new_n496), .A2(new_n502), .A3(new_n888), .ZN(new_n889));
  INV_X1    g464(.A(new_n889), .ZN(new_n890));
  AOI21_X1  g465(.A(new_n888), .B1(new_n496), .B2(new_n502), .ZN(new_n891));
  NOR2_X1   g466(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  INV_X1    g467(.A(new_n892), .ZN(new_n893));
  INV_X1    g468(.A(new_n803), .ZN(new_n894));
  AND3_X1   g469(.A1(new_n830), .A2(KEYINPUT107), .A3(new_n894), .ZN(new_n895));
  AOI21_X1  g470(.A(new_n894), .B1(new_n830), .B2(KEYINPUT107), .ZN(new_n896));
  NOR3_X1   g471(.A1(new_n895), .A2(new_n896), .A3(new_n780), .ZN(new_n897));
  AOI21_X1  g472(.A(new_n820), .B1(new_n819), .B2(new_n826), .ZN(new_n898));
  NOR3_X1   g473(.A1(new_n828), .A2(new_n825), .A3(KEYINPUT99), .ZN(new_n899));
  OAI21_X1  g474(.A(KEYINPUT107), .B1(new_n898), .B2(new_n899), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n900), .A2(new_n803), .ZN(new_n901));
  NAND3_X1  g476(.A1(new_n830), .A2(KEYINPUT107), .A3(new_n894), .ZN(new_n902));
  AOI21_X1  g477(.A(new_n779), .B1(new_n901), .B2(new_n902), .ZN(new_n903));
  OAI21_X1  g478(.A(new_n893), .B1(new_n897), .B2(new_n903), .ZN(new_n904));
  OAI21_X1  g479(.A(new_n780), .B1(new_n895), .B2(new_n896), .ZN(new_n905));
  NAND3_X1  g480(.A1(new_n901), .A2(new_n779), .A3(new_n902), .ZN(new_n906));
  NAND3_X1  g481(.A1(new_n905), .A2(new_n906), .A3(new_n892), .ZN(new_n907));
  AOI21_X1  g482(.A(new_n887), .B1(new_n904), .B2(new_n907), .ZN(new_n908));
  INV_X1    g483(.A(KEYINPUT108), .ZN(new_n909));
  NAND3_X1  g484(.A1(new_n904), .A2(new_n887), .A3(new_n907), .ZN(new_n910));
  AOI21_X1  g485(.A(new_n908), .B1(new_n909), .B2(new_n910), .ZN(new_n911));
  AOI211_X1 g486(.A(KEYINPUT108), .B(new_n887), .C1(new_n904), .C2(new_n907), .ZN(new_n912));
  OAI21_X1  g487(.A(new_n877), .B1(new_n911), .B2(new_n912), .ZN(new_n913));
  NOR2_X1   g488(.A1(new_n908), .A2(new_n877), .ZN(new_n914));
  AOI21_X1  g489(.A(G37), .B1(new_n914), .B2(new_n910), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n913), .A2(new_n915), .ZN(new_n916));
  XNOR2_X1  g491(.A(new_n916), .B(KEYINPUT40), .ZN(G395));
  INV_X1    g492(.A(KEYINPUT110), .ZN(new_n918));
  INV_X1    g493(.A(KEYINPUT109), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n607), .A2(new_n608), .ZN(new_n920));
  INV_X1    g495(.A(new_n604), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  AOI21_X1  g497(.A(new_n919), .B1(new_n922), .B2(new_n846), .ZN(new_n923));
  NOR3_X1   g498(.A1(new_n609), .A2(KEYINPUT109), .A3(G299), .ZN(new_n924));
  OAI21_X1  g499(.A(new_n918), .B1(new_n923), .B2(new_n924), .ZN(new_n925));
  INV_X1    g500(.A(KEYINPUT41), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n609), .A2(G299), .ZN(new_n927));
  NAND3_X1  g502(.A1(new_n922), .A2(new_n919), .A3(new_n846), .ZN(new_n928));
  OAI21_X1  g503(.A(KEYINPUT109), .B1(new_n609), .B2(G299), .ZN(new_n929));
  NAND3_X1  g504(.A1(new_n928), .A2(new_n929), .A3(KEYINPUT110), .ZN(new_n930));
  NAND4_X1  g505(.A1(new_n925), .A2(new_n926), .A3(new_n927), .A4(new_n930), .ZN(new_n931));
  NAND3_X1  g506(.A1(new_n928), .A2(new_n929), .A3(new_n927), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n932), .A2(KEYINPUT41), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n931), .A2(new_n933), .ZN(new_n934));
  XOR2_X1   g509(.A(new_n618), .B(new_n866), .Z(new_n935));
  OR2_X1    g510(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n935), .A2(new_n932), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n938), .A2(KEYINPUT42), .ZN(new_n939));
  XOR2_X1   g514(.A(G166), .B(G288), .Z(new_n940));
  INV_X1    g515(.A(new_n940), .ZN(new_n941));
  NAND2_X1  g516(.A1(G290), .A2(G305), .ZN(new_n942));
  OAI21_X1  g517(.A(new_n599), .B1(new_n589), .B2(new_n590), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n941), .A2(new_n944), .ZN(new_n945));
  NAND3_X1  g520(.A1(new_n940), .A2(new_n942), .A3(new_n943), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n945), .A2(new_n946), .ZN(new_n947));
  INV_X1    g522(.A(new_n947), .ZN(new_n948));
  INV_X1    g523(.A(KEYINPUT42), .ZN(new_n949));
  NAND3_X1  g524(.A1(new_n936), .A2(new_n949), .A3(new_n937), .ZN(new_n950));
  AND3_X1   g525(.A1(new_n939), .A2(new_n948), .A3(new_n950), .ZN(new_n951));
  AOI21_X1  g526(.A(new_n948), .B1(new_n939), .B2(new_n950), .ZN(new_n952));
  OAI21_X1  g527(.A(G868), .B1(new_n951), .B2(new_n952), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n864), .A2(new_n616), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n953), .A2(new_n954), .ZN(G295));
  NAND2_X1  g530(.A1(new_n953), .A2(new_n954), .ZN(G331));
  NAND2_X1  g531(.A1(G301), .A2(new_n544), .ZN(new_n957));
  OAI211_X1 g532(.A(new_n866), .B(new_n957), .C1(G286), .C2(G301), .ZN(new_n958));
  AOI21_X1  g533(.A(G301), .B1(new_n573), .B2(new_n575), .ZN(new_n959));
  INV_X1    g534(.A(new_n957), .ZN(new_n960));
  OAI211_X1 g535(.A(new_n865), .B(new_n863), .C1(new_n959), .C2(new_n960), .ZN(new_n961));
  AND2_X1   g536(.A1(new_n958), .A2(new_n961), .ZN(new_n962));
  NOR2_X1   g537(.A1(new_n962), .A2(new_n932), .ZN(new_n963));
  AOI21_X1  g538(.A(new_n963), .B1(new_n934), .B2(new_n962), .ZN(new_n964));
  AOI21_X1  g539(.A(G37), .B1(new_n964), .B2(new_n947), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n958), .A2(new_n961), .ZN(new_n966));
  AOI21_X1  g541(.A(new_n966), .B1(new_n931), .B2(new_n933), .ZN(new_n967));
  OAI21_X1  g542(.A(new_n948), .B1(new_n967), .B2(new_n963), .ZN(new_n968));
  AOI21_X1  g543(.A(KEYINPUT43), .B1(new_n965), .B2(new_n968), .ZN(new_n969));
  NAND3_X1  g544(.A1(new_n958), .A2(new_n961), .A3(KEYINPUT41), .ZN(new_n970));
  INV_X1    g545(.A(new_n932), .ZN(new_n971));
  AOI22_X1  g546(.A1(new_n945), .A2(new_n946), .B1(new_n970), .B2(new_n971), .ZN(new_n972));
  NAND3_X1  g547(.A1(new_n925), .A2(new_n927), .A3(new_n930), .ZN(new_n973));
  NAND3_X1  g548(.A1(new_n973), .A2(KEYINPUT41), .A3(new_n962), .ZN(new_n974));
  AOI21_X1  g549(.A(G37), .B1(new_n972), .B2(new_n974), .ZN(new_n975));
  AND3_X1   g550(.A1(new_n968), .A2(new_n975), .A3(KEYINPUT43), .ZN(new_n976));
  OAI21_X1  g551(.A(KEYINPUT44), .B1(new_n969), .B2(new_n976), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n934), .A2(new_n962), .ZN(new_n978));
  INV_X1    g553(.A(new_n963), .ZN(new_n979));
  NAND3_X1  g554(.A1(new_n978), .A2(new_n947), .A3(new_n979), .ZN(new_n980));
  INV_X1    g555(.A(G37), .ZN(new_n981));
  NAND3_X1  g556(.A1(new_n980), .A2(new_n968), .A3(new_n981), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n982), .A2(KEYINPUT43), .ZN(new_n983));
  INV_X1    g558(.A(KEYINPUT43), .ZN(new_n984));
  NAND3_X1  g559(.A1(new_n968), .A2(new_n975), .A3(new_n984), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n983), .A2(new_n985), .ZN(new_n986));
  INV_X1    g561(.A(new_n986), .ZN(new_n987));
  OAI21_X1  g562(.A(new_n977), .B1(new_n987), .B2(KEYINPUT44), .ZN(G397));
  INV_X1    g563(.A(KEYINPUT45), .ZN(new_n989));
  XNOR2_X1  g564(.A(KEYINPUT111), .B(G1384), .ZN(new_n990));
  INV_X1    g565(.A(new_n990), .ZN(new_n991));
  OAI21_X1  g566(.A(new_n989), .B1(new_n893), .B2(new_n991), .ZN(new_n992));
  NAND2_X1  g567(.A1(new_n482), .A2(G40), .ZN(new_n993));
  NOR2_X1   g568(.A1(new_n992), .A2(new_n993), .ZN(new_n994));
  INV_X1    g569(.A(G2067), .ZN(new_n995));
  XNOR2_X1  g570(.A(new_n779), .B(new_n995), .ZN(new_n996));
  INV_X1    g571(.A(new_n996), .ZN(new_n997));
  OAI21_X1  g572(.A(new_n994), .B1(new_n894), .B2(new_n997), .ZN(new_n998));
  INV_X1    g573(.A(G1996), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n994), .A2(new_n999), .ZN(new_n1000));
  AND2_X1   g575(.A1(new_n1000), .A2(KEYINPUT46), .ZN(new_n1001));
  NOR2_X1   g576(.A1(new_n1000), .A2(KEYINPUT46), .ZN(new_n1002));
  OAI21_X1  g577(.A(new_n998), .B1(new_n1001), .B2(new_n1002), .ZN(new_n1003));
  XOR2_X1   g578(.A(new_n1003), .B(KEYINPUT47), .Z(new_n1004));
  XNOR2_X1  g579(.A(new_n803), .B(G1996), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n1005), .A2(new_n996), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n730), .A2(new_n733), .ZN(new_n1007));
  OAI22_X1  g582(.A1(new_n1006), .A2(new_n1007), .B1(G2067), .B2(new_n779), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n1008), .A2(new_n994), .ZN(new_n1009));
  NOR2_X1   g584(.A1(G290), .A2(G1986), .ZN(new_n1010));
  NAND3_X1  g585(.A1(new_n994), .A2(new_n1010), .A3(KEYINPUT48), .ZN(new_n1011));
  OR2_X1    g586(.A1(new_n730), .A2(new_n733), .ZN(new_n1012));
  NAND4_X1  g587(.A1(new_n1005), .A2(new_n996), .A3(new_n1007), .A4(new_n1012), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n994), .A2(new_n1013), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n1011), .A2(new_n1014), .ZN(new_n1015));
  AOI21_X1  g590(.A(KEYINPUT48), .B1(new_n994), .B2(new_n1010), .ZN(new_n1016));
  OAI21_X1  g591(.A(new_n1009), .B1(new_n1015), .B2(new_n1016), .ZN(new_n1017));
  NOR2_X1   g592(.A1(new_n1004), .A2(new_n1017), .ZN(new_n1018));
  INV_X1    g593(.A(G8), .ZN(new_n1019));
  NOR2_X1   g594(.A1(G166), .A2(new_n1019), .ZN(new_n1020));
  XNOR2_X1  g595(.A(KEYINPUT115), .B(KEYINPUT55), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n1020), .A2(new_n1021), .ZN(new_n1022));
  NAND2_X1  g597(.A1(KEYINPUT115), .A2(KEYINPUT55), .ZN(new_n1023));
  OAI21_X1  g598(.A(new_n1023), .B1(G166), .B2(new_n1019), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n1022), .A2(new_n1024), .ZN(new_n1025));
  INV_X1    g600(.A(new_n1025), .ZN(new_n1026));
  AOI211_X1 g601(.A(KEYINPUT50), .B(G1384), .C1(new_n496), .C2(new_n502), .ZN(new_n1027));
  NOR2_X1   g602(.A1(new_n1027), .A2(new_n993), .ZN(new_n1028));
  AOI21_X1  g603(.A(G1384), .B1(new_n496), .B2(new_n502), .ZN(new_n1029));
  INV_X1    g604(.A(new_n1029), .ZN(new_n1030));
  NAND2_X1  g605(.A1(new_n1030), .A2(KEYINPUT50), .ZN(new_n1031));
  AND3_X1   g606(.A1(new_n1028), .A2(new_n765), .A3(new_n1031), .ZN(new_n1032));
  INV_X1    g607(.A(G40), .ZN(new_n1033));
  NOR3_X1   g608(.A1(new_n474), .A2(new_n481), .A3(new_n1033), .ZN(new_n1034));
  OAI21_X1  g609(.A(new_n1034), .B1(new_n1029), .B2(KEYINPUT45), .ZN(new_n1035));
  INV_X1    g610(.A(new_n1035), .ZN(new_n1036));
  INV_X1    g611(.A(KEYINPUT112), .ZN(new_n1037));
  NOR2_X1   g612(.A1(new_n991), .A2(new_n989), .ZN(new_n1038));
  AOI21_X1  g613(.A(new_n1037), .B1(new_n892), .B2(new_n1038), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n503), .A2(KEYINPUT106), .ZN(new_n1040));
  NAND3_X1  g615(.A1(new_n1040), .A2(new_n889), .A3(new_n1038), .ZN(new_n1041));
  NOR2_X1   g616(.A1(new_n1041), .A2(KEYINPUT112), .ZN(new_n1042));
  OAI21_X1  g617(.A(new_n1036), .B1(new_n1039), .B2(new_n1042), .ZN(new_n1043));
  INV_X1    g618(.A(G1971), .ZN(new_n1044));
  AOI21_X1  g619(.A(new_n1032), .B1(new_n1043), .B2(new_n1044), .ZN(new_n1045));
  OAI21_X1  g620(.A(new_n1026), .B1(new_n1045), .B2(new_n1019), .ZN(new_n1046));
  AOI21_X1  g621(.A(new_n1019), .B1(new_n1034), .B2(new_n1029), .ZN(new_n1047));
  INV_X1    g622(.A(G1976), .ZN(new_n1048));
  OAI21_X1  g623(.A(new_n1047), .B1(G288), .B2(new_n1048), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n1049), .A2(KEYINPUT52), .ZN(new_n1050));
  INV_X1    g625(.A(KEYINPUT52), .ZN(new_n1051));
  OAI21_X1  g626(.A(new_n1051), .B1(new_n740), .B2(G1976), .ZN(new_n1052));
  OAI21_X1  g627(.A(new_n1050), .B1(new_n1052), .B2(new_n1049), .ZN(new_n1053));
  INV_X1    g628(.A(KEYINPUT118), .ZN(new_n1054));
  INV_X1    g629(.A(G1981), .ZN(new_n1055));
  NAND3_X1  g630(.A1(new_n586), .A2(new_n1055), .A3(new_n588), .ZN(new_n1056));
  NAND4_X1  g631(.A1(new_n510), .A2(new_n514), .A3(G48), .A4(G543), .ZN(new_n1057));
  NAND4_X1  g632(.A1(new_n531), .A2(G86), .A3(new_n510), .A4(new_n514), .ZN(new_n1058));
  AOI22_X1  g633(.A1(new_n531), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n1059));
  OAI211_X1 g634(.A(new_n1057), .B(new_n1058), .C1(new_n1059), .C2(new_n508), .ZN(new_n1060));
  INV_X1    g635(.A(KEYINPUT117), .ZN(new_n1061));
  NAND3_X1  g636(.A1(new_n1060), .A2(new_n1061), .A3(G1981), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n1056), .A2(new_n1062), .ZN(new_n1063));
  AOI21_X1  g638(.A(new_n1061), .B1(new_n1060), .B2(G1981), .ZN(new_n1064));
  NOR2_X1   g639(.A1(new_n1063), .A2(new_n1064), .ZN(new_n1065));
  OAI21_X1  g640(.A(new_n1054), .B1(new_n1065), .B2(KEYINPUT49), .ZN(new_n1066));
  INV_X1    g641(.A(KEYINPUT49), .ZN(new_n1067));
  OAI211_X1 g642(.A(KEYINPUT118), .B(new_n1067), .C1(new_n1063), .C2(new_n1064), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n1066), .A2(new_n1068), .ZN(new_n1069));
  INV_X1    g644(.A(new_n1047), .ZN(new_n1070));
  AOI21_X1  g645(.A(new_n1070), .B1(new_n1065), .B2(KEYINPUT49), .ZN(new_n1071));
  AOI21_X1  g646(.A(new_n1053), .B1(new_n1069), .B2(new_n1071), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n1046), .A2(new_n1072), .ZN(new_n1073));
  NAND3_X1  g648(.A1(new_n1030), .A2(KEYINPUT113), .A3(KEYINPUT50), .ZN(new_n1074));
  INV_X1    g649(.A(KEYINPUT113), .ZN(new_n1075));
  INV_X1    g650(.A(KEYINPUT50), .ZN(new_n1076));
  OAI21_X1  g651(.A(new_n1075), .B1(new_n1029), .B2(new_n1076), .ZN(new_n1077));
  NAND3_X1  g652(.A1(new_n1028), .A2(new_n1074), .A3(new_n1077), .ZN(new_n1078));
  OAI21_X1  g653(.A(KEYINPUT114), .B1(new_n1078), .B2(G2090), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n1029), .A2(new_n1076), .ZN(new_n1080));
  AND3_X1   g655(.A1(new_n1077), .A2(new_n1034), .A3(new_n1080), .ZN(new_n1081));
  INV_X1    g656(.A(KEYINPUT114), .ZN(new_n1082));
  NAND4_X1  g657(.A1(new_n1081), .A2(new_n1082), .A3(new_n765), .A4(new_n1074), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n1079), .A2(new_n1083), .ZN(new_n1084));
  NAND3_X1  g659(.A1(new_n892), .A2(new_n1037), .A3(new_n1038), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n1041), .A2(KEYINPUT112), .ZN(new_n1086));
  AOI21_X1  g661(.A(new_n1035), .B1(new_n1085), .B2(new_n1086), .ZN(new_n1087));
  NOR2_X1   g662(.A1(new_n1087), .A2(G1971), .ZN(new_n1088));
  OAI211_X1 g663(.A(G8), .B(new_n1025), .C1(new_n1084), .C2(new_n1088), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n1089), .A2(KEYINPUT116), .ZN(new_n1090));
  OAI211_X1 g665(.A(new_n1079), .B(new_n1083), .C1(G1971), .C2(new_n1087), .ZN(new_n1091));
  INV_X1    g666(.A(KEYINPUT116), .ZN(new_n1092));
  NAND4_X1  g667(.A1(new_n1091), .A2(new_n1092), .A3(G8), .A4(new_n1025), .ZN(new_n1093));
  AOI21_X1  g668(.A(new_n1073), .B1(new_n1090), .B2(new_n1093), .ZN(new_n1094));
  INV_X1    g669(.A(G2084), .ZN(new_n1095));
  NAND4_X1  g670(.A1(new_n1028), .A2(new_n1074), .A3(new_n1095), .A4(new_n1077), .ZN(new_n1096));
  INV_X1    g671(.A(G1966), .ZN(new_n1097));
  NOR2_X1   g672(.A1(new_n1030), .A2(new_n989), .ZN(new_n1098));
  OAI21_X1  g673(.A(new_n1097), .B1(new_n1098), .B2(new_n1035), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n1096), .A2(new_n1099), .ZN(new_n1100));
  INV_X1    g675(.A(KEYINPUT124), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n1100), .A2(new_n1101), .ZN(new_n1102));
  NAND3_X1  g677(.A1(new_n1096), .A2(KEYINPUT124), .A3(new_n1099), .ZN(new_n1103));
  NAND3_X1  g678(.A1(new_n1102), .A2(G168), .A3(new_n1103), .ZN(new_n1104));
  INV_X1    g679(.A(KEYINPUT51), .ZN(new_n1105));
  NOR2_X1   g680(.A1(new_n1105), .A2(new_n1019), .ZN(new_n1106));
  NAND2_X1  g681(.A1(new_n1104), .A2(new_n1106), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n1100), .A2(G8), .ZN(new_n1108));
  AOI21_X1  g683(.A(KEYINPUT51), .B1(new_n544), .B2(G8), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n1108), .A2(new_n1109), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n1107), .A2(new_n1110), .ZN(new_n1111));
  INV_X1    g686(.A(KEYINPUT62), .ZN(new_n1112));
  INV_X1    g687(.A(new_n1103), .ZN(new_n1113));
  AOI21_X1  g688(.A(KEYINPUT124), .B1(new_n1096), .B2(new_n1099), .ZN(new_n1114));
  NOR2_X1   g689(.A1(new_n1113), .A2(new_n1114), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n544), .A2(G8), .ZN(new_n1116));
  OR2_X1    g691(.A1(new_n1115), .A2(new_n1116), .ZN(new_n1117));
  NAND3_X1  g692(.A1(new_n1111), .A2(new_n1112), .A3(new_n1117), .ZN(new_n1118));
  AOI22_X1  g693(.A1(new_n1104), .A2(new_n1106), .B1(new_n1108), .B2(new_n1109), .ZN(new_n1119));
  NOR2_X1   g694(.A1(new_n1115), .A2(new_n1116), .ZN(new_n1120));
  OAI21_X1  g695(.A(KEYINPUT62), .B1(new_n1119), .B2(new_n1120), .ZN(new_n1121));
  INV_X1    g696(.A(KEYINPUT53), .ZN(new_n1122));
  OAI21_X1  g697(.A(new_n1122), .B1(new_n1043), .B2(G2078), .ZN(new_n1123));
  NOR2_X1   g698(.A1(new_n1098), .A2(new_n1035), .ZN(new_n1124));
  NOR2_X1   g699(.A1(new_n1122), .A2(G2078), .ZN(new_n1125));
  AOI22_X1  g700(.A1(new_n1078), .A2(new_n786), .B1(new_n1124), .B2(new_n1125), .ZN(new_n1126));
  AOI21_X1  g701(.A(G301), .B1(new_n1123), .B2(new_n1126), .ZN(new_n1127));
  NAND4_X1  g702(.A1(new_n1094), .A2(new_n1118), .A3(new_n1121), .A4(new_n1127), .ZN(new_n1128));
  AND2_X1   g703(.A1(new_n1090), .A2(new_n1093), .ZN(new_n1129));
  INV_X1    g704(.A(KEYINPUT63), .ZN(new_n1130));
  NOR2_X1   g705(.A1(new_n1108), .A2(G286), .ZN(new_n1131));
  AND3_X1   g706(.A1(new_n1046), .A2(new_n1130), .A3(new_n1131), .ZN(new_n1132));
  OAI21_X1  g707(.A(new_n1072), .B1(new_n1129), .B2(new_n1132), .ZN(new_n1133));
  NAND2_X1  g708(.A1(new_n1069), .A2(new_n1071), .ZN(new_n1134));
  NAND3_X1  g709(.A1(new_n1134), .A2(new_n1048), .A3(new_n740), .ZN(new_n1135));
  AOI21_X1  g710(.A(new_n1070), .B1(new_n1135), .B2(new_n1056), .ZN(new_n1136));
  AND2_X1   g711(.A1(new_n1091), .A2(G8), .ZN(new_n1137));
  OAI211_X1 g712(.A(new_n1072), .B(new_n1131), .C1(new_n1137), .C2(new_n1025), .ZN(new_n1138));
  AOI21_X1  g713(.A(new_n1136), .B1(new_n1138), .B2(KEYINPUT63), .ZN(new_n1139));
  NAND3_X1  g714(.A1(new_n1128), .A2(new_n1133), .A3(new_n1139), .ZN(new_n1140));
  XOR2_X1   g715(.A(new_n481), .B(KEYINPUT125), .Z(new_n1141));
  OR3_X1    g716(.A1(new_n1141), .A2(new_n1033), .A3(new_n474), .ZN(new_n1142));
  AOI211_X1 g717(.A(new_n1122), .B(G2078), .C1(new_n1142), .C2(KEYINPUT126), .ZN(new_n1143));
  NAND2_X1  g718(.A1(new_n1085), .A2(new_n1086), .ZN(new_n1144));
  OR2_X1    g719(.A1(new_n1142), .A2(KEYINPUT126), .ZN(new_n1145));
  NAND4_X1  g720(.A1(new_n1143), .A2(new_n1144), .A3(new_n992), .A4(new_n1145), .ZN(new_n1146));
  XNOR2_X1  g721(.A(G301), .B(KEYINPUT54), .ZN(new_n1147));
  AOI21_X1  g722(.A(new_n1147), .B1(new_n1078), .B2(new_n786), .ZN(new_n1148));
  AND2_X1   g723(.A1(new_n1146), .A2(new_n1148), .ZN(new_n1149));
  NAND2_X1  g724(.A1(new_n1123), .A2(new_n1126), .ZN(new_n1150));
  AOI22_X1  g725(.A1(new_n1149), .A2(new_n1123), .B1(new_n1150), .B2(new_n1147), .ZN(new_n1151));
  NAND2_X1  g726(.A1(new_n1111), .A2(new_n1117), .ZN(new_n1152));
  NAND3_X1  g727(.A1(new_n1094), .A2(new_n1151), .A3(new_n1152), .ZN(new_n1153));
  XNOR2_X1  g728(.A(KEYINPUT56), .B(G2072), .ZN(new_n1154));
  NAND3_X1  g729(.A1(new_n1144), .A2(new_n1036), .A3(new_n1154), .ZN(new_n1155));
  AOI21_X1  g730(.A(G1956), .B1(new_n1028), .B2(new_n1031), .ZN(new_n1156));
  INV_X1    g731(.A(new_n1156), .ZN(new_n1157));
  NAND2_X1  g732(.A1(new_n1155), .A2(new_n1157), .ZN(new_n1158));
  INV_X1    g733(.A(KEYINPUT121), .ZN(new_n1159));
  XOR2_X1   g734(.A(G299), .B(KEYINPUT57), .Z(new_n1160));
  INV_X1    g735(.A(new_n1160), .ZN(new_n1161));
  NAND3_X1  g736(.A1(new_n1158), .A2(new_n1159), .A3(new_n1161), .ZN(new_n1162));
  AOI21_X1  g737(.A(new_n1156), .B1(new_n1087), .B2(new_n1154), .ZN(new_n1163));
  OAI21_X1  g738(.A(KEYINPUT121), .B1(new_n1163), .B2(new_n1160), .ZN(new_n1164));
  NAND3_X1  g739(.A1(new_n1034), .A2(new_n1029), .A3(new_n995), .ZN(new_n1165));
  NAND2_X1  g740(.A1(new_n1165), .A2(KEYINPUT120), .ZN(new_n1166));
  INV_X1    g741(.A(KEYINPUT120), .ZN(new_n1167));
  NAND4_X1  g742(.A1(new_n1034), .A2(new_n1029), .A3(new_n1167), .A4(new_n995), .ZN(new_n1168));
  NAND2_X1  g743(.A1(new_n1166), .A2(new_n1168), .ZN(new_n1169));
  INV_X1    g744(.A(G1348), .ZN(new_n1170));
  AOI21_X1  g745(.A(new_n1169), .B1(new_n1170), .B2(new_n1078), .ZN(new_n1171));
  OAI211_X1 g746(.A(new_n1162), .B(new_n1164), .C1(new_n922), .C2(new_n1171), .ZN(new_n1172));
  INV_X1    g747(.A(KEYINPUT119), .ZN(new_n1173));
  OAI21_X1  g748(.A(new_n1173), .B1(new_n1158), .B2(new_n1161), .ZN(new_n1174));
  NAND3_X1  g749(.A1(new_n1163), .A2(KEYINPUT119), .A3(new_n1160), .ZN(new_n1175));
  NAND2_X1  g750(.A1(new_n1174), .A2(new_n1175), .ZN(new_n1176));
  NAND2_X1  g751(.A1(new_n1172), .A2(new_n1176), .ZN(new_n1177));
  INV_X1    g752(.A(KEYINPUT122), .ZN(new_n1178));
  AOI21_X1  g753(.A(new_n1178), .B1(new_n1158), .B2(new_n1161), .ZN(new_n1179));
  NOR3_X1   g754(.A1(new_n1163), .A2(KEYINPUT122), .A3(new_n1160), .ZN(new_n1180));
  NOR2_X1   g755(.A1(new_n1179), .A2(new_n1180), .ZN(new_n1181));
  AOI21_X1  g756(.A(KEYINPUT61), .B1(new_n1181), .B2(new_n1176), .ZN(new_n1182));
  INV_X1    g757(.A(KEYINPUT61), .ZN(new_n1183));
  AOI21_X1  g758(.A(new_n1183), .B1(new_n1163), .B2(new_n1160), .ZN(new_n1184));
  NAND3_X1  g759(.A1(new_n1164), .A2(new_n1162), .A3(new_n1184), .ZN(new_n1185));
  AOI21_X1  g760(.A(G1348), .B1(new_n1081), .B2(new_n1074), .ZN(new_n1186));
  INV_X1    g761(.A(KEYINPUT60), .ZN(new_n1187));
  NOR4_X1   g762(.A1(new_n1186), .A2(new_n1187), .A3(new_n609), .A4(new_n1169), .ZN(new_n1188));
  AOI21_X1  g763(.A(new_n922), .B1(new_n1171), .B2(KEYINPUT60), .ZN(new_n1189));
  OAI21_X1  g764(.A(new_n1187), .B1(new_n1186), .B2(new_n1169), .ZN(new_n1190));
  AOI21_X1  g765(.A(new_n1188), .B1(new_n1189), .B2(new_n1190), .ZN(new_n1191));
  INV_X1    g766(.A(KEYINPUT59), .ZN(new_n1192));
  NOR2_X1   g767(.A1(new_n1043), .A2(G1996), .ZN(new_n1193));
  XNOR2_X1  g768(.A(KEYINPUT58), .B(G1341), .ZN(new_n1194));
  AOI21_X1  g769(.A(new_n1194), .B1(new_n1034), .B2(new_n1029), .ZN(new_n1195));
  OAI211_X1 g770(.A(new_n1192), .B(new_n557), .C1(new_n1193), .C2(new_n1195), .ZN(new_n1196));
  AOI21_X1  g771(.A(new_n1195), .B1(new_n1087), .B2(new_n999), .ZN(new_n1197));
  OAI21_X1  g772(.A(KEYINPUT59), .B1(new_n1197), .B2(new_n556), .ZN(new_n1198));
  NAND2_X1  g773(.A1(new_n1196), .A2(new_n1198), .ZN(new_n1199));
  NAND3_X1  g774(.A1(new_n1185), .A2(new_n1191), .A3(new_n1199), .ZN(new_n1200));
  OAI21_X1  g775(.A(new_n1177), .B1(new_n1182), .B2(new_n1200), .ZN(new_n1201));
  INV_X1    g776(.A(KEYINPUT123), .ZN(new_n1202));
  AOI21_X1  g777(.A(new_n1153), .B1(new_n1201), .B2(new_n1202), .ZN(new_n1203));
  OAI211_X1 g778(.A(KEYINPUT123), .B(new_n1177), .C1(new_n1182), .C2(new_n1200), .ZN(new_n1204));
  AOI21_X1  g779(.A(new_n1140), .B1(new_n1203), .B2(new_n1204), .ZN(new_n1205));
  AOI21_X1  g780(.A(new_n1013), .B1(G1986), .B2(G290), .ZN(new_n1206));
  INV_X1    g781(.A(new_n1010), .ZN(new_n1207));
  AOI211_X1 g782(.A(new_n993), .B(new_n992), .C1(new_n1206), .C2(new_n1207), .ZN(new_n1208));
  OAI21_X1  g783(.A(new_n1018), .B1(new_n1205), .B2(new_n1208), .ZN(G329));
  assign    G231 = 1'b0;
  AND3_X1   g784(.A1(new_n675), .A2(new_n657), .A3(G319), .ZN(new_n1211));
  OAI21_X1  g785(.A(new_n1211), .B1(new_n714), .B2(new_n715), .ZN(new_n1212));
  AOI21_X1  g786(.A(new_n1212), .B1(new_n913), .B2(new_n915), .ZN(new_n1213));
  AOI21_X1  g787(.A(KEYINPUT127), .B1(new_n986), .B2(new_n1213), .ZN(new_n1214));
  AOI21_X1  g788(.A(new_n984), .B1(new_n965), .B2(new_n968), .ZN(new_n1215));
  INV_X1    g789(.A(new_n985), .ZN(new_n1216));
  OAI211_X1 g790(.A(KEYINPUT127), .B(new_n1213), .C1(new_n1215), .C2(new_n1216), .ZN(new_n1217));
  INV_X1    g791(.A(new_n1217), .ZN(new_n1218));
  NOR2_X1   g792(.A1(new_n1214), .A2(new_n1218), .ZN(G308));
  NAND2_X1  g793(.A1(new_n986), .A2(new_n1213), .ZN(G225));
endmodule


