//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 0 0 1 0 1 0 0 1 1 1 1 0 0 0 1 1 1 1 0 0 0 1 1 0 1 1 1 1 1 1 1 0 1 1 1 1 1 1 0 0 1 1 0 0 1 0 1 1 1 0 1 0 0 1 0 1 1 1 0 0 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:28:16 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n448, new_n451, new_n452, new_n453, new_n456, new_n457,
    new_n458, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n484, new_n485, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n528, new_n529, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n536, new_n537, new_n538, new_n539, new_n540,
    new_n541, new_n542, new_n545, new_n546, new_n547, new_n548, new_n549,
    new_n550, new_n551, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n564, new_n565, new_n567, new_n568,
    new_n569, new_n570, new_n571, new_n572, new_n573, new_n574, new_n575,
    new_n576, new_n577, new_n579, new_n580, new_n581, new_n583, new_n584,
    new_n585, new_n586, new_n587, new_n588, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n612, new_n613, new_n616, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n844, new_n845, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1169, new_n1170, new_n1171, new_n1172,
    new_n1173, new_n1174, new_n1175;
  XOR2_X1   g000(.A(KEYINPUT64), .B(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  XNOR2_X1  g004(.A(KEYINPUT65), .B(G1083), .ZN(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  XNOR2_X1  g011(.A(KEYINPUT66), .B(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(new_n448));
  XOR2_X1   g023(.A(new_n448), .B(KEYINPUT67), .Z(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G220), .A2(G221), .A3(G218), .A4(G219), .ZN(new_n451));
  XOR2_X1   g026(.A(new_n451), .B(KEYINPUT2), .Z(new_n452));
  NAND4_X1  g027(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n453));
  NOR2_X1   g028(.A1(new_n452), .A2(new_n453), .ZN(G325));
  INV_X1    g029(.A(G325), .ZN(G261));
  NAND2_X1  g030(.A1(new_n452), .A2(G2106), .ZN(new_n456));
  NAND2_X1  g031(.A1(new_n453), .A2(G567), .ZN(new_n457));
  NAND2_X1  g032(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  INV_X1    g033(.A(new_n458), .ZN(G319));
  AND2_X1   g034(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n460));
  NOR2_X1   g035(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n461));
  NOR2_X1   g036(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  INV_X1    g037(.A(G125), .ZN(new_n463));
  NOR2_X1   g038(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n464), .A2(KEYINPUT68), .ZN(new_n465));
  INV_X1    g040(.A(new_n465), .ZN(new_n466));
  NAND2_X1  g041(.A1(G113), .A2(G2104), .ZN(new_n467));
  OAI21_X1  g042(.A(new_n467), .B1(new_n464), .B2(KEYINPUT68), .ZN(new_n468));
  OAI21_X1  g043(.A(G2105), .B1(new_n466), .B2(new_n468), .ZN(new_n469));
  INV_X1    g044(.A(KEYINPUT69), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  OR2_X1    g046(.A1(new_n460), .A2(new_n461), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n472), .A2(G125), .ZN(new_n473));
  INV_X1    g048(.A(KEYINPUT68), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  NAND3_X1  g050(.A1(new_n475), .A2(new_n465), .A3(new_n467), .ZN(new_n476));
  NAND3_X1  g051(.A1(new_n476), .A2(KEYINPUT69), .A3(G2105), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n471), .A2(new_n477), .ZN(new_n478));
  INV_X1    g053(.A(G2105), .ZN(new_n479));
  OAI211_X1 g054(.A(G137), .B(new_n479), .C1(new_n460), .C2(new_n461), .ZN(new_n480));
  NAND3_X1  g055(.A1(new_n479), .A2(G101), .A3(G2104), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  INV_X1    g057(.A(KEYINPUT70), .ZN(new_n483));
  XNOR2_X1  g058(.A(new_n482), .B(new_n483), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n478), .A2(new_n484), .ZN(new_n485));
  INV_X1    g060(.A(new_n485), .ZN(G160));
  NOR2_X1   g061(.A1(new_n462), .A2(G2105), .ZN(new_n487));
  NAND2_X1  g062(.A1(new_n487), .A2(G136), .ZN(new_n488));
  NOR2_X1   g063(.A1(new_n462), .A2(new_n479), .ZN(new_n489));
  NAND2_X1  g064(.A1(new_n489), .A2(G124), .ZN(new_n490));
  INV_X1    g065(.A(G100), .ZN(new_n491));
  AND3_X1   g066(.A1(new_n491), .A2(new_n479), .A3(KEYINPUT71), .ZN(new_n492));
  AOI21_X1  g067(.A(KEYINPUT71), .B1(new_n491), .B2(new_n479), .ZN(new_n493));
  OAI221_X1 g068(.A(G2104), .B1(G112), .B2(new_n479), .C1(new_n492), .C2(new_n493), .ZN(new_n494));
  AND3_X1   g069(.A1(new_n488), .A2(new_n490), .A3(new_n494), .ZN(G162));
  OAI211_X1 g070(.A(G138), .B(new_n479), .C1(new_n460), .C2(new_n461), .ZN(new_n496));
  INV_X1    g071(.A(KEYINPUT4), .ZN(new_n497));
  OR2_X1    g072(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  NAND2_X1  g073(.A1(new_n489), .A2(G126), .ZN(new_n499));
  NAND2_X1  g074(.A1(new_n496), .A2(new_n497), .ZN(new_n500));
  OR2_X1    g075(.A1(G102), .A2(G2105), .ZN(new_n501));
  OAI211_X1 g076(.A(new_n501), .B(G2104), .C1(G114), .C2(new_n479), .ZN(new_n502));
  NAND4_X1  g077(.A1(new_n498), .A2(new_n499), .A3(new_n500), .A4(new_n502), .ZN(new_n503));
  INV_X1    g078(.A(new_n503), .ZN(G164));
  AND3_X1   g079(.A1(KEYINPUT73), .A2(KEYINPUT5), .A3(G543), .ZN(new_n505));
  AOI21_X1  g080(.A(KEYINPUT5), .B1(KEYINPUT73), .B2(G543), .ZN(new_n506));
  NOR2_X1   g081(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  INV_X1    g082(.A(KEYINPUT72), .ZN(new_n508));
  NOR2_X1   g083(.A1(new_n508), .A2(G651), .ZN(new_n509));
  INV_X1    g084(.A(G651), .ZN(new_n510));
  NOR2_X1   g085(.A1(new_n510), .A2(KEYINPUT72), .ZN(new_n511));
  OAI21_X1  g086(.A(KEYINPUT6), .B1(new_n509), .B2(new_n511), .ZN(new_n512));
  NOR2_X1   g087(.A1(KEYINPUT6), .A2(G651), .ZN(new_n513));
  INV_X1    g088(.A(new_n513), .ZN(new_n514));
  AOI21_X1  g089(.A(new_n507), .B1(new_n512), .B2(new_n514), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n515), .A2(G88), .ZN(new_n516));
  INV_X1    g091(.A(G543), .ZN(new_n517));
  AOI21_X1  g092(.A(new_n517), .B1(new_n512), .B2(new_n514), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n518), .A2(G50), .ZN(new_n519));
  NAND2_X1  g094(.A1(G75), .A2(G543), .ZN(new_n520));
  INV_X1    g095(.A(G62), .ZN(new_n521));
  OAI21_X1  g096(.A(new_n520), .B1(new_n507), .B2(new_n521), .ZN(new_n522));
  XNOR2_X1  g097(.A(KEYINPUT72), .B(G651), .ZN(new_n523));
  INV_X1    g098(.A(new_n523), .ZN(new_n524));
  NAND2_X1  g099(.A1(new_n522), .A2(new_n524), .ZN(new_n525));
  NAND3_X1  g100(.A1(new_n516), .A2(new_n519), .A3(new_n525), .ZN(G303));
  INV_X1    g101(.A(G303), .ZN(G166));
  INV_X1    g102(.A(KEYINPUT6), .ZN(new_n528));
  NAND2_X1  g103(.A1(new_n510), .A2(KEYINPUT72), .ZN(new_n529));
  NAND2_X1  g104(.A1(new_n508), .A2(G651), .ZN(new_n530));
  AOI21_X1  g105(.A(new_n528), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  OAI211_X1 g106(.A(G51), .B(G543), .C1(new_n531), .C2(new_n513), .ZN(new_n532));
  INV_X1    g107(.A(new_n506), .ZN(new_n533));
  NAND3_X1  g108(.A1(KEYINPUT73), .A2(KEYINPUT5), .A3(G543), .ZN(new_n534));
  NAND2_X1  g109(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  OAI211_X1 g110(.A(new_n535), .B(G89), .C1(new_n531), .C2(new_n513), .ZN(new_n536));
  AND2_X1   g111(.A1(G63), .A2(G651), .ZN(new_n537));
  NAND3_X1  g112(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n538));
  NAND2_X1  g113(.A1(new_n538), .A2(KEYINPUT7), .ZN(new_n539));
  INV_X1    g114(.A(KEYINPUT7), .ZN(new_n540));
  NAND4_X1  g115(.A1(new_n540), .A2(G76), .A3(G543), .A4(G651), .ZN(new_n541));
  AOI22_X1  g116(.A1(new_n535), .A2(new_n537), .B1(new_n539), .B2(new_n541), .ZN(new_n542));
  NAND3_X1  g117(.A1(new_n532), .A2(new_n536), .A3(new_n542), .ZN(G286));
  INV_X1    g118(.A(G286), .ZN(G168));
  OAI21_X1  g119(.A(new_n514), .B1(new_n523), .B2(new_n528), .ZN(new_n545));
  NAND3_X1  g120(.A1(new_n545), .A2(G52), .A3(G543), .ZN(new_n546));
  NAND3_X1  g121(.A1(new_n545), .A2(G90), .A3(new_n535), .ZN(new_n547));
  INV_X1    g122(.A(G64), .ZN(new_n548));
  AOI21_X1  g123(.A(new_n548), .B1(new_n533), .B2(new_n534), .ZN(new_n549));
  AND2_X1   g124(.A1(G77), .A2(G543), .ZN(new_n550));
  OAI21_X1  g125(.A(new_n524), .B1(new_n549), .B2(new_n550), .ZN(new_n551));
  NAND3_X1  g126(.A1(new_n546), .A2(new_n547), .A3(new_n551), .ZN(G301));
  INV_X1    g127(.A(G301), .ZN(G171));
  NAND3_X1  g128(.A1(new_n545), .A2(G43), .A3(G543), .ZN(new_n554));
  XNOR2_X1  g129(.A(KEYINPUT74), .B(G81), .ZN(new_n555));
  NAND3_X1  g130(.A1(new_n545), .A2(new_n535), .A3(new_n555), .ZN(new_n556));
  INV_X1    g131(.A(G56), .ZN(new_n557));
  AOI21_X1  g132(.A(new_n557), .B1(new_n533), .B2(new_n534), .ZN(new_n558));
  AND2_X1   g133(.A1(G68), .A2(G543), .ZN(new_n559));
  OAI21_X1  g134(.A(new_n524), .B1(new_n558), .B2(new_n559), .ZN(new_n560));
  AND3_X1   g135(.A1(new_n554), .A2(new_n556), .A3(new_n560), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n561), .A2(G860), .ZN(G153));
  NAND4_X1  g137(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g138(.A1(G1), .A2(G3), .ZN(new_n564));
  XNOR2_X1  g139(.A(new_n564), .B(KEYINPUT8), .ZN(new_n565));
  NAND4_X1  g140(.A1(G319), .A2(G483), .A3(G661), .A4(new_n565), .ZN(G188));
  OAI211_X1 g141(.A(G53), .B(G543), .C1(new_n531), .C2(new_n513), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n567), .A2(KEYINPUT9), .ZN(new_n568));
  INV_X1    g143(.A(KEYINPUT9), .ZN(new_n569));
  NAND4_X1  g144(.A1(new_n545), .A2(new_n569), .A3(G53), .A4(G543), .ZN(new_n570));
  NAND2_X1  g145(.A1(new_n568), .A2(new_n570), .ZN(new_n571));
  NAND2_X1  g146(.A1(G78), .A2(G543), .ZN(new_n572));
  INV_X1    g147(.A(G65), .ZN(new_n573));
  OAI21_X1  g148(.A(new_n572), .B1(new_n507), .B2(new_n573), .ZN(new_n574));
  AOI22_X1  g149(.A1(new_n515), .A2(G91), .B1(new_n574), .B2(G651), .ZN(new_n575));
  AND3_X1   g150(.A1(new_n571), .A2(KEYINPUT75), .A3(new_n575), .ZN(new_n576));
  AOI21_X1  g151(.A(KEYINPUT75), .B1(new_n571), .B2(new_n575), .ZN(new_n577));
  NOR2_X1   g152(.A1(new_n576), .A2(new_n577), .ZN(G299));
  NAND2_X1  g153(.A1(new_n518), .A2(G49), .ZN(new_n579));
  NAND2_X1  g154(.A1(new_n515), .A2(G87), .ZN(new_n580));
  OAI21_X1  g155(.A(G651), .B1(new_n535), .B2(G74), .ZN(new_n581));
  NAND3_X1  g156(.A1(new_n579), .A2(new_n580), .A3(new_n581), .ZN(G288));
  NAND2_X1  g157(.A1(new_n515), .A2(G86), .ZN(new_n583));
  NAND2_X1  g158(.A1(new_n518), .A2(G48), .ZN(new_n584));
  NAND2_X1  g159(.A1(G73), .A2(G543), .ZN(new_n585));
  INV_X1    g160(.A(G61), .ZN(new_n586));
  OAI21_X1  g161(.A(new_n585), .B1(new_n507), .B2(new_n586), .ZN(new_n587));
  NAND2_X1  g162(.A1(new_n587), .A2(new_n524), .ZN(new_n588));
  NAND3_X1  g163(.A1(new_n583), .A2(new_n584), .A3(new_n588), .ZN(G305));
  NAND2_X1  g164(.A1(new_n518), .A2(G47), .ZN(new_n590));
  NAND2_X1  g165(.A1(new_n515), .A2(G85), .ZN(new_n591));
  NAND2_X1  g166(.A1(G72), .A2(G543), .ZN(new_n592));
  INV_X1    g167(.A(G60), .ZN(new_n593));
  OAI21_X1  g168(.A(new_n592), .B1(new_n507), .B2(new_n593), .ZN(new_n594));
  NAND2_X1  g169(.A1(new_n594), .A2(new_n524), .ZN(new_n595));
  NAND3_X1  g170(.A1(new_n590), .A2(new_n591), .A3(new_n595), .ZN(G290));
  NAND2_X1  g171(.A1(G301), .A2(G868), .ZN(new_n597));
  NAND2_X1  g172(.A1(G79), .A2(G543), .ZN(new_n598));
  INV_X1    g173(.A(KEYINPUT76), .ZN(new_n599));
  XNOR2_X1  g174(.A(new_n598), .B(new_n599), .ZN(new_n600));
  AOI21_X1  g175(.A(new_n600), .B1(G66), .B2(new_n535), .ZN(new_n601));
  INV_X1    g176(.A(G54), .ZN(new_n602));
  OAI21_X1  g177(.A(G543), .B1(new_n531), .B2(new_n513), .ZN(new_n603));
  OAI22_X1  g178(.A1(new_n601), .A2(new_n510), .B1(new_n602), .B2(new_n603), .ZN(new_n604));
  OAI211_X1 g179(.A(new_n535), .B(G92), .C1(new_n531), .C2(new_n513), .ZN(new_n605));
  INV_X1    g180(.A(KEYINPUT10), .ZN(new_n606));
  NAND2_X1  g181(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  NAND3_X1  g182(.A1(new_n515), .A2(KEYINPUT10), .A3(G92), .ZN(new_n608));
  AOI21_X1  g183(.A(new_n604), .B1(new_n607), .B2(new_n608), .ZN(new_n609));
  OAI21_X1  g184(.A(new_n597), .B1(new_n609), .B2(G868), .ZN(G321));
  XOR2_X1   g185(.A(G321), .B(KEYINPUT77), .Z(G284));
  INV_X1    g186(.A(G868), .ZN(new_n612));
  NAND2_X1  g187(.A1(G299), .A2(new_n612), .ZN(new_n613));
  OAI21_X1  g188(.A(new_n613), .B1(new_n612), .B2(G168), .ZN(G297));
  OAI21_X1  g189(.A(new_n613), .B1(new_n612), .B2(G168), .ZN(G280));
  INV_X1    g190(.A(G559), .ZN(new_n616));
  OAI21_X1  g191(.A(new_n609), .B1(new_n616), .B2(G860), .ZN(G148));
  NAND3_X1  g192(.A1(new_n554), .A2(new_n556), .A3(new_n560), .ZN(new_n618));
  NAND2_X1  g193(.A1(new_n608), .A2(new_n607), .ZN(new_n619));
  OR2_X1    g194(.A1(new_n601), .A2(new_n510), .ZN(new_n620));
  NAND2_X1  g195(.A1(new_n518), .A2(G54), .ZN(new_n621));
  NAND3_X1  g196(.A1(new_n619), .A2(new_n620), .A3(new_n621), .ZN(new_n622));
  NOR2_X1   g197(.A1(new_n622), .A2(G559), .ZN(new_n623));
  XNOR2_X1  g198(.A(new_n623), .B(KEYINPUT78), .ZN(new_n624));
  MUX2_X1   g199(.A(new_n618), .B(new_n624), .S(G868), .Z(G323));
  XNOR2_X1  g200(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND3_X1  g201(.A1(new_n479), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n627));
  XNOR2_X1  g202(.A(new_n627), .B(KEYINPUT12), .ZN(new_n628));
  XNOR2_X1  g203(.A(KEYINPUT79), .B(KEYINPUT13), .ZN(new_n629));
  XNOR2_X1  g204(.A(new_n628), .B(new_n629), .ZN(new_n630));
  INV_X1    g205(.A(new_n630), .ZN(new_n631));
  INV_X1    g206(.A(G2100), .ZN(new_n632));
  NAND2_X1  g207(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  XNOR2_X1  g208(.A(new_n633), .B(KEYINPUT80), .ZN(new_n634));
  AOI22_X1  g209(.A1(G123), .A2(new_n489), .B1(new_n487), .B2(G135), .ZN(new_n635));
  INV_X1    g210(.A(KEYINPUT81), .ZN(new_n636));
  NOR3_X1   g211(.A1(new_n636), .A2(new_n479), .A3(G111), .ZN(new_n637));
  OAI21_X1  g212(.A(new_n636), .B1(new_n479), .B2(G111), .ZN(new_n638));
  OAI211_X1 g213(.A(new_n638), .B(G2104), .C1(G99), .C2(G2105), .ZN(new_n639));
  OAI21_X1  g214(.A(new_n635), .B1(new_n637), .B2(new_n639), .ZN(new_n640));
  XOR2_X1   g215(.A(KEYINPUT82), .B(G2096), .Z(new_n641));
  XNOR2_X1  g216(.A(new_n640), .B(new_n641), .ZN(new_n642));
  OAI211_X1 g217(.A(new_n634), .B(new_n642), .C1(new_n632), .C2(new_n631), .ZN(G156));
  XNOR2_X1  g218(.A(G2427), .B(G2438), .ZN(new_n644));
  XNOR2_X1  g219(.A(new_n644), .B(G2430), .ZN(new_n645));
  XNOR2_X1  g220(.A(KEYINPUT15), .B(G2435), .ZN(new_n646));
  OR2_X1    g221(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  NAND2_X1  g222(.A1(new_n645), .A2(new_n646), .ZN(new_n648));
  NAND3_X1  g223(.A1(new_n647), .A2(KEYINPUT14), .A3(new_n648), .ZN(new_n649));
  XNOR2_X1  g224(.A(G2451), .B(G2454), .ZN(new_n650));
  XNOR2_X1  g225(.A(new_n650), .B(KEYINPUT16), .ZN(new_n651));
  XNOR2_X1  g226(.A(new_n649), .B(new_n651), .ZN(new_n652));
  XNOR2_X1  g227(.A(G2443), .B(G2446), .ZN(new_n653));
  XOR2_X1   g228(.A(new_n652), .B(new_n653), .Z(new_n654));
  XNOR2_X1  g229(.A(G1341), .B(G1348), .ZN(new_n655));
  INV_X1    g230(.A(new_n655), .ZN(new_n656));
  OAI21_X1  g231(.A(G14), .B1(new_n654), .B2(new_n656), .ZN(new_n657));
  XNOR2_X1  g232(.A(new_n652), .B(new_n653), .ZN(new_n658));
  OAI21_X1  g233(.A(KEYINPUT83), .B1(new_n658), .B2(new_n655), .ZN(new_n659));
  INV_X1    g234(.A(KEYINPUT83), .ZN(new_n660));
  NAND3_X1  g235(.A1(new_n654), .A2(new_n660), .A3(new_n656), .ZN(new_n661));
  AOI21_X1  g236(.A(new_n657), .B1(new_n659), .B2(new_n661), .ZN(G401));
  INV_X1    g237(.A(KEYINPUT18), .ZN(new_n663));
  XOR2_X1   g238(.A(G2084), .B(G2090), .Z(new_n664));
  XNOR2_X1  g239(.A(G2067), .B(G2678), .ZN(new_n665));
  NAND2_X1  g240(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  NAND2_X1  g241(.A1(new_n666), .A2(KEYINPUT17), .ZN(new_n667));
  NOR2_X1   g242(.A1(new_n664), .A2(new_n665), .ZN(new_n668));
  OAI21_X1  g243(.A(new_n663), .B1(new_n667), .B2(new_n668), .ZN(new_n669));
  XNOR2_X1  g244(.A(new_n669), .B(new_n632), .ZN(new_n670));
  XOR2_X1   g245(.A(G2072), .B(G2078), .Z(new_n671));
  AOI21_X1  g246(.A(new_n671), .B1(new_n666), .B2(KEYINPUT18), .ZN(new_n672));
  XOR2_X1   g247(.A(new_n672), .B(G2096), .Z(new_n673));
  XNOR2_X1  g248(.A(new_n670), .B(new_n673), .ZN(G227));
  XNOR2_X1  g249(.A(G1971), .B(G1976), .ZN(new_n675));
  XNOR2_X1  g250(.A(KEYINPUT84), .B(KEYINPUT19), .ZN(new_n676));
  XNOR2_X1  g251(.A(new_n675), .B(new_n676), .ZN(new_n677));
  XNOR2_X1  g252(.A(G1956), .B(G2474), .ZN(new_n678));
  XNOR2_X1  g253(.A(G1961), .B(G1966), .ZN(new_n679));
  NAND3_X1  g254(.A1(new_n677), .A2(new_n678), .A3(new_n679), .ZN(new_n680));
  XNOR2_X1  g255(.A(new_n678), .B(new_n679), .ZN(new_n681));
  NOR2_X1   g256(.A1(new_n678), .A2(new_n679), .ZN(new_n682));
  NAND2_X1  g257(.A1(new_n677), .A2(new_n682), .ZN(new_n683));
  AND2_X1   g258(.A1(new_n683), .A2(KEYINPUT20), .ZN(new_n684));
  NOR2_X1   g259(.A1(new_n683), .A2(KEYINPUT20), .ZN(new_n685));
  OAI221_X1 g260(.A(new_n680), .B1(new_n677), .B2(new_n681), .C1(new_n684), .C2(new_n685), .ZN(new_n686));
  XNOR2_X1  g261(.A(G1981), .B(G1986), .ZN(new_n687));
  XNOR2_X1  g262(.A(new_n686), .B(new_n687), .ZN(new_n688));
  XNOR2_X1  g263(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n689));
  XNOR2_X1  g264(.A(new_n689), .B(KEYINPUT85), .ZN(new_n690));
  XNOR2_X1  g265(.A(new_n688), .B(new_n690), .ZN(new_n691));
  XNOR2_X1  g266(.A(G1991), .B(G1996), .ZN(new_n692));
  XNOR2_X1  g267(.A(new_n691), .B(new_n692), .ZN(new_n693));
  INV_X1    g268(.A(new_n693), .ZN(G229));
  INV_X1    g269(.A(G29), .ZN(new_n695));
  NAND2_X1  g270(.A1(new_n472), .A2(G127), .ZN(new_n696));
  NAND2_X1  g271(.A1(G115), .A2(G2104), .ZN(new_n697));
  AOI21_X1  g272(.A(new_n479), .B1(new_n696), .B2(new_n697), .ZN(new_n698));
  NAND3_X1  g273(.A1(new_n479), .A2(G103), .A3(G2104), .ZN(new_n699));
  XNOR2_X1  g274(.A(new_n699), .B(KEYINPUT93), .ZN(new_n700));
  XOR2_X1   g275(.A(KEYINPUT92), .B(KEYINPUT25), .Z(new_n701));
  XNOR2_X1  g276(.A(new_n700), .B(new_n701), .ZN(new_n702));
  NAND2_X1  g277(.A1(new_n487), .A2(G139), .ZN(new_n703));
  NAND2_X1  g278(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  INV_X1    g279(.A(KEYINPUT94), .ZN(new_n705));
  NAND2_X1  g280(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  NAND3_X1  g281(.A1(new_n702), .A2(KEYINPUT94), .A3(new_n703), .ZN(new_n707));
  AOI21_X1  g282(.A(new_n698), .B1(new_n706), .B2(new_n707), .ZN(new_n708));
  INV_X1    g283(.A(KEYINPUT95), .ZN(new_n709));
  NOR2_X1   g284(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  INV_X1    g285(.A(new_n710), .ZN(new_n711));
  NAND2_X1  g286(.A1(new_n708), .A2(new_n709), .ZN(new_n712));
  AOI21_X1  g287(.A(new_n695), .B1(new_n711), .B2(new_n712), .ZN(new_n713));
  INV_X1    g288(.A(G33), .ZN(new_n714));
  NOR2_X1   g289(.A1(new_n714), .A2(G29), .ZN(new_n715));
  OR3_X1    g290(.A1(new_n713), .A2(KEYINPUT96), .A3(new_n715), .ZN(new_n716));
  OAI21_X1  g291(.A(KEYINPUT96), .B1(new_n713), .B2(new_n715), .ZN(new_n717));
  NAND2_X1  g292(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  OR2_X1    g293(.A1(new_n718), .A2(G2072), .ZN(new_n719));
  NAND2_X1  g294(.A1(new_n718), .A2(G2072), .ZN(new_n720));
  XNOR2_X1  g295(.A(KEYINPUT31), .B(G11), .ZN(new_n721));
  XNOR2_X1  g296(.A(new_n721), .B(KEYINPUT99), .ZN(new_n722));
  INV_X1    g297(.A(KEYINPUT30), .ZN(new_n723));
  AND2_X1   g298(.A1(new_n723), .A2(G28), .ZN(new_n724));
  OAI21_X1  g299(.A(new_n695), .B1(new_n723), .B2(G28), .ZN(new_n725));
  OAI221_X1 g300(.A(new_n722), .B1(new_n724), .B2(new_n725), .C1(new_n640), .C2(new_n695), .ZN(new_n726));
  XNOR2_X1  g301(.A(new_n726), .B(KEYINPUT100), .ZN(new_n727));
  NAND2_X1  g302(.A1(G164), .A2(G29), .ZN(new_n728));
  OAI21_X1  g303(.A(new_n728), .B1(G27), .B2(G29), .ZN(new_n729));
  INV_X1    g304(.A(G2078), .ZN(new_n730));
  NOR2_X1   g305(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  AND2_X1   g306(.A1(new_n729), .A2(new_n730), .ZN(new_n732));
  NOR3_X1   g307(.A1(new_n727), .A2(new_n731), .A3(new_n732), .ZN(new_n733));
  NAND2_X1  g308(.A1(new_n695), .A2(G32), .ZN(new_n734));
  XOR2_X1   g309(.A(KEYINPUT98), .B(KEYINPUT26), .Z(new_n735));
  NAND3_X1  g310(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n736));
  XNOR2_X1  g311(.A(new_n735), .B(new_n736), .ZN(new_n737));
  NAND2_X1  g312(.A1(new_n489), .A2(G129), .ZN(new_n738));
  NAND2_X1  g313(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  NAND3_X1  g314(.A1(new_n479), .A2(G105), .A3(G2104), .ZN(new_n740));
  XOR2_X1   g315(.A(new_n740), .B(KEYINPUT97), .Z(new_n741));
  NAND2_X1  g316(.A1(new_n487), .A2(G141), .ZN(new_n742));
  NAND2_X1  g317(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  NOR2_X1   g318(.A1(new_n739), .A2(new_n743), .ZN(new_n744));
  OAI21_X1  g319(.A(new_n734), .B1(new_n744), .B2(new_n695), .ZN(new_n745));
  XOR2_X1   g320(.A(KEYINPUT27), .B(G1996), .Z(new_n746));
  XNOR2_X1  g321(.A(new_n745), .B(new_n746), .ZN(new_n747));
  NOR2_X1   g322(.A1(G29), .A2(G35), .ZN(new_n748));
  AOI21_X1  g323(.A(new_n748), .B1(G162), .B2(G29), .ZN(new_n749));
  XNOR2_X1  g324(.A(KEYINPUT29), .B(G2090), .ZN(new_n750));
  XNOR2_X1  g325(.A(new_n749), .B(new_n750), .ZN(new_n751));
  NOR2_X1   g326(.A1(new_n747), .A2(new_n751), .ZN(new_n752));
  NOR2_X1   g327(.A1(G5), .A2(G16), .ZN(new_n753));
  AOI21_X1  g328(.A(new_n753), .B1(G171), .B2(G16), .ZN(new_n754));
  OR2_X1    g329(.A1(new_n754), .A2(G1961), .ZN(new_n755));
  INV_X1    g330(.A(G16), .ZN(new_n756));
  NAND2_X1  g331(.A1(new_n756), .A2(G19), .ZN(new_n757));
  XNOR2_X1  g332(.A(new_n757), .B(KEYINPUT88), .ZN(new_n758));
  OAI21_X1  g333(.A(new_n758), .B1(new_n561), .B2(new_n756), .ZN(new_n759));
  XOR2_X1   g334(.A(KEYINPUT89), .B(G1341), .Z(new_n760));
  AOI22_X1  g335(.A1(new_n754), .A2(G1961), .B1(new_n759), .B2(new_n760), .ZN(new_n761));
  NAND4_X1  g336(.A1(new_n733), .A2(new_n752), .A3(new_n755), .A4(new_n761), .ZN(new_n762));
  NAND2_X1  g337(.A1(new_n695), .A2(G26), .ZN(new_n763));
  XOR2_X1   g338(.A(new_n763), .B(KEYINPUT28), .Z(new_n764));
  NAND2_X1  g339(.A1(new_n489), .A2(G128), .ZN(new_n765));
  XNOR2_X1  g340(.A(new_n765), .B(KEYINPUT90), .ZN(new_n766));
  NAND2_X1  g341(.A1(new_n487), .A2(G140), .ZN(new_n767));
  NOR2_X1   g342(.A1(new_n479), .A2(G116), .ZN(new_n768));
  OAI21_X1  g343(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n769));
  OAI211_X1 g344(.A(new_n766), .B(new_n767), .C1(new_n768), .C2(new_n769), .ZN(new_n770));
  AOI21_X1  g345(.A(new_n764), .B1(new_n770), .B2(G29), .ZN(new_n771));
  XNOR2_X1  g346(.A(KEYINPUT91), .B(G2067), .ZN(new_n772));
  XNOR2_X1  g347(.A(new_n771), .B(new_n772), .ZN(new_n773));
  NAND2_X1  g348(.A1(new_n756), .A2(G4), .ZN(new_n774));
  OAI21_X1  g349(.A(new_n774), .B1(new_n609), .B2(new_n756), .ZN(new_n775));
  INV_X1    g350(.A(G1348), .ZN(new_n776));
  XNOR2_X1  g351(.A(new_n775), .B(new_n776), .ZN(new_n777));
  NAND2_X1  g352(.A1(new_n756), .A2(G21), .ZN(new_n778));
  OAI21_X1  g353(.A(new_n778), .B1(G168), .B2(new_n756), .ZN(new_n779));
  NAND2_X1  g354(.A1(new_n779), .A2(G1966), .ZN(new_n780));
  OR2_X1    g355(.A1(new_n759), .A2(new_n760), .ZN(new_n781));
  NAND4_X1  g356(.A1(new_n773), .A2(new_n777), .A3(new_n780), .A4(new_n781), .ZN(new_n782));
  NOR2_X1   g357(.A1(new_n779), .A2(G1966), .ZN(new_n783));
  XOR2_X1   g358(.A(new_n783), .B(KEYINPUT101), .Z(new_n784));
  INV_X1    g359(.A(G2084), .ZN(new_n785));
  OAI21_X1  g360(.A(new_n695), .B1(KEYINPUT24), .B2(G34), .ZN(new_n786));
  AOI21_X1  g361(.A(new_n786), .B1(KEYINPUT24), .B2(G34), .ZN(new_n787));
  AOI21_X1  g362(.A(new_n787), .B1(new_n485), .B2(G29), .ZN(new_n788));
  OAI21_X1  g363(.A(new_n784), .B1(new_n785), .B2(new_n788), .ZN(new_n789));
  NOR3_X1   g364(.A1(new_n762), .A2(new_n782), .A3(new_n789), .ZN(new_n790));
  NAND2_X1  g365(.A1(new_n788), .A2(new_n785), .ZN(new_n791));
  XOR2_X1   g366(.A(new_n791), .B(KEYINPUT102), .Z(new_n792));
  NAND2_X1  g367(.A1(new_n756), .A2(G20), .ZN(new_n793));
  XOR2_X1   g368(.A(new_n793), .B(KEYINPUT23), .Z(new_n794));
  AOI21_X1  g369(.A(new_n794), .B1(G299), .B2(G16), .ZN(new_n795));
  XOR2_X1   g370(.A(new_n795), .B(G1956), .Z(new_n796));
  NOR2_X1   g371(.A1(new_n792), .A2(new_n796), .ZN(new_n797));
  NAND4_X1  g372(.A1(new_n719), .A2(new_n720), .A3(new_n790), .A4(new_n797), .ZN(new_n798));
  NAND2_X1  g373(.A1(new_n487), .A2(G131), .ZN(new_n799));
  NAND2_X1  g374(.A1(new_n489), .A2(G119), .ZN(new_n800));
  NOR2_X1   g375(.A1(new_n479), .A2(G107), .ZN(new_n801));
  OAI21_X1  g376(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n802));
  OAI211_X1 g377(.A(new_n799), .B(new_n800), .C1(new_n801), .C2(new_n802), .ZN(new_n803));
  MUX2_X1   g378(.A(G25), .B(new_n803), .S(G29), .Z(new_n804));
  XOR2_X1   g379(.A(KEYINPUT35), .B(G1991), .Z(new_n805));
  INV_X1    g380(.A(new_n805), .ZN(new_n806));
  XNOR2_X1  g381(.A(new_n804), .B(new_n806), .ZN(new_n807));
  AND2_X1   g382(.A1(new_n756), .A2(G24), .ZN(new_n808));
  AOI21_X1  g383(.A(new_n808), .B1(G290), .B2(G16), .ZN(new_n809));
  INV_X1    g384(.A(G1986), .ZN(new_n810));
  AND2_X1   g385(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  NOR2_X1   g386(.A1(new_n809), .A2(new_n810), .ZN(new_n812));
  NOR3_X1   g387(.A1(new_n807), .A2(new_n811), .A3(new_n812), .ZN(new_n813));
  INV_X1    g388(.A(new_n813), .ZN(new_n814));
  NAND2_X1  g389(.A1(new_n756), .A2(G23), .ZN(new_n815));
  INV_X1    g390(.A(G288), .ZN(new_n816));
  OAI21_X1  g391(.A(new_n815), .B1(new_n816), .B2(new_n756), .ZN(new_n817));
  OR2_X1    g392(.A1(new_n817), .A2(KEYINPUT86), .ZN(new_n818));
  NAND2_X1  g393(.A1(new_n817), .A2(KEYINPUT86), .ZN(new_n819));
  NAND2_X1  g394(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  XOR2_X1   g395(.A(KEYINPUT33), .B(G1976), .Z(new_n821));
  INV_X1    g396(.A(new_n821), .ZN(new_n822));
  NAND2_X1  g397(.A1(new_n820), .A2(new_n822), .ZN(new_n823));
  MUX2_X1   g398(.A(G6), .B(G305), .S(G16), .Z(new_n824));
  XOR2_X1   g399(.A(KEYINPUT32), .B(G1981), .Z(new_n825));
  XNOR2_X1  g400(.A(new_n824), .B(new_n825), .ZN(new_n826));
  NAND3_X1  g401(.A1(new_n818), .A2(new_n821), .A3(new_n819), .ZN(new_n827));
  NAND2_X1  g402(.A1(new_n756), .A2(G22), .ZN(new_n828));
  OAI21_X1  g403(.A(new_n828), .B1(G166), .B2(new_n756), .ZN(new_n829));
  INV_X1    g404(.A(G1971), .ZN(new_n830));
  XNOR2_X1  g405(.A(new_n829), .B(new_n830), .ZN(new_n831));
  NAND4_X1  g406(.A1(new_n823), .A2(new_n826), .A3(new_n827), .A4(new_n831), .ZN(new_n832));
  INV_X1    g407(.A(KEYINPUT87), .ZN(new_n833));
  XNOR2_X1  g408(.A(new_n832), .B(new_n833), .ZN(new_n834));
  INV_X1    g409(.A(KEYINPUT34), .ZN(new_n835));
  AOI21_X1  g410(.A(new_n814), .B1(new_n834), .B2(new_n835), .ZN(new_n836));
  XNOR2_X1  g411(.A(new_n832), .B(KEYINPUT87), .ZN(new_n837));
  NAND2_X1  g412(.A1(new_n837), .A2(KEYINPUT34), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n836), .A2(new_n838), .ZN(new_n839));
  NAND2_X1  g414(.A1(new_n839), .A2(KEYINPUT36), .ZN(new_n840));
  INV_X1    g415(.A(KEYINPUT36), .ZN(new_n841));
  NAND3_X1  g416(.A1(new_n836), .A2(new_n841), .A3(new_n838), .ZN(new_n842));
  AOI21_X1  g417(.A(new_n798), .B1(new_n840), .B2(new_n842), .ZN(G311));
  NAND2_X1  g418(.A1(new_n840), .A2(new_n842), .ZN(new_n844));
  INV_X1    g419(.A(new_n798), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n844), .A2(new_n845), .ZN(G150));
  NOR2_X1   g421(.A1(new_n622), .A2(new_n616), .ZN(new_n847));
  XNOR2_X1  g422(.A(new_n847), .B(KEYINPUT38), .ZN(new_n848));
  OAI211_X1 g423(.A(new_n535), .B(G93), .C1(new_n531), .C2(new_n513), .ZN(new_n849));
  OAI211_X1 g424(.A(G55), .B(G543), .C1(new_n531), .C2(new_n513), .ZN(new_n850));
  OAI21_X1  g425(.A(G67), .B1(new_n505), .B2(new_n506), .ZN(new_n851));
  NAND2_X1  g426(.A1(G80), .A2(G543), .ZN(new_n852));
  AOI21_X1  g427(.A(new_n523), .B1(new_n851), .B2(new_n852), .ZN(new_n853));
  OAI211_X1 g428(.A(new_n849), .B(new_n850), .C1(new_n853), .C2(KEYINPUT103), .ZN(new_n854));
  AND2_X1   g429(.A1(new_n853), .A2(KEYINPUT103), .ZN(new_n855));
  NOR2_X1   g430(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  NAND2_X1  g431(.A1(new_n856), .A2(new_n561), .ZN(new_n857));
  OAI21_X1  g432(.A(new_n618), .B1(new_n854), .B2(new_n855), .ZN(new_n858));
  NAND2_X1  g433(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  XNOR2_X1  g434(.A(new_n848), .B(new_n859), .ZN(new_n860));
  OR2_X1    g435(.A1(new_n860), .A2(KEYINPUT39), .ZN(new_n861));
  INV_X1    g436(.A(G860), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n860), .A2(KEYINPUT39), .ZN(new_n863));
  NAND3_X1  g438(.A1(new_n861), .A2(new_n862), .A3(new_n863), .ZN(new_n864));
  NOR2_X1   g439(.A1(new_n856), .A2(new_n862), .ZN(new_n865));
  XNOR2_X1  g440(.A(new_n865), .B(KEYINPUT37), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n864), .A2(new_n866), .ZN(G145));
  XNOR2_X1  g442(.A(new_n485), .B(new_n640), .ZN(new_n868));
  XOR2_X1   g443(.A(new_n868), .B(G162), .Z(new_n869));
  INV_X1    g444(.A(new_n744), .ZN(new_n870));
  INV_X1    g445(.A(new_n712), .ZN(new_n871));
  OAI21_X1  g446(.A(new_n870), .B1(new_n871), .B2(new_n710), .ZN(new_n872));
  NAND3_X1  g447(.A1(new_n711), .A2(new_n712), .A3(new_n744), .ZN(new_n873));
  AOI22_X1  g448(.A1(G130), .A2(new_n489), .B1(new_n487), .B2(G142), .ZN(new_n874));
  NOR3_X1   g449(.A1(new_n479), .A2(KEYINPUT104), .A3(G118), .ZN(new_n875));
  OAI21_X1  g450(.A(KEYINPUT104), .B1(new_n479), .B2(G118), .ZN(new_n876));
  OAI211_X1 g451(.A(new_n876), .B(G2104), .C1(G106), .C2(G2105), .ZN(new_n877));
  OAI21_X1  g452(.A(new_n874), .B1(new_n875), .B2(new_n877), .ZN(new_n878));
  XNOR2_X1  g453(.A(new_n878), .B(KEYINPUT106), .ZN(new_n879));
  XNOR2_X1  g454(.A(new_n879), .B(new_n803), .ZN(new_n880));
  INV_X1    g455(.A(new_n880), .ZN(new_n881));
  NAND3_X1  g456(.A1(new_n872), .A2(new_n873), .A3(new_n881), .ZN(new_n882));
  INV_X1    g457(.A(new_n882), .ZN(new_n883));
  AOI21_X1  g458(.A(new_n881), .B1(new_n872), .B2(new_n873), .ZN(new_n884));
  XNOR2_X1  g459(.A(new_n770), .B(new_n503), .ZN(new_n885));
  XNOR2_X1  g460(.A(new_n628), .B(KEYINPUT105), .ZN(new_n886));
  XNOR2_X1  g461(.A(new_n885), .B(new_n886), .ZN(new_n887));
  INV_X1    g462(.A(new_n887), .ZN(new_n888));
  NOR3_X1   g463(.A1(new_n883), .A2(new_n884), .A3(new_n888), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n872), .A2(new_n873), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n890), .A2(new_n880), .ZN(new_n891));
  AOI21_X1  g466(.A(new_n887), .B1(new_n891), .B2(new_n882), .ZN(new_n892));
  OAI21_X1  g467(.A(new_n869), .B1(new_n889), .B2(new_n892), .ZN(new_n893));
  INV_X1    g468(.A(G37), .ZN(new_n894));
  OAI21_X1  g469(.A(new_n888), .B1(new_n883), .B2(new_n884), .ZN(new_n895));
  INV_X1    g470(.A(new_n869), .ZN(new_n896));
  NAND3_X1  g471(.A1(new_n891), .A2(new_n887), .A3(new_n882), .ZN(new_n897));
  NAND3_X1  g472(.A1(new_n895), .A2(new_n896), .A3(new_n897), .ZN(new_n898));
  NAND3_X1  g473(.A1(new_n893), .A2(new_n894), .A3(new_n898), .ZN(new_n899));
  XNOR2_X1  g474(.A(new_n899), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g475(.A1(new_n816), .A2(G303), .ZN(new_n901));
  NAND2_X1  g476(.A1(G166), .A2(G288), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  NAND4_X1  g478(.A1(G305), .A2(new_n595), .A3(new_n590), .A4(new_n591), .ZN(new_n904));
  NAND4_X1  g479(.A1(G290), .A2(new_n588), .A3(new_n583), .A4(new_n584), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  NAND2_X1  g481(.A1(new_n903), .A2(new_n906), .ZN(new_n907));
  NAND4_X1  g482(.A1(new_n901), .A2(new_n902), .A3(new_n904), .A4(new_n905), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  XOR2_X1   g484(.A(new_n909), .B(KEYINPUT42), .Z(new_n910));
  INV_X1    g485(.A(KEYINPUT108), .ZN(new_n911));
  NOR2_X1   g486(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  XNOR2_X1  g487(.A(new_n624), .B(new_n859), .ZN(new_n913));
  INV_X1    g488(.A(KEYINPUT107), .ZN(new_n914));
  NOR3_X1   g489(.A1(new_n576), .A2(new_n622), .A3(new_n577), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n571), .A2(new_n575), .ZN(new_n916));
  INV_X1    g491(.A(KEYINPUT75), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  NAND3_X1  g493(.A1(new_n571), .A2(KEYINPUT75), .A3(new_n575), .ZN(new_n919));
  AOI21_X1  g494(.A(new_n609), .B1(new_n918), .B2(new_n919), .ZN(new_n920));
  OAI21_X1  g495(.A(new_n914), .B1(new_n915), .B2(new_n920), .ZN(new_n921));
  OAI21_X1  g496(.A(new_n622), .B1(new_n576), .B2(new_n577), .ZN(new_n922));
  NAND3_X1  g497(.A1(new_n918), .A2(new_n919), .A3(new_n609), .ZN(new_n923));
  NAND3_X1  g498(.A1(new_n922), .A2(new_n923), .A3(KEYINPUT107), .ZN(new_n924));
  NAND3_X1  g499(.A1(new_n913), .A2(new_n921), .A3(new_n924), .ZN(new_n925));
  AND3_X1   g500(.A1(new_n922), .A2(new_n923), .A3(KEYINPUT41), .ZN(new_n926));
  AOI21_X1  g501(.A(KEYINPUT41), .B1(new_n922), .B2(new_n923), .ZN(new_n927));
  NOR2_X1   g502(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  OAI21_X1  g503(.A(new_n925), .B1(new_n913), .B2(new_n928), .ZN(new_n929));
  AND2_X1   g504(.A1(new_n910), .A2(new_n911), .ZN(new_n930));
  AOI21_X1  g505(.A(new_n912), .B1(new_n929), .B2(new_n930), .ZN(new_n931));
  OAI21_X1  g506(.A(new_n931), .B1(new_n930), .B2(new_n929), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n932), .A2(G868), .ZN(new_n933));
  OAI21_X1  g508(.A(new_n933), .B1(G868), .B2(new_n856), .ZN(G295));
  OAI21_X1  g509(.A(new_n933), .B1(G868), .B2(new_n856), .ZN(G331));
  INV_X1    g510(.A(KEYINPUT44), .ZN(new_n936));
  NAND2_X1  g511(.A1(G168), .A2(G301), .ZN(new_n937));
  NAND4_X1  g512(.A1(G286), .A2(new_n551), .A3(new_n546), .A4(new_n547), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  INV_X1    g514(.A(new_n858), .ZN(new_n940));
  NOR3_X1   g515(.A1(new_n618), .A2(new_n854), .A3(new_n855), .ZN(new_n941));
  OAI21_X1  g516(.A(new_n939), .B1(new_n940), .B2(new_n941), .ZN(new_n942));
  NAND4_X1  g517(.A1(new_n857), .A2(new_n858), .A3(new_n938), .A4(new_n937), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  INV_X1    g519(.A(KEYINPUT41), .ZN(new_n945));
  OAI21_X1  g520(.A(new_n945), .B1(new_n915), .B2(new_n920), .ZN(new_n946));
  NAND3_X1  g521(.A1(new_n922), .A2(new_n923), .A3(KEYINPUT41), .ZN(new_n947));
  AOI21_X1  g522(.A(new_n944), .B1(new_n946), .B2(new_n947), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n922), .A2(new_n923), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n944), .A2(new_n949), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n950), .A2(new_n909), .ZN(new_n951));
  OAI21_X1  g526(.A(KEYINPUT110), .B1(new_n948), .B2(new_n951), .ZN(new_n952));
  INV_X1    g527(.A(new_n944), .ZN(new_n953));
  OAI21_X1  g528(.A(new_n953), .B1(new_n926), .B2(new_n927), .ZN(new_n954));
  INV_X1    g529(.A(KEYINPUT110), .ZN(new_n955));
  NAND4_X1  g530(.A1(new_n954), .A2(new_n955), .A3(new_n909), .A4(new_n950), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n952), .A2(new_n956), .ZN(new_n957));
  NAND3_X1  g532(.A1(new_n921), .A2(new_n924), .A3(new_n944), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n954), .A2(new_n958), .ZN(new_n959));
  AND3_X1   g534(.A1(new_n907), .A2(KEYINPUT109), .A3(new_n908), .ZN(new_n960));
  AOI21_X1  g535(.A(KEYINPUT109), .B1(new_n907), .B2(new_n908), .ZN(new_n961));
  NOR2_X1   g536(.A1(new_n960), .A2(new_n961), .ZN(new_n962));
  AOI21_X1  g537(.A(G37), .B1(new_n959), .B2(new_n962), .ZN(new_n963));
  INV_X1    g538(.A(KEYINPUT43), .ZN(new_n964));
  AND3_X1   g539(.A1(new_n957), .A2(new_n963), .A3(new_n964), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n954), .A2(new_n950), .ZN(new_n966));
  AOI21_X1  g541(.A(G37), .B1(new_n966), .B2(new_n962), .ZN(new_n967));
  AOI21_X1  g542(.A(new_n964), .B1(new_n957), .B2(new_n967), .ZN(new_n968));
  OAI21_X1  g543(.A(new_n936), .B1(new_n965), .B2(new_n968), .ZN(new_n969));
  NAND3_X1  g544(.A1(new_n957), .A2(new_n967), .A3(new_n964), .ZN(new_n970));
  AOI21_X1  g545(.A(new_n964), .B1(new_n957), .B2(new_n963), .ZN(new_n971));
  INV_X1    g546(.A(KEYINPUT111), .ZN(new_n972));
  OAI211_X1 g547(.A(KEYINPUT44), .B(new_n970), .C1(new_n971), .C2(new_n972), .ZN(new_n973));
  AOI211_X1 g548(.A(KEYINPUT111), .B(new_n964), .C1(new_n957), .C2(new_n963), .ZN(new_n974));
  OAI21_X1  g549(.A(new_n969), .B1(new_n973), .B2(new_n974), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n975), .A2(KEYINPUT112), .ZN(new_n976));
  INV_X1    g551(.A(KEYINPUT112), .ZN(new_n977));
  OAI211_X1 g552(.A(new_n977), .B(new_n969), .C1(new_n973), .C2(new_n974), .ZN(new_n978));
  NAND2_X1  g553(.A1(new_n976), .A2(new_n978), .ZN(G397));
  XNOR2_X1  g554(.A(new_n770), .B(G2067), .ZN(new_n980));
  AOI21_X1  g555(.A(new_n980), .B1(G1996), .B2(new_n870), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n484), .A2(G40), .ZN(new_n982));
  AOI21_X1  g557(.A(new_n982), .B1(new_n471), .B2(new_n477), .ZN(new_n983));
  INV_X1    g558(.A(G1384), .ZN(new_n984));
  AOI21_X1  g559(.A(KEYINPUT45), .B1(new_n503), .B2(new_n984), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n983), .A2(new_n985), .ZN(new_n986));
  NOR2_X1   g561(.A1(new_n981), .A2(new_n986), .ZN(new_n987));
  INV_X1    g562(.A(new_n986), .ZN(new_n988));
  INV_X1    g563(.A(G1996), .ZN(new_n989));
  NAND3_X1  g564(.A1(new_n988), .A2(KEYINPUT113), .A3(new_n989), .ZN(new_n990));
  INV_X1    g565(.A(KEYINPUT113), .ZN(new_n991));
  OAI21_X1  g566(.A(new_n991), .B1(new_n986), .B2(G1996), .ZN(new_n992));
  AOI21_X1  g567(.A(new_n870), .B1(new_n990), .B2(new_n992), .ZN(new_n993));
  NOR2_X1   g568(.A1(new_n987), .A2(new_n993), .ZN(new_n994));
  XNOR2_X1  g569(.A(new_n803), .B(new_n805), .ZN(new_n995));
  OAI21_X1  g570(.A(new_n994), .B1(new_n986), .B2(new_n995), .ZN(new_n996));
  XNOR2_X1  g571(.A(G290), .B(G1986), .ZN(new_n997));
  AOI21_X1  g572(.A(new_n996), .B1(new_n988), .B2(new_n997), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n503), .A2(new_n984), .ZN(new_n999));
  INV_X1    g574(.A(KEYINPUT45), .ZN(new_n1000));
  NOR2_X1   g575(.A1(new_n999), .A2(new_n1000), .ZN(new_n1001));
  NOR2_X1   g576(.A1(new_n1001), .A2(new_n985), .ZN(new_n1002));
  NAND3_X1  g577(.A1(new_n1002), .A2(new_n983), .A3(new_n730), .ZN(new_n1003));
  XOR2_X1   g578(.A(KEYINPUT122), .B(KEYINPUT53), .Z(new_n1004));
  NAND2_X1  g579(.A1(new_n999), .A2(KEYINPUT50), .ZN(new_n1005));
  INV_X1    g580(.A(KEYINPUT50), .ZN(new_n1006));
  NAND3_X1  g581(.A1(new_n503), .A2(new_n1006), .A3(new_n984), .ZN(new_n1007));
  NAND3_X1  g582(.A1(new_n983), .A2(new_n1005), .A3(new_n1007), .ZN(new_n1008));
  INV_X1    g583(.A(G1961), .ZN(new_n1009));
  AOI22_X1  g584(.A1(new_n1003), .A2(new_n1004), .B1(new_n1008), .B2(new_n1009), .ZN(new_n1010));
  INV_X1    g585(.A(new_n983), .ZN(new_n1011));
  XNOR2_X1  g586(.A(new_n999), .B(new_n1000), .ZN(new_n1012));
  NOR2_X1   g587(.A1(new_n1011), .A2(new_n1012), .ZN(new_n1013));
  NAND3_X1  g588(.A1(new_n1013), .A2(KEYINPUT53), .A3(new_n730), .ZN(new_n1014));
  NAND3_X1  g589(.A1(new_n1010), .A2(new_n1014), .A3(G301), .ZN(new_n1015));
  AND2_X1   g590(.A1(new_n1015), .A2(KEYINPUT54), .ZN(new_n1016));
  NOR2_X1   g591(.A1(new_n730), .A2(KEYINPUT124), .ZN(new_n1017));
  INV_X1    g592(.A(KEYINPUT124), .ZN(new_n1018));
  OAI21_X1  g593(.A(KEYINPUT53), .B1(new_n1018), .B2(G2078), .ZN(new_n1019));
  NOR3_X1   g594(.A1(new_n1001), .A2(new_n1017), .A3(new_n1019), .ZN(new_n1020));
  AOI21_X1  g595(.A(new_n982), .B1(G2105), .B2(new_n476), .ZN(new_n1021));
  INV_X1    g596(.A(new_n985), .ZN(new_n1022));
  AOI21_X1  g597(.A(KEYINPUT123), .B1(new_n1021), .B2(new_n1022), .ZN(new_n1023));
  INV_X1    g598(.A(new_n982), .ZN(new_n1024));
  AND4_X1   g599(.A1(KEYINPUT123), .A2(new_n1022), .A3(new_n469), .A4(new_n1024), .ZN(new_n1025));
  OAI21_X1  g600(.A(new_n1020), .B1(new_n1023), .B2(new_n1025), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n1010), .A2(new_n1026), .ZN(new_n1027));
  AOI21_X1  g602(.A(KEYINPUT125), .B1(new_n1027), .B2(G171), .ZN(new_n1028));
  INV_X1    g603(.A(KEYINPUT125), .ZN(new_n1029));
  AOI211_X1 g604(.A(new_n1029), .B(G301), .C1(new_n1010), .C2(new_n1026), .ZN(new_n1030));
  OAI21_X1  g605(.A(new_n1016), .B1(new_n1028), .B2(new_n1030), .ZN(new_n1031));
  INV_X1    g606(.A(KEYINPUT54), .ZN(new_n1032));
  NOR2_X1   g607(.A1(new_n1027), .A2(G171), .ZN(new_n1033));
  AOI21_X1  g608(.A(G301), .B1(new_n1010), .B2(new_n1014), .ZN(new_n1034));
  OAI21_X1  g609(.A(new_n1032), .B1(new_n1033), .B2(new_n1034), .ZN(new_n1035));
  NAND3_X1  g610(.A1(new_n983), .A2(new_n984), .A3(new_n503), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n816), .A2(G1976), .ZN(new_n1037));
  NAND3_X1  g612(.A1(new_n1036), .A2(G8), .A3(new_n1037), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n1038), .A2(KEYINPUT52), .ZN(new_n1039));
  INV_X1    g614(.A(G1976), .ZN(new_n1040));
  AOI21_X1  g615(.A(KEYINPUT52), .B1(G288), .B2(new_n1040), .ZN(new_n1041));
  NAND4_X1  g616(.A1(new_n1036), .A2(G8), .A3(new_n1037), .A4(new_n1041), .ZN(new_n1042));
  OR2_X1    g617(.A1(G305), .A2(G1981), .ZN(new_n1043));
  NAND2_X1  g618(.A1(G305), .A2(G1981), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n1043), .A2(new_n1044), .ZN(new_n1045));
  INV_X1    g620(.A(KEYINPUT49), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n1045), .A2(new_n1046), .ZN(new_n1047));
  NAND3_X1  g622(.A1(new_n1043), .A2(KEYINPUT49), .A3(new_n1044), .ZN(new_n1048));
  NAND4_X1  g623(.A1(new_n1047), .A2(new_n1036), .A3(G8), .A4(new_n1048), .ZN(new_n1049));
  AND3_X1   g624(.A1(new_n1039), .A2(new_n1042), .A3(new_n1049), .ZN(new_n1050));
  XOR2_X1   g625(.A(KEYINPUT114), .B(G2090), .Z(new_n1051));
  NAND4_X1  g626(.A1(new_n983), .A2(new_n1005), .A3(new_n1007), .A4(new_n1051), .ZN(new_n1052));
  INV_X1    g627(.A(new_n1052), .ZN(new_n1053));
  AOI21_X1  g628(.A(G1971), .B1(new_n1002), .B2(new_n983), .ZN(new_n1054));
  OAI21_X1  g629(.A(G8), .B1(new_n1053), .B2(new_n1054), .ZN(new_n1055));
  NAND2_X1  g630(.A1(G303), .A2(G8), .ZN(new_n1056));
  XNOR2_X1  g631(.A(new_n1056), .B(KEYINPUT55), .ZN(new_n1057));
  NAND2_X1  g632(.A1(new_n1055), .A2(new_n1057), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n1002), .A2(new_n983), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n1059), .A2(new_n830), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n1060), .A2(new_n1052), .ZN(new_n1061));
  INV_X1    g636(.A(new_n1057), .ZN(new_n1062));
  NAND3_X1  g637(.A1(new_n1061), .A2(G8), .A3(new_n1062), .ZN(new_n1063));
  AND3_X1   g638(.A1(new_n1050), .A2(new_n1058), .A3(new_n1063), .ZN(new_n1064));
  INV_X1    g639(.A(G8), .ZN(new_n1065));
  INV_X1    g640(.A(G1966), .ZN(new_n1066));
  OAI21_X1  g641(.A(new_n1066), .B1(new_n1011), .B2(new_n1012), .ZN(new_n1067));
  XOR2_X1   g642(.A(KEYINPUT116), .B(G2084), .Z(new_n1068));
  NAND4_X1  g643(.A1(new_n983), .A2(new_n1005), .A3(new_n1007), .A4(new_n1068), .ZN(new_n1069));
  AOI21_X1  g644(.A(new_n1065), .B1(new_n1067), .B2(new_n1069), .ZN(new_n1070));
  NAND2_X1  g645(.A1(G286), .A2(G8), .ZN(new_n1071));
  XNOR2_X1  g646(.A(new_n1071), .B(KEYINPUT121), .ZN(new_n1072));
  INV_X1    g647(.A(new_n1072), .ZN(new_n1073));
  NOR3_X1   g648(.A1(new_n1070), .A2(KEYINPUT51), .A3(new_n1073), .ZN(new_n1074));
  AND3_X1   g649(.A1(new_n983), .A2(new_n1005), .A3(new_n1007), .ZN(new_n1075));
  AOI22_X1  g650(.A1(new_n1075), .A2(new_n1068), .B1(new_n1059), .B2(new_n1066), .ZN(new_n1076));
  OAI21_X1  g651(.A(new_n1072), .B1(new_n1076), .B2(new_n1065), .ZN(new_n1077));
  INV_X1    g652(.A(KEYINPUT51), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n1067), .A2(new_n1069), .ZN(new_n1079));
  AOI21_X1  g654(.A(new_n1078), .B1(new_n1079), .B2(new_n1073), .ZN(new_n1080));
  AOI21_X1  g655(.A(new_n1074), .B1(new_n1077), .B2(new_n1080), .ZN(new_n1081));
  NAND4_X1  g656(.A1(new_n1031), .A2(new_n1035), .A3(new_n1064), .A4(new_n1081), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n1013), .A2(new_n989), .ZN(new_n1083));
  XOR2_X1   g658(.A(KEYINPUT58), .B(G1341), .Z(new_n1084));
  NAND2_X1  g659(.A1(new_n1036), .A2(new_n1084), .ZN(new_n1085));
  AOI21_X1  g660(.A(new_n618), .B1(new_n1083), .B2(new_n1085), .ZN(new_n1086));
  INV_X1    g661(.A(KEYINPUT119), .ZN(new_n1087));
  NOR3_X1   g662(.A1(new_n1086), .A2(new_n1087), .A3(KEYINPUT59), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n1086), .A2(new_n1087), .ZN(new_n1089));
  INV_X1    g664(.A(KEYINPUT59), .ZN(new_n1090));
  INV_X1    g665(.A(new_n1085), .ZN(new_n1091));
  NOR2_X1   g666(.A1(new_n1059), .A2(G1996), .ZN(new_n1092));
  OAI21_X1  g667(.A(new_n561), .B1(new_n1091), .B2(new_n1092), .ZN(new_n1093));
  AOI21_X1  g668(.A(new_n1090), .B1(new_n1093), .B2(KEYINPUT119), .ZN(new_n1094));
  AOI21_X1  g669(.A(new_n1088), .B1(new_n1089), .B2(new_n1094), .ZN(new_n1095));
  OAI22_X1  g670(.A1(new_n1075), .A2(G1348), .B1(G2067), .B2(new_n1036), .ZN(new_n1096));
  INV_X1    g671(.A(KEYINPUT60), .ZN(new_n1097));
  OR3_X1    g672(.A1(new_n1096), .A2(KEYINPUT120), .A3(new_n1097), .ZN(new_n1098));
  OAI21_X1  g673(.A(KEYINPUT120), .B1(new_n1096), .B2(new_n1097), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n1098), .A2(new_n1099), .ZN(new_n1100));
  AOI21_X1  g675(.A(new_n622), .B1(new_n1096), .B2(new_n1097), .ZN(new_n1101));
  INV_X1    g676(.A(new_n1101), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n1100), .A2(new_n1102), .ZN(new_n1103));
  XNOR2_X1  g678(.A(KEYINPUT56), .B(G2072), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n1013), .A2(new_n1104), .ZN(new_n1105));
  XOR2_X1   g680(.A(new_n916), .B(KEYINPUT57), .Z(new_n1106));
  XNOR2_X1  g681(.A(KEYINPUT118), .B(G1956), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n1008), .A2(new_n1107), .ZN(new_n1108));
  NAND3_X1  g683(.A1(new_n1105), .A2(new_n1106), .A3(new_n1108), .ZN(new_n1109));
  INV_X1    g684(.A(new_n1109), .ZN(new_n1110));
  AOI21_X1  g685(.A(new_n1106), .B1(new_n1105), .B2(new_n1108), .ZN(new_n1111));
  OAI21_X1  g686(.A(KEYINPUT61), .B1(new_n1110), .B2(new_n1111), .ZN(new_n1112));
  INV_X1    g687(.A(new_n1111), .ZN(new_n1113));
  INV_X1    g688(.A(KEYINPUT61), .ZN(new_n1114));
  NAND3_X1  g689(.A1(new_n1113), .A2(new_n1114), .A3(new_n1109), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n1112), .A2(new_n1115), .ZN(new_n1116));
  NAND3_X1  g691(.A1(new_n1098), .A2(new_n1101), .A3(new_n1099), .ZN(new_n1117));
  NAND4_X1  g692(.A1(new_n1095), .A2(new_n1103), .A3(new_n1116), .A4(new_n1117), .ZN(new_n1118));
  AND2_X1   g693(.A1(new_n1096), .A2(new_n609), .ZN(new_n1119));
  AOI21_X1  g694(.A(new_n1111), .B1(new_n1119), .B2(new_n1109), .ZN(new_n1120));
  AOI21_X1  g695(.A(new_n1082), .B1(new_n1118), .B2(new_n1120), .ZN(new_n1121));
  AOI211_X1 g696(.A(new_n1065), .B(G286), .C1(new_n1067), .C2(new_n1069), .ZN(new_n1122));
  NAND4_X1  g697(.A1(new_n1050), .A2(new_n1058), .A3(new_n1063), .A4(new_n1122), .ZN(new_n1123));
  XOR2_X1   g698(.A(KEYINPUT117), .B(KEYINPUT63), .Z(new_n1124));
  NAND2_X1  g699(.A1(new_n1123), .A2(new_n1124), .ZN(new_n1125));
  AOI21_X1  g700(.A(new_n1062), .B1(new_n1061), .B2(G8), .ZN(new_n1126));
  AOI211_X1 g701(.A(new_n1065), .B(new_n1057), .C1(new_n1060), .C2(new_n1052), .ZN(new_n1127));
  NOR2_X1   g702(.A1(new_n1126), .A2(new_n1127), .ZN(new_n1128));
  NOR2_X1   g703(.A1(KEYINPUT117), .A2(KEYINPUT63), .ZN(new_n1129));
  NAND4_X1  g704(.A1(new_n1128), .A2(new_n1050), .A3(new_n1122), .A4(new_n1129), .ZN(new_n1130));
  NAND3_X1  g705(.A1(new_n1049), .A2(new_n1040), .A3(new_n816), .ZN(new_n1131));
  NAND2_X1  g706(.A1(new_n1131), .A2(new_n1043), .ZN(new_n1132));
  NAND2_X1  g707(.A1(new_n1036), .A2(G8), .ZN(new_n1133));
  XNOR2_X1  g708(.A(new_n1133), .B(KEYINPUT115), .ZN(new_n1134));
  AOI22_X1  g709(.A1(new_n1050), .A2(new_n1127), .B1(new_n1132), .B2(new_n1134), .ZN(new_n1135));
  AND3_X1   g710(.A1(new_n1125), .A2(new_n1130), .A3(new_n1135), .ZN(new_n1136));
  OAI211_X1 g711(.A(new_n1078), .B(new_n1072), .C1(new_n1076), .C2(new_n1065), .ZN(new_n1137));
  NOR2_X1   g712(.A1(new_n1070), .A2(new_n1073), .ZN(new_n1138));
  OAI21_X1  g713(.A(KEYINPUT51), .B1(new_n1076), .B2(new_n1072), .ZN(new_n1139));
  OAI211_X1 g714(.A(KEYINPUT62), .B(new_n1137), .C1(new_n1138), .C2(new_n1139), .ZN(new_n1140));
  NAND2_X1  g715(.A1(new_n1140), .A2(KEYINPUT126), .ZN(new_n1141));
  OAI21_X1  g716(.A(new_n1137), .B1(new_n1138), .B2(new_n1139), .ZN(new_n1142));
  INV_X1    g717(.A(KEYINPUT62), .ZN(new_n1143));
  NAND2_X1  g718(.A1(new_n1142), .A2(new_n1143), .ZN(new_n1144));
  NAND2_X1  g719(.A1(new_n1077), .A2(new_n1080), .ZN(new_n1145));
  INV_X1    g720(.A(KEYINPUT126), .ZN(new_n1146));
  NAND4_X1  g721(.A1(new_n1145), .A2(new_n1146), .A3(KEYINPUT62), .A4(new_n1137), .ZN(new_n1147));
  AND4_X1   g722(.A1(new_n1034), .A2(new_n1050), .A3(new_n1058), .A4(new_n1063), .ZN(new_n1148));
  NAND4_X1  g723(.A1(new_n1141), .A2(new_n1144), .A3(new_n1147), .A4(new_n1148), .ZN(new_n1149));
  NAND2_X1  g724(.A1(new_n1136), .A2(new_n1149), .ZN(new_n1150));
  OAI21_X1  g725(.A(new_n998), .B1(new_n1121), .B2(new_n1150), .ZN(new_n1151));
  NOR4_X1   g726(.A1(new_n987), .A2(new_n993), .A3(new_n806), .A4(new_n803), .ZN(new_n1152));
  NOR2_X1   g727(.A1(new_n770), .A2(G2067), .ZN(new_n1153));
  OAI21_X1  g728(.A(new_n988), .B1(new_n1152), .B2(new_n1153), .ZN(new_n1154));
  NOR3_X1   g729(.A1(new_n986), .A2(G1986), .A3(G290), .ZN(new_n1155));
  XNOR2_X1  g730(.A(new_n1155), .B(KEYINPUT48), .ZN(new_n1156));
  NAND2_X1  g731(.A1(new_n990), .A2(new_n992), .ZN(new_n1157));
  INV_X1    g732(.A(KEYINPUT46), .ZN(new_n1158));
  XNOR2_X1  g733(.A(new_n1157), .B(new_n1158), .ZN(new_n1159));
  INV_X1    g734(.A(KEYINPUT47), .ZN(new_n1160));
  OAI21_X1  g735(.A(new_n988), .B1(new_n980), .B2(new_n870), .ZN(new_n1161));
  NAND3_X1  g736(.A1(new_n1159), .A2(new_n1160), .A3(new_n1161), .ZN(new_n1162));
  INV_X1    g737(.A(new_n1162), .ZN(new_n1163));
  AOI21_X1  g738(.A(new_n1160), .B1(new_n1159), .B2(new_n1161), .ZN(new_n1164));
  OAI221_X1 g739(.A(new_n1154), .B1(new_n996), .B2(new_n1156), .C1(new_n1163), .C2(new_n1164), .ZN(new_n1165));
  INV_X1    g740(.A(new_n1165), .ZN(new_n1166));
  NAND2_X1  g741(.A1(new_n1151), .A2(new_n1166), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g742(.A(KEYINPUT127), .ZN(new_n1169));
  NOR2_X1   g743(.A1(G227), .A2(new_n458), .ZN(new_n1170));
  INV_X1    g744(.A(new_n1170), .ZN(new_n1171));
  OAI21_X1  g745(.A(new_n1169), .B1(G401), .B2(new_n1171), .ZN(new_n1172));
  AND2_X1   g746(.A1(new_n661), .A2(new_n659), .ZN(new_n1173));
  OAI211_X1 g747(.A(KEYINPUT127), .B(new_n1170), .C1(new_n1173), .C2(new_n657), .ZN(new_n1174));
  AND3_X1   g748(.A1(new_n1172), .A2(new_n1174), .A3(new_n693), .ZN(new_n1175));
  OAI211_X1 g749(.A(new_n1175), .B(new_n899), .C1(new_n968), .C2(new_n965), .ZN(G225));
  INV_X1    g750(.A(G225), .ZN(G308));
endmodule


