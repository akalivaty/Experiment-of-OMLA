

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584;

  XNOR2_X1 U323 ( .A(n394), .B(n393), .ZN(n529) );
  XNOR2_X1 U324 ( .A(n432), .B(KEYINPUT119), .ZN(n433) );
  XNOR2_X1 U325 ( .A(n324), .B(n323), .ZN(n325) );
  NOR2_X1 U326 ( .A1(n384), .A2(n382), .ZN(n383) );
  XOR2_X1 U327 ( .A(G99GAT), .B(G85GAT), .Z(n344) );
  XNOR2_X1 U328 ( .A(n349), .B(KEYINPUT72), .ZN(n350) );
  XNOR2_X1 U329 ( .A(n309), .B(KEYINPUT66), .ZN(n310) );
  XNOR2_X1 U330 ( .A(n392), .B(KEYINPUT109), .ZN(n393) );
  XNOR2_X1 U331 ( .A(n351), .B(n350), .ZN(n355) );
  XNOR2_X1 U332 ( .A(n311), .B(n310), .ZN(n314) );
  XNOR2_X1 U333 ( .A(n407), .B(KEYINPUT54), .ZN(n408) );
  XNOR2_X1 U334 ( .A(n326), .B(n325), .ZN(n384) );
  XNOR2_X1 U335 ( .A(n454), .B(KEYINPUT121), .ZN(n563) );
  XNOR2_X1 U336 ( .A(n457), .B(KEYINPUT122), .ZN(n458) );
  XNOR2_X1 U337 ( .A(n459), .B(n458), .ZN(G1351GAT) );
  XOR2_X1 U338 ( .A(KEYINPUT6), .B(KEYINPUT1), .Z(n292) );
  XNOR2_X1 U339 ( .A(G127GAT), .B(G148GAT), .ZN(n291) );
  XNOR2_X1 U340 ( .A(n292), .B(n291), .ZN(n307) );
  XOR2_X1 U341 ( .A(G113GAT), .B(G1GAT), .Z(n333) );
  XOR2_X1 U342 ( .A(G85GAT), .B(G155GAT), .Z(n294) );
  XNOR2_X1 U343 ( .A(G29GAT), .B(G162GAT), .ZN(n293) );
  XNOR2_X1 U344 ( .A(n294), .B(n293), .ZN(n295) );
  XOR2_X1 U345 ( .A(n333), .B(n295), .Z(n297) );
  NAND2_X1 U346 ( .A1(G225GAT), .A2(G233GAT), .ZN(n296) );
  XNOR2_X1 U347 ( .A(n297), .B(n296), .ZN(n301) );
  XOR2_X1 U348 ( .A(G57GAT), .B(KEYINPUT4), .Z(n299) );
  XNOR2_X1 U349 ( .A(KEYINPUT94), .B(KEYINPUT5), .ZN(n298) );
  XNOR2_X1 U350 ( .A(n299), .B(n298), .ZN(n300) );
  XOR2_X1 U351 ( .A(n301), .B(n300), .Z(n305) );
  XNOR2_X1 U352 ( .A(G134GAT), .B(G120GAT), .ZN(n302) );
  XNOR2_X1 U353 ( .A(n302), .B(KEYINPUT0), .ZN(n447) );
  XNOR2_X1 U354 ( .A(G141GAT), .B(KEYINPUT3), .ZN(n303) );
  XNOR2_X1 U355 ( .A(n303), .B(KEYINPUT2), .ZN(n426) );
  XNOR2_X1 U356 ( .A(n447), .B(n426), .ZN(n304) );
  XNOR2_X1 U357 ( .A(n305), .B(n304), .ZN(n306) );
  XNOR2_X1 U358 ( .A(n307), .B(n306), .ZN(n530) );
  XNOR2_X1 U359 ( .A(G36GAT), .B(G190GAT), .ZN(n308) );
  XNOR2_X1 U360 ( .A(n308), .B(G218GAT), .ZN(n397) );
  XOR2_X1 U361 ( .A(n397), .B(n344), .Z(n311) );
  NAND2_X1 U362 ( .A1(G232GAT), .A2(G233GAT), .ZN(n309) );
  XNOR2_X1 U363 ( .A(G50GAT), .B(KEYINPUT75), .ZN(n312) );
  XNOR2_X1 U364 ( .A(n312), .B(G162GAT), .ZN(n413) );
  XOR2_X1 U365 ( .A(n413), .B(KEYINPUT11), .Z(n313) );
  XNOR2_X1 U366 ( .A(n314), .B(n313), .ZN(n326) );
  XOR2_X1 U367 ( .A(KEYINPUT69), .B(KEYINPUT7), .Z(n316) );
  XNOR2_X1 U368 ( .A(G43GAT), .B(G29GAT), .ZN(n315) );
  XNOR2_X1 U369 ( .A(n316), .B(n315), .ZN(n317) );
  XOR2_X1 U370 ( .A(KEYINPUT8), .B(n317), .Z(n330) );
  XOR2_X1 U371 ( .A(KEYINPUT67), .B(KEYINPUT76), .Z(n319) );
  XNOR2_X1 U372 ( .A(G106GAT), .B(G92GAT), .ZN(n318) );
  XNOR2_X1 U373 ( .A(n319), .B(n318), .ZN(n320) );
  XOR2_X1 U374 ( .A(n330), .B(n320), .Z(n324) );
  XOR2_X1 U375 ( .A(KEYINPUT77), .B(KEYINPUT10), .Z(n322) );
  XNOR2_X1 U376 ( .A(G134GAT), .B(KEYINPUT9), .ZN(n321) );
  XNOR2_X1 U377 ( .A(n322), .B(n321), .ZN(n323) );
  XOR2_X1 U378 ( .A(G15GAT), .B(G22GAT), .Z(n328) );
  XNOR2_X1 U379 ( .A(G197GAT), .B(G141GAT), .ZN(n327) );
  XNOR2_X1 U380 ( .A(n328), .B(n327), .ZN(n329) );
  XNOR2_X1 U381 ( .A(n330), .B(n329), .ZN(n341) );
  XOR2_X1 U382 ( .A(KEYINPUT30), .B(KEYINPUT68), .Z(n332) );
  XNOR2_X1 U383 ( .A(G169GAT), .B(G8GAT), .ZN(n331) );
  XNOR2_X1 U384 ( .A(n332), .B(n331), .ZN(n337) );
  XOR2_X1 U385 ( .A(G36GAT), .B(G50GAT), .Z(n335) );
  XNOR2_X1 U386 ( .A(n333), .B(KEYINPUT29), .ZN(n334) );
  XNOR2_X1 U387 ( .A(n335), .B(n334), .ZN(n336) );
  XOR2_X1 U388 ( .A(n337), .B(n336), .Z(n339) );
  NAND2_X1 U389 ( .A1(G229GAT), .A2(G233GAT), .ZN(n338) );
  XNOR2_X1 U390 ( .A(n339), .B(n338), .ZN(n340) );
  XNOR2_X1 U391 ( .A(n341), .B(n340), .ZN(n570) );
  XOR2_X1 U392 ( .A(KEYINPUT32), .B(KEYINPUT33), .Z(n343) );
  XNOR2_X1 U393 ( .A(KEYINPUT74), .B(KEYINPUT73), .ZN(n342) );
  XNOR2_X1 U394 ( .A(n343), .B(n342), .ZN(n348) );
  XOR2_X1 U395 ( .A(KEYINPUT31), .B(n344), .Z(n346) );
  XOR2_X1 U396 ( .A(G106GAT), .B(G148GAT), .Z(n421) );
  XNOR2_X1 U397 ( .A(G120GAT), .B(n421), .ZN(n345) );
  XNOR2_X1 U398 ( .A(n346), .B(n345), .ZN(n347) );
  XOR2_X1 U399 ( .A(n348), .B(n347), .Z(n351) );
  NAND2_X1 U400 ( .A1(G230GAT), .A2(G233GAT), .ZN(n349) );
  XOR2_X1 U401 ( .A(G64GAT), .B(G92GAT), .Z(n353) );
  XNOR2_X1 U402 ( .A(G176GAT), .B(G204GAT), .ZN(n352) );
  XNOR2_X1 U403 ( .A(n353), .B(n352), .ZN(n401) );
  XOR2_X1 U404 ( .A(n401), .B(KEYINPUT71), .Z(n354) );
  XNOR2_X1 U405 ( .A(n355), .B(n354), .ZN(n359) );
  XOR2_X1 U406 ( .A(KEYINPUT70), .B(KEYINPUT13), .Z(n357) );
  XNOR2_X1 U407 ( .A(G71GAT), .B(G78GAT), .ZN(n356) );
  XNOR2_X1 U408 ( .A(n357), .B(n356), .ZN(n358) );
  XNOR2_X1 U409 ( .A(G57GAT), .B(n358), .ZN(n379) );
  XNOR2_X1 U410 ( .A(n359), .B(n379), .ZN(n386) );
  XOR2_X1 U411 ( .A(KEYINPUT41), .B(KEYINPUT65), .Z(n360) );
  XNOR2_X1 U412 ( .A(n386), .B(n360), .ZN(n460) );
  NOR2_X1 U413 ( .A1(n570), .A2(n460), .ZN(n362) );
  XNOR2_X1 U414 ( .A(KEYINPUT46), .B(KEYINPUT107), .ZN(n361) );
  XNOR2_X1 U415 ( .A(n362), .B(n361), .ZN(n381) );
  XOR2_X1 U416 ( .A(KEYINPUT82), .B(KEYINPUT14), .Z(n364) );
  XNOR2_X1 U417 ( .A(G1GAT), .B(G64GAT), .ZN(n363) );
  XNOR2_X1 U418 ( .A(n364), .B(n363), .ZN(n368) );
  XOR2_X1 U419 ( .A(KEYINPUT84), .B(KEYINPUT15), .Z(n366) );
  XNOR2_X1 U420 ( .A(KEYINPUT12), .B(KEYINPUT81), .ZN(n365) );
  XNOR2_X1 U421 ( .A(n366), .B(n365), .ZN(n367) );
  XOR2_X1 U422 ( .A(n368), .B(n367), .Z(n373) );
  XOR2_X1 U423 ( .A(KEYINPUT80), .B(KEYINPUT83), .Z(n370) );
  NAND2_X1 U424 ( .A1(G231GAT), .A2(G233GAT), .ZN(n369) );
  XNOR2_X1 U425 ( .A(n370), .B(n369), .ZN(n371) );
  XNOR2_X1 U426 ( .A(KEYINPUT79), .B(n371), .ZN(n372) );
  XNOR2_X1 U427 ( .A(n373), .B(n372), .ZN(n376) );
  XOR2_X1 U428 ( .A(KEYINPUT78), .B(G211GAT), .Z(n375) );
  XNOR2_X1 U429 ( .A(G8GAT), .B(G183GAT), .ZN(n374) );
  XNOR2_X1 U430 ( .A(n375), .B(n374), .ZN(n398) );
  XOR2_X1 U431 ( .A(n376), .B(n398), .Z(n378) );
  XOR2_X1 U432 ( .A(G15GAT), .B(G127GAT), .Z(n440) );
  XOR2_X1 U433 ( .A(G22GAT), .B(G155GAT), .Z(n424) );
  XNOR2_X1 U434 ( .A(n440), .B(n424), .ZN(n377) );
  XNOR2_X1 U435 ( .A(n378), .B(n377), .ZN(n380) );
  XNOR2_X1 U436 ( .A(n380), .B(n379), .ZN(n579) );
  XNOR2_X1 U437 ( .A(n579), .B(KEYINPUT106), .ZN(n565) );
  NAND2_X1 U438 ( .A1(n381), .A2(n565), .ZN(n382) );
  XNOR2_X1 U439 ( .A(n383), .B(KEYINPUT47), .ZN(n391) );
  XOR2_X1 U440 ( .A(KEYINPUT36), .B(n384), .Z(n582) );
  NOR2_X1 U441 ( .A1(n582), .A2(n579), .ZN(n385) );
  XOR2_X1 U442 ( .A(KEYINPUT45), .B(n385), .Z(n387) );
  NOR2_X1 U443 ( .A1(n387), .A2(n386), .ZN(n388) );
  XNOR2_X1 U444 ( .A(n388), .B(KEYINPUT108), .ZN(n389) );
  NAND2_X1 U445 ( .A1(n389), .A2(n570), .ZN(n390) );
  NAND2_X1 U446 ( .A1(n391), .A2(n390), .ZN(n394) );
  XNOR2_X1 U447 ( .A(KEYINPUT48), .B(KEYINPUT64), .ZN(n392) );
  XOR2_X1 U448 ( .A(G197GAT), .B(KEYINPUT21), .Z(n427) );
  XOR2_X1 U449 ( .A(KEYINPUT95), .B(n427), .Z(n396) );
  NAND2_X1 U450 ( .A1(G226GAT), .A2(G233GAT), .ZN(n395) );
  XNOR2_X1 U451 ( .A(n396), .B(n395), .ZN(n405) );
  XOR2_X1 U452 ( .A(n398), .B(n397), .Z(n403) );
  XOR2_X1 U453 ( .A(KEYINPUT19), .B(KEYINPUT17), .Z(n400) );
  XNOR2_X1 U454 ( .A(G169GAT), .B(KEYINPUT18), .ZN(n399) );
  XNOR2_X1 U455 ( .A(n400), .B(n399), .ZN(n448) );
  XNOR2_X1 U456 ( .A(n448), .B(n401), .ZN(n402) );
  XNOR2_X1 U457 ( .A(n403), .B(n402), .ZN(n404) );
  XOR2_X1 U458 ( .A(n405), .B(n404), .Z(n495) );
  XNOR2_X1 U459 ( .A(n495), .B(KEYINPUT117), .ZN(n406) );
  NOR2_X1 U460 ( .A1(n529), .A2(n406), .ZN(n409) );
  INV_X1 U461 ( .A(KEYINPUT118), .ZN(n407) );
  XNOR2_X1 U462 ( .A(n409), .B(n408), .ZN(n410) );
  NOR2_X1 U463 ( .A1(n530), .A2(n410), .ZN(n569) );
  XOR2_X1 U464 ( .A(KEYINPUT90), .B(KEYINPUT91), .Z(n412) );
  XNOR2_X1 U465 ( .A(KEYINPUT24), .B(KEYINPUT92), .ZN(n411) );
  XNOR2_X1 U466 ( .A(n412), .B(n411), .ZN(n417) );
  XOR2_X1 U467 ( .A(G78GAT), .B(n413), .Z(n415) );
  NAND2_X1 U468 ( .A1(G228GAT), .A2(G233GAT), .ZN(n414) );
  XNOR2_X1 U469 ( .A(n415), .B(n414), .ZN(n416) );
  XNOR2_X1 U470 ( .A(n417), .B(n416), .ZN(n431) );
  XOR2_X1 U471 ( .A(KEYINPUT93), .B(KEYINPUT23), .Z(n419) );
  XNOR2_X1 U472 ( .A(G211GAT), .B(G204GAT), .ZN(n418) );
  XNOR2_X1 U473 ( .A(n419), .B(n418), .ZN(n420) );
  XOR2_X1 U474 ( .A(n420), .B(KEYINPUT22), .Z(n423) );
  XNOR2_X1 U475 ( .A(n421), .B(G218GAT), .ZN(n422) );
  XNOR2_X1 U476 ( .A(n423), .B(n422), .ZN(n425) );
  XOR2_X1 U477 ( .A(n425), .B(n424), .Z(n429) );
  XNOR2_X1 U478 ( .A(n427), .B(n426), .ZN(n428) );
  XNOR2_X1 U479 ( .A(n429), .B(n428), .ZN(n430) );
  XNOR2_X1 U480 ( .A(n431), .B(n430), .ZN(n470) );
  NAND2_X1 U481 ( .A1(n569), .A2(n470), .ZN(n434) );
  XOR2_X1 U482 ( .A(KEYINPUT120), .B(KEYINPUT55), .Z(n432) );
  XNOR2_X1 U483 ( .A(n434), .B(n433), .ZN(n453) );
  XOR2_X1 U484 ( .A(KEYINPUT86), .B(KEYINPUT87), .Z(n436) );
  XNOR2_X1 U485 ( .A(KEYINPUT89), .B(G71GAT), .ZN(n435) );
  XNOR2_X1 U486 ( .A(n436), .B(n435), .ZN(n452) );
  XOR2_X1 U487 ( .A(KEYINPUT88), .B(G99GAT), .Z(n438) );
  XNOR2_X1 U488 ( .A(G43GAT), .B(G190GAT), .ZN(n437) );
  XNOR2_X1 U489 ( .A(n438), .B(n437), .ZN(n439) );
  XOR2_X1 U490 ( .A(n440), .B(n439), .Z(n442) );
  NAND2_X1 U491 ( .A1(G227GAT), .A2(G233GAT), .ZN(n441) );
  XNOR2_X1 U492 ( .A(n442), .B(n441), .ZN(n446) );
  XOR2_X1 U493 ( .A(G176GAT), .B(G183GAT), .Z(n444) );
  XNOR2_X1 U494 ( .A(G113GAT), .B(KEYINPUT20), .ZN(n443) );
  XNOR2_X1 U495 ( .A(n444), .B(n443), .ZN(n445) );
  XOR2_X1 U496 ( .A(n446), .B(n445), .Z(n450) );
  XNOR2_X1 U497 ( .A(n448), .B(n447), .ZN(n449) );
  XNOR2_X1 U498 ( .A(n450), .B(n449), .ZN(n451) );
  XNOR2_X1 U499 ( .A(n452), .B(n451), .ZN(n535) );
  NAND2_X1 U500 ( .A1(n453), .A2(n535), .ZN(n454) );
  NAND2_X1 U501 ( .A1(n563), .A2(n384), .ZN(n459) );
  XOR2_X1 U502 ( .A(KEYINPUT123), .B(KEYINPUT124), .Z(n456) );
  XNOR2_X1 U503 ( .A(G190GAT), .B(KEYINPUT58), .ZN(n455) );
  XNOR2_X1 U504 ( .A(n456), .B(n455), .ZN(n457) );
  INV_X1 U505 ( .A(n460), .ZN(n553) );
  NAND2_X1 U506 ( .A1(n563), .A2(n553), .ZN(n463) );
  XOR2_X1 U507 ( .A(KEYINPUT56), .B(KEYINPUT57), .Z(n461) );
  XNOR2_X1 U508 ( .A(n461), .B(G176GAT), .ZN(n462) );
  XNOR2_X1 U509 ( .A(n463), .B(n462), .ZN(G1349GAT) );
  INV_X1 U510 ( .A(n530), .ZN(n515) );
  NOR2_X1 U511 ( .A1(n570), .A2(n386), .ZN(n491) );
  XNOR2_X1 U512 ( .A(KEYINPUT85), .B(KEYINPUT16), .ZN(n465) );
  NOR2_X1 U513 ( .A1(n384), .A2(n579), .ZN(n464) );
  XNOR2_X1 U514 ( .A(n465), .B(n464), .ZN(n477) );
  INV_X1 U515 ( .A(n535), .ZN(n520) );
  XOR2_X1 U516 ( .A(n470), .B(KEYINPUT28), .Z(n533) );
  XOR2_X1 U517 ( .A(n495), .B(KEYINPUT27), .Z(n528) );
  NOR2_X1 U518 ( .A1(n533), .A2(n528), .ZN(n466) );
  NAND2_X1 U519 ( .A1(n520), .A2(n466), .ZN(n467) );
  NAND2_X1 U520 ( .A1(n530), .A2(n467), .ZN(n476) );
  NAND2_X1 U521 ( .A1(n495), .A2(n535), .ZN(n468) );
  NAND2_X1 U522 ( .A1(n470), .A2(n468), .ZN(n469) );
  XOR2_X1 U523 ( .A(KEYINPUT25), .B(n469), .Z(n474) );
  NOR2_X1 U524 ( .A1(n535), .A2(n470), .ZN(n471) );
  XOR2_X1 U525 ( .A(n471), .B(KEYINPUT26), .Z(n567) );
  NOR2_X1 U526 ( .A1(n528), .A2(n567), .ZN(n472) );
  NOR2_X1 U527 ( .A1(n472), .A2(n530), .ZN(n473) );
  NAND2_X1 U528 ( .A1(n474), .A2(n473), .ZN(n475) );
  NAND2_X1 U529 ( .A1(n476), .A2(n475), .ZN(n488) );
  NOR2_X1 U530 ( .A1(n477), .A2(n488), .ZN(n504) );
  NAND2_X1 U531 ( .A1(n491), .A2(n504), .ZN(n486) );
  NOR2_X1 U532 ( .A1(n515), .A2(n486), .ZN(n479) );
  XNOR2_X1 U533 ( .A(KEYINPUT96), .B(KEYINPUT34), .ZN(n478) );
  XNOR2_X1 U534 ( .A(n479), .B(n478), .ZN(n480) );
  XOR2_X1 U535 ( .A(G1GAT), .B(n480), .Z(G1324GAT) );
  INV_X1 U536 ( .A(n495), .ZN(n517) );
  NOR2_X1 U537 ( .A1(n517), .A2(n486), .ZN(n481) );
  XOR2_X1 U538 ( .A(G8GAT), .B(n481), .Z(G1325GAT) );
  NOR2_X1 U539 ( .A1(n486), .A2(n520), .ZN(n485) );
  XOR2_X1 U540 ( .A(KEYINPUT97), .B(KEYINPUT98), .Z(n483) );
  XNOR2_X1 U541 ( .A(G15GAT), .B(KEYINPUT35), .ZN(n482) );
  XNOR2_X1 U542 ( .A(n483), .B(n482), .ZN(n484) );
  XNOR2_X1 U543 ( .A(n485), .B(n484), .ZN(G1326GAT) );
  INV_X1 U544 ( .A(n533), .ZN(n524) );
  NOR2_X1 U545 ( .A1(n524), .A2(n486), .ZN(n487) );
  XOR2_X1 U546 ( .A(G22GAT), .B(n487), .Z(G1327GAT) );
  XOR2_X1 U547 ( .A(G29GAT), .B(KEYINPUT39), .Z(n494) );
  NOR2_X1 U548 ( .A1(n582), .A2(n488), .ZN(n489) );
  NAND2_X1 U549 ( .A1(n489), .A2(n579), .ZN(n490) );
  XNOR2_X1 U550 ( .A(n490), .B(KEYINPUT37), .ZN(n514) );
  NAND2_X1 U551 ( .A1(n491), .A2(n514), .ZN(n492) );
  XOR2_X1 U552 ( .A(KEYINPUT38), .B(n492), .Z(n500) );
  NAND2_X1 U553 ( .A1(n500), .A2(n530), .ZN(n493) );
  XNOR2_X1 U554 ( .A(n494), .B(n493), .ZN(G1328GAT) );
  NAND2_X1 U555 ( .A1(n500), .A2(n495), .ZN(n496) );
  XNOR2_X1 U556 ( .A(n496), .B(G36GAT), .ZN(G1329GAT) );
  XOR2_X1 U557 ( .A(KEYINPUT40), .B(KEYINPUT99), .Z(n498) );
  NAND2_X1 U558 ( .A1(n500), .A2(n535), .ZN(n497) );
  XNOR2_X1 U559 ( .A(n498), .B(n497), .ZN(n499) );
  XNOR2_X1 U560 ( .A(G43GAT), .B(n499), .ZN(G1330GAT) );
  NAND2_X1 U561 ( .A1(n500), .A2(n533), .ZN(n501) );
  XNOR2_X1 U562 ( .A(n501), .B(G50GAT), .ZN(G1331GAT) );
  XOR2_X1 U563 ( .A(KEYINPUT101), .B(KEYINPUT42), .Z(n503) );
  XNOR2_X1 U564 ( .A(G57GAT), .B(KEYINPUT100), .ZN(n502) );
  XNOR2_X1 U565 ( .A(n503), .B(n502), .ZN(n506) );
  INV_X1 U566 ( .A(n570), .ZN(n561) );
  NOR2_X1 U567 ( .A1(n561), .A2(n460), .ZN(n513) );
  NAND2_X1 U568 ( .A1(n513), .A2(n504), .ZN(n509) );
  NOR2_X1 U569 ( .A1(n515), .A2(n509), .ZN(n505) );
  XOR2_X1 U570 ( .A(n506), .B(n505), .Z(G1332GAT) );
  NOR2_X1 U571 ( .A1(n517), .A2(n509), .ZN(n507) );
  XOR2_X1 U572 ( .A(G64GAT), .B(n507), .Z(G1333GAT) );
  NOR2_X1 U573 ( .A1(n520), .A2(n509), .ZN(n508) );
  XOR2_X1 U574 ( .A(G71GAT), .B(n508), .Z(G1334GAT) );
  NOR2_X1 U575 ( .A1(n524), .A2(n509), .ZN(n511) );
  XNOR2_X1 U576 ( .A(KEYINPUT43), .B(KEYINPUT102), .ZN(n510) );
  XNOR2_X1 U577 ( .A(n511), .B(n510), .ZN(n512) );
  XNOR2_X1 U578 ( .A(G78GAT), .B(n512), .ZN(G1335GAT) );
  NAND2_X1 U579 ( .A1(n514), .A2(n513), .ZN(n523) );
  NOR2_X1 U580 ( .A1(n515), .A2(n523), .ZN(n516) );
  XOR2_X1 U581 ( .A(G85GAT), .B(n516), .Z(G1336GAT) );
  NOR2_X1 U582 ( .A1(n517), .A2(n523), .ZN(n519) );
  XNOR2_X1 U583 ( .A(G92GAT), .B(KEYINPUT103), .ZN(n518) );
  XNOR2_X1 U584 ( .A(n519), .B(n518), .ZN(G1337GAT) );
  NOR2_X1 U585 ( .A1(n520), .A2(n523), .ZN(n521) );
  XOR2_X1 U586 ( .A(KEYINPUT104), .B(n521), .Z(n522) );
  XNOR2_X1 U587 ( .A(G99GAT), .B(n522), .ZN(G1338GAT) );
  NOR2_X1 U588 ( .A1(n524), .A2(n523), .ZN(n526) );
  XNOR2_X1 U589 ( .A(KEYINPUT44), .B(KEYINPUT105), .ZN(n525) );
  XNOR2_X1 U590 ( .A(n526), .B(n525), .ZN(n527) );
  XNOR2_X1 U591 ( .A(G106GAT), .B(n527), .ZN(G1339GAT) );
  NOR2_X1 U592 ( .A1(n529), .A2(n528), .ZN(n531) );
  NAND2_X1 U593 ( .A1(n531), .A2(n530), .ZN(n532) );
  XNOR2_X1 U594 ( .A(KEYINPUT110), .B(n532), .ZN(n548) );
  NOR2_X1 U595 ( .A1(n548), .A2(n533), .ZN(n534) );
  NAND2_X1 U596 ( .A1(n535), .A2(n534), .ZN(n536) );
  XNOR2_X1 U597 ( .A(n536), .B(KEYINPUT111), .ZN(n544) );
  NAND2_X1 U598 ( .A1(n544), .A2(n561), .ZN(n537) );
  XNOR2_X1 U599 ( .A(G113GAT), .B(n537), .ZN(G1340GAT) );
  XOR2_X1 U600 ( .A(G120GAT), .B(KEYINPUT49), .Z(n539) );
  NAND2_X1 U601 ( .A1(n544), .A2(n553), .ZN(n538) );
  XNOR2_X1 U602 ( .A(n539), .B(n538), .ZN(G1341GAT) );
  INV_X1 U603 ( .A(n544), .ZN(n540) );
  NOR2_X1 U604 ( .A1(n565), .A2(n540), .ZN(n542) );
  XNOR2_X1 U605 ( .A(KEYINPUT50), .B(KEYINPUT112), .ZN(n541) );
  XNOR2_X1 U606 ( .A(n542), .B(n541), .ZN(n543) );
  XOR2_X1 U607 ( .A(G127GAT), .B(n543), .Z(G1342GAT) );
  XOR2_X1 U608 ( .A(KEYINPUT51), .B(KEYINPUT113), .Z(n546) );
  NAND2_X1 U609 ( .A1(n544), .A2(n384), .ZN(n545) );
  XNOR2_X1 U610 ( .A(n546), .B(n545), .ZN(n547) );
  XOR2_X1 U611 ( .A(G134GAT), .B(n547), .Z(G1343GAT) );
  NOR2_X1 U612 ( .A1(n548), .A2(n567), .ZN(n559) );
  NAND2_X1 U613 ( .A1(n559), .A2(n561), .ZN(n549) );
  XNOR2_X1 U614 ( .A(G141GAT), .B(n549), .ZN(G1344GAT) );
  XOR2_X1 U615 ( .A(KEYINPUT53), .B(KEYINPUT115), .Z(n551) );
  XNOR2_X1 U616 ( .A(G148GAT), .B(KEYINPUT52), .ZN(n550) );
  XNOR2_X1 U617 ( .A(n551), .B(n550), .ZN(n552) );
  XOR2_X1 U618 ( .A(KEYINPUT114), .B(n552), .Z(n555) );
  NAND2_X1 U619 ( .A1(n559), .A2(n553), .ZN(n554) );
  XNOR2_X1 U620 ( .A(n555), .B(n554), .ZN(G1345GAT) );
  XNOR2_X1 U621 ( .A(G155GAT), .B(KEYINPUT116), .ZN(n558) );
  INV_X1 U622 ( .A(n579), .ZN(n556) );
  NAND2_X1 U623 ( .A1(n559), .A2(n556), .ZN(n557) );
  XNOR2_X1 U624 ( .A(n558), .B(n557), .ZN(G1346GAT) );
  NAND2_X1 U625 ( .A1(n559), .A2(n384), .ZN(n560) );
  XNOR2_X1 U626 ( .A(n560), .B(G162GAT), .ZN(G1347GAT) );
  NAND2_X1 U627 ( .A1(n561), .A2(n563), .ZN(n562) );
  XNOR2_X1 U628 ( .A(n562), .B(G169GAT), .ZN(G1348GAT) );
  INV_X1 U629 ( .A(n563), .ZN(n564) );
  NOR2_X1 U630 ( .A1(n565), .A2(n564), .ZN(n566) );
  XOR2_X1 U631 ( .A(G183GAT), .B(n566), .Z(G1350GAT) );
  INV_X1 U632 ( .A(n567), .ZN(n568) );
  NAND2_X1 U633 ( .A1(n569), .A2(n568), .ZN(n581) );
  NOR2_X1 U634 ( .A1(n581), .A2(n570), .ZN(n574) );
  XOR2_X1 U635 ( .A(KEYINPUT60), .B(KEYINPUT59), .Z(n572) );
  XNOR2_X1 U636 ( .A(G197GAT), .B(KEYINPUT125), .ZN(n571) );
  XNOR2_X1 U637 ( .A(n572), .B(n571), .ZN(n573) );
  XNOR2_X1 U638 ( .A(n574), .B(n573), .ZN(G1352GAT) );
  XOR2_X1 U639 ( .A(KEYINPUT61), .B(KEYINPUT126), .Z(n577) );
  INV_X1 U640 ( .A(n581), .ZN(n575) );
  NAND2_X1 U641 ( .A1(n575), .A2(n386), .ZN(n576) );
  XNOR2_X1 U642 ( .A(n577), .B(n576), .ZN(n578) );
  XNOR2_X1 U643 ( .A(G204GAT), .B(n578), .ZN(G1353GAT) );
  NOR2_X1 U644 ( .A1(n579), .A2(n581), .ZN(n580) );
  XOR2_X1 U645 ( .A(G211GAT), .B(n580), .Z(G1354GAT) );
  NOR2_X1 U646 ( .A1(n582), .A2(n581), .ZN(n583) );
  XOR2_X1 U647 ( .A(KEYINPUT62), .B(n583), .Z(n584) );
  XNOR2_X1 U648 ( .A(G218GAT), .B(n584), .ZN(G1355GAT) );
endmodule

