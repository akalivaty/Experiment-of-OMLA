//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 1 1 1 0 0 0 0 0 0 1 0 0 1 0 1 1 0 1 1 1 0 0 0 1 0 0 1 0 0 1 0 1 1 0 1 1 0 0 0 0 1 1 1 0 1 0 0 1 1 1 1 0 0 1 0 0 1 1 0 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:18:25 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n712, new_n713, new_n714,
    new_n715, new_n716, new_n717, new_n718, new_n720, new_n721, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n741, new_n742, new_n743, new_n744, new_n745,
    new_n746, new_n747, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n774, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n782, new_n783, new_n784,
    new_n785, new_n787, new_n788, new_n789, new_n791, new_n792, new_n793,
    new_n795, new_n796, new_n797, new_n798, new_n799, new_n800, new_n801,
    new_n802, new_n803, new_n804, new_n805, new_n806, new_n807, new_n808,
    new_n809, new_n810, new_n811, new_n812, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n824,
    new_n825, new_n826, new_n827, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n885, new_n886, new_n888, new_n889, new_n890, new_n892,
    new_n893, new_n894, new_n895, new_n896, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n949, new_n950,
    new_n951, new_n952, new_n953, new_n954, new_n955, new_n956, new_n957,
    new_n958, new_n959, new_n960, new_n961, new_n962, new_n963, new_n964,
    new_n965, new_n967, new_n968, new_n969, new_n971, new_n972, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n993, new_n994, new_n996, new_n997,
    new_n998, new_n1000, new_n1001, new_n1002, new_n1004, new_n1005,
    new_n1006, new_n1007, new_n1008, new_n1009, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1021, new_n1022, new_n1023, new_n1024, new_n1025,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032;
  INV_X1    g000(.A(KEYINPUT17), .ZN(new_n202));
  INV_X1    g001(.A(G43gat), .ZN(new_n203));
  NOR2_X1   g002(.A1(new_n203), .A2(G50gat), .ZN(new_n204));
  INV_X1    g003(.A(G50gat), .ZN(new_n205));
  NOR2_X1   g004(.A1(new_n205), .A2(G43gat), .ZN(new_n206));
  OAI21_X1  g005(.A(KEYINPUT89), .B1(new_n204), .B2(new_n206), .ZN(new_n207));
  NAND2_X1  g006(.A1(new_n205), .A2(G43gat), .ZN(new_n208));
  NAND2_X1  g007(.A1(new_n203), .A2(G50gat), .ZN(new_n209));
  INV_X1    g008(.A(KEYINPUT89), .ZN(new_n210));
  NAND3_X1  g009(.A1(new_n208), .A2(new_n209), .A3(new_n210), .ZN(new_n211));
  NAND3_X1  g010(.A1(new_n207), .A2(KEYINPUT15), .A3(new_n211), .ZN(new_n212));
  INV_X1    g011(.A(G29gat), .ZN(new_n213));
  INV_X1    g012(.A(G36gat), .ZN(new_n214));
  NAND3_X1  g013(.A1(new_n213), .A2(new_n214), .A3(KEYINPUT90), .ZN(new_n215));
  INV_X1    g014(.A(KEYINPUT90), .ZN(new_n216));
  OAI21_X1  g015(.A(new_n216), .B1(G29gat), .B2(G36gat), .ZN(new_n217));
  NAND3_X1  g016(.A1(new_n215), .A2(new_n217), .A3(KEYINPUT14), .ZN(new_n218));
  NAND2_X1  g017(.A1(G29gat), .A2(G36gat), .ZN(new_n219));
  INV_X1    g018(.A(KEYINPUT14), .ZN(new_n220));
  OAI211_X1 g019(.A(new_n216), .B(new_n220), .C1(G29gat), .C2(G36gat), .ZN(new_n221));
  NAND3_X1  g020(.A1(new_n218), .A2(new_n219), .A3(new_n221), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n212), .A2(new_n222), .ZN(new_n223));
  INV_X1    g022(.A(KEYINPUT15), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n208), .A2(new_n209), .ZN(new_n225));
  AOI21_X1  g024(.A(new_n224), .B1(new_n225), .B2(KEYINPUT89), .ZN(new_n226));
  XNOR2_X1  g025(.A(KEYINPUT91), .B(G50gat), .ZN(new_n227));
  OAI21_X1  g026(.A(new_n208), .B1(new_n227), .B2(G43gat), .ZN(new_n228));
  AOI22_X1  g027(.A1(new_n211), .A2(new_n226), .B1(new_n228), .B2(new_n224), .ZN(new_n229));
  OAI211_X1 g028(.A(new_n202), .B(new_n223), .C1(new_n229), .C2(new_n222), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n205), .A2(KEYINPUT91), .ZN(new_n231));
  INV_X1    g030(.A(KEYINPUT91), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n232), .A2(G50gat), .ZN(new_n233));
  AOI21_X1  g032(.A(G43gat), .B1(new_n231), .B2(new_n233), .ZN(new_n234));
  OAI21_X1  g033(.A(new_n224), .B1(new_n234), .B2(new_n204), .ZN(new_n235));
  AOI21_X1  g034(.A(new_n222), .B1(new_n212), .B2(new_n235), .ZN(new_n236));
  AND2_X1   g035(.A1(new_n221), .A2(new_n219), .ZN(new_n237));
  AOI22_X1  g036(.A1(new_n226), .A2(new_n211), .B1(new_n237), .B2(new_n218), .ZN(new_n238));
  OAI21_X1  g037(.A(KEYINPUT17), .B1(new_n236), .B2(new_n238), .ZN(new_n239));
  XOR2_X1   g038(.A(G15gat), .B(G22gat), .Z(new_n240));
  INV_X1    g039(.A(G1gat), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n240), .A2(new_n241), .ZN(new_n242));
  XNOR2_X1  g041(.A(G15gat), .B(G22gat), .ZN(new_n243));
  INV_X1    g042(.A(KEYINPUT16), .ZN(new_n244));
  OAI21_X1  g043(.A(new_n243), .B1(new_n244), .B2(G1gat), .ZN(new_n245));
  INV_X1    g044(.A(G8gat), .ZN(new_n246));
  OR2_X1    g045(.A1(new_n246), .A2(KEYINPUT92), .ZN(new_n247));
  NAND3_X1  g046(.A1(new_n242), .A2(new_n245), .A3(new_n247), .ZN(new_n248));
  NAND3_X1  g047(.A1(new_n248), .A2(KEYINPUT92), .A3(new_n246), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n246), .A2(KEYINPUT92), .ZN(new_n250));
  NAND4_X1  g049(.A1(new_n242), .A2(new_n245), .A3(new_n250), .A4(new_n247), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n249), .A2(new_n251), .ZN(new_n252));
  NAND3_X1  g051(.A1(new_n230), .A2(new_n239), .A3(new_n252), .ZN(new_n253));
  INV_X1    g052(.A(KEYINPUT93), .ZN(new_n254));
  NAND2_X1  g053(.A1(new_n253), .A2(new_n254), .ZN(new_n255));
  NAND4_X1  g054(.A1(new_n230), .A2(new_n239), .A3(KEYINPUT93), .A4(new_n252), .ZN(new_n256));
  NAND2_X1  g055(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  NAND2_X1  g056(.A1(G229gat), .A2(G233gat), .ZN(new_n258));
  OAI21_X1  g057(.A(new_n223), .B1(new_n229), .B2(new_n222), .ZN(new_n259));
  OAI21_X1  g058(.A(new_n258), .B1(new_n259), .B2(new_n252), .ZN(new_n260));
  INV_X1    g059(.A(new_n260), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n257), .A2(new_n261), .ZN(new_n262));
  INV_X1    g061(.A(KEYINPUT94), .ZN(new_n263));
  INV_X1    g062(.A(KEYINPUT18), .ZN(new_n264));
  NAND3_X1  g063(.A1(new_n262), .A2(new_n263), .A3(new_n264), .ZN(new_n265));
  AOI21_X1  g064(.A(new_n260), .B1(new_n255), .B2(new_n256), .ZN(new_n266));
  OAI21_X1  g065(.A(KEYINPUT94), .B1(new_n266), .B2(KEYINPUT18), .ZN(new_n267));
  XOR2_X1   g066(.A(new_n258), .B(KEYINPUT13), .Z(new_n268));
  INV_X1    g067(.A(new_n268), .ZN(new_n269));
  INV_X1    g068(.A(new_n252), .ZN(new_n270));
  NOR2_X1   g069(.A1(new_n236), .A2(new_n238), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n259), .A2(new_n252), .ZN(new_n273));
  AOI21_X1  g072(.A(new_n269), .B1(new_n272), .B2(new_n273), .ZN(new_n274));
  AOI21_X1  g073(.A(new_n274), .B1(new_n266), .B2(KEYINPUT18), .ZN(new_n275));
  XNOR2_X1  g074(.A(G113gat), .B(G141gat), .ZN(new_n276));
  INV_X1    g075(.A(KEYINPUT11), .ZN(new_n277));
  XNOR2_X1  g076(.A(new_n276), .B(new_n277), .ZN(new_n278));
  XNOR2_X1  g077(.A(new_n278), .B(G169gat), .ZN(new_n279));
  INV_X1    g078(.A(G197gat), .ZN(new_n280));
  XNOR2_X1  g079(.A(new_n279), .B(new_n280), .ZN(new_n281));
  INV_X1    g080(.A(KEYINPUT12), .ZN(new_n282));
  XNOR2_X1  g081(.A(new_n281), .B(new_n282), .ZN(new_n283));
  NAND4_X1  g082(.A1(new_n265), .A2(new_n267), .A3(new_n275), .A4(new_n283), .ZN(new_n284));
  INV_X1    g083(.A(new_n283), .ZN(new_n285));
  NAND3_X1  g084(.A1(new_n257), .A2(KEYINPUT18), .A3(new_n261), .ZN(new_n286));
  INV_X1    g085(.A(new_n274), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  NOR2_X1   g087(.A1(new_n266), .A2(KEYINPUT18), .ZN(new_n289));
  OAI21_X1  g088(.A(new_n285), .B1(new_n288), .B2(new_n289), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n284), .A2(new_n290), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n291), .A2(KEYINPUT95), .ZN(new_n292));
  INV_X1    g091(.A(KEYINPUT95), .ZN(new_n293));
  NAND3_X1  g092(.A1(new_n284), .A2(new_n290), .A3(new_n293), .ZN(new_n294));
  NAND2_X1  g093(.A1(new_n292), .A2(new_n294), .ZN(new_n295));
  INV_X1    g094(.A(new_n295), .ZN(new_n296));
  INV_X1    g095(.A(G190gat), .ZN(new_n297));
  INV_X1    g096(.A(KEYINPUT67), .ZN(new_n298));
  INV_X1    g097(.A(G183gat), .ZN(new_n299));
  OAI21_X1  g098(.A(new_n298), .B1(new_n299), .B2(KEYINPUT27), .ZN(new_n300));
  XNOR2_X1  g099(.A(KEYINPUT27), .B(G183gat), .ZN(new_n301));
  OAI211_X1 g100(.A(new_n297), .B(new_n300), .C1(new_n301), .C2(new_n298), .ZN(new_n302));
  INV_X1    g101(.A(KEYINPUT68), .ZN(new_n303));
  OR2_X1    g102(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  AOI21_X1  g103(.A(KEYINPUT28), .B1(new_n302), .B2(new_n303), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  AND2_X1   g105(.A1(new_n297), .A2(KEYINPUT28), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n301), .A2(new_n307), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n306), .A2(new_n308), .ZN(new_n309));
  NOR2_X1   g108(.A1(G169gat), .A2(G176gat), .ZN(new_n310));
  INV_X1    g109(.A(KEYINPUT26), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  OAI21_X1  g111(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n313));
  NAND2_X1  g112(.A1(G169gat), .A2(G176gat), .ZN(new_n314));
  NAND3_X1  g113(.A1(new_n312), .A2(new_n313), .A3(new_n314), .ZN(new_n315));
  NAND2_X1  g114(.A1(G183gat), .A2(G190gat), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n315), .A2(new_n316), .ZN(new_n317));
  INV_X1    g116(.A(new_n317), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n309), .A2(new_n318), .ZN(new_n319));
  INV_X1    g118(.A(G113gat), .ZN(new_n320));
  INV_X1    g119(.A(G120gat), .ZN(new_n321));
  AOI21_X1  g120(.A(KEYINPUT1), .B1(new_n320), .B2(new_n321), .ZN(new_n322));
  OAI21_X1  g121(.A(new_n322), .B1(new_n320), .B2(new_n321), .ZN(new_n323));
  XNOR2_X1  g122(.A(G127gat), .B(G134gat), .ZN(new_n324));
  XNOR2_X1  g123(.A(new_n323), .B(new_n324), .ZN(new_n325));
  NOR2_X1   g124(.A1(G183gat), .A2(G190gat), .ZN(new_n326));
  INV_X1    g125(.A(KEYINPUT64), .ZN(new_n327));
  XNOR2_X1  g126(.A(new_n326), .B(new_n327), .ZN(new_n328));
  XNOR2_X1  g127(.A(new_n316), .B(KEYINPUT24), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n328), .A2(new_n329), .ZN(new_n330));
  INV_X1    g129(.A(KEYINPUT23), .ZN(new_n331));
  OAI21_X1  g130(.A(new_n331), .B1(G169gat), .B2(G176gat), .ZN(new_n332));
  XOR2_X1   g131(.A(KEYINPUT65), .B(G169gat), .Z(new_n333));
  INV_X1    g132(.A(G176gat), .ZN(new_n334));
  NAND3_X1  g133(.A1(new_n333), .A2(KEYINPUT23), .A3(new_n334), .ZN(new_n335));
  AOI21_X1  g134(.A(KEYINPUT25), .B1(G169gat), .B2(G176gat), .ZN(new_n336));
  NAND4_X1  g135(.A1(new_n330), .A2(new_n332), .A3(new_n335), .A4(new_n336), .ZN(new_n337));
  INV_X1    g136(.A(KEYINPUT25), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n310), .A2(KEYINPUT23), .ZN(new_n339));
  NAND3_X1  g138(.A1(new_n339), .A2(new_n314), .A3(new_n332), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n316), .A2(KEYINPUT66), .ZN(new_n341));
  OR2_X1    g140(.A1(new_n341), .A2(KEYINPUT24), .ZN(new_n342));
  AOI21_X1  g141(.A(new_n326), .B1(new_n341), .B2(KEYINPUT24), .ZN(new_n343));
  AOI21_X1  g142(.A(new_n340), .B1(new_n342), .B2(new_n343), .ZN(new_n344));
  OAI21_X1  g143(.A(new_n337), .B1(new_n338), .B2(new_n344), .ZN(new_n345));
  INV_X1    g144(.A(new_n345), .ZN(new_n346));
  NAND3_X1  g145(.A1(new_n319), .A2(new_n325), .A3(new_n346), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n347), .A2(KEYINPUT69), .ZN(new_n348));
  AOI21_X1  g147(.A(new_n317), .B1(new_n306), .B2(new_n308), .ZN(new_n349));
  NOR2_X1   g148(.A1(new_n349), .A2(new_n345), .ZN(new_n350));
  INV_X1    g149(.A(KEYINPUT69), .ZN(new_n351));
  NAND3_X1  g150(.A1(new_n350), .A2(new_n351), .A3(new_n325), .ZN(new_n352));
  NAND2_X1  g151(.A1(G227gat), .A2(G233gat), .ZN(new_n353));
  INV_X1    g152(.A(new_n325), .ZN(new_n354));
  OAI21_X1  g153(.A(new_n354), .B1(new_n349), .B2(new_n345), .ZN(new_n355));
  NAND4_X1  g154(.A1(new_n348), .A2(new_n352), .A3(new_n353), .A4(new_n355), .ZN(new_n356));
  INV_X1    g155(.A(KEYINPUT34), .ZN(new_n357));
  XNOR2_X1  g156(.A(new_n356), .B(new_n357), .ZN(new_n358));
  INV_X1    g157(.A(new_n358), .ZN(new_n359));
  INV_X1    g158(.A(KEYINPUT32), .ZN(new_n360));
  NAND3_X1  g159(.A1(new_n348), .A2(new_n352), .A3(new_n355), .ZN(new_n361));
  INV_X1    g160(.A(new_n353), .ZN(new_n362));
  AOI21_X1  g161(.A(new_n360), .B1(new_n361), .B2(new_n362), .ZN(new_n363));
  AOI21_X1  g162(.A(KEYINPUT33), .B1(new_n361), .B2(new_n362), .ZN(new_n364));
  XNOR2_X1  g163(.A(KEYINPUT70), .B(G71gat), .ZN(new_n365));
  XNOR2_X1  g164(.A(new_n365), .B(G99gat), .ZN(new_n366));
  XOR2_X1   g165(.A(G15gat), .B(G43gat), .Z(new_n367));
  XOR2_X1   g166(.A(new_n366), .B(new_n367), .Z(new_n368));
  INV_X1    g167(.A(new_n368), .ZN(new_n369));
  NOR3_X1   g168(.A1(new_n363), .A2(new_n364), .A3(new_n369), .ZN(new_n370));
  AOI221_X4 g169(.A(new_n360), .B1(KEYINPUT33), .B2(new_n368), .C1(new_n361), .C2(new_n362), .ZN(new_n371));
  OAI21_X1  g170(.A(new_n359), .B1(new_n370), .B2(new_n371), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n372), .A2(KEYINPUT71), .ZN(new_n373));
  AOI21_X1  g172(.A(new_n351), .B1(new_n350), .B2(new_n325), .ZN(new_n374));
  INV_X1    g173(.A(new_n355), .ZN(new_n375));
  NOR4_X1   g174(.A1(new_n349), .A2(KEYINPUT69), .A3(new_n345), .A4(new_n354), .ZN(new_n376));
  NOR3_X1   g175(.A1(new_n374), .A2(new_n375), .A3(new_n376), .ZN(new_n377));
  OAI21_X1  g176(.A(KEYINPUT32), .B1(new_n377), .B2(new_n353), .ZN(new_n378));
  INV_X1    g177(.A(KEYINPUT33), .ZN(new_n379));
  OAI21_X1  g178(.A(new_n379), .B1(new_n377), .B2(new_n353), .ZN(new_n380));
  NAND3_X1  g179(.A1(new_n378), .A2(new_n380), .A3(new_n368), .ZN(new_n381));
  OAI21_X1  g180(.A(new_n363), .B1(new_n364), .B2(new_n369), .ZN(new_n382));
  AOI21_X1  g181(.A(new_n358), .B1(new_n381), .B2(new_n382), .ZN(new_n383));
  INV_X1    g182(.A(KEYINPUT71), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n373), .A2(new_n385), .ZN(new_n386));
  XNOR2_X1  g185(.A(G64gat), .B(G92gat), .ZN(new_n387));
  XNOR2_X1  g186(.A(new_n387), .B(KEYINPUT78), .ZN(new_n388));
  XNOR2_X1  g187(.A(G8gat), .B(G36gat), .ZN(new_n389));
  XOR2_X1   g188(.A(new_n388), .B(new_n389), .Z(new_n390));
  OAI21_X1  g189(.A(KEYINPUT76), .B1(new_n349), .B2(new_n345), .ZN(new_n391));
  INV_X1    g190(.A(KEYINPUT76), .ZN(new_n392));
  AOI22_X1  g191(.A1(new_n304), .A2(new_n305), .B1(new_n301), .B2(new_n307), .ZN(new_n393));
  OAI211_X1 g192(.A(new_n346), .B(new_n392), .C1(new_n393), .C2(new_n317), .ZN(new_n394));
  NAND2_X1  g193(.A1(G226gat), .A2(G233gat), .ZN(new_n395));
  XOR2_X1   g194(.A(new_n395), .B(KEYINPUT75), .Z(new_n396));
  NAND3_X1  g195(.A1(new_n391), .A2(new_n394), .A3(new_n396), .ZN(new_n397));
  OAI21_X1  g196(.A(new_n395), .B1(new_n350), .B2(KEYINPUT29), .ZN(new_n398));
  XNOR2_X1  g197(.A(G211gat), .B(G218gat), .ZN(new_n399));
  INV_X1    g198(.A(KEYINPUT73), .ZN(new_n400));
  XNOR2_X1  g199(.A(new_n399), .B(new_n400), .ZN(new_n401));
  INV_X1    g200(.A(KEYINPUT74), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n401), .A2(new_n402), .ZN(new_n403));
  XNOR2_X1  g202(.A(new_n399), .B(KEYINPUT73), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n404), .A2(KEYINPUT74), .ZN(new_n405));
  XNOR2_X1  g204(.A(KEYINPUT72), .B(G218gat), .ZN(new_n406));
  INV_X1    g205(.A(G211gat), .ZN(new_n407));
  NOR2_X1   g206(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  OR2_X1    g207(.A1(new_n408), .A2(KEYINPUT22), .ZN(new_n409));
  XNOR2_X1  g208(.A(G197gat), .B(G204gat), .ZN(new_n410));
  NAND4_X1  g209(.A1(new_n403), .A2(new_n405), .A3(new_n409), .A4(new_n410), .ZN(new_n411));
  OAI21_X1  g210(.A(new_n410), .B1(new_n408), .B2(KEYINPUT22), .ZN(new_n412));
  NAND3_X1  g211(.A1(new_n412), .A2(new_n401), .A3(new_n402), .ZN(new_n413));
  AND2_X1   g212(.A1(new_n411), .A2(new_n413), .ZN(new_n414));
  NAND3_X1  g213(.A1(new_n397), .A2(new_n398), .A3(new_n414), .ZN(new_n415));
  NOR2_X1   g214(.A1(new_n350), .A2(new_n395), .ZN(new_n416));
  XNOR2_X1  g215(.A(KEYINPUT77), .B(KEYINPUT29), .ZN(new_n417));
  NAND3_X1  g216(.A1(new_n391), .A2(new_n394), .A3(new_n417), .ZN(new_n418));
  INV_X1    g217(.A(new_n396), .ZN(new_n419));
  AOI21_X1  g218(.A(new_n416), .B1(new_n418), .B2(new_n419), .ZN(new_n420));
  OAI211_X1 g219(.A(new_n390), .B(new_n415), .C1(new_n420), .C2(new_n414), .ZN(new_n421));
  INV_X1    g220(.A(new_n421), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n422), .A2(KEYINPUT30), .ZN(new_n423));
  INV_X1    g222(.A(KEYINPUT30), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n421), .A2(new_n424), .ZN(new_n425));
  OAI21_X1  g224(.A(new_n415), .B1(new_n420), .B2(new_n414), .ZN(new_n426));
  INV_X1    g225(.A(new_n390), .ZN(new_n427));
  AND3_X1   g226(.A1(new_n426), .A2(KEYINPUT79), .A3(new_n427), .ZN(new_n428));
  AOI21_X1  g227(.A(KEYINPUT79), .B1(new_n426), .B2(new_n427), .ZN(new_n429));
  OAI211_X1 g228(.A(new_n423), .B(new_n425), .C1(new_n428), .C2(new_n429), .ZN(new_n430));
  INV_X1    g229(.A(KEYINPUT85), .ZN(new_n431));
  INV_X1    g230(.A(KEYINPUT29), .ZN(new_n432));
  NAND3_X1  g231(.A1(new_n411), .A2(new_n432), .A3(new_n413), .ZN(new_n433));
  INV_X1    g232(.A(KEYINPUT3), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n433), .A2(new_n434), .ZN(new_n435));
  XOR2_X1   g234(.A(G141gat), .B(G148gat), .Z(new_n436));
  INV_X1    g235(.A(KEYINPUT2), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n436), .A2(new_n437), .ZN(new_n438));
  INV_X1    g237(.A(G155gat), .ZN(new_n439));
  INV_X1    g238(.A(G162gat), .ZN(new_n440));
  NAND3_X1  g239(.A1(new_n439), .A2(new_n440), .A3(KEYINPUT80), .ZN(new_n441));
  INV_X1    g240(.A(KEYINPUT80), .ZN(new_n442));
  OAI21_X1  g241(.A(new_n442), .B1(G155gat), .B2(G162gat), .ZN(new_n443));
  NAND2_X1  g242(.A1(G155gat), .A2(G162gat), .ZN(new_n444));
  AND2_X1   g243(.A1(new_n443), .A2(new_n444), .ZN(new_n445));
  NAND3_X1  g244(.A1(new_n438), .A2(new_n441), .A3(new_n445), .ZN(new_n446));
  NAND3_X1  g245(.A1(new_n437), .A2(new_n439), .A3(new_n440), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n447), .A2(new_n444), .ZN(new_n448));
  INV_X1    g247(.A(KEYINPUT81), .ZN(new_n449));
  NAND3_X1  g248(.A1(new_n436), .A2(new_n448), .A3(new_n449), .ZN(new_n450));
  INV_X1    g249(.A(new_n450), .ZN(new_n451));
  AOI21_X1  g250(.A(new_n449), .B1(new_n436), .B2(new_n448), .ZN(new_n452));
  OAI21_X1  g251(.A(new_n446), .B1(new_n451), .B2(new_n452), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n453), .A2(KEYINPUT82), .ZN(new_n454));
  INV_X1    g253(.A(KEYINPUT82), .ZN(new_n455));
  OAI211_X1 g254(.A(new_n455), .B(new_n446), .C1(new_n451), .C2(new_n452), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n454), .A2(new_n456), .ZN(new_n457));
  INV_X1    g256(.A(new_n457), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n435), .A2(new_n458), .ZN(new_n459));
  INV_X1    g258(.A(KEYINPUT84), .ZN(new_n460));
  NOR2_X1   g259(.A1(new_n453), .A2(KEYINPUT3), .ZN(new_n461));
  INV_X1    g260(.A(new_n417), .ZN(new_n462));
  NOR2_X1   g261(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  OAI21_X1  g262(.A(new_n460), .B1(new_n414), .B2(new_n463), .ZN(new_n464));
  INV_X1    g263(.A(G228gat), .ZN(new_n465));
  INV_X1    g264(.A(G233gat), .ZN(new_n466));
  NOR2_X1   g265(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n411), .A2(new_n413), .ZN(new_n468));
  OAI211_X1 g267(.A(new_n468), .B(KEYINPUT84), .C1(new_n461), .C2(new_n462), .ZN(new_n469));
  NAND4_X1  g268(.A1(new_n459), .A2(new_n464), .A3(new_n467), .A4(new_n469), .ZN(new_n470));
  NOR2_X1   g269(.A1(new_n414), .A2(new_n463), .ZN(new_n471));
  INV_X1    g270(.A(new_n453), .ZN(new_n472));
  NAND3_X1  g271(.A1(new_n411), .A2(new_n417), .A3(new_n413), .ZN(new_n473));
  AOI21_X1  g272(.A(new_n472), .B1(new_n473), .B2(new_n434), .ZN(new_n474));
  OAI22_X1  g273(.A1(new_n471), .A2(new_n474), .B1(new_n465), .B2(new_n466), .ZN(new_n475));
  INV_X1    g274(.A(G22gat), .ZN(new_n476));
  NAND3_X1  g275(.A1(new_n470), .A2(new_n475), .A3(new_n476), .ZN(new_n477));
  INV_X1    g276(.A(new_n477), .ZN(new_n478));
  AOI21_X1  g277(.A(new_n476), .B1(new_n470), .B2(new_n475), .ZN(new_n479));
  OAI21_X1  g278(.A(new_n431), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n470), .A2(new_n475), .ZN(new_n481));
  NAND2_X1  g280(.A1(new_n481), .A2(G22gat), .ZN(new_n482));
  NAND3_X1  g281(.A1(new_n482), .A2(KEYINPUT85), .A3(new_n477), .ZN(new_n483));
  XNOR2_X1  g282(.A(G78gat), .B(G106gat), .ZN(new_n484));
  XNOR2_X1  g283(.A(KEYINPUT31), .B(G50gat), .ZN(new_n485));
  XOR2_X1   g284(.A(new_n484), .B(new_n485), .Z(new_n486));
  INV_X1    g285(.A(new_n486), .ZN(new_n487));
  NAND3_X1  g286(.A1(new_n480), .A2(new_n483), .A3(new_n487), .ZN(new_n488));
  NAND3_X1  g287(.A1(new_n381), .A2(new_n358), .A3(new_n382), .ZN(new_n489));
  NAND4_X1  g288(.A1(new_n482), .A2(KEYINPUT85), .A3(new_n477), .A4(new_n486), .ZN(new_n490));
  NAND3_X1  g289(.A1(new_n488), .A2(new_n489), .A3(new_n490), .ZN(new_n491));
  NOR3_X1   g290(.A1(new_n386), .A2(new_n430), .A3(new_n491), .ZN(new_n492));
  INV_X1    g291(.A(KEYINPUT35), .ZN(new_n493));
  INV_X1    g292(.A(KEYINPUT5), .ZN(new_n494));
  NOR2_X1   g293(.A1(new_n354), .A2(new_n453), .ZN(new_n495));
  INV_X1    g294(.A(new_n495), .ZN(new_n496));
  OAI21_X1  g295(.A(new_n496), .B1(new_n457), .B2(new_n325), .ZN(new_n497));
  NAND2_X1  g296(.A1(G225gat), .A2(G233gat), .ZN(new_n498));
  INV_X1    g297(.A(new_n498), .ZN(new_n499));
  AOI21_X1  g298(.A(new_n494), .B1(new_n497), .B2(new_n499), .ZN(new_n500));
  NOR2_X1   g299(.A1(new_n495), .A2(KEYINPUT4), .ZN(new_n501));
  INV_X1    g300(.A(KEYINPUT4), .ZN(new_n502));
  NOR3_X1   g301(.A1(new_n354), .A2(new_n453), .A3(new_n502), .ZN(new_n503));
  NOR2_X1   g302(.A1(new_n501), .A2(new_n503), .ZN(new_n504));
  INV_X1    g303(.A(new_n461), .ZN(new_n505));
  OAI211_X1 g304(.A(new_n354), .B(new_n505), .C1(new_n457), .C2(new_n434), .ZN(new_n506));
  NAND2_X1  g305(.A1(new_n504), .A2(new_n506), .ZN(new_n507));
  NOR2_X1   g306(.A1(new_n495), .A2(new_n498), .ZN(new_n508));
  OAI21_X1  g307(.A(new_n500), .B1(new_n507), .B2(new_n508), .ZN(new_n509));
  NAND4_X1  g308(.A1(new_n504), .A2(new_n506), .A3(new_n494), .A4(new_n498), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  XNOR2_X1  g310(.A(G1gat), .B(G29gat), .ZN(new_n512));
  XNOR2_X1  g311(.A(new_n512), .B(KEYINPUT0), .ZN(new_n513));
  XNOR2_X1  g312(.A(new_n513), .B(G57gat), .ZN(new_n514));
  INV_X1    g313(.A(G85gat), .ZN(new_n515));
  XNOR2_X1  g314(.A(new_n514), .B(new_n515), .ZN(new_n516));
  INV_X1    g315(.A(new_n516), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n511), .A2(new_n517), .ZN(new_n518));
  INV_X1    g317(.A(KEYINPUT6), .ZN(new_n519));
  NOR2_X1   g318(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  INV_X1    g319(.A(new_n520), .ZN(new_n521));
  NAND3_X1  g320(.A1(new_n509), .A2(new_n516), .A3(new_n510), .ZN(new_n522));
  INV_X1    g321(.A(KEYINPUT83), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  NAND4_X1  g323(.A1(new_n509), .A2(KEYINPUT83), .A3(new_n516), .A4(new_n510), .ZN(new_n525));
  NAND4_X1  g324(.A1(new_n524), .A2(new_n518), .A3(new_n519), .A4(new_n525), .ZN(new_n526));
  AOI21_X1  g325(.A(new_n493), .B1(new_n521), .B2(new_n526), .ZN(new_n527));
  AND3_X1   g326(.A1(new_n524), .A2(new_n519), .A3(new_n525), .ZN(new_n528));
  NAND3_X1  g327(.A1(new_n509), .A2(KEYINPUT87), .A3(new_n510), .ZN(new_n529));
  INV_X1    g328(.A(new_n529), .ZN(new_n530));
  AOI21_X1  g329(.A(KEYINPUT87), .B1(new_n509), .B2(new_n510), .ZN(new_n531));
  OAI21_X1  g330(.A(new_n517), .B1(new_n530), .B2(new_n531), .ZN(new_n532));
  AOI21_X1  g331(.A(new_n520), .B1(new_n528), .B2(new_n532), .ZN(new_n533));
  INV_X1    g332(.A(new_n533), .ZN(new_n534));
  AND3_X1   g333(.A1(new_n488), .A2(new_n490), .A3(new_n489), .ZN(new_n535));
  INV_X1    g334(.A(new_n430), .ZN(new_n536));
  NAND4_X1  g335(.A1(new_n534), .A2(new_n535), .A3(new_n536), .A4(new_n372), .ZN(new_n537));
  AOI22_X1  g336(.A1(new_n492), .A2(new_n527), .B1(new_n537), .B2(new_n493), .ZN(new_n538));
  AND2_X1   g337(.A1(new_n426), .A2(KEYINPUT37), .ZN(new_n539));
  INV_X1    g338(.A(KEYINPUT37), .ZN(new_n540));
  OAI211_X1 g339(.A(new_n540), .B(new_n415), .C1(new_n420), .C2(new_n414), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n541), .A2(new_n427), .ZN(new_n542));
  OAI21_X1  g341(.A(KEYINPUT38), .B1(new_n539), .B2(new_n542), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n543), .A2(KEYINPUT88), .ZN(new_n544));
  INV_X1    g343(.A(KEYINPUT88), .ZN(new_n545));
  OAI211_X1 g344(.A(new_n545), .B(KEYINPUT38), .C1(new_n539), .C2(new_n542), .ZN(new_n546));
  INV_X1    g345(.A(new_n542), .ZN(new_n547));
  OR2_X1    g346(.A1(new_n420), .A2(new_n468), .ZN(new_n548));
  NAND3_X1  g347(.A1(new_n397), .A2(new_n398), .A3(new_n468), .ZN(new_n549));
  AND2_X1   g348(.A1(new_n549), .A2(KEYINPUT37), .ZN(new_n550));
  AOI21_X1  g349(.A(KEYINPUT38), .B1(new_n548), .B2(new_n550), .ZN(new_n551));
  AOI21_X1  g350(.A(new_n422), .B1(new_n547), .B2(new_n551), .ZN(new_n552));
  NAND4_X1  g351(.A1(new_n533), .A2(new_n544), .A3(new_n546), .A4(new_n552), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n488), .A2(new_n490), .ZN(new_n554));
  INV_X1    g353(.A(KEYINPUT39), .ZN(new_n555));
  NAND3_X1  g354(.A1(new_n507), .A2(new_n555), .A3(new_n499), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n507), .A2(new_n499), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n557), .A2(KEYINPUT39), .ZN(new_n558));
  OAI211_X1 g357(.A(new_n496), .B(new_n498), .C1(new_n457), .C2(new_n325), .ZN(new_n559));
  XNOR2_X1  g358(.A(new_n559), .B(KEYINPUT86), .ZN(new_n560));
  OAI211_X1 g359(.A(new_n516), .B(new_n556), .C1(new_n558), .C2(new_n560), .ZN(new_n561));
  INV_X1    g360(.A(KEYINPUT40), .ZN(new_n562));
  NAND2_X1  g361(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  AND2_X1   g362(.A1(new_n556), .A2(new_n516), .ZN(new_n564));
  OAI211_X1 g363(.A(new_n564), .B(KEYINPUT40), .C1(new_n558), .C2(new_n560), .ZN(new_n565));
  AND3_X1   g364(.A1(new_n532), .A2(new_n563), .A3(new_n565), .ZN(new_n566));
  AOI21_X1  g365(.A(new_n554), .B1(new_n566), .B2(new_n430), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n553), .A2(new_n567), .ZN(new_n568));
  NAND4_X1  g367(.A1(new_n373), .A2(new_n385), .A3(KEYINPUT36), .A4(new_n489), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n372), .A2(new_n489), .ZN(new_n570));
  INV_X1    g369(.A(KEYINPUT36), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  NAND2_X1  g371(.A1(new_n569), .A2(new_n572), .ZN(new_n573));
  NAND2_X1  g372(.A1(new_n521), .A2(new_n526), .ZN(new_n574));
  INV_X1    g373(.A(new_n574), .ZN(new_n575));
  OAI21_X1  g374(.A(new_n554), .B1(new_n575), .B2(new_n430), .ZN(new_n576));
  NAND3_X1  g375(.A1(new_n568), .A2(new_n573), .A3(new_n576), .ZN(new_n577));
  AOI21_X1  g376(.A(new_n296), .B1(new_n538), .B2(new_n577), .ZN(new_n578));
  XNOR2_X1  g377(.A(KEYINPUT98), .B(G183gat), .ZN(new_n579));
  INV_X1    g378(.A(new_n579), .ZN(new_n580));
  XNOR2_X1  g379(.A(G71gat), .B(G78gat), .ZN(new_n581));
  INV_X1    g380(.A(new_n581), .ZN(new_n582));
  AOI21_X1  g381(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n583));
  AND2_X1   g382(.A1(G57gat), .A2(G64gat), .ZN(new_n584));
  NOR2_X1   g383(.A1(G57gat), .A2(G64gat), .ZN(new_n585));
  NOR3_X1   g384(.A1(new_n583), .A2(new_n584), .A3(new_n585), .ZN(new_n586));
  OAI21_X1  g385(.A(KEYINPUT96), .B1(G71gat), .B2(G78gat), .ZN(new_n587));
  INV_X1    g386(.A(new_n587), .ZN(new_n588));
  OAI21_X1  g387(.A(new_n582), .B1(new_n586), .B2(new_n588), .ZN(new_n589));
  NAND2_X1  g388(.A1(G71gat), .A2(G78gat), .ZN(new_n590));
  INV_X1    g389(.A(KEYINPUT9), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  OR2_X1    g391(.A1(G57gat), .A2(G64gat), .ZN(new_n593));
  NAND2_X1  g392(.A1(G57gat), .A2(G64gat), .ZN(new_n594));
  NAND3_X1  g393(.A1(new_n592), .A2(new_n593), .A3(new_n594), .ZN(new_n595));
  NAND3_X1  g394(.A1(new_n595), .A2(new_n581), .A3(new_n587), .ZN(new_n596));
  NAND2_X1  g395(.A1(new_n589), .A2(new_n596), .ZN(new_n597));
  NOR2_X1   g396(.A1(new_n597), .A2(KEYINPUT21), .ZN(new_n598));
  XNOR2_X1  g397(.A(G127gat), .B(G155gat), .ZN(new_n599));
  INV_X1    g398(.A(new_n599), .ZN(new_n600));
  NOR2_X1   g399(.A1(new_n598), .A2(new_n600), .ZN(new_n601));
  INV_X1    g400(.A(new_n601), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n598), .A2(new_n600), .ZN(new_n603));
  AOI21_X1  g402(.A(new_n407), .B1(new_n602), .B2(new_n603), .ZN(new_n604));
  INV_X1    g403(.A(new_n603), .ZN(new_n605));
  NOR3_X1   g404(.A1(new_n605), .A2(G211gat), .A3(new_n601), .ZN(new_n606));
  NOR2_X1   g405(.A1(new_n604), .A2(new_n606), .ZN(new_n607));
  NAND2_X1  g406(.A1(G231gat), .A2(G233gat), .ZN(new_n608));
  XNOR2_X1  g407(.A(new_n608), .B(KEYINPUT97), .ZN(new_n609));
  XNOR2_X1  g408(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n610));
  XOR2_X1   g409(.A(new_n609), .B(new_n610), .Z(new_n611));
  NAND2_X1  g410(.A1(new_n607), .A2(new_n611), .ZN(new_n612));
  AOI21_X1  g411(.A(new_n270), .B1(KEYINPUT21), .B2(new_n597), .ZN(new_n613));
  INV_X1    g412(.A(new_n613), .ZN(new_n614));
  INV_X1    g413(.A(new_n611), .ZN(new_n615));
  OAI21_X1  g414(.A(new_n615), .B1(new_n604), .B2(new_n606), .ZN(new_n616));
  AND3_X1   g415(.A1(new_n612), .A2(new_n614), .A3(new_n616), .ZN(new_n617));
  AOI21_X1  g416(.A(new_n614), .B1(new_n612), .B2(new_n616), .ZN(new_n618));
  OAI21_X1  g417(.A(new_n580), .B1(new_n617), .B2(new_n618), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n612), .A2(new_n616), .ZN(new_n620));
  NAND2_X1  g419(.A1(new_n620), .A2(new_n613), .ZN(new_n621));
  NAND3_X1  g420(.A1(new_n612), .A2(new_n614), .A3(new_n616), .ZN(new_n622));
  NAND3_X1  g421(.A1(new_n621), .A2(new_n579), .A3(new_n622), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n619), .A2(new_n623), .ZN(new_n624));
  INV_X1    g423(.A(KEYINPUT99), .ZN(new_n625));
  NAND2_X1  g424(.A1(G99gat), .A2(G106gat), .ZN(new_n626));
  NAND2_X1  g425(.A1(new_n626), .A2(KEYINPUT8), .ZN(new_n627));
  NAND2_X1  g426(.A1(G85gat), .A2(G92gat), .ZN(new_n628));
  INV_X1    g427(.A(KEYINPUT7), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  INV_X1    g429(.A(G92gat), .ZN(new_n631));
  NAND2_X1  g430(.A1(new_n515), .A2(new_n631), .ZN(new_n632));
  NAND3_X1  g431(.A1(KEYINPUT7), .A2(G85gat), .A3(G92gat), .ZN(new_n633));
  NAND4_X1  g432(.A1(new_n627), .A2(new_n630), .A3(new_n632), .A4(new_n633), .ZN(new_n634));
  XNOR2_X1  g433(.A(G99gat), .B(G106gat), .ZN(new_n635));
  INV_X1    g434(.A(new_n635), .ZN(new_n636));
  NOR2_X1   g435(.A1(new_n634), .A2(new_n636), .ZN(new_n637));
  AND3_X1   g436(.A1(KEYINPUT7), .A2(G85gat), .A3(G92gat), .ZN(new_n638));
  AOI21_X1  g437(.A(KEYINPUT7), .B1(G85gat), .B2(G92gat), .ZN(new_n639));
  NOR2_X1   g438(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  AOI22_X1  g439(.A1(KEYINPUT8), .A2(new_n626), .B1(new_n515), .B2(new_n631), .ZN(new_n641));
  AOI21_X1  g440(.A(new_n635), .B1(new_n640), .B2(new_n641), .ZN(new_n642));
  OAI21_X1  g441(.A(new_n625), .B1(new_n637), .B2(new_n642), .ZN(new_n643));
  NAND2_X1  g442(.A1(new_n634), .A2(new_n636), .ZN(new_n644));
  NAND3_X1  g443(.A1(new_n640), .A2(new_n635), .A3(new_n641), .ZN(new_n645));
  NAND3_X1  g444(.A1(new_n644), .A2(KEYINPUT99), .A3(new_n645), .ZN(new_n646));
  NAND2_X1  g445(.A1(new_n643), .A2(new_n646), .ZN(new_n647));
  NOR2_X1   g446(.A1(new_n259), .A2(new_n647), .ZN(new_n648));
  AND2_X1   g447(.A1(G232gat), .A2(G233gat), .ZN(new_n649));
  AOI21_X1  g448(.A(new_n648), .B1(KEYINPUT41), .B2(new_n649), .ZN(new_n650));
  XOR2_X1   g449(.A(G190gat), .B(G218gat), .Z(new_n651));
  XNOR2_X1  g450(.A(new_n651), .B(KEYINPUT100), .ZN(new_n652));
  NAND3_X1  g451(.A1(new_n230), .A2(new_n239), .A3(new_n647), .ZN(new_n653));
  AND3_X1   g452(.A1(new_n650), .A2(new_n652), .A3(new_n653), .ZN(new_n654));
  AOI21_X1  g453(.A(new_n652), .B1(new_n650), .B2(new_n653), .ZN(new_n655));
  XOR2_X1   g454(.A(G134gat), .B(G162gat), .Z(new_n656));
  NOR2_X1   g455(.A1(new_n649), .A2(KEYINPUT41), .ZN(new_n657));
  XNOR2_X1  g456(.A(new_n656), .B(new_n657), .ZN(new_n658));
  OR3_X1    g457(.A1(new_n654), .A2(new_n655), .A3(new_n658), .ZN(new_n659));
  OAI21_X1  g458(.A(new_n658), .B1(new_n654), .B2(new_n655), .ZN(new_n660));
  NAND2_X1  g459(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  OAI21_X1  g460(.A(KEYINPUT101), .B1(new_n624), .B2(new_n661), .ZN(new_n662));
  INV_X1    g461(.A(new_n661), .ZN(new_n663));
  INV_X1    g462(.A(KEYINPUT101), .ZN(new_n664));
  NAND4_X1  g463(.A1(new_n663), .A2(new_n619), .A3(new_n623), .A4(new_n664), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n662), .A2(new_n665), .ZN(new_n666));
  NAND2_X1  g465(.A1(G230gat), .A2(G233gat), .ZN(new_n667));
  XNOR2_X1  g466(.A(new_n667), .B(KEYINPUT104), .ZN(new_n668));
  INV_X1    g467(.A(KEYINPUT10), .ZN(new_n669));
  AOI21_X1  g468(.A(new_n669), .B1(new_n589), .B2(new_n596), .ZN(new_n670));
  NAND3_X1  g469(.A1(new_n670), .A2(new_n643), .A3(new_n646), .ZN(new_n671));
  INV_X1    g470(.A(KEYINPUT103), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  NAND4_X1  g472(.A1(new_n670), .A2(new_n643), .A3(KEYINPUT103), .A4(new_n646), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  INV_X1    g474(.A(KEYINPUT102), .ZN(new_n676));
  OAI21_X1  g475(.A(new_n676), .B1(new_n637), .B2(new_n642), .ZN(new_n677));
  AND3_X1   g476(.A1(new_n595), .A2(new_n581), .A3(new_n587), .ZN(new_n678));
  AOI21_X1  g477(.A(new_n581), .B1(new_n595), .B2(new_n587), .ZN(new_n679));
  NOR2_X1   g478(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  NAND3_X1  g479(.A1(new_n644), .A2(KEYINPUT102), .A3(new_n645), .ZN(new_n681));
  NAND3_X1  g480(.A1(new_n677), .A2(new_n680), .A3(new_n681), .ZN(new_n682));
  NAND2_X1  g481(.A1(new_n644), .A2(new_n645), .ZN(new_n683));
  NAND3_X1  g482(.A1(new_n597), .A2(new_n676), .A3(new_n683), .ZN(new_n684));
  NAND2_X1  g483(.A1(new_n682), .A2(new_n684), .ZN(new_n685));
  NAND2_X1  g484(.A1(new_n685), .A2(new_n669), .ZN(new_n686));
  AOI21_X1  g485(.A(new_n668), .B1(new_n675), .B2(new_n686), .ZN(new_n687));
  INV_X1    g486(.A(new_n687), .ZN(new_n688));
  NAND3_X1  g487(.A1(new_n682), .A2(new_n668), .A3(new_n684), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  XNOR2_X1  g489(.A(G120gat), .B(G148gat), .ZN(new_n691));
  XNOR2_X1  g490(.A(new_n691), .B(G176gat), .ZN(new_n692));
  XOR2_X1   g491(.A(new_n692), .B(G204gat), .Z(new_n693));
  INV_X1    g492(.A(new_n693), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n690), .A2(new_n694), .ZN(new_n695));
  NAND3_X1  g494(.A1(new_n688), .A2(new_n689), .A3(new_n693), .ZN(new_n696));
  NAND2_X1  g495(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  NOR2_X1   g496(.A1(new_n666), .A2(new_n697), .ZN(new_n698));
  NAND2_X1  g497(.A1(new_n578), .A2(new_n698), .ZN(new_n699));
  NOR2_X1   g498(.A1(new_n699), .A2(new_n574), .ZN(new_n700));
  XNOR2_X1  g499(.A(KEYINPUT105), .B(G1gat), .ZN(new_n701));
  XNOR2_X1  g500(.A(new_n700), .B(new_n701), .ZN(G1324gat));
  INV_X1    g501(.A(KEYINPUT42), .ZN(new_n703));
  INV_X1    g502(.A(new_n699), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n704), .A2(new_n430), .ZN(new_n705));
  XOR2_X1   g504(.A(KEYINPUT16), .B(G8gat), .Z(new_n706));
  INV_X1    g505(.A(new_n706), .ZN(new_n707));
  OAI21_X1  g506(.A(new_n703), .B1(new_n705), .B2(new_n707), .ZN(new_n708));
  NAND4_X1  g507(.A1(new_n704), .A2(KEYINPUT42), .A3(new_n430), .A4(new_n706), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n705), .A2(G8gat), .ZN(new_n710));
  NAND3_X1  g509(.A1(new_n708), .A2(new_n709), .A3(new_n710), .ZN(G1325gat));
  NAND2_X1  g510(.A1(new_n573), .A2(KEYINPUT106), .ZN(new_n712));
  INV_X1    g511(.A(KEYINPUT106), .ZN(new_n713));
  NAND3_X1  g512(.A1(new_n569), .A2(new_n713), .A3(new_n572), .ZN(new_n714));
  AND2_X1   g513(.A1(new_n712), .A2(new_n714), .ZN(new_n715));
  INV_X1    g514(.A(new_n715), .ZN(new_n716));
  OAI21_X1  g515(.A(G15gat), .B1(new_n699), .B2(new_n716), .ZN(new_n717));
  OR2_X1    g516(.A1(new_n570), .A2(G15gat), .ZN(new_n718));
  OAI21_X1  g517(.A(new_n717), .B1(new_n699), .B2(new_n718), .ZN(G1326gat));
  NAND2_X1  g518(.A1(new_n704), .A2(new_n554), .ZN(new_n720));
  XNOR2_X1  g519(.A(KEYINPUT43), .B(G22gat), .ZN(new_n721));
  XNOR2_X1  g520(.A(new_n720), .B(new_n721), .ZN(G1327gat));
  INV_X1    g521(.A(new_n624), .ZN(new_n723));
  NOR2_X1   g522(.A1(new_n723), .A2(new_n697), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n724), .A2(new_n661), .ZN(new_n725));
  INV_X1    g524(.A(new_n725), .ZN(new_n726));
  NAND4_X1  g525(.A1(new_n578), .A2(new_n213), .A3(new_n575), .A4(new_n726), .ZN(new_n727));
  XNOR2_X1  g526(.A(new_n727), .B(KEYINPUT45), .ZN(new_n728));
  NAND2_X1  g527(.A1(new_n724), .A2(new_n291), .ZN(new_n729));
  INV_X1    g528(.A(new_n729), .ZN(new_n730));
  INV_X1    g529(.A(KEYINPUT44), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n538), .A2(new_n577), .ZN(new_n732));
  AOI21_X1  g531(.A(new_n731), .B1(new_n732), .B2(new_n661), .ZN(new_n733));
  AOI211_X1 g532(.A(KEYINPUT44), .B(new_n663), .C1(new_n538), .C2(new_n577), .ZN(new_n734));
  OAI211_X1 g533(.A(new_n575), .B(new_n730), .C1(new_n733), .C2(new_n734), .ZN(new_n735));
  INV_X1    g534(.A(new_n735), .ZN(new_n736));
  OAI21_X1  g535(.A(G29gat), .B1(new_n736), .B2(KEYINPUT107), .ZN(new_n737));
  INV_X1    g536(.A(KEYINPUT107), .ZN(new_n738));
  NOR2_X1   g537(.A1(new_n735), .A2(new_n738), .ZN(new_n739));
  OAI21_X1  g538(.A(new_n728), .B1(new_n737), .B2(new_n739), .ZN(G1328gat));
  NAND4_X1  g539(.A1(new_n578), .A2(new_n214), .A3(new_n430), .A4(new_n726), .ZN(new_n741));
  XOR2_X1   g540(.A(new_n741), .B(KEYINPUT46), .Z(new_n742));
  OAI211_X1 g541(.A(new_n430), .B(new_n730), .C1(new_n733), .C2(new_n734), .ZN(new_n743));
  INV_X1    g542(.A(new_n743), .ZN(new_n744));
  OAI21_X1  g543(.A(G36gat), .B1(new_n744), .B2(KEYINPUT108), .ZN(new_n745));
  INV_X1    g544(.A(KEYINPUT108), .ZN(new_n746));
  NOR2_X1   g545(.A1(new_n743), .A2(new_n746), .ZN(new_n747));
  OAI21_X1  g546(.A(new_n742), .B1(new_n745), .B2(new_n747), .ZN(G1329gat));
  INV_X1    g547(.A(new_n570), .ZN(new_n749));
  AND4_X1   g548(.A1(new_n203), .A2(new_n578), .A3(new_n749), .A4(new_n726), .ZN(new_n750));
  OAI211_X1 g549(.A(new_n715), .B(new_n730), .C1(new_n733), .C2(new_n734), .ZN(new_n751));
  AOI21_X1  g550(.A(new_n750), .B1(new_n751), .B2(G43gat), .ZN(new_n752));
  AND3_X1   g551(.A1(new_n568), .A2(new_n573), .A3(new_n576), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n537), .A2(new_n493), .ZN(new_n754));
  XNOR2_X1  g553(.A(new_n383), .B(KEYINPUT71), .ZN(new_n755));
  NAND4_X1  g554(.A1(new_n755), .A2(new_n536), .A3(new_n535), .A4(new_n527), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n754), .A2(new_n756), .ZN(new_n757));
  OAI21_X1  g556(.A(new_n661), .B1(new_n753), .B2(new_n757), .ZN(new_n758));
  NAND2_X1  g557(.A1(new_n758), .A2(KEYINPUT44), .ZN(new_n759));
  NAND3_X1  g558(.A1(new_n732), .A2(new_n731), .A3(new_n661), .ZN(new_n760));
  AOI21_X1  g559(.A(new_n729), .B1(new_n759), .B2(new_n760), .ZN(new_n761));
  INV_X1    g560(.A(new_n573), .ZN(new_n762));
  AOI21_X1  g561(.A(new_n203), .B1(new_n761), .B2(new_n762), .ZN(new_n763));
  INV_X1    g562(.A(KEYINPUT47), .ZN(new_n764));
  OR2_X1    g563(.A1(new_n750), .A2(new_n764), .ZN(new_n765));
  OAI22_X1  g564(.A1(new_n752), .A2(KEYINPUT47), .B1(new_n763), .B2(new_n765), .ZN(G1330gat));
  INV_X1    g565(.A(KEYINPUT48), .ZN(new_n767));
  AOI21_X1  g566(.A(new_n227), .B1(new_n761), .B2(new_n554), .ZN(new_n768));
  NAND4_X1  g567(.A1(new_n578), .A2(new_n554), .A3(new_n227), .A4(new_n726), .ZN(new_n769));
  INV_X1    g568(.A(new_n769), .ZN(new_n770));
  OAI21_X1  g569(.A(new_n767), .B1(new_n768), .B2(new_n770), .ZN(new_n771));
  OAI211_X1 g570(.A(new_n554), .B(new_n730), .C1(new_n733), .C2(new_n734), .ZN(new_n772));
  INV_X1    g571(.A(new_n772), .ZN(new_n773));
  OAI211_X1 g572(.A(KEYINPUT48), .B(new_n769), .C1(new_n773), .C2(new_n227), .ZN(new_n774));
  NAND2_X1  g573(.A1(new_n771), .A2(new_n774), .ZN(G1331gat));
  INV_X1    g574(.A(new_n697), .ZN(new_n776));
  NOR3_X1   g575(.A1(new_n666), .A2(new_n291), .A3(new_n776), .ZN(new_n777));
  NAND2_X1  g576(.A1(new_n732), .A2(new_n777), .ZN(new_n778));
  NOR2_X1   g577(.A1(new_n778), .A2(new_n574), .ZN(new_n779));
  XNOR2_X1  g578(.A(KEYINPUT109), .B(G57gat), .ZN(new_n780));
  XNOR2_X1  g579(.A(new_n779), .B(new_n780), .ZN(G1332gat));
  NOR2_X1   g580(.A1(new_n778), .A2(new_n536), .ZN(new_n782));
  NOR2_X1   g581(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n783));
  AND2_X1   g582(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n784));
  OAI21_X1  g583(.A(new_n782), .B1(new_n783), .B2(new_n784), .ZN(new_n785));
  OAI21_X1  g584(.A(new_n785), .B1(new_n782), .B2(new_n783), .ZN(G1333gat));
  OAI21_X1  g585(.A(G71gat), .B1(new_n778), .B2(new_n716), .ZN(new_n787));
  OR2_X1    g586(.A1(new_n570), .A2(G71gat), .ZN(new_n788));
  OAI21_X1  g587(.A(new_n787), .B1(new_n778), .B2(new_n788), .ZN(new_n789));
  XOR2_X1   g588(.A(new_n789), .B(KEYINPUT50), .Z(G1334gat));
  INV_X1    g589(.A(new_n554), .ZN(new_n791));
  NOR2_X1   g590(.A1(new_n778), .A2(new_n791), .ZN(new_n792));
  XOR2_X1   g591(.A(KEYINPUT110), .B(G78gat), .Z(new_n793));
  XNOR2_X1  g592(.A(new_n792), .B(new_n793), .ZN(G1335gat));
  INV_X1    g593(.A(KEYINPUT111), .ZN(new_n795));
  NOR2_X1   g594(.A1(new_n723), .A2(new_n291), .ZN(new_n796));
  INV_X1    g595(.A(new_n796), .ZN(new_n797));
  NOR2_X1   g596(.A1(new_n797), .A2(new_n776), .ZN(new_n798));
  INV_X1    g597(.A(new_n798), .ZN(new_n799));
  AOI21_X1  g598(.A(new_n799), .B1(new_n759), .B2(new_n760), .ZN(new_n800));
  AOI21_X1  g599(.A(new_n515), .B1(new_n800), .B2(new_n575), .ZN(new_n801));
  OAI21_X1  g600(.A(KEYINPUT51), .B1(new_n758), .B2(new_n797), .ZN(new_n802));
  INV_X1    g601(.A(KEYINPUT51), .ZN(new_n803));
  NAND4_X1  g602(.A1(new_n732), .A2(new_n803), .A3(new_n661), .A4(new_n796), .ZN(new_n804));
  NOR2_X1   g603(.A1(new_n574), .A2(G85gat), .ZN(new_n805));
  AND4_X1   g604(.A1(new_n697), .A2(new_n802), .A3(new_n804), .A4(new_n805), .ZN(new_n806));
  OAI21_X1  g605(.A(new_n795), .B1(new_n801), .B2(new_n806), .ZN(new_n807));
  OAI211_X1 g606(.A(new_n575), .B(new_n798), .C1(new_n733), .C2(new_n734), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n808), .A2(G85gat), .ZN(new_n809));
  NAND3_X1  g608(.A1(new_n802), .A2(new_n697), .A3(new_n804), .ZN(new_n810));
  INV_X1    g609(.A(new_n805), .ZN(new_n811));
  OAI211_X1 g610(.A(new_n809), .B(KEYINPUT111), .C1(new_n810), .C2(new_n811), .ZN(new_n812));
  NAND2_X1  g611(.A1(new_n807), .A2(new_n812), .ZN(G1336gat));
  AOI21_X1  g612(.A(new_n631), .B1(new_n800), .B2(new_n430), .ZN(new_n814));
  NOR2_X1   g613(.A1(new_n536), .A2(G92gat), .ZN(new_n815));
  AND4_X1   g614(.A1(new_n697), .A2(new_n802), .A3(new_n804), .A4(new_n815), .ZN(new_n816));
  OAI21_X1  g615(.A(KEYINPUT52), .B1(new_n814), .B2(new_n816), .ZN(new_n817));
  OAI211_X1 g616(.A(new_n430), .B(new_n798), .C1(new_n733), .C2(new_n734), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n818), .A2(G92gat), .ZN(new_n819));
  INV_X1    g618(.A(KEYINPUT52), .ZN(new_n820));
  INV_X1    g619(.A(new_n815), .ZN(new_n821));
  OAI211_X1 g620(.A(new_n819), .B(new_n820), .C1(new_n810), .C2(new_n821), .ZN(new_n822));
  NAND2_X1  g621(.A1(new_n817), .A2(new_n822), .ZN(G1337gat));
  NAND2_X1  g622(.A1(new_n800), .A2(new_n715), .ZN(new_n824));
  INV_X1    g623(.A(new_n824), .ZN(new_n825));
  XNOR2_X1  g624(.A(KEYINPUT112), .B(G99gat), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n749), .A2(new_n826), .ZN(new_n827));
  OAI22_X1  g626(.A1(new_n825), .A2(new_n826), .B1(new_n810), .B2(new_n827), .ZN(G1338gat));
  INV_X1    g627(.A(G106gat), .ZN(new_n829));
  AOI21_X1  g628(.A(new_n829), .B1(new_n800), .B2(new_n554), .ZN(new_n830));
  NOR2_X1   g629(.A1(new_n791), .A2(G106gat), .ZN(new_n831));
  AND4_X1   g630(.A1(new_n697), .A2(new_n802), .A3(new_n804), .A4(new_n831), .ZN(new_n832));
  OAI21_X1  g631(.A(KEYINPUT53), .B1(new_n830), .B2(new_n832), .ZN(new_n833));
  OAI211_X1 g632(.A(new_n554), .B(new_n798), .C1(new_n733), .C2(new_n734), .ZN(new_n834));
  NAND2_X1  g633(.A1(new_n834), .A2(G106gat), .ZN(new_n835));
  INV_X1    g634(.A(KEYINPUT53), .ZN(new_n836));
  INV_X1    g635(.A(new_n831), .ZN(new_n837));
  OAI211_X1 g636(.A(new_n835), .B(new_n836), .C1(new_n810), .C2(new_n837), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n833), .A2(new_n838), .ZN(G1339gat));
  INV_X1    g638(.A(KEYINPUT54), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n675), .A2(new_n686), .ZN(new_n841));
  INV_X1    g640(.A(new_n668), .ZN(new_n842));
  AOI21_X1  g641(.A(new_n840), .B1(new_n841), .B2(new_n842), .ZN(new_n843));
  NAND3_X1  g642(.A1(new_n675), .A2(new_n686), .A3(new_n668), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  INV_X1    g644(.A(KEYINPUT113), .ZN(new_n846));
  AOI211_X1 g645(.A(new_n846), .B(new_n693), .C1(new_n687), .C2(new_n840), .ZN(new_n847));
  NAND3_X1  g646(.A1(new_n841), .A2(new_n840), .A3(new_n842), .ZN(new_n848));
  AOI21_X1  g647(.A(KEYINPUT113), .B1(new_n848), .B2(new_n694), .ZN(new_n849));
  OAI21_X1  g648(.A(new_n845), .B1(new_n847), .B2(new_n849), .ZN(new_n850));
  INV_X1    g649(.A(KEYINPUT55), .ZN(new_n851));
  NAND2_X1  g650(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  INV_X1    g651(.A(new_n696), .ZN(new_n853));
  AOI211_X1 g652(.A(KEYINPUT54), .B(new_n668), .C1(new_n675), .C2(new_n686), .ZN(new_n854));
  OAI21_X1  g653(.A(new_n846), .B1(new_n854), .B2(new_n693), .ZN(new_n855));
  NAND3_X1  g654(.A1(new_n848), .A2(KEYINPUT113), .A3(new_n694), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n855), .A2(new_n856), .ZN(new_n857));
  AOI21_X1  g656(.A(new_n851), .B1(new_n843), .B2(new_n844), .ZN(new_n858));
  AOI21_X1  g657(.A(new_n853), .B1(new_n857), .B2(new_n858), .ZN(new_n859));
  NAND3_X1  g658(.A1(new_n852), .A2(new_n859), .A3(new_n291), .ZN(new_n860));
  INV_X1    g659(.A(new_n281), .ZN(new_n861));
  AOI21_X1  g660(.A(new_n258), .B1(new_n257), .B2(new_n272), .ZN(new_n862));
  AND3_X1   g661(.A1(new_n272), .A2(new_n273), .A3(new_n269), .ZN(new_n863));
  OAI21_X1  g662(.A(new_n861), .B1(new_n862), .B2(new_n863), .ZN(new_n864));
  NAND3_X1  g663(.A1(new_n697), .A2(new_n284), .A3(new_n864), .ZN(new_n865));
  AOI21_X1  g664(.A(new_n661), .B1(new_n860), .B2(new_n865), .ZN(new_n866));
  OAI21_X1  g665(.A(new_n858), .B1(new_n847), .B2(new_n849), .ZN(new_n867));
  AND3_X1   g666(.A1(new_n675), .A2(new_n686), .A3(new_n668), .ZN(new_n868));
  NOR3_X1   g667(.A1(new_n868), .A2(new_n687), .A3(new_n840), .ZN(new_n869));
  AOI21_X1  g668(.A(new_n869), .B1(new_n855), .B2(new_n856), .ZN(new_n870));
  OAI211_X1 g669(.A(new_n696), .B(new_n867), .C1(new_n870), .C2(KEYINPUT55), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n284), .A2(new_n864), .ZN(new_n872));
  NOR3_X1   g671(.A1(new_n871), .A2(new_n663), .A3(new_n872), .ZN(new_n873));
  OAI21_X1  g672(.A(new_n624), .B1(new_n866), .B2(new_n873), .ZN(new_n874));
  INV_X1    g673(.A(new_n291), .ZN(new_n875));
  NAND4_X1  g674(.A1(new_n662), .A2(new_n665), .A3(new_n875), .A4(new_n776), .ZN(new_n876));
  AOI21_X1  g675(.A(new_n574), .B1(new_n874), .B2(new_n876), .ZN(new_n877));
  NAND4_X1  g676(.A1(new_n877), .A2(new_n536), .A3(new_n372), .A4(new_n535), .ZN(new_n878));
  OAI21_X1  g677(.A(G113gat), .B1(new_n878), .B2(new_n296), .ZN(new_n879));
  AND2_X1   g678(.A1(new_n877), .A2(new_n492), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n291), .A2(new_n320), .ZN(new_n881));
  XOR2_X1   g680(.A(new_n881), .B(KEYINPUT114), .Z(new_n882));
  NAND2_X1  g681(.A1(new_n880), .A2(new_n882), .ZN(new_n883));
  NAND2_X1  g682(.A1(new_n879), .A2(new_n883), .ZN(G1340gat));
  NOR3_X1   g683(.A1(new_n878), .A2(new_n321), .A3(new_n776), .ZN(new_n885));
  AOI21_X1  g684(.A(G120gat), .B1(new_n880), .B2(new_n697), .ZN(new_n886));
  NOR2_X1   g685(.A1(new_n885), .A2(new_n886), .ZN(G1341gat));
  OAI21_X1  g686(.A(G127gat), .B1(new_n878), .B2(new_n624), .ZN(new_n888));
  INV_X1    g687(.A(G127gat), .ZN(new_n889));
  NAND3_X1  g688(.A1(new_n880), .A2(new_n889), .A3(new_n723), .ZN(new_n890));
  NAND2_X1  g689(.A1(new_n888), .A2(new_n890), .ZN(G1342gat));
  INV_X1    g690(.A(G134gat), .ZN(new_n892));
  NAND3_X1  g691(.A1(new_n880), .A2(new_n892), .A3(new_n661), .ZN(new_n893));
  OR2_X1    g692(.A1(new_n893), .A2(KEYINPUT56), .ZN(new_n894));
  OAI21_X1  g693(.A(G134gat), .B1(new_n878), .B2(new_n663), .ZN(new_n895));
  NAND2_X1  g694(.A1(new_n893), .A2(KEYINPUT56), .ZN(new_n896));
  NAND3_X1  g695(.A1(new_n894), .A2(new_n895), .A3(new_n896), .ZN(G1343gat));
  AOI21_X1  g696(.A(new_n791), .B1(new_n712), .B2(new_n714), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n898), .A2(new_n877), .ZN(new_n899));
  NAND2_X1  g698(.A1(new_n899), .A2(KEYINPUT121), .ZN(new_n900));
  INV_X1    g699(.A(KEYINPUT121), .ZN(new_n901));
  NAND3_X1  g700(.A1(new_n898), .A2(new_n901), .A3(new_n877), .ZN(new_n902));
  AOI21_X1  g701(.A(new_n430), .B1(new_n900), .B2(new_n902), .ZN(new_n903));
  NOR2_X1   g702(.A1(new_n296), .A2(G141gat), .ZN(new_n904));
  XOR2_X1   g703(.A(new_n904), .B(KEYINPUT120), .Z(new_n905));
  NAND2_X1  g704(.A1(new_n903), .A2(new_n905), .ZN(new_n906));
  INV_X1    g705(.A(KEYINPUT58), .ZN(new_n907));
  INV_X1    g706(.A(KEYINPUT122), .ZN(new_n908));
  NOR3_X1   g707(.A1(new_n762), .A2(new_n574), .A3(new_n430), .ZN(new_n909));
  NAND2_X1  g708(.A1(new_n554), .A2(KEYINPUT57), .ZN(new_n910));
  XNOR2_X1  g709(.A(KEYINPUT117), .B(KEYINPUT55), .ZN(new_n911));
  INV_X1    g710(.A(new_n911), .ZN(new_n912));
  OAI211_X1 g711(.A(new_n696), .B(new_n867), .C1(new_n870), .C2(new_n912), .ZN(new_n913));
  INV_X1    g712(.A(KEYINPUT118), .ZN(new_n914));
  NAND2_X1  g713(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  NAND2_X1  g714(.A1(new_n850), .A2(new_n911), .ZN(new_n916));
  NAND3_X1  g715(.A1(new_n916), .A2(new_n859), .A3(KEYINPUT118), .ZN(new_n917));
  NAND3_X1  g716(.A1(new_n295), .A2(new_n915), .A3(new_n917), .ZN(new_n918));
  XNOR2_X1  g717(.A(new_n865), .B(KEYINPUT116), .ZN(new_n919));
  AOI21_X1  g718(.A(new_n661), .B1(new_n918), .B2(new_n919), .ZN(new_n920));
  OAI21_X1  g719(.A(new_n624), .B1(new_n920), .B2(new_n873), .ZN(new_n921));
  AOI21_X1  g720(.A(new_n910), .B1(new_n921), .B2(new_n876), .ZN(new_n922));
  XOR2_X1   g721(.A(KEYINPUT115), .B(KEYINPUT57), .Z(new_n923));
  INV_X1    g722(.A(new_n923), .ZN(new_n924));
  NAND2_X1  g723(.A1(new_n874), .A2(new_n876), .ZN(new_n925));
  AOI21_X1  g724(.A(new_n924), .B1(new_n925), .B2(new_n554), .ZN(new_n926));
  OAI21_X1  g725(.A(new_n909), .B1(new_n922), .B2(new_n926), .ZN(new_n927));
  OAI21_X1  g726(.A(new_n908), .B1(new_n927), .B2(new_n296), .ZN(new_n928));
  NAND2_X1  g727(.A1(new_n928), .A2(G141gat), .ZN(new_n929));
  NOR3_X1   g728(.A1(new_n927), .A2(new_n908), .A3(new_n296), .ZN(new_n930));
  OAI211_X1 g729(.A(new_n906), .B(new_n907), .C1(new_n929), .C2(new_n930), .ZN(new_n931));
  AND4_X1   g730(.A1(new_n536), .A2(new_n898), .A3(new_n877), .A4(new_n905), .ZN(new_n932));
  AOI21_X1  g731(.A(new_n293), .B1(new_n284), .B2(new_n290), .ZN(new_n933));
  AND3_X1   g732(.A1(new_n284), .A2(new_n290), .A3(new_n293), .ZN(new_n934));
  OAI22_X1  g733(.A1(new_n933), .A2(new_n934), .B1(new_n913), .B2(new_n914), .ZN(new_n935));
  AOI21_X1  g734(.A(KEYINPUT118), .B1(new_n916), .B2(new_n859), .ZN(new_n936));
  OAI21_X1  g735(.A(new_n919), .B1(new_n935), .B2(new_n936), .ZN(new_n937));
  AOI21_X1  g736(.A(new_n873), .B1(new_n937), .B2(new_n663), .ZN(new_n938));
  OAI21_X1  g737(.A(new_n876), .B1(new_n938), .B2(new_n723), .ZN(new_n939));
  INV_X1    g738(.A(new_n910), .ZN(new_n940));
  AOI21_X1  g739(.A(new_n926), .B1(new_n939), .B2(new_n940), .ZN(new_n941));
  INV_X1    g740(.A(new_n909), .ZN(new_n942));
  OAI21_X1  g741(.A(KEYINPUT119), .B1(new_n941), .B2(new_n942), .ZN(new_n943));
  INV_X1    g742(.A(KEYINPUT119), .ZN(new_n944));
  OAI211_X1 g743(.A(new_n944), .B(new_n909), .C1(new_n922), .C2(new_n926), .ZN(new_n945));
  NAND3_X1  g744(.A1(new_n943), .A2(new_n291), .A3(new_n945), .ZN(new_n946));
  AOI21_X1  g745(.A(new_n932), .B1(new_n946), .B2(G141gat), .ZN(new_n947));
  OAI21_X1  g746(.A(new_n931), .B1(new_n907), .B2(new_n947), .ZN(G1344gat));
  INV_X1    g747(.A(KEYINPUT59), .ZN(new_n949));
  OR2_X1    g748(.A1(new_n949), .A2(G148gat), .ZN(new_n950));
  AOI21_X1  g749(.A(new_n950), .B1(new_n903), .B2(new_n697), .ZN(new_n951));
  NAND3_X1  g750(.A1(new_n943), .A2(new_n697), .A3(new_n945), .ZN(new_n952));
  NAND2_X1  g751(.A1(new_n952), .A2(new_n949), .ZN(new_n953));
  OAI21_X1  g752(.A(KEYINPUT123), .B1(new_n871), .B2(new_n663), .ZN(new_n954));
  NAND3_X1  g753(.A1(new_n954), .A2(new_n284), .A3(new_n864), .ZN(new_n955));
  NOR3_X1   g754(.A1(new_n871), .A2(KEYINPUT123), .A3(new_n663), .ZN(new_n956));
  NOR2_X1   g755(.A1(new_n955), .A2(new_n956), .ZN(new_n957));
  OAI21_X1  g756(.A(new_n624), .B1(new_n957), .B2(new_n920), .ZN(new_n958));
  NAND2_X1  g757(.A1(new_n698), .A2(new_n296), .ZN(new_n959));
  NAND2_X1  g758(.A1(new_n958), .A2(new_n959), .ZN(new_n960));
  AOI21_X1  g759(.A(KEYINPUT57), .B1(new_n960), .B2(new_n554), .ZN(new_n961));
  AOI211_X1 g760(.A(new_n791), .B(new_n923), .C1(new_n874), .C2(new_n876), .ZN(new_n962));
  OR2_X1    g761(.A1(new_n961), .A2(new_n962), .ZN(new_n963));
  NAND4_X1  g762(.A1(new_n963), .A2(KEYINPUT59), .A3(new_n697), .A4(new_n909), .ZN(new_n964));
  NAND2_X1  g763(.A1(new_n953), .A2(new_n964), .ZN(new_n965));
  AOI21_X1  g764(.A(new_n951), .B1(new_n965), .B2(G148gat), .ZN(G1345gat));
  NAND2_X1  g765(.A1(new_n943), .A2(new_n945), .ZN(new_n967));
  OAI21_X1  g766(.A(G155gat), .B1(new_n967), .B2(new_n624), .ZN(new_n968));
  NAND3_X1  g767(.A1(new_n903), .A2(new_n439), .A3(new_n723), .ZN(new_n969));
  NAND2_X1  g768(.A1(new_n968), .A2(new_n969), .ZN(G1346gat));
  OAI21_X1  g769(.A(G162gat), .B1(new_n967), .B2(new_n663), .ZN(new_n971));
  NAND3_X1  g770(.A1(new_n903), .A2(new_n440), .A3(new_n661), .ZN(new_n972));
  NAND2_X1  g771(.A1(new_n971), .A2(new_n972), .ZN(G1347gat));
  AOI21_X1  g772(.A(new_n575), .B1(new_n874), .B2(new_n876), .ZN(new_n974));
  NOR3_X1   g773(.A1(new_n536), .A2(new_n491), .A3(new_n383), .ZN(new_n975));
  AND2_X1   g774(.A1(new_n974), .A2(new_n975), .ZN(new_n976));
  INV_X1    g775(.A(new_n976), .ZN(new_n977));
  OAI21_X1  g776(.A(G169gat), .B1(new_n977), .B2(new_n296), .ZN(new_n978));
  INV_X1    g777(.A(KEYINPUT125), .ZN(new_n979));
  INV_X1    g778(.A(new_n974), .ZN(new_n980));
  INV_X1    g779(.A(KEYINPUT124), .ZN(new_n981));
  AOI21_X1  g780(.A(new_n536), .B1(new_n980), .B2(new_n981), .ZN(new_n982));
  NAND2_X1  g781(.A1(new_n974), .A2(KEYINPUT124), .ZN(new_n983));
  AND2_X1   g782(.A1(new_n982), .A2(new_n983), .ZN(new_n984));
  NOR2_X1   g783(.A1(new_n386), .A2(new_n491), .ZN(new_n985));
  NAND2_X1  g784(.A1(new_n984), .A2(new_n985), .ZN(new_n986));
  INV_X1    g785(.A(new_n986), .ZN(new_n987));
  INV_X1    g786(.A(new_n333), .ZN(new_n988));
  NOR2_X1   g787(.A1(new_n875), .A2(new_n988), .ZN(new_n989));
  AOI21_X1  g788(.A(new_n979), .B1(new_n987), .B2(new_n989), .ZN(new_n990));
  NOR4_X1   g789(.A1(new_n986), .A2(KEYINPUT125), .A3(new_n988), .A4(new_n875), .ZN(new_n991));
  OAI21_X1  g790(.A(new_n978), .B1(new_n990), .B2(new_n991), .ZN(G1348gat));
  OAI21_X1  g791(.A(G176gat), .B1(new_n977), .B2(new_n776), .ZN(new_n993));
  NAND2_X1  g792(.A1(new_n697), .A2(new_n334), .ZN(new_n994));
  OAI21_X1  g793(.A(new_n993), .B1(new_n986), .B2(new_n994), .ZN(G1349gat));
  OAI21_X1  g794(.A(G183gat), .B1(new_n977), .B2(new_n624), .ZN(new_n996));
  NAND2_X1  g795(.A1(new_n723), .A2(new_n301), .ZN(new_n997));
  OAI21_X1  g796(.A(new_n996), .B1(new_n986), .B2(new_n997), .ZN(new_n998));
  XNOR2_X1  g797(.A(new_n998), .B(KEYINPUT60), .ZN(G1350gat));
  AOI21_X1  g798(.A(new_n297), .B1(new_n976), .B2(new_n661), .ZN(new_n1000));
  XOR2_X1   g799(.A(new_n1000), .B(KEYINPUT61), .Z(new_n1001));
  NAND2_X1  g800(.A1(new_n661), .A2(new_n297), .ZN(new_n1002));
  OAI21_X1  g801(.A(new_n1001), .B1(new_n986), .B2(new_n1002), .ZN(G1351gat));
  NAND2_X1  g802(.A1(new_n984), .A2(new_n898), .ZN(new_n1004));
  INV_X1    g803(.A(new_n1004), .ZN(new_n1005));
  AOI21_X1  g804(.A(G197gat), .B1(new_n1005), .B2(new_n291), .ZN(new_n1006));
  NOR3_X1   g805(.A1(new_n715), .A2(new_n575), .A3(new_n536), .ZN(new_n1007));
  AND2_X1   g806(.A1(new_n963), .A2(new_n1007), .ZN(new_n1008));
  NOR2_X1   g807(.A1(new_n296), .A2(new_n280), .ZN(new_n1009));
  AOI21_X1  g808(.A(new_n1006), .B1(new_n1008), .B2(new_n1009), .ZN(G1352gat));
  NAND3_X1  g809(.A1(new_n963), .A2(new_n697), .A3(new_n1007), .ZN(new_n1011));
  NAND2_X1  g810(.A1(new_n1011), .A2(G204gat), .ZN(new_n1012));
  OR2_X1    g811(.A1(new_n776), .A2(G204gat), .ZN(new_n1013));
  OR3_X1    g812(.A1(new_n1004), .A2(KEYINPUT62), .A3(new_n1013), .ZN(new_n1014));
  OAI21_X1  g813(.A(KEYINPUT62), .B1(new_n1004), .B2(new_n1013), .ZN(new_n1015));
  NAND3_X1  g814(.A1(new_n1012), .A2(new_n1014), .A3(new_n1015), .ZN(G1353gat));
  OAI211_X1 g815(.A(new_n1007), .B(new_n723), .C1(new_n961), .C2(new_n962), .ZN(new_n1017));
  NAND2_X1  g816(.A1(new_n1017), .A2(G211gat), .ZN(new_n1018));
  NAND2_X1  g817(.A1(new_n1018), .A2(KEYINPUT63), .ZN(new_n1019));
  INV_X1    g818(.A(KEYINPUT63), .ZN(new_n1020));
  NAND3_X1  g819(.A1(new_n1017), .A2(new_n1020), .A3(G211gat), .ZN(new_n1021));
  INV_X1    g820(.A(KEYINPUT126), .ZN(new_n1022));
  NOR2_X1   g821(.A1(new_n624), .A2(G211gat), .ZN(new_n1023));
  AOI21_X1  g822(.A(new_n1022), .B1(new_n1005), .B2(new_n1023), .ZN(new_n1024));
  NOR4_X1   g823(.A1(new_n1004), .A2(KEYINPUT126), .A3(G211gat), .A4(new_n624), .ZN(new_n1025));
  OAI211_X1 g824(.A(new_n1019), .B(new_n1021), .C1(new_n1024), .C2(new_n1025), .ZN(G1354gat));
  NOR2_X1   g825(.A1(new_n663), .A2(new_n406), .ZN(new_n1027));
  OAI211_X1 g826(.A(new_n1007), .B(new_n1027), .C1(new_n961), .C2(new_n962), .ZN(new_n1028));
  NAND4_X1  g827(.A1(new_n982), .A2(new_n661), .A3(new_n898), .A4(new_n983), .ZN(new_n1029));
  INV_X1    g828(.A(G218gat), .ZN(new_n1030));
  NAND2_X1  g829(.A1(new_n1029), .A2(new_n1030), .ZN(new_n1031));
  NAND2_X1  g830(.A1(new_n1028), .A2(new_n1031), .ZN(new_n1032));
  XNOR2_X1  g831(.A(new_n1032), .B(KEYINPUT127), .ZN(G1355gat));
endmodule


