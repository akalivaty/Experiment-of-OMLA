//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 1 0 0 0 1 0 0 0 1 0 1 1 0 1 0 1 0 1 0 0 1 1 1 0 0 1 1 1 1 0 1 1 1 1 1 1 1 1 0 0 1 0 1 1 1 1 1 1 0 0 1 0 0 0 0 0 0 1 0 1 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:29:41 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n456, new_n457,
    new_n458, new_n459, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n529, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n536, new_n537, new_n540, new_n541, new_n542,
    new_n543, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n553, new_n555, new_n556, new_n558, new_n559, new_n560, new_n561,
    new_n562, new_n563, new_n564, new_n565, new_n566, new_n567, new_n568,
    new_n570, new_n571, new_n572, new_n573, new_n575, new_n576, new_n577,
    new_n578, new_n579, new_n580, new_n581, new_n582, new_n583, new_n585,
    new_n586, new_n587, new_n588, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n602,
    new_n603, new_n606, new_n607, new_n609, new_n610, new_n611, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1133, new_n1134, new_n1135;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  XOR2_X1   g011(.A(KEYINPUT64), .B(G96), .Z(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G221), .A2(G220), .A3(G218), .A4(G219), .ZN(new_n450));
  XOR2_X1   g025(.A(KEYINPUT65), .B(KEYINPUT2), .Z(new_n451));
  XNOR2_X1  g026(.A(new_n450), .B(new_n451), .ZN(new_n452));
  NAND4_X1  g027(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n453));
  NOR2_X1   g028(.A1(new_n452), .A2(new_n453), .ZN(G325));
  INV_X1    g029(.A(G325), .ZN(G261));
  NAND2_X1  g030(.A1(new_n453), .A2(G567), .ZN(new_n456));
  NAND2_X1  g031(.A1(new_n452), .A2(G2106), .ZN(new_n457));
  INV_X1    g032(.A(KEYINPUT66), .ZN(new_n458));
  OAI21_X1  g033(.A(new_n456), .B1(new_n457), .B2(new_n458), .ZN(new_n459));
  AOI21_X1  g034(.A(new_n459), .B1(new_n458), .B2(new_n457), .ZN(G319));
  INV_X1    g035(.A(KEYINPUT68), .ZN(new_n461));
  AND2_X1   g036(.A1(KEYINPUT67), .A2(KEYINPUT3), .ZN(new_n462));
  NOR2_X1   g037(.A1(KEYINPUT67), .A2(KEYINPUT3), .ZN(new_n463));
  OAI211_X1 g038(.A(new_n461), .B(G2104), .C1(new_n462), .C2(new_n463), .ZN(new_n464));
  INV_X1    g039(.A(G2105), .ZN(new_n465));
  INV_X1    g040(.A(G2104), .ZN(new_n466));
  INV_X1    g041(.A(KEYINPUT67), .ZN(new_n467));
  INV_X1    g042(.A(KEYINPUT3), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  NAND2_X1  g044(.A1(KEYINPUT67), .A2(KEYINPUT3), .ZN(new_n470));
  AOI21_X1  g045(.A(new_n466), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  AOI21_X1  g046(.A(KEYINPUT68), .B1(new_n466), .B2(KEYINPUT3), .ZN(new_n472));
  OAI211_X1 g047(.A(new_n464), .B(new_n465), .C1(new_n471), .C2(new_n472), .ZN(new_n473));
  INV_X1    g048(.A(new_n473), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n474), .A2(G137), .ZN(new_n475));
  NAND2_X1  g050(.A1(G113), .A2(G2104), .ZN(new_n476));
  XOR2_X1   g051(.A(KEYINPUT3), .B(G2104), .Z(new_n477));
  INV_X1    g052(.A(G125), .ZN(new_n478));
  OAI21_X1  g053(.A(new_n476), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  NOR2_X1   g054(.A1(new_n466), .A2(G2105), .ZN(new_n480));
  AOI22_X1  g055(.A1(new_n479), .A2(G2105), .B1(G101), .B2(new_n480), .ZN(new_n481));
  AND2_X1   g056(.A1(new_n475), .A2(new_n481), .ZN(G160));
  NAND2_X1  g057(.A1(new_n474), .A2(G136), .ZN(new_n483));
  OAI211_X1 g058(.A(new_n464), .B(G2105), .C1(new_n471), .C2(new_n472), .ZN(new_n484));
  INV_X1    g059(.A(new_n484), .ZN(new_n485));
  NAND2_X1  g060(.A1(new_n485), .A2(G124), .ZN(new_n486));
  MUX2_X1   g061(.A(G100), .B(G112), .S(G2105), .Z(new_n487));
  NAND2_X1  g062(.A1(new_n487), .A2(G2104), .ZN(new_n488));
  NAND3_X1  g063(.A1(new_n483), .A2(new_n486), .A3(new_n488), .ZN(new_n489));
  INV_X1    g064(.A(new_n489), .ZN(G162));
  INV_X1    g065(.A(G138), .ZN(new_n491));
  NOR4_X1   g066(.A1(new_n477), .A2(KEYINPUT4), .A3(new_n491), .A4(G2105), .ZN(new_n492));
  OAI21_X1  g067(.A(G2104), .B1(new_n462), .B2(new_n463), .ZN(new_n493));
  INV_X1    g068(.A(new_n472), .ZN(new_n494));
  NAND2_X1  g069(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  NAND4_X1  g070(.A1(new_n495), .A2(G138), .A3(new_n465), .A4(new_n464), .ZN(new_n496));
  AOI21_X1  g071(.A(new_n492), .B1(new_n496), .B2(KEYINPUT4), .ZN(new_n497));
  INV_X1    g072(.A(G114), .ZN(new_n498));
  AND3_X1   g073(.A1(new_n498), .A2(KEYINPUT69), .A3(G2105), .ZN(new_n499));
  AOI21_X1  g074(.A(KEYINPUT69), .B1(new_n498), .B2(G2105), .ZN(new_n500));
  OAI221_X1 g075(.A(G2104), .B1(G102), .B2(G2105), .C1(new_n499), .C2(new_n500), .ZN(new_n501));
  INV_X1    g076(.A(G126), .ZN(new_n502));
  OAI21_X1  g077(.A(new_n501), .B1(new_n484), .B2(new_n502), .ZN(new_n503));
  NOR2_X1   g078(.A1(new_n497), .A2(new_n503), .ZN(G164));
  NAND2_X1  g079(.A1(G75), .A2(G543), .ZN(new_n505));
  INV_X1    g080(.A(KEYINPUT5), .ZN(new_n506));
  INV_X1    g081(.A(G543), .ZN(new_n507));
  OR3_X1    g082(.A1(new_n506), .A2(new_n507), .A3(KEYINPUT71), .ZN(new_n508));
  OAI21_X1  g083(.A(new_n507), .B1(new_n506), .B2(KEYINPUT71), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  INV_X1    g085(.A(new_n510), .ZN(new_n511));
  INV_X1    g086(.A(G62), .ZN(new_n512));
  OAI21_X1  g087(.A(new_n505), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n513), .A2(G651), .ZN(new_n514));
  INV_X1    g089(.A(KEYINPUT6), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n515), .A2(G651), .ZN(new_n516));
  XNOR2_X1  g091(.A(new_n516), .B(KEYINPUT70), .ZN(new_n517));
  INV_X1    g092(.A(G651), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n518), .A2(KEYINPUT6), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n517), .A2(new_n519), .ZN(new_n520));
  INV_X1    g095(.A(new_n520), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n521), .A2(new_n510), .ZN(new_n522));
  INV_X1    g097(.A(G88), .ZN(new_n523));
  INV_X1    g098(.A(G50), .ZN(new_n524));
  NOR2_X1   g099(.A1(new_n520), .A2(new_n507), .ZN(new_n525));
  INV_X1    g100(.A(new_n525), .ZN(new_n526));
  OAI221_X1 g101(.A(new_n514), .B1(new_n522), .B2(new_n523), .C1(new_n524), .C2(new_n526), .ZN(G303));
  INV_X1    g102(.A(G303), .ZN(G166));
  NAND2_X1  g103(.A1(new_n525), .A2(G51), .ZN(new_n529));
  NOR2_X1   g104(.A1(new_n520), .A2(new_n511), .ZN(new_n530));
  XOR2_X1   g105(.A(KEYINPUT72), .B(G89), .Z(new_n531));
  NAND2_X1  g106(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  AND2_X1   g107(.A1(G63), .A2(G651), .ZN(new_n533));
  NAND3_X1  g108(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n534));
  NAND2_X1  g109(.A1(new_n534), .A2(KEYINPUT7), .ZN(new_n535));
  OR2_X1    g110(.A1(new_n534), .A2(KEYINPUT7), .ZN(new_n536));
  AOI22_X1  g111(.A1(new_n510), .A2(new_n533), .B1(new_n535), .B2(new_n536), .ZN(new_n537));
  NAND3_X1  g112(.A1(new_n529), .A2(new_n532), .A3(new_n537), .ZN(G286));
  INV_X1    g113(.A(G286), .ZN(G168));
  AOI22_X1  g114(.A1(new_n510), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n540));
  OR2_X1    g115(.A1(new_n540), .A2(new_n518), .ZN(new_n541));
  NAND2_X1  g116(.A1(new_n530), .A2(G90), .ZN(new_n542));
  NAND2_X1  g117(.A1(new_n525), .A2(G52), .ZN(new_n543));
  NAND3_X1  g118(.A1(new_n541), .A2(new_n542), .A3(new_n543), .ZN(G301));
  INV_X1    g119(.A(G301), .ZN(G171));
  AOI22_X1  g120(.A1(G43), .A2(new_n525), .B1(new_n530), .B2(G81), .ZN(new_n546));
  INV_X1    g121(.A(KEYINPUT73), .ZN(new_n547));
  XNOR2_X1  g122(.A(new_n546), .B(new_n547), .ZN(new_n548));
  AOI22_X1  g123(.A1(new_n510), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n549));
  OR2_X1    g124(.A1(new_n549), .A2(new_n518), .ZN(new_n550));
  AND2_X1   g125(.A1(new_n548), .A2(new_n550), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n551), .A2(G860), .ZN(G153));
  AND3_X1   g127(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n553), .A2(G36), .ZN(G176));
  NAND2_X1  g129(.A1(G1), .A2(G3), .ZN(new_n555));
  XNOR2_X1  g130(.A(new_n555), .B(KEYINPUT8), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n553), .A2(new_n556), .ZN(G188));
  NAND2_X1  g132(.A1(new_n525), .A2(G53), .ZN(new_n558));
  INV_X1    g133(.A(KEYINPUT74), .ZN(new_n559));
  NOR2_X1   g134(.A1(new_n559), .A2(KEYINPUT9), .ZN(new_n560));
  OR2_X1    g135(.A1(new_n558), .A2(new_n560), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n558), .A2(new_n560), .ZN(new_n562));
  AOI22_X1  g137(.A1(new_n561), .A2(new_n562), .B1(new_n559), .B2(KEYINPUT9), .ZN(new_n563));
  AOI22_X1  g138(.A1(new_n510), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n564));
  INV_X1    g139(.A(new_n564), .ZN(new_n565));
  AOI22_X1  g140(.A1(G651), .A2(new_n565), .B1(new_n530), .B2(G91), .ZN(new_n566));
  INV_X1    g141(.A(new_n566), .ZN(new_n567));
  NOR2_X1   g142(.A1(new_n563), .A2(new_n567), .ZN(new_n568));
  INV_X1    g143(.A(new_n568), .ZN(G299));
  NAND2_X1  g144(.A1(new_n530), .A2(G87), .ZN(new_n570));
  NAND2_X1  g145(.A1(new_n525), .A2(G49), .ZN(new_n571));
  OAI21_X1  g146(.A(G651), .B1(new_n510), .B2(G74), .ZN(new_n572));
  NAND3_X1  g147(.A1(new_n570), .A2(new_n571), .A3(new_n572), .ZN(new_n573));
  XOR2_X1   g148(.A(new_n573), .B(KEYINPUT75), .Z(G288));
  INV_X1    g149(.A(G48), .ZN(new_n575));
  OAI21_X1  g150(.A(KEYINPUT76), .B1(new_n526), .B2(new_n575), .ZN(new_n576));
  INV_X1    g151(.A(KEYINPUT76), .ZN(new_n577));
  NAND3_X1  g152(.A1(new_n525), .A2(new_n577), .A3(G48), .ZN(new_n578));
  NAND2_X1  g153(.A1(new_n576), .A2(new_n578), .ZN(new_n579));
  NAND2_X1  g154(.A1(G73), .A2(G543), .ZN(new_n580));
  INV_X1    g155(.A(G61), .ZN(new_n581));
  OAI21_X1  g156(.A(new_n580), .B1(new_n511), .B2(new_n581), .ZN(new_n582));
  AOI22_X1  g157(.A1(G86), .A2(new_n530), .B1(new_n582), .B2(G651), .ZN(new_n583));
  NAND2_X1  g158(.A1(new_n579), .A2(new_n583), .ZN(G305));
  AOI22_X1  g159(.A1(new_n510), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n585));
  OR2_X1    g160(.A1(new_n585), .A2(new_n518), .ZN(new_n586));
  NAND2_X1  g161(.A1(new_n530), .A2(G85), .ZN(new_n587));
  NAND2_X1  g162(.A1(new_n525), .A2(G47), .ZN(new_n588));
  NAND3_X1  g163(.A1(new_n586), .A2(new_n587), .A3(new_n588), .ZN(G290));
  NAND2_X1  g164(.A1(G301), .A2(G868), .ZN(new_n590));
  XNOR2_X1  g165(.A(new_n590), .B(KEYINPUT77), .ZN(new_n591));
  NAND2_X1  g166(.A1(new_n525), .A2(G54), .ZN(new_n592));
  AOI22_X1  g167(.A1(new_n510), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n593));
  NAND2_X1  g168(.A1(new_n530), .A2(G92), .ZN(new_n594));
  INV_X1    g169(.A(KEYINPUT10), .ZN(new_n595));
  NOR2_X1   g170(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  AOI21_X1  g171(.A(KEYINPUT10), .B1(new_n530), .B2(G92), .ZN(new_n597));
  OAI221_X1 g172(.A(new_n592), .B1(new_n518), .B2(new_n593), .C1(new_n596), .C2(new_n597), .ZN(new_n598));
  XNOR2_X1  g173(.A(new_n598), .B(KEYINPUT78), .ZN(new_n599));
  OAI21_X1  g174(.A(new_n591), .B1(new_n599), .B2(G868), .ZN(G284));
  OAI21_X1  g175(.A(new_n591), .B1(new_n599), .B2(G868), .ZN(G321));
  INV_X1    g176(.A(G868), .ZN(new_n602));
  NOR2_X1   g177(.A1(G286), .A2(new_n602), .ZN(new_n603));
  AOI21_X1  g178(.A(new_n603), .B1(new_n568), .B2(new_n602), .ZN(G297));
  AOI21_X1  g179(.A(new_n603), .B1(new_n568), .B2(new_n602), .ZN(G280));
  INV_X1    g180(.A(G559), .ZN(new_n606));
  OAI21_X1  g181(.A(new_n599), .B1(new_n606), .B2(G860), .ZN(new_n607));
  XNOR2_X1  g182(.A(new_n607), .B(KEYINPUT79), .ZN(G148));
  NAND2_X1  g183(.A1(new_n551), .A2(new_n602), .ZN(new_n609));
  NAND2_X1  g184(.A1(new_n599), .A2(new_n606), .ZN(new_n610));
  OAI21_X1  g185(.A(new_n609), .B1(new_n610), .B2(new_n602), .ZN(new_n611));
  XNOR2_X1  g186(.A(new_n611), .B(KEYINPUT80), .ZN(G323));
  XNOR2_X1  g187(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g188(.A1(new_n474), .A2(G135), .ZN(new_n614));
  NAND2_X1  g189(.A1(new_n485), .A2(G123), .ZN(new_n615));
  AND2_X1   g190(.A1(G111), .A2(G2105), .ZN(new_n616));
  AOI21_X1  g191(.A(new_n616), .B1(G99), .B2(new_n465), .ZN(new_n617));
  OAI211_X1 g192(.A(new_n614), .B(new_n615), .C1(new_n466), .C2(new_n617), .ZN(new_n618));
  OR2_X1    g193(.A1(new_n618), .A2(G2096), .ZN(new_n619));
  NAND2_X1  g194(.A1(new_n618), .A2(G2096), .ZN(new_n620));
  XNOR2_X1  g195(.A(KEYINPUT81), .B(KEYINPUT13), .ZN(new_n621));
  XNOR2_X1  g196(.A(new_n621), .B(G2100), .ZN(new_n622));
  NAND3_X1  g197(.A1(new_n465), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n623));
  XOR2_X1   g198(.A(new_n623), .B(KEYINPUT12), .Z(new_n624));
  XOR2_X1   g199(.A(new_n622), .B(new_n624), .Z(new_n625));
  NAND3_X1  g200(.A1(new_n619), .A2(new_n620), .A3(new_n625), .ZN(G156));
  INV_X1    g201(.A(G14), .ZN(new_n627));
  XOR2_X1   g202(.A(KEYINPUT15), .B(G2435), .Z(new_n628));
  XNOR2_X1  g203(.A(new_n628), .B(G2438), .ZN(new_n629));
  XNOR2_X1  g204(.A(new_n629), .B(G2427), .ZN(new_n630));
  INV_X1    g205(.A(G2430), .ZN(new_n631));
  OR2_X1    g206(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  NAND2_X1  g207(.A1(new_n630), .A2(new_n631), .ZN(new_n633));
  NAND3_X1  g208(.A1(new_n632), .A2(KEYINPUT14), .A3(new_n633), .ZN(new_n634));
  XNOR2_X1  g209(.A(G2451), .B(G2454), .ZN(new_n635));
  XNOR2_X1  g210(.A(new_n635), .B(KEYINPUT16), .ZN(new_n636));
  XOR2_X1   g211(.A(G2443), .B(G2446), .Z(new_n637));
  XNOR2_X1  g212(.A(new_n636), .B(new_n637), .ZN(new_n638));
  XNOR2_X1  g213(.A(new_n634), .B(new_n638), .ZN(new_n639));
  XNOR2_X1  g214(.A(G1341), .B(G1348), .ZN(new_n640));
  INV_X1    g215(.A(new_n640), .ZN(new_n641));
  NOR2_X1   g216(.A1(new_n639), .A2(new_n641), .ZN(new_n642));
  XOR2_X1   g217(.A(new_n642), .B(KEYINPUT82), .Z(new_n643));
  AOI211_X1 g218(.A(new_n627), .B(new_n643), .C1(new_n639), .C2(new_n641), .ZN(G401));
  XOR2_X1   g219(.A(G2072), .B(G2078), .Z(new_n645));
  XOR2_X1   g220(.A(new_n645), .B(KEYINPUT17), .Z(new_n646));
  XOR2_X1   g221(.A(G2084), .B(G2090), .Z(new_n647));
  INV_X1    g222(.A(new_n647), .ZN(new_n648));
  XNOR2_X1  g223(.A(G2067), .B(G2678), .ZN(new_n649));
  NOR3_X1   g224(.A1(new_n646), .A2(new_n648), .A3(new_n649), .ZN(new_n650));
  XNOR2_X1  g225(.A(new_n650), .B(KEYINPUT84), .ZN(new_n651));
  NAND2_X1  g226(.A1(new_n646), .A2(new_n649), .ZN(new_n652));
  INV_X1    g227(.A(new_n645), .ZN(new_n653));
  OAI211_X1 g228(.A(new_n652), .B(new_n648), .C1(new_n653), .C2(new_n649), .ZN(new_n654));
  NAND3_X1  g229(.A1(new_n653), .A2(new_n647), .A3(new_n649), .ZN(new_n655));
  XOR2_X1   g230(.A(KEYINPUT83), .B(KEYINPUT18), .Z(new_n656));
  XNOR2_X1  g231(.A(new_n655), .B(new_n656), .ZN(new_n657));
  NAND3_X1  g232(.A1(new_n651), .A2(new_n654), .A3(new_n657), .ZN(new_n658));
  XOR2_X1   g233(.A(new_n658), .B(G2096), .Z(new_n659));
  XOR2_X1   g234(.A(KEYINPUT85), .B(G2100), .Z(new_n660));
  XNOR2_X1  g235(.A(new_n659), .B(new_n660), .ZN(G227));
  XOR2_X1   g236(.A(G1971), .B(G1976), .Z(new_n662));
  XNOR2_X1  g237(.A(new_n662), .B(KEYINPUT19), .ZN(new_n663));
  XNOR2_X1  g238(.A(G1956), .B(G2474), .ZN(new_n664));
  XNOR2_X1  g239(.A(G1961), .B(G1966), .ZN(new_n665));
  NOR2_X1   g240(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  AND2_X1   g241(.A1(new_n664), .A2(new_n665), .ZN(new_n667));
  NOR3_X1   g242(.A1(new_n663), .A2(new_n666), .A3(new_n667), .ZN(new_n668));
  NAND2_X1  g243(.A1(new_n663), .A2(new_n666), .ZN(new_n669));
  XOR2_X1   g244(.A(new_n669), .B(KEYINPUT20), .Z(new_n670));
  AOI211_X1 g245(.A(new_n668), .B(new_n670), .C1(new_n663), .C2(new_n667), .ZN(new_n671));
  XOR2_X1   g246(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n672));
  XOR2_X1   g247(.A(new_n671), .B(new_n672), .Z(new_n673));
  XNOR2_X1  g248(.A(G1991), .B(G1996), .ZN(new_n674));
  XNOR2_X1  g249(.A(G1981), .B(G1986), .ZN(new_n675));
  XNOR2_X1  g250(.A(new_n674), .B(new_n675), .ZN(new_n676));
  XNOR2_X1  g251(.A(new_n673), .B(new_n676), .ZN(new_n677));
  INV_X1    g252(.A(new_n677), .ZN(G229));
  MUX2_X1   g253(.A(G6), .B(G305), .S(G16), .Z(new_n679));
  XNOR2_X1  g254(.A(KEYINPUT32), .B(G1981), .ZN(new_n680));
  XNOR2_X1  g255(.A(new_n679), .B(new_n680), .ZN(new_n681));
  INV_X1    g256(.A(G16), .ZN(new_n682));
  NAND2_X1  g257(.A1(new_n682), .A2(G23), .ZN(new_n683));
  INV_X1    g258(.A(new_n573), .ZN(new_n684));
  OAI21_X1  g259(.A(new_n683), .B1(new_n684), .B2(new_n682), .ZN(new_n685));
  XOR2_X1   g260(.A(KEYINPUT33), .B(G1976), .Z(new_n686));
  XNOR2_X1  g261(.A(new_n685), .B(new_n686), .ZN(new_n687));
  NAND2_X1  g262(.A1(new_n682), .A2(G22), .ZN(new_n688));
  XOR2_X1   g263(.A(new_n688), .B(KEYINPUT90), .Z(new_n689));
  OAI21_X1  g264(.A(new_n689), .B1(G166), .B2(new_n682), .ZN(new_n690));
  XNOR2_X1  g265(.A(KEYINPUT91), .B(G1971), .ZN(new_n691));
  XNOR2_X1  g266(.A(new_n690), .B(new_n691), .ZN(new_n692));
  NOR3_X1   g267(.A1(new_n681), .A2(new_n687), .A3(new_n692), .ZN(new_n693));
  INV_X1    g268(.A(KEYINPUT34), .ZN(new_n694));
  OR2_X1    g269(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  INV_X1    g270(.A(G29), .ZN(new_n696));
  NAND2_X1  g271(.A1(new_n696), .A2(G25), .ZN(new_n697));
  XNOR2_X1  g272(.A(new_n697), .B(KEYINPUT86), .ZN(new_n698));
  NAND2_X1  g273(.A1(new_n474), .A2(G131), .ZN(new_n699));
  XNOR2_X1  g274(.A(new_n699), .B(KEYINPUT87), .ZN(new_n700));
  NAND2_X1  g275(.A1(new_n485), .A2(G119), .ZN(new_n701));
  OAI21_X1  g276(.A(KEYINPUT88), .B1(G95), .B2(G2105), .ZN(new_n702));
  INV_X1    g277(.A(new_n702), .ZN(new_n703));
  NOR3_X1   g278(.A1(KEYINPUT88), .A2(G95), .A3(G2105), .ZN(new_n704));
  OAI221_X1 g279(.A(G2104), .B1(G107), .B2(new_n465), .C1(new_n703), .C2(new_n704), .ZN(new_n705));
  AND2_X1   g280(.A1(new_n701), .A2(new_n705), .ZN(new_n706));
  NAND2_X1  g281(.A1(new_n700), .A2(new_n706), .ZN(new_n707));
  INV_X1    g282(.A(new_n707), .ZN(new_n708));
  OAI21_X1  g283(.A(new_n698), .B1(new_n708), .B2(new_n696), .ZN(new_n709));
  XNOR2_X1  g284(.A(new_n709), .B(KEYINPUT89), .ZN(new_n710));
  XOR2_X1   g285(.A(KEYINPUT35), .B(G1991), .Z(new_n711));
  INV_X1    g286(.A(new_n711), .ZN(new_n712));
  XNOR2_X1  g287(.A(new_n710), .B(new_n712), .ZN(new_n713));
  NAND2_X1  g288(.A1(new_n693), .A2(new_n694), .ZN(new_n714));
  OR2_X1    g289(.A1(G16), .A2(G24), .ZN(new_n715));
  OAI21_X1  g290(.A(new_n715), .B1(G290), .B2(new_n682), .ZN(new_n716));
  INV_X1    g291(.A(G1986), .ZN(new_n717));
  OAI21_X1  g292(.A(KEYINPUT92), .B1(new_n716), .B2(new_n717), .ZN(new_n718));
  AOI21_X1  g293(.A(new_n718), .B1(new_n717), .B2(new_n716), .ZN(new_n719));
  NAND4_X1  g294(.A1(new_n695), .A2(new_n713), .A3(new_n714), .A4(new_n719), .ZN(new_n720));
  INV_X1    g295(.A(new_n720), .ZN(new_n721));
  OR2_X1    g296(.A1(new_n721), .A2(KEYINPUT36), .ZN(new_n722));
  NAND2_X1  g297(.A1(new_n721), .A2(KEYINPUT36), .ZN(new_n723));
  NOR2_X1   g298(.A1(G171), .A2(new_n682), .ZN(new_n724));
  AOI21_X1  g299(.A(new_n724), .B1(G5), .B2(new_n682), .ZN(new_n725));
  INV_X1    g300(.A(G1961), .ZN(new_n726));
  NAND2_X1  g301(.A1(new_n682), .A2(G21), .ZN(new_n727));
  OAI21_X1  g302(.A(new_n727), .B1(G168), .B2(new_n682), .ZN(new_n728));
  OAI22_X1  g303(.A1(new_n725), .A2(new_n726), .B1(new_n728), .B2(G1966), .ZN(new_n729));
  NAND2_X1  g304(.A1(new_n725), .A2(new_n726), .ZN(new_n730));
  XOR2_X1   g305(.A(KEYINPUT31), .B(G11), .Z(new_n731));
  INV_X1    g306(.A(KEYINPUT30), .ZN(new_n732));
  OAI21_X1  g307(.A(new_n696), .B1(new_n732), .B2(G28), .ZN(new_n733));
  NOR2_X1   g308(.A1(new_n733), .A2(KEYINPUT98), .ZN(new_n734));
  AOI21_X1  g309(.A(new_n734), .B1(new_n732), .B2(G28), .ZN(new_n735));
  NAND2_X1  g310(.A1(new_n733), .A2(KEYINPUT98), .ZN(new_n736));
  AOI21_X1  g311(.A(new_n731), .B1(new_n735), .B2(new_n736), .ZN(new_n737));
  OAI211_X1 g312(.A(new_n730), .B(new_n737), .C1(new_n696), .C2(new_n618), .ZN(new_n738));
  XOR2_X1   g313(.A(KEYINPUT27), .B(G1996), .Z(new_n739));
  XNOR2_X1  g314(.A(new_n739), .B(KEYINPUT96), .ZN(new_n740));
  NAND3_X1  g315(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n741));
  INV_X1    g316(.A(KEYINPUT26), .ZN(new_n742));
  OR2_X1    g317(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  NAND2_X1  g318(.A1(new_n741), .A2(new_n742), .ZN(new_n744));
  AOI22_X1  g319(.A1(new_n743), .A2(new_n744), .B1(G105), .B2(new_n480), .ZN(new_n745));
  INV_X1    g320(.A(G141), .ZN(new_n746));
  INV_X1    g321(.A(G129), .ZN(new_n747));
  OAI221_X1 g322(.A(new_n745), .B1(new_n473), .B2(new_n746), .C1(new_n747), .C2(new_n484), .ZN(new_n748));
  MUX2_X1   g323(.A(G32), .B(new_n748), .S(G29), .Z(new_n749));
  AOI211_X1 g324(.A(new_n729), .B(new_n738), .C1(new_n740), .C2(new_n749), .ZN(new_n750));
  NOR2_X1   g325(.A1(G29), .A2(G35), .ZN(new_n751));
  AOI21_X1  g326(.A(new_n751), .B1(G162), .B2(G29), .ZN(new_n752));
  XNOR2_X1  g327(.A(KEYINPUT100), .B(KEYINPUT29), .ZN(new_n753));
  XNOR2_X1  g328(.A(new_n752), .B(new_n753), .ZN(new_n754));
  NAND2_X1  g329(.A1(new_n754), .A2(G2090), .ZN(new_n755));
  OR2_X1    g330(.A1(new_n754), .A2(G2090), .ZN(new_n756));
  NOR2_X1   g331(.A1(new_n749), .A2(new_n740), .ZN(new_n757));
  XOR2_X1   g332(.A(new_n757), .B(KEYINPUT97), .Z(new_n758));
  NAND4_X1  g333(.A1(new_n750), .A2(new_n755), .A3(new_n756), .A4(new_n758), .ZN(new_n759));
  NAND2_X1  g334(.A1(new_n474), .A2(G139), .ZN(new_n760));
  AOI21_X1  g335(.A(KEYINPUT25), .B1(new_n480), .B2(G103), .ZN(new_n761));
  AND3_X1   g336(.A1(new_n480), .A2(KEYINPUT25), .A3(G103), .ZN(new_n762));
  INV_X1    g337(.A(G127), .ZN(new_n763));
  NOR2_X1   g338(.A1(new_n477), .A2(new_n763), .ZN(new_n764));
  AOI21_X1  g339(.A(new_n764), .B1(G115), .B2(G2104), .ZN(new_n765));
  OAI221_X1 g340(.A(new_n760), .B1(new_n761), .B2(new_n762), .C1(new_n465), .C2(new_n765), .ZN(new_n766));
  MUX2_X1   g341(.A(G33), .B(new_n766), .S(G29), .Z(new_n767));
  XNOR2_X1  g342(.A(new_n767), .B(KEYINPUT95), .ZN(new_n768));
  XNOR2_X1  g343(.A(new_n768), .B(G2072), .ZN(new_n769));
  NAND2_X1  g344(.A1(new_n682), .A2(G19), .ZN(new_n770));
  XOR2_X1   g345(.A(new_n770), .B(KEYINPUT93), .Z(new_n771));
  NAND2_X1  g346(.A1(new_n548), .A2(new_n550), .ZN(new_n772));
  AOI21_X1  g347(.A(new_n771), .B1(new_n772), .B2(G16), .ZN(new_n773));
  XNOR2_X1  g348(.A(new_n773), .B(G1341), .ZN(new_n774));
  NOR2_X1   g349(.A1(G27), .A2(G29), .ZN(new_n775));
  AOI21_X1  g350(.A(new_n775), .B1(G164), .B2(G29), .ZN(new_n776));
  XOR2_X1   g351(.A(KEYINPUT99), .B(G2078), .Z(new_n777));
  XNOR2_X1  g352(.A(new_n776), .B(new_n777), .ZN(new_n778));
  NAND3_X1  g353(.A1(new_n769), .A2(new_n774), .A3(new_n778), .ZN(new_n779));
  NAND2_X1  g354(.A1(new_n728), .A2(G1966), .ZN(new_n780));
  INV_X1    g355(.A(G2084), .ZN(new_n781));
  AND2_X1   g356(.A1(KEYINPUT24), .A2(G34), .ZN(new_n782));
  NOR2_X1   g357(.A1(KEYINPUT24), .A2(G34), .ZN(new_n783));
  OAI21_X1  g358(.A(new_n696), .B1(new_n782), .B2(new_n783), .ZN(new_n784));
  INV_X1    g359(.A(G160), .ZN(new_n785));
  OAI21_X1  g360(.A(new_n784), .B1(new_n785), .B2(new_n696), .ZN(new_n786));
  OAI21_X1  g361(.A(new_n780), .B1(new_n781), .B2(new_n786), .ZN(new_n787));
  NAND2_X1  g362(.A1(new_n682), .A2(G20), .ZN(new_n788));
  XNOR2_X1  g363(.A(new_n788), .B(KEYINPUT23), .ZN(new_n789));
  OAI21_X1  g364(.A(new_n789), .B1(new_n568), .B2(new_n682), .ZN(new_n790));
  XNOR2_X1  g365(.A(KEYINPUT101), .B(G1956), .ZN(new_n791));
  NOR2_X1   g366(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  AOI211_X1 g367(.A(new_n787), .B(new_n792), .C1(new_n781), .C2(new_n786), .ZN(new_n793));
  NOR2_X1   g368(.A1(G4), .A2(G16), .ZN(new_n794));
  AOI21_X1  g369(.A(new_n794), .B1(new_n599), .B2(G16), .ZN(new_n795));
  INV_X1    g370(.A(G1348), .ZN(new_n796));
  XNOR2_X1  g371(.A(new_n795), .B(new_n796), .ZN(new_n797));
  MUX2_X1   g372(.A(G104), .B(G116), .S(G2105), .Z(new_n798));
  AOI22_X1  g373(.A1(new_n485), .A2(G128), .B1(G2104), .B2(new_n798), .ZN(new_n799));
  INV_X1    g374(.A(G140), .ZN(new_n800));
  OAI21_X1  g375(.A(new_n799), .B1(new_n800), .B2(new_n473), .ZN(new_n801));
  NAND2_X1  g376(.A1(new_n801), .A2(G29), .ZN(new_n802));
  NAND2_X1  g377(.A1(new_n696), .A2(G26), .ZN(new_n803));
  XNOR2_X1  g378(.A(new_n803), .B(KEYINPUT94), .ZN(new_n804));
  XNOR2_X1  g379(.A(new_n804), .B(KEYINPUT28), .ZN(new_n805));
  NAND2_X1  g380(.A1(new_n802), .A2(new_n805), .ZN(new_n806));
  XNOR2_X1  g381(.A(new_n806), .B(G2067), .ZN(new_n807));
  AOI21_X1  g382(.A(new_n807), .B1(new_n790), .B2(new_n791), .ZN(new_n808));
  NAND3_X1  g383(.A1(new_n793), .A2(new_n797), .A3(new_n808), .ZN(new_n809));
  NOR3_X1   g384(.A1(new_n759), .A2(new_n779), .A3(new_n809), .ZN(new_n810));
  NAND3_X1  g385(.A1(new_n722), .A2(new_n723), .A3(new_n810), .ZN(G150));
  INV_X1    g386(.A(G150), .ZN(G311));
  NAND2_X1  g387(.A1(new_n530), .A2(G93), .ZN(new_n813));
  NAND2_X1  g388(.A1(new_n525), .A2(G55), .ZN(new_n814));
  AOI22_X1  g389(.A1(new_n510), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n815));
  OAI211_X1 g390(.A(new_n813), .B(new_n814), .C1(new_n518), .C2(new_n815), .ZN(new_n816));
  NAND2_X1  g391(.A1(new_n816), .A2(G860), .ZN(new_n817));
  XOR2_X1   g392(.A(new_n817), .B(KEYINPUT37), .Z(new_n818));
  OR2_X1    g393(.A1(new_n816), .A2(KEYINPUT102), .ZN(new_n819));
  NAND2_X1  g394(.A1(new_n816), .A2(KEYINPUT102), .ZN(new_n820));
  NAND3_X1  g395(.A1(new_n551), .A2(new_n819), .A3(new_n820), .ZN(new_n821));
  NAND3_X1  g396(.A1(new_n772), .A2(KEYINPUT102), .A3(new_n816), .ZN(new_n822));
  NAND2_X1  g397(.A1(new_n821), .A2(new_n822), .ZN(new_n823));
  INV_X1    g398(.A(new_n823), .ZN(new_n824));
  INV_X1    g399(.A(KEYINPUT78), .ZN(new_n825));
  XNOR2_X1  g400(.A(new_n598), .B(new_n825), .ZN(new_n826));
  OAI21_X1  g401(.A(KEYINPUT38), .B1(new_n826), .B2(new_n606), .ZN(new_n827));
  INV_X1    g402(.A(KEYINPUT38), .ZN(new_n828));
  NAND3_X1  g403(.A1(new_n599), .A2(new_n828), .A3(G559), .ZN(new_n829));
  AND3_X1   g404(.A1(new_n824), .A2(new_n827), .A3(new_n829), .ZN(new_n830));
  AOI21_X1  g405(.A(new_n824), .B1(new_n827), .B2(new_n829), .ZN(new_n831));
  NOR2_X1   g406(.A1(new_n830), .A2(new_n831), .ZN(new_n832));
  OAI21_X1  g407(.A(KEYINPUT103), .B1(new_n832), .B2(KEYINPUT39), .ZN(new_n833));
  INV_X1    g408(.A(KEYINPUT103), .ZN(new_n834));
  INV_X1    g409(.A(KEYINPUT39), .ZN(new_n835));
  OAI211_X1 g410(.A(new_n834), .B(new_n835), .C1(new_n830), .C2(new_n831), .ZN(new_n836));
  NAND2_X1  g411(.A1(new_n833), .A2(new_n836), .ZN(new_n837));
  AOI21_X1  g412(.A(G860), .B1(new_n832), .B2(KEYINPUT39), .ZN(new_n838));
  AND3_X1   g413(.A1(new_n837), .A2(KEYINPUT104), .A3(new_n838), .ZN(new_n839));
  AOI21_X1  g414(.A(KEYINPUT104), .B1(new_n837), .B2(new_n838), .ZN(new_n840));
  OAI21_X1  g415(.A(new_n818), .B1(new_n839), .B2(new_n840), .ZN(new_n841));
  INV_X1    g416(.A(KEYINPUT105), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  OAI211_X1 g418(.A(KEYINPUT105), .B(new_n818), .C1(new_n839), .C2(new_n840), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n843), .A2(new_n844), .ZN(G145));
  MUX2_X1   g420(.A(G106), .B(G118), .S(G2105), .Z(new_n846));
  AOI22_X1  g421(.A1(new_n485), .A2(G130), .B1(G2104), .B2(new_n846), .ZN(new_n847));
  INV_X1    g422(.A(G142), .ZN(new_n848));
  OAI21_X1  g423(.A(new_n847), .B1(new_n848), .B2(new_n473), .ZN(new_n849));
  XNOR2_X1  g424(.A(new_n849), .B(new_n624), .ZN(new_n850));
  XNOR2_X1  g425(.A(new_n850), .B(new_n708), .ZN(new_n851));
  XOR2_X1   g426(.A(new_n851), .B(KEYINPUT108), .Z(new_n852));
  NAND2_X1  g427(.A1(new_n496), .A2(KEYINPUT4), .ZN(new_n853));
  INV_X1    g428(.A(new_n492), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n503), .A2(KEYINPUT106), .ZN(new_n856));
  INV_X1    g431(.A(KEYINPUT106), .ZN(new_n857));
  OAI211_X1 g432(.A(new_n857), .B(new_n501), .C1(new_n484), .C2(new_n502), .ZN(new_n858));
  NAND3_X1  g433(.A1(new_n855), .A2(new_n856), .A3(new_n858), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n859), .A2(KEYINPUT107), .ZN(new_n860));
  INV_X1    g435(.A(KEYINPUT107), .ZN(new_n861));
  NAND4_X1  g436(.A1(new_n855), .A2(new_n856), .A3(new_n861), .A4(new_n858), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n860), .A2(new_n862), .ZN(new_n863));
  XNOR2_X1  g438(.A(new_n863), .B(new_n801), .ZN(new_n864));
  XOR2_X1   g439(.A(new_n766), .B(new_n748), .Z(new_n865));
  XNOR2_X1  g440(.A(new_n864), .B(new_n865), .ZN(new_n866));
  INV_X1    g441(.A(new_n866), .ZN(new_n867));
  XNOR2_X1  g442(.A(new_n852), .B(new_n867), .ZN(new_n868));
  XOR2_X1   g443(.A(G160), .B(new_n489), .Z(new_n869));
  XNOR2_X1  g444(.A(new_n869), .B(new_n618), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n868), .A2(new_n870), .ZN(new_n871));
  INV_X1    g446(.A(G37), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n852), .A2(new_n867), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n866), .A2(new_n851), .ZN(new_n874));
  XOR2_X1   g449(.A(new_n870), .B(KEYINPUT109), .Z(new_n875));
  NAND3_X1  g450(.A1(new_n873), .A2(new_n874), .A3(new_n875), .ZN(new_n876));
  NAND3_X1  g451(.A1(new_n871), .A2(new_n872), .A3(new_n876), .ZN(new_n877));
  XNOR2_X1  g452(.A(new_n877), .B(KEYINPUT40), .ZN(G395));
  NOR2_X1   g453(.A1(new_n816), .A2(G868), .ZN(new_n879));
  XNOR2_X1  g454(.A(new_n823), .B(new_n610), .ZN(new_n880));
  OR2_X1    g455(.A1(new_n568), .A2(new_n598), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n568), .A2(new_n598), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n880), .A2(new_n883), .ZN(new_n884));
  XOR2_X1   g459(.A(KEYINPUT111), .B(KEYINPUT41), .Z(new_n885));
  NOR2_X1   g460(.A1(new_n883), .A2(new_n885), .ZN(new_n886));
  INV_X1    g461(.A(KEYINPUT41), .ZN(new_n887));
  INV_X1    g462(.A(KEYINPUT110), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n882), .A2(new_n888), .ZN(new_n889));
  NAND3_X1  g464(.A1(new_n568), .A2(KEYINPUT110), .A3(new_n598), .ZN(new_n890));
  NAND3_X1  g465(.A1(new_n889), .A2(new_n890), .A3(new_n881), .ZN(new_n891));
  AOI21_X1  g466(.A(new_n886), .B1(new_n887), .B2(new_n891), .ZN(new_n892));
  OAI21_X1  g467(.A(new_n884), .B1(new_n892), .B2(new_n880), .ZN(new_n893));
  XNOR2_X1  g468(.A(new_n893), .B(KEYINPUT42), .ZN(new_n894));
  XNOR2_X1  g469(.A(G305), .B(G303), .ZN(new_n895));
  XNOR2_X1  g470(.A(G290), .B(new_n573), .ZN(new_n896));
  XNOR2_X1  g471(.A(new_n895), .B(new_n896), .ZN(new_n897));
  XNOR2_X1  g472(.A(new_n894), .B(new_n897), .ZN(new_n898));
  AOI21_X1  g473(.A(new_n879), .B1(new_n898), .B2(G868), .ZN(G295));
  AOI21_X1  g474(.A(new_n879), .B1(new_n898), .B2(G868), .ZN(G331));
  INV_X1    g475(.A(KEYINPUT43), .ZN(new_n901));
  XOR2_X1   g476(.A(G301), .B(G286), .Z(new_n902));
  XNOR2_X1  g477(.A(new_n823), .B(new_n902), .ZN(new_n903));
  OR3_X1    g478(.A1(new_n903), .A2(new_n887), .A3(new_n891), .ZN(new_n904));
  OAI21_X1  g479(.A(new_n883), .B1(new_n903), .B2(new_n885), .ZN(new_n905));
  AOI21_X1  g480(.A(new_n897), .B1(new_n904), .B2(new_n905), .ZN(new_n906));
  NAND2_X1  g481(.A1(new_n903), .A2(new_n883), .ZN(new_n907));
  OAI211_X1 g482(.A(new_n907), .B(new_n897), .C1(new_n892), .C2(new_n903), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n908), .A2(new_n872), .ZN(new_n909));
  OAI21_X1  g484(.A(new_n901), .B1(new_n906), .B2(new_n909), .ZN(new_n910));
  OAI21_X1  g485(.A(new_n907), .B1(new_n892), .B2(new_n903), .ZN(new_n911));
  INV_X1    g486(.A(new_n897), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  NAND4_X1  g488(.A1(new_n913), .A2(KEYINPUT43), .A3(new_n872), .A4(new_n908), .ZN(new_n914));
  AOI21_X1  g489(.A(KEYINPUT44), .B1(new_n910), .B2(new_n914), .ZN(new_n915));
  OAI21_X1  g490(.A(KEYINPUT43), .B1(new_n906), .B2(new_n909), .ZN(new_n916));
  NAND3_X1  g491(.A1(new_n913), .A2(new_n872), .A3(new_n908), .ZN(new_n917));
  OAI21_X1  g492(.A(new_n916), .B1(new_n917), .B2(KEYINPUT43), .ZN(new_n918));
  AOI21_X1  g493(.A(new_n915), .B1(KEYINPUT44), .B2(new_n918), .ZN(G397));
  INV_X1    g494(.A(KEYINPUT45), .ZN(new_n920));
  OAI21_X1  g495(.A(new_n920), .B1(new_n863), .B2(G1384), .ZN(new_n921));
  NAND2_X1  g496(.A1(G160), .A2(G40), .ZN(new_n922));
  NOR2_X1   g497(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n708), .A2(new_n711), .ZN(new_n924));
  INV_X1    g499(.A(G2067), .ZN(new_n925));
  XNOR2_X1  g500(.A(new_n801), .B(new_n925), .ZN(new_n926));
  INV_X1    g501(.A(G1996), .ZN(new_n927));
  XNOR2_X1  g502(.A(new_n748), .B(new_n927), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n707), .A2(new_n712), .ZN(new_n929));
  NAND4_X1  g504(.A1(new_n924), .A2(new_n926), .A3(new_n928), .A4(new_n929), .ZN(new_n930));
  NAND2_X1  g505(.A1(G290), .A2(G1986), .ZN(new_n931));
  NOR2_X1   g506(.A1(new_n931), .A2(KEYINPUT112), .ZN(new_n932));
  AND2_X1   g507(.A1(new_n931), .A2(KEYINPUT112), .ZN(new_n933));
  NOR2_X1   g508(.A1(G290), .A2(G1986), .ZN(new_n934));
  INV_X1    g509(.A(new_n934), .ZN(new_n935));
  AOI21_X1  g510(.A(new_n932), .B1(new_n933), .B2(new_n935), .ZN(new_n936));
  OAI21_X1  g511(.A(new_n923), .B1(new_n930), .B2(new_n936), .ZN(new_n937));
  INV_X1    g512(.A(KEYINPUT122), .ZN(new_n938));
  AND2_X1   g513(.A1(G160), .A2(G40), .ZN(new_n939));
  XOR2_X1   g514(.A(KEYINPUT116), .B(G2084), .Z(new_n940));
  INV_X1    g515(.A(G1384), .ZN(new_n941));
  AOI21_X1  g516(.A(KEYINPUT50), .B1(new_n859), .B2(new_n941), .ZN(new_n942));
  OAI211_X1 g517(.A(KEYINPUT50), .B(new_n941), .C1(new_n497), .C2(new_n503), .ZN(new_n943));
  INV_X1    g518(.A(new_n943), .ZN(new_n944));
  OAI211_X1 g519(.A(new_n939), .B(new_n940), .C1(new_n942), .C2(new_n944), .ZN(new_n945));
  INV_X1    g520(.A(new_n945), .ZN(new_n946));
  NAND3_X1  g521(.A1(new_n859), .A2(new_n920), .A3(new_n941), .ZN(new_n947));
  OAI21_X1  g522(.A(new_n941), .B1(new_n497), .B2(new_n503), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n948), .A2(KEYINPUT45), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n947), .A2(new_n949), .ZN(new_n950));
  AOI21_X1  g525(.A(G1966), .B1(new_n950), .B2(new_n939), .ZN(new_n951));
  OAI21_X1  g526(.A(new_n938), .B1(new_n946), .B2(new_n951), .ZN(new_n952));
  AOI21_X1  g527(.A(new_n922), .B1(new_n947), .B2(new_n949), .ZN(new_n953));
  OAI211_X1 g528(.A(new_n945), .B(KEYINPUT122), .C1(G1966), .C2(new_n953), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n952), .A2(new_n954), .ZN(new_n955));
  OAI211_X1 g530(.A(KEYINPUT51), .B(G8), .C1(new_n955), .C2(G286), .ZN(new_n956));
  OAI21_X1  g531(.A(G8), .B1(new_n946), .B2(new_n951), .ZN(new_n957));
  INV_X1    g532(.A(KEYINPUT51), .ZN(new_n958));
  NAND2_X1  g533(.A1(G286), .A2(G8), .ZN(new_n959));
  NAND3_X1  g534(.A1(new_n957), .A2(new_n958), .A3(new_n959), .ZN(new_n960));
  NAND2_X1  g535(.A1(new_n956), .A2(new_n960), .ZN(new_n961));
  AOI21_X1  g536(.A(new_n959), .B1(new_n952), .B2(new_n954), .ZN(new_n962));
  INV_X1    g537(.A(new_n962), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n961), .A2(new_n963), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n964), .A2(KEYINPUT123), .ZN(new_n965));
  INV_X1    g540(.A(KEYINPUT62), .ZN(new_n966));
  INV_X1    g541(.A(KEYINPUT123), .ZN(new_n967));
  NAND3_X1  g542(.A1(new_n961), .A2(new_n967), .A3(new_n963), .ZN(new_n968));
  NAND3_X1  g543(.A1(new_n965), .A2(new_n966), .A3(new_n968), .ZN(new_n969));
  AOI21_X1  g544(.A(new_n967), .B1(new_n961), .B2(new_n963), .ZN(new_n970));
  AOI211_X1 g545(.A(KEYINPUT123), .B(new_n962), .C1(new_n956), .C2(new_n960), .ZN(new_n971));
  OAI21_X1  g546(.A(KEYINPUT62), .B1(new_n970), .B2(new_n971), .ZN(new_n972));
  INV_X1    g547(.A(KEYINPUT127), .ZN(new_n973));
  NAND3_X1  g548(.A1(new_n939), .A2(new_n941), .A3(new_n859), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n974), .A2(G8), .ZN(new_n975));
  AOI21_X1  g550(.A(new_n975), .B1(G1976), .B2(new_n684), .ZN(new_n976));
  INV_X1    g551(.A(G1976), .ZN(new_n977));
  AOI21_X1  g552(.A(KEYINPUT52), .B1(G288), .B2(new_n977), .ZN(new_n978));
  NAND2_X1  g553(.A1(new_n976), .A2(new_n978), .ZN(new_n979));
  INV_X1    g554(.A(KEYINPUT49), .ZN(new_n980));
  INV_X1    g555(.A(G1981), .ZN(new_n981));
  NAND3_X1  g556(.A1(new_n579), .A2(new_n981), .A3(new_n583), .ZN(new_n982));
  INV_X1    g557(.A(new_n982), .ZN(new_n983));
  AOI21_X1  g558(.A(new_n981), .B1(new_n579), .B2(new_n583), .ZN(new_n984));
  OAI21_X1  g559(.A(new_n980), .B1(new_n983), .B2(new_n984), .ZN(new_n985));
  INV_X1    g560(.A(new_n984), .ZN(new_n986));
  NAND3_X1  g561(.A1(new_n986), .A2(KEYINPUT49), .A3(new_n982), .ZN(new_n987));
  INV_X1    g562(.A(new_n975), .ZN(new_n988));
  NAND3_X1  g563(.A1(new_n985), .A2(new_n987), .A3(new_n988), .ZN(new_n989));
  INV_X1    g564(.A(KEYINPUT52), .ZN(new_n990));
  OAI211_X1 g565(.A(new_n979), .B(new_n989), .C1(new_n990), .C2(new_n976), .ZN(new_n991));
  NAND2_X1  g566(.A1(G303), .A2(G8), .ZN(new_n992));
  XNOR2_X1  g567(.A(KEYINPUT113), .B(KEYINPUT55), .ZN(new_n993));
  XOR2_X1   g568(.A(new_n992), .B(new_n993), .Z(new_n994));
  NAND4_X1  g569(.A1(new_n860), .A2(KEYINPUT45), .A3(new_n941), .A4(new_n862), .ZN(new_n995));
  AOI21_X1  g570(.A(new_n922), .B1(new_n920), .B2(new_n948), .ZN(new_n996));
  AOI21_X1  g571(.A(G1971), .B1(new_n995), .B2(new_n996), .ZN(new_n997));
  INV_X1    g572(.A(G2090), .ZN(new_n998));
  OAI211_X1 g573(.A(new_n998), .B(new_n939), .C1(new_n942), .C2(new_n944), .ZN(new_n999));
  INV_X1    g574(.A(new_n999), .ZN(new_n1000));
  OAI211_X1 g575(.A(new_n994), .B(G8), .C1(new_n997), .C2(new_n1000), .ZN(new_n1001));
  INV_X1    g576(.A(KEYINPUT114), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n1001), .A2(new_n1002), .ZN(new_n1003));
  OR2_X1    g578(.A1(new_n1000), .A2(new_n997), .ZN(new_n1004));
  NAND4_X1  g579(.A1(new_n1004), .A2(KEYINPUT114), .A3(G8), .A4(new_n994), .ZN(new_n1005));
  AOI21_X1  g580(.A(new_n991), .B1(new_n1003), .B2(new_n1005), .ZN(new_n1006));
  INV_X1    g581(.A(KEYINPUT53), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n995), .A2(new_n996), .ZN(new_n1008));
  OAI21_X1  g583(.A(new_n1007), .B1(new_n1008), .B2(G2078), .ZN(new_n1009));
  OAI21_X1  g584(.A(new_n939), .B1(new_n942), .B2(new_n944), .ZN(new_n1010));
  XNOR2_X1  g585(.A(KEYINPUT124), .B(G1961), .ZN(new_n1011));
  NOR2_X1   g586(.A1(new_n1007), .A2(G2078), .ZN(new_n1012));
  AOI22_X1  g587(.A1(new_n1010), .A2(new_n1011), .B1(new_n953), .B2(new_n1012), .ZN(new_n1013));
  AOI21_X1  g588(.A(G301), .B1(new_n1009), .B2(new_n1013), .ZN(new_n1014));
  INV_X1    g589(.A(KEYINPUT50), .ZN(new_n1015));
  NAND2_X1  g590(.A1(new_n948), .A2(new_n1015), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n859), .A2(new_n941), .ZN(new_n1017));
  OAI21_X1  g592(.A(new_n1016), .B1(new_n1017), .B2(new_n1015), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n1018), .A2(new_n939), .ZN(new_n1019));
  NOR2_X1   g594(.A1(new_n1019), .A2(G2090), .ZN(new_n1020));
  OAI21_X1  g595(.A(G8), .B1(new_n1020), .B2(new_n997), .ZN(new_n1021));
  INV_X1    g596(.A(new_n994), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n1021), .A2(new_n1022), .ZN(new_n1023));
  NAND3_X1  g598(.A1(new_n1006), .A2(new_n1014), .A3(new_n1023), .ZN(new_n1024));
  INV_X1    g599(.A(new_n1024), .ZN(new_n1025));
  NAND4_X1  g600(.A1(new_n969), .A2(new_n972), .A3(new_n973), .A4(new_n1025), .ZN(new_n1026));
  INV_X1    g601(.A(KEYINPUT61), .ZN(new_n1027));
  INV_X1    g602(.A(KEYINPUT119), .ZN(new_n1028));
  XOR2_X1   g603(.A(KEYINPUT117), .B(KEYINPUT57), .Z(new_n1029));
  INV_X1    g604(.A(new_n1029), .ZN(new_n1030));
  NAND2_X1  g605(.A1(new_n561), .A2(new_n562), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n559), .A2(KEYINPUT9), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n1031), .A2(new_n1032), .ZN(new_n1033));
  AOI21_X1  g608(.A(new_n1030), .B1(new_n1033), .B2(new_n566), .ZN(new_n1034));
  NOR3_X1   g609(.A1(new_n563), .A2(new_n567), .A3(new_n1029), .ZN(new_n1035));
  OAI21_X1  g610(.A(new_n1028), .B1(new_n1034), .B2(new_n1035), .ZN(new_n1036));
  NAND3_X1  g611(.A1(new_n1033), .A2(new_n566), .A3(new_n1030), .ZN(new_n1037));
  OAI21_X1  g612(.A(new_n1029), .B1(new_n563), .B2(new_n567), .ZN(new_n1038));
  NAND3_X1  g613(.A1(new_n1037), .A2(new_n1038), .A3(KEYINPUT119), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n1036), .A2(new_n1039), .ZN(new_n1040));
  XNOR2_X1  g615(.A(KEYINPUT56), .B(G2072), .ZN(new_n1041));
  NAND3_X1  g616(.A1(new_n995), .A2(new_n996), .A3(new_n1041), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n1042), .A2(KEYINPUT118), .ZN(new_n1043));
  INV_X1    g618(.A(KEYINPUT118), .ZN(new_n1044));
  NAND4_X1  g619(.A1(new_n995), .A2(new_n1044), .A3(new_n996), .A4(new_n1041), .ZN(new_n1045));
  INV_X1    g620(.A(G1956), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n1019), .A2(new_n1046), .ZN(new_n1047));
  NAND3_X1  g622(.A1(new_n1043), .A2(new_n1045), .A3(new_n1047), .ZN(new_n1048));
  AOI21_X1  g623(.A(new_n1027), .B1(new_n1040), .B2(new_n1048), .ZN(new_n1049));
  AND2_X1   g624(.A1(new_n1047), .A2(new_n1045), .ZN(new_n1050));
  NOR2_X1   g625(.A1(new_n1034), .A2(new_n1035), .ZN(new_n1051));
  NAND3_X1  g626(.A1(new_n1050), .A2(new_n1043), .A3(new_n1051), .ZN(new_n1052));
  AND3_X1   g627(.A1(new_n1049), .A2(KEYINPUT120), .A3(new_n1052), .ZN(new_n1053));
  AOI21_X1  g628(.A(KEYINPUT120), .B1(new_n1049), .B2(new_n1052), .ZN(new_n1054));
  NOR2_X1   g629(.A1(new_n1053), .A2(new_n1054), .ZN(new_n1055));
  NOR2_X1   g630(.A1(new_n1017), .A2(new_n922), .ZN(new_n1056));
  AOI22_X1  g631(.A1(new_n1010), .A2(new_n796), .B1(new_n925), .B2(new_n1056), .ZN(new_n1057));
  NOR2_X1   g632(.A1(new_n826), .A2(new_n1057), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n1010), .A2(new_n796), .ZN(new_n1059));
  OAI21_X1  g634(.A(new_n1059), .B1(G2067), .B2(new_n974), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n1060), .A2(KEYINPUT60), .ZN(new_n1061));
  AOI21_X1  g636(.A(new_n1058), .B1(new_n1061), .B2(new_n826), .ZN(new_n1062));
  XOR2_X1   g637(.A(KEYINPUT121), .B(KEYINPUT60), .Z(new_n1063));
  INV_X1    g638(.A(new_n1063), .ZN(new_n1064));
  XNOR2_X1  g639(.A(KEYINPUT58), .B(G1341), .ZN(new_n1065));
  OAI22_X1  g640(.A1(new_n1008), .A2(G1996), .B1(new_n1056), .B2(new_n1065), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n1066), .A2(new_n551), .ZN(new_n1067));
  NAND2_X1  g642(.A1(new_n1067), .A2(KEYINPUT59), .ZN(new_n1068));
  INV_X1    g643(.A(KEYINPUT59), .ZN(new_n1069));
  NAND3_X1  g644(.A1(new_n1066), .A2(new_n1069), .A3(new_n551), .ZN(new_n1070));
  AOI22_X1  g645(.A1(new_n1062), .A2(new_n1064), .B1(new_n1068), .B2(new_n1070), .ZN(new_n1071));
  NOR3_X1   g646(.A1(new_n1048), .A2(new_n1035), .A3(new_n1034), .ZN(new_n1072));
  AOI21_X1  g647(.A(new_n1051), .B1(new_n1050), .B2(new_n1043), .ZN(new_n1073));
  OAI21_X1  g648(.A(new_n1027), .B1(new_n1072), .B2(new_n1073), .ZN(new_n1074));
  AOI21_X1  g649(.A(new_n599), .B1(new_n1060), .B2(KEYINPUT60), .ZN(new_n1075));
  OAI21_X1  g650(.A(new_n1063), .B1(new_n1075), .B2(new_n1058), .ZN(new_n1076));
  NAND3_X1  g651(.A1(new_n1071), .A2(new_n1074), .A3(new_n1076), .ZN(new_n1077));
  AOI21_X1  g652(.A(new_n1058), .B1(new_n1040), .B2(new_n1048), .ZN(new_n1078));
  OAI22_X1  g653(.A1(new_n1055), .A2(new_n1077), .B1(new_n1078), .B2(new_n1072), .ZN(new_n1079));
  INV_X1    g654(.A(KEYINPUT54), .ZN(new_n1080));
  NAND4_X1  g655(.A1(new_n921), .A2(new_n939), .A3(new_n995), .A4(new_n1012), .ZN(new_n1081));
  NAND2_X1  g656(.A1(new_n1010), .A2(new_n1011), .ZN(new_n1082));
  NAND3_X1  g657(.A1(new_n1009), .A2(new_n1081), .A3(new_n1082), .ZN(new_n1083));
  NOR2_X1   g658(.A1(new_n1083), .A2(G171), .ZN(new_n1084));
  OAI21_X1  g659(.A(new_n1080), .B1(new_n1084), .B2(new_n1014), .ZN(new_n1085));
  NAND3_X1  g660(.A1(new_n1006), .A2(new_n1023), .A3(new_n1085), .ZN(new_n1086));
  AND2_X1   g661(.A1(new_n1009), .A2(new_n1013), .ZN(new_n1087));
  AOI21_X1  g662(.A(new_n1080), .B1(new_n1087), .B2(G301), .ZN(new_n1088));
  INV_X1    g663(.A(KEYINPUT125), .ZN(new_n1089));
  AND3_X1   g664(.A1(new_n1083), .A2(new_n1089), .A3(G171), .ZN(new_n1090));
  AOI21_X1  g665(.A(new_n1089), .B1(new_n1083), .B2(G171), .ZN(new_n1091));
  OAI21_X1  g666(.A(new_n1088), .B1(new_n1090), .B2(new_n1091), .ZN(new_n1092));
  NAND2_X1  g667(.A1(new_n1092), .A2(KEYINPUT126), .ZN(new_n1093));
  INV_X1    g668(.A(KEYINPUT126), .ZN(new_n1094));
  OAI211_X1 g669(.A(new_n1094), .B(new_n1088), .C1(new_n1090), .C2(new_n1091), .ZN(new_n1095));
  AOI21_X1  g670(.A(new_n1086), .B1(new_n1093), .B2(new_n1095), .ZN(new_n1096));
  NAND2_X1  g671(.A1(new_n965), .A2(new_n968), .ZN(new_n1097));
  NAND3_X1  g672(.A1(new_n1079), .A2(new_n1096), .A3(new_n1097), .ZN(new_n1098));
  XNOR2_X1  g673(.A(new_n975), .B(KEYINPUT115), .ZN(new_n1099));
  NOR2_X1   g674(.A1(G288), .A2(G1976), .ZN(new_n1100));
  AND2_X1   g675(.A1(new_n989), .A2(new_n1100), .ZN(new_n1101));
  OAI21_X1  g676(.A(new_n1099), .B1(new_n1101), .B2(new_n983), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n1003), .A2(new_n1005), .ZN(new_n1103));
  OAI21_X1  g678(.A(new_n1102), .B1(new_n1103), .B2(new_n991), .ZN(new_n1104));
  INV_X1    g679(.A(KEYINPUT63), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n1006), .A2(new_n1023), .ZN(new_n1106));
  OR2_X1    g681(.A1(new_n957), .A2(G286), .ZN(new_n1107));
  OAI21_X1  g682(.A(new_n1105), .B1(new_n1106), .B2(new_n1107), .ZN(new_n1108));
  AOI21_X1  g683(.A(new_n994), .B1(new_n1004), .B2(G8), .ZN(new_n1109));
  NOR3_X1   g684(.A1(new_n1109), .A2(new_n1107), .A3(new_n1105), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n1006), .A2(new_n1110), .ZN(new_n1111));
  AOI21_X1  g686(.A(new_n1104), .B1(new_n1108), .B2(new_n1111), .ZN(new_n1112));
  NAND3_X1  g687(.A1(new_n1026), .A2(new_n1098), .A3(new_n1112), .ZN(new_n1113));
  NOR2_X1   g688(.A1(new_n970), .A2(new_n971), .ZN(new_n1114));
  AOI21_X1  g689(.A(new_n1024), .B1(new_n1114), .B2(new_n966), .ZN(new_n1115));
  AOI21_X1  g690(.A(new_n973), .B1(new_n1115), .B2(new_n972), .ZN(new_n1116));
  OAI21_X1  g691(.A(new_n937), .B1(new_n1113), .B2(new_n1116), .ZN(new_n1117));
  AOI21_X1  g692(.A(KEYINPUT48), .B1(new_n923), .B2(new_n934), .ZN(new_n1118));
  AND3_X1   g693(.A1(new_n923), .A2(KEYINPUT48), .A3(new_n934), .ZN(new_n1119));
  AOI211_X1 g694(.A(new_n1118), .B(new_n1119), .C1(new_n923), .C2(new_n930), .ZN(new_n1120));
  INV_X1    g695(.A(new_n926), .ZN(new_n1121));
  OAI21_X1  g696(.A(new_n923), .B1(new_n748), .B2(new_n1121), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n923), .A2(new_n927), .ZN(new_n1123));
  AND2_X1   g698(.A1(new_n1123), .A2(KEYINPUT46), .ZN(new_n1124));
  NOR2_X1   g699(.A1(new_n1123), .A2(KEYINPUT46), .ZN(new_n1125));
  OAI21_X1  g700(.A(new_n1122), .B1(new_n1124), .B2(new_n1125), .ZN(new_n1126));
  XOR2_X1   g701(.A(new_n1126), .B(KEYINPUT47), .Z(new_n1127));
  NAND2_X1  g702(.A1(new_n926), .A2(new_n928), .ZN(new_n1128));
  OAI22_X1  g703(.A1(new_n1128), .A2(new_n924), .B1(G2067), .B2(new_n801), .ZN(new_n1129));
  AOI211_X1 g704(.A(new_n1120), .B(new_n1127), .C1(new_n923), .C2(new_n1129), .ZN(new_n1130));
  NAND2_X1  g705(.A1(new_n1117), .A2(new_n1130), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g706(.A(G227), .ZN(new_n1133));
  NAND3_X1  g707(.A1(new_n677), .A2(G319), .A3(new_n1133), .ZN(new_n1134));
  NOR2_X1   g708(.A1(G401), .A2(new_n1134), .ZN(new_n1135));
  NAND4_X1  g709(.A1(new_n910), .A2(new_n877), .A3(new_n914), .A4(new_n1135), .ZN(G225));
  INV_X1    g710(.A(G225), .ZN(G308));
endmodule


