//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 0 1 1 0 0 1 0 0 1 1 0 0 1 1 0 1 1 0 0 1 1 0 1 1 0 1 0 1 0 0 0 0 1 1 0 1 1 1 0 0 1 0 1 1 0 0 0 0 1 1 1 0 1 0 1 1 0 0 1 1 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:22:43 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n727, new_n728, new_n729, new_n730, new_n731,
    new_n732, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n741, new_n743, new_n744, new_n745, new_n746, new_n747, new_n749,
    new_n750, new_n751, new_n752, new_n753, new_n754, new_n755, new_n756,
    new_n757, new_n759, new_n760, new_n761, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n791, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n820, new_n821, new_n822, new_n823, new_n824,
    new_n825, new_n826, new_n827, new_n828, new_n829, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n925, new_n926, new_n927, new_n928, new_n929, new_n930, new_n931,
    new_n932, new_n933, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n948, new_n949, new_n950, new_n951, new_n953, new_n954, new_n955,
    new_n956, new_n957, new_n958, new_n959, new_n960, new_n961, new_n962,
    new_n963, new_n964, new_n965, new_n966, new_n968, new_n969, new_n970,
    new_n971, new_n972, new_n973, new_n975, new_n976, new_n977, new_n978,
    new_n979, new_n980, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1021;
  INV_X1    g000(.A(G217), .ZN(new_n187));
  INV_X1    g001(.A(G902), .ZN(new_n188));
  AOI21_X1  g002(.A(new_n187), .B1(G234), .B2(new_n188), .ZN(new_n189));
  INV_X1    g003(.A(new_n189), .ZN(new_n190));
  INV_X1    g004(.A(KEYINPUT67), .ZN(new_n191));
  INV_X1    g005(.A(G119), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n191), .A2(new_n192), .ZN(new_n193));
  NAND2_X1  g007(.A1(KEYINPUT67), .A2(G119), .ZN(new_n194));
  NAND3_X1  g008(.A1(new_n193), .A2(G128), .A3(new_n194), .ZN(new_n195));
  NOR2_X1   g009(.A1(new_n192), .A2(G128), .ZN(new_n196));
  INV_X1    g010(.A(new_n196), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n195), .A2(new_n197), .ZN(new_n198));
  XNOR2_X1  g012(.A(KEYINPUT24), .B(G110), .ZN(new_n199));
  NOR2_X1   g013(.A1(new_n198), .A2(new_n199), .ZN(new_n200));
  INV_X1    g014(.A(G140), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n201), .A2(G125), .ZN(new_n202));
  INV_X1    g016(.A(G125), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n203), .A2(G140), .ZN(new_n204));
  NAND3_X1  g018(.A1(new_n202), .A2(new_n204), .A3(KEYINPUT75), .ZN(new_n205));
  OR3_X1    g019(.A1(new_n203), .A2(KEYINPUT75), .A3(G140), .ZN(new_n206));
  NAND3_X1  g020(.A1(new_n205), .A2(new_n206), .A3(KEYINPUT16), .ZN(new_n207));
  INV_X1    g021(.A(KEYINPUT16), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n202), .A2(new_n208), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n207), .A2(new_n209), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n210), .A2(G146), .ZN(new_n211));
  INV_X1    g025(.A(G146), .ZN(new_n212));
  NAND3_X1  g026(.A1(new_n207), .A2(new_n212), .A3(new_n209), .ZN(new_n213));
  AOI21_X1  g027(.A(new_n200), .B1(new_n211), .B2(new_n213), .ZN(new_n214));
  INV_X1    g028(.A(KEYINPUT74), .ZN(new_n215));
  INV_X1    g029(.A(G128), .ZN(new_n216));
  AND2_X1   g030(.A1(KEYINPUT67), .A2(G119), .ZN(new_n217));
  NOR2_X1   g031(.A1(KEYINPUT67), .A2(G119), .ZN(new_n218));
  OAI21_X1  g032(.A(new_n216), .B1(new_n217), .B2(new_n218), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n219), .A2(KEYINPUT73), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n195), .A2(KEYINPUT23), .ZN(new_n221));
  INV_X1    g035(.A(KEYINPUT73), .ZN(new_n222));
  OAI211_X1 g036(.A(new_n222), .B(new_n216), .C1(new_n217), .C2(new_n218), .ZN(new_n223));
  NAND3_X1  g037(.A1(new_n220), .A2(new_n221), .A3(new_n223), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n196), .A2(KEYINPUT23), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  AOI21_X1  g040(.A(new_n215), .B1(new_n226), .B2(G110), .ZN(new_n227));
  INV_X1    g041(.A(G110), .ZN(new_n228));
  AOI211_X1 g042(.A(KEYINPUT74), .B(new_n228), .C1(new_n224), .C2(new_n225), .ZN(new_n229));
  OAI21_X1  g043(.A(new_n214), .B1(new_n227), .B2(new_n229), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n198), .A2(new_n199), .ZN(new_n231));
  OAI21_X1  g045(.A(new_n231), .B1(new_n226), .B2(G110), .ZN(new_n232));
  XNOR2_X1  g046(.A(G125), .B(G140), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n233), .A2(new_n212), .ZN(new_n234));
  INV_X1    g048(.A(KEYINPUT76), .ZN(new_n235));
  XNOR2_X1  g049(.A(new_n234), .B(new_n235), .ZN(new_n236));
  AND2_X1   g050(.A1(new_n211), .A2(new_n236), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n232), .A2(new_n237), .ZN(new_n238));
  INV_X1    g052(.A(G953), .ZN(new_n239));
  NAND3_X1  g053(.A1(new_n239), .A2(G221), .A3(G234), .ZN(new_n240));
  XNOR2_X1  g054(.A(new_n240), .B(KEYINPUT77), .ZN(new_n241));
  XNOR2_X1  g055(.A(KEYINPUT22), .B(G137), .ZN(new_n242));
  XNOR2_X1  g056(.A(new_n241), .B(new_n242), .ZN(new_n243));
  AND3_X1   g057(.A1(new_n230), .A2(new_n238), .A3(new_n243), .ZN(new_n244));
  AOI21_X1  g058(.A(new_n243), .B1(new_n230), .B2(new_n238), .ZN(new_n245));
  OAI21_X1  g059(.A(new_n188), .B1(new_n244), .B2(new_n245), .ZN(new_n246));
  INV_X1    g060(.A(KEYINPUT25), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n246), .A2(new_n247), .ZN(new_n248));
  INV_X1    g062(.A(new_n243), .ZN(new_n249));
  INV_X1    g063(.A(new_n213), .ZN(new_n250));
  AOI21_X1  g064(.A(new_n212), .B1(new_n207), .B2(new_n209), .ZN(new_n251));
  OAI22_X1  g065(.A1(new_n250), .A2(new_n251), .B1(new_n198), .B2(new_n199), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n226), .A2(G110), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n253), .A2(KEYINPUT74), .ZN(new_n254));
  NAND3_X1  g068(.A1(new_n226), .A2(new_n215), .A3(G110), .ZN(new_n255));
  AOI21_X1  g069(.A(new_n252), .B1(new_n254), .B2(new_n255), .ZN(new_n256));
  AND2_X1   g070(.A1(new_n232), .A2(new_n237), .ZN(new_n257));
  OAI21_X1  g071(.A(new_n249), .B1(new_n256), .B2(new_n257), .ZN(new_n258));
  NAND3_X1  g072(.A1(new_n230), .A2(new_n238), .A3(new_n243), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  NAND3_X1  g074(.A1(new_n260), .A2(KEYINPUT25), .A3(new_n188), .ZN(new_n261));
  AOI21_X1  g075(.A(new_n190), .B1(new_n248), .B2(new_n261), .ZN(new_n262));
  NOR2_X1   g076(.A1(new_n189), .A2(G902), .ZN(new_n263));
  AND2_X1   g077(.A1(new_n260), .A2(new_n263), .ZN(new_n264));
  NOR2_X1   g078(.A1(new_n262), .A2(new_n264), .ZN(new_n265));
  INV_X1    g079(.A(new_n265), .ZN(new_n266));
  INV_X1    g080(.A(G134), .ZN(new_n267));
  OAI21_X1  g081(.A(KEYINPUT11), .B1(new_n267), .B2(G137), .ZN(new_n268));
  INV_X1    g082(.A(KEYINPUT11), .ZN(new_n269));
  INV_X1    g083(.A(G137), .ZN(new_n270));
  NAND3_X1  g084(.A1(new_n269), .A2(new_n270), .A3(G134), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n268), .A2(new_n271), .ZN(new_n272));
  INV_X1    g086(.A(G131), .ZN(new_n273));
  OAI21_X1  g087(.A(KEYINPUT66), .B1(new_n270), .B2(G134), .ZN(new_n274));
  INV_X1    g088(.A(KEYINPUT66), .ZN(new_n275));
  NAND3_X1  g089(.A1(new_n275), .A2(new_n267), .A3(G137), .ZN(new_n276));
  NAND4_X1  g090(.A1(new_n272), .A2(new_n273), .A3(new_n274), .A4(new_n276), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n212), .A2(G143), .ZN(new_n278));
  INV_X1    g092(.A(G143), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n279), .A2(G146), .ZN(new_n280));
  OAI211_X1 g094(.A(new_n278), .B(new_n280), .C1(KEYINPUT1), .C2(new_n216), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n278), .A2(new_n280), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n278), .A2(KEYINPUT1), .ZN(new_n283));
  NAND3_X1  g097(.A1(new_n282), .A2(new_n283), .A3(G128), .ZN(new_n284));
  NOR2_X1   g098(.A1(new_n267), .A2(G137), .ZN(new_n285));
  NOR2_X1   g099(.A1(new_n270), .A2(G134), .ZN(new_n286));
  OAI21_X1  g100(.A(G131), .B1(new_n285), .B2(new_n286), .ZN(new_n287));
  NAND4_X1  g101(.A1(new_n277), .A2(new_n281), .A3(new_n284), .A4(new_n287), .ZN(new_n288));
  NAND3_X1  g102(.A1(new_n193), .A2(G116), .A3(new_n194), .ZN(new_n289));
  INV_X1    g103(.A(G116), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n290), .A2(G119), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n289), .A2(new_n291), .ZN(new_n292));
  XNOR2_X1  g106(.A(KEYINPUT2), .B(G113), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  INV_X1    g108(.A(new_n293), .ZN(new_n295));
  NAND3_X1  g109(.A1(new_n295), .A2(new_n289), .A3(new_n291), .ZN(new_n296));
  AND2_X1   g110(.A1(new_n294), .A2(new_n296), .ZN(new_n297));
  AND2_X1   g111(.A1(new_n268), .A2(new_n271), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n274), .A2(new_n276), .ZN(new_n299));
  OAI21_X1  g113(.A(G131), .B1(new_n298), .B2(new_n299), .ZN(new_n300));
  AND2_X1   g114(.A1(new_n300), .A2(new_n277), .ZN(new_n301));
  NAND4_X1  g115(.A1(new_n278), .A2(new_n280), .A3(KEYINPUT0), .A4(G128), .ZN(new_n302));
  NOR2_X1   g116(.A1(KEYINPUT0), .A2(G128), .ZN(new_n303));
  AOI21_X1  g117(.A(new_n303), .B1(new_n278), .B2(new_n280), .ZN(new_n304));
  AND3_X1   g118(.A1(KEYINPUT64), .A2(KEYINPUT0), .A3(G128), .ZN(new_n305));
  AOI21_X1  g119(.A(KEYINPUT64), .B1(KEYINPUT0), .B2(G128), .ZN(new_n306));
  NOR2_X1   g120(.A1(new_n305), .A2(new_n306), .ZN(new_n307));
  AND3_X1   g121(.A1(new_n304), .A2(KEYINPUT65), .A3(new_n307), .ZN(new_n308));
  AOI21_X1  g122(.A(KEYINPUT65), .B1(new_n304), .B2(new_n307), .ZN(new_n309));
  OAI21_X1  g123(.A(new_n302), .B1(new_n308), .B2(new_n309), .ZN(new_n310));
  OAI211_X1 g124(.A(new_n288), .B(new_n297), .C1(new_n301), .C2(new_n310), .ZN(new_n311));
  XNOR2_X1  g125(.A(KEYINPUT26), .B(G101), .ZN(new_n312));
  XNOR2_X1  g126(.A(KEYINPUT68), .B(KEYINPUT27), .ZN(new_n313));
  XNOR2_X1  g127(.A(new_n312), .B(new_n313), .ZN(new_n314));
  NOR2_X1   g128(.A1(G237), .A2(G953), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n315), .A2(G210), .ZN(new_n316));
  XNOR2_X1  g130(.A(new_n316), .B(KEYINPUT69), .ZN(new_n317));
  AND2_X1   g131(.A1(new_n314), .A2(new_n317), .ZN(new_n318));
  NOR2_X1   g132(.A1(new_n314), .A2(new_n317), .ZN(new_n319));
  NOR2_X1   g133(.A1(new_n318), .A2(new_n319), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n311), .A2(new_n320), .ZN(new_n321));
  OAI21_X1  g135(.A(new_n288), .B1(new_n301), .B2(new_n310), .ZN(new_n322));
  INV_X1    g136(.A(KEYINPUT30), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  AND2_X1   g138(.A1(new_n288), .A2(KEYINPUT30), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n300), .A2(new_n277), .ZN(new_n326));
  INV_X1    g140(.A(KEYINPUT65), .ZN(new_n327));
  INV_X1    g141(.A(new_n303), .ZN(new_n328));
  NOR2_X1   g142(.A1(new_n279), .A2(G146), .ZN(new_n329));
  NOR2_X1   g143(.A1(new_n212), .A2(G143), .ZN(new_n330));
  OAI21_X1  g144(.A(new_n328), .B1(new_n329), .B2(new_n330), .ZN(new_n331));
  INV_X1    g145(.A(new_n306), .ZN(new_n332));
  NAND3_X1  g146(.A1(KEYINPUT64), .A2(KEYINPUT0), .A3(G128), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  OAI21_X1  g148(.A(new_n327), .B1(new_n331), .B2(new_n334), .ZN(new_n335));
  NAND3_X1  g149(.A1(new_n304), .A2(new_n307), .A3(KEYINPUT65), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n335), .A2(new_n336), .ZN(new_n337));
  NAND3_X1  g151(.A1(new_n326), .A2(new_n337), .A3(new_n302), .ZN(new_n338));
  AOI21_X1  g152(.A(new_n297), .B1(new_n325), .B2(new_n338), .ZN(new_n339));
  AOI21_X1  g153(.A(new_n321), .B1(new_n324), .B2(new_n339), .ZN(new_n340));
  INV_X1    g154(.A(KEYINPUT31), .ZN(new_n341));
  OAI21_X1  g155(.A(KEYINPUT70), .B1(new_n340), .B2(new_n341), .ZN(new_n342));
  XNOR2_X1  g156(.A(new_n314), .B(new_n317), .ZN(new_n343));
  INV_X1    g157(.A(KEYINPUT28), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n294), .A2(new_n296), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n322), .A2(new_n345), .ZN(new_n346));
  AOI21_X1  g160(.A(new_n344), .B1(new_n346), .B2(new_n311), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n311), .A2(new_n344), .ZN(new_n348));
  INV_X1    g162(.A(new_n348), .ZN(new_n349));
  OAI21_X1  g163(.A(new_n343), .B1(new_n347), .B2(new_n349), .ZN(new_n350));
  INV_X1    g164(.A(new_n302), .ZN(new_n351));
  AOI21_X1  g165(.A(new_n351), .B1(new_n335), .B2(new_n336), .ZN(new_n352));
  AND2_X1   g166(.A1(new_n277), .A2(new_n287), .ZN(new_n353));
  AND2_X1   g167(.A1(new_n284), .A2(new_n281), .ZN(new_n354));
  AOI22_X1  g168(.A1(new_n352), .A2(new_n326), .B1(new_n353), .B2(new_n354), .ZN(new_n355));
  AOI21_X1  g169(.A(new_n343), .B1(new_n355), .B2(new_n297), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n325), .A2(new_n338), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n357), .A2(new_n345), .ZN(new_n358));
  NOR2_X1   g172(.A1(new_n355), .A2(KEYINPUT30), .ZN(new_n359));
  OAI21_X1  g173(.A(new_n356), .B1(new_n358), .B2(new_n359), .ZN(new_n360));
  INV_X1    g174(.A(KEYINPUT70), .ZN(new_n361));
  NAND3_X1  g175(.A1(new_n360), .A2(new_n361), .A3(KEYINPUT31), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n340), .A2(new_n341), .ZN(new_n363));
  NAND4_X1  g177(.A1(new_n342), .A2(new_n350), .A3(new_n362), .A4(new_n363), .ZN(new_n364));
  NOR2_X1   g178(.A1(G472), .A2(G902), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  INV_X1    g180(.A(KEYINPUT71), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n366), .A2(new_n367), .ZN(new_n368));
  INV_X1    g182(.A(KEYINPUT32), .ZN(new_n369));
  NAND3_X1  g183(.A1(new_n364), .A2(KEYINPUT71), .A3(new_n365), .ZN(new_n370));
  NAND3_X1  g184(.A1(new_n368), .A2(new_n369), .A3(new_n370), .ZN(new_n371));
  AND2_X1   g185(.A1(new_n364), .A2(new_n365), .ZN(new_n372));
  NOR3_X1   g186(.A1(new_n347), .A2(new_n349), .A3(new_n343), .ZN(new_n373));
  INV_X1    g187(.A(KEYINPUT29), .ZN(new_n374));
  AOI22_X1  g188(.A1(new_n324), .A2(new_n339), .B1(new_n355), .B2(new_n297), .ZN(new_n375));
  OAI21_X1  g189(.A(new_n374), .B1(new_n375), .B2(new_n320), .ZN(new_n376));
  OAI21_X1  g190(.A(KEYINPUT72), .B1(new_n373), .B2(new_n376), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n346), .A2(new_n311), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n378), .A2(KEYINPUT28), .ZN(new_n379));
  NAND3_X1  g193(.A1(new_n379), .A2(new_n348), .A3(new_n320), .ZN(new_n380));
  OAI21_X1  g194(.A(new_n311), .B1(new_n358), .B2(new_n359), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n381), .A2(new_n343), .ZN(new_n382));
  INV_X1    g196(.A(KEYINPUT72), .ZN(new_n383));
  NAND4_X1  g197(.A1(new_n380), .A2(new_n382), .A3(new_n383), .A4(new_n374), .ZN(new_n384));
  AOI21_X1  g198(.A(G902), .B1(new_n373), .B2(KEYINPUT29), .ZN(new_n385));
  NAND3_X1  g199(.A1(new_n377), .A2(new_n384), .A3(new_n385), .ZN(new_n386));
  AOI22_X1  g200(.A1(new_n372), .A2(KEYINPUT32), .B1(new_n386), .B2(G472), .ZN(new_n387));
  AOI21_X1  g201(.A(new_n266), .B1(new_n371), .B2(new_n387), .ZN(new_n388));
  XNOR2_X1  g202(.A(G113), .B(G122), .ZN(new_n389));
  INV_X1    g203(.A(G104), .ZN(new_n390));
  XNOR2_X1  g204(.A(new_n389), .B(new_n390), .ZN(new_n391));
  NAND3_X1  g205(.A1(new_n205), .A2(new_n206), .A3(G146), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n236), .A2(new_n392), .ZN(new_n393));
  OR2_X1    g207(.A1(KEYINPUT89), .A2(G143), .ZN(new_n394));
  NAND2_X1  g208(.A1(KEYINPUT89), .A2(G143), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n394), .A2(new_n395), .ZN(new_n396));
  NAND3_X1  g210(.A1(new_n396), .A2(G214), .A3(new_n315), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n315), .A2(G214), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n398), .A2(new_n395), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n397), .A2(new_n399), .ZN(new_n400));
  NAND3_X1  g214(.A1(new_n400), .A2(KEYINPUT18), .A3(G131), .ZN(new_n401));
  NAND2_X1  g215(.A1(KEYINPUT18), .A2(G131), .ZN(new_n402));
  NAND3_X1  g216(.A1(new_n397), .A2(new_n399), .A3(new_n402), .ZN(new_n403));
  NAND3_X1  g217(.A1(new_n393), .A2(new_n401), .A3(new_n403), .ZN(new_n404));
  NOR2_X1   g218(.A1(new_n250), .A2(new_n251), .ZN(new_n405));
  AOI21_X1  g219(.A(new_n398), .B1(new_n394), .B2(new_n395), .ZN(new_n406));
  AND2_X1   g220(.A1(new_n398), .A2(new_n395), .ZN(new_n407));
  OAI211_X1 g221(.A(KEYINPUT17), .B(G131), .C1(new_n406), .C2(new_n407), .ZN(new_n408));
  AOI21_X1  g222(.A(KEYINPUT90), .B1(new_n405), .B2(new_n408), .ZN(new_n409));
  NAND4_X1  g223(.A1(new_n211), .A2(KEYINPUT90), .A3(new_n213), .A4(new_n408), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n400), .A2(G131), .ZN(new_n411));
  INV_X1    g225(.A(KEYINPUT17), .ZN(new_n412));
  NAND3_X1  g226(.A1(new_n397), .A2(new_n273), .A3(new_n399), .ZN(new_n413));
  NAND3_X1  g227(.A1(new_n411), .A2(new_n412), .A3(new_n413), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n410), .A2(new_n414), .ZN(new_n415));
  OAI211_X1 g229(.A(new_n391), .B(new_n404), .C1(new_n409), .C2(new_n415), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n411), .A2(new_n413), .ZN(new_n417));
  INV_X1    g231(.A(KEYINPUT19), .ZN(new_n418));
  AOI21_X1  g232(.A(new_n418), .B1(new_n205), .B2(new_n206), .ZN(new_n419));
  NOR2_X1   g233(.A1(new_n233), .A2(KEYINPUT19), .ZN(new_n420));
  NOR2_X1   g234(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  OAI211_X1 g235(.A(new_n417), .B(new_n211), .C1(G146), .C2(new_n421), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n422), .A2(new_n404), .ZN(new_n423));
  INV_X1    g237(.A(new_n391), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n423), .A2(new_n424), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n416), .A2(new_n425), .ZN(new_n426));
  NOR2_X1   g240(.A1(G475), .A2(G902), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n426), .A2(new_n427), .ZN(new_n428));
  NAND3_X1  g242(.A1(new_n428), .A2(KEYINPUT91), .A3(KEYINPUT20), .ZN(new_n429));
  INV_X1    g243(.A(KEYINPUT91), .ZN(new_n430));
  INV_X1    g244(.A(new_n427), .ZN(new_n431));
  AOI21_X1  g245(.A(new_n431), .B1(new_n416), .B2(new_n425), .ZN(new_n432));
  INV_X1    g246(.A(KEYINPUT20), .ZN(new_n433));
  OAI21_X1  g247(.A(new_n430), .B1(new_n432), .B2(new_n433), .ZN(new_n434));
  INV_X1    g248(.A(KEYINPUT92), .ZN(new_n435));
  AOI21_X1  g249(.A(KEYINPUT20), .B1(new_n431), .B2(new_n435), .ZN(new_n436));
  OAI211_X1 g250(.A(new_n426), .B(new_n436), .C1(new_n435), .C2(new_n431), .ZN(new_n437));
  NAND3_X1  g251(.A1(new_n429), .A2(new_n434), .A3(new_n437), .ZN(new_n438));
  OAI21_X1  g252(.A(new_n404), .B1(new_n409), .B2(new_n415), .ZN(new_n439));
  AND2_X1   g253(.A1(new_n439), .A2(new_n424), .ZN(new_n440));
  INV_X1    g254(.A(new_n416), .ZN(new_n441));
  OAI21_X1  g255(.A(new_n188), .B1(new_n440), .B2(new_n441), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n442), .A2(G475), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n438), .A2(new_n443), .ZN(new_n444));
  INV_X1    g258(.A(G478), .ZN(new_n445));
  NOR2_X1   g259(.A1(new_n445), .A2(KEYINPUT15), .ZN(new_n446));
  INV_X1    g260(.A(new_n446), .ZN(new_n447));
  OR2_X1    g261(.A1(KEYINPUT78), .A2(G107), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n290), .A2(G122), .ZN(new_n449));
  INV_X1    g263(.A(G122), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n450), .A2(G116), .ZN(new_n451));
  NAND2_X1  g265(.A1(KEYINPUT78), .A2(G107), .ZN(new_n452));
  AND4_X1   g266(.A1(new_n448), .A2(new_n449), .A3(new_n451), .A4(new_n452), .ZN(new_n453));
  INV_X1    g267(.A(KEYINPUT14), .ZN(new_n454));
  NOR2_X1   g268(.A1(new_n449), .A2(new_n454), .ZN(new_n455));
  INV_X1    g269(.A(G107), .ZN(new_n456));
  NOR2_X1   g270(.A1(new_n455), .A2(new_n456), .ZN(new_n457));
  XNOR2_X1  g271(.A(G116), .B(G122), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n458), .A2(new_n454), .ZN(new_n459));
  AOI21_X1  g273(.A(new_n453), .B1(new_n457), .B2(new_n459), .ZN(new_n460));
  OAI21_X1  g274(.A(KEYINPUT93), .B1(new_n216), .B2(G143), .ZN(new_n461));
  INV_X1    g275(.A(KEYINPUT93), .ZN(new_n462));
  NAND3_X1  g276(.A1(new_n462), .A2(new_n279), .A3(G128), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n461), .A2(new_n463), .ZN(new_n464));
  NOR2_X1   g278(.A1(new_n279), .A2(G128), .ZN(new_n465));
  INV_X1    g279(.A(new_n465), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n464), .A2(new_n466), .ZN(new_n467));
  NOR2_X1   g281(.A1(new_n467), .A2(G134), .ZN(new_n468));
  AOI21_X1  g282(.A(new_n267), .B1(new_n464), .B2(new_n466), .ZN(new_n469));
  OAI21_X1  g283(.A(new_n460), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  INV_X1    g284(.A(KEYINPUT95), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  OAI211_X1 g286(.A(new_n460), .B(KEYINPUT95), .C1(new_n468), .C2(new_n469), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  INV_X1    g288(.A(KEYINPUT13), .ZN(new_n475));
  AOI21_X1  g289(.A(new_n465), .B1(new_n464), .B2(new_n475), .ZN(new_n476));
  NAND3_X1  g290(.A1(new_n461), .A2(new_n463), .A3(KEYINPUT13), .ZN(new_n477));
  AOI21_X1  g291(.A(new_n267), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  AOI21_X1  g292(.A(new_n458), .B1(new_n448), .B2(new_n452), .ZN(new_n479));
  OAI22_X1  g293(.A1(new_n479), .A2(new_n453), .B1(new_n467), .B2(G134), .ZN(new_n480));
  OR3_X1    g294(.A1(new_n478), .A2(new_n480), .A3(KEYINPUT94), .ZN(new_n481));
  OAI21_X1  g295(.A(KEYINPUT94), .B1(new_n478), .B2(new_n480), .ZN(new_n482));
  NAND3_X1  g296(.A1(new_n474), .A2(new_n481), .A3(new_n482), .ZN(new_n483));
  XNOR2_X1  g297(.A(KEYINPUT9), .B(G234), .ZN(new_n484));
  NOR3_X1   g298(.A1(new_n484), .A2(new_n187), .A3(G953), .ZN(new_n485));
  INV_X1    g299(.A(new_n485), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n483), .A2(new_n486), .ZN(new_n487));
  NAND4_X1  g301(.A1(new_n474), .A2(new_n481), .A3(new_n482), .A4(new_n485), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  AOI21_X1  g303(.A(new_n447), .B1(new_n489), .B2(new_n188), .ZN(new_n490));
  AOI211_X1 g304(.A(G902), .B(new_n446), .C1(new_n487), .C2(new_n488), .ZN(new_n491));
  NOR2_X1   g305(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  INV_X1    g306(.A(new_n492), .ZN(new_n493));
  NOR2_X1   g307(.A1(new_n444), .A2(new_n493), .ZN(new_n494));
  OAI21_X1  g308(.A(G221), .B1(new_n484), .B2(G902), .ZN(new_n495));
  INV_X1    g309(.A(G469), .ZN(new_n496));
  XNOR2_X1  g310(.A(G110), .B(G140), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n239), .A2(G227), .ZN(new_n498));
  XOR2_X1   g312(.A(new_n497), .B(new_n498), .Z(new_n499));
  OAI21_X1  g313(.A(KEYINPUT3), .B1(new_n390), .B2(G107), .ZN(new_n500));
  AOI21_X1  g314(.A(G101), .B1(new_n390), .B2(G107), .ZN(new_n501));
  XNOR2_X1  g315(.A(KEYINPUT78), .B(G107), .ZN(new_n502));
  OR2_X1    g316(.A1(new_n390), .A2(KEYINPUT3), .ZN(new_n503));
  OAI211_X1 g317(.A(new_n500), .B(new_n501), .C1(new_n502), .C2(new_n503), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n390), .A2(G107), .ZN(new_n505));
  OAI211_X1 g319(.A(new_n500), .B(new_n505), .C1(new_n502), .C2(new_n503), .ZN(new_n506));
  AOI22_X1  g320(.A1(KEYINPUT4), .A2(new_n504), .B1(new_n506), .B2(G101), .ZN(new_n507));
  AND3_X1   g321(.A1(new_n506), .A2(KEYINPUT4), .A3(G101), .ZN(new_n508));
  OAI21_X1  g322(.A(new_n352), .B1(new_n507), .B2(new_n508), .ZN(new_n509));
  AOI21_X1  g323(.A(G104), .B1(new_n448), .B2(new_n452), .ZN(new_n510));
  INV_X1    g324(.A(KEYINPUT79), .ZN(new_n511));
  OAI21_X1  g325(.A(new_n511), .B1(new_n390), .B2(G107), .ZN(new_n512));
  NAND3_X1  g326(.A1(new_n456), .A2(KEYINPUT79), .A3(G104), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  OAI21_X1  g328(.A(G101), .B1(new_n510), .B2(new_n514), .ZN(new_n515));
  NAND4_X1  g329(.A1(new_n515), .A2(new_n281), .A3(new_n284), .A4(new_n504), .ZN(new_n516));
  INV_X1    g330(.A(KEYINPUT10), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  NAND4_X1  g332(.A1(new_n354), .A2(KEYINPUT10), .A3(new_n504), .A4(new_n515), .ZN(new_n519));
  NAND4_X1  g333(.A1(new_n509), .A2(new_n301), .A3(new_n518), .A4(new_n519), .ZN(new_n520));
  INV_X1    g334(.A(KEYINPUT80), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  AND2_X1   g336(.A1(new_n518), .A2(new_n519), .ZN(new_n523));
  NAND4_X1  g337(.A1(new_n523), .A2(KEYINPUT80), .A3(new_n301), .A4(new_n509), .ZN(new_n524));
  AND2_X1   g338(.A1(new_n522), .A2(new_n524), .ZN(new_n525));
  INV_X1    g339(.A(new_n516), .ZN(new_n526));
  AOI22_X1  g340(.A1(new_n515), .A2(new_n504), .B1(new_n281), .B2(new_n284), .ZN(new_n527));
  OAI211_X1 g341(.A(KEYINPUT81), .B(new_n326), .C1(new_n526), .C2(new_n527), .ZN(new_n528));
  NAND3_X1  g342(.A1(new_n528), .A2(KEYINPUT82), .A3(KEYINPUT12), .ZN(new_n529));
  INV_X1    g343(.A(KEYINPUT12), .ZN(new_n530));
  OAI21_X1  g344(.A(new_n326), .B1(new_n526), .B2(new_n527), .ZN(new_n531));
  OAI21_X1  g345(.A(new_n530), .B1(new_n531), .B2(KEYINPUT82), .ZN(new_n532));
  INV_X1    g346(.A(KEYINPUT82), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n515), .A2(new_n504), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n284), .A2(new_n281), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  AOI21_X1  g350(.A(new_n301), .B1(new_n516), .B2(new_n536), .ZN(new_n537));
  AOI21_X1  g351(.A(new_n533), .B1(new_n537), .B2(KEYINPUT81), .ZN(new_n538));
  OAI21_X1  g352(.A(new_n529), .B1(new_n532), .B2(new_n538), .ZN(new_n539));
  OAI21_X1  g353(.A(new_n499), .B1(new_n525), .B2(new_n539), .ZN(new_n540));
  AOI21_X1  g354(.A(new_n499), .B1(new_n522), .B2(new_n524), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n523), .A2(new_n509), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n542), .A2(new_n326), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n541), .A2(new_n543), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n540), .A2(new_n544), .ZN(new_n545));
  AOI21_X1  g359(.A(new_n496), .B1(new_n545), .B2(new_n188), .ZN(new_n546));
  XOR2_X1   g360(.A(KEYINPUT83), .B(G469), .Z(new_n547));
  NAND2_X1  g361(.A1(new_n522), .A2(new_n524), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n548), .A2(new_n543), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n549), .A2(new_n499), .ZN(new_n550));
  AOI21_X1  g364(.A(KEYINPUT12), .B1(new_n537), .B2(new_n533), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n528), .A2(KEYINPUT82), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  INV_X1    g367(.A(new_n499), .ZN(new_n554));
  NAND4_X1  g368(.A1(new_n548), .A2(new_n553), .A3(new_n529), .A4(new_n554), .ZN(new_n555));
  AOI211_X1 g369(.A(G902), .B(new_n547), .C1(new_n550), .C2(new_n555), .ZN(new_n556));
  OAI21_X1  g370(.A(new_n495), .B1(new_n546), .B2(new_n556), .ZN(new_n557));
  OAI21_X1  g371(.A(G210), .B1(G237), .B2(G902), .ZN(new_n558));
  XOR2_X1   g372(.A(new_n558), .B(KEYINPUT88), .Z(new_n559));
  AOI21_X1  g373(.A(KEYINPUT86), .B1(new_n535), .B2(new_n203), .ZN(new_n560));
  INV_X1    g374(.A(KEYINPUT86), .ZN(new_n561));
  AOI211_X1 g375(.A(new_n561), .B(G125), .C1(new_n284), .C2(new_n281), .ZN(new_n562));
  NOR2_X1   g376(.A1(new_n560), .A2(new_n562), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n310), .A2(G125), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  NAND3_X1  g379(.A1(new_n565), .A2(G224), .A3(new_n239), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n239), .A2(G224), .ZN(new_n567));
  NAND3_X1  g381(.A1(new_n563), .A2(new_n564), .A3(new_n567), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n566), .A2(new_n568), .ZN(new_n569));
  NAND2_X1  g383(.A1(KEYINPUT85), .A2(KEYINPUT6), .ZN(new_n570));
  INV_X1    g384(.A(new_n570), .ZN(new_n571));
  XNOR2_X1  g385(.A(G110), .B(G122), .ZN(new_n572));
  XNOR2_X1  g386(.A(new_n572), .B(KEYINPUT84), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n506), .A2(G101), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n504), .A2(KEYINPUT4), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  NAND3_X1  g390(.A1(new_n506), .A2(KEYINPUT4), .A3(G101), .ZN(new_n577));
  AOI21_X1  g391(.A(new_n297), .B1(new_n576), .B2(new_n577), .ZN(new_n578));
  AND3_X1   g392(.A1(new_n289), .A2(KEYINPUT5), .A3(new_n291), .ZN(new_n579));
  OAI21_X1  g393(.A(G113), .B1(new_n289), .B2(KEYINPUT5), .ZN(new_n580));
  OAI21_X1  g394(.A(new_n296), .B1(new_n579), .B2(new_n580), .ZN(new_n581));
  NOR2_X1   g395(.A1(new_n581), .A2(new_n534), .ZN(new_n582));
  OAI211_X1 g396(.A(new_n571), .B(new_n573), .C1(new_n578), .C2(new_n582), .ZN(new_n583));
  INV_X1    g397(.A(new_n582), .ZN(new_n584));
  OAI21_X1  g398(.A(new_n345), .B1(new_n507), .B2(new_n508), .ZN(new_n585));
  NAND4_X1  g399(.A1(new_n584), .A2(new_n585), .A3(KEYINPUT6), .A4(new_n572), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n583), .A2(new_n586), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n584), .A2(new_n585), .ZN(new_n588));
  AOI21_X1  g402(.A(new_n571), .B1(new_n588), .B2(new_n573), .ZN(new_n589));
  OAI21_X1  g403(.A(new_n569), .B1(new_n587), .B2(new_n589), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n567), .A2(KEYINPUT7), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n565), .A2(new_n591), .ZN(new_n592));
  NAND3_X1  g406(.A1(new_n584), .A2(new_n585), .A3(new_n572), .ZN(new_n593));
  NAND4_X1  g407(.A1(new_n563), .A2(new_n564), .A3(KEYINPUT7), .A4(new_n567), .ZN(new_n594));
  XNOR2_X1  g408(.A(new_n572), .B(KEYINPUT8), .ZN(new_n595));
  AND2_X1   g409(.A1(new_n581), .A2(new_n534), .ZN(new_n596));
  OAI21_X1  g410(.A(new_n595), .B1(new_n596), .B2(new_n582), .ZN(new_n597));
  NAND4_X1  g411(.A1(new_n592), .A2(new_n593), .A3(new_n594), .A4(new_n597), .ZN(new_n598));
  NAND3_X1  g412(.A1(new_n598), .A2(KEYINPUT87), .A3(new_n188), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n590), .A2(new_n599), .ZN(new_n600));
  AOI21_X1  g414(.A(KEYINPUT87), .B1(new_n598), .B2(new_n188), .ZN(new_n601));
  OAI21_X1  g415(.A(new_n559), .B1(new_n600), .B2(new_n601), .ZN(new_n602));
  INV_X1    g416(.A(new_n601), .ZN(new_n603));
  INV_X1    g417(.A(new_n559), .ZN(new_n604));
  NAND4_X1  g418(.A1(new_n603), .A2(new_n604), .A3(new_n590), .A4(new_n599), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n602), .A2(new_n605), .ZN(new_n606));
  NAND2_X1  g420(.A1(G234), .A2(G237), .ZN(new_n607));
  NAND3_X1  g421(.A1(new_n607), .A2(G952), .A3(new_n239), .ZN(new_n608));
  INV_X1    g422(.A(new_n608), .ZN(new_n609));
  NAND3_X1  g423(.A1(new_n607), .A2(G902), .A3(G953), .ZN(new_n610));
  INV_X1    g424(.A(new_n610), .ZN(new_n611));
  XNOR2_X1  g425(.A(KEYINPUT21), .B(G898), .ZN(new_n612));
  AOI21_X1  g426(.A(new_n609), .B1(new_n611), .B2(new_n612), .ZN(new_n613));
  OAI21_X1  g427(.A(G214), .B1(G237), .B2(G902), .ZN(new_n614));
  INV_X1    g428(.A(new_n614), .ZN(new_n615));
  NOR2_X1   g429(.A1(new_n613), .A2(new_n615), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n606), .A2(new_n616), .ZN(new_n617));
  NOR2_X1   g431(.A1(new_n557), .A2(new_n617), .ZN(new_n618));
  NAND3_X1  g432(.A1(new_n388), .A2(new_n494), .A3(new_n618), .ZN(new_n619));
  XNOR2_X1  g433(.A(new_n619), .B(G101), .ZN(G3));
  NOR2_X1   g434(.A1(new_n557), .A2(new_n266), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n364), .A2(new_n188), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n622), .A2(G472), .ZN(new_n623));
  AND3_X1   g437(.A1(new_n368), .A2(new_n623), .A3(new_n370), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n621), .A2(new_n624), .ZN(new_n625));
  INV_X1    g439(.A(KEYINPUT98), .ZN(new_n626));
  NOR3_X1   g440(.A1(new_n600), .A2(new_n559), .A3(new_n601), .ZN(new_n627));
  AOI21_X1  g441(.A(new_n615), .B1(new_n627), .B2(KEYINPUT96), .ZN(new_n628));
  INV_X1    g442(.A(new_n613), .ZN(new_n629));
  INV_X1    g443(.A(KEYINPUT96), .ZN(new_n630));
  NAND3_X1  g444(.A1(new_n602), .A2(new_n605), .A3(new_n630), .ZN(new_n631));
  NAND3_X1  g445(.A1(new_n628), .A2(new_n629), .A3(new_n631), .ZN(new_n632));
  NAND2_X1  g446(.A1(new_n483), .A2(KEYINPUT97), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n633), .A2(KEYINPUT33), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n489), .A2(new_n634), .ZN(new_n635));
  NAND4_X1  g449(.A1(new_n487), .A2(new_n633), .A3(KEYINPUT33), .A4(new_n488), .ZN(new_n636));
  AOI21_X1  g450(.A(new_n445), .B1(new_n635), .B2(new_n636), .ZN(new_n637));
  NAND3_X1  g451(.A1(new_n489), .A2(new_n445), .A3(new_n188), .ZN(new_n638));
  NAND2_X1  g452(.A1(G478), .A2(G902), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  NOR2_X1   g454(.A1(new_n637), .A2(new_n640), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n444), .A2(new_n641), .ZN(new_n642));
  OAI21_X1  g456(.A(new_n626), .B1(new_n632), .B2(new_n642), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n627), .A2(KEYINPUT96), .ZN(new_n644));
  AND3_X1   g458(.A1(new_n631), .A2(new_n644), .A3(new_n614), .ZN(new_n645));
  AND2_X1   g459(.A1(new_n444), .A2(new_n641), .ZN(new_n646));
  NAND4_X1  g460(.A1(new_n645), .A2(new_n646), .A3(KEYINPUT98), .A4(new_n629), .ZN(new_n647));
  AOI21_X1  g461(.A(new_n625), .B1(new_n643), .B2(new_n647), .ZN(new_n648));
  XNOR2_X1  g462(.A(KEYINPUT34), .B(G104), .ZN(new_n649));
  XNOR2_X1  g463(.A(new_n648), .B(new_n649), .ZN(G6));
  NAND2_X1  g464(.A1(new_n493), .A2(new_n443), .ZN(new_n651));
  NAND3_X1  g465(.A1(new_n426), .A2(new_n433), .A3(new_n427), .ZN(new_n652));
  XNOR2_X1  g466(.A(new_n652), .B(KEYINPUT100), .ZN(new_n653));
  INV_X1    g467(.A(KEYINPUT99), .ZN(new_n654));
  AOI21_X1  g468(.A(KEYINPUT91), .B1(new_n428), .B2(KEYINPUT20), .ZN(new_n655));
  NOR3_X1   g469(.A1(new_n432), .A2(new_n430), .A3(new_n433), .ZN(new_n656));
  OAI21_X1  g470(.A(new_n654), .B1(new_n655), .B2(new_n656), .ZN(new_n657));
  NAND3_X1  g471(.A1(new_n429), .A2(KEYINPUT99), .A3(new_n434), .ZN(new_n658));
  AOI21_X1  g472(.A(new_n653), .B1(new_n657), .B2(new_n658), .ZN(new_n659));
  NOR3_X1   g473(.A1(new_n632), .A2(new_n651), .A3(new_n659), .ZN(new_n660));
  NAND3_X1  g474(.A1(new_n660), .A2(new_n624), .A3(new_n621), .ZN(new_n661));
  XOR2_X1   g475(.A(KEYINPUT35), .B(G107), .Z(new_n662));
  XNOR2_X1  g476(.A(new_n661), .B(new_n662), .ZN(G9));
  AOI21_X1  g477(.A(KEYINPUT25), .B1(new_n260), .B2(new_n188), .ZN(new_n664));
  AOI211_X1 g478(.A(new_n247), .B(G902), .C1(new_n258), .C2(new_n259), .ZN(new_n665));
  OAI21_X1  g479(.A(new_n189), .B1(new_n664), .B2(new_n665), .ZN(new_n666));
  NAND2_X1  g480(.A1(new_n230), .A2(new_n238), .ZN(new_n667));
  NOR2_X1   g481(.A1(new_n243), .A2(KEYINPUT36), .ZN(new_n668));
  XNOR2_X1  g482(.A(new_n667), .B(new_n668), .ZN(new_n669));
  NAND2_X1  g483(.A1(new_n669), .A2(new_n263), .ZN(new_n670));
  NAND2_X1  g484(.A1(new_n666), .A2(new_n670), .ZN(new_n671));
  NAND4_X1  g485(.A1(new_n618), .A2(new_n494), .A3(new_n624), .A4(new_n671), .ZN(new_n672));
  XOR2_X1   g486(.A(KEYINPUT37), .B(G110), .Z(new_n673));
  XNOR2_X1  g487(.A(new_n672), .B(new_n673), .ZN(G12));
  NAND2_X1  g488(.A1(new_n371), .A2(new_n387), .ZN(new_n675));
  INV_X1    g489(.A(new_n547), .ZN(new_n676));
  AND4_X1   g490(.A1(new_n548), .A2(new_n553), .A3(new_n529), .A4(new_n554), .ZN(new_n677));
  AOI21_X1  g491(.A(new_n554), .B1(new_n548), .B2(new_n543), .ZN(new_n678));
  OAI211_X1 g492(.A(new_n188), .B(new_n676), .C1(new_n677), .C2(new_n678), .ZN(new_n679));
  AOI21_X1  g493(.A(G902), .B1(new_n540), .B2(new_n544), .ZN(new_n680));
  OAI21_X1  g494(.A(new_n679), .B1(new_n680), .B2(new_n496), .ZN(new_n681));
  AND3_X1   g495(.A1(new_n681), .A2(new_n495), .A3(new_n671), .ZN(new_n682));
  NAND3_X1  g496(.A1(new_n675), .A2(new_n682), .A3(new_n645), .ZN(new_n683));
  OR2_X1    g497(.A1(new_n610), .A2(G900), .ZN(new_n684));
  NAND2_X1  g498(.A1(new_n684), .A2(new_n608), .ZN(new_n685));
  INV_X1    g499(.A(new_n685), .ZN(new_n686));
  OR3_X1    g500(.A1(new_n659), .A2(new_n651), .A3(new_n686), .ZN(new_n687));
  OAI21_X1  g501(.A(KEYINPUT101), .B1(new_n683), .B2(new_n687), .ZN(new_n688));
  NAND3_X1  g502(.A1(new_n681), .A2(new_n671), .A3(new_n495), .ZN(new_n689));
  AOI21_X1  g503(.A(new_n689), .B1(new_n371), .B2(new_n387), .ZN(new_n690));
  INV_X1    g504(.A(KEYINPUT101), .ZN(new_n691));
  NOR3_X1   g505(.A1(new_n659), .A2(new_n651), .A3(new_n686), .ZN(new_n692));
  NAND4_X1  g506(.A1(new_n690), .A2(new_n691), .A3(new_n645), .A4(new_n692), .ZN(new_n693));
  NAND2_X1  g507(.A1(new_n688), .A2(new_n693), .ZN(new_n694));
  XNOR2_X1  g508(.A(new_n694), .B(G128), .ZN(G30));
  INV_X1    g509(.A(new_n495), .ZN(new_n696));
  AND2_X1   g510(.A1(new_n520), .A2(new_n521), .ZN(new_n697));
  NOR2_X1   g511(.A1(new_n520), .A2(new_n521), .ZN(new_n698));
  OAI211_X1 g512(.A(new_n553), .B(new_n529), .C1(new_n697), .C2(new_n698), .ZN(new_n699));
  AOI22_X1  g513(.A1(new_n699), .A2(new_n499), .B1(new_n541), .B2(new_n543), .ZN(new_n700));
  OAI21_X1  g514(.A(G469), .B1(new_n700), .B2(G902), .ZN(new_n701));
  AOI21_X1  g515(.A(new_n696), .B1(new_n701), .B2(new_n679), .ZN(new_n702));
  XNOR2_X1  g516(.A(new_n685), .B(KEYINPUT39), .ZN(new_n703));
  NAND2_X1  g517(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  INV_X1    g518(.A(new_n704), .ZN(new_n705));
  NAND2_X1  g519(.A1(new_n705), .A2(KEYINPUT40), .ZN(new_n706));
  INV_X1    g520(.A(KEYINPUT40), .ZN(new_n707));
  NAND2_X1  g521(.A1(new_n704), .A2(new_n707), .ZN(new_n708));
  NAND2_X1  g522(.A1(new_n706), .A2(new_n708), .ZN(new_n709));
  NAND2_X1  g523(.A1(new_n709), .A2(KEYINPUT104), .ZN(new_n710));
  INV_X1    g524(.A(KEYINPUT104), .ZN(new_n711));
  NAND3_X1  g525(.A1(new_n706), .A2(new_n711), .A3(new_n708), .ZN(new_n712));
  INV_X1    g526(.A(KEYINPUT102), .ZN(new_n713));
  XNOR2_X1  g527(.A(new_n606), .B(new_n713), .ZN(new_n714));
  XOR2_X1   g528(.A(KEYINPUT103), .B(KEYINPUT38), .Z(new_n715));
  XNOR2_X1  g529(.A(new_n714), .B(new_n715), .ZN(new_n716));
  AOI21_X1  g530(.A(new_n320), .B1(new_n346), .B2(new_n311), .ZN(new_n717));
  OAI21_X1  g531(.A(new_n188), .B1(new_n340), .B2(new_n717), .ZN(new_n718));
  AOI22_X1  g532(.A1(new_n372), .A2(KEYINPUT32), .B1(G472), .B2(new_n718), .ZN(new_n719));
  NAND2_X1  g533(.A1(new_n371), .A2(new_n719), .ZN(new_n720));
  INV_X1    g534(.A(new_n670), .ZN(new_n721));
  NOR2_X1   g535(.A1(new_n262), .A2(new_n721), .ZN(new_n722));
  AOI21_X1  g536(.A(new_n492), .B1(new_n438), .B2(new_n443), .ZN(new_n723));
  AND4_X1   g537(.A1(new_n614), .A2(new_n720), .A3(new_n722), .A4(new_n723), .ZN(new_n724));
  NAND4_X1  g538(.A1(new_n710), .A2(new_n712), .A3(new_n716), .A4(new_n724), .ZN(new_n725));
  XNOR2_X1  g539(.A(new_n725), .B(G143), .ZN(G45));
  AND3_X1   g540(.A1(new_n444), .A2(new_n641), .A3(new_n685), .ZN(new_n727));
  NAND4_X1  g541(.A1(new_n690), .A2(KEYINPUT105), .A3(new_n645), .A4(new_n727), .ZN(new_n728));
  NAND4_X1  g542(.A1(new_n675), .A2(new_n682), .A3(new_n645), .A4(new_n727), .ZN(new_n729));
  INV_X1    g543(.A(KEYINPUT105), .ZN(new_n730));
  NAND2_X1  g544(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  NAND2_X1  g545(.A1(new_n728), .A2(new_n731), .ZN(new_n732));
  XNOR2_X1  g546(.A(new_n732), .B(G146), .ZN(G48));
  NOR2_X1   g547(.A1(new_n677), .A2(new_n678), .ZN(new_n734));
  OAI21_X1  g548(.A(G469), .B1(new_n734), .B2(G902), .ZN(new_n735));
  AND3_X1   g549(.A1(new_n735), .A2(new_n495), .A3(new_n679), .ZN(new_n736));
  NAND2_X1  g550(.A1(new_n388), .A2(new_n736), .ZN(new_n737));
  AOI21_X1  g551(.A(new_n737), .B1(new_n643), .B2(new_n647), .ZN(new_n738));
  XOR2_X1   g552(.A(KEYINPUT41), .B(G113), .Z(new_n739));
  XNOR2_X1  g553(.A(new_n738), .B(new_n739), .ZN(G15));
  NAND3_X1  g554(.A1(new_n660), .A2(new_n388), .A3(new_n736), .ZN(new_n741));
  XNOR2_X1  g555(.A(new_n741), .B(G116), .ZN(G18));
  NAND2_X1  g556(.A1(new_n628), .A2(new_n631), .ZN(new_n743));
  NAND3_X1  g557(.A1(new_n735), .A2(new_n495), .A3(new_n679), .ZN(new_n744));
  NOR2_X1   g558(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  NOR2_X1   g559(.A1(new_n722), .A2(new_n613), .ZN(new_n746));
  NAND4_X1  g560(.A1(new_n745), .A2(new_n675), .A3(new_n494), .A4(new_n746), .ZN(new_n747));
  XNOR2_X1  g561(.A(new_n747), .B(G119), .ZN(G21));
  AND3_X1   g562(.A1(new_n628), .A2(new_n723), .A3(new_n631), .ZN(new_n749));
  NAND2_X1  g563(.A1(new_n360), .A2(KEYINPUT31), .ZN(new_n750));
  INV_X1    g564(.A(KEYINPUT106), .ZN(new_n751));
  NAND3_X1  g565(.A1(new_n350), .A2(new_n750), .A3(new_n751), .ZN(new_n752));
  NAND2_X1  g566(.A1(new_n752), .A2(new_n363), .ZN(new_n753));
  AOI21_X1  g567(.A(new_n751), .B1(new_n350), .B2(new_n750), .ZN(new_n754));
  OAI21_X1  g568(.A(new_n365), .B1(new_n753), .B2(new_n754), .ZN(new_n755));
  AND3_X1   g569(.A1(new_n265), .A2(new_n623), .A3(new_n755), .ZN(new_n756));
  NAND4_X1  g570(.A1(new_n749), .A2(new_n756), .A3(new_n629), .A4(new_n736), .ZN(new_n757));
  XNOR2_X1  g571(.A(new_n757), .B(G122), .ZN(G24));
  AND3_X1   g572(.A1(new_n671), .A2(new_n623), .A3(new_n755), .ZN(new_n759));
  NAND4_X1  g573(.A1(new_n759), .A2(new_n645), .A3(new_n727), .A4(new_n736), .ZN(new_n760));
  XOR2_X1   g574(.A(KEYINPUT107), .B(G125), .Z(new_n761));
  XNOR2_X1  g575(.A(new_n760), .B(new_n761), .ZN(G27));
  INV_X1    g576(.A(KEYINPUT110), .ZN(new_n763));
  NAND2_X1  g577(.A1(new_n386), .A2(G472), .ZN(new_n764));
  NAND2_X1  g578(.A1(new_n366), .A2(new_n369), .ZN(new_n765));
  NAND3_X1  g579(.A1(new_n364), .A2(KEYINPUT32), .A3(new_n365), .ZN(new_n766));
  NAND3_X1  g580(.A1(new_n764), .A2(new_n765), .A3(new_n766), .ZN(new_n767));
  NAND4_X1  g581(.A1(new_n727), .A2(KEYINPUT42), .A3(new_n265), .A4(new_n767), .ZN(new_n768));
  INV_X1    g582(.A(new_n768), .ZN(new_n769));
  NAND3_X1  g583(.A1(new_n602), .A2(new_n605), .A3(new_n614), .ZN(new_n770));
  INV_X1    g584(.A(new_n770), .ZN(new_n771));
  INV_X1    g585(.A(KEYINPUT108), .ZN(new_n772));
  OAI21_X1  g586(.A(new_n771), .B1(new_n702), .B2(new_n772), .ZN(new_n773));
  AOI211_X1 g587(.A(KEYINPUT108), .B(new_n696), .C1(new_n701), .C2(new_n679), .ZN(new_n774));
  NOR2_X1   g588(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  AOI21_X1  g589(.A(new_n763), .B1(new_n769), .B2(new_n775), .ZN(new_n776));
  NAND2_X1  g590(.A1(new_n557), .A2(KEYINPUT108), .ZN(new_n777));
  NAND2_X1  g591(.A1(new_n702), .A2(new_n772), .ZN(new_n778));
  NAND3_X1  g592(.A1(new_n777), .A2(new_n778), .A3(new_n771), .ZN(new_n779));
  NOR3_X1   g593(.A1(new_n779), .A2(new_n768), .A3(KEYINPUT110), .ZN(new_n780));
  NOR2_X1   g594(.A1(new_n776), .A2(new_n780), .ZN(new_n781));
  AOI21_X1  g595(.A(new_n770), .B1(new_n557), .B2(KEYINPUT108), .ZN(new_n782));
  NAND4_X1  g596(.A1(new_n388), .A2(new_n782), .A3(new_n727), .A4(new_n778), .ZN(new_n783));
  INV_X1    g597(.A(KEYINPUT109), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  NAND4_X1  g599(.A1(new_n775), .A2(KEYINPUT109), .A3(new_n388), .A4(new_n727), .ZN(new_n786));
  INV_X1    g600(.A(KEYINPUT42), .ZN(new_n787));
  NAND3_X1  g601(.A1(new_n785), .A2(new_n786), .A3(new_n787), .ZN(new_n788));
  NAND2_X1  g602(.A1(new_n781), .A2(new_n788), .ZN(new_n789));
  XNOR2_X1  g603(.A(new_n789), .B(G131), .ZN(G33));
  NAND3_X1  g604(.A1(new_n775), .A2(new_n388), .A3(new_n692), .ZN(new_n791));
  XNOR2_X1  g605(.A(new_n791), .B(G134), .ZN(G36));
  AND2_X1   g606(.A1(new_n438), .A2(new_n443), .ZN(new_n793));
  NAND2_X1  g607(.A1(new_n793), .A2(new_n641), .ZN(new_n794));
  XNOR2_X1  g608(.A(new_n794), .B(KEYINPUT43), .ZN(new_n795));
  INV_X1    g609(.A(KEYINPUT112), .ZN(new_n796));
  NAND2_X1  g610(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  NOR2_X1   g611(.A1(new_n624), .A2(new_n722), .ZN(new_n798));
  NAND2_X1  g612(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  NOR2_X1   g613(.A1(new_n795), .A2(new_n796), .ZN(new_n800));
  INV_X1    g614(.A(KEYINPUT44), .ZN(new_n801));
  NOR3_X1   g615(.A1(new_n799), .A2(new_n800), .A3(new_n801), .ZN(new_n802));
  INV_X1    g616(.A(new_n802), .ZN(new_n803));
  OAI21_X1  g617(.A(new_n801), .B1(new_n799), .B2(new_n800), .ZN(new_n804));
  INV_X1    g618(.A(KEYINPUT45), .ZN(new_n805));
  AOI21_X1  g619(.A(new_n496), .B1(new_n545), .B2(new_n805), .ZN(new_n806));
  OR2_X1    g620(.A1(new_n806), .A2(KEYINPUT111), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n700), .A2(KEYINPUT45), .ZN(new_n808));
  NAND2_X1  g622(.A1(new_n806), .A2(KEYINPUT111), .ZN(new_n809));
  NAND3_X1  g623(.A1(new_n807), .A2(new_n808), .A3(new_n809), .ZN(new_n810));
  NAND2_X1  g624(.A1(G469), .A2(G902), .ZN(new_n811));
  AOI21_X1  g625(.A(KEYINPUT46), .B1(new_n810), .B2(new_n811), .ZN(new_n812));
  INV_X1    g626(.A(new_n812), .ZN(new_n813));
  NAND3_X1  g627(.A1(new_n810), .A2(KEYINPUT46), .A3(new_n811), .ZN(new_n814));
  NAND3_X1  g628(.A1(new_n813), .A2(new_n679), .A3(new_n814), .ZN(new_n815));
  AND3_X1   g629(.A1(new_n815), .A2(new_n495), .A3(new_n703), .ZN(new_n816));
  NAND4_X1  g630(.A1(new_n803), .A2(new_n771), .A3(new_n804), .A4(new_n816), .ZN(new_n817));
  XOR2_X1   g631(.A(KEYINPUT113), .B(G137), .Z(new_n818));
  XNOR2_X1  g632(.A(new_n817), .B(new_n818), .ZN(G39));
  INV_X1    g633(.A(KEYINPUT47), .ZN(new_n820));
  AND3_X1   g634(.A1(new_n810), .A2(KEYINPUT46), .A3(new_n811), .ZN(new_n821));
  NOR3_X1   g635(.A1(new_n821), .A2(new_n812), .A3(new_n556), .ZN(new_n822));
  OAI21_X1  g636(.A(new_n820), .B1(new_n822), .B2(new_n696), .ZN(new_n823));
  NAND3_X1  g637(.A1(new_n815), .A2(KEYINPUT47), .A3(new_n495), .ZN(new_n824));
  NAND2_X1  g638(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  INV_X1    g639(.A(new_n675), .ZN(new_n826));
  NAND4_X1  g640(.A1(new_n826), .A2(new_n266), .A3(new_n727), .A4(new_n771), .ZN(new_n827));
  INV_X1    g641(.A(new_n827), .ZN(new_n828));
  NAND2_X1  g642(.A1(new_n825), .A2(new_n828), .ZN(new_n829));
  XNOR2_X1  g643(.A(new_n829), .B(G140), .ZN(G42));
  INV_X1    g644(.A(new_n716), .ZN(new_n831));
  NAND2_X1  g645(.A1(new_n831), .A2(new_n615), .ZN(new_n832));
  NOR2_X1   g646(.A1(new_n795), .A2(new_n608), .ZN(new_n833));
  NAND3_X1  g647(.A1(new_n833), .A2(new_n736), .A3(new_n756), .ZN(new_n834));
  INV_X1    g648(.A(KEYINPUT50), .ZN(new_n835));
  OR3_X1    g649(.A1(new_n832), .A2(new_n834), .A3(new_n835), .ZN(new_n836));
  OAI21_X1  g650(.A(new_n835), .B1(new_n832), .B2(new_n834), .ZN(new_n837));
  NAND2_X1  g651(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  NAND2_X1  g652(.A1(new_n735), .A2(new_n679), .ZN(new_n839));
  NOR2_X1   g653(.A1(new_n839), .A2(new_n495), .ZN(new_n840));
  INV_X1    g654(.A(new_n840), .ZN(new_n841));
  NAND3_X1  g655(.A1(new_n823), .A2(new_n824), .A3(new_n841), .ZN(new_n842));
  AND3_X1   g656(.A1(new_n833), .A2(new_n756), .A3(new_n771), .ZN(new_n843));
  NAND2_X1  g657(.A1(new_n842), .A2(new_n843), .ZN(new_n844));
  NOR2_X1   g658(.A1(new_n744), .A2(new_n770), .ZN(new_n845));
  AND2_X1   g659(.A1(new_n833), .A2(new_n845), .ZN(new_n846));
  NAND2_X1  g660(.A1(new_n846), .A2(new_n759), .ZN(new_n847));
  INV_X1    g661(.A(new_n720), .ZN(new_n848));
  NAND4_X1  g662(.A1(new_n848), .A2(new_n265), .A3(new_n609), .A4(new_n845), .ZN(new_n849));
  OR3_X1    g663(.A1(new_n849), .A2(new_n444), .A3(new_n641), .ZN(new_n850));
  NAND2_X1  g664(.A1(new_n847), .A2(new_n850), .ZN(new_n851));
  INV_X1    g665(.A(new_n851), .ZN(new_n852));
  NAND4_X1  g666(.A1(new_n838), .A2(new_n844), .A3(KEYINPUT51), .A4(new_n852), .ZN(new_n853));
  INV_X1    g667(.A(KEYINPUT117), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  AOI21_X1  g669(.A(new_n851), .B1(new_n842), .B2(new_n843), .ZN(new_n856));
  NAND4_X1  g670(.A1(new_n856), .A2(KEYINPUT117), .A3(KEYINPUT51), .A4(new_n838), .ZN(new_n857));
  NAND2_X1  g671(.A1(new_n855), .A2(new_n857), .ZN(new_n858));
  AOI21_X1  g672(.A(KEYINPUT51), .B1(new_n856), .B2(new_n838), .ZN(new_n859));
  OR2_X1    g673(.A1(new_n834), .A2(new_n743), .ZN(new_n860));
  AOI21_X1  g674(.A(new_n266), .B1(new_n387), .B2(new_n765), .ZN(new_n861));
  NAND2_X1  g675(.A1(new_n846), .A2(new_n861), .ZN(new_n862));
  AND2_X1   g676(.A1(new_n862), .A2(KEYINPUT48), .ZN(new_n863));
  NOR2_X1   g677(.A1(new_n862), .A2(KEYINPUT48), .ZN(new_n864));
  OAI221_X1 g678(.A(new_n860), .B1(new_n642), .B2(new_n849), .C1(new_n863), .C2(new_n864), .ZN(new_n865));
  NOR2_X1   g679(.A1(new_n859), .A2(new_n865), .ZN(new_n866));
  AND4_X1   g680(.A1(new_n495), .A2(new_n681), .A3(new_n722), .A4(new_n685), .ZN(new_n867));
  NAND3_X1  g681(.A1(new_n867), .A2(new_n749), .A3(new_n720), .ZN(new_n868));
  NAND2_X1  g682(.A1(new_n868), .A2(new_n760), .ZN(new_n869));
  INV_X1    g683(.A(new_n869), .ZN(new_n870));
  AND4_X1   g684(.A1(KEYINPUT52), .A2(new_n694), .A3(new_n732), .A4(new_n870), .ZN(new_n871));
  AOI21_X1  g685(.A(new_n869), .B1(new_n731), .B2(new_n728), .ZN(new_n872));
  AOI21_X1  g686(.A(KEYINPUT52), .B1(new_n872), .B2(new_n694), .ZN(new_n873));
  NOR2_X1   g687(.A1(new_n871), .A2(new_n873), .ZN(new_n874));
  NAND4_X1  g688(.A1(new_n782), .A2(new_n727), .A3(new_n759), .A4(new_n778), .ZN(new_n875));
  NAND3_X1  g689(.A1(new_n492), .A2(new_n443), .A3(new_n685), .ZN(new_n876));
  NOR3_X1   g690(.A1(new_n659), .A2(new_n770), .A3(new_n876), .ZN(new_n877));
  NAND2_X1  g691(.A1(new_n690), .A2(new_n877), .ZN(new_n878));
  NAND3_X1  g692(.A1(new_n791), .A2(new_n875), .A3(new_n878), .ZN(new_n879));
  INV_X1    g693(.A(KEYINPUT115), .ZN(new_n880));
  NAND4_X1  g694(.A1(new_n646), .A2(new_n880), .A3(new_n606), .A4(new_n616), .ZN(new_n881));
  OAI21_X1  g695(.A(KEYINPUT115), .B1(new_n642), .B2(new_n617), .ZN(new_n882));
  NAND4_X1  g696(.A1(new_n881), .A2(new_n624), .A3(new_n882), .A4(new_n621), .ZN(new_n883));
  NAND3_X1  g697(.A1(new_n493), .A2(new_n443), .A3(new_n438), .ZN(new_n884));
  NOR2_X1   g698(.A1(new_n617), .A2(new_n884), .ZN(new_n885));
  NAND3_X1  g699(.A1(new_n621), .A2(new_n624), .A3(new_n885), .ZN(new_n886));
  NAND4_X1  g700(.A1(new_n883), .A2(new_n672), .A3(new_n619), .A4(new_n886), .ZN(new_n887));
  NOR2_X1   g701(.A1(new_n879), .A2(new_n887), .ZN(new_n888));
  NAND3_X1  g702(.A1(new_n741), .A2(new_n747), .A3(new_n757), .ZN(new_n889));
  OAI21_X1  g703(.A(KEYINPUT114), .B1(new_n889), .B2(new_n738), .ZN(new_n890));
  AND2_X1   g704(.A1(new_n747), .A2(new_n757), .ZN(new_n891));
  NAND2_X1  g705(.A1(new_n647), .A2(new_n643), .ZN(new_n892));
  NAND3_X1  g706(.A1(new_n892), .A2(new_n388), .A3(new_n736), .ZN(new_n893));
  INV_X1    g707(.A(KEYINPUT114), .ZN(new_n894));
  NAND4_X1  g708(.A1(new_n891), .A2(new_n893), .A3(new_n894), .A4(new_n741), .ZN(new_n895));
  NAND4_X1  g709(.A1(new_n789), .A2(new_n888), .A3(new_n890), .A4(new_n895), .ZN(new_n896));
  OAI21_X1  g710(.A(KEYINPUT53), .B1(new_n874), .B2(new_n896), .ZN(new_n897));
  NAND3_X1  g711(.A1(new_n694), .A2(new_n732), .A3(new_n870), .ZN(new_n898));
  INV_X1    g712(.A(KEYINPUT52), .ZN(new_n899));
  NAND3_X1  g713(.A1(new_n898), .A2(KEYINPUT116), .A3(new_n899), .ZN(new_n900));
  NAND3_X1  g714(.A1(new_n872), .A2(KEYINPUT52), .A3(new_n694), .ZN(new_n901));
  NAND2_X1  g715(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  NOR2_X1   g716(.A1(new_n873), .A2(KEYINPUT116), .ZN(new_n903));
  NOR2_X1   g717(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  AND2_X1   g718(.A1(new_n890), .A2(new_n895), .ZN(new_n905));
  INV_X1    g719(.A(KEYINPUT53), .ZN(new_n906));
  NAND4_X1  g720(.A1(new_n905), .A2(new_n906), .A3(new_n789), .A4(new_n888), .ZN(new_n907));
  OAI211_X1 g721(.A(new_n897), .B(KEYINPUT54), .C1(new_n904), .C2(new_n907), .ZN(new_n908));
  NOR3_X1   g722(.A1(new_n889), .A2(new_n738), .A3(new_n906), .ZN(new_n909));
  AND3_X1   g723(.A1(new_n789), .A2(new_n888), .A3(new_n909), .ZN(new_n910));
  OAI21_X1  g724(.A(new_n910), .B1(new_n902), .B2(new_n903), .ZN(new_n911));
  OAI21_X1  g725(.A(new_n906), .B1(new_n874), .B2(new_n896), .ZN(new_n912));
  INV_X1    g726(.A(KEYINPUT54), .ZN(new_n913));
  NAND3_X1  g727(.A1(new_n911), .A2(new_n912), .A3(new_n913), .ZN(new_n914));
  NAND4_X1  g728(.A1(new_n858), .A2(new_n866), .A3(new_n908), .A4(new_n914), .ZN(new_n915));
  INV_X1    g729(.A(KEYINPUT118), .ZN(new_n916));
  OAI211_X1 g730(.A(G952), .B(new_n239), .C1(new_n915), .C2(new_n916), .ZN(new_n917));
  OAI21_X1  g731(.A(G953), .B1(new_n915), .B2(KEYINPUT118), .ZN(new_n918));
  AND2_X1   g732(.A1(new_n839), .A2(KEYINPUT49), .ZN(new_n919));
  NOR2_X1   g733(.A1(new_n839), .A2(KEYINPUT49), .ZN(new_n920));
  NAND4_X1  g734(.A1(new_n265), .A2(new_n641), .A3(new_n495), .A4(new_n614), .ZN(new_n921));
  NOR3_X1   g735(.A1(new_n919), .A2(new_n920), .A3(new_n921), .ZN(new_n922));
  NAND4_X1  g736(.A1(new_n831), .A2(new_n793), .A3(new_n848), .A4(new_n922), .ZN(new_n923));
  NAND3_X1  g737(.A1(new_n917), .A2(new_n918), .A3(new_n923), .ZN(G75));
  NOR2_X1   g738(.A1(new_n239), .A2(G952), .ZN(new_n925));
  INV_X1    g739(.A(new_n925), .ZN(new_n926));
  AOI21_X1  g740(.A(new_n188), .B1(new_n911), .B2(new_n912), .ZN(new_n927));
  AOI21_X1  g741(.A(KEYINPUT56), .B1(new_n927), .B2(new_n559), .ZN(new_n928));
  NOR2_X1   g742(.A1(new_n587), .A2(new_n589), .ZN(new_n929));
  XOR2_X1   g743(.A(new_n929), .B(new_n569), .Z(new_n930));
  XNOR2_X1  g744(.A(new_n930), .B(KEYINPUT55), .ZN(new_n931));
  INV_X1    g745(.A(new_n931), .ZN(new_n932));
  OAI21_X1  g746(.A(new_n926), .B1(new_n928), .B2(new_n932), .ZN(new_n933));
  AOI21_X1  g747(.A(new_n933), .B1(new_n928), .B2(new_n932), .ZN(G51));
  XNOR2_X1  g748(.A(new_n811), .B(KEYINPUT119), .ZN(new_n935));
  XNOR2_X1  g749(.A(new_n935), .B(KEYINPUT57), .ZN(new_n936));
  AND3_X1   g750(.A1(new_n911), .A2(new_n912), .A3(new_n913), .ZN(new_n937));
  AOI21_X1  g751(.A(new_n913), .B1(new_n911), .B2(new_n912), .ZN(new_n938));
  OAI21_X1  g752(.A(new_n936), .B1(new_n937), .B2(new_n938), .ZN(new_n939));
  INV_X1    g753(.A(KEYINPUT120), .ZN(new_n940));
  NAND2_X1  g754(.A1(new_n939), .A2(new_n940), .ZN(new_n941));
  INV_X1    g755(.A(new_n734), .ZN(new_n942));
  OAI211_X1 g756(.A(KEYINPUT120), .B(new_n936), .C1(new_n937), .C2(new_n938), .ZN(new_n943));
  NAND3_X1  g757(.A1(new_n941), .A2(new_n942), .A3(new_n943), .ZN(new_n944));
  INV_X1    g758(.A(new_n810), .ZN(new_n945));
  NAND2_X1  g759(.A1(new_n927), .A2(new_n945), .ZN(new_n946));
  AOI21_X1  g760(.A(new_n925), .B1(new_n944), .B2(new_n946), .ZN(G54));
  NAND3_X1  g761(.A1(new_n927), .A2(KEYINPUT58), .A3(G475), .ZN(new_n948));
  INV_X1    g762(.A(new_n426), .ZN(new_n949));
  AND2_X1   g763(.A1(new_n948), .A2(new_n949), .ZN(new_n950));
  NOR2_X1   g764(.A1(new_n948), .A2(new_n949), .ZN(new_n951));
  NOR3_X1   g765(.A1(new_n950), .A2(new_n951), .A3(new_n925), .ZN(G60));
  NAND2_X1  g766(.A1(new_n908), .A2(new_n914), .ZN(new_n953));
  XNOR2_X1  g767(.A(new_n639), .B(KEYINPUT59), .ZN(new_n954));
  NAND2_X1  g768(.A1(new_n953), .A2(new_n954), .ZN(new_n955));
  AND2_X1   g769(.A1(new_n635), .A2(new_n636), .ZN(new_n956));
  XNOR2_X1  g770(.A(new_n956), .B(KEYINPUT121), .ZN(new_n957));
  INV_X1    g771(.A(new_n957), .ZN(new_n958));
  NAND2_X1  g772(.A1(new_n955), .A2(new_n958), .ZN(new_n959));
  INV_X1    g773(.A(KEYINPUT122), .ZN(new_n960));
  AND2_X1   g774(.A1(new_n957), .A2(new_n954), .ZN(new_n961));
  OAI21_X1  g775(.A(new_n961), .B1(new_n937), .B2(new_n938), .ZN(new_n962));
  NAND4_X1  g776(.A1(new_n959), .A2(new_n960), .A3(new_n926), .A4(new_n962), .ZN(new_n963));
  NAND2_X1  g777(.A1(new_n962), .A2(new_n926), .ZN(new_n964));
  AOI21_X1  g778(.A(new_n957), .B1(new_n953), .B2(new_n954), .ZN(new_n965));
  OAI21_X1  g779(.A(KEYINPUT122), .B1(new_n964), .B2(new_n965), .ZN(new_n966));
  NAND2_X1  g780(.A1(new_n963), .A2(new_n966), .ZN(G63));
  NAND2_X1  g781(.A1(G217), .A2(G902), .ZN(new_n968));
  XNOR2_X1  g782(.A(new_n968), .B(KEYINPUT60), .ZN(new_n969));
  AOI21_X1  g783(.A(new_n969), .B1(new_n911), .B2(new_n912), .ZN(new_n970));
  NAND2_X1  g784(.A1(new_n970), .A2(new_n669), .ZN(new_n971));
  OAI211_X1 g785(.A(new_n971), .B(new_n926), .C1(new_n260), .C2(new_n970), .ZN(new_n972));
  AOI21_X1  g786(.A(KEYINPUT61), .B1(new_n971), .B2(KEYINPUT123), .ZN(new_n973));
  XNOR2_X1  g787(.A(new_n972), .B(new_n973), .ZN(G66));
  INV_X1    g788(.A(new_n612), .ZN(new_n975));
  AOI21_X1  g789(.A(new_n239), .B1(new_n975), .B2(G224), .ZN(new_n976));
  INV_X1    g790(.A(new_n887), .ZN(new_n977));
  NAND2_X1  g791(.A1(new_n905), .A2(new_n977), .ZN(new_n978));
  AOI21_X1  g792(.A(new_n976), .B1(new_n978), .B2(new_n239), .ZN(new_n979));
  OAI21_X1  g793(.A(new_n929), .B1(G898), .B2(new_n239), .ZN(new_n980));
  XOR2_X1   g794(.A(new_n979), .B(new_n980), .Z(G69));
  NAND2_X1  g795(.A1(new_n642), .A2(new_n884), .ZN(new_n982));
  AND3_X1   g796(.A1(new_n388), .A2(new_n705), .A3(new_n771), .ZN(new_n983));
  AOI22_X1  g797(.A1(new_n825), .A2(new_n828), .B1(new_n982), .B2(new_n983), .ZN(new_n984));
  AND2_X1   g798(.A1(new_n732), .A2(new_n760), .ZN(new_n985));
  NAND3_X1  g799(.A1(new_n985), .A2(new_n694), .A3(new_n725), .ZN(new_n986));
  NAND2_X1  g800(.A1(new_n986), .A2(KEYINPUT62), .ZN(new_n987));
  INV_X1    g801(.A(KEYINPUT62), .ZN(new_n988));
  NAND4_X1  g802(.A1(new_n985), .A2(new_n725), .A3(new_n988), .A4(new_n694), .ZN(new_n989));
  NAND4_X1  g803(.A1(new_n984), .A2(new_n817), .A3(new_n987), .A4(new_n989), .ZN(new_n990));
  NAND2_X1  g804(.A1(new_n990), .A2(new_n239), .ZN(new_n991));
  NAND2_X1  g805(.A1(new_n324), .A2(new_n357), .ZN(new_n992));
  XOR2_X1   g806(.A(new_n992), .B(new_n421), .Z(new_n993));
  NAND2_X1  g807(.A1(new_n991), .A2(new_n993), .ZN(new_n994));
  AOI21_X1  g808(.A(new_n993), .B1(G900), .B2(G953), .ZN(new_n995));
  AND2_X1   g809(.A1(new_n861), .A2(new_n749), .ZN(new_n996));
  NAND4_X1  g810(.A1(new_n815), .A2(new_n495), .A3(new_n703), .A4(new_n996), .ZN(new_n997));
  NAND4_X1  g811(.A1(new_n997), .A2(new_n985), .A3(new_n694), .A4(new_n791), .ZN(new_n998));
  INV_X1    g812(.A(new_n998), .ZN(new_n999));
  NAND4_X1  g813(.A1(new_n999), .A2(new_n789), .A3(new_n829), .A4(new_n817), .ZN(new_n1000));
  OAI21_X1  g814(.A(new_n995), .B1(new_n1000), .B2(G953), .ZN(new_n1001));
  NAND3_X1  g815(.A1(new_n994), .A2(KEYINPUT124), .A3(new_n1001), .ZN(new_n1002));
  AOI21_X1  g816(.A(new_n239), .B1(G227), .B2(G900), .ZN(new_n1003));
  XNOR2_X1  g817(.A(new_n1002), .B(new_n1003), .ZN(G72));
  XNOR2_X1  g818(.A(KEYINPUT125), .B(KEYINPUT63), .ZN(new_n1005));
  NAND2_X1  g819(.A1(G472), .A2(G902), .ZN(new_n1006));
  XNOR2_X1  g820(.A(new_n1005), .B(new_n1006), .ZN(new_n1007));
  INV_X1    g821(.A(new_n1007), .ZN(new_n1008));
  OAI21_X1  g822(.A(new_n1008), .B1(new_n990), .B2(new_n978), .ZN(new_n1009));
  XNOR2_X1  g823(.A(new_n381), .B(KEYINPUT126), .ZN(new_n1010));
  NAND3_X1  g824(.A1(new_n1009), .A2(new_n320), .A3(new_n1010), .ZN(new_n1011));
  OAI21_X1  g825(.A(new_n1008), .B1(new_n1000), .B2(new_n978), .ZN(new_n1012));
  NOR2_X1   g826(.A1(new_n1010), .A2(new_n320), .ZN(new_n1013));
  NAND2_X1  g827(.A1(new_n1012), .A2(new_n1013), .ZN(new_n1014));
  AOI21_X1  g828(.A(new_n1007), .B1(new_n382), .B2(new_n360), .ZN(new_n1015));
  OAI211_X1 g829(.A(new_n897), .B(new_n1015), .C1(new_n904), .C2(new_n907), .ZN(new_n1016));
  AND2_X1   g830(.A1(new_n1016), .A2(new_n926), .ZN(new_n1017));
  NAND3_X1  g831(.A1(new_n1011), .A2(new_n1014), .A3(new_n1017), .ZN(new_n1018));
  INV_X1    g832(.A(KEYINPUT127), .ZN(new_n1019));
  NAND2_X1  g833(.A1(new_n1018), .A2(new_n1019), .ZN(new_n1020));
  NAND4_X1  g834(.A1(new_n1011), .A2(new_n1014), .A3(new_n1017), .A4(KEYINPUT127), .ZN(new_n1021));
  NAND2_X1  g835(.A1(new_n1020), .A2(new_n1021), .ZN(G57));
endmodule


