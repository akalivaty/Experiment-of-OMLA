

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302,
         n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313,
         n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324,
         n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335,
         n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346,
         n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590, n591, n592;

  XOR2_X1 U324 ( .A(KEYINPUT62), .B(n592), .Z(n292) );
  XNOR2_X1 U325 ( .A(n302), .B(n301), .ZN(n304) );
  XNOR2_X1 U326 ( .A(n330), .B(KEYINPUT9), .ZN(n331) );
  XNOR2_X1 U327 ( .A(n332), .B(n331), .ZN(n335) );
  XOR2_X1 U328 ( .A(KEYINPUT34), .B(KEYINPUT98), .Z(n453) );
  XOR2_X1 U329 ( .A(G113GAT), .B(G15GAT), .Z(n434) );
  XNOR2_X1 U330 ( .A(G1GAT), .B(KEYINPUT67), .ZN(n293) );
  XNOR2_X1 U331 ( .A(n293), .B(G8GAT), .ZN(n345) );
  XOR2_X1 U332 ( .A(n434), .B(n345), .Z(n295) );
  NAND2_X1 U333 ( .A1(G229GAT), .A2(G233GAT), .ZN(n294) );
  XNOR2_X1 U334 ( .A(n295), .B(n294), .ZN(n296) );
  XOR2_X1 U335 ( .A(n296), .B(G197GAT), .Z(n298) );
  XOR2_X1 U336 ( .A(G141GAT), .B(G22GAT), .Z(n364) );
  XNOR2_X1 U337 ( .A(G169GAT), .B(n364), .ZN(n297) );
  XNOR2_X1 U338 ( .A(n298), .B(n297), .ZN(n309) );
  XNOR2_X1 U339 ( .A(KEYINPUT66), .B(G50GAT), .ZN(n300) );
  INV_X1 U340 ( .A(KEYINPUT7), .ZN(n299) );
  XNOR2_X1 U341 ( .A(n300), .B(n299), .ZN(n302) );
  XOR2_X1 U342 ( .A(G43GAT), .B(G29GAT), .Z(n301) );
  XNOR2_X1 U343 ( .A(G36GAT), .B(KEYINPUT8), .ZN(n303) );
  XNOR2_X1 U344 ( .A(n304), .B(n303), .ZN(n327) );
  XOR2_X1 U345 ( .A(KEYINPUT30), .B(KEYINPUT65), .Z(n306) );
  XNOR2_X1 U346 ( .A(KEYINPUT64), .B(KEYINPUT29), .ZN(n305) );
  XNOR2_X1 U347 ( .A(n306), .B(n305), .ZN(n307) );
  XOR2_X1 U348 ( .A(n327), .B(n307), .Z(n308) );
  XOR2_X1 U349 ( .A(n309), .B(n308), .Z(n533) );
  XOR2_X1 U350 ( .A(KEYINPUT68), .B(n533), .Z(n554) );
  INV_X1 U351 ( .A(n554), .ZN(n519) );
  XOR2_X1 U352 ( .A(G92GAT), .B(G85GAT), .Z(n311) );
  XNOR2_X1 U353 ( .A(G99GAT), .B(G106GAT), .ZN(n310) );
  XNOR2_X1 U354 ( .A(n311), .B(n310), .ZN(n333) );
  XOR2_X1 U355 ( .A(KEYINPUT70), .B(KEYINPUT33), .Z(n313) );
  XNOR2_X1 U356 ( .A(G176GAT), .B(KEYINPUT69), .ZN(n312) );
  XNOR2_X1 U357 ( .A(n313), .B(n312), .ZN(n314) );
  XOR2_X1 U358 ( .A(n333), .B(n314), .Z(n316) );
  XOR2_X1 U359 ( .A(G120GAT), .B(G71GAT), .Z(n427) );
  XOR2_X1 U360 ( .A(G148GAT), .B(G78GAT), .Z(n370) );
  XNOR2_X1 U361 ( .A(n427), .B(n370), .ZN(n315) );
  XNOR2_X1 U362 ( .A(n316), .B(n315), .ZN(n323) );
  XOR2_X1 U363 ( .A(KEYINPUT71), .B(KEYINPUT32), .Z(n318) );
  NAND2_X1 U364 ( .A1(G230GAT), .A2(G233GAT), .ZN(n317) );
  XNOR2_X1 U365 ( .A(n318), .B(n317), .ZN(n319) );
  XOR2_X1 U366 ( .A(n319), .B(KEYINPUT31), .Z(n321) );
  XOR2_X1 U367 ( .A(G57GAT), .B(KEYINPUT13), .Z(n341) );
  XOR2_X1 U368 ( .A(G204GAT), .B(G64GAT), .Z(n415) );
  XNOR2_X1 U369 ( .A(n341), .B(n415), .ZN(n320) );
  XNOR2_X1 U370 ( .A(n321), .B(n320), .ZN(n322) );
  XNOR2_X1 U371 ( .A(n323), .B(n322), .ZN(n583) );
  NAND2_X1 U372 ( .A1(n519), .A2(n583), .ZN(n466) );
  XNOR2_X1 U373 ( .A(KEYINPUT11), .B(KEYINPUT72), .ZN(n324) );
  XOR2_X1 U374 ( .A(G218GAT), .B(G162GAT), .Z(n371) );
  XOR2_X1 U375 ( .A(n324), .B(n371), .Z(n337) );
  INV_X1 U376 ( .A(n327), .ZN(n326) );
  XOR2_X1 U377 ( .A(G190GAT), .B(G134GAT), .Z(n428) );
  INV_X1 U378 ( .A(n428), .ZN(n325) );
  NAND2_X1 U379 ( .A1(n326), .A2(n325), .ZN(n329) );
  NAND2_X1 U380 ( .A1(n327), .A2(n428), .ZN(n328) );
  NAND2_X1 U381 ( .A1(n329), .A2(n328), .ZN(n332) );
  AND2_X1 U382 ( .A1(G232GAT), .A2(G233GAT), .ZN(n330) );
  XOR2_X1 U383 ( .A(n333), .B(KEYINPUT10), .Z(n334) );
  XNOR2_X1 U384 ( .A(n335), .B(n334), .ZN(n336) );
  XNOR2_X1 U385 ( .A(n337), .B(n336), .ZN(n543) );
  XOR2_X1 U386 ( .A(KEYINPUT73), .B(n543), .Z(n461) );
  INV_X1 U387 ( .A(n461), .ZN(n566) );
  XOR2_X1 U388 ( .A(G71GAT), .B(G127GAT), .Z(n339) );
  XNOR2_X1 U389 ( .A(G15GAT), .B(G183GAT), .ZN(n338) );
  XNOR2_X1 U390 ( .A(n339), .B(n338), .ZN(n340) );
  XOR2_X1 U391 ( .A(n341), .B(n340), .Z(n343) );
  NAND2_X1 U392 ( .A1(G231GAT), .A2(G233GAT), .ZN(n342) );
  XNOR2_X1 U393 ( .A(n343), .B(n342), .ZN(n344) );
  XOR2_X1 U394 ( .A(n344), .B(KEYINPUT79), .Z(n347) );
  XNOR2_X1 U395 ( .A(n345), .B(KEYINPUT78), .ZN(n346) );
  XNOR2_X1 U396 ( .A(n347), .B(n346), .ZN(n351) );
  XOR2_X1 U397 ( .A(G211GAT), .B(G78GAT), .Z(n349) );
  XNOR2_X1 U398 ( .A(G22GAT), .B(G155GAT), .ZN(n348) );
  XNOR2_X1 U399 ( .A(n349), .B(n348), .ZN(n350) );
  XOR2_X1 U400 ( .A(n351), .B(n350), .Z(n359) );
  XOR2_X1 U401 ( .A(KEYINPUT15), .B(KEYINPUT14), .Z(n353) );
  XNOR2_X1 U402 ( .A(G64GAT), .B(KEYINPUT77), .ZN(n352) );
  XNOR2_X1 U403 ( .A(n353), .B(n352), .ZN(n357) );
  XOR2_X1 U404 ( .A(KEYINPUT12), .B(KEYINPUT76), .Z(n355) );
  XNOR2_X1 U405 ( .A(KEYINPUT75), .B(KEYINPUT74), .ZN(n354) );
  XNOR2_X1 U406 ( .A(n355), .B(n354), .ZN(n356) );
  XNOR2_X1 U407 ( .A(n357), .B(n356), .ZN(n358) );
  XOR2_X1 U408 ( .A(n359), .B(n358), .Z(n541) );
  INV_X1 U409 ( .A(n541), .ZN(n588) );
  NOR2_X1 U410 ( .A1(n461), .A2(n588), .ZN(n360) );
  XNOR2_X1 U411 ( .A(n360), .B(KEYINPUT16), .ZN(n451) );
  XOR2_X1 U412 ( .A(KEYINPUT90), .B(KEYINPUT24), .Z(n362) );
  XNOR2_X1 U413 ( .A(G204GAT), .B(KEYINPUT92), .ZN(n361) );
  XNOR2_X1 U414 ( .A(n362), .B(n361), .ZN(n363) );
  XOR2_X1 U415 ( .A(n363), .B(G106GAT), .Z(n366) );
  XNOR2_X1 U416 ( .A(G50GAT), .B(n364), .ZN(n365) );
  XNOR2_X1 U417 ( .A(n366), .B(n365), .ZN(n369) );
  XOR2_X1 U418 ( .A(G211GAT), .B(KEYINPUT21), .Z(n368) );
  XNOR2_X1 U419 ( .A(G197GAT), .B(KEYINPUT89), .ZN(n367) );
  XNOR2_X1 U420 ( .A(n368), .B(n367), .ZN(n414) );
  XOR2_X1 U421 ( .A(n369), .B(n414), .Z(n373) );
  XNOR2_X1 U422 ( .A(n371), .B(n370), .ZN(n372) );
  XNOR2_X1 U423 ( .A(n373), .B(n372), .ZN(n382) );
  XOR2_X1 U424 ( .A(KEYINPUT23), .B(KEYINPUT22), .Z(n375) );
  XNOR2_X1 U425 ( .A(KEYINPUT88), .B(KEYINPUT87), .ZN(n374) );
  XNOR2_X1 U426 ( .A(n375), .B(n374), .ZN(n380) );
  XNOR2_X1 U427 ( .A(G155GAT), .B(KEYINPUT3), .ZN(n376) );
  XNOR2_X1 U428 ( .A(n376), .B(KEYINPUT2), .ZN(n386) );
  XOR2_X1 U429 ( .A(KEYINPUT91), .B(n386), .Z(n378) );
  NAND2_X1 U430 ( .A1(G228GAT), .A2(G233GAT), .ZN(n377) );
  XNOR2_X1 U431 ( .A(n378), .B(n377), .ZN(n379) );
  XOR2_X1 U432 ( .A(n380), .B(n379), .Z(n381) );
  XNOR2_X1 U433 ( .A(n382), .B(n381), .ZN(n551) );
  XOR2_X1 U434 ( .A(KEYINPUT28), .B(n551), .Z(n497) );
  INV_X1 U435 ( .A(n497), .ZN(n517) );
  XOR2_X1 U436 ( .A(KEYINPUT4), .B(KEYINPUT93), .Z(n384) );
  XNOR2_X1 U437 ( .A(G1GAT), .B(G57GAT), .ZN(n383) );
  XNOR2_X1 U438 ( .A(n384), .B(n383), .ZN(n401) );
  XNOR2_X1 U439 ( .A(G127GAT), .B(KEYINPUT0), .ZN(n385) );
  XNOR2_X1 U440 ( .A(n385), .B(KEYINPUT80), .ZN(n423) );
  XNOR2_X1 U441 ( .A(n423), .B(n386), .ZN(n399) );
  XOR2_X1 U442 ( .A(G85GAT), .B(G162GAT), .Z(n388) );
  XNOR2_X1 U443 ( .A(G29GAT), .B(G134GAT), .ZN(n387) );
  XNOR2_X1 U444 ( .A(n388), .B(n387), .ZN(n392) );
  XOR2_X1 U445 ( .A(G148GAT), .B(G120GAT), .Z(n390) );
  XNOR2_X1 U446 ( .A(G141GAT), .B(G113GAT), .ZN(n389) );
  XNOR2_X1 U447 ( .A(n390), .B(n389), .ZN(n391) );
  XOR2_X1 U448 ( .A(n392), .B(n391), .Z(n397) );
  XOR2_X1 U449 ( .A(KEYINPUT6), .B(KEYINPUT1), .Z(n394) );
  NAND2_X1 U450 ( .A1(G225GAT), .A2(G233GAT), .ZN(n393) );
  XNOR2_X1 U451 ( .A(n394), .B(n393), .ZN(n395) );
  XNOR2_X1 U452 ( .A(KEYINPUT5), .B(n395), .ZN(n396) );
  XNOR2_X1 U453 ( .A(n397), .B(n396), .ZN(n398) );
  XNOR2_X1 U454 ( .A(n399), .B(n398), .ZN(n400) );
  XOR2_X1 U455 ( .A(n401), .B(n400), .Z(n550) );
  INV_X1 U456 ( .A(n550), .ZN(n573) );
  XOR2_X1 U457 ( .A(G176GAT), .B(G183GAT), .Z(n403) );
  XNOR2_X1 U458 ( .A(G169GAT), .B(KEYINPUT18), .ZN(n402) );
  XNOR2_X1 U459 ( .A(n403), .B(n402), .ZN(n407) );
  XOR2_X1 U460 ( .A(KEYINPUT19), .B(KEYINPUT84), .Z(n405) );
  XNOR2_X1 U461 ( .A(KEYINPUT17), .B(KEYINPUT83), .ZN(n404) );
  XNOR2_X1 U462 ( .A(n405), .B(n404), .ZN(n406) );
  XOR2_X1 U463 ( .A(n407), .B(n406), .Z(n433) );
  XOR2_X1 U464 ( .A(KEYINPUT72), .B(G218GAT), .Z(n409) );
  XNOR2_X1 U465 ( .A(G36GAT), .B(G190GAT), .ZN(n408) );
  XNOR2_X1 U466 ( .A(n409), .B(n408), .ZN(n413) );
  XOR2_X1 U467 ( .A(KEYINPUT94), .B(KEYINPUT95), .Z(n411) );
  XNOR2_X1 U468 ( .A(G8GAT), .B(G92GAT), .ZN(n410) );
  XNOR2_X1 U469 ( .A(n411), .B(n410), .ZN(n412) );
  XNOR2_X1 U470 ( .A(n413), .B(n412), .ZN(n419) );
  XOR2_X1 U471 ( .A(n415), .B(n414), .Z(n417) );
  NAND2_X1 U472 ( .A1(G226GAT), .A2(G233GAT), .ZN(n416) );
  XNOR2_X1 U473 ( .A(n417), .B(n416), .ZN(n418) );
  XNOR2_X1 U474 ( .A(n419), .B(n418), .ZN(n420) );
  XOR2_X1 U475 ( .A(n433), .B(n420), .Z(n546) );
  XNOR2_X1 U476 ( .A(KEYINPUT27), .B(n546), .ZN(n443) );
  NAND2_X1 U477 ( .A1(n573), .A2(n443), .ZN(n515) );
  XOR2_X1 U478 ( .A(KEYINPUT85), .B(KEYINPUT82), .Z(n426) );
  XOR2_X1 U479 ( .A(KEYINPUT81), .B(KEYINPUT20), .Z(n422) );
  XNOR2_X1 U480 ( .A(G43GAT), .B(G99GAT), .ZN(n421) );
  XNOR2_X1 U481 ( .A(n422), .B(n421), .ZN(n424) );
  XNOR2_X1 U482 ( .A(n424), .B(n423), .ZN(n425) );
  XNOR2_X1 U483 ( .A(n426), .B(n425), .ZN(n432) );
  XOR2_X1 U484 ( .A(n428), .B(n427), .Z(n430) );
  NAND2_X1 U485 ( .A1(G227GAT), .A2(G233GAT), .ZN(n429) );
  XNOR2_X1 U486 ( .A(n430), .B(n429), .ZN(n431) );
  XOR2_X1 U487 ( .A(n432), .B(n431), .Z(n436) );
  XNOR2_X1 U488 ( .A(n434), .B(n433), .ZN(n435) );
  XNOR2_X1 U489 ( .A(n436), .B(n435), .ZN(n564) );
  XNOR2_X1 U490 ( .A(KEYINPUT86), .B(n564), .ZN(n437) );
  NOR2_X1 U491 ( .A1(n515), .A2(n437), .ZN(n438) );
  NAND2_X1 U492 ( .A1(n517), .A2(n438), .ZN(n450) );
  NOR2_X1 U493 ( .A1(n564), .A2(n551), .ZN(n440) );
  XNOR2_X1 U494 ( .A(KEYINPUT97), .B(KEYINPUT26), .ZN(n439) );
  XNOR2_X1 U495 ( .A(n440), .B(n439), .ZN(n441) );
  XNOR2_X1 U496 ( .A(KEYINPUT96), .B(n441), .ZN(n572) );
  INV_X1 U497 ( .A(n572), .ZN(n442) );
  NAND2_X1 U498 ( .A1(n443), .A2(n442), .ZN(n447) );
  NAND2_X1 U499 ( .A1(n564), .A2(n546), .ZN(n444) );
  NAND2_X1 U500 ( .A1(n551), .A2(n444), .ZN(n445) );
  XOR2_X1 U501 ( .A(KEYINPUT25), .B(n445), .Z(n446) );
  NAND2_X1 U502 ( .A1(n447), .A2(n446), .ZN(n448) );
  NAND2_X1 U503 ( .A1(n448), .A2(n550), .ZN(n449) );
  NAND2_X1 U504 ( .A1(n450), .A2(n449), .ZN(n462) );
  NAND2_X1 U505 ( .A1(n451), .A2(n462), .ZN(n479) );
  NOR2_X1 U506 ( .A1(n466), .A2(n479), .ZN(n459) );
  NAND2_X1 U507 ( .A1(n459), .A2(n573), .ZN(n452) );
  XNOR2_X1 U508 ( .A(n453), .B(n452), .ZN(n454) );
  XOR2_X1 U509 ( .A(G1GAT), .B(n454), .Z(G1324GAT) );
  NAND2_X1 U510 ( .A1(n459), .A2(n546), .ZN(n455) );
  XNOR2_X1 U511 ( .A(n455), .B(G8GAT), .ZN(G1325GAT) );
  XOR2_X1 U512 ( .A(KEYINPUT99), .B(KEYINPUT35), .Z(n457) );
  NAND2_X1 U513 ( .A1(n459), .A2(n564), .ZN(n456) );
  XNOR2_X1 U514 ( .A(n457), .B(n456), .ZN(n458) );
  XOR2_X1 U515 ( .A(G15GAT), .B(n458), .Z(G1326GAT) );
  NAND2_X1 U516 ( .A1(n497), .A2(n459), .ZN(n460) );
  XNOR2_X1 U517 ( .A(n460), .B(G22GAT), .ZN(G1327GAT) );
  XOR2_X1 U518 ( .A(KEYINPUT100), .B(KEYINPUT39), .Z(n469) );
  XNOR2_X1 U519 ( .A(KEYINPUT101), .B(KEYINPUT37), .ZN(n465) );
  XOR2_X1 U520 ( .A(KEYINPUT36), .B(n461), .Z(n591) );
  NOR2_X1 U521 ( .A1(n591), .A2(n541), .ZN(n463) );
  NAND2_X1 U522 ( .A1(n463), .A2(n462), .ZN(n464) );
  XNOR2_X1 U523 ( .A(n465), .B(n464), .ZN(n492) );
  NOR2_X1 U524 ( .A1(n466), .A2(n492), .ZN(n467) );
  XNOR2_X1 U525 ( .A(n467), .B(KEYINPUT38), .ZN(n477) );
  NAND2_X1 U526 ( .A1(n477), .A2(n573), .ZN(n468) );
  XNOR2_X1 U527 ( .A(n469), .B(n468), .ZN(n470) );
  XNOR2_X1 U528 ( .A(G29GAT), .B(n470), .ZN(G1328GAT) );
  NAND2_X1 U529 ( .A1(n477), .A2(n546), .ZN(n471) );
  XNOR2_X1 U530 ( .A(n471), .B(KEYINPUT102), .ZN(n472) );
  XNOR2_X1 U531 ( .A(G36GAT), .B(n472), .ZN(G1329GAT) );
  XNOR2_X1 U532 ( .A(G43GAT), .B(KEYINPUT104), .ZN(n476) );
  XOR2_X1 U533 ( .A(KEYINPUT103), .B(KEYINPUT40), .Z(n474) );
  NAND2_X1 U534 ( .A1(n564), .A2(n477), .ZN(n473) );
  XNOR2_X1 U535 ( .A(n474), .B(n473), .ZN(n475) );
  XNOR2_X1 U536 ( .A(n476), .B(n475), .ZN(G1330GAT) );
  NAND2_X1 U537 ( .A1(n497), .A2(n477), .ZN(n478) );
  XNOR2_X1 U538 ( .A(G50GAT), .B(n478), .ZN(G1331GAT) );
  XOR2_X1 U539 ( .A(KEYINPUT106), .B(KEYINPUT42), .Z(n482) );
  XOR2_X1 U540 ( .A(KEYINPUT41), .B(n583), .Z(n558) );
  INV_X1 U541 ( .A(n558), .ZN(n536) );
  INV_X1 U542 ( .A(n533), .ZN(n577) );
  NAND2_X1 U543 ( .A1(n536), .A2(n577), .ZN(n491) );
  NOR2_X1 U544 ( .A1(n491), .A2(n479), .ZN(n480) );
  XOR2_X1 U545 ( .A(KEYINPUT105), .B(n480), .Z(n487) );
  NAND2_X1 U546 ( .A1(n487), .A2(n573), .ZN(n481) );
  XNOR2_X1 U547 ( .A(n482), .B(n481), .ZN(n483) );
  XOR2_X1 U548 ( .A(G57GAT), .B(n483), .Z(G1332GAT) );
  XOR2_X1 U549 ( .A(G64GAT), .B(KEYINPUT107), .Z(n485) );
  NAND2_X1 U550 ( .A1(n487), .A2(n546), .ZN(n484) );
  XNOR2_X1 U551 ( .A(n485), .B(n484), .ZN(G1333GAT) );
  NAND2_X1 U552 ( .A1(n487), .A2(n564), .ZN(n486) );
  XNOR2_X1 U553 ( .A(n486), .B(G71GAT), .ZN(G1334GAT) );
  XOR2_X1 U554 ( .A(KEYINPUT108), .B(KEYINPUT43), .Z(n489) );
  NAND2_X1 U555 ( .A1(n487), .A2(n497), .ZN(n488) );
  XNOR2_X1 U556 ( .A(n489), .B(n488), .ZN(n490) );
  XNOR2_X1 U557 ( .A(G78GAT), .B(n490), .ZN(G1335GAT) );
  NOR2_X1 U558 ( .A1(n492), .A2(n491), .ZN(n493) );
  XOR2_X1 U559 ( .A(KEYINPUT109), .B(n493), .Z(n498) );
  NAND2_X1 U560 ( .A1(n498), .A2(n573), .ZN(n494) );
  XNOR2_X1 U561 ( .A(G85GAT), .B(n494), .ZN(G1336GAT) );
  NAND2_X1 U562 ( .A1(n498), .A2(n546), .ZN(n495) );
  XNOR2_X1 U563 ( .A(n495), .B(G92GAT), .ZN(G1337GAT) );
  NAND2_X1 U564 ( .A1(n498), .A2(n564), .ZN(n496) );
  XNOR2_X1 U565 ( .A(n496), .B(G99GAT), .ZN(G1338GAT) );
  XNOR2_X1 U566 ( .A(G106GAT), .B(KEYINPUT110), .ZN(n502) );
  XOR2_X1 U567 ( .A(KEYINPUT111), .B(KEYINPUT44), .Z(n500) );
  NAND2_X1 U568 ( .A1(n498), .A2(n497), .ZN(n499) );
  XNOR2_X1 U569 ( .A(n500), .B(n499), .ZN(n501) );
  XNOR2_X1 U570 ( .A(n502), .B(n501), .ZN(G1339GAT) );
  NOR2_X1 U571 ( .A1(n591), .A2(n588), .ZN(n503) );
  XNOR2_X1 U572 ( .A(n503), .B(KEYINPUT45), .ZN(n506) );
  INV_X1 U573 ( .A(n583), .ZN(n504) );
  NOR2_X1 U574 ( .A1(n519), .A2(n504), .ZN(n505) );
  NAND2_X1 U575 ( .A1(n506), .A2(n505), .ZN(n513) );
  NAND2_X1 U576 ( .A1(n533), .A2(n536), .ZN(n507) );
  XNOR2_X1 U577 ( .A(KEYINPUT46), .B(n507), .ZN(n508) );
  NAND2_X1 U578 ( .A1(n508), .A2(n588), .ZN(n509) );
  NOR2_X1 U579 ( .A1(n543), .A2(n509), .ZN(n510) );
  XOR2_X1 U580 ( .A(KEYINPUT47), .B(n510), .Z(n511) );
  XOR2_X1 U581 ( .A(n511), .B(KEYINPUT112), .Z(n512) );
  AND2_X1 U582 ( .A1(n513), .A2(n512), .ZN(n514) );
  XNOR2_X1 U583 ( .A(n514), .B(KEYINPUT48), .ZN(n548) );
  NOR2_X1 U584 ( .A1(n515), .A2(n548), .ZN(n516) );
  XNOR2_X1 U585 ( .A(n516), .B(KEYINPUT113), .ZN(n532) );
  NAND2_X1 U586 ( .A1(n564), .A2(n517), .ZN(n518) );
  NOR2_X1 U587 ( .A1(n532), .A2(n518), .ZN(n529) );
  NAND2_X1 U588 ( .A1(n519), .A2(n529), .ZN(n520) );
  XNOR2_X1 U589 ( .A(n520), .B(KEYINPUT114), .ZN(n521) );
  XNOR2_X1 U590 ( .A(G113GAT), .B(n521), .ZN(G1340GAT) );
  XOR2_X1 U591 ( .A(KEYINPUT116), .B(KEYINPUT49), .Z(n523) );
  NAND2_X1 U592 ( .A1(n529), .A2(n536), .ZN(n522) );
  XNOR2_X1 U593 ( .A(n523), .B(n522), .ZN(n525) );
  XOR2_X1 U594 ( .A(G120GAT), .B(KEYINPUT115), .Z(n524) );
  XNOR2_X1 U595 ( .A(n525), .B(n524), .ZN(G1341GAT) );
  XOR2_X1 U596 ( .A(KEYINPUT50), .B(KEYINPUT117), .Z(n527) );
  NAND2_X1 U597 ( .A1(n529), .A2(n541), .ZN(n526) );
  XNOR2_X1 U598 ( .A(n527), .B(n526), .ZN(n528) );
  XNOR2_X1 U599 ( .A(G127GAT), .B(n528), .ZN(G1342GAT) );
  XOR2_X1 U600 ( .A(G134GAT), .B(KEYINPUT51), .Z(n531) );
  NAND2_X1 U601 ( .A1(n529), .A2(n461), .ZN(n530) );
  XNOR2_X1 U602 ( .A(n531), .B(n530), .ZN(G1343GAT) );
  XNOR2_X1 U603 ( .A(G141GAT), .B(KEYINPUT118), .ZN(n535) );
  NOR2_X1 U604 ( .A1(n572), .A2(n532), .ZN(n544) );
  NAND2_X1 U605 ( .A1(n533), .A2(n544), .ZN(n534) );
  XNOR2_X1 U606 ( .A(n535), .B(n534), .ZN(G1344GAT) );
  XOR2_X1 U607 ( .A(KEYINPUT52), .B(KEYINPUT119), .Z(n538) );
  NAND2_X1 U608 ( .A1(n544), .A2(n536), .ZN(n537) );
  XNOR2_X1 U609 ( .A(n538), .B(n537), .ZN(n540) );
  XOR2_X1 U610 ( .A(G148GAT), .B(KEYINPUT53), .Z(n539) );
  XNOR2_X1 U611 ( .A(n540), .B(n539), .ZN(G1345GAT) );
  NAND2_X1 U612 ( .A1(n541), .A2(n544), .ZN(n542) );
  XNOR2_X1 U613 ( .A(n542), .B(G155GAT), .ZN(G1346GAT) );
  NAND2_X1 U614 ( .A1(n544), .A2(n543), .ZN(n545) );
  XNOR2_X1 U615 ( .A(n545), .B(G162GAT), .ZN(G1347GAT) );
  INV_X1 U616 ( .A(n546), .ZN(n547) );
  NOR2_X1 U617 ( .A1(n548), .A2(n547), .ZN(n549) );
  XNOR2_X1 U618 ( .A(n549), .B(KEYINPUT54), .ZN(n575) );
  AND2_X1 U619 ( .A1(n575), .A2(n550), .ZN(n552) );
  NAND2_X1 U620 ( .A1(n552), .A2(n551), .ZN(n553) );
  XNOR2_X1 U621 ( .A(KEYINPUT55), .B(n553), .ZN(n568) );
  NAND2_X1 U622 ( .A1(n568), .A2(n564), .ZN(n561) );
  NOR2_X1 U623 ( .A1(n554), .A2(n561), .ZN(n555) );
  XOR2_X1 U624 ( .A(G169GAT), .B(n555), .Z(G1348GAT) );
  XOR2_X1 U625 ( .A(KEYINPUT56), .B(KEYINPUT120), .Z(n557) );
  XNOR2_X1 U626 ( .A(G176GAT), .B(KEYINPUT57), .ZN(n556) );
  XNOR2_X1 U627 ( .A(n557), .B(n556), .ZN(n560) );
  NOR2_X1 U628 ( .A1(n558), .A2(n561), .ZN(n559) );
  XOR2_X1 U629 ( .A(n560), .B(n559), .Z(G1349GAT) );
  NOR2_X1 U630 ( .A1(n588), .A2(n561), .ZN(n563) );
  XNOR2_X1 U631 ( .A(G183GAT), .B(KEYINPUT121), .ZN(n562) );
  XNOR2_X1 U632 ( .A(n563), .B(n562), .ZN(G1350GAT) );
  INV_X1 U633 ( .A(n564), .ZN(n565) );
  NOR2_X1 U634 ( .A1(n566), .A2(n565), .ZN(n567) );
  AND2_X1 U635 ( .A1(n568), .A2(n567), .ZN(n570) );
  XNOR2_X1 U636 ( .A(KEYINPUT58), .B(KEYINPUT122), .ZN(n569) );
  XNOR2_X1 U637 ( .A(n570), .B(n569), .ZN(n571) );
  XOR2_X1 U638 ( .A(G190GAT), .B(n571), .Z(G1351GAT) );
  XNOR2_X1 U639 ( .A(KEYINPUT125), .B(KEYINPUT124), .ZN(n579) );
  NOR2_X1 U640 ( .A1(n573), .A2(n572), .ZN(n574) );
  AND2_X1 U641 ( .A1(n575), .A2(n574), .ZN(n576) );
  XNOR2_X1 U642 ( .A(n576), .B(KEYINPUT123), .ZN(n590) );
  NOR2_X1 U643 ( .A1(n590), .A2(n577), .ZN(n578) );
  XNOR2_X1 U644 ( .A(n579), .B(n578), .ZN(n580) );
  XOR2_X1 U645 ( .A(n580), .B(KEYINPUT59), .Z(n582) );
  XNOR2_X1 U646 ( .A(G197GAT), .B(KEYINPUT60), .ZN(n581) );
  XNOR2_X1 U647 ( .A(n582), .B(n581), .ZN(G1352GAT) );
  NOR2_X1 U648 ( .A1(n590), .A2(n583), .ZN(n587) );
  XOR2_X1 U649 ( .A(KEYINPUT126), .B(KEYINPUT61), .Z(n585) );
  XNOR2_X1 U650 ( .A(G204GAT), .B(KEYINPUT127), .ZN(n584) );
  XNOR2_X1 U651 ( .A(n585), .B(n584), .ZN(n586) );
  XNOR2_X1 U652 ( .A(n587), .B(n586), .ZN(G1353GAT) );
  NOR2_X1 U653 ( .A1(n588), .A2(n590), .ZN(n589) );
  XOR2_X1 U654 ( .A(G211GAT), .B(n589), .Z(G1354GAT) );
  NOR2_X1 U655 ( .A1(n591), .A2(n590), .ZN(n592) );
  XNOR2_X1 U656 ( .A(G218GAT), .B(n292), .ZN(G1355GAT) );
endmodule

