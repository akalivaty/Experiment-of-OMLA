//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 1 1 1 0 1 0 0 1 0 0 0 1 0 0 1 1 0 1 1 0 0 1 0 1 0 0 1 1 1 0 0 0 1 1 1 0 1 1 0 1 0 1 1 0 0 0 1 0 1 1 1 1 1 1 1 0 0 0 0 1 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:31:42 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n447, new_n451, new_n452, new_n453, new_n454, new_n457,
    new_n458, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n495, new_n496,
    new_n497, new_n498, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n517, new_n518, new_n519,
    new_n520, new_n521, new_n522, new_n523, new_n524, new_n527, new_n528,
    new_n529, new_n530, new_n531, new_n532, new_n533, new_n534, new_n535,
    new_n536, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n559,
    new_n560, new_n562, new_n563, new_n564, new_n565, new_n566, new_n567,
    new_n568, new_n569, new_n570, new_n571, new_n572, new_n573, new_n576,
    new_n577, new_n578, new_n580, new_n581, new_n582, new_n583, new_n584,
    new_n585, new_n586, new_n587, new_n588, new_n589, new_n590, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n619, new_n620, new_n623, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1197, new_n1198, new_n1199, new_n1200, new_n1201, new_n1202;
  BUF_X1    g000(.A(G452), .Z(G350));
  XNOR2_X1  g001(.A(KEYINPUT64), .B(G452), .ZN(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  XNOR2_X1  g009(.A(KEYINPUT65), .B(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  XOR2_X1   g014(.A(KEYINPUT66), .B(G57), .Z(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  AND2_X1   g016(.A1(G2072), .A2(G2078), .ZN(new_n442));
  NAND3_X1  g017(.A1(new_n442), .A2(G2084), .A3(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G219), .A2(G220), .A3(G218), .A4(G221), .ZN(new_n451));
  XOR2_X1   g026(.A(KEYINPUT67), .B(KEYINPUT2), .Z(new_n452));
  XNOR2_X1  g027(.A(new_n451), .B(new_n452), .ZN(new_n453));
  OR4_X1    g028(.A1(G235), .A2(G237), .A3(G238), .A4(G236), .ZN(new_n454));
  NOR2_X1   g029(.A1(new_n453), .A2(new_n454), .ZN(G325));
  INV_X1    g030(.A(G325), .ZN(G261));
  NAND2_X1  g031(.A1(new_n453), .A2(G2106), .ZN(new_n457));
  NAND2_X1  g032(.A1(new_n454), .A2(G567), .ZN(new_n458));
  AND2_X1   g033(.A1(new_n457), .A2(new_n458), .ZN(G319));
  INV_X1    g034(.A(G2105), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n460), .A2(G2104), .ZN(new_n461));
  INV_X1    g036(.A(KEYINPUT68), .ZN(new_n462));
  XNOR2_X1  g037(.A(new_n461), .B(new_n462), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n463), .A2(G101), .ZN(new_n464));
  INV_X1    g039(.A(G137), .ZN(new_n465));
  AND2_X1   g040(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n466));
  NOR2_X1   g041(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n467));
  NOR2_X1   g042(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  INV_X1    g043(.A(new_n468), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n469), .A2(new_n460), .ZN(new_n470));
  OAI21_X1  g045(.A(new_n464), .B1(new_n465), .B2(new_n470), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n469), .A2(G125), .ZN(new_n472));
  NAND2_X1  g047(.A1(G113), .A2(G2104), .ZN(new_n473));
  AOI21_X1  g048(.A(new_n460), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  NOR2_X1   g049(.A1(new_n471), .A2(new_n474), .ZN(G160));
  NOR2_X1   g050(.A1(new_n468), .A2(G2105), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n476), .A2(G136), .ZN(new_n477));
  NOR2_X1   g052(.A1(new_n468), .A2(new_n460), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n478), .A2(G124), .ZN(new_n479));
  OR2_X1    g054(.A1(G100), .A2(G2105), .ZN(new_n480));
  OAI211_X1 g055(.A(new_n480), .B(G2104), .C1(G112), .C2(new_n460), .ZN(new_n481));
  NAND3_X1  g056(.A1(new_n477), .A2(new_n479), .A3(new_n481), .ZN(new_n482));
  INV_X1    g057(.A(new_n482), .ZN(G162));
  OAI21_X1  g058(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n484));
  INV_X1    g059(.A(G114), .ZN(new_n485));
  AOI21_X1  g060(.A(new_n484), .B1(new_n485), .B2(G2105), .ZN(new_n486));
  OAI211_X1 g061(.A(G138), .B(new_n460), .C1(new_n466), .C2(new_n467), .ZN(new_n487));
  OR2_X1    g062(.A1(new_n487), .A2(KEYINPUT4), .ZN(new_n488));
  NAND2_X1  g063(.A1(new_n487), .A2(KEYINPUT4), .ZN(new_n489));
  AOI21_X1  g064(.A(new_n486), .B1(new_n488), .B2(new_n489), .ZN(new_n490));
  OAI211_X1 g065(.A(G126), .B(G2105), .C1(new_n466), .C2(new_n467), .ZN(new_n491));
  XOR2_X1   g066(.A(new_n491), .B(KEYINPUT69), .Z(new_n492));
  NAND2_X1  g067(.A1(new_n490), .A2(new_n492), .ZN(new_n493));
  INV_X1    g068(.A(new_n493), .ZN(G164));
  AND2_X1   g069(.A1(KEYINPUT5), .A2(G543), .ZN(new_n495));
  NOR2_X1   g070(.A1(KEYINPUT5), .A2(G543), .ZN(new_n496));
  NOR2_X1   g071(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  INV_X1    g072(.A(G62), .ZN(new_n498));
  NOR2_X1   g073(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  AND2_X1   g074(.A1(G75), .A2(G543), .ZN(new_n500));
  OAI21_X1  g075(.A(G651), .B1(new_n499), .B2(new_n500), .ZN(new_n501));
  INV_X1    g076(.A(G651), .ZN(new_n502));
  OAI21_X1  g077(.A(KEYINPUT70), .B1(new_n502), .B2(KEYINPUT6), .ZN(new_n503));
  INV_X1    g078(.A(KEYINPUT70), .ZN(new_n504));
  INV_X1    g079(.A(KEYINPUT6), .ZN(new_n505));
  NAND3_X1  g080(.A1(new_n504), .A2(new_n505), .A3(G651), .ZN(new_n506));
  AOI22_X1  g081(.A1(new_n503), .A2(new_n506), .B1(KEYINPUT6), .B2(new_n502), .ZN(new_n507));
  NAND3_X1  g082(.A1(new_n507), .A2(G50), .A3(G543), .ZN(new_n508));
  INV_X1    g083(.A(KEYINPUT5), .ZN(new_n509));
  INV_X1    g084(.A(G543), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  NAND2_X1  g086(.A1(KEYINPUT5), .A2(G543), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  NAND3_X1  g088(.A1(new_n507), .A2(G88), .A3(new_n513), .ZN(new_n514));
  NAND3_X1  g089(.A1(new_n501), .A2(new_n508), .A3(new_n514), .ZN(G303));
  INV_X1    g090(.A(G303), .ZN(G166));
  NAND3_X1  g091(.A1(new_n507), .A2(G89), .A3(new_n513), .ZN(new_n517));
  NAND3_X1  g092(.A1(new_n507), .A2(G51), .A3(G543), .ZN(new_n518));
  NAND3_X1  g093(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n519));
  XNOR2_X1  g094(.A(new_n519), .B(KEYINPUT7), .ZN(new_n520));
  OAI21_X1  g095(.A(KEYINPUT71), .B1(new_n495), .B2(new_n496), .ZN(new_n521));
  INV_X1    g096(.A(KEYINPUT71), .ZN(new_n522));
  NAND3_X1  g097(.A1(new_n511), .A2(new_n522), .A3(new_n512), .ZN(new_n523));
  NAND4_X1  g098(.A1(new_n521), .A2(new_n523), .A3(G63), .A4(G651), .ZN(new_n524));
  NAND4_X1  g099(.A1(new_n517), .A2(new_n518), .A3(new_n520), .A4(new_n524), .ZN(G286));
  INV_X1    g100(.A(G286), .ZN(G168));
  NAND2_X1  g101(.A1(new_n507), .A2(new_n513), .ZN(new_n527));
  XNOR2_X1  g102(.A(KEYINPUT72), .B(G90), .ZN(new_n528));
  NAND2_X1  g103(.A1(new_n503), .A2(new_n506), .ZN(new_n529));
  NAND2_X1  g104(.A1(new_n502), .A2(KEYINPUT6), .ZN(new_n530));
  NAND3_X1  g105(.A1(new_n529), .A2(G543), .A3(new_n530), .ZN(new_n531));
  INV_X1    g106(.A(G52), .ZN(new_n532));
  OAI22_X1  g107(.A1(new_n527), .A2(new_n528), .B1(new_n531), .B2(new_n532), .ZN(new_n533));
  NAND3_X1  g108(.A1(new_n521), .A2(new_n523), .A3(G64), .ZN(new_n534));
  NAND2_X1  g109(.A1(G77), .A2(G543), .ZN(new_n535));
  AOI21_X1  g110(.A(new_n502), .B1(new_n534), .B2(new_n535), .ZN(new_n536));
  NOR2_X1   g111(.A1(new_n533), .A2(new_n536), .ZN(G171));
  INV_X1    g112(.A(KEYINPUT74), .ZN(new_n538));
  NAND3_X1  g113(.A1(new_n521), .A2(new_n523), .A3(G56), .ZN(new_n539));
  NAND2_X1  g114(.A1(G68), .A2(G543), .ZN(new_n540));
  AND3_X1   g115(.A1(new_n539), .A2(KEYINPUT73), .A3(new_n540), .ZN(new_n541));
  AOI21_X1  g116(.A(KEYINPUT73), .B1(new_n539), .B2(new_n540), .ZN(new_n542));
  NOR3_X1   g117(.A1(new_n541), .A2(new_n542), .A3(new_n502), .ZN(new_n543));
  INV_X1    g118(.A(G81), .ZN(new_n544));
  INV_X1    g119(.A(G43), .ZN(new_n545));
  OAI22_X1  g120(.A1(new_n527), .A2(new_n544), .B1(new_n531), .B2(new_n545), .ZN(new_n546));
  OAI21_X1  g121(.A(new_n538), .B1(new_n543), .B2(new_n546), .ZN(new_n547));
  NAND2_X1  g122(.A1(new_n539), .A2(new_n540), .ZN(new_n548));
  INV_X1    g123(.A(KEYINPUT73), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  NAND3_X1  g125(.A1(new_n539), .A2(KEYINPUT73), .A3(new_n540), .ZN(new_n551));
  NAND3_X1  g126(.A1(new_n550), .A2(G651), .A3(new_n551), .ZN(new_n552));
  INV_X1    g127(.A(new_n546), .ZN(new_n553));
  NAND3_X1  g128(.A1(new_n552), .A2(KEYINPUT74), .A3(new_n553), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n547), .A2(new_n554), .ZN(new_n555));
  INV_X1    g130(.A(new_n555), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n556), .A2(G860), .ZN(G153));
  NAND4_X1  g132(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g133(.A1(G1), .A2(G3), .ZN(new_n559));
  XNOR2_X1  g134(.A(new_n559), .B(KEYINPUT8), .ZN(new_n560));
  NAND4_X1  g135(.A1(G319), .A2(G483), .A3(G661), .A4(new_n560), .ZN(G188));
  NAND4_X1  g136(.A1(new_n529), .A2(G53), .A3(G543), .A4(new_n530), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n562), .A2(KEYINPUT9), .ZN(new_n563));
  INV_X1    g138(.A(KEYINPUT9), .ZN(new_n564));
  NAND4_X1  g139(.A1(new_n507), .A2(new_n564), .A3(G53), .A4(G543), .ZN(new_n565));
  NAND2_X1  g140(.A1(new_n563), .A2(new_n565), .ZN(new_n566));
  INV_X1    g141(.A(G65), .ZN(new_n567));
  AOI21_X1  g142(.A(new_n567), .B1(new_n511), .B2(new_n512), .ZN(new_n568));
  AND2_X1   g143(.A1(G78), .A2(G543), .ZN(new_n569));
  OAI21_X1  g144(.A(G651), .B1(new_n568), .B2(new_n569), .ZN(new_n570));
  NAND4_X1  g145(.A1(new_n529), .A2(G91), .A3(new_n530), .A4(new_n513), .ZN(new_n571));
  NAND2_X1  g146(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  INV_X1    g147(.A(new_n572), .ZN(new_n573));
  NAND2_X1  g148(.A1(new_n566), .A2(new_n573), .ZN(G299));
  INV_X1    g149(.A(G171), .ZN(G301));
  NAND4_X1  g150(.A1(new_n529), .A2(G87), .A3(new_n530), .A4(new_n513), .ZN(new_n576));
  NAND4_X1  g151(.A1(new_n529), .A2(G49), .A3(G543), .A4(new_n530), .ZN(new_n577));
  AOI21_X1  g152(.A(G74), .B1(new_n521), .B2(new_n523), .ZN(new_n578));
  OAI211_X1 g153(.A(new_n576), .B(new_n577), .C1(new_n578), .C2(new_n502), .ZN(G288));
  NAND4_X1  g154(.A1(new_n529), .A2(G86), .A3(new_n530), .A4(new_n513), .ZN(new_n580));
  INV_X1    g155(.A(KEYINPUT76), .ZN(new_n581));
  XNOR2_X1  g156(.A(new_n580), .B(new_n581), .ZN(new_n582));
  INV_X1    g157(.A(G61), .ZN(new_n583));
  OAI21_X1  g158(.A(KEYINPUT75), .B1(new_n497), .B2(new_n583), .ZN(new_n584));
  INV_X1    g159(.A(KEYINPUT75), .ZN(new_n585));
  NAND3_X1  g160(.A1(new_n513), .A2(new_n585), .A3(G61), .ZN(new_n586));
  NAND2_X1  g161(.A1(G73), .A2(G543), .ZN(new_n587));
  NAND3_X1  g162(.A1(new_n584), .A2(new_n586), .A3(new_n587), .ZN(new_n588));
  INV_X1    g163(.A(new_n531), .ZN(new_n589));
  AOI22_X1  g164(.A1(new_n588), .A2(G651), .B1(new_n589), .B2(G48), .ZN(new_n590));
  NAND2_X1  g165(.A1(new_n582), .A2(new_n590), .ZN(G305));
  XOR2_X1   g166(.A(KEYINPUT78), .B(G85), .Z(new_n592));
  NAND3_X1  g167(.A1(new_n507), .A2(new_n513), .A3(new_n592), .ZN(new_n593));
  INV_X1    g168(.A(G47), .ZN(new_n594));
  OAI21_X1  g169(.A(new_n593), .B1(new_n594), .B2(new_n531), .ZN(new_n595));
  NAND3_X1  g170(.A1(new_n521), .A2(new_n523), .A3(G60), .ZN(new_n596));
  NAND2_X1  g171(.A1(G72), .A2(G543), .ZN(new_n597));
  NAND2_X1  g172(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  NAND2_X1  g173(.A1(new_n598), .A2(G651), .ZN(new_n599));
  NAND2_X1  g174(.A1(new_n599), .A2(KEYINPUT77), .ZN(new_n600));
  INV_X1    g175(.A(KEYINPUT77), .ZN(new_n601));
  NAND3_X1  g176(.A1(new_n598), .A2(new_n601), .A3(G651), .ZN(new_n602));
  AOI21_X1  g177(.A(new_n595), .B1(new_n600), .B2(new_n602), .ZN(new_n603));
  INV_X1    g178(.A(new_n603), .ZN(G290));
  NAND2_X1  g179(.A1(G301), .A2(G868), .ZN(new_n605));
  NAND4_X1  g180(.A1(new_n529), .A2(G92), .A3(new_n530), .A4(new_n513), .ZN(new_n606));
  XNOR2_X1  g181(.A(new_n606), .B(KEYINPUT10), .ZN(new_n607));
  OAI21_X1  g182(.A(G66), .B1(new_n495), .B2(new_n496), .ZN(new_n608));
  NAND2_X1  g183(.A1(G79), .A2(G543), .ZN(new_n609));
  NAND2_X1  g184(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  OAI21_X1  g185(.A(G651), .B1(new_n610), .B2(KEYINPUT79), .ZN(new_n611));
  INV_X1    g186(.A(KEYINPUT79), .ZN(new_n612));
  AOI21_X1  g187(.A(new_n612), .B1(new_n608), .B2(new_n609), .ZN(new_n613));
  INV_X1    g188(.A(G54), .ZN(new_n614));
  OAI22_X1  g189(.A1(new_n611), .A2(new_n613), .B1(new_n614), .B2(new_n531), .ZN(new_n615));
  NOR2_X1   g190(.A1(new_n607), .A2(new_n615), .ZN(new_n616));
  OAI21_X1  g191(.A(new_n605), .B1(G868), .B2(new_n616), .ZN(G284));
  OAI21_X1  g192(.A(new_n605), .B1(G868), .B2(new_n616), .ZN(G321));
  NAND2_X1  g193(.A1(G286), .A2(G868), .ZN(new_n619));
  AOI21_X1  g194(.A(new_n572), .B1(new_n563), .B2(new_n565), .ZN(new_n620));
  OAI21_X1  g195(.A(new_n619), .B1(new_n620), .B2(G868), .ZN(G297));
  OAI21_X1  g196(.A(new_n619), .B1(new_n620), .B2(G868), .ZN(G280));
  INV_X1    g197(.A(G559), .ZN(new_n623));
  OAI21_X1  g198(.A(new_n616), .B1(new_n623), .B2(G860), .ZN(G148));
  INV_X1    g199(.A(KEYINPUT81), .ZN(new_n625));
  NAND2_X1  g200(.A1(new_n616), .A2(new_n623), .ZN(new_n626));
  XNOR2_X1  g201(.A(new_n626), .B(KEYINPUT80), .ZN(new_n627));
  AOI21_X1  g202(.A(new_n625), .B1(new_n627), .B2(G868), .ZN(new_n628));
  OAI21_X1  g203(.A(new_n628), .B1(G868), .B2(new_n556), .ZN(new_n629));
  NAND3_X1  g204(.A1(new_n627), .A2(new_n625), .A3(G868), .ZN(new_n630));
  AND2_X1   g205(.A1(new_n629), .A2(new_n630), .ZN(G323));
  XNOR2_X1  g206(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g207(.A1(new_n478), .A2(G123), .ZN(new_n633));
  NOR2_X1   g208(.A1(new_n460), .A2(G111), .ZN(new_n634));
  OAI21_X1  g209(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n635));
  OAI21_X1  g210(.A(new_n633), .B1(new_n634), .B2(new_n635), .ZN(new_n636));
  AOI21_X1  g211(.A(new_n636), .B1(G135), .B2(new_n476), .ZN(new_n637));
  XNOR2_X1  g212(.A(new_n637), .B(KEYINPUT82), .ZN(new_n638));
  XOR2_X1   g213(.A(new_n638), .B(G2096), .Z(new_n639));
  NAND2_X1  g214(.A1(new_n463), .A2(new_n469), .ZN(new_n640));
  XNOR2_X1  g215(.A(new_n640), .B(KEYINPUT12), .ZN(new_n641));
  XNOR2_X1  g216(.A(new_n641), .B(KEYINPUT13), .ZN(new_n642));
  XNOR2_X1  g217(.A(new_n642), .B(G2100), .ZN(new_n643));
  NAND2_X1  g218(.A1(new_n639), .A2(new_n643), .ZN(G156));
  XNOR2_X1  g219(.A(G2427), .B(G2438), .ZN(new_n645));
  XNOR2_X1  g220(.A(new_n645), .B(G2430), .ZN(new_n646));
  XNOR2_X1  g221(.A(KEYINPUT15), .B(G2435), .ZN(new_n647));
  OR2_X1    g222(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  NAND2_X1  g223(.A1(new_n646), .A2(new_n647), .ZN(new_n649));
  NAND3_X1  g224(.A1(new_n648), .A2(new_n649), .A3(KEYINPUT14), .ZN(new_n650));
  XOR2_X1   g225(.A(G1341), .B(G1348), .Z(new_n651));
  XNOR2_X1  g226(.A(G2443), .B(G2446), .ZN(new_n652));
  XNOR2_X1  g227(.A(new_n651), .B(new_n652), .ZN(new_n653));
  XNOR2_X1  g228(.A(new_n650), .B(new_n653), .ZN(new_n654));
  XOR2_X1   g229(.A(G2451), .B(G2454), .Z(new_n655));
  XNOR2_X1  g230(.A(KEYINPUT83), .B(KEYINPUT16), .ZN(new_n656));
  XNOR2_X1  g231(.A(new_n655), .B(new_n656), .ZN(new_n657));
  OR2_X1    g232(.A1(new_n654), .A2(new_n657), .ZN(new_n658));
  NAND2_X1  g233(.A1(new_n654), .A2(new_n657), .ZN(new_n659));
  AND3_X1   g234(.A1(new_n658), .A2(G14), .A3(new_n659), .ZN(G401));
  XOR2_X1   g235(.A(G2067), .B(G2678), .Z(new_n661));
  XNOR2_X1  g236(.A(new_n661), .B(KEYINPUT84), .ZN(new_n662));
  NOR2_X1   g237(.A1(G2072), .A2(G2078), .ZN(new_n663));
  NOR2_X1   g238(.A1(new_n442), .A2(new_n663), .ZN(new_n664));
  XOR2_X1   g239(.A(G2084), .B(G2090), .Z(new_n665));
  INV_X1    g240(.A(new_n665), .ZN(new_n666));
  NOR3_X1   g241(.A1(new_n662), .A2(new_n664), .A3(new_n666), .ZN(new_n667));
  XNOR2_X1  g242(.A(new_n667), .B(KEYINPUT18), .ZN(new_n668));
  NAND2_X1  g243(.A1(new_n662), .A2(new_n664), .ZN(new_n669));
  XNOR2_X1  g244(.A(new_n664), .B(KEYINPUT17), .ZN(new_n670));
  OAI211_X1 g245(.A(new_n669), .B(new_n666), .C1(new_n662), .C2(new_n670), .ZN(new_n671));
  NAND3_X1  g246(.A1(new_n662), .A2(new_n665), .A3(new_n670), .ZN(new_n672));
  NAND3_X1  g247(.A1(new_n668), .A2(new_n671), .A3(new_n672), .ZN(new_n673));
  XOR2_X1   g248(.A(G2096), .B(G2100), .Z(new_n674));
  XNOR2_X1  g249(.A(new_n673), .B(new_n674), .ZN(G227));
  XNOR2_X1  g250(.A(G1991), .B(G1996), .ZN(new_n676));
  INV_X1    g251(.A(new_n676), .ZN(new_n677));
  XNOR2_X1  g252(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n678));
  XNOR2_X1  g253(.A(new_n678), .B(KEYINPUT89), .ZN(new_n679));
  XOR2_X1   g254(.A(G1971), .B(G1976), .Z(new_n680));
  XNOR2_X1  g255(.A(KEYINPUT85), .B(KEYINPUT19), .ZN(new_n681));
  XNOR2_X1  g256(.A(new_n680), .B(new_n681), .ZN(new_n682));
  XOR2_X1   g257(.A(G1961), .B(G1966), .Z(new_n683));
  XNOR2_X1  g258(.A(new_n683), .B(KEYINPUT87), .ZN(new_n684));
  XNOR2_X1  g259(.A(G1956), .B(G2474), .ZN(new_n685));
  XNOR2_X1  g260(.A(new_n685), .B(KEYINPUT86), .ZN(new_n686));
  NAND3_X1  g261(.A1(new_n682), .A2(new_n684), .A3(new_n686), .ZN(new_n687));
  OAI21_X1  g262(.A(new_n687), .B1(new_n686), .B2(new_n684), .ZN(new_n688));
  INV_X1    g263(.A(KEYINPUT88), .ZN(new_n689));
  NAND2_X1  g264(.A1(new_n682), .A2(new_n689), .ZN(new_n690));
  XOR2_X1   g265(.A(new_n688), .B(new_n690), .Z(new_n691));
  NAND2_X1  g266(.A1(new_n684), .A2(new_n686), .ZN(new_n692));
  NOR2_X1   g267(.A1(new_n692), .A2(new_n682), .ZN(new_n693));
  XOR2_X1   g268(.A(new_n693), .B(KEYINPUT20), .Z(new_n694));
  NAND2_X1  g269(.A1(new_n691), .A2(new_n694), .ZN(new_n695));
  INV_X1    g270(.A(G1981), .ZN(new_n696));
  XNOR2_X1  g271(.A(new_n695), .B(new_n696), .ZN(new_n697));
  AND2_X1   g272(.A1(new_n697), .A2(G1986), .ZN(new_n698));
  NOR2_X1   g273(.A1(new_n697), .A2(G1986), .ZN(new_n699));
  OAI21_X1  g274(.A(new_n679), .B1(new_n698), .B2(new_n699), .ZN(new_n700));
  INV_X1    g275(.A(new_n700), .ZN(new_n701));
  NOR3_X1   g276(.A1(new_n698), .A2(new_n699), .A3(new_n679), .ZN(new_n702));
  OAI21_X1  g277(.A(new_n677), .B1(new_n701), .B2(new_n702), .ZN(new_n703));
  INV_X1    g278(.A(new_n702), .ZN(new_n704));
  NAND3_X1  g279(.A1(new_n704), .A2(new_n676), .A3(new_n700), .ZN(new_n705));
  NAND2_X1  g280(.A1(new_n703), .A2(new_n705), .ZN(G229));
  NOR2_X1   g281(.A1(G16), .A2(G23), .ZN(new_n707));
  OR2_X1    g282(.A1(G288), .A2(KEYINPUT92), .ZN(new_n708));
  NAND2_X1  g283(.A1(G288), .A2(KEYINPUT92), .ZN(new_n709));
  AND2_X1   g284(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  AOI21_X1  g285(.A(new_n707), .B1(new_n710), .B2(G16), .ZN(new_n711));
  XOR2_X1   g286(.A(KEYINPUT33), .B(G1976), .Z(new_n712));
  XNOR2_X1  g287(.A(new_n711), .B(new_n712), .ZN(new_n713));
  INV_X1    g288(.A(G16), .ZN(new_n714));
  NAND2_X1  g289(.A1(new_n714), .A2(G6), .ZN(new_n715));
  INV_X1    g290(.A(G305), .ZN(new_n716));
  OAI21_X1  g291(.A(new_n715), .B1(new_n716), .B2(new_n714), .ZN(new_n717));
  XNOR2_X1  g292(.A(KEYINPUT32), .B(G1981), .ZN(new_n718));
  NOR2_X1   g293(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  AND2_X1   g294(.A1(new_n717), .A2(new_n718), .ZN(new_n720));
  NAND2_X1  g295(.A1(new_n714), .A2(G22), .ZN(new_n721));
  OAI21_X1  g296(.A(new_n721), .B1(G166), .B2(new_n714), .ZN(new_n722));
  XNOR2_X1  g297(.A(new_n722), .B(G1971), .ZN(new_n723));
  NOR4_X1   g298(.A1(new_n713), .A2(new_n719), .A3(new_n720), .A4(new_n723), .ZN(new_n724));
  INV_X1    g299(.A(KEYINPUT34), .ZN(new_n725));
  NAND2_X1  g300(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  NAND2_X1  g301(.A1(new_n714), .A2(G24), .ZN(new_n727));
  OAI21_X1  g302(.A(new_n727), .B1(new_n603), .B2(new_n714), .ZN(new_n728));
  XNOR2_X1  g303(.A(new_n728), .B(KEYINPUT91), .ZN(new_n729));
  XNOR2_X1  g304(.A(new_n729), .B(G1986), .ZN(new_n730));
  NAND2_X1  g305(.A1(new_n726), .A2(new_n730), .ZN(new_n731));
  INV_X1    g306(.A(G29), .ZN(new_n732));
  NAND2_X1  g307(.A1(new_n732), .A2(G25), .ZN(new_n733));
  NAND2_X1  g308(.A1(new_n478), .A2(G119), .ZN(new_n734));
  INV_X1    g309(.A(G131), .ZN(new_n735));
  OAI21_X1  g310(.A(new_n734), .B1(new_n735), .B2(new_n470), .ZN(new_n736));
  OR2_X1    g311(.A1(G95), .A2(G2105), .ZN(new_n737));
  OAI211_X1 g312(.A(new_n737), .B(G2104), .C1(G107), .C2(new_n460), .ZN(new_n738));
  XNOR2_X1  g313(.A(new_n738), .B(KEYINPUT90), .ZN(new_n739));
  NOR2_X1   g314(.A1(new_n736), .A2(new_n739), .ZN(new_n740));
  OAI21_X1  g315(.A(new_n733), .B1(new_n740), .B2(new_n732), .ZN(new_n741));
  XNOR2_X1  g316(.A(KEYINPUT35), .B(G1991), .ZN(new_n742));
  XOR2_X1   g317(.A(new_n741), .B(new_n742), .Z(new_n743));
  OAI21_X1  g318(.A(new_n743), .B1(new_n724), .B2(new_n725), .ZN(new_n744));
  NOR2_X1   g319(.A1(new_n731), .A2(new_n744), .ZN(new_n745));
  XNOR2_X1  g320(.A(new_n745), .B(KEYINPUT36), .ZN(new_n746));
  NOR2_X1   g321(.A1(new_n556), .A2(new_n714), .ZN(new_n747));
  AOI21_X1  g322(.A(new_n747), .B1(new_n714), .B2(G19), .ZN(new_n748));
  XOR2_X1   g323(.A(KEYINPUT94), .B(G1341), .Z(new_n749));
  NAND2_X1  g324(.A1(new_n714), .A2(G20), .ZN(new_n750));
  XOR2_X1   g325(.A(new_n750), .B(KEYINPUT23), .Z(new_n751));
  AOI21_X1  g326(.A(new_n751), .B1(G299), .B2(G16), .ZN(new_n752));
  XNOR2_X1  g327(.A(new_n752), .B(G1956), .ZN(new_n753));
  NAND2_X1  g328(.A1(new_n732), .A2(G35), .ZN(new_n754));
  OAI21_X1  g329(.A(new_n754), .B1(G162), .B2(new_n732), .ZN(new_n755));
  XOR2_X1   g330(.A(new_n755), .B(KEYINPUT29), .Z(new_n756));
  INV_X1    g331(.A(G2090), .ZN(new_n757));
  OAI21_X1  g332(.A(new_n753), .B1(new_n756), .B2(new_n757), .ZN(new_n758));
  AOI22_X1  g333(.A1(new_n748), .A2(new_n749), .B1(new_n758), .B2(KEYINPUT102), .ZN(new_n759));
  OAI21_X1  g334(.A(new_n759), .B1(new_n748), .B2(new_n749), .ZN(new_n760));
  INV_X1    g335(.A(G34), .ZN(new_n761));
  AOI21_X1  g336(.A(G29), .B1(new_n761), .B2(KEYINPUT24), .ZN(new_n762));
  OAI21_X1  g337(.A(new_n762), .B1(KEYINPUT24), .B2(new_n761), .ZN(new_n763));
  INV_X1    g338(.A(G160), .ZN(new_n764));
  OAI21_X1  g339(.A(new_n763), .B1(new_n764), .B2(new_n732), .ZN(new_n765));
  INV_X1    g340(.A(G2084), .ZN(new_n766));
  NAND2_X1  g341(.A1(new_n732), .A2(G33), .ZN(new_n767));
  AND2_X1   g342(.A1(new_n469), .A2(G127), .ZN(new_n768));
  AND2_X1   g343(.A1(G115), .A2(G2104), .ZN(new_n769));
  OAI21_X1  g344(.A(G2105), .B1(new_n768), .B2(new_n769), .ZN(new_n770));
  INV_X1    g345(.A(KEYINPUT25), .ZN(new_n771));
  NAND2_X1  g346(.A1(G103), .A2(G2104), .ZN(new_n772));
  OAI21_X1  g347(.A(new_n771), .B1(new_n772), .B2(G2105), .ZN(new_n773));
  NAND4_X1  g348(.A1(new_n460), .A2(KEYINPUT25), .A3(G103), .A4(G2104), .ZN(new_n774));
  AOI22_X1  g349(.A1(new_n476), .A2(G139), .B1(new_n773), .B2(new_n774), .ZN(new_n775));
  AND2_X1   g350(.A1(new_n770), .A2(new_n775), .ZN(new_n776));
  OAI21_X1  g351(.A(new_n767), .B1(new_n776), .B2(new_n732), .ZN(new_n777));
  OAI22_X1  g352(.A1(new_n765), .A2(new_n766), .B1(G2072), .B2(new_n777), .ZN(new_n778));
  AOI21_X1  g353(.A(new_n778), .B1(G2072), .B2(new_n777), .ZN(new_n779));
  XNOR2_X1  g354(.A(KEYINPUT27), .B(G1996), .ZN(new_n780));
  XNOR2_X1  g355(.A(new_n780), .B(KEYINPUT96), .ZN(new_n781));
  AND2_X1   g356(.A1(new_n732), .A2(G32), .ZN(new_n782));
  AOI22_X1  g357(.A1(G105), .A2(new_n463), .B1(new_n476), .B2(G141), .ZN(new_n783));
  NAND3_X1  g358(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n784));
  XNOR2_X1  g359(.A(new_n784), .B(KEYINPUT26), .ZN(new_n785));
  AOI21_X1  g360(.A(new_n785), .B1(G129), .B2(new_n478), .ZN(new_n786));
  NAND2_X1  g361(.A1(new_n783), .A2(new_n786), .ZN(new_n787));
  INV_X1    g362(.A(KEYINPUT95), .ZN(new_n788));
  NAND2_X1  g363(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  NAND3_X1  g364(.A1(new_n783), .A2(KEYINPUT95), .A3(new_n786), .ZN(new_n790));
  NAND2_X1  g365(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  AOI21_X1  g366(.A(new_n782), .B1(new_n791), .B2(G29), .ZN(new_n792));
  INV_X1    g367(.A(new_n792), .ZN(new_n793));
  OAI21_X1  g368(.A(new_n779), .B1(new_n781), .B2(new_n793), .ZN(new_n794));
  XNOR2_X1  g369(.A(new_n794), .B(KEYINPUT97), .ZN(new_n795));
  NAND2_X1  g370(.A1(new_n714), .A2(G5), .ZN(new_n796));
  OAI21_X1  g371(.A(new_n796), .B1(G171), .B2(new_n714), .ZN(new_n797));
  XNOR2_X1  g372(.A(new_n797), .B(KEYINPUT100), .ZN(new_n798));
  INV_X1    g373(.A(G1961), .ZN(new_n799));
  XNOR2_X1  g374(.A(new_n798), .B(new_n799), .ZN(new_n800));
  NAND2_X1  g375(.A1(new_n732), .A2(G27), .ZN(new_n801));
  XNOR2_X1  g376(.A(new_n801), .B(KEYINPUT101), .ZN(new_n802));
  AOI21_X1  g377(.A(new_n802), .B1(new_n493), .B2(G29), .ZN(new_n803));
  XNOR2_X1  g378(.A(new_n803), .B(G2078), .ZN(new_n804));
  NAND2_X1  g379(.A1(new_n732), .A2(G26), .ZN(new_n805));
  XNOR2_X1  g380(.A(new_n805), .B(KEYINPUT28), .ZN(new_n806));
  NAND2_X1  g381(.A1(new_n476), .A2(G140), .ZN(new_n807));
  NAND2_X1  g382(.A1(new_n478), .A2(G128), .ZN(new_n808));
  OR2_X1    g383(.A1(G104), .A2(G2105), .ZN(new_n809));
  OAI211_X1 g384(.A(new_n809), .B(G2104), .C1(G116), .C2(new_n460), .ZN(new_n810));
  NAND3_X1  g385(.A1(new_n807), .A2(new_n808), .A3(new_n810), .ZN(new_n811));
  INV_X1    g386(.A(new_n811), .ZN(new_n812));
  OAI21_X1  g387(.A(new_n806), .B1(new_n812), .B2(new_n732), .ZN(new_n813));
  INV_X1    g388(.A(G2067), .ZN(new_n814));
  XNOR2_X1  g389(.A(new_n813), .B(new_n814), .ZN(new_n815));
  XNOR2_X1  g390(.A(KEYINPUT31), .B(G11), .ZN(new_n816));
  XOR2_X1   g391(.A(KEYINPUT99), .B(G28), .Z(new_n817));
  NOR2_X1   g392(.A1(new_n817), .A2(KEYINPUT30), .ZN(new_n818));
  NAND2_X1  g393(.A1(new_n817), .A2(KEYINPUT30), .ZN(new_n819));
  NAND2_X1  g394(.A1(new_n819), .A2(new_n732), .ZN(new_n820));
  OAI221_X1 g395(.A(new_n816), .B1(new_n818), .B2(new_n820), .C1(new_n638), .C2(new_n732), .ZN(new_n821));
  AOI21_X1  g396(.A(new_n821), .B1(new_n766), .B2(new_n765), .ZN(new_n822));
  NAND2_X1  g397(.A1(new_n756), .A2(new_n757), .ZN(new_n823));
  NAND2_X1  g398(.A1(new_n793), .A2(new_n781), .ZN(new_n824));
  AND4_X1   g399(.A1(new_n815), .A2(new_n822), .A3(new_n823), .A4(new_n824), .ZN(new_n825));
  NAND4_X1  g400(.A1(new_n795), .A2(new_n800), .A3(new_n804), .A4(new_n825), .ZN(new_n826));
  NAND2_X1  g401(.A1(new_n714), .A2(G21), .ZN(new_n827));
  OAI21_X1  g402(.A(new_n827), .B1(G168), .B2(new_n714), .ZN(new_n828));
  XNOR2_X1  g403(.A(new_n828), .B(KEYINPUT98), .ZN(new_n829));
  INV_X1    g404(.A(G1966), .ZN(new_n830));
  XNOR2_X1  g405(.A(new_n829), .B(new_n830), .ZN(new_n831));
  NAND2_X1  g406(.A1(new_n714), .A2(G4), .ZN(new_n832));
  OAI21_X1  g407(.A(new_n832), .B1(new_n616), .B2(new_n714), .ZN(new_n833));
  XOR2_X1   g408(.A(KEYINPUT93), .B(G1348), .Z(new_n834));
  XNOR2_X1  g409(.A(new_n833), .B(new_n834), .ZN(new_n835));
  OAI211_X1 g410(.A(new_n831), .B(new_n835), .C1(KEYINPUT102), .C2(new_n758), .ZN(new_n836));
  NOR4_X1   g411(.A1(new_n746), .A2(new_n760), .A3(new_n826), .A4(new_n836), .ZN(G311));
  OR4_X1    g412(.A1(new_n746), .A2(new_n760), .A3(new_n826), .A4(new_n836), .ZN(G150));
  INV_X1    g413(.A(G93), .ZN(new_n839));
  INV_X1    g414(.A(G55), .ZN(new_n840));
  OAI22_X1  g415(.A1(new_n527), .A2(new_n839), .B1(new_n531), .B2(new_n840), .ZN(new_n841));
  NAND3_X1  g416(.A1(new_n521), .A2(new_n523), .A3(G67), .ZN(new_n842));
  INV_X1    g417(.A(G80), .ZN(new_n843));
  OAI21_X1  g418(.A(new_n842), .B1(new_n843), .B2(new_n510), .ZN(new_n844));
  AOI21_X1  g419(.A(new_n841), .B1(new_n844), .B2(G651), .ZN(new_n845));
  NAND3_X1  g420(.A1(new_n845), .A2(new_n552), .A3(new_n553), .ZN(new_n846));
  INV_X1    g421(.A(new_n846), .ZN(new_n847));
  INV_X1    g422(.A(new_n845), .ZN(new_n848));
  AOI21_X1  g423(.A(new_n847), .B1(new_n555), .B2(new_n848), .ZN(new_n849));
  XNOR2_X1  g424(.A(new_n849), .B(KEYINPUT38), .ZN(new_n850));
  INV_X1    g425(.A(new_n616), .ZN(new_n851));
  NOR2_X1   g426(.A1(new_n851), .A2(new_n623), .ZN(new_n852));
  XNOR2_X1  g427(.A(new_n850), .B(new_n852), .ZN(new_n853));
  INV_X1    g428(.A(KEYINPUT39), .ZN(new_n854));
  NOR2_X1   g429(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  XOR2_X1   g430(.A(new_n855), .B(KEYINPUT103), .Z(new_n856));
  AOI21_X1  g431(.A(G860), .B1(new_n853), .B2(new_n854), .ZN(new_n857));
  NAND2_X1  g432(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  NAND2_X1  g433(.A1(new_n848), .A2(G860), .ZN(new_n859));
  XOR2_X1   g434(.A(new_n859), .B(KEYINPUT37), .Z(new_n860));
  NAND2_X1  g435(.A1(new_n858), .A2(new_n860), .ZN(G145));
  XNOR2_X1  g436(.A(G164), .B(new_n776), .ZN(new_n862));
  XNOR2_X1  g437(.A(new_n641), .B(new_n740), .ZN(new_n863));
  XOR2_X1   g438(.A(new_n862), .B(new_n863), .Z(new_n864));
  NOR2_X1   g439(.A1(new_n791), .A2(new_n811), .ZN(new_n865));
  INV_X1    g440(.A(new_n865), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n476), .A2(G142), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n478), .A2(G130), .ZN(new_n868));
  OR2_X1    g443(.A1(G106), .A2(G2105), .ZN(new_n869));
  OAI211_X1 g444(.A(new_n869), .B(G2104), .C1(G118), .C2(new_n460), .ZN(new_n870));
  NAND3_X1  g445(.A1(new_n867), .A2(new_n868), .A3(new_n870), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n791), .A2(new_n811), .ZN(new_n872));
  NAND3_X1  g447(.A1(new_n866), .A2(new_n871), .A3(new_n872), .ZN(new_n873));
  INV_X1    g448(.A(new_n873), .ZN(new_n874));
  AOI21_X1  g449(.A(new_n871), .B1(new_n866), .B2(new_n872), .ZN(new_n875));
  OAI21_X1  g450(.A(new_n864), .B1(new_n874), .B2(new_n875), .ZN(new_n876));
  XNOR2_X1  g451(.A(new_n862), .B(new_n863), .ZN(new_n877));
  INV_X1    g452(.A(new_n875), .ZN(new_n878));
  NAND3_X1  g453(.A1(new_n877), .A2(new_n878), .A3(new_n873), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n876), .A2(new_n879), .ZN(new_n880));
  XNOR2_X1  g455(.A(new_n638), .B(new_n764), .ZN(new_n881));
  XNOR2_X1  g456(.A(new_n881), .B(G162), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n880), .A2(new_n882), .ZN(new_n883));
  INV_X1    g458(.A(G37), .ZN(new_n884));
  XNOR2_X1  g459(.A(new_n881), .B(new_n482), .ZN(new_n885));
  NAND3_X1  g460(.A1(new_n885), .A2(new_n879), .A3(new_n876), .ZN(new_n886));
  NAND3_X1  g461(.A1(new_n883), .A2(new_n884), .A3(new_n886), .ZN(new_n887));
  INV_X1    g462(.A(KEYINPUT104), .ZN(new_n888));
  XNOR2_X1  g463(.A(new_n887), .B(new_n888), .ZN(new_n889));
  XNOR2_X1  g464(.A(KEYINPUT105), .B(KEYINPUT40), .ZN(new_n890));
  XNOR2_X1  g465(.A(new_n889), .B(new_n890), .ZN(G395));
  AND3_X1   g466(.A1(new_n552), .A2(KEYINPUT74), .A3(new_n553), .ZN(new_n892));
  AOI21_X1  g467(.A(KEYINPUT74), .B1(new_n552), .B2(new_n553), .ZN(new_n893));
  OAI21_X1  g468(.A(new_n848), .B1(new_n892), .B2(new_n893), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n894), .A2(new_n846), .ZN(new_n895));
  OR2_X1    g470(.A1(new_n627), .A2(new_n895), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n627), .A2(new_n895), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  AOI22_X1  g473(.A1(new_n513), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n899));
  AOI21_X1  g474(.A(new_n502), .B1(new_n899), .B2(new_n612), .ZN(new_n900));
  INV_X1    g475(.A(new_n613), .ZN(new_n901));
  AOI22_X1  g476(.A1(new_n900), .A2(new_n901), .B1(new_n589), .B2(G54), .ZN(new_n902));
  INV_X1    g477(.A(KEYINPUT10), .ZN(new_n903));
  XNOR2_X1  g478(.A(new_n606), .B(new_n903), .ZN(new_n904));
  NAND3_X1  g479(.A1(G299), .A2(new_n902), .A3(new_n904), .ZN(new_n905));
  OAI21_X1  g480(.A(new_n620), .B1(new_n607), .B2(new_n615), .ZN(new_n906));
  NAND2_X1  g481(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n898), .A2(new_n907), .ZN(new_n908));
  AND3_X1   g483(.A1(new_n905), .A2(new_n906), .A3(KEYINPUT41), .ZN(new_n909));
  AOI21_X1  g484(.A(KEYINPUT41), .B1(new_n905), .B2(new_n906), .ZN(new_n910));
  NOR2_X1   g485(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  INV_X1    g486(.A(new_n911), .ZN(new_n912));
  NAND3_X1  g487(.A1(new_n896), .A2(new_n912), .A3(new_n897), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n908), .A2(new_n913), .ZN(new_n914));
  INV_X1    g489(.A(KEYINPUT42), .ZN(new_n915));
  NAND3_X1  g490(.A1(new_n914), .A2(KEYINPUT108), .A3(new_n915), .ZN(new_n916));
  NAND3_X1  g491(.A1(G166), .A2(new_n590), .A3(new_n582), .ZN(new_n917));
  INV_X1    g492(.A(new_n917), .ZN(new_n918));
  AOI21_X1  g493(.A(G166), .B1(new_n590), .B2(new_n582), .ZN(new_n919));
  OAI21_X1  g494(.A(KEYINPUT107), .B1(new_n918), .B2(new_n919), .ZN(new_n920));
  NAND2_X1  g495(.A1(G305), .A2(G303), .ZN(new_n921));
  INV_X1    g496(.A(KEYINPUT107), .ZN(new_n922));
  NAND3_X1  g497(.A1(new_n921), .A2(new_n922), .A3(new_n917), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n920), .A2(new_n923), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n708), .A2(new_n709), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n925), .A2(KEYINPUT106), .ZN(new_n926));
  INV_X1    g501(.A(KEYINPUT106), .ZN(new_n927));
  NAND3_X1  g502(.A1(new_n708), .A2(new_n927), .A3(new_n709), .ZN(new_n928));
  NAND3_X1  g503(.A1(new_n926), .A2(G290), .A3(new_n928), .ZN(new_n929));
  AND3_X1   g504(.A1(new_n708), .A2(new_n927), .A3(new_n709), .ZN(new_n930));
  AOI21_X1  g505(.A(new_n927), .B1(new_n708), .B2(new_n709), .ZN(new_n931));
  OAI21_X1  g506(.A(new_n603), .B1(new_n930), .B2(new_n931), .ZN(new_n932));
  AOI21_X1  g507(.A(new_n924), .B1(new_n929), .B2(new_n932), .ZN(new_n933));
  AOI21_X1  g508(.A(new_n922), .B1(new_n921), .B2(new_n917), .ZN(new_n934));
  AND3_X1   g509(.A1(new_n932), .A2(new_n929), .A3(new_n934), .ZN(new_n935));
  NOR2_X1   g510(.A1(new_n933), .A2(new_n935), .ZN(new_n936));
  INV_X1    g511(.A(KEYINPUT108), .ZN(new_n937));
  AOI21_X1  g512(.A(new_n936), .B1(new_n937), .B2(KEYINPUT42), .ZN(new_n938));
  OAI211_X1 g513(.A(new_n908), .B(new_n913), .C1(new_n937), .C2(KEYINPUT42), .ZN(new_n939));
  AND3_X1   g514(.A1(new_n916), .A2(new_n938), .A3(new_n939), .ZN(new_n940));
  AOI21_X1  g515(.A(new_n938), .B1(new_n916), .B2(new_n939), .ZN(new_n941));
  OAI21_X1  g516(.A(G868), .B1(new_n940), .B2(new_n941), .ZN(new_n942));
  INV_X1    g517(.A(KEYINPUT109), .ZN(new_n943));
  OR2_X1    g518(.A1(new_n845), .A2(G868), .ZN(new_n944));
  AND3_X1   g519(.A1(new_n942), .A2(new_n943), .A3(new_n944), .ZN(new_n945));
  AOI21_X1  g520(.A(new_n943), .B1(new_n942), .B2(new_n944), .ZN(new_n946));
  NOR2_X1   g521(.A1(new_n945), .A2(new_n946), .ZN(G295));
  NAND2_X1  g522(.A1(new_n942), .A2(new_n944), .ZN(G331));
  INV_X1    g523(.A(KEYINPUT44), .ZN(new_n949));
  INV_X1    g524(.A(KEYINPUT110), .ZN(new_n950));
  XNOR2_X1  g525(.A(G171), .B(G168), .ZN(new_n951));
  AOI21_X1  g526(.A(new_n845), .B1(new_n547), .B2(new_n554), .ZN(new_n952));
  OAI21_X1  g527(.A(new_n951), .B1(new_n952), .B2(new_n847), .ZN(new_n953));
  XNOR2_X1  g528(.A(G171), .B(G286), .ZN(new_n954));
  NAND3_X1  g529(.A1(new_n894), .A2(new_n846), .A3(new_n954), .ZN(new_n955));
  AOI211_X1 g530(.A(new_n950), .B(new_n911), .C1(new_n953), .C2(new_n955), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n953), .A2(new_n955), .ZN(new_n957));
  AOI21_X1  g532(.A(KEYINPUT110), .B1(new_n957), .B2(new_n912), .ZN(new_n958));
  NOR2_X1   g533(.A1(new_n956), .A2(new_n958), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n955), .A2(KEYINPUT111), .ZN(new_n960));
  INV_X1    g535(.A(KEYINPUT111), .ZN(new_n961));
  NAND3_X1  g536(.A1(new_n849), .A2(new_n961), .A3(new_n954), .ZN(new_n962));
  NAND4_X1  g537(.A1(new_n960), .A2(new_n962), .A3(new_n907), .A4(new_n953), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n936), .A2(new_n963), .ZN(new_n964));
  OAI21_X1  g539(.A(new_n884), .B1(new_n959), .B2(new_n964), .ZN(new_n965));
  NOR3_X1   g540(.A1(new_n952), .A2(new_n847), .A3(new_n951), .ZN(new_n966));
  AOI21_X1  g541(.A(new_n954), .B1(new_n894), .B2(new_n846), .ZN(new_n967));
  OAI21_X1  g542(.A(new_n912), .B1(new_n966), .B2(new_n967), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n968), .A2(new_n950), .ZN(new_n969));
  NAND3_X1  g544(.A1(new_n957), .A2(KEYINPUT110), .A3(new_n912), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n969), .A2(new_n970), .ZN(new_n971));
  AOI21_X1  g546(.A(new_n936), .B1(new_n971), .B2(new_n963), .ZN(new_n972));
  NOR2_X1   g547(.A1(new_n965), .A2(new_n972), .ZN(new_n973));
  INV_X1    g548(.A(KEYINPUT43), .ZN(new_n974));
  NOR2_X1   g549(.A1(new_n973), .A2(new_n974), .ZN(new_n975));
  NAND3_X1  g550(.A1(new_n932), .A2(new_n929), .A3(new_n934), .ZN(new_n976));
  AND2_X1   g551(.A1(new_n932), .A2(new_n929), .ZN(new_n977));
  OAI21_X1  g552(.A(new_n976), .B1(new_n977), .B2(new_n924), .ZN(new_n978));
  AND2_X1   g553(.A1(new_n960), .A2(new_n962), .ZN(new_n979));
  AND2_X1   g554(.A1(new_n953), .A2(new_n907), .ZN(new_n980));
  AOI21_X1  g555(.A(new_n978), .B1(new_n979), .B2(new_n980), .ZN(new_n981));
  AOI21_X1  g556(.A(G37), .B1(new_n981), .B2(new_n971), .ZN(new_n982));
  NAND3_X1  g557(.A1(new_n960), .A2(new_n962), .A3(new_n953), .ZN(new_n983));
  NAND2_X1  g558(.A1(new_n983), .A2(new_n912), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n980), .A2(new_n955), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n984), .A2(new_n985), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n986), .A2(new_n978), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n982), .A2(new_n987), .ZN(new_n988));
  NOR2_X1   g563(.A1(new_n988), .A2(KEYINPUT43), .ZN(new_n989));
  OAI21_X1  g564(.A(new_n949), .B1(new_n975), .B2(new_n989), .ZN(new_n990));
  AOI21_X1  g565(.A(new_n949), .B1(new_n973), .B2(new_n974), .ZN(new_n991));
  INV_X1    g566(.A(KEYINPUT112), .ZN(new_n992));
  AOI21_X1  g567(.A(new_n992), .B1(new_n988), .B2(KEYINPUT43), .ZN(new_n993));
  AOI211_X1 g568(.A(KEYINPUT112), .B(new_n974), .C1(new_n982), .C2(new_n987), .ZN(new_n994));
  OAI211_X1 g569(.A(new_n991), .B(KEYINPUT113), .C1(new_n993), .C2(new_n994), .ZN(new_n995));
  INV_X1    g570(.A(new_n995), .ZN(new_n996));
  AOI21_X1  g571(.A(new_n936), .B1(new_n984), .B2(new_n985), .ZN(new_n997));
  OAI21_X1  g572(.A(KEYINPUT43), .B1(new_n965), .B2(new_n997), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n998), .A2(KEYINPUT112), .ZN(new_n999));
  NAND3_X1  g574(.A1(new_n988), .A2(new_n992), .A3(KEYINPUT43), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n999), .A2(new_n1000), .ZN(new_n1001));
  AOI21_X1  g576(.A(KEYINPUT113), .B1(new_n1001), .B2(new_n991), .ZN(new_n1002));
  OAI21_X1  g577(.A(new_n990), .B1(new_n996), .B2(new_n1002), .ZN(G397));
  INV_X1    g578(.A(G1384), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n493), .A2(new_n1004), .ZN(new_n1005));
  XOR2_X1   g580(.A(KEYINPUT114), .B(KEYINPUT45), .Z(new_n1006));
  NAND2_X1  g581(.A1(new_n1005), .A2(new_n1006), .ZN(new_n1007));
  NAND2_X1  g582(.A1(G160), .A2(G40), .ZN(new_n1008));
  NOR2_X1   g583(.A1(new_n1007), .A2(new_n1008), .ZN(new_n1009));
  XNOR2_X1  g584(.A(new_n811), .B(G2067), .ZN(new_n1010));
  AND2_X1   g585(.A1(new_n1009), .A2(new_n1010), .ZN(new_n1011));
  INV_X1    g586(.A(new_n1009), .ZN(new_n1012));
  XOR2_X1   g587(.A(new_n791), .B(G1996), .Z(new_n1013));
  OAI22_X1  g588(.A1(new_n1011), .A2(KEYINPUT115), .B1(new_n1012), .B2(new_n1013), .ZN(new_n1014));
  AOI21_X1  g589(.A(new_n1014), .B1(KEYINPUT115), .B2(new_n1011), .ZN(new_n1015));
  XNOR2_X1  g590(.A(new_n740), .B(new_n742), .ZN(new_n1016));
  OAI21_X1  g591(.A(new_n1015), .B1(new_n1012), .B2(new_n1016), .ZN(new_n1017));
  INV_X1    g592(.A(G1986), .ZN(new_n1018));
  XNOR2_X1  g593(.A(new_n603), .B(new_n1018), .ZN(new_n1019));
  AOI21_X1  g594(.A(new_n1017), .B1(new_n1009), .B2(new_n1019), .ZN(new_n1020));
  XNOR2_X1  g595(.A(new_n1020), .B(KEYINPUT116), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n710), .A2(G1976), .ZN(new_n1022));
  INV_X1    g597(.A(G8), .ZN(new_n1023));
  INV_X1    g598(.A(G40), .ZN(new_n1024));
  NOR3_X1   g599(.A1(new_n471), .A2(new_n474), .A3(new_n1024), .ZN(new_n1025));
  AOI21_X1  g600(.A(G1384), .B1(new_n490), .B2(new_n492), .ZN(new_n1026));
  AOI21_X1  g601(.A(new_n1023), .B1(new_n1025), .B2(new_n1026), .ZN(new_n1027));
  INV_X1    g602(.A(G1976), .ZN(new_n1028));
  AOI21_X1  g603(.A(KEYINPUT52), .B1(G288), .B2(new_n1028), .ZN(new_n1029));
  NAND3_X1  g604(.A1(new_n1022), .A2(new_n1027), .A3(new_n1029), .ZN(new_n1030));
  NAND2_X1  g605(.A1(new_n1025), .A2(new_n1026), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n1031), .A2(G8), .ZN(new_n1032));
  AOI21_X1  g607(.A(new_n1032), .B1(G1976), .B2(new_n710), .ZN(new_n1033));
  INV_X1    g608(.A(KEYINPUT52), .ZN(new_n1034));
  OAI21_X1  g609(.A(new_n1030), .B1(new_n1033), .B2(new_n1034), .ZN(new_n1035));
  INV_X1    g610(.A(KEYINPUT118), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n588), .A2(G651), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n589), .A2(G48), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n1037), .A2(new_n1038), .ZN(new_n1039));
  INV_X1    g614(.A(new_n580), .ZN(new_n1040));
  OAI21_X1  g615(.A(G1981), .B1(new_n1039), .B2(new_n1040), .ZN(new_n1041));
  OAI21_X1  g616(.A(new_n1041), .B1(G1981), .B2(G305), .ZN(new_n1042));
  INV_X1    g617(.A(KEYINPUT49), .ZN(new_n1043));
  AOI21_X1  g618(.A(new_n1036), .B1(new_n1042), .B2(new_n1043), .ZN(new_n1044));
  INV_X1    g619(.A(new_n1044), .ZN(new_n1045));
  NAND3_X1  g620(.A1(new_n1042), .A2(new_n1036), .A3(new_n1043), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n1045), .A2(new_n1046), .ZN(new_n1047));
  NOR2_X1   g622(.A1(new_n1042), .A2(new_n1043), .ZN(new_n1048));
  NOR2_X1   g623(.A1(new_n1048), .A2(new_n1032), .ZN(new_n1049));
  AOI21_X1  g624(.A(new_n1035), .B1(new_n1047), .B2(new_n1049), .ZN(new_n1050));
  NAND2_X1  g625(.A1(G303), .A2(G8), .ZN(new_n1051));
  XNOR2_X1  g626(.A(new_n1051), .B(KEYINPUT55), .ZN(new_n1052));
  INV_X1    g627(.A(KEYINPUT50), .ZN(new_n1053));
  OAI21_X1  g628(.A(new_n1025), .B1(new_n1026), .B2(new_n1053), .ZN(new_n1054));
  INV_X1    g629(.A(new_n1054), .ZN(new_n1055));
  INV_X1    g630(.A(KEYINPUT117), .ZN(new_n1056));
  NAND3_X1  g631(.A1(new_n1026), .A2(new_n1056), .A3(new_n1053), .ZN(new_n1057));
  INV_X1    g632(.A(new_n1057), .ZN(new_n1058));
  AOI21_X1  g633(.A(new_n1056), .B1(new_n1026), .B2(new_n1053), .ZN(new_n1059));
  OAI211_X1 g634(.A(new_n1055), .B(new_n757), .C1(new_n1058), .C2(new_n1059), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n1026), .A2(KEYINPUT45), .ZN(new_n1061));
  NAND3_X1  g636(.A1(new_n1007), .A2(new_n1061), .A3(new_n1025), .ZN(new_n1062));
  INV_X1    g637(.A(G1971), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n1062), .A2(new_n1063), .ZN(new_n1064));
  AOI211_X1 g639(.A(new_n1023), .B(new_n1052), .C1(new_n1060), .C2(new_n1064), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n1050), .A2(new_n1065), .ZN(new_n1066));
  INV_X1    g641(.A(new_n1046), .ZN(new_n1067));
  OAI21_X1  g642(.A(new_n1049), .B1(new_n1067), .B2(new_n1044), .ZN(new_n1068));
  NOR2_X1   g643(.A1(G288), .A2(G1976), .ZN(new_n1069));
  AOI22_X1  g644(.A1(new_n1068), .A2(new_n1069), .B1(new_n696), .B2(new_n716), .ZN(new_n1070));
  OAI21_X1  g645(.A(new_n1066), .B1(new_n1032), .B2(new_n1070), .ZN(new_n1071));
  INV_X1    g646(.A(KEYINPUT45), .ZN(new_n1072));
  AOI21_X1  g647(.A(new_n1008), .B1(new_n1072), .B2(new_n1005), .ZN(new_n1073));
  OR2_X1    g648(.A1(new_n1005), .A2(new_n1006), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n1073), .A2(new_n1074), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n1075), .A2(new_n830), .ZN(new_n1076));
  OAI211_X1 g651(.A(new_n1055), .B(new_n766), .C1(new_n1058), .C2(new_n1059), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n1076), .A2(new_n1077), .ZN(new_n1078));
  OAI21_X1  g653(.A(G8), .B1(new_n1078), .B2(G286), .ZN(new_n1079));
  AOI21_X1  g654(.A(new_n1079), .B1(G286), .B2(new_n1078), .ZN(new_n1080));
  AOI21_X1  g655(.A(new_n1023), .B1(new_n1076), .B2(new_n1077), .ZN(new_n1081));
  OAI21_X1  g656(.A(KEYINPUT51), .B1(new_n1081), .B2(KEYINPUT125), .ZN(new_n1082));
  MUX2_X1   g657(.A(new_n1080), .B(new_n1079), .S(new_n1082), .Z(new_n1083));
  INV_X1    g658(.A(new_n1052), .ZN(new_n1084));
  INV_X1    g659(.A(KEYINPUT119), .ZN(new_n1085));
  NAND3_X1  g660(.A1(new_n1026), .A2(new_n1085), .A3(new_n1053), .ZN(new_n1086));
  INV_X1    g661(.A(new_n1086), .ZN(new_n1087));
  AOI21_X1  g662(.A(new_n1085), .B1(new_n1026), .B2(new_n1053), .ZN(new_n1088));
  OAI21_X1  g663(.A(new_n1055), .B1(new_n1087), .B2(new_n1088), .ZN(new_n1089));
  OAI21_X1  g664(.A(new_n1064), .B1(new_n1089), .B2(G2090), .ZN(new_n1090));
  AOI21_X1  g665(.A(new_n1084), .B1(new_n1090), .B2(G8), .ZN(new_n1091));
  NOR2_X1   g666(.A1(new_n1091), .A2(new_n1065), .ZN(new_n1092));
  OAI21_X1  g667(.A(new_n1055), .B1(new_n1058), .B2(new_n1059), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1093), .A2(new_n799), .ZN(new_n1094));
  INV_X1    g669(.A(KEYINPUT53), .ZN(new_n1095));
  OAI21_X1  g670(.A(new_n1095), .B1(new_n1062), .B2(G2078), .ZN(new_n1096));
  INV_X1    g671(.A(G2078), .ZN(new_n1097));
  NAND4_X1  g672(.A1(new_n1073), .A2(new_n1074), .A3(KEYINPUT53), .A4(new_n1097), .ZN(new_n1098));
  NAND3_X1  g673(.A1(new_n1094), .A2(new_n1096), .A3(new_n1098), .ZN(new_n1099));
  NAND4_X1  g674(.A1(new_n1092), .A2(G171), .A3(new_n1050), .A4(new_n1099), .ZN(new_n1100));
  INV_X1    g675(.A(KEYINPUT62), .ZN(new_n1101));
  NOR2_X1   g676(.A1(new_n1100), .A2(new_n1101), .ZN(new_n1102));
  AOI21_X1  g677(.A(new_n1071), .B1(new_n1083), .B2(new_n1102), .ZN(new_n1103));
  NOR2_X1   g678(.A1(new_n1100), .A2(KEYINPUT62), .ZN(new_n1104));
  INV_X1    g679(.A(KEYINPUT124), .ZN(new_n1105));
  OR2_X1    g680(.A1(new_n573), .A2(KEYINPUT123), .ZN(new_n1106));
  NAND2_X1  g681(.A1(new_n573), .A2(KEYINPUT123), .ZN(new_n1107));
  NAND3_X1  g682(.A1(new_n1106), .A2(new_n566), .A3(new_n1107), .ZN(new_n1108));
  XNOR2_X1  g683(.A(KEYINPUT122), .B(KEYINPUT57), .ZN(new_n1109));
  AOI22_X1  g684(.A1(new_n1108), .A2(new_n1109), .B1(KEYINPUT57), .B2(new_n620), .ZN(new_n1110));
  INV_X1    g685(.A(new_n1110), .ZN(new_n1111));
  AOI21_X1  g686(.A(new_n1008), .B1(new_n1005), .B2(new_n1006), .ZN(new_n1112));
  XNOR2_X1  g687(.A(KEYINPUT56), .B(G2072), .ZN(new_n1113));
  NAND3_X1  g688(.A1(new_n1112), .A2(new_n1061), .A3(new_n1113), .ZN(new_n1114));
  INV_X1    g689(.A(new_n1088), .ZN(new_n1115));
  AOI21_X1  g690(.A(new_n1054), .B1(new_n1115), .B2(new_n1086), .ZN(new_n1116));
  OAI211_X1 g691(.A(new_n1111), .B(new_n1114), .C1(new_n1116), .C2(G1956), .ZN(new_n1117));
  NOR2_X1   g692(.A1(new_n1031), .A2(G2067), .ZN(new_n1118));
  AOI21_X1  g693(.A(new_n1118), .B1(new_n1093), .B2(new_n834), .ZN(new_n1119));
  NOR2_X1   g694(.A1(new_n1119), .A2(new_n851), .ZN(new_n1120));
  INV_X1    g695(.A(G1956), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n1089), .A2(new_n1121), .ZN(new_n1122));
  AOI21_X1  g697(.A(new_n1111), .B1(new_n1122), .B2(new_n1114), .ZN(new_n1123));
  OAI211_X1 g698(.A(new_n1105), .B(new_n1117), .C1(new_n1120), .C2(new_n1123), .ZN(new_n1124));
  OAI21_X1  g699(.A(new_n1117), .B1(new_n1120), .B2(new_n1123), .ZN(new_n1125));
  NAND2_X1  g700(.A1(new_n1125), .A2(KEYINPUT124), .ZN(new_n1126));
  INV_X1    g701(.A(new_n1123), .ZN(new_n1127));
  NAND3_X1  g702(.A1(new_n1127), .A2(KEYINPUT61), .A3(new_n1117), .ZN(new_n1128));
  INV_X1    g703(.A(KEYINPUT61), .ZN(new_n1129));
  INV_X1    g704(.A(new_n1117), .ZN(new_n1130));
  OAI21_X1  g705(.A(new_n1129), .B1(new_n1130), .B2(new_n1123), .ZN(new_n1131));
  NAND2_X1  g706(.A1(new_n1128), .A2(new_n1131), .ZN(new_n1132));
  XOR2_X1   g707(.A(KEYINPUT58), .B(G1341), .Z(new_n1133));
  NAND2_X1  g708(.A1(new_n1031), .A2(new_n1133), .ZN(new_n1134));
  OAI21_X1  g709(.A(new_n1134), .B1(new_n1062), .B2(G1996), .ZN(new_n1135));
  AND3_X1   g710(.A1(new_n1135), .A2(KEYINPUT59), .A3(new_n556), .ZN(new_n1136));
  AOI21_X1  g711(.A(KEYINPUT59), .B1(new_n1135), .B2(new_n556), .ZN(new_n1137));
  NOR2_X1   g712(.A1(new_n1136), .A2(new_n1137), .ZN(new_n1138));
  NAND3_X1  g713(.A1(new_n1119), .A2(KEYINPUT60), .A3(new_n851), .ZN(new_n1139));
  NOR2_X1   g714(.A1(new_n1119), .A2(KEYINPUT60), .ZN(new_n1140));
  NAND2_X1  g715(.A1(new_n1093), .A2(new_n834), .ZN(new_n1141));
  NAND3_X1  g716(.A1(new_n1025), .A2(new_n1026), .A3(new_n814), .ZN(new_n1142));
  NAND3_X1  g717(.A1(new_n1141), .A2(KEYINPUT60), .A3(new_n1142), .ZN(new_n1143));
  NAND2_X1  g718(.A1(new_n1143), .A2(new_n616), .ZN(new_n1144));
  OAI211_X1 g719(.A(new_n1138), .B(new_n1139), .C1(new_n1140), .C2(new_n1144), .ZN(new_n1145));
  OAI211_X1 g720(.A(new_n1124), .B(new_n1126), .C1(new_n1132), .C2(new_n1145), .ZN(new_n1146));
  NAND4_X1  g721(.A1(new_n1112), .A2(KEYINPUT53), .A3(new_n1097), .A4(new_n1061), .ZN(new_n1147));
  NAND3_X1  g722(.A1(new_n1094), .A2(new_n1096), .A3(new_n1147), .ZN(new_n1148));
  NAND2_X1  g723(.A1(new_n1148), .A2(G171), .ZN(new_n1149));
  NAND2_X1  g724(.A1(new_n1149), .A2(KEYINPUT54), .ZN(new_n1150));
  NOR2_X1   g725(.A1(new_n1099), .A2(G171), .ZN(new_n1151));
  NOR2_X1   g726(.A1(new_n1150), .A2(new_n1151), .ZN(new_n1152));
  XOR2_X1   g727(.A(KEYINPUT126), .B(KEYINPUT54), .Z(new_n1153));
  NAND2_X1  g728(.A1(new_n1099), .A2(G171), .ZN(new_n1154));
  NAND4_X1  g729(.A1(new_n1094), .A2(G301), .A3(new_n1096), .A4(new_n1147), .ZN(new_n1155));
  AOI21_X1  g730(.A(new_n1153), .B1(new_n1154), .B2(new_n1155), .ZN(new_n1156));
  AOI22_X1  g731(.A1(new_n1116), .A2(new_n757), .B1(new_n1063), .B2(new_n1062), .ZN(new_n1157));
  OAI21_X1  g732(.A(new_n1052), .B1(new_n1157), .B2(new_n1023), .ZN(new_n1158));
  AOI21_X1  g733(.A(new_n1023), .B1(new_n1060), .B2(new_n1064), .ZN(new_n1159));
  NAND2_X1  g734(.A1(new_n1159), .A2(new_n1084), .ZN(new_n1160));
  NAND3_X1  g735(.A1(new_n1050), .A2(new_n1158), .A3(new_n1160), .ZN(new_n1161));
  NOR3_X1   g736(.A1(new_n1152), .A2(new_n1156), .A3(new_n1161), .ZN(new_n1162));
  AOI21_X1  g737(.A(new_n1104), .B1(new_n1146), .B2(new_n1162), .ZN(new_n1163));
  OAI21_X1  g738(.A(new_n1103), .B1(new_n1163), .B2(new_n1083), .ZN(new_n1164));
  AOI21_X1  g739(.A(new_n1034), .B1(new_n1022), .B2(new_n1027), .ZN(new_n1165));
  AOI21_X1  g740(.A(new_n1165), .B1(new_n1033), .B2(new_n1029), .ZN(new_n1166));
  AND3_X1   g741(.A1(new_n1068), .A2(new_n1166), .A3(G168), .ZN(new_n1167));
  NAND4_X1  g742(.A1(new_n1167), .A2(new_n1092), .A3(KEYINPUT120), .A4(new_n1081), .ZN(new_n1168));
  INV_X1    g743(.A(KEYINPUT120), .ZN(new_n1169));
  NAND2_X1  g744(.A1(new_n1158), .A2(new_n1160), .ZN(new_n1170));
  NAND4_X1  g745(.A1(new_n1068), .A2(new_n1081), .A3(new_n1166), .A4(G168), .ZN(new_n1171));
  OAI21_X1  g746(.A(new_n1169), .B1(new_n1170), .B2(new_n1171), .ZN(new_n1172));
  INV_X1    g747(.A(KEYINPUT63), .ZN(new_n1173));
  NAND3_X1  g748(.A1(new_n1168), .A2(new_n1172), .A3(new_n1173), .ZN(new_n1174));
  NAND2_X1  g749(.A1(new_n1174), .A2(KEYINPUT121), .ZN(new_n1175));
  INV_X1    g750(.A(KEYINPUT121), .ZN(new_n1176));
  NAND4_X1  g751(.A1(new_n1168), .A2(new_n1172), .A3(new_n1176), .A4(new_n1173), .ZN(new_n1177));
  NOR2_X1   g752(.A1(new_n1159), .A2(new_n1084), .ZN(new_n1178));
  OR4_X1    g753(.A1(new_n1173), .A2(new_n1171), .A3(new_n1065), .A4(new_n1178), .ZN(new_n1179));
  AND3_X1   g754(.A1(new_n1175), .A2(new_n1177), .A3(new_n1179), .ZN(new_n1180));
  OAI21_X1  g755(.A(new_n1021), .B1(new_n1164), .B2(new_n1180), .ZN(new_n1181));
  NAND3_X1  g756(.A1(new_n1009), .A2(new_n1018), .A3(new_n603), .ZN(new_n1182));
  XOR2_X1   g757(.A(new_n1182), .B(KEYINPUT48), .Z(new_n1183));
  NOR2_X1   g758(.A1(new_n1017), .A2(new_n1183), .ZN(new_n1184));
  NOR3_X1   g759(.A1(new_n736), .A2(new_n739), .A3(new_n742), .ZN(new_n1185));
  NAND2_X1  g760(.A1(new_n1015), .A2(new_n1185), .ZN(new_n1186));
  NAND2_X1  g761(.A1(new_n812), .A2(new_n814), .ZN(new_n1187));
  AOI21_X1  g762(.A(new_n1012), .B1(new_n1186), .B2(new_n1187), .ZN(new_n1188));
  OR3_X1    g763(.A1(new_n1012), .A2(KEYINPUT46), .A3(G1996), .ZN(new_n1189));
  OAI21_X1  g764(.A(KEYINPUT46), .B1(new_n1012), .B2(G1996), .ZN(new_n1190));
  OR2_X1    g765(.A1(new_n791), .A2(new_n1010), .ZN(new_n1191));
  AOI22_X1  g766(.A1(new_n1189), .A2(new_n1190), .B1(new_n1009), .B2(new_n1191), .ZN(new_n1192));
  XNOR2_X1  g767(.A(new_n1192), .B(KEYINPUT47), .ZN(new_n1193));
  NOR3_X1   g768(.A1(new_n1184), .A2(new_n1188), .A3(new_n1193), .ZN(new_n1194));
  NAND2_X1  g769(.A1(new_n1181), .A2(new_n1194), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g770(.A(G319), .ZN(new_n1197));
  NOR2_X1   g771(.A1(G227), .A2(new_n1197), .ZN(new_n1198));
  XNOR2_X1  g772(.A(new_n1198), .B(KEYINPUT127), .ZN(new_n1199));
  NOR2_X1   g773(.A1(new_n1199), .A2(G401), .ZN(new_n1200));
  NAND4_X1  g774(.A1(new_n889), .A2(new_n705), .A3(new_n703), .A4(new_n1200), .ZN(new_n1201));
  NOR2_X1   g775(.A1(new_n975), .A2(new_n989), .ZN(new_n1202));
  NOR2_X1   g776(.A1(new_n1201), .A2(new_n1202), .ZN(G308));
  OR2_X1    g777(.A1(new_n1201), .A2(new_n1202), .ZN(G225));
endmodule


