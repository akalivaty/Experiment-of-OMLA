//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 0 0 1 1 1 0 1 0 0 0 0 0 1 0 1 1 0 0 0 1 0 1 0 0 1 0 0 0 1 1 1 0 1 1 1 0 1 0 1 1 1 0 1 1 1 1 0 0 1 0 0 1 1 1 1 0 1 1 1 0 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:38:58 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n206, new_n207, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1198, new_n1199,
    new_n1200, new_n1201, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1219, new_n1220, new_n1221, new_n1222, new_n1223, new_n1224,
    new_n1225, new_n1226, new_n1227, new_n1228, new_n1229, new_n1230,
    new_n1231, new_n1232, new_n1233, new_n1234, new_n1235, new_n1237,
    new_n1238, new_n1239, new_n1240, new_n1241, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1300, new_n1301, new_n1302, new_n1303, new_n1304, new_n1305,
    new_n1306, new_n1307;
  INV_X1    g0000(.A(G50), .ZN(new_n201));
  INV_X1    g0001(.A(G58), .ZN(new_n202));
  INV_X1    g0002(.A(G68), .ZN(new_n203));
  NAND3_X1  g0003(.A1(new_n201), .A2(new_n202), .A3(new_n203), .ZN(new_n204));
  NOR2_X1   g0004(.A1(new_n204), .A2(G77), .ZN(G353));
  NOR2_X1   g0005(.A1(G97), .A2(G107), .ZN(new_n206));
  INV_X1    g0006(.A(new_n206), .ZN(new_n207));
  NAND2_X1  g0007(.A1(new_n207), .A2(G87), .ZN(G355));
  NAND2_X1  g0008(.A1(G1), .A2(G20), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n209), .A2(G13), .ZN(new_n210));
  OAI211_X1 g0010(.A(new_n210), .B(G250), .C1(G257), .C2(G264), .ZN(new_n211));
  XOR2_X1   g0011(.A(new_n211), .B(KEYINPUT0), .Z(new_n212));
  AOI22_X1  g0012(.A1(G77), .A2(G244), .B1(G97), .B2(G257), .ZN(new_n213));
  INV_X1    g0013(.A(G87), .ZN(new_n214));
  INV_X1    g0014(.A(G250), .ZN(new_n215));
  OAI21_X1  g0015(.A(new_n213), .B1(new_n214), .B2(new_n215), .ZN(new_n216));
  AOI21_X1  g0016(.A(new_n216), .B1(G116), .B2(G270), .ZN(new_n217));
  NAND2_X1  g0017(.A1(G58), .A2(G232), .ZN(new_n218));
  NAND2_X1  g0018(.A1(G107), .A2(G264), .ZN(new_n219));
  NAND2_X1  g0019(.A1(G50), .A2(G226), .ZN(new_n220));
  NAND4_X1  g0020(.A1(new_n217), .A2(new_n218), .A3(new_n219), .A4(new_n220), .ZN(new_n221));
  INV_X1    g0021(.A(G238), .ZN(new_n222));
  NOR2_X1   g0022(.A1(new_n203), .A2(new_n222), .ZN(new_n223));
  OAI21_X1  g0023(.A(new_n209), .B1(new_n221), .B2(new_n223), .ZN(new_n224));
  XNOR2_X1  g0024(.A(new_n224), .B(KEYINPUT1), .ZN(new_n225));
  NAND2_X1  g0025(.A1(G1), .A2(G13), .ZN(new_n226));
  INV_X1    g0026(.A(G20), .ZN(new_n227));
  NOR2_X1   g0027(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  OAI21_X1  g0028(.A(G50), .B1(G58), .B2(G68), .ZN(new_n229));
  XOR2_X1   g0029(.A(new_n229), .B(KEYINPUT64), .Z(new_n230));
  AOI211_X1 g0030(.A(new_n212), .B(new_n225), .C1(new_n228), .C2(new_n230), .ZN(G361));
  XOR2_X1   g0031(.A(KEYINPUT65), .B(KEYINPUT2), .Z(new_n232));
  XNOR2_X1  g0032(.A(G238), .B(G244), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n232), .B(new_n233), .ZN(new_n234));
  XNOR2_X1  g0034(.A(G226), .B(G232), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XOR2_X1   g0036(.A(G250), .B(G257), .Z(new_n237));
  XNOR2_X1  g0037(.A(G264), .B(G270), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XOR2_X1   g0039(.A(new_n236), .B(new_n239), .Z(G358));
  XNOR2_X1  g0040(.A(G50), .B(G58), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n241), .B(KEYINPUT66), .ZN(new_n242));
  XOR2_X1   g0042(.A(G68), .B(G77), .Z(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n244), .B(KEYINPUT67), .ZN(new_n245));
  XOR2_X1   g0045(.A(G87), .B(G97), .Z(new_n246));
  XNOR2_X1  g0046(.A(G107), .B(G116), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n246), .B(new_n247), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n245), .B(new_n248), .ZN(G351));
  INV_X1    g0049(.A(G1), .ZN(new_n250));
  NAND3_X1  g0050(.A1(new_n250), .A2(G13), .A3(G20), .ZN(new_n251));
  NOR2_X1   g0051(.A1(new_n251), .A2(G77), .ZN(new_n252));
  XNOR2_X1  g0052(.A(KEYINPUT8), .B(G58), .ZN(new_n253));
  INV_X1    g0053(.A(KEYINPUT70), .ZN(new_n254));
  XNOR2_X1  g0054(.A(new_n253), .B(new_n254), .ZN(new_n255));
  NOR2_X1   g0055(.A1(G20), .A2(G33), .ZN(new_n256));
  AOI22_X1  g0056(.A1(new_n255), .A2(new_n256), .B1(G20), .B2(G77), .ZN(new_n257));
  OR2_X1    g0057(.A1(new_n257), .A2(KEYINPUT71), .ZN(new_n258));
  XOR2_X1   g0058(.A(KEYINPUT15), .B(G87), .Z(new_n259));
  NAND3_X1  g0059(.A1(new_n259), .A2(new_n227), .A3(G33), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n257), .A2(KEYINPUT71), .ZN(new_n261));
  NAND3_X1  g0061(.A1(new_n258), .A2(new_n260), .A3(new_n261), .ZN(new_n262));
  NAND3_X1  g0062(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n263), .A2(new_n226), .ZN(new_n264));
  AOI21_X1  g0064(.A(new_n252), .B1(new_n262), .B2(new_n264), .ZN(new_n265));
  OAI211_X1 g0065(.A(new_n263), .B(new_n226), .C1(G1), .C2(new_n227), .ZN(new_n266));
  INV_X1    g0066(.A(new_n266), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n267), .A2(G77), .ZN(new_n268));
  XNOR2_X1  g0068(.A(new_n268), .B(KEYINPUT72), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n265), .A2(new_n269), .ZN(new_n270));
  AND2_X1   g0070(.A1(G33), .A2(G41), .ZN(new_n271));
  OAI21_X1  g0071(.A(KEYINPUT68), .B1(new_n271), .B2(new_n226), .ZN(new_n272));
  NAND2_X1  g0072(.A1(G33), .A2(G41), .ZN(new_n273));
  INV_X1    g0073(.A(KEYINPUT68), .ZN(new_n274));
  NAND4_X1  g0074(.A1(new_n273), .A2(new_n274), .A3(G1), .A4(G13), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n272), .A2(new_n275), .ZN(new_n276));
  INV_X1    g0076(.A(G41), .ZN(new_n277));
  INV_X1    g0077(.A(G45), .ZN(new_n278));
  AOI21_X1  g0078(.A(G1), .B1(new_n277), .B2(new_n278), .ZN(new_n279));
  INV_X1    g0079(.A(new_n279), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n276), .A2(new_n280), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n281), .A2(KEYINPUT69), .ZN(new_n282));
  AOI21_X1  g0082(.A(new_n279), .B1(new_n272), .B2(new_n275), .ZN(new_n283));
  INV_X1    g0083(.A(KEYINPUT69), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  NAND3_X1  g0085(.A1(new_n282), .A2(G244), .A3(new_n285), .ZN(new_n286));
  INV_X1    g0086(.A(G274), .ZN(new_n287));
  AOI21_X1  g0087(.A(new_n287), .B1(new_n272), .B2(new_n275), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n288), .A2(new_n279), .ZN(new_n289));
  OR2_X1    g0089(.A1(KEYINPUT3), .A2(G33), .ZN(new_n290));
  NAND2_X1  g0090(.A1(KEYINPUT3), .A2(G33), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  INV_X1    g0092(.A(G1698), .ZN(new_n293));
  NAND3_X1  g0093(.A1(new_n292), .A2(G232), .A3(new_n293), .ZN(new_n294));
  NAND3_X1  g0094(.A1(new_n292), .A2(G238), .A3(G1698), .ZN(new_n295));
  INV_X1    g0095(.A(G107), .ZN(new_n296));
  OAI211_X1 g0096(.A(new_n294), .B(new_n295), .C1(new_n296), .C2(new_n292), .ZN(new_n297));
  NOR2_X1   g0097(.A1(new_n271), .A2(new_n226), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n297), .A2(new_n298), .ZN(new_n299));
  NAND3_X1  g0099(.A1(new_n286), .A2(new_n289), .A3(new_n299), .ZN(new_n300));
  INV_X1    g0100(.A(G169), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  OR2_X1    g0102(.A1(new_n300), .A2(G179), .ZN(new_n303));
  NAND3_X1  g0103(.A1(new_n270), .A2(new_n302), .A3(new_n303), .ZN(new_n304));
  INV_X1    g0104(.A(G190), .ZN(new_n305));
  OR2_X1    g0105(.A1(new_n300), .A2(new_n305), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n300), .A2(G200), .ZN(new_n307));
  NAND4_X1  g0107(.A1(new_n265), .A2(new_n306), .A3(new_n269), .A4(new_n307), .ZN(new_n308));
  AND2_X1   g0108(.A1(new_n304), .A2(new_n308), .ZN(new_n309));
  INV_X1    g0109(.A(KEYINPUT74), .ZN(new_n310));
  INV_X1    g0110(.A(new_n289), .ZN(new_n311));
  OAI21_X1  g0111(.A(new_n292), .B1(G232), .B2(new_n293), .ZN(new_n312));
  NOR2_X1   g0112(.A1(G226), .A2(G1698), .ZN(new_n313));
  INV_X1    g0113(.A(G33), .ZN(new_n314));
  INV_X1    g0114(.A(G97), .ZN(new_n315));
  OAI22_X1  g0115(.A1(new_n312), .A2(new_n313), .B1(new_n314), .B2(new_n315), .ZN(new_n316));
  AOI21_X1  g0116(.A(new_n311), .B1(new_n298), .B2(new_n316), .ZN(new_n317));
  NAND3_X1  g0117(.A1(new_n282), .A2(G238), .A3(new_n285), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n317), .A2(new_n318), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n319), .A2(KEYINPUT13), .ZN(new_n320));
  INV_X1    g0120(.A(KEYINPUT13), .ZN(new_n321));
  NAND3_X1  g0121(.A1(new_n317), .A2(new_n321), .A3(new_n318), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n320), .A2(new_n322), .ZN(new_n323));
  AOI21_X1  g0123(.A(new_n310), .B1(new_n323), .B2(G200), .ZN(new_n324));
  INV_X1    g0124(.A(G200), .ZN(new_n325));
  AOI211_X1 g0125(.A(KEYINPUT74), .B(new_n325), .C1(new_n320), .C2(new_n322), .ZN(new_n326));
  NOR2_X1   g0126(.A1(new_n324), .A2(new_n326), .ZN(new_n327));
  INV_X1    g0127(.A(new_n256), .ZN(new_n328));
  OAI22_X1  g0128(.A1(new_n328), .A2(new_n201), .B1(new_n227), .B2(G68), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n227), .A2(G33), .ZN(new_n330));
  INV_X1    g0130(.A(G77), .ZN(new_n331));
  NOR2_X1   g0131(.A1(new_n330), .A2(new_n331), .ZN(new_n332));
  OAI21_X1  g0132(.A(new_n264), .B1(new_n329), .B2(new_n332), .ZN(new_n333));
  XOR2_X1   g0133(.A(new_n333), .B(KEYINPUT11), .Z(new_n334));
  NOR2_X1   g0134(.A1(new_n266), .A2(new_n203), .ZN(new_n335));
  INV_X1    g0135(.A(new_n251), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n336), .A2(new_n203), .ZN(new_n337));
  INV_X1    g0137(.A(KEYINPUT12), .ZN(new_n338));
  XNOR2_X1  g0138(.A(new_n337), .B(new_n338), .ZN(new_n339));
  NOR3_X1   g0139(.A1(new_n334), .A2(new_n335), .A3(new_n339), .ZN(new_n340));
  OAI21_X1  g0140(.A(new_n340), .B1(new_n323), .B2(new_n305), .ZN(new_n341));
  INV_X1    g0141(.A(new_n341), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n327), .A2(new_n342), .ZN(new_n343));
  INV_X1    g0143(.A(new_n322), .ZN(new_n344));
  AOI21_X1  g0144(.A(new_n321), .B1(new_n317), .B2(new_n318), .ZN(new_n345));
  OAI21_X1  g0145(.A(G169), .B1(new_n344), .B2(new_n345), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n346), .A2(KEYINPUT14), .ZN(new_n347));
  INV_X1    g0147(.A(KEYINPUT14), .ZN(new_n348));
  NAND3_X1  g0148(.A1(new_n323), .A2(new_n348), .A3(G169), .ZN(new_n349));
  NOR2_X1   g0149(.A1(new_n344), .A2(new_n345), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n350), .A2(G179), .ZN(new_n351));
  NAND3_X1  g0151(.A1(new_n347), .A2(new_n349), .A3(new_n351), .ZN(new_n352));
  INV_X1    g0152(.A(new_n340), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n352), .A2(new_n353), .ZN(new_n354));
  NAND3_X1  g0154(.A1(new_n309), .A2(new_n343), .A3(new_n354), .ZN(new_n355));
  NOR2_X1   g0155(.A1(new_n251), .A2(G50), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n204), .A2(G20), .ZN(new_n357));
  INV_X1    g0157(.A(G150), .ZN(new_n358));
  OAI221_X1 g0158(.A(new_n357), .B1(new_n358), .B2(new_n328), .C1(new_n330), .C2(new_n253), .ZN(new_n359));
  AOI21_X1  g0159(.A(new_n356), .B1(new_n359), .B2(new_n264), .ZN(new_n360));
  NOR2_X1   g0160(.A1(new_n266), .A2(new_n201), .ZN(new_n361));
  INV_X1    g0161(.A(new_n361), .ZN(new_n362));
  AND2_X1   g0162(.A1(new_n360), .A2(new_n362), .ZN(new_n363));
  INV_X1    g0163(.A(KEYINPUT73), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n363), .A2(new_n364), .ZN(new_n365));
  AOI21_X1  g0165(.A(new_n364), .B1(new_n360), .B2(new_n362), .ZN(new_n366));
  INV_X1    g0166(.A(new_n366), .ZN(new_n367));
  NAND3_X1  g0167(.A1(new_n365), .A2(new_n367), .A3(KEYINPUT9), .ZN(new_n368));
  INV_X1    g0168(.A(KEYINPUT9), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n360), .A2(new_n362), .ZN(new_n370));
  NOR2_X1   g0170(.A1(new_n370), .A2(KEYINPUT73), .ZN(new_n371));
  OAI21_X1  g0171(.A(new_n369), .B1(new_n371), .B2(new_n366), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n368), .A2(new_n372), .ZN(new_n373));
  AND2_X1   g0173(.A1(KEYINPUT3), .A2(G33), .ZN(new_n374));
  NOR2_X1   g0174(.A1(KEYINPUT3), .A2(G33), .ZN(new_n375));
  NOR2_X1   g0175(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n376), .A2(new_n331), .ZN(new_n377));
  INV_X1    g0177(.A(new_n298), .ZN(new_n378));
  OR2_X1    g0178(.A1(G222), .A2(G1698), .ZN(new_n379));
  OAI21_X1  g0179(.A(new_n379), .B1(G223), .B2(new_n293), .ZN(new_n380));
  AOI21_X1  g0180(.A(new_n378), .B1(new_n292), .B2(new_n380), .ZN(new_n381));
  AOI21_X1  g0181(.A(new_n311), .B1(new_n377), .B2(new_n381), .ZN(new_n382));
  NAND3_X1  g0182(.A1(new_n282), .A2(G226), .A3(new_n285), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n382), .A2(new_n383), .ZN(new_n384));
  INV_X1    g0184(.A(new_n384), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n385), .A2(G190), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n384), .A2(G200), .ZN(new_n387));
  NAND3_X1  g0187(.A1(new_n373), .A2(new_n386), .A3(new_n387), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n388), .A2(KEYINPUT10), .ZN(new_n389));
  INV_X1    g0189(.A(KEYINPUT10), .ZN(new_n390));
  NAND4_X1  g0190(.A1(new_n373), .A2(new_n390), .A3(new_n386), .A4(new_n387), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n389), .A2(new_n391), .ZN(new_n392));
  NOR2_X1   g0192(.A1(new_n384), .A2(G179), .ZN(new_n393));
  AOI211_X1 g0193(.A(new_n363), .B(new_n393), .C1(new_n301), .C2(new_n384), .ZN(new_n394));
  INV_X1    g0194(.A(new_n394), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n253), .A2(new_n251), .ZN(new_n396));
  OAI21_X1  g0196(.A(new_n396), .B1(new_n267), .B2(new_n253), .ZN(new_n397));
  XNOR2_X1  g0197(.A(new_n397), .B(KEYINPUT76), .ZN(new_n398));
  AOI21_X1  g0198(.A(KEYINPUT7), .B1(new_n376), .B2(new_n227), .ZN(new_n399));
  INV_X1    g0199(.A(KEYINPUT7), .ZN(new_n400));
  NOR4_X1   g0200(.A1(new_n374), .A2(new_n375), .A3(new_n400), .A4(G20), .ZN(new_n401));
  OAI21_X1  g0201(.A(G68), .B1(new_n399), .B2(new_n401), .ZN(new_n402));
  INV_X1    g0202(.A(KEYINPUT16), .ZN(new_n403));
  NOR2_X1   g0203(.A1(new_n202), .A2(new_n203), .ZN(new_n404));
  NOR2_X1   g0204(.A1(G58), .A2(G68), .ZN(new_n405));
  OAI21_X1  g0205(.A(G20), .B1(new_n404), .B2(new_n405), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n256), .A2(G159), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  INV_X1    g0208(.A(new_n408), .ZN(new_n409));
  NAND4_X1  g0209(.A1(new_n402), .A2(KEYINPUT75), .A3(new_n403), .A4(new_n409), .ZN(new_n410));
  AND2_X1   g0210(.A1(new_n410), .A2(new_n264), .ZN(new_n411));
  NAND3_X1  g0211(.A1(new_n290), .A2(new_n227), .A3(new_n291), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n412), .A2(new_n400), .ZN(new_n413));
  NAND4_X1  g0213(.A1(new_n290), .A2(KEYINPUT7), .A3(new_n227), .A4(new_n291), .ZN(new_n414));
  AOI21_X1  g0214(.A(new_n203), .B1(new_n413), .B2(new_n414), .ZN(new_n415));
  OAI21_X1  g0215(.A(KEYINPUT16), .B1(new_n415), .B2(new_n408), .ZN(new_n416));
  NAND3_X1  g0216(.A1(new_n402), .A2(new_n403), .A3(new_n409), .ZN(new_n417));
  NAND3_X1  g0217(.A1(new_n409), .A2(KEYINPUT75), .A3(new_n403), .ZN(new_n418));
  NAND3_X1  g0218(.A1(new_n416), .A2(new_n417), .A3(new_n418), .ZN(new_n419));
  AOI21_X1  g0219(.A(new_n398), .B1(new_n411), .B2(new_n419), .ZN(new_n420));
  OR2_X1    g0220(.A1(G223), .A2(G1698), .ZN(new_n421));
  OAI221_X1 g0221(.A(new_n421), .B1(G226), .B2(new_n293), .C1(new_n374), .C2(new_n375), .ZN(new_n422));
  OAI21_X1  g0222(.A(new_n422), .B1(new_n314), .B2(new_n214), .ZN(new_n423));
  AOI22_X1  g0223(.A1(new_n423), .A2(new_n298), .B1(G232), .B2(new_n283), .ZN(new_n424));
  NAND3_X1  g0224(.A1(new_n424), .A2(new_n305), .A3(new_n289), .ZN(new_n425));
  OR2_X1    g0225(.A1(new_n425), .A2(KEYINPUT78), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n423), .A2(new_n298), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n283), .A2(G232), .ZN(new_n428));
  NAND3_X1  g0228(.A1(new_n427), .A2(new_n289), .A3(new_n428), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n429), .A2(new_n325), .ZN(new_n430));
  NAND3_X1  g0230(.A1(new_n430), .A2(KEYINPUT78), .A3(new_n425), .ZN(new_n431));
  NAND3_X1  g0231(.A1(new_n420), .A2(new_n426), .A3(new_n431), .ZN(new_n432));
  INV_X1    g0232(.A(KEYINPUT17), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n432), .A2(new_n433), .ZN(new_n434));
  NAND4_X1  g0234(.A1(new_n420), .A2(KEYINPUT17), .A3(new_n426), .A4(new_n431), .ZN(new_n435));
  AND2_X1   g0235(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  NAND3_X1  g0236(.A1(new_n419), .A2(new_n264), .A3(new_n410), .ZN(new_n437));
  INV_X1    g0237(.A(new_n398), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n437), .A2(new_n438), .ZN(new_n439));
  INV_X1    g0239(.A(G179), .ZN(new_n440));
  NOR2_X1   g0240(.A1(new_n429), .A2(new_n440), .ZN(new_n441));
  AOI21_X1  g0241(.A(new_n301), .B1(new_n424), .B2(new_n289), .ZN(new_n442));
  OAI21_X1  g0242(.A(KEYINPUT77), .B1(new_n441), .B2(new_n442), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n429), .A2(G169), .ZN(new_n444));
  INV_X1    g0244(.A(KEYINPUT77), .ZN(new_n445));
  OAI211_X1 g0245(.A(new_n444), .B(new_n445), .C1(new_n440), .C2(new_n429), .ZN(new_n446));
  NAND3_X1  g0246(.A1(new_n439), .A2(new_n443), .A3(new_n446), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n447), .A2(KEYINPUT18), .ZN(new_n448));
  INV_X1    g0248(.A(KEYINPUT18), .ZN(new_n449));
  NAND4_X1  g0249(.A1(new_n439), .A2(new_n449), .A3(new_n443), .A4(new_n446), .ZN(new_n450));
  AND2_X1   g0250(.A1(new_n448), .A2(new_n450), .ZN(new_n451));
  NAND4_X1  g0251(.A1(new_n392), .A2(new_n395), .A3(new_n436), .A4(new_n451), .ZN(new_n452));
  NOR2_X1   g0252(.A1(new_n355), .A2(new_n452), .ZN(new_n453));
  INV_X1    g0253(.A(new_n453), .ZN(new_n454));
  INV_X1    g0254(.A(G116), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n336), .A2(new_n455), .ZN(new_n456));
  AND2_X1   g0256(.A1(new_n263), .A2(new_n226), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n250), .A2(G33), .ZN(new_n458));
  NAND4_X1  g0258(.A1(new_n457), .A2(G116), .A3(new_n458), .A4(new_n251), .ZN(new_n459));
  AOI22_X1  g0259(.A1(new_n263), .A2(new_n226), .B1(G20), .B2(new_n455), .ZN(new_n460));
  NAND2_X1  g0260(.A1(G33), .A2(G283), .ZN(new_n461));
  OAI211_X1 g0261(.A(new_n461), .B(new_n227), .C1(G33), .C2(new_n315), .ZN(new_n462));
  AND3_X1   g0262(.A1(new_n460), .A2(KEYINPUT20), .A3(new_n462), .ZN(new_n463));
  AOI21_X1  g0263(.A(KEYINPUT20), .B1(new_n460), .B2(new_n462), .ZN(new_n464));
  OAI211_X1 g0264(.A(new_n456), .B(new_n459), .C1(new_n463), .C2(new_n464), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n465), .A2(G179), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n277), .A2(KEYINPUT5), .ZN(new_n467));
  INV_X1    g0267(.A(KEYINPUT5), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n468), .A2(G41), .ZN(new_n469));
  NAND4_X1  g0269(.A1(new_n469), .A2(KEYINPUT83), .A3(new_n250), .A4(G45), .ZN(new_n470));
  OAI211_X1 g0270(.A(new_n250), .B(G45), .C1(new_n277), .C2(KEYINPUT5), .ZN(new_n471));
  INV_X1    g0271(.A(KEYINPUT83), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  NAND4_X1  g0273(.A1(new_n288), .A2(new_n467), .A3(new_n470), .A4(new_n473), .ZN(new_n474));
  NAND3_X1  g0274(.A1(new_n473), .A2(new_n467), .A3(new_n470), .ZN(new_n475));
  NAND3_X1  g0275(.A1(new_n475), .A2(G270), .A3(new_n276), .ZN(new_n476));
  OAI211_X1 g0276(.A(G257), .B(new_n293), .C1(new_n374), .C2(new_n375), .ZN(new_n477));
  OAI211_X1 g0277(.A(G264), .B(G1698), .C1(new_n374), .C2(new_n375), .ZN(new_n478));
  NAND3_X1  g0278(.A1(new_n290), .A2(G303), .A3(new_n291), .ZN(new_n479));
  NAND3_X1  g0279(.A1(new_n477), .A2(new_n478), .A3(new_n479), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n480), .A2(new_n298), .ZN(new_n481));
  NAND3_X1  g0281(.A1(new_n474), .A2(new_n476), .A3(new_n481), .ZN(new_n482));
  NOR2_X1   g0282(.A1(new_n466), .A2(new_n482), .ZN(new_n483));
  NAND3_X1  g0283(.A1(new_n482), .A2(G169), .A3(new_n465), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n484), .A2(KEYINPUT21), .ZN(new_n485));
  INV_X1    g0285(.A(KEYINPUT21), .ZN(new_n486));
  NAND4_X1  g0286(.A1(new_n482), .A2(new_n486), .A3(G169), .A4(new_n465), .ZN(new_n487));
  AOI21_X1  g0287(.A(new_n483), .B1(new_n485), .B2(new_n487), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n482), .A2(G200), .ZN(new_n489));
  OAI21_X1  g0289(.A(new_n489), .B1(new_n305), .B2(new_n482), .ZN(new_n490));
  OAI21_X1  g0290(.A(new_n488), .B1(new_n465), .B2(new_n490), .ZN(new_n491));
  OAI21_X1  g0291(.A(G107), .B1(new_n399), .B2(new_n401), .ZN(new_n492));
  INV_X1    g0292(.A(KEYINPUT6), .ZN(new_n493));
  NOR2_X1   g0293(.A1(new_n315), .A2(new_n296), .ZN(new_n494));
  OAI21_X1  g0294(.A(new_n493), .B1(new_n494), .B2(new_n206), .ZN(new_n495));
  NAND3_X1  g0295(.A1(new_n296), .A2(KEYINPUT6), .A3(G97), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n497), .A2(G20), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n256), .A2(G77), .ZN(new_n499));
  XOR2_X1   g0299(.A(new_n499), .B(KEYINPUT79), .Z(new_n500));
  NAND3_X1  g0300(.A1(new_n492), .A2(new_n498), .A3(new_n500), .ZN(new_n501));
  AND3_X1   g0301(.A1(new_n501), .A2(KEYINPUT80), .A3(new_n264), .ZN(new_n502));
  AOI21_X1  g0302(.A(KEYINPUT80), .B1(new_n501), .B2(new_n264), .ZN(new_n503));
  NOR2_X1   g0303(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  NOR2_X1   g0304(.A1(new_n336), .A2(G97), .ZN(new_n505));
  NAND3_X1  g0305(.A1(new_n457), .A2(new_n458), .A3(new_n251), .ZN(new_n506));
  AOI21_X1  g0306(.A(new_n505), .B1(new_n506), .B2(G97), .ZN(new_n507));
  INV_X1    g0307(.A(KEYINPUT81), .ZN(new_n508));
  XNOR2_X1  g0308(.A(new_n507), .B(new_n508), .ZN(new_n509));
  OAI211_X1 g0309(.A(G244), .B(new_n293), .C1(new_n374), .C2(new_n375), .ZN(new_n510));
  INV_X1    g0310(.A(KEYINPUT4), .ZN(new_n511));
  AOI22_X1  g0311(.A1(new_n510), .A2(new_n511), .B1(G33), .B2(G283), .ZN(new_n512));
  NAND4_X1  g0312(.A1(new_n292), .A2(KEYINPUT4), .A3(G244), .A4(new_n293), .ZN(new_n513));
  OAI211_X1 g0313(.A(G250), .B(G1698), .C1(new_n374), .C2(new_n375), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n514), .A2(KEYINPUT82), .ZN(new_n515));
  INV_X1    g0315(.A(KEYINPUT82), .ZN(new_n516));
  NAND4_X1  g0316(.A1(new_n292), .A2(new_n516), .A3(G250), .A4(G1698), .ZN(new_n517));
  NAND4_X1  g0317(.A1(new_n512), .A2(new_n513), .A3(new_n515), .A4(new_n517), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n518), .A2(new_n298), .ZN(new_n519));
  NAND3_X1  g0319(.A1(new_n475), .A2(G257), .A3(new_n276), .ZN(new_n520));
  NAND3_X1  g0320(.A1(new_n519), .A2(new_n520), .A3(new_n474), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n521), .A2(G200), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n276), .A2(G274), .ZN(new_n523));
  NOR2_X1   g0323(.A1(new_n523), .A2(new_n475), .ZN(new_n524));
  AOI21_X1  g0324(.A(new_n524), .B1(new_n518), .B2(new_n298), .ZN(new_n525));
  NAND3_X1  g0325(.A1(new_n525), .A2(G190), .A3(new_n520), .ZN(new_n526));
  NAND4_X1  g0326(.A1(new_n504), .A2(new_n509), .A3(new_n522), .A4(new_n526), .ZN(new_n527));
  NAND3_X1  g0327(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n528), .A2(new_n227), .ZN(new_n529));
  OAI21_X1  g0329(.A(new_n529), .B1(new_n207), .B2(G87), .ZN(new_n530));
  OAI211_X1 g0330(.A(new_n227), .B(G68), .C1(new_n374), .C2(new_n375), .ZN(new_n531));
  INV_X1    g0331(.A(KEYINPUT19), .ZN(new_n532));
  OAI21_X1  g0332(.A(new_n532), .B1(new_n330), .B2(new_n315), .ZN(new_n533));
  NAND3_X1  g0333(.A1(new_n530), .A2(new_n531), .A3(new_n533), .ZN(new_n534));
  INV_X1    g0334(.A(new_n259), .ZN(new_n535));
  AOI22_X1  g0335(.A1(new_n534), .A2(new_n264), .B1(new_n535), .B2(new_n336), .ZN(new_n536));
  INV_X1    g0336(.A(new_n506), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n537), .A2(new_n259), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n536), .A2(new_n538), .ZN(new_n539));
  AOI21_X1  g0339(.A(G250), .B1(new_n250), .B2(G45), .ZN(new_n540));
  AOI21_X1  g0340(.A(new_n540), .B1(new_n272), .B2(new_n275), .ZN(new_n541));
  NOR3_X1   g0341(.A1(new_n278), .A2(G1), .A3(G274), .ZN(new_n542));
  INV_X1    g0342(.A(new_n542), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n541), .A2(new_n543), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n222), .A2(new_n293), .ZN(new_n545));
  INV_X1    g0345(.A(G244), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n546), .A2(G1698), .ZN(new_n547));
  OAI211_X1 g0347(.A(new_n545), .B(new_n547), .C1(new_n374), .C2(new_n375), .ZN(new_n548));
  NAND2_X1  g0348(.A1(G33), .A2(G116), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n550), .A2(new_n298), .ZN(new_n551));
  NAND3_X1  g0351(.A1(new_n544), .A2(new_n551), .A3(new_n440), .ZN(new_n552));
  AOI211_X1 g0352(.A(new_n540), .B(new_n542), .C1(new_n272), .C2(new_n275), .ZN(new_n553));
  AOI21_X1  g0353(.A(new_n378), .B1(new_n548), .B2(new_n549), .ZN(new_n554));
  OAI21_X1  g0354(.A(new_n301), .B1(new_n553), .B2(new_n554), .ZN(new_n555));
  NAND3_X1  g0355(.A1(new_n539), .A2(new_n552), .A3(new_n555), .ZN(new_n556));
  OAI21_X1  g0356(.A(G200), .B1(new_n553), .B2(new_n554), .ZN(new_n557));
  NAND3_X1  g0357(.A1(new_n544), .A2(new_n551), .A3(G190), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n537), .A2(G87), .ZN(new_n559));
  NAND4_X1  g0359(.A1(new_n557), .A2(new_n558), .A3(new_n536), .A4(new_n559), .ZN(new_n560));
  AND2_X1   g0360(.A1(new_n556), .A2(new_n560), .ZN(new_n561));
  INV_X1    g0361(.A(KEYINPUT80), .ZN(new_n562));
  AOI21_X1  g0362(.A(new_n296), .B1(new_n413), .B2(new_n414), .ZN(new_n563));
  AOI21_X1  g0363(.A(new_n227), .B1(new_n495), .B2(new_n496), .ZN(new_n564));
  XNOR2_X1  g0364(.A(new_n499), .B(KEYINPUT79), .ZN(new_n565));
  NOR3_X1   g0365(.A1(new_n563), .A2(new_n564), .A3(new_n565), .ZN(new_n566));
  OAI21_X1  g0366(.A(new_n562), .B1(new_n566), .B2(new_n457), .ZN(new_n567));
  NAND3_X1  g0367(.A1(new_n501), .A2(KEYINPUT80), .A3(new_n264), .ZN(new_n568));
  NAND3_X1  g0368(.A1(new_n567), .A2(new_n509), .A3(new_n568), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n521), .A2(new_n301), .ZN(new_n570));
  NAND3_X1  g0370(.A1(new_n525), .A2(new_n440), .A3(new_n520), .ZN(new_n571));
  NAND3_X1  g0371(.A1(new_n569), .A2(new_n570), .A3(new_n571), .ZN(new_n572));
  NAND3_X1  g0372(.A1(new_n527), .A2(new_n561), .A3(new_n572), .ZN(new_n573));
  INV_X1    g0373(.A(KEYINPUT84), .ZN(new_n574));
  AOI21_X1  g0374(.A(new_n491), .B1(new_n573), .B2(new_n574), .ZN(new_n575));
  NAND4_X1  g0375(.A1(new_n527), .A2(new_n572), .A3(KEYINPUT84), .A4(new_n561), .ZN(new_n576));
  INV_X1    g0376(.A(KEYINPUT24), .ZN(new_n577));
  OAI211_X1 g0377(.A(new_n227), .B(G87), .C1(new_n374), .C2(new_n375), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n578), .A2(KEYINPUT22), .ZN(new_n579));
  INV_X1    g0379(.A(KEYINPUT22), .ZN(new_n580));
  NAND4_X1  g0380(.A1(new_n292), .A2(new_n580), .A3(new_n227), .A4(G87), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n579), .A2(new_n581), .ZN(new_n582));
  INV_X1    g0382(.A(KEYINPUT85), .ZN(new_n583));
  NOR2_X1   g0383(.A1(new_n330), .A2(new_n455), .ZN(new_n584));
  INV_X1    g0384(.A(KEYINPUT23), .ZN(new_n585));
  OAI21_X1  g0385(.A(new_n585), .B1(new_n227), .B2(G107), .ZN(new_n586));
  NAND3_X1  g0386(.A1(new_n296), .A2(KEYINPUT23), .A3(G20), .ZN(new_n587));
  AOI21_X1  g0387(.A(new_n584), .B1(new_n586), .B2(new_n587), .ZN(new_n588));
  AND3_X1   g0388(.A1(new_n582), .A2(new_n583), .A3(new_n588), .ZN(new_n589));
  AOI21_X1  g0389(.A(new_n583), .B1(new_n582), .B2(new_n588), .ZN(new_n590));
  OAI21_X1  g0390(.A(new_n577), .B1(new_n589), .B2(new_n590), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n582), .A2(new_n588), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n592), .A2(KEYINPUT85), .ZN(new_n593));
  NAND3_X1  g0393(.A1(new_n582), .A2(new_n583), .A3(new_n588), .ZN(new_n594));
  NAND3_X1  g0394(.A1(new_n593), .A2(KEYINPUT24), .A3(new_n594), .ZN(new_n595));
  NAND3_X1  g0395(.A1(new_n591), .A2(new_n595), .A3(new_n264), .ZN(new_n596));
  INV_X1    g0396(.A(KEYINPUT25), .ZN(new_n597));
  OAI21_X1  g0397(.A(new_n597), .B1(new_n251), .B2(G107), .ZN(new_n598));
  NAND3_X1  g0398(.A1(new_n336), .A2(KEYINPUT25), .A3(new_n296), .ZN(new_n599));
  AOI22_X1  g0399(.A1(new_n537), .A2(G107), .B1(new_n598), .B2(new_n599), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n596), .A2(new_n600), .ZN(new_n601));
  NAND3_X1  g0401(.A1(new_n475), .A2(G264), .A3(new_n276), .ZN(new_n602));
  OAI211_X1 g0402(.A(G257), .B(G1698), .C1(new_n374), .C2(new_n375), .ZN(new_n603));
  OAI211_X1 g0403(.A(G250), .B(new_n293), .C1(new_n374), .C2(new_n375), .ZN(new_n604));
  NAND2_X1  g0404(.A1(G33), .A2(G294), .ZN(new_n605));
  NAND3_X1  g0405(.A1(new_n603), .A2(new_n604), .A3(new_n605), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n606), .A2(new_n298), .ZN(new_n607));
  NAND3_X1  g0407(.A1(new_n474), .A2(new_n602), .A3(new_n607), .ZN(new_n608));
  AND2_X1   g0408(.A1(new_n608), .A2(G169), .ZN(new_n609));
  NOR2_X1   g0409(.A1(new_n608), .A2(new_n440), .ZN(new_n610));
  OAI21_X1  g0410(.A(KEYINPUT86), .B1(new_n609), .B2(new_n610), .ZN(new_n611));
  AND3_X1   g0411(.A1(new_n474), .A2(new_n602), .A3(new_n607), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n612), .A2(G179), .ZN(new_n613));
  INV_X1    g0413(.A(KEYINPUT86), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n608), .A2(G169), .ZN(new_n615));
  NAND3_X1  g0415(.A1(new_n613), .A2(new_n614), .A3(new_n615), .ZN(new_n616));
  NAND3_X1  g0416(.A1(new_n601), .A2(new_n611), .A3(new_n616), .ZN(new_n617));
  INV_X1    g0417(.A(KEYINPUT88), .ZN(new_n618));
  NAND3_X1  g0418(.A1(new_n612), .A2(KEYINPUT87), .A3(new_n305), .ZN(new_n619));
  INV_X1    g0419(.A(KEYINPUT87), .ZN(new_n620));
  AOI21_X1  g0420(.A(new_n620), .B1(new_n608), .B2(new_n325), .ZN(new_n621));
  NOR2_X1   g0421(.A1(new_n608), .A2(G190), .ZN(new_n622));
  OAI21_X1  g0422(.A(new_n619), .B1(new_n621), .B2(new_n622), .ZN(new_n623));
  NAND3_X1  g0423(.A1(new_n623), .A2(new_n596), .A3(new_n600), .ZN(new_n624));
  AND3_X1   g0424(.A1(new_n617), .A2(new_n618), .A3(new_n624), .ZN(new_n625));
  AOI21_X1  g0425(.A(new_n618), .B1(new_n617), .B2(new_n624), .ZN(new_n626));
  OAI211_X1 g0426(.A(new_n575), .B(new_n576), .C1(new_n625), .C2(new_n626), .ZN(new_n627));
  NOR2_X1   g0427(.A1(new_n454), .A2(new_n627), .ZN(G372));
  INV_X1    g0428(.A(new_n392), .ZN(new_n629));
  OAI21_X1  g0429(.A(new_n444), .B1(new_n440), .B2(new_n429), .ZN(new_n630));
  AND3_X1   g0430(.A1(new_n439), .A2(KEYINPUT18), .A3(new_n630), .ZN(new_n631));
  AOI21_X1  g0431(.A(KEYINPUT18), .B1(new_n439), .B2(new_n630), .ZN(new_n632));
  NOR2_X1   g0432(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  NOR3_X1   g0433(.A1(new_n341), .A2(new_n324), .A3(new_n326), .ZN(new_n634));
  AOI21_X1  g0434(.A(new_n634), .B1(new_n354), .B2(new_n304), .ZN(new_n635));
  AOI21_X1  g0435(.A(new_n633), .B1(new_n635), .B2(new_n436), .ZN(new_n636));
  AOI21_X1  g0436(.A(new_n629), .B1(new_n636), .B2(KEYINPUT90), .ZN(new_n637));
  INV_X1    g0437(.A(KEYINPUT90), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n354), .A2(new_n304), .ZN(new_n639));
  AND3_X1   g0439(.A1(new_n639), .A2(new_n343), .A3(new_n436), .ZN(new_n640));
  OAI21_X1  g0440(.A(new_n638), .B1(new_n640), .B2(new_n633), .ZN(new_n641));
  AOI21_X1  g0441(.A(new_n394), .B1(new_n637), .B2(new_n641), .ZN(new_n642));
  AND2_X1   g0442(.A1(new_n569), .A2(new_n570), .ZN(new_n643));
  NAND4_X1  g0443(.A1(new_n643), .A2(KEYINPUT26), .A3(new_n561), .A4(new_n571), .ZN(new_n644));
  NAND4_X1  g0444(.A1(new_n561), .A2(new_n569), .A3(new_n570), .A4(new_n571), .ZN(new_n645));
  INV_X1    g0445(.A(KEYINPUT26), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n644), .A2(new_n647), .ZN(new_n648));
  NOR2_X1   g0448(.A1(new_n488), .A2(KEYINPUT89), .ZN(new_n649));
  INV_X1    g0449(.A(KEYINPUT89), .ZN(new_n650));
  AOI211_X1 g0450(.A(new_n650), .B(new_n483), .C1(new_n485), .C2(new_n487), .ZN(new_n651));
  AOI22_X1  g0451(.A1(new_n596), .A2(new_n600), .B1(new_n615), .B2(new_n613), .ZN(new_n652));
  NOR3_X1   g0452(.A1(new_n649), .A2(new_n651), .A3(new_n652), .ZN(new_n653));
  NAND4_X1  g0453(.A1(new_n624), .A2(new_n527), .A3(new_n560), .A4(new_n572), .ZN(new_n654));
  OAI211_X1 g0454(.A(new_n648), .B(new_n556), .C1(new_n653), .C2(new_n654), .ZN(new_n655));
  INV_X1    g0455(.A(new_n655), .ZN(new_n656));
  OAI21_X1  g0456(.A(new_n642), .B1(new_n454), .B2(new_n656), .ZN(G369));
  INV_X1    g0457(.A(G13), .ZN(new_n658));
  NOR2_X1   g0458(.A1(new_n658), .A2(G20), .ZN(new_n659));
  INV_X1    g0459(.A(new_n659), .ZN(new_n660));
  OR3_X1    g0460(.A1(new_n660), .A2(KEYINPUT27), .A3(G1), .ZN(new_n661));
  OAI21_X1  g0461(.A(KEYINPUT27), .B1(new_n660), .B2(G1), .ZN(new_n662));
  NAND3_X1  g0462(.A1(new_n661), .A2(G213), .A3(new_n662), .ZN(new_n663));
  INV_X1    g0463(.A(G343), .ZN(new_n664));
  NOR2_X1   g0464(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n601), .A2(new_n665), .ZN(new_n666));
  XNOR2_X1  g0466(.A(new_n666), .B(KEYINPUT91), .ZN(new_n667));
  NAND3_X1  g0467(.A1(new_n617), .A2(new_n618), .A3(new_n624), .ZN(new_n668));
  AND2_X1   g0468(.A1(new_n596), .A2(new_n600), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n611), .A2(new_n616), .ZN(new_n670));
  OAI21_X1  g0470(.A(new_n624), .B1(new_n669), .B2(new_n670), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n671), .A2(KEYINPUT88), .ZN(new_n672));
  AOI21_X1  g0472(.A(new_n667), .B1(new_n668), .B2(new_n672), .ZN(new_n673));
  INV_X1    g0473(.A(new_n665), .ZN(new_n674));
  NOR2_X1   g0474(.A1(new_n617), .A2(new_n674), .ZN(new_n675));
  NOR2_X1   g0475(.A1(new_n673), .A2(new_n675), .ZN(new_n676));
  AND2_X1   g0476(.A1(new_n665), .A2(new_n465), .ZN(new_n677));
  OR2_X1    g0477(.A1(new_n491), .A2(new_n677), .ZN(new_n678));
  OAI21_X1  g0478(.A(new_n677), .B1(new_n649), .B2(new_n651), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n680), .A2(G330), .ZN(new_n681));
  NOR2_X1   g0481(.A1(new_n676), .A2(new_n681), .ZN(new_n682));
  NOR2_X1   g0482(.A1(new_n488), .A2(new_n665), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n673), .A2(new_n683), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n652), .A2(new_n674), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  NOR2_X1   g0486(.A1(new_n682), .A2(new_n686), .ZN(new_n687));
  XNOR2_X1  g0487(.A(new_n687), .B(KEYINPUT92), .ZN(G399));
  INV_X1    g0488(.A(new_n210), .ZN(new_n689));
  NOR2_X1   g0489(.A1(new_n689), .A2(G41), .ZN(new_n690));
  INV_X1    g0490(.A(new_n690), .ZN(new_n691));
  NOR3_X1   g0491(.A1(new_n207), .A2(G87), .A3(G116), .ZN(new_n692));
  NAND3_X1  g0492(.A1(new_n691), .A2(G1), .A3(new_n692), .ZN(new_n693));
  INV_X1    g0493(.A(new_n230), .ZN(new_n694));
  OAI21_X1  g0494(.A(new_n693), .B1(new_n694), .B2(new_n691), .ZN(new_n695));
  XOR2_X1   g0495(.A(KEYINPUT93), .B(KEYINPUT28), .Z(new_n696));
  XNOR2_X1  g0496(.A(new_n695), .B(new_n696), .ZN(new_n697));
  NOR2_X1   g0497(.A1(new_n553), .A2(new_n554), .ZN(new_n698));
  AND2_X1   g0498(.A1(new_n476), .A2(new_n481), .ZN(new_n699));
  NAND4_X1  g0499(.A1(new_n612), .A2(G179), .A3(new_n698), .A4(new_n699), .ZN(new_n700));
  OAI21_X1  g0500(.A(KEYINPUT94), .B1(new_n700), .B2(new_n521), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n701), .A2(KEYINPUT30), .ZN(new_n702));
  INV_X1    g0502(.A(KEYINPUT30), .ZN(new_n703));
  OAI211_X1 g0503(.A(KEYINPUT94), .B(new_n703), .C1(new_n700), .C2(new_n521), .ZN(new_n704));
  AOI22_X1  g0504(.A1(new_n525), .A2(new_n520), .B1(new_n699), .B2(new_n474), .ZN(new_n705));
  INV_X1    g0505(.A(new_n698), .ZN(new_n706));
  NAND4_X1  g0506(.A1(new_n705), .A2(new_n440), .A3(new_n706), .A4(new_n608), .ZN(new_n707));
  NAND3_X1  g0507(.A1(new_n702), .A2(new_n704), .A3(new_n707), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n708), .A2(new_n665), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n709), .A2(KEYINPUT31), .ZN(new_n710));
  INV_X1    g0510(.A(KEYINPUT31), .ZN(new_n711));
  NAND3_X1  g0511(.A1(new_n708), .A2(new_n711), .A3(new_n665), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n710), .A2(new_n712), .ZN(new_n713));
  OAI21_X1  g0513(.A(new_n713), .B1(new_n627), .B2(new_n665), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n714), .A2(G330), .ZN(new_n715));
  OR3_X1    g0515(.A1(new_n645), .A2(KEYINPUT95), .A3(new_n646), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n617), .A2(new_n488), .ZN(new_n717));
  INV_X1    g0517(.A(new_n717), .ZN(new_n718));
  OAI21_X1  g0518(.A(new_n716), .B1(new_n718), .B2(new_n654), .ZN(new_n719));
  NAND3_X1  g0519(.A1(new_n644), .A2(new_n647), .A3(KEYINPUT95), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n720), .A2(new_n556), .ZN(new_n721));
  OAI21_X1  g0521(.A(new_n674), .B1(new_n719), .B2(new_n721), .ZN(new_n722));
  NAND2_X1  g0522(.A1(new_n722), .A2(KEYINPUT29), .ZN(new_n723));
  INV_X1    g0523(.A(new_n654), .ZN(new_n724));
  AND2_X1   g0524(.A1(new_n485), .A2(new_n487), .ZN(new_n725));
  OAI21_X1  g0525(.A(new_n650), .B1(new_n725), .B2(new_n483), .ZN(new_n726));
  INV_X1    g0526(.A(new_n652), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n488), .A2(KEYINPUT89), .ZN(new_n728));
  NAND3_X1  g0528(.A1(new_n726), .A2(new_n727), .A3(new_n728), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n724), .A2(new_n729), .ZN(new_n730));
  INV_X1    g0530(.A(new_n556), .ZN(new_n731));
  AOI21_X1  g0531(.A(new_n731), .B1(new_n644), .B2(new_n647), .ZN(new_n732));
  AOI21_X1  g0532(.A(new_n665), .B1(new_n730), .B2(new_n732), .ZN(new_n733));
  INV_X1    g0533(.A(KEYINPUT29), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  NAND3_X1  g0535(.A1(new_n715), .A2(new_n723), .A3(new_n735), .ZN(new_n736));
  INV_X1    g0536(.A(new_n736), .ZN(new_n737));
  OAI21_X1  g0537(.A(new_n697), .B1(new_n737), .B2(G1), .ZN(G364));
  INV_X1    g0538(.A(new_n680), .ZN(new_n739));
  INV_X1    g0539(.A(G330), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  AOI21_X1  g0541(.A(new_n250), .B1(new_n659), .B2(G45), .ZN(new_n742));
  INV_X1    g0542(.A(new_n742), .ZN(new_n743));
  NOR2_X1   g0543(.A1(new_n690), .A2(new_n743), .ZN(new_n744));
  INV_X1    g0544(.A(new_n744), .ZN(new_n745));
  NAND3_X1  g0545(.A1(new_n741), .A2(new_n681), .A3(new_n745), .ZN(new_n746));
  XNOR2_X1  g0546(.A(new_n746), .B(KEYINPUT96), .ZN(new_n747));
  NOR2_X1   g0547(.A1(G13), .A2(G33), .ZN(new_n748));
  INV_X1    g0548(.A(new_n748), .ZN(new_n749));
  NOR2_X1   g0549(.A1(new_n749), .A2(G20), .ZN(new_n750));
  AOI21_X1  g0550(.A(new_n745), .B1(new_n739), .B2(new_n750), .ZN(new_n751));
  NOR2_X1   g0551(.A1(new_n227), .A2(new_n305), .ZN(new_n752));
  NOR2_X1   g0552(.A1(new_n440), .A2(G200), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  INV_X1    g0554(.A(new_n754), .ZN(new_n755));
  NOR2_X1   g0555(.A1(new_n227), .A2(G190), .ZN(new_n756));
  NOR2_X1   g0556(.A1(G179), .A2(G200), .ZN(new_n757));
  NAND2_X1  g0557(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  INV_X1    g0558(.A(new_n758), .ZN(new_n759));
  AOI22_X1  g0559(.A1(G322), .A2(new_n755), .B1(new_n759), .B2(G329), .ZN(new_n760));
  NAND2_X1  g0560(.A1(new_n760), .A2(new_n376), .ZN(new_n761));
  NOR2_X1   g0561(.A1(new_n440), .A2(new_n325), .ZN(new_n762));
  NAND2_X1  g0562(.A1(new_n752), .A2(new_n762), .ZN(new_n763));
  INV_X1    g0563(.A(new_n763), .ZN(new_n764));
  AOI21_X1  g0564(.A(new_n761), .B1(G326), .B2(new_n764), .ZN(new_n765));
  NOR2_X1   g0565(.A1(new_n325), .A2(G179), .ZN(new_n766));
  NAND2_X1  g0566(.A1(new_n752), .A2(new_n766), .ZN(new_n767));
  INV_X1    g0567(.A(new_n767), .ZN(new_n768));
  NAND2_X1  g0568(.A1(new_n768), .A2(G303), .ZN(new_n769));
  NAND2_X1  g0569(.A1(new_n757), .A2(G190), .ZN(new_n770));
  NAND2_X1  g0570(.A1(new_n770), .A2(G20), .ZN(new_n771));
  NAND2_X1  g0571(.A1(new_n771), .A2(G294), .ZN(new_n772));
  XOR2_X1   g0572(.A(KEYINPUT33), .B(G317), .Z(new_n773));
  NAND2_X1  g0573(.A1(new_n762), .A2(new_n756), .ZN(new_n774));
  NAND2_X1  g0574(.A1(new_n756), .A2(new_n753), .ZN(new_n775));
  INV_X1    g0575(.A(G311), .ZN(new_n776));
  OAI22_X1  g0576(.A1(new_n773), .A2(new_n774), .B1(new_n775), .B2(new_n776), .ZN(new_n777));
  NAND2_X1  g0577(.A1(new_n756), .A2(new_n766), .ZN(new_n778));
  INV_X1    g0578(.A(new_n778), .ZN(new_n779));
  AOI21_X1  g0579(.A(new_n777), .B1(G283), .B2(new_n779), .ZN(new_n780));
  NAND4_X1  g0580(.A1(new_n765), .A2(new_n769), .A3(new_n772), .A4(new_n780), .ZN(new_n781));
  INV_X1    g0581(.A(new_n771), .ZN(new_n782));
  NOR2_X1   g0582(.A1(new_n782), .A2(new_n315), .ZN(new_n783));
  INV_X1    g0583(.A(new_n774), .ZN(new_n784));
  AOI21_X1  g0584(.A(new_n783), .B1(G68), .B2(new_n784), .ZN(new_n785));
  XNOR2_X1  g0585(.A(new_n785), .B(KEYINPUT98), .ZN(new_n786));
  OAI22_X1  g0586(.A1(new_n754), .A2(new_n202), .B1(new_n778), .B2(new_n296), .ZN(new_n787));
  AOI21_X1  g0587(.A(new_n787), .B1(G87), .B2(new_n768), .ZN(new_n788));
  INV_X1    g0588(.A(new_n775), .ZN(new_n789));
  AOI21_X1  g0589(.A(new_n376), .B1(new_n789), .B2(G77), .ZN(new_n790));
  NAND2_X1  g0590(.A1(new_n759), .A2(G159), .ZN(new_n791));
  AOI22_X1  g0591(.A1(new_n791), .A2(KEYINPUT32), .B1(G50), .B2(new_n764), .ZN(new_n792));
  NAND4_X1  g0592(.A1(new_n786), .A2(new_n788), .A3(new_n790), .A4(new_n792), .ZN(new_n793));
  NOR2_X1   g0593(.A1(new_n791), .A2(KEYINPUT32), .ZN(new_n794));
  OAI21_X1  g0594(.A(new_n781), .B1(new_n793), .B2(new_n794), .ZN(new_n795));
  AOI21_X1  g0595(.A(new_n226), .B1(G20), .B2(new_n301), .ZN(new_n796));
  NAND2_X1  g0596(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  NAND2_X1  g0597(.A1(new_n244), .A2(G45), .ZN(new_n798));
  XOR2_X1   g0598(.A(new_n798), .B(KEYINPUT97), .Z(new_n799));
  NOR2_X1   g0599(.A1(new_n689), .A2(new_n292), .ZN(new_n800));
  OAI211_X1 g0600(.A(new_n799), .B(new_n800), .C1(G45), .C2(new_n694), .ZN(new_n801));
  INV_X1    g0601(.A(G355), .ZN(new_n802));
  NAND2_X1  g0602(.A1(new_n292), .A2(new_n210), .ZN(new_n803));
  OAI221_X1 g0603(.A(new_n801), .B1(G116), .B2(new_n210), .C1(new_n802), .C2(new_n803), .ZN(new_n804));
  NOR2_X1   g0604(.A1(new_n750), .A2(new_n796), .ZN(new_n805));
  NAND2_X1  g0605(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  NAND3_X1  g0606(.A1(new_n751), .A2(new_n797), .A3(new_n806), .ZN(new_n807));
  NAND2_X1  g0607(.A1(new_n747), .A2(new_n807), .ZN(G396));
  NOR2_X1   g0608(.A1(new_n304), .A2(new_n665), .ZN(new_n809));
  INV_X1    g0609(.A(new_n809), .ZN(new_n810));
  NAND2_X1  g0610(.A1(new_n270), .A2(new_n665), .ZN(new_n811));
  NAND2_X1  g0611(.A1(new_n811), .A2(new_n308), .ZN(new_n812));
  NAND2_X1  g0612(.A1(new_n812), .A2(new_n304), .ZN(new_n813));
  NAND2_X1  g0613(.A1(new_n810), .A2(new_n813), .ZN(new_n814));
  INV_X1    g0614(.A(KEYINPUT100), .ZN(new_n815));
  OAI211_X1 g0615(.A(new_n814), .B(new_n815), .C1(new_n656), .C2(new_n665), .ZN(new_n816));
  AOI21_X1  g0616(.A(new_n809), .B1(new_n304), .B2(new_n812), .ZN(new_n817));
  OAI21_X1  g0617(.A(KEYINPUT100), .B1(new_n817), .B2(new_n733), .ZN(new_n818));
  NAND2_X1  g0618(.A1(new_n816), .A2(new_n818), .ZN(new_n819));
  INV_X1    g0619(.A(new_n715), .ZN(new_n820));
  NAND3_X1  g0620(.A1(new_n655), .A2(new_n309), .A3(new_n674), .ZN(new_n821));
  INV_X1    g0621(.A(KEYINPUT101), .ZN(new_n822));
  NAND2_X1  g0622(.A1(new_n821), .A2(new_n822), .ZN(new_n823));
  NAND3_X1  g0623(.A1(new_n733), .A2(KEYINPUT101), .A3(new_n309), .ZN(new_n824));
  NAND2_X1  g0624(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  NAND3_X1  g0625(.A1(new_n819), .A2(new_n820), .A3(new_n825), .ZN(new_n826));
  NAND2_X1  g0626(.A1(new_n826), .A2(new_n745), .ZN(new_n827));
  NAND2_X1  g0627(.A1(new_n827), .A2(KEYINPUT102), .ZN(new_n828));
  INV_X1    g0628(.A(KEYINPUT102), .ZN(new_n829));
  NAND3_X1  g0629(.A1(new_n826), .A2(new_n829), .A3(new_n745), .ZN(new_n830));
  AND2_X1   g0630(.A1(new_n819), .A2(new_n825), .ZN(new_n831));
  OAI211_X1 g0631(.A(new_n828), .B(new_n830), .C1(new_n820), .C2(new_n831), .ZN(new_n832));
  INV_X1    g0632(.A(new_n796), .ZN(new_n833));
  INV_X1    g0633(.A(G132), .ZN(new_n834));
  NOR2_X1   g0634(.A1(new_n758), .A2(new_n834), .ZN(new_n835));
  XNOR2_X1  g0635(.A(KEYINPUT99), .B(G143), .ZN(new_n836));
  AOI22_X1  g0636(.A1(new_n755), .A2(new_n836), .B1(new_n789), .B2(G159), .ZN(new_n837));
  INV_X1    g0637(.A(G137), .ZN(new_n838));
  OAI221_X1 g0638(.A(new_n837), .B1(new_n838), .B2(new_n763), .C1(new_n358), .C2(new_n774), .ZN(new_n839));
  XOR2_X1   g0639(.A(new_n839), .B(KEYINPUT34), .Z(new_n840));
  AOI211_X1 g0640(.A(new_n835), .B(new_n840), .C1(G58), .C2(new_n771), .ZN(new_n841));
  NOR2_X1   g0641(.A1(new_n778), .A2(new_n203), .ZN(new_n842));
  INV_X1    g0642(.A(new_n842), .ZN(new_n843));
  NAND2_X1  g0643(.A1(new_n768), .A2(G50), .ZN(new_n844));
  NAND4_X1  g0644(.A1(new_n841), .A2(new_n292), .A3(new_n843), .A4(new_n844), .ZN(new_n845));
  NOR2_X1   g0645(.A1(new_n767), .A2(new_n296), .ZN(new_n846));
  AOI211_X1 g0646(.A(new_n846), .B(new_n783), .C1(G116), .C2(new_n789), .ZN(new_n847));
  NAND2_X1  g0647(.A1(new_n755), .A2(G294), .ZN(new_n848));
  NOR2_X1   g0648(.A1(new_n778), .A2(new_n214), .ZN(new_n849));
  INV_X1    g0649(.A(G283), .ZN(new_n850));
  OAI21_X1  g0650(.A(new_n376), .B1(new_n774), .B2(new_n850), .ZN(new_n851));
  AOI211_X1 g0651(.A(new_n849), .B(new_n851), .C1(G303), .C2(new_n764), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n759), .A2(G311), .ZN(new_n853));
  NAND4_X1  g0653(.A1(new_n847), .A2(new_n848), .A3(new_n852), .A4(new_n853), .ZN(new_n854));
  AOI21_X1  g0654(.A(new_n833), .B1(new_n845), .B2(new_n854), .ZN(new_n855));
  AOI211_X1 g0655(.A(new_n745), .B(new_n855), .C1(new_n748), .C2(new_n814), .ZN(new_n856));
  NOR2_X1   g0656(.A1(new_n796), .A2(new_n748), .ZN(new_n857));
  INV_X1    g0657(.A(new_n857), .ZN(new_n858));
  OAI21_X1  g0658(.A(new_n856), .B1(G77), .B2(new_n858), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n832), .A2(new_n859), .ZN(G384));
  INV_X1    g0660(.A(KEYINPUT40), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n714), .A2(KEYINPUT108), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n672), .A2(new_n668), .ZN(new_n863));
  NAND4_X1  g0663(.A1(new_n863), .A2(new_n575), .A3(new_n576), .A4(new_n674), .ZN(new_n864));
  INV_X1    g0664(.A(KEYINPUT108), .ZN(new_n865));
  NAND3_X1  g0665(.A1(new_n864), .A2(new_n865), .A3(new_n713), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n862), .A2(new_n866), .ZN(new_n867));
  NAND4_X1  g0667(.A1(new_n448), .A2(new_n434), .A3(new_n435), .A4(new_n450), .ZN(new_n868));
  INV_X1    g0668(.A(new_n663), .ZN(new_n869));
  AND2_X1   g0669(.A1(new_n416), .A2(new_n417), .ZN(new_n870));
  OAI21_X1  g0670(.A(new_n438), .B1(new_n870), .B2(new_n457), .ZN(new_n871));
  NAND3_X1  g0671(.A1(new_n868), .A2(new_n869), .A3(new_n871), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n439), .A2(new_n869), .ZN(new_n873));
  INV_X1    g0673(.A(KEYINPUT37), .ZN(new_n874));
  NAND4_X1  g0674(.A1(new_n447), .A2(new_n873), .A3(new_n874), .A4(new_n432), .ZN(new_n875));
  OAI21_X1  g0675(.A(new_n871), .B1(new_n630), .B2(new_n869), .ZN(new_n876));
  AND2_X1   g0676(.A1(new_n432), .A2(new_n876), .ZN(new_n877));
  OAI21_X1  g0677(.A(new_n875), .B1(new_n877), .B2(new_n874), .ZN(new_n878));
  AND3_X1   g0678(.A1(new_n872), .A2(KEYINPUT38), .A3(new_n878), .ZN(new_n879));
  AOI21_X1  g0679(.A(KEYINPUT38), .B1(new_n872), .B2(new_n878), .ZN(new_n880));
  OR2_X1    g0680(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n353), .A2(new_n665), .ZN(new_n882));
  NAND3_X1  g0682(.A1(new_n343), .A2(new_n354), .A3(new_n882), .ZN(new_n883));
  NAND3_X1  g0683(.A1(new_n352), .A2(new_n353), .A3(new_n665), .ZN(new_n884));
  AND2_X1   g0684(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  INV_X1    g0685(.A(new_n885), .ZN(new_n886));
  NAND4_X1  g0686(.A1(new_n867), .A2(new_n881), .A3(new_n817), .A4(new_n886), .ZN(new_n887));
  AOI211_X1 g0687(.A(new_n814), .B(new_n885), .C1(new_n862), .C2(new_n866), .ZN(new_n888));
  INV_X1    g0688(.A(KEYINPUT105), .ZN(new_n889));
  INV_X1    g0689(.A(new_n873), .ZN(new_n890));
  OAI211_X1 g0690(.A(new_n434), .B(new_n435), .C1(new_n631), .C2(new_n632), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n439), .A2(new_n630), .ZN(new_n892));
  NAND3_X1  g0692(.A1(new_n892), .A2(new_n873), .A3(new_n432), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n893), .A2(KEYINPUT37), .ZN(new_n894));
  AOI22_X1  g0694(.A1(new_n890), .A2(new_n891), .B1(new_n894), .B2(new_n875), .ZN(new_n895));
  OAI21_X1  g0695(.A(new_n889), .B1(new_n895), .B2(KEYINPUT38), .ZN(new_n896));
  INV_X1    g0696(.A(KEYINPUT38), .ZN(new_n897));
  AND2_X1   g0697(.A1(new_n891), .A2(new_n890), .ZN(new_n898));
  AND3_X1   g0698(.A1(new_n873), .A2(new_n432), .A3(new_n874), .ZN(new_n899));
  AOI22_X1  g0699(.A1(new_n899), .A2(new_n447), .B1(new_n893), .B2(KEYINPUT37), .ZN(new_n900));
  OAI211_X1 g0700(.A(KEYINPUT105), .B(new_n897), .C1(new_n898), .C2(new_n900), .ZN(new_n901));
  NAND3_X1  g0701(.A1(new_n872), .A2(KEYINPUT38), .A3(new_n878), .ZN(new_n902));
  NAND3_X1  g0702(.A1(new_n896), .A2(new_n901), .A3(new_n902), .ZN(new_n903));
  AND2_X1   g0703(.A1(new_n903), .A2(KEYINPUT40), .ZN(new_n904));
  AOI22_X1  g0704(.A1(new_n861), .A2(new_n887), .B1(new_n888), .B2(new_n904), .ZN(new_n905));
  NAND3_X1  g0705(.A1(new_n905), .A2(new_n453), .A3(new_n867), .ZN(new_n906));
  AND3_X1   g0706(.A1(new_n864), .A2(new_n865), .A3(new_n713), .ZN(new_n907));
  AOI21_X1  g0707(.A(new_n865), .B1(new_n864), .B2(new_n713), .ZN(new_n908));
  OAI211_X1 g0708(.A(new_n886), .B(new_n817), .C1(new_n907), .C2(new_n908), .ZN(new_n909));
  NOR2_X1   g0709(.A1(new_n879), .A2(new_n880), .ZN(new_n910));
  OAI21_X1  g0710(.A(new_n861), .B1(new_n909), .B2(new_n910), .ZN(new_n911));
  AOI21_X1  g0711(.A(new_n814), .B1(new_n862), .B2(new_n866), .ZN(new_n912));
  NAND4_X1  g0712(.A1(new_n912), .A2(KEYINPUT40), .A3(new_n886), .A4(new_n903), .ZN(new_n913));
  NAND3_X1  g0713(.A1(new_n911), .A2(G330), .A3(new_n913), .ZN(new_n914));
  NAND3_X1  g0714(.A1(new_n867), .A2(G330), .A3(new_n453), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n906), .A2(new_n916), .ZN(new_n917));
  XNOR2_X1  g0717(.A(new_n917), .B(KEYINPUT107), .ZN(new_n918));
  INV_X1    g0718(.A(KEYINPUT39), .ZN(new_n919));
  NOR3_X1   g0719(.A1(new_n879), .A2(new_n880), .A3(new_n919), .ZN(new_n920));
  AOI21_X1  g0720(.A(new_n920), .B1(new_n919), .B2(new_n903), .ZN(new_n921));
  NOR2_X1   g0721(.A1(new_n354), .A2(new_n665), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  NOR2_X1   g0723(.A1(new_n821), .A2(new_n822), .ZN(new_n924));
  AOI21_X1  g0724(.A(KEYINPUT101), .B1(new_n733), .B2(new_n309), .ZN(new_n925));
  OAI21_X1  g0725(.A(new_n810), .B1(new_n924), .B2(new_n925), .ZN(new_n926));
  NAND3_X1  g0726(.A1(new_n926), .A2(new_n881), .A3(new_n886), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n633), .A2(new_n663), .ZN(new_n928));
  NAND3_X1  g0728(.A1(new_n923), .A2(new_n927), .A3(new_n928), .ZN(new_n929));
  XNOR2_X1  g0729(.A(new_n918), .B(new_n929), .ZN(new_n930));
  INV_X1    g0730(.A(KEYINPUT106), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n723), .A2(new_n735), .ZN(new_n932));
  AOI21_X1  g0732(.A(new_n931), .B1(new_n932), .B2(new_n453), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n724), .A2(new_n717), .ZN(new_n934));
  NAND4_X1  g0734(.A1(new_n934), .A2(new_n556), .A3(new_n716), .A4(new_n720), .ZN(new_n935));
  AOI21_X1  g0735(.A(new_n734), .B1(new_n935), .B2(new_n674), .ZN(new_n936));
  AOI211_X1 g0736(.A(KEYINPUT29), .B(new_n665), .C1(new_n730), .C2(new_n732), .ZN(new_n937));
  OAI211_X1 g0737(.A(new_n453), .B(new_n931), .C1(new_n936), .C2(new_n937), .ZN(new_n938));
  INV_X1    g0738(.A(new_n938), .ZN(new_n939));
  OAI21_X1  g0739(.A(new_n642), .B1(new_n933), .B2(new_n939), .ZN(new_n940));
  XNOR2_X1  g0740(.A(new_n930), .B(new_n940), .ZN(new_n941));
  OAI21_X1  g0741(.A(new_n941), .B1(new_n250), .B2(new_n659), .ZN(new_n942));
  NOR3_X1   g0742(.A1(new_n694), .A2(new_n331), .A3(new_n404), .ZN(new_n943));
  NOR2_X1   g0743(.A1(new_n203), .A2(G50), .ZN(new_n944));
  OAI211_X1 g0744(.A(G1), .B(new_n658), .C1(new_n943), .C2(new_n944), .ZN(new_n945));
  OAI211_X1 g0745(.A(G116), .B(new_n228), .C1(new_n497), .C2(KEYINPUT35), .ZN(new_n946));
  XNOR2_X1  g0746(.A(new_n946), .B(KEYINPUT103), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n497), .A2(KEYINPUT35), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  XNOR2_X1  g0749(.A(new_n949), .B(KEYINPUT104), .ZN(new_n950));
  XNOR2_X1  g0750(.A(new_n950), .B(KEYINPUT36), .ZN(new_n951));
  NAND3_X1  g0751(.A1(new_n942), .A2(new_n945), .A3(new_n951), .ZN(G367));
  NAND2_X1  g0752(.A1(new_n569), .A2(new_n665), .ZN(new_n953));
  NAND3_X1  g0753(.A1(new_n527), .A2(new_n572), .A3(new_n953), .ZN(new_n954));
  NOR2_X1   g0754(.A1(new_n684), .A2(new_n954), .ZN(new_n955));
  XNOR2_X1  g0755(.A(KEYINPUT110), .B(KEYINPUT42), .ZN(new_n956));
  XNOR2_X1  g0756(.A(new_n955), .B(new_n956), .ZN(new_n957));
  OAI21_X1  g0757(.A(new_n572), .B1(new_n954), .B2(new_n617), .ZN(new_n958));
  XOR2_X1   g0758(.A(new_n958), .B(KEYINPUT109), .Z(new_n959));
  OAI21_X1  g0759(.A(new_n957), .B1(new_n665), .B2(new_n959), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n536), .A2(new_n559), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n961), .A2(new_n665), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n561), .A2(new_n962), .ZN(new_n963));
  OR2_X1    g0763(.A1(new_n556), .A2(new_n962), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n963), .A2(new_n964), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n965), .A2(KEYINPUT43), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n960), .A2(new_n966), .ZN(new_n967));
  NOR2_X1   g0767(.A1(new_n965), .A2(KEYINPUT43), .ZN(new_n968));
  OR2_X1    g0768(.A1(new_n967), .A2(new_n968), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n967), .A2(new_n968), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n969), .A2(new_n970), .ZN(new_n971));
  INV_X1    g0771(.A(new_n682), .ZN(new_n972));
  NAND3_X1  g0772(.A1(new_n643), .A2(new_n571), .A3(new_n665), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n973), .A2(new_n954), .ZN(new_n974));
  INV_X1    g0774(.A(new_n974), .ZN(new_n975));
  OAI21_X1  g0775(.A(new_n971), .B1(new_n972), .B2(new_n975), .ZN(new_n976));
  NAND4_X1  g0776(.A1(new_n970), .A2(new_n682), .A3(new_n974), .A4(new_n969), .ZN(new_n977));
  XNOR2_X1  g0777(.A(KEYINPUT111), .B(KEYINPUT41), .ZN(new_n978));
  XOR2_X1   g0778(.A(new_n690), .B(new_n978), .Z(new_n979));
  NAND3_X1  g0779(.A1(new_n684), .A2(new_n685), .A3(new_n974), .ZN(new_n980));
  AND2_X1   g0780(.A1(new_n980), .A2(KEYINPUT112), .ZN(new_n981));
  NOR2_X1   g0781(.A1(new_n980), .A2(KEYINPUT112), .ZN(new_n982));
  INV_X1    g0782(.A(KEYINPUT45), .ZN(new_n983));
  OR3_X1    g0783(.A1(new_n981), .A2(new_n982), .A3(new_n983), .ZN(new_n984));
  AOI21_X1  g0784(.A(new_n974), .B1(new_n684), .B2(new_n685), .ZN(new_n985));
  XNOR2_X1  g0785(.A(new_n985), .B(KEYINPUT44), .ZN(new_n986));
  OAI21_X1  g0786(.A(new_n983), .B1(new_n981), .B2(new_n982), .ZN(new_n987));
  NAND3_X1  g0787(.A1(new_n984), .A2(new_n986), .A3(new_n987), .ZN(new_n988));
  NAND2_X1  g0788(.A1(new_n988), .A2(new_n682), .ZN(new_n989));
  NAND4_X1  g0789(.A1(new_n984), .A2(new_n972), .A3(new_n986), .A4(new_n987), .ZN(new_n990));
  OAI21_X1  g0790(.A(new_n676), .B1(new_n488), .B2(new_n665), .ZN(new_n991));
  NAND2_X1  g0791(.A1(new_n991), .A2(new_n684), .ZN(new_n992));
  XNOR2_X1  g0792(.A(new_n992), .B(new_n681), .ZN(new_n993));
  NOR2_X1   g0793(.A1(new_n993), .A2(new_n736), .ZN(new_n994));
  NAND3_X1  g0794(.A1(new_n989), .A2(new_n990), .A3(new_n994), .ZN(new_n995));
  AOI21_X1  g0795(.A(new_n979), .B1(new_n995), .B2(new_n737), .ZN(new_n996));
  OAI211_X1 g0796(.A(new_n976), .B(new_n977), .C1(new_n996), .C2(new_n743), .ZN(new_n997));
  OAI21_X1  g0797(.A(new_n292), .B1(new_n758), .B2(new_n838), .ZN(new_n998));
  AOI22_X1  g0798(.A1(G159), .A2(new_n784), .B1(new_n789), .B2(G50), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n771), .A2(G68), .ZN(new_n1000));
  INV_X1    g0800(.A(new_n836), .ZN(new_n1001));
  OAI211_X1 g0801(.A(new_n999), .B(new_n1000), .C1(new_n763), .C2(new_n1001), .ZN(new_n1002));
  AOI211_X1 g0802(.A(new_n998), .B(new_n1002), .C1(G58), .C2(new_n768), .ZN(new_n1003));
  OAI221_X1 g0803(.A(new_n1003), .B1(new_n331), .B2(new_n778), .C1(new_n358), .C2(new_n754), .ZN(new_n1004));
  INV_X1    g0804(.A(G294), .ZN(new_n1005));
  NOR2_X1   g0805(.A1(new_n774), .A2(new_n1005), .ZN(new_n1006));
  OAI21_X1  g0806(.A(KEYINPUT114), .B1(new_n767), .B2(new_n455), .ZN(new_n1007));
  XOR2_X1   g0807(.A(new_n1007), .B(KEYINPUT46), .Z(new_n1008));
  XNOR2_X1  g0808(.A(KEYINPUT113), .B(G311), .ZN(new_n1009));
  OAI221_X1 g0809(.A(new_n1008), .B1(new_n296), .B2(new_n782), .C1(new_n763), .C2(new_n1009), .ZN(new_n1010));
  AOI211_X1 g0810(.A(new_n1006), .B(new_n1010), .C1(G317), .C2(new_n759), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n779), .A2(G97), .ZN(new_n1012));
  NAND2_X1  g0812(.A1(new_n755), .A2(G303), .ZN(new_n1013));
  NAND3_X1  g0813(.A1(new_n1011), .A2(new_n1012), .A3(new_n1013), .ZN(new_n1014));
  OAI21_X1  g0814(.A(new_n376), .B1(new_n775), .B2(new_n850), .ZN(new_n1015));
  OAI21_X1  g0815(.A(new_n1004), .B1(new_n1014), .B2(new_n1015), .ZN(new_n1016));
  XNOR2_X1  g0816(.A(new_n1016), .B(KEYINPUT47), .ZN(new_n1017));
  NAND2_X1  g0817(.A1(new_n1017), .A2(new_n796), .ZN(new_n1018));
  NAND3_X1  g0818(.A1(new_n963), .A2(new_n750), .A3(new_n964), .ZN(new_n1019));
  INV_X1    g0819(.A(new_n800), .ZN(new_n1020));
  OAI221_X1 g0820(.A(new_n805), .B1(new_n210), .B2(new_n535), .C1(new_n239), .C2(new_n1020), .ZN(new_n1021));
  NAND4_X1  g0821(.A1(new_n1018), .A2(new_n744), .A3(new_n1019), .A4(new_n1021), .ZN(new_n1022));
  NAND2_X1  g0822(.A1(new_n997), .A2(new_n1022), .ZN(G387));
  INV_X1    g0823(.A(new_n994), .ZN(new_n1024));
  AOI21_X1  g0824(.A(new_n691), .B1(new_n993), .B2(new_n736), .ZN(new_n1025));
  NAND2_X1  g0825(.A1(new_n1024), .A2(new_n1025), .ZN(new_n1026));
  OAI21_X1  g0826(.A(new_n1012), .B1(new_n203), .B2(new_n775), .ZN(new_n1027));
  AOI211_X1 g0827(.A(new_n376), .B(new_n1027), .C1(G150), .C2(new_n759), .ZN(new_n1028));
  NAND2_X1  g0828(.A1(new_n771), .A2(new_n259), .ZN(new_n1029));
  NAND2_X1  g0829(.A1(new_n764), .A2(G159), .ZN(new_n1030));
  OR2_X1    g0830(.A1(new_n1030), .A2(KEYINPUT116), .ZN(new_n1031));
  NOR2_X1   g0831(.A1(new_n767), .A2(new_n331), .ZN(new_n1032));
  OAI22_X1  g0832(.A1(new_n201), .A2(new_n754), .B1(new_n774), .B2(new_n253), .ZN(new_n1033));
  AOI211_X1 g0833(.A(new_n1032), .B(new_n1033), .C1(KEYINPUT116), .C2(new_n1030), .ZN(new_n1034));
  NAND4_X1  g0834(.A1(new_n1028), .A2(new_n1029), .A3(new_n1031), .A4(new_n1034), .ZN(new_n1035));
  AOI22_X1  g0835(.A1(new_n764), .A2(G322), .B1(new_n789), .B2(G303), .ZN(new_n1036));
  INV_X1    g0836(.A(G317), .ZN(new_n1037));
  OAI221_X1 g0837(.A(new_n1036), .B1(new_n1037), .B2(new_n754), .C1(new_n774), .C2(new_n1009), .ZN(new_n1038));
  XNOR2_X1  g0838(.A(new_n1038), .B(KEYINPUT48), .ZN(new_n1039));
  OAI221_X1 g0839(.A(new_n1039), .B1(new_n850), .B2(new_n782), .C1(new_n1005), .C2(new_n767), .ZN(new_n1040));
  XOR2_X1   g0840(.A(new_n1040), .B(KEYINPUT49), .Z(new_n1041));
  AOI21_X1  g0841(.A(new_n292), .B1(new_n759), .B2(G326), .ZN(new_n1042));
  OAI21_X1  g0842(.A(new_n1042), .B1(new_n455), .B2(new_n778), .ZN(new_n1043));
  OAI21_X1  g0843(.A(new_n1035), .B1(new_n1041), .B2(new_n1043), .ZN(new_n1044));
  NAND2_X1  g0844(.A1(new_n1044), .A2(new_n796), .ZN(new_n1045));
  AND2_X1   g0845(.A1(new_n236), .A2(G45), .ZN(new_n1046));
  OAI22_X1  g0846(.A1(new_n1046), .A2(new_n1020), .B1(new_n692), .B2(new_n803), .ZN(new_n1047));
  NAND2_X1  g0847(.A1(new_n255), .A2(new_n201), .ZN(new_n1048));
  XOR2_X1   g0848(.A(new_n1048), .B(KEYINPUT50), .Z(new_n1049));
  AOI21_X1  g0849(.A(G45), .B1(G68), .B2(G77), .ZN(new_n1050));
  NAND3_X1  g0850(.A1(new_n1049), .A2(new_n692), .A3(new_n1050), .ZN(new_n1051));
  AOI22_X1  g0851(.A1(new_n1047), .A2(new_n1051), .B1(new_n296), .B2(new_n689), .ZN(new_n1052));
  INV_X1    g0852(.A(new_n805), .ZN(new_n1053));
  OAI21_X1  g0853(.A(new_n744), .B1(new_n1052), .B2(new_n1053), .ZN(new_n1054));
  XNOR2_X1  g0854(.A(new_n1054), .B(KEYINPUT115), .ZN(new_n1055));
  NAND2_X1  g0855(.A1(new_n1045), .A2(new_n1055), .ZN(new_n1056));
  OR2_X1    g0856(.A1(new_n1056), .A2(KEYINPUT117), .ZN(new_n1057));
  NAND2_X1  g0857(.A1(new_n676), .A2(new_n750), .ZN(new_n1058));
  NAND2_X1  g0858(.A1(new_n1056), .A2(KEYINPUT117), .ZN(new_n1059));
  NAND3_X1  g0859(.A1(new_n1057), .A2(new_n1058), .A3(new_n1059), .ZN(new_n1060));
  OAI211_X1 g0860(.A(new_n1026), .B(new_n1060), .C1(new_n742), .C2(new_n993), .ZN(G393));
  NAND2_X1  g0861(.A1(new_n989), .A2(new_n990), .ZN(new_n1062));
  NAND2_X1  g0862(.A1(new_n1062), .A2(new_n1024), .ZN(new_n1063));
  NAND3_X1  g0863(.A1(new_n1063), .A2(new_n690), .A3(new_n995), .ZN(new_n1064));
  NAND3_X1  g0864(.A1(new_n989), .A2(new_n743), .A3(new_n990), .ZN(new_n1065));
  AOI21_X1  g0865(.A(new_n745), .B1(new_n975), .B2(new_n750), .ZN(new_n1066));
  OAI221_X1 g0866(.A(new_n805), .B1(new_n315), .B2(new_n210), .C1(new_n248), .C2(new_n1020), .ZN(new_n1067));
  NAND2_X1  g0867(.A1(new_n255), .A2(new_n789), .ZN(new_n1068));
  OAI21_X1  g0868(.A(new_n1068), .B1(new_n758), .B2(new_n1001), .ZN(new_n1069));
  AOI21_X1  g0869(.A(new_n1069), .B1(G68), .B2(new_n768), .ZN(new_n1070));
  NAND2_X1  g0870(.A1(new_n771), .A2(G77), .ZN(new_n1071));
  INV_X1    g0871(.A(G159), .ZN(new_n1072));
  OAI22_X1  g0872(.A1(new_n763), .A2(new_n358), .B1(new_n754), .B2(new_n1072), .ZN(new_n1073));
  XNOR2_X1  g0873(.A(new_n1073), .B(KEYINPUT51), .ZN(new_n1074));
  AOI211_X1 g0874(.A(new_n376), .B(new_n849), .C1(G50), .C2(new_n784), .ZN(new_n1075));
  NAND4_X1  g0875(.A1(new_n1070), .A2(new_n1071), .A3(new_n1074), .A4(new_n1075), .ZN(new_n1076));
  OAI22_X1  g0876(.A1(new_n763), .A2(new_n1037), .B1(new_n754), .B2(new_n776), .ZN(new_n1077));
  XNOR2_X1  g0877(.A(new_n1077), .B(KEYINPUT52), .ZN(new_n1078));
  OAI22_X1  g0878(.A1(new_n782), .A2(new_n455), .B1(new_n767), .B2(new_n850), .ZN(new_n1079));
  AOI21_X1  g0879(.A(new_n1079), .B1(G294), .B2(new_n789), .ZN(new_n1080));
  AOI21_X1  g0880(.A(new_n292), .B1(new_n759), .B2(G322), .ZN(new_n1081));
  AOI22_X1  g0881(.A1(G303), .A2(new_n784), .B1(new_n779), .B2(G107), .ZN(new_n1082));
  NAND4_X1  g0882(.A1(new_n1078), .A2(new_n1080), .A3(new_n1081), .A4(new_n1082), .ZN(new_n1083));
  AND2_X1   g0883(.A1(new_n1076), .A2(new_n1083), .ZN(new_n1084));
  OAI211_X1 g0884(.A(new_n1066), .B(new_n1067), .C1(new_n833), .C2(new_n1084), .ZN(new_n1085));
  AND2_X1   g0885(.A1(new_n1065), .A2(new_n1085), .ZN(new_n1086));
  NAND2_X1  g0886(.A1(new_n1064), .A2(new_n1086), .ZN(G390));
  INV_X1    g0887(.A(new_n309), .ZN(new_n1088));
  OAI21_X1  g0888(.A(new_n810), .B1(new_n722), .B2(new_n1088), .ZN(new_n1089));
  NAND2_X1  g0889(.A1(new_n1089), .A2(new_n886), .ZN(new_n1090));
  INV_X1    g0890(.A(new_n922), .ZN(new_n1091));
  NAND3_X1  g0891(.A1(new_n1090), .A2(new_n1091), .A3(new_n903), .ZN(new_n1092));
  AOI21_X1  g0892(.A(new_n922), .B1(new_n926), .B2(new_n886), .ZN(new_n1093));
  OAI21_X1  g0893(.A(new_n1092), .B1(new_n1093), .B2(new_n921), .ZN(new_n1094));
  NOR2_X1   g0894(.A1(new_n909), .A2(new_n740), .ZN(new_n1095));
  INV_X1    g0895(.A(new_n1095), .ZN(new_n1096));
  NAND2_X1  g0896(.A1(new_n1094), .A2(new_n1096), .ZN(new_n1097));
  NOR3_X1   g0897(.A1(new_n715), .A2(new_n814), .A3(new_n885), .ZN(new_n1098));
  OAI211_X1 g0898(.A(new_n1092), .B(new_n1098), .C1(new_n1093), .C2(new_n921), .ZN(new_n1099));
  INV_X1    g0899(.A(new_n1089), .ZN(new_n1100));
  OAI211_X1 g0900(.A(G330), .B(new_n817), .C1(new_n907), .C2(new_n908), .ZN(new_n1101));
  AOI21_X1  g0901(.A(new_n1098), .B1(new_n1101), .B2(new_n885), .ZN(new_n1102));
  OAI21_X1  g0902(.A(new_n885), .B1(new_n715), .B2(new_n814), .ZN(new_n1103));
  OAI21_X1  g0903(.A(new_n1103), .B1(new_n909), .B2(new_n740), .ZN(new_n1104));
  AOI22_X1  g0904(.A1(new_n1100), .A2(new_n1102), .B1(new_n1104), .B2(new_n926), .ZN(new_n1105));
  OAI211_X1 g0905(.A(new_n642), .B(new_n915), .C1(new_n933), .C2(new_n939), .ZN(new_n1106));
  OAI211_X1 g0906(.A(new_n1097), .B(new_n1099), .C1(new_n1105), .C2(new_n1106), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n903), .A2(new_n919), .ZN(new_n1108));
  INV_X1    g0908(.A(new_n920), .ZN(new_n1109));
  NAND2_X1  g0909(.A1(new_n1108), .A2(new_n1109), .ZN(new_n1110));
  AOI21_X1  g0910(.A(new_n809), .B1(new_n823), .B2(new_n824), .ZN(new_n1111));
  OAI21_X1  g0911(.A(new_n1091), .B1(new_n1111), .B2(new_n885), .ZN(new_n1112));
  AND2_X1   g0912(.A1(new_n903), .A2(new_n1091), .ZN(new_n1113));
  AOI22_X1  g0913(.A1(new_n1110), .A2(new_n1112), .B1(new_n1090), .B2(new_n1113), .ZN(new_n1114));
  OAI21_X1  g0914(.A(new_n1099), .B1(new_n1114), .B2(new_n1095), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n1104), .A2(new_n926), .ZN(new_n1116));
  NAND2_X1  g0916(.A1(new_n1101), .A2(new_n885), .ZN(new_n1117));
  INV_X1    g0917(.A(new_n1098), .ZN(new_n1118));
  NAND3_X1  g0918(.A1(new_n1117), .A2(new_n1100), .A3(new_n1118), .ZN(new_n1119));
  AOI21_X1  g0919(.A(new_n1106), .B1(new_n1116), .B2(new_n1119), .ZN(new_n1120));
  NAND2_X1  g0920(.A1(new_n1115), .A2(new_n1120), .ZN(new_n1121));
  NAND3_X1  g0921(.A1(new_n1107), .A2(new_n1121), .A3(new_n690), .ZN(new_n1122));
  OAI21_X1  g0922(.A(new_n744), .B1(new_n921), .B2(new_n749), .ZN(new_n1123));
  AND2_X1   g0923(.A1(new_n857), .A2(new_n253), .ZN(new_n1124));
  INV_X1    g0924(.A(G128), .ZN(new_n1125));
  OAI22_X1  g0925(.A1(new_n763), .A2(new_n1125), .B1(new_n754), .B2(new_n834), .ZN(new_n1126));
  INV_X1    g0926(.A(KEYINPUT53), .ZN(new_n1127));
  AOI21_X1  g0927(.A(new_n1127), .B1(new_n768), .B2(G150), .ZN(new_n1128));
  XOR2_X1   g0928(.A(KEYINPUT54), .B(G143), .Z(new_n1129));
  AOI211_X1 g0929(.A(new_n1126), .B(new_n1128), .C1(new_n789), .C2(new_n1129), .ZN(new_n1130));
  INV_X1    g0930(.A(G125), .ZN(new_n1131));
  OAI22_X1  g0931(.A1(new_n774), .A2(new_n838), .B1(new_n758), .B2(new_n1131), .ZN(new_n1132));
  AOI211_X1 g0932(.A(new_n376), .B(new_n1132), .C1(G50), .C2(new_n779), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n771), .A2(G159), .ZN(new_n1134));
  NAND3_X1  g0934(.A1(new_n768), .A2(new_n1127), .A3(G150), .ZN(new_n1135));
  NAND4_X1  g0935(.A1(new_n1130), .A2(new_n1133), .A3(new_n1134), .A4(new_n1135), .ZN(new_n1136));
  OAI21_X1  g0936(.A(new_n376), .B1(new_n767), .B2(new_n214), .ZN(new_n1137));
  XOR2_X1   g0937(.A(new_n1137), .B(KEYINPUT118), .Z(new_n1138));
  OAI22_X1  g0938(.A1(new_n754), .A2(new_n455), .B1(new_n758), .B2(new_n1005), .ZN(new_n1139));
  AOI211_X1 g0939(.A(new_n842), .B(new_n1139), .C1(G107), .C2(new_n784), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n789), .A2(G97), .ZN(new_n1141));
  AOI22_X1  g0941(.A1(new_n764), .A2(G283), .B1(new_n771), .B2(G77), .ZN(new_n1142));
  NAND4_X1  g0942(.A1(new_n1138), .A2(new_n1140), .A3(new_n1141), .A4(new_n1142), .ZN(new_n1143));
  AOI21_X1  g0943(.A(new_n833), .B1(new_n1136), .B2(new_n1143), .ZN(new_n1144));
  NOR3_X1   g0944(.A1(new_n1123), .A2(new_n1124), .A3(new_n1144), .ZN(new_n1145));
  AOI21_X1  g0945(.A(new_n1145), .B1(new_n1115), .B2(new_n743), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n1122), .A2(new_n1146), .ZN(G378));
  NAND2_X1  g0947(.A1(new_n392), .A2(new_n395), .ZN(new_n1148));
  NOR3_X1   g0948(.A1(new_n371), .A2(new_n366), .A3(new_n663), .ZN(new_n1149));
  XNOR2_X1  g0949(.A(new_n1148), .B(new_n1149), .ZN(new_n1150));
  XNOR2_X1  g0950(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1151));
  XOR2_X1   g0951(.A(new_n1150), .B(new_n1151), .Z(new_n1152));
  INV_X1    g0952(.A(new_n1152), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n1153), .A2(new_n748), .ZN(new_n1154));
  NAND2_X1  g0954(.A1(new_n779), .A2(G58), .ZN(new_n1155));
  XNOR2_X1  g0955(.A(new_n1155), .B(KEYINPUT119), .ZN(new_n1156));
  OAI211_X1 g0956(.A(new_n1156), .B(new_n277), .C1(new_n331), .C2(new_n767), .ZN(new_n1157));
  AOI21_X1  g0957(.A(new_n1157), .B1(G97), .B2(new_n784), .ZN(new_n1158));
  OAI221_X1 g0958(.A(new_n1000), .B1(new_n296), .B2(new_n754), .C1(new_n455), .C2(new_n763), .ZN(new_n1159));
  AOI211_X1 g0959(.A(new_n292), .B(new_n1159), .C1(new_n259), .C2(new_n789), .ZN(new_n1160));
  OAI211_X1 g0960(.A(new_n1158), .B(new_n1160), .C1(new_n850), .C2(new_n758), .ZN(new_n1161));
  XOR2_X1   g0961(.A(new_n1161), .B(KEYINPUT58), .Z(new_n1162));
  OAI21_X1  g0962(.A(new_n201), .B1(new_n374), .B2(G41), .ZN(new_n1163));
  OAI22_X1  g0963(.A1(new_n782), .A2(new_n358), .B1(new_n763), .B2(new_n1131), .ZN(new_n1164));
  AOI22_X1  g0964(.A1(G132), .A2(new_n784), .B1(new_n789), .B2(G137), .ZN(new_n1165));
  OAI21_X1  g0965(.A(new_n1165), .B1(new_n1125), .B2(new_n754), .ZN(new_n1166));
  AOI211_X1 g0966(.A(new_n1164), .B(new_n1166), .C1(new_n768), .C2(new_n1129), .ZN(new_n1167));
  INV_X1    g0967(.A(KEYINPUT59), .ZN(new_n1168));
  AOI21_X1  g0968(.A(G33), .B1(new_n1167), .B2(new_n1168), .ZN(new_n1169));
  AOI21_X1  g0969(.A(G41), .B1(new_n759), .B2(G124), .ZN(new_n1170));
  OAI211_X1 g0970(.A(new_n1169), .B(new_n1170), .C1(new_n1072), .C2(new_n778), .ZN(new_n1171));
  NOR2_X1   g0971(.A1(new_n1167), .A2(new_n1168), .ZN(new_n1172));
  OAI21_X1  g0972(.A(new_n1163), .B1(new_n1171), .B2(new_n1172), .ZN(new_n1173));
  OAI21_X1  g0973(.A(new_n796), .B1(new_n1162), .B2(new_n1173), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n857), .A2(new_n201), .ZN(new_n1175));
  NAND4_X1  g0975(.A1(new_n1154), .A2(new_n744), .A3(new_n1174), .A4(new_n1175), .ZN(new_n1176));
  INV_X1    g0976(.A(new_n1176), .ZN(new_n1177));
  AOI21_X1  g0977(.A(new_n1152), .B1(new_n905), .B2(G330), .ZN(new_n1178));
  AND4_X1   g0978(.A1(G330), .A2(new_n911), .A3(new_n1152), .A4(new_n913), .ZN(new_n1179));
  OAI21_X1  g0979(.A(new_n929), .B1(new_n1178), .B2(new_n1179), .ZN(new_n1180));
  INV_X1    g0980(.A(new_n929), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n914), .A2(new_n1153), .ZN(new_n1182));
  NAND4_X1  g0982(.A1(new_n911), .A2(new_n1152), .A3(G330), .A4(new_n913), .ZN(new_n1183));
  NAND3_X1  g0983(.A1(new_n1181), .A2(new_n1182), .A3(new_n1183), .ZN(new_n1184));
  NAND2_X1  g0984(.A1(new_n1180), .A2(new_n1184), .ZN(new_n1185));
  AOI21_X1  g0985(.A(new_n1177), .B1(new_n1185), .B2(new_n743), .ZN(new_n1186));
  INV_X1    g0986(.A(new_n1106), .ZN(new_n1187));
  AOI22_X1  g0987(.A1(new_n1180), .A2(new_n1184), .B1(new_n1121), .B2(new_n1187), .ZN(new_n1188));
  OAI21_X1  g0988(.A(new_n690), .B1(new_n1188), .B2(KEYINPUT57), .ZN(new_n1189));
  NAND3_X1  g0989(.A1(new_n1180), .A2(KEYINPUT120), .A3(new_n1184), .ZN(new_n1190));
  AOI21_X1  g0990(.A(new_n1181), .B1(new_n1182), .B2(new_n1183), .ZN(new_n1191));
  INV_X1    g0991(.A(KEYINPUT120), .ZN(new_n1192));
  NAND2_X1  g0992(.A1(new_n1191), .A2(new_n1192), .ZN(new_n1193));
  INV_X1    g0993(.A(KEYINPUT57), .ZN(new_n1194));
  AOI21_X1  g0994(.A(new_n1194), .B1(new_n1121), .B2(new_n1187), .ZN(new_n1195));
  AND3_X1   g0995(.A1(new_n1190), .A2(new_n1193), .A3(new_n1195), .ZN(new_n1196));
  OAI21_X1  g0996(.A(new_n1186), .B1(new_n1189), .B2(new_n1196), .ZN(G375));
  NAND2_X1  g0997(.A1(new_n1116), .A2(new_n1119), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(new_n1198), .A2(new_n1187), .ZN(new_n1199));
  INV_X1    g0999(.A(new_n979), .ZN(new_n1200));
  NAND3_X1  g1000(.A1(new_n1116), .A2(new_n1106), .A3(new_n1119), .ZN(new_n1201));
  NAND3_X1  g1001(.A1(new_n1199), .A2(new_n1200), .A3(new_n1201), .ZN(new_n1202));
  OAI221_X1 g1002(.A(new_n1156), .B1(new_n201), .B2(new_n782), .C1(new_n834), .C2(new_n763), .ZN(new_n1203));
  AND2_X1   g1003(.A1(new_n784), .A2(new_n1129), .ZN(new_n1204));
  OAI22_X1  g1004(.A1(new_n775), .A2(new_n358), .B1(new_n758), .B2(new_n1125), .ZN(new_n1205));
  OAI221_X1 g1005(.A(new_n292), .B1(new_n754), .B2(new_n838), .C1(new_n1072), .C2(new_n767), .ZN(new_n1206));
  NOR4_X1   g1006(.A1(new_n1203), .A2(new_n1204), .A3(new_n1205), .A4(new_n1206), .ZN(new_n1207));
  AOI21_X1  g1007(.A(new_n292), .B1(new_n759), .B2(G303), .ZN(new_n1208));
  OAI221_X1 g1008(.A(new_n1208), .B1(new_n331), .B2(new_n778), .C1(new_n455), .C2(new_n774), .ZN(new_n1209));
  NOR2_X1   g1009(.A1(new_n767), .A2(new_n315), .ZN(new_n1210));
  OAI22_X1  g1010(.A1(new_n754), .A2(new_n850), .B1(new_n775), .B2(new_n296), .ZN(new_n1211));
  OAI21_X1  g1011(.A(new_n1029), .B1(new_n1005), .B2(new_n763), .ZN(new_n1212));
  NOR4_X1   g1012(.A1(new_n1209), .A2(new_n1210), .A3(new_n1211), .A4(new_n1212), .ZN(new_n1213));
  OAI21_X1  g1013(.A(new_n796), .B1(new_n1207), .B2(new_n1213), .ZN(new_n1214));
  OAI211_X1 g1014(.A(new_n744), .B(new_n1214), .C1(new_n886), .C2(new_n749), .ZN(new_n1215));
  AOI21_X1  g1015(.A(new_n1215), .B1(new_n203), .B2(new_n857), .ZN(new_n1216));
  AOI21_X1  g1016(.A(new_n1216), .B1(new_n1198), .B2(new_n743), .ZN(new_n1217));
  NAND2_X1  g1017(.A1(new_n1202), .A2(new_n1217), .ZN(G381));
  NAND2_X1  g1018(.A1(new_n1185), .A2(new_n743), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(new_n1219), .A2(new_n1176), .ZN(new_n1220));
  NAND2_X1  g1020(.A1(new_n1121), .A2(new_n1187), .ZN(new_n1221));
  NOR3_X1   g1021(.A1(new_n1178), .A2(new_n1179), .A3(new_n929), .ZN(new_n1222));
  OAI21_X1  g1022(.A(new_n1221), .B1(new_n1222), .B2(new_n1191), .ZN(new_n1223));
  AOI21_X1  g1023(.A(new_n691), .B1(new_n1223), .B2(new_n1194), .ZN(new_n1224));
  NAND3_X1  g1024(.A1(new_n1190), .A2(new_n1193), .A3(new_n1195), .ZN(new_n1225));
  AOI21_X1  g1025(.A(new_n1220), .B1(new_n1224), .B2(new_n1225), .ZN(new_n1226));
  INV_X1    g1026(.A(KEYINPUT122), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(G378), .A2(new_n1227), .ZN(new_n1228));
  NAND3_X1  g1028(.A1(new_n1122), .A2(KEYINPUT122), .A3(new_n1146), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n1228), .A2(new_n1229), .ZN(new_n1230));
  AND2_X1   g1030(.A1(new_n1226), .A2(new_n1230), .ZN(new_n1231));
  NOR3_X1   g1031(.A1(G393), .A2(G396), .A3(G384), .ZN(new_n1232));
  XOR2_X1   g1032(.A(new_n1232), .B(KEYINPUT121), .Z(new_n1233));
  INV_X1    g1033(.A(G387), .ZN(new_n1234));
  NOR2_X1   g1034(.A1(G390), .A2(G381), .ZN(new_n1235));
  NAND4_X1  g1035(.A1(new_n1231), .A2(new_n1233), .A3(new_n1234), .A4(new_n1235), .ZN(G407));
  NAND2_X1  g1036(.A1(new_n664), .A2(G213), .ZN(new_n1237));
  INV_X1    g1037(.A(new_n1237), .ZN(new_n1238));
  NAND3_X1  g1038(.A1(new_n1231), .A2(KEYINPUT123), .A3(new_n1238), .ZN(new_n1239));
  NAND3_X1  g1039(.A1(G407), .A2(G213), .A3(new_n1239), .ZN(new_n1240));
  AOI21_X1  g1040(.A(KEYINPUT123), .B1(new_n1231), .B2(new_n1238), .ZN(new_n1241));
  OR2_X1    g1041(.A1(new_n1240), .A2(new_n1241), .ZN(G409));
  OAI211_X1 g1042(.A(G378), .B(new_n1186), .C1(new_n1189), .C2(new_n1196), .ZN(new_n1243));
  NAND3_X1  g1043(.A1(new_n1190), .A2(new_n743), .A3(new_n1193), .ZN(new_n1244));
  NAND3_X1  g1044(.A1(new_n1185), .A2(new_n1200), .A3(new_n1221), .ZN(new_n1245));
  NAND3_X1  g1045(.A1(new_n1244), .A2(new_n1176), .A3(new_n1245), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(new_n1230), .A2(new_n1246), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n1243), .A2(new_n1247), .ZN(new_n1248));
  INV_X1    g1048(.A(KEYINPUT60), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n1201), .A2(new_n1249), .ZN(new_n1250));
  NAND4_X1  g1050(.A1(new_n1116), .A2(new_n1119), .A3(new_n1106), .A4(KEYINPUT60), .ZN(new_n1251));
  NAND4_X1  g1051(.A1(new_n1250), .A2(new_n1199), .A3(new_n690), .A4(new_n1251), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(new_n1252), .A2(new_n1217), .ZN(new_n1253));
  INV_X1    g1053(.A(KEYINPUT124), .ZN(new_n1254));
  NAND2_X1  g1054(.A1(G384), .A2(new_n1254), .ZN(new_n1255));
  INV_X1    g1055(.A(G384), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(new_n1256), .A2(KEYINPUT124), .ZN(new_n1257));
  NAND3_X1  g1057(.A1(new_n1253), .A2(new_n1255), .A3(new_n1257), .ZN(new_n1258));
  NAND4_X1  g1058(.A1(new_n1252), .A2(KEYINPUT124), .A3(new_n1256), .A4(new_n1217), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(new_n1258), .A2(new_n1259), .ZN(new_n1260));
  NAND3_X1  g1060(.A1(new_n1248), .A2(new_n1237), .A3(new_n1260), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(new_n1261), .A2(KEYINPUT62), .ZN(new_n1262));
  INV_X1    g1062(.A(KEYINPUT61), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n1238), .A2(G2897), .ZN(new_n1264));
  XOR2_X1   g1064(.A(new_n1264), .B(KEYINPUT125), .Z(new_n1265));
  NAND2_X1  g1065(.A1(new_n1260), .A2(new_n1265), .ZN(new_n1266));
  INV_X1    g1066(.A(new_n1265), .ZN(new_n1267));
  NAND3_X1  g1067(.A1(new_n1258), .A2(new_n1259), .A3(new_n1267), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1266), .A2(new_n1268), .ZN(new_n1269));
  INV_X1    g1069(.A(new_n1269), .ZN(new_n1270));
  AOI22_X1  g1070(.A1(new_n1226), .A2(G378), .B1(new_n1230), .B2(new_n1246), .ZN(new_n1271));
  OAI21_X1  g1071(.A(new_n1270), .B1(new_n1271), .B2(new_n1238), .ZN(new_n1272));
  AOI21_X1  g1072(.A(new_n1238), .B1(new_n1243), .B2(new_n1247), .ZN(new_n1273));
  INV_X1    g1073(.A(KEYINPUT62), .ZN(new_n1274));
  NAND3_X1  g1074(.A1(new_n1273), .A2(new_n1274), .A3(new_n1260), .ZN(new_n1275));
  NAND4_X1  g1075(.A1(new_n1262), .A2(new_n1263), .A3(new_n1272), .A4(new_n1275), .ZN(new_n1276));
  INV_X1    g1076(.A(G390), .ZN(new_n1277));
  INV_X1    g1077(.A(G396), .ZN(new_n1278));
  XNOR2_X1  g1078(.A(G393), .B(new_n1278), .ZN(new_n1279));
  AOI21_X1  g1079(.A(new_n1279), .B1(G387), .B2(KEYINPUT126), .ZN(new_n1280));
  XNOR2_X1  g1080(.A(G393), .B(G396), .ZN(new_n1281));
  AOI21_X1  g1081(.A(new_n1281), .B1(new_n997), .B2(new_n1022), .ZN(new_n1282));
  OAI21_X1  g1082(.A(new_n1277), .B1(new_n1280), .B2(new_n1282), .ZN(new_n1283));
  NAND2_X1  g1083(.A1(G387), .A2(new_n1279), .ZN(new_n1284));
  INV_X1    g1084(.A(KEYINPUT126), .ZN(new_n1285));
  AOI21_X1  g1085(.A(new_n1285), .B1(new_n997), .B2(new_n1022), .ZN(new_n1286));
  OAI211_X1 g1086(.A(new_n1284), .B(G390), .C1(new_n1279), .C2(new_n1286), .ZN(new_n1287));
  NAND2_X1  g1087(.A1(new_n1283), .A2(new_n1287), .ZN(new_n1288));
  INV_X1    g1088(.A(new_n1288), .ZN(new_n1289));
  NAND2_X1  g1089(.A1(new_n1276), .A2(new_n1289), .ZN(new_n1290));
  AOI21_X1  g1090(.A(new_n1269), .B1(new_n1248), .B2(new_n1237), .ZN(new_n1291));
  INV_X1    g1091(.A(KEYINPUT63), .ZN(new_n1292));
  OAI21_X1  g1092(.A(new_n1261), .B1(new_n1291), .B2(new_n1292), .ZN(new_n1293));
  AOI21_X1  g1093(.A(KEYINPUT61), .B1(new_n1283), .B2(new_n1287), .ZN(new_n1294));
  INV_X1    g1094(.A(KEYINPUT127), .ZN(new_n1295));
  OAI21_X1  g1095(.A(new_n1295), .B1(new_n1261), .B2(new_n1292), .ZN(new_n1296));
  NAND4_X1  g1096(.A1(new_n1273), .A2(KEYINPUT127), .A3(KEYINPUT63), .A4(new_n1260), .ZN(new_n1297));
  NAND4_X1  g1097(.A1(new_n1293), .A2(new_n1294), .A3(new_n1296), .A4(new_n1297), .ZN(new_n1298));
  NAND2_X1  g1098(.A1(new_n1290), .A2(new_n1298), .ZN(G405));
  NAND2_X1  g1099(.A1(G375), .A2(new_n1230), .ZN(new_n1300));
  AND2_X1   g1100(.A1(new_n1300), .A2(new_n1243), .ZN(new_n1301));
  NOR2_X1   g1101(.A1(new_n1301), .A2(new_n1260), .ZN(new_n1302));
  INV_X1    g1102(.A(new_n1302), .ZN(new_n1303));
  NAND3_X1  g1103(.A1(new_n1300), .A2(new_n1243), .A3(new_n1260), .ZN(new_n1304));
  NAND3_X1  g1104(.A1(new_n1303), .A2(new_n1289), .A3(new_n1304), .ZN(new_n1305));
  INV_X1    g1105(.A(new_n1304), .ZN(new_n1306));
  OAI21_X1  g1106(.A(new_n1288), .B1(new_n1302), .B2(new_n1306), .ZN(new_n1307));
  NAND2_X1  g1107(.A1(new_n1305), .A2(new_n1307), .ZN(G402));
endmodule


