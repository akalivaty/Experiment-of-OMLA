

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
         n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706,
         n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717,
         n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
         n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739,
         n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750,
         n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761,
         n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772,
         n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783,
         n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n794,
         n795, n796, n797, n798, n799, n800, n801, n802, n803, n804, n805,
         n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n816,
         n817, n818, n819, n820, n821, n822, n823, n824, n825, n826, n827,
         n828, n829, n830, n831, n832, n833, n834, n835, n836, n837, n838,
         n839, n840, n841, n842, n843, n844, n845, n846, n847, n848, n849,
         n850, n851, n852, n853, n854, n855, n856, n857, n858, n859, n860,
         n861, n862, n863, n864, n865, n866, n867, n868, n869, n870, n871,
         n872, n873, n874, n875, n876, n877, n878, n879, n880, n881, n882,
         n883, n884, n885, n886, n887, n888, n889, n890, n891, n892, n893,
         n894, n895, n896, n897, n898, n899, n900, n901, n902, n903, n904,
         n905, n906, n907, n908, n909, n910, n911, n912, n913, n914, n915,
         n916, n917, n918, n919, n920, n921, n922, n923, n924, n925, n926,
         n927, n928, n929, n930, n931, n932, n933, n934, n935, n936, n937,
         n938, n939, n940, n941, n942, n943, n944, n945, n946, n947, n948,
         n949, n950, n951, n952, n953, n954, n955, n956, n957, n958, n959,
         n960, n961, n962, n963, n964, n965, n966, n967, n968, n969, n970,
         n971, n972, n973, n974, n975, n976, n977, n978, n979, n980, n981,
         n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, n992,
         n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003,
         n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013,
         n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023,
         n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033,
         n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  AND2_X1 U561 ( .A1(n537), .A2(G2105), .ZN(n901) );
  AND2_X1 U562 ( .A1(n776), .A2(n531), .ZN(n777) );
  NAND2_X1 U563 ( .A1(n659), .A2(n658), .ZN(n692) );
  XNOR2_X1 U564 ( .A(n695), .B(n694), .ZN(n697) );
  XNOR2_X1 U565 ( .A(n693), .B(KEYINPUT97), .ZN(n694) );
  NOR2_X1 U566 ( .A1(n985), .A2(n674), .ZN(n689) );
  INV_X1 U567 ( .A(n692), .ZN(n706) );
  XNOR2_X1 U568 ( .A(n704), .B(n703), .ZN(n711) );
  NOR2_X1 U569 ( .A1(G2084), .A2(n726), .ZN(n734) );
  AND2_X1 U570 ( .A1(n732), .A2(n731), .ZN(n733) );
  XOR2_X1 U571 ( .A(n701), .B(KEYINPUT28), .Z(n527) );
  OR2_X1 U572 ( .A1(G1971), .A2(G303), .ZN(n528) );
  NAND2_X1 U573 ( .A1(G29), .A2(n983), .ZN(n529) );
  AND2_X1 U574 ( .A1(n774), .A2(n987), .ZN(n530) );
  NOR2_X1 U575 ( .A1(n775), .A2(n530), .ZN(n531) );
  XOR2_X1 U576 ( .A(KEYINPUT30), .B(n716), .Z(n532) );
  NOR2_X1 U577 ( .A1(n692), .A2(n669), .ZN(n670) );
  XNOR2_X1 U578 ( .A(KEYINPUT26), .B(n670), .ZN(n671) );
  INV_X1 U579 ( .A(KEYINPUT27), .ZN(n693) );
  INV_X1 U580 ( .A(G8), .ZN(n714) );
  NOR2_X1 U581 ( .A1(n734), .A2(n714), .ZN(n715) );
  AND2_X1 U582 ( .A1(n735), .A2(n715), .ZN(n716) );
  INV_X1 U583 ( .A(KEYINPUT29), .ZN(n703) );
  INV_X1 U584 ( .A(KEYINPUT31), .ZN(n721) );
  INV_X1 U585 ( .A(KEYINPUT94), .ZN(n712) );
  INV_X1 U586 ( .A(KEYINPUT105), .ZN(n765) );
  NOR2_X1 U587 ( .A1(G2105), .A2(G2104), .ZN(n533) );
  NOR2_X1 U588 ( .A1(n537), .A2(G2105), .ZN(n617) );
  INV_X1 U589 ( .A(n534), .ZN(n896) );
  NOR2_X1 U590 ( .A1(G651), .A2(G543), .ZN(n806) );
  INV_X1 U591 ( .A(KEYINPUT64), .ZN(n552) );
  XNOR2_X1 U592 ( .A(n553), .B(n552), .ZN(n616) );
  XOR2_X1 U593 ( .A(KEYINPUT17), .B(n533), .Z(n543) );
  INV_X1 U594 ( .A(n543), .ZN(n534) );
  NAND2_X1 U595 ( .A1(G138), .A2(n896), .ZN(n536) );
  XNOR2_X1 U596 ( .A(KEYINPUT65), .B(G2104), .ZN(n537) );
  NAND2_X1 U597 ( .A1(G126), .A2(n901), .ZN(n535) );
  NAND2_X1 U598 ( .A1(n536), .A2(n535), .ZN(n542) );
  NAND2_X1 U599 ( .A1(G102), .A2(n617), .ZN(n538) );
  XNOR2_X1 U600 ( .A(n538), .B(KEYINPUT88), .ZN(n540) );
  AND2_X1 U601 ( .A1(G2105), .A2(G2104), .ZN(n900) );
  NAND2_X1 U602 ( .A1(n900), .A2(G114), .ZN(n539) );
  NAND2_X1 U603 ( .A1(n540), .A2(n539), .ZN(n541) );
  NOR2_X1 U604 ( .A1(n542), .A2(n541), .ZN(G164) );
  NAND2_X1 U605 ( .A1(G137), .A2(n543), .ZN(n544) );
  XNOR2_X1 U606 ( .A(n544), .B(KEYINPUT66), .ZN(n551) );
  NAND2_X1 U607 ( .A1(G113), .A2(n900), .ZN(n546) );
  NAND2_X1 U608 ( .A1(G125), .A2(n901), .ZN(n545) );
  NAND2_X1 U609 ( .A1(n546), .A2(n545), .ZN(n549) );
  NAND2_X1 U610 ( .A1(n617), .A2(G101), .ZN(n547) );
  XNOR2_X1 U611 ( .A(n547), .B(KEYINPUT23), .ZN(n548) );
  NOR2_X1 U612 ( .A1(n549), .A2(n548), .ZN(n550) );
  NAND2_X1 U613 ( .A1(n551), .A2(n550), .ZN(n553) );
  BUF_X1 U614 ( .A(n616), .Z(G160) );
  XOR2_X1 U615 ( .A(G543), .B(KEYINPUT0), .Z(n610) );
  NOR2_X2 U616 ( .A1(G651), .A2(n610), .ZN(n808) );
  NAND2_X1 U617 ( .A1(G52), .A2(n808), .ZN(n556) );
  INV_X1 U618 ( .A(G651), .ZN(n558) );
  NOR2_X1 U619 ( .A1(G543), .A2(n558), .ZN(n554) );
  XOR2_X1 U620 ( .A(KEYINPUT1), .B(n554), .Z(n812) );
  NAND2_X1 U621 ( .A1(G64), .A2(n812), .ZN(n555) );
  NAND2_X1 U622 ( .A1(n556), .A2(n555), .ZN(n563) );
  NAND2_X1 U623 ( .A1(n806), .A2(G90), .ZN(n557) );
  XOR2_X1 U624 ( .A(KEYINPUT69), .B(n557), .Z(n560) );
  NOR2_X1 U625 ( .A1(n610), .A2(n558), .ZN(n809) );
  NAND2_X1 U626 ( .A1(n809), .A2(G77), .ZN(n559) );
  NAND2_X1 U627 ( .A1(n560), .A2(n559), .ZN(n561) );
  XOR2_X1 U628 ( .A(KEYINPUT9), .B(n561), .Z(n562) );
  NOR2_X1 U629 ( .A1(n563), .A2(n562), .ZN(G171) );
  AND2_X1 U630 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U631 ( .A(G57), .ZN(G237) );
  INV_X1 U632 ( .A(G132), .ZN(G219) );
  INV_X1 U633 ( .A(G82), .ZN(G220) );
  NAND2_X1 U634 ( .A1(G75), .A2(n809), .ZN(n565) );
  NAND2_X1 U635 ( .A1(G88), .A2(n806), .ZN(n564) );
  NAND2_X1 U636 ( .A1(n565), .A2(n564), .ZN(n569) );
  NAND2_X1 U637 ( .A1(G50), .A2(n808), .ZN(n567) );
  NAND2_X1 U638 ( .A1(G62), .A2(n812), .ZN(n566) );
  NAND2_X1 U639 ( .A1(n567), .A2(n566), .ZN(n568) );
  NOR2_X1 U640 ( .A1(n569), .A2(n568), .ZN(G166) );
  NAND2_X1 U641 ( .A1(n808), .A2(G51), .ZN(n570) );
  XOR2_X1 U642 ( .A(KEYINPUT75), .B(n570), .Z(n572) );
  NAND2_X1 U643 ( .A1(n812), .A2(G63), .ZN(n571) );
  NAND2_X1 U644 ( .A1(n572), .A2(n571), .ZN(n573) );
  XNOR2_X1 U645 ( .A(KEYINPUT6), .B(n573), .ZN(n580) );
  NAND2_X1 U646 ( .A1(G89), .A2(n806), .ZN(n574) );
  XNOR2_X1 U647 ( .A(n574), .B(KEYINPUT74), .ZN(n575) );
  XNOR2_X1 U648 ( .A(n575), .B(KEYINPUT4), .ZN(n577) );
  NAND2_X1 U649 ( .A1(G76), .A2(n809), .ZN(n576) );
  NAND2_X1 U650 ( .A1(n577), .A2(n576), .ZN(n578) );
  XOR2_X1 U651 ( .A(n578), .B(KEYINPUT5), .Z(n579) );
  NOR2_X1 U652 ( .A1(n580), .A2(n579), .ZN(n581) );
  XOR2_X1 U653 ( .A(KEYINPUT76), .B(n581), .Z(n582) );
  XNOR2_X1 U654 ( .A(KEYINPUT7), .B(n582), .ZN(G168) );
  XNOR2_X1 U655 ( .A(KEYINPUT77), .B(KEYINPUT8), .ZN(n583) );
  XNOR2_X1 U656 ( .A(n583), .B(G168), .ZN(G286) );
  NAND2_X1 U657 ( .A1(G47), .A2(n808), .ZN(n584) );
  XNOR2_X1 U658 ( .A(n584), .B(KEYINPUT68), .ZN(n586) );
  NAND2_X1 U659 ( .A1(n812), .A2(G60), .ZN(n585) );
  NAND2_X1 U660 ( .A1(n586), .A2(n585), .ZN(n589) );
  NAND2_X1 U661 ( .A1(G72), .A2(n809), .ZN(n587) );
  XNOR2_X1 U662 ( .A(KEYINPUT67), .B(n587), .ZN(n588) );
  NOR2_X1 U663 ( .A1(n589), .A2(n588), .ZN(n591) );
  NAND2_X1 U664 ( .A1(n806), .A2(G85), .ZN(n590) );
  NAND2_X1 U665 ( .A1(n591), .A2(n590), .ZN(G290) );
  NAND2_X1 U666 ( .A1(G78), .A2(n809), .ZN(n593) );
  NAND2_X1 U667 ( .A1(G91), .A2(n806), .ZN(n592) );
  NAND2_X1 U668 ( .A1(n593), .A2(n592), .ZN(n594) );
  XOR2_X1 U669 ( .A(KEYINPUT70), .B(n594), .Z(n600) );
  NAND2_X1 U670 ( .A1(n812), .A2(G65), .ZN(n595) );
  XOR2_X1 U671 ( .A(KEYINPUT71), .B(n595), .Z(n597) );
  NAND2_X1 U672 ( .A1(n808), .A2(G53), .ZN(n596) );
  NAND2_X1 U673 ( .A1(n597), .A2(n596), .ZN(n598) );
  XOR2_X1 U674 ( .A(KEYINPUT72), .B(n598), .Z(n599) );
  NAND2_X1 U675 ( .A1(n600), .A2(n599), .ZN(G299) );
  INV_X1 U676 ( .A(G166), .ZN(G303) );
  NAND2_X1 U677 ( .A1(G61), .A2(n812), .ZN(n602) );
  NAND2_X1 U678 ( .A1(G86), .A2(n806), .ZN(n601) );
  NAND2_X1 U679 ( .A1(n602), .A2(n601), .ZN(n605) );
  NAND2_X1 U680 ( .A1(n809), .A2(G73), .ZN(n603) );
  XOR2_X1 U681 ( .A(KEYINPUT2), .B(n603), .Z(n604) );
  NOR2_X1 U682 ( .A1(n605), .A2(n604), .ZN(n606) );
  XOR2_X1 U683 ( .A(KEYINPUT83), .B(n606), .Z(n608) );
  NAND2_X1 U684 ( .A1(n808), .A2(G48), .ZN(n607) );
  NAND2_X1 U685 ( .A1(n608), .A2(n607), .ZN(G305) );
  NAND2_X1 U686 ( .A1(G74), .A2(G651), .ZN(n609) );
  XNOR2_X1 U687 ( .A(n609), .B(KEYINPUT82), .ZN(n615) );
  NAND2_X1 U688 ( .A1(G49), .A2(n808), .ZN(n612) );
  NAND2_X1 U689 ( .A1(G87), .A2(n610), .ZN(n611) );
  NAND2_X1 U690 ( .A1(n612), .A2(n611), .ZN(n613) );
  NOR2_X1 U691 ( .A1(n812), .A2(n613), .ZN(n614) );
  NAND2_X1 U692 ( .A1(n615), .A2(n614), .ZN(G288) );
  INV_X1 U693 ( .A(KEYINPUT40), .ZN(n781) );
  NOR2_X1 U694 ( .A1(G164), .A2(G1384), .ZN(n658) );
  NAND2_X1 U695 ( .A1(n616), .A2(G40), .ZN(n657) );
  NOR2_X1 U696 ( .A1(n658), .A2(n657), .ZN(n774) );
  XOR2_X1 U697 ( .A(KEYINPUT92), .B(KEYINPUT38), .Z(n619) );
  BUF_X1 U698 ( .A(n617), .Z(n897) );
  NAND2_X1 U699 ( .A1(G105), .A2(n897), .ZN(n618) );
  XNOR2_X1 U700 ( .A(n619), .B(n618), .ZN(n623) );
  NAND2_X1 U701 ( .A1(G141), .A2(n896), .ZN(n621) );
  NAND2_X1 U702 ( .A1(G117), .A2(n900), .ZN(n620) );
  NAND2_X1 U703 ( .A1(n621), .A2(n620), .ZN(n622) );
  NOR2_X1 U704 ( .A1(n623), .A2(n622), .ZN(n625) );
  NAND2_X1 U705 ( .A1(n901), .A2(G129), .ZN(n624) );
  NAND2_X1 U706 ( .A1(n625), .A2(n624), .ZN(n891) );
  NOR2_X1 U707 ( .A1(G1996), .A2(n891), .ZN(n959) );
  NAND2_X1 U708 ( .A1(G107), .A2(n900), .ZN(n627) );
  NAND2_X1 U709 ( .A1(G119), .A2(n901), .ZN(n626) );
  NAND2_X1 U710 ( .A1(n627), .A2(n626), .ZN(n632) );
  NAND2_X1 U711 ( .A1(G131), .A2(n896), .ZN(n629) );
  NAND2_X1 U712 ( .A1(G95), .A2(n897), .ZN(n628) );
  NAND2_X1 U713 ( .A1(n629), .A2(n628), .ZN(n630) );
  XOR2_X1 U714 ( .A(KEYINPUT91), .B(n630), .Z(n631) );
  NOR2_X1 U715 ( .A1(n632), .A2(n631), .ZN(n886) );
  INV_X1 U716 ( .A(G1991), .ZN(n636) );
  NOR2_X1 U717 ( .A1(n886), .A2(n636), .ZN(n634) );
  AND2_X1 U718 ( .A1(n891), .A2(G1996), .ZN(n633) );
  NOR2_X1 U719 ( .A1(n634), .A2(n633), .ZN(n974) );
  INV_X1 U720 ( .A(n774), .ZN(n635) );
  NOR2_X1 U721 ( .A1(n974), .A2(n635), .ZN(n770) );
  NOR2_X1 U722 ( .A1(G1986), .A2(G290), .ZN(n637) );
  AND2_X1 U723 ( .A1(n636), .A2(n886), .ZN(n963) );
  NOR2_X1 U724 ( .A1(n637), .A2(n963), .ZN(n638) );
  NOR2_X1 U725 ( .A1(n770), .A2(n638), .ZN(n639) );
  NOR2_X1 U726 ( .A1(n959), .A2(n639), .ZN(n640) );
  XNOR2_X1 U727 ( .A(n640), .B(KEYINPUT39), .ZN(n652) );
  NAND2_X1 U728 ( .A1(G140), .A2(n896), .ZN(n642) );
  NAND2_X1 U729 ( .A1(G104), .A2(n897), .ZN(n641) );
  NAND2_X1 U730 ( .A1(n642), .A2(n641), .ZN(n644) );
  XOR2_X1 U731 ( .A(KEYINPUT34), .B(KEYINPUT89), .Z(n643) );
  XNOR2_X1 U732 ( .A(n644), .B(n643), .ZN(n650) );
  NAND2_X1 U733 ( .A1(n901), .A2(G128), .ZN(n645) );
  XNOR2_X1 U734 ( .A(n645), .B(KEYINPUT90), .ZN(n647) );
  NAND2_X1 U735 ( .A1(G116), .A2(n900), .ZN(n646) );
  NAND2_X1 U736 ( .A1(n647), .A2(n646), .ZN(n648) );
  XOR2_X1 U737 ( .A(KEYINPUT35), .B(n648), .Z(n649) );
  NOR2_X1 U738 ( .A1(n650), .A2(n649), .ZN(n651) );
  XNOR2_X1 U739 ( .A(KEYINPUT36), .B(n651), .ZN(n892) );
  XNOR2_X1 U740 ( .A(G2067), .B(KEYINPUT37), .ZN(n653) );
  NOR2_X1 U741 ( .A1(n892), .A2(n653), .ZN(n980) );
  NAND2_X1 U742 ( .A1(n774), .A2(n980), .ZN(n772) );
  NAND2_X1 U743 ( .A1(n652), .A2(n772), .ZN(n654) );
  NAND2_X1 U744 ( .A1(n892), .A2(n653), .ZN(n973) );
  NAND2_X1 U745 ( .A1(n654), .A2(n973), .ZN(n655) );
  NAND2_X1 U746 ( .A1(n774), .A2(n655), .ZN(n656) );
  XNOR2_X1 U747 ( .A(KEYINPUT109), .B(n656), .ZN(n779) );
  INV_X1 U748 ( .A(n657), .ZN(n659) );
  NAND2_X1 U749 ( .A1(G8), .A2(n692), .ZN(n758) );
  NAND2_X1 U750 ( .A1(G56), .A2(n812), .ZN(n660) );
  XOR2_X1 U751 ( .A(KEYINPUT14), .B(n660), .Z(n666) );
  NAND2_X1 U752 ( .A1(n806), .A2(G81), .ZN(n661) );
  XNOR2_X1 U753 ( .A(n661), .B(KEYINPUT12), .ZN(n663) );
  NAND2_X1 U754 ( .A1(G68), .A2(n809), .ZN(n662) );
  NAND2_X1 U755 ( .A1(n663), .A2(n662), .ZN(n664) );
  XOR2_X1 U756 ( .A(KEYINPUT13), .B(n664), .Z(n665) );
  NOR2_X1 U757 ( .A1(n666), .A2(n665), .ZN(n668) );
  NAND2_X1 U758 ( .A1(n808), .A2(G43), .ZN(n667) );
  NAND2_X1 U759 ( .A1(n668), .A2(n667), .ZN(n985) );
  INV_X1 U760 ( .A(G1996), .ZN(n669) );
  INV_X1 U761 ( .A(n671), .ZN(n673) );
  BUF_X2 U762 ( .A(n692), .Z(n726) );
  NAND2_X1 U763 ( .A1(n726), .A2(G1341), .ZN(n672) );
  NAND2_X1 U764 ( .A1(n673), .A2(n672), .ZN(n674) );
  NAND2_X1 U765 ( .A1(G66), .A2(n812), .ZN(n676) );
  NAND2_X1 U766 ( .A1(G92), .A2(n806), .ZN(n675) );
  NAND2_X1 U767 ( .A1(n676), .A2(n675), .ZN(n681) );
  NAND2_X1 U768 ( .A1(G54), .A2(n808), .ZN(n678) );
  NAND2_X1 U769 ( .A1(G79), .A2(n809), .ZN(n677) );
  NAND2_X1 U770 ( .A1(n678), .A2(n677), .ZN(n679) );
  XOR2_X1 U771 ( .A(KEYINPUT73), .B(n679), .Z(n680) );
  NOR2_X1 U772 ( .A1(n681), .A2(n680), .ZN(n682) );
  XOR2_X1 U773 ( .A(KEYINPUT15), .B(n682), .Z(n913) );
  NAND2_X1 U774 ( .A1(n689), .A2(n913), .ZN(n687) );
  INV_X1 U775 ( .A(G2067), .ZN(n938) );
  NOR2_X1 U776 ( .A1(n726), .A2(n938), .ZN(n683) );
  XNOR2_X1 U777 ( .A(n683), .B(KEYINPUT99), .ZN(n685) );
  NAND2_X1 U778 ( .A1(n726), .A2(G1348), .ZN(n684) );
  NAND2_X1 U779 ( .A1(n685), .A2(n684), .ZN(n686) );
  NAND2_X1 U780 ( .A1(n687), .A2(n686), .ZN(n688) );
  XNOR2_X1 U781 ( .A(n688), .B(KEYINPUT100), .ZN(n691) );
  OR2_X1 U782 ( .A1(n689), .A2(n913), .ZN(n690) );
  NAND2_X1 U783 ( .A1(n691), .A2(n690), .ZN(n699) );
  INV_X1 U784 ( .A(G299), .ZN(n819) );
  NAND2_X1 U785 ( .A1(G2072), .A2(n706), .ZN(n695) );
  XOR2_X1 U786 ( .A(G1956), .B(KEYINPUT98), .Z(n1012) );
  NOR2_X1 U787 ( .A1(n706), .A2(n1012), .ZN(n696) );
  NOR2_X1 U788 ( .A1(n697), .A2(n696), .ZN(n700) );
  NAND2_X1 U789 ( .A1(n819), .A2(n700), .ZN(n698) );
  NAND2_X1 U790 ( .A1(n699), .A2(n698), .ZN(n702) );
  NOR2_X1 U791 ( .A1(n819), .A2(n700), .ZN(n701) );
  NAND2_X1 U792 ( .A1(n702), .A2(n527), .ZN(n704) );
  XOR2_X1 U793 ( .A(KEYINPUT25), .B(G2078), .Z(n942) );
  NOR2_X1 U794 ( .A1(n942), .A2(n726), .ZN(n705) );
  XOR2_X1 U795 ( .A(KEYINPUT96), .B(n705), .Z(n709) );
  NOR2_X1 U796 ( .A1(n706), .A2(G1961), .ZN(n707) );
  XNOR2_X1 U797 ( .A(KEYINPUT95), .B(n707), .ZN(n708) );
  NAND2_X1 U798 ( .A1(n709), .A2(n708), .ZN(n717) );
  NAND2_X1 U799 ( .A1(n717), .A2(G171), .ZN(n710) );
  NAND2_X1 U800 ( .A1(n711), .A2(n710), .ZN(n724) );
  NOR2_X1 U801 ( .A1(G1966), .A2(n758), .ZN(n713) );
  XNOR2_X1 U802 ( .A(n713), .B(n712), .ZN(n735) );
  NOR2_X1 U803 ( .A1(G168), .A2(n532), .ZN(n720) );
  NOR2_X1 U804 ( .A1(G171), .A2(n717), .ZN(n718) );
  XOR2_X1 U805 ( .A(KEYINPUT101), .B(n718), .Z(n719) );
  NOR2_X1 U806 ( .A1(n720), .A2(n719), .ZN(n722) );
  XNOR2_X1 U807 ( .A(n722), .B(n721), .ZN(n723) );
  NAND2_X1 U808 ( .A1(n724), .A2(n723), .ZN(n736) );
  AND2_X1 U809 ( .A1(G286), .A2(G8), .ZN(n725) );
  NAND2_X1 U810 ( .A1(n736), .A2(n725), .ZN(n732) );
  NOR2_X1 U811 ( .A1(G1971), .A2(n758), .ZN(n728) );
  NOR2_X1 U812 ( .A1(G2090), .A2(n726), .ZN(n727) );
  NOR2_X1 U813 ( .A1(n728), .A2(n727), .ZN(n729) );
  NAND2_X1 U814 ( .A1(n729), .A2(G303), .ZN(n730) );
  OR2_X1 U815 ( .A1(n714), .A2(n730), .ZN(n731) );
  XNOR2_X1 U816 ( .A(n733), .B(KEYINPUT32), .ZN(n740) );
  NAND2_X1 U817 ( .A1(G8), .A2(n734), .ZN(n738) );
  AND2_X1 U818 ( .A1(n736), .A2(n735), .ZN(n737) );
  NAND2_X1 U819 ( .A1(n738), .A2(n737), .ZN(n739) );
  NAND2_X1 U820 ( .A1(n740), .A2(n739), .ZN(n749) );
  NOR2_X1 U821 ( .A1(G2090), .A2(G303), .ZN(n741) );
  NAND2_X1 U822 ( .A1(G8), .A2(n741), .ZN(n742) );
  NAND2_X1 U823 ( .A1(n749), .A2(n742), .ZN(n743) );
  NAND2_X1 U824 ( .A1(n758), .A2(n743), .ZN(n744) );
  XNOR2_X1 U825 ( .A(n744), .B(KEYINPUT106), .ZN(n748) );
  INV_X1 U826 ( .A(n758), .ZN(n755) );
  NOR2_X1 U827 ( .A1(G1981), .A2(G305), .ZN(n745) );
  XNOR2_X1 U828 ( .A(n745), .B(KEYINPUT24), .ZN(n746) );
  NAND2_X1 U829 ( .A1(n755), .A2(n746), .ZN(n747) );
  NAND2_X1 U830 ( .A1(n748), .A2(n747), .ZN(n768) );
  AND2_X1 U831 ( .A1(n749), .A2(n528), .ZN(n753) );
  NOR2_X1 U832 ( .A1(G1976), .A2(G288), .ZN(n750) );
  XOR2_X1 U833 ( .A(KEYINPUT102), .B(n750), .Z(n997) );
  INV_X1 U834 ( .A(KEYINPUT33), .ZN(n751) );
  AND2_X1 U835 ( .A1(n997), .A2(n751), .ZN(n752) );
  AND2_X1 U836 ( .A1(n753), .A2(n752), .ZN(n764) );
  NAND2_X1 U837 ( .A1(G288), .A2(G1976), .ZN(n754) );
  XOR2_X1 U838 ( .A(KEYINPUT103), .B(n754), .Z(n993) );
  AND2_X1 U839 ( .A1(n755), .A2(n993), .ZN(n756) );
  OR2_X1 U840 ( .A1(KEYINPUT33), .A2(n756), .ZN(n762) );
  XOR2_X1 U841 ( .A(KEYINPUT104), .B(G1981), .Z(n757) );
  XNOR2_X1 U842 ( .A(G305), .B(n757), .ZN(n1000) );
  NOR2_X1 U843 ( .A1(n997), .A2(n758), .ZN(n759) );
  NAND2_X1 U844 ( .A1(KEYINPUT33), .A2(n759), .ZN(n760) );
  AND2_X1 U845 ( .A1(n1000), .A2(n760), .ZN(n761) );
  NAND2_X1 U846 ( .A1(n762), .A2(n761), .ZN(n763) );
  NOR2_X2 U847 ( .A1(n764), .A2(n763), .ZN(n766) );
  XNOR2_X1 U848 ( .A(n766), .B(n765), .ZN(n767) );
  NOR2_X1 U849 ( .A1(n768), .A2(n767), .ZN(n769) );
  XNOR2_X1 U850 ( .A(n769), .B(KEYINPUT107), .ZN(n776) );
  INV_X1 U851 ( .A(n770), .ZN(n771) );
  NAND2_X1 U852 ( .A1(n772), .A2(n771), .ZN(n773) );
  XOR2_X1 U853 ( .A(KEYINPUT93), .B(n773), .Z(n775) );
  XNOR2_X1 U854 ( .A(G1986), .B(G290), .ZN(n987) );
  XNOR2_X1 U855 ( .A(n777), .B(KEYINPUT108), .ZN(n778) );
  NOR2_X1 U856 ( .A1(n779), .A2(n778), .ZN(n780) );
  XNOR2_X1 U857 ( .A(n781), .B(n780), .ZN(G329) );
  NAND2_X1 U858 ( .A1(G7), .A2(G661), .ZN(n782) );
  XNOR2_X1 U859 ( .A(n782), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U860 ( .A(G223), .ZN(n847) );
  NAND2_X1 U861 ( .A1(n847), .A2(G567), .ZN(n783) );
  XOR2_X1 U862 ( .A(KEYINPUT11), .B(n783), .Z(G234) );
  INV_X1 U863 ( .A(G860), .ZN(n805) );
  OR2_X1 U864 ( .A1(n985), .A2(n805), .ZN(G153) );
  INV_X1 U865 ( .A(G171), .ZN(G301) );
  NAND2_X1 U866 ( .A1(G868), .A2(G301), .ZN(n785) );
  INV_X1 U867 ( .A(n913), .ZN(n990) );
  INV_X1 U868 ( .A(G868), .ZN(n828) );
  NAND2_X1 U869 ( .A1(n990), .A2(n828), .ZN(n784) );
  NAND2_X1 U870 ( .A1(n785), .A2(n784), .ZN(G284) );
  NAND2_X1 U871 ( .A1(G868), .A2(G286), .ZN(n787) );
  NAND2_X1 U872 ( .A1(G299), .A2(n828), .ZN(n786) );
  NAND2_X1 U873 ( .A1(n787), .A2(n786), .ZN(G297) );
  NAND2_X1 U874 ( .A1(n805), .A2(G559), .ZN(n788) );
  NAND2_X1 U875 ( .A1(n788), .A2(n913), .ZN(n789) );
  XNOR2_X1 U876 ( .A(n789), .B(KEYINPUT16), .ZN(G148) );
  NAND2_X1 U877 ( .A1(n913), .A2(G868), .ZN(n790) );
  NOR2_X1 U878 ( .A1(G559), .A2(n790), .ZN(n791) );
  XNOR2_X1 U879 ( .A(n791), .B(KEYINPUT78), .ZN(n793) );
  NOR2_X1 U880 ( .A1(n985), .A2(G868), .ZN(n792) );
  NOR2_X1 U881 ( .A1(n793), .A2(n792), .ZN(G282) );
  NAND2_X1 U882 ( .A1(G135), .A2(n896), .ZN(n795) );
  NAND2_X1 U883 ( .A1(G111), .A2(n900), .ZN(n794) );
  NAND2_X1 U884 ( .A1(n795), .A2(n794), .ZN(n800) );
  NAND2_X1 U885 ( .A1(n901), .A2(G123), .ZN(n796) );
  XNOR2_X1 U886 ( .A(n796), .B(KEYINPUT18), .ZN(n798) );
  NAND2_X1 U887 ( .A1(G99), .A2(n897), .ZN(n797) );
  NAND2_X1 U888 ( .A1(n798), .A2(n797), .ZN(n799) );
  NOR2_X1 U889 ( .A1(n800), .A2(n799), .ZN(n962) );
  XNOR2_X1 U890 ( .A(G2096), .B(n962), .ZN(n802) );
  INV_X1 U891 ( .A(G2100), .ZN(n801) );
  NAND2_X1 U892 ( .A1(n802), .A2(n801), .ZN(G156) );
  XNOR2_X1 U893 ( .A(n985), .B(KEYINPUT79), .ZN(n804) );
  NAND2_X1 U894 ( .A1(n913), .A2(G559), .ZN(n803) );
  XNOR2_X1 U895 ( .A(n804), .B(n803), .ZN(n826) );
  NAND2_X1 U896 ( .A1(n805), .A2(n826), .ZN(n818) );
  NAND2_X1 U897 ( .A1(G93), .A2(n806), .ZN(n807) );
  XNOR2_X1 U898 ( .A(n807), .B(KEYINPUT80), .ZN(n817) );
  NAND2_X1 U899 ( .A1(G55), .A2(n808), .ZN(n811) );
  NAND2_X1 U900 ( .A1(G80), .A2(n809), .ZN(n810) );
  NAND2_X1 U901 ( .A1(n811), .A2(n810), .ZN(n815) );
  NAND2_X1 U902 ( .A1(G67), .A2(n812), .ZN(n813) );
  XNOR2_X1 U903 ( .A(KEYINPUT81), .B(n813), .ZN(n814) );
  NOR2_X1 U904 ( .A1(n815), .A2(n814), .ZN(n816) );
  NAND2_X1 U905 ( .A1(n817), .A2(n816), .ZN(n829) );
  XNOR2_X1 U906 ( .A(n818), .B(n829), .ZN(G145) );
  XNOR2_X1 U907 ( .A(n819), .B(G305), .ZN(n825) );
  XNOR2_X1 U908 ( .A(KEYINPUT19), .B(KEYINPUT84), .ZN(n821) );
  XNOR2_X1 U909 ( .A(G290), .B(G166), .ZN(n820) );
  XNOR2_X1 U910 ( .A(n821), .B(n820), .ZN(n822) );
  XOR2_X1 U911 ( .A(n822), .B(G288), .Z(n823) );
  XNOR2_X1 U912 ( .A(n829), .B(n823), .ZN(n824) );
  XNOR2_X1 U913 ( .A(n825), .B(n824), .ZN(n912) );
  XOR2_X1 U914 ( .A(n912), .B(n826), .Z(n827) );
  NOR2_X1 U915 ( .A1(n828), .A2(n827), .ZN(n831) );
  NOR2_X1 U916 ( .A1(G868), .A2(n829), .ZN(n830) );
  NOR2_X1 U917 ( .A1(n831), .A2(n830), .ZN(n832) );
  XOR2_X1 U918 ( .A(KEYINPUT85), .B(n832), .Z(G295) );
  NAND2_X1 U919 ( .A1(G2078), .A2(G2084), .ZN(n834) );
  XOR2_X1 U920 ( .A(KEYINPUT86), .B(KEYINPUT20), .Z(n833) );
  XNOR2_X1 U921 ( .A(n834), .B(n833), .ZN(n835) );
  NAND2_X1 U922 ( .A1(G2090), .A2(n835), .ZN(n836) );
  XNOR2_X1 U923 ( .A(KEYINPUT21), .B(n836), .ZN(n837) );
  NAND2_X1 U924 ( .A1(n837), .A2(G2072), .ZN(n838) );
  XOR2_X1 U925 ( .A(KEYINPUT87), .B(n838), .Z(G158) );
  XNOR2_X1 U926 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U927 ( .A1(G220), .A2(G219), .ZN(n839) );
  XOR2_X1 U928 ( .A(KEYINPUT22), .B(n839), .Z(n840) );
  NOR2_X1 U929 ( .A1(G218), .A2(n840), .ZN(n841) );
  NAND2_X1 U930 ( .A1(G96), .A2(n841), .ZN(n934) );
  NAND2_X1 U931 ( .A1(n934), .A2(G2106), .ZN(n845) );
  NAND2_X1 U932 ( .A1(G69), .A2(G120), .ZN(n842) );
  NOR2_X1 U933 ( .A1(G237), .A2(n842), .ZN(n843) );
  NAND2_X1 U934 ( .A1(G108), .A2(n843), .ZN(n935) );
  NAND2_X1 U935 ( .A1(n935), .A2(G567), .ZN(n844) );
  NAND2_X1 U936 ( .A1(n845), .A2(n844), .ZN(n853) );
  NAND2_X1 U937 ( .A1(G483), .A2(G661), .ZN(n846) );
  NOR2_X1 U938 ( .A1(n853), .A2(n846), .ZN(n852) );
  NAND2_X1 U939 ( .A1(n852), .A2(G36), .ZN(G176) );
  NAND2_X1 U940 ( .A1(n847), .A2(G2106), .ZN(n848) );
  XNOR2_X1 U941 ( .A(n848), .B(KEYINPUT110), .ZN(G217) );
  AND2_X1 U942 ( .A1(G15), .A2(G2), .ZN(n849) );
  NAND2_X1 U943 ( .A1(G661), .A2(n849), .ZN(G259) );
  NAND2_X1 U944 ( .A1(G3), .A2(G1), .ZN(n850) );
  XOR2_X1 U945 ( .A(KEYINPUT111), .B(n850), .Z(n851) );
  NAND2_X1 U946 ( .A1(n852), .A2(n851), .ZN(G188) );
  INV_X1 U947 ( .A(n853), .ZN(G319) );
  XOR2_X1 U948 ( .A(G2096), .B(KEYINPUT43), .Z(n855) );
  XNOR2_X1 U949 ( .A(G2090), .B(G2678), .ZN(n854) );
  XNOR2_X1 U950 ( .A(n855), .B(n854), .ZN(n856) );
  XOR2_X1 U951 ( .A(n856), .B(KEYINPUT112), .Z(n858) );
  XNOR2_X1 U952 ( .A(G2067), .B(G2072), .ZN(n857) );
  XNOR2_X1 U953 ( .A(n858), .B(n857), .ZN(n862) );
  XOR2_X1 U954 ( .A(KEYINPUT42), .B(G2100), .Z(n860) );
  XNOR2_X1 U955 ( .A(G2078), .B(G2084), .ZN(n859) );
  XNOR2_X1 U956 ( .A(n860), .B(n859), .ZN(n861) );
  XNOR2_X1 U957 ( .A(n862), .B(n861), .ZN(G227) );
  XOR2_X1 U958 ( .A(G1966), .B(G1971), .Z(n864) );
  XNOR2_X1 U959 ( .A(G1981), .B(G1976), .ZN(n863) );
  XNOR2_X1 U960 ( .A(n864), .B(n863), .ZN(n865) );
  XOR2_X1 U961 ( .A(n865), .B(G2474), .Z(n867) );
  XNOR2_X1 U962 ( .A(G1986), .B(G1956), .ZN(n866) );
  XNOR2_X1 U963 ( .A(n867), .B(n866), .ZN(n871) );
  XOR2_X1 U964 ( .A(KEYINPUT41), .B(G1961), .Z(n869) );
  XNOR2_X1 U965 ( .A(G1996), .B(G1991), .ZN(n868) );
  XNOR2_X1 U966 ( .A(n869), .B(n868), .ZN(n870) );
  XNOR2_X1 U967 ( .A(n871), .B(n870), .ZN(G229) );
  NAND2_X1 U968 ( .A1(G136), .A2(n896), .ZN(n873) );
  NAND2_X1 U969 ( .A1(G112), .A2(n900), .ZN(n872) );
  NAND2_X1 U970 ( .A1(n873), .A2(n872), .ZN(n878) );
  NAND2_X1 U971 ( .A1(n901), .A2(G124), .ZN(n874) );
  XNOR2_X1 U972 ( .A(n874), .B(KEYINPUT44), .ZN(n876) );
  NAND2_X1 U973 ( .A1(G100), .A2(n897), .ZN(n875) );
  NAND2_X1 U974 ( .A1(n876), .A2(n875), .ZN(n877) );
  NOR2_X1 U975 ( .A1(n878), .A2(n877), .ZN(G162) );
  NAND2_X1 U976 ( .A1(G118), .A2(n900), .ZN(n880) );
  NAND2_X1 U977 ( .A1(G130), .A2(n901), .ZN(n879) );
  NAND2_X1 U978 ( .A1(n880), .A2(n879), .ZN(n885) );
  NAND2_X1 U979 ( .A1(G142), .A2(n896), .ZN(n882) );
  NAND2_X1 U980 ( .A1(G106), .A2(n897), .ZN(n881) );
  NAND2_X1 U981 ( .A1(n882), .A2(n881), .ZN(n883) );
  XOR2_X1 U982 ( .A(n883), .B(KEYINPUT45), .Z(n884) );
  NOR2_X1 U983 ( .A1(n885), .A2(n884), .ZN(n887) );
  XOR2_X1 U984 ( .A(n887), .B(n886), .Z(n910) );
  XOR2_X1 U985 ( .A(KEYINPUT48), .B(KEYINPUT46), .Z(n889) );
  XNOR2_X1 U986 ( .A(G164), .B(KEYINPUT113), .ZN(n888) );
  XNOR2_X1 U987 ( .A(n889), .B(n888), .ZN(n890) );
  XNOR2_X1 U988 ( .A(G162), .B(n890), .ZN(n894) );
  XOR2_X1 U989 ( .A(n892), .B(n891), .Z(n893) );
  XNOR2_X1 U990 ( .A(n894), .B(n893), .ZN(n895) );
  XNOR2_X1 U991 ( .A(n962), .B(n895), .ZN(n908) );
  NAND2_X1 U992 ( .A1(G139), .A2(n896), .ZN(n899) );
  NAND2_X1 U993 ( .A1(G103), .A2(n897), .ZN(n898) );
  NAND2_X1 U994 ( .A1(n899), .A2(n898), .ZN(n906) );
  NAND2_X1 U995 ( .A1(G115), .A2(n900), .ZN(n903) );
  NAND2_X1 U996 ( .A1(G127), .A2(n901), .ZN(n902) );
  NAND2_X1 U997 ( .A1(n903), .A2(n902), .ZN(n904) );
  XOR2_X1 U998 ( .A(KEYINPUT47), .B(n904), .Z(n905) );
  NOR2_X1 U999 ( .A1(n906), .A2(n905), .ZN(n967) );
  XNOR2_X1 U1000 ( .A(G160), .B(n967), .ZN(n907) );
  XNOR2_X1 U1001 ( .A(n908), .B(n907), .ZN(n909) );
  XOR2_X1 U1002 ( .A(n910), .B(n909), .Z(n911) );
  NOR2_X1 U1003 ( .A1(G37), .A2(n911), .ZN(G395) );
  XNOR2_X1 U1004 ( .A(n985), .B(n912), .ZN(n915) );
  XNOR2_X1 U1005 ( .A(G171), .B(n913), .ZN(n914) );
  XNOR2_X1 U1006 ( .A(n915), .B(n914), .ZN(n916) );
  XOR2_X1 U1007 ( .A(n916), .B(G286), .Z(n917) );
  NOR2_X1 U1008 ( .A1(G37), .A2(n917), .ZN(n918) );
  XNOR2_X1 U1009 ( .A(KEYINPUT114), .B(n918), .ZN(G397) );
  XOR2_X1 U1010 ( .A(G2451), .B(G2430), .Z(n920) );
  XNOR2_X1 U1011 ( .A(G2438), .B(G2443), .ZN(n919) );
  XNOR2_X1 U1012 ( .A(n920), .B(n919), .ZN(n926) );
  XOR2_X1 U1013 ( .A(G2435), .B(G2454), .Z(n922) );
  XNOR2_X1 U1014 ( .A(G1341), .B(G1348), .ZN(n921) );
  XNOR2_X1 U1015 ( .A(n922), .B(n921), .ZN(n924) );
  XOR2_X1 U1016 ( .A(G2446), .B(G2427), .Z(n923) );
  XNOR2_X1 U1017 ( .A(n924), .B(n923), .ZN(n925) );
  XOR2_X1 U1018 ( .A(n926), .B(n925), .Z(n927) );
  NAND2_X1 U1019 ( .A1(G14), .A2(n927), .ZN(n936) );
  NAND2_X1 U1020 ( .A1(G319), .A2(n936), .ZN(n931) );
  NOR2_X1 U1021 ( .A1(G227), .A2(G229), .ZN(n928) );
  XOR2_X1 U1022 ( .A(KEYINPUT115), .B(n928), .Z(n929) );
  XNOR2_X1 U1023 ( .A(n929), .B(KEYINPUT49), .ZN(n930) );
  NOR2_X1 U1024 ( .A1(n931), .A2(n930), .ZN(n933) );
  NOR2_X1 U1025 ( .A1(G395), .A2(G397), .ZN(n932) );
  NAND2_X1 U1026 ( .A1(n933), .A2(n932), .ZN(G225) );
  XOR2_X1 U1027 ( .A(KEYINPUT116), .B(G225), .Z(G308) );
  INV_X1 U1029 ( .A(G120), .ZN(G236) );
  INV_X1 U1030 ( .A(G96), .ZN(G221) );
  INV_X1 U1031 ( .A(G69), .ZN(G235) );
  NOR2_X1 U1032 ( .A1(n935), .A2(n934), .ZN(G325) );
  INV_X1 U1033 ( .A(G325), .ZN(G261) );
  INV_X1 U1034 ( .A(G108), .ZN(G238) );
  INV_X1 U1035 ( .A(n936), .ZN(G401) );
  XOR2_X1 U1036 ( .A(KEYINPUT55), .B(KEYINPUT120), .Z(n957) );
  XOR2_X1 U1037 ( .A(KEYINPUT54), .B(G34), .Z(n937) );
  XNOR2_X1 U1038 ( .A(n937), .B(G2084), .ZN(n953) );
  XNOR2_X1 U1039 ( .A(G2090), .B(G35), .ZN(n951) );
  XNOR2_X1 U1040 ( .A(G26), .B(n938), .ZN(n939) );
  NAND2_X1 U1041 ( .A1(n939), .A2(G28), .ZN(n948) );
  XNOR2_X1 U1042 ( .A(G1996), .B(G32), .ZN(n941) );
  XNOR2_X1 U1043 ( .A(G33), .B(G2072), .ZN(n940) );
  NOR2_X1 U1044 ( .A1(n941), .A2(n940), .ZN(n946) );
  XNOR2_X1 U1045 ( .A(G1991), .B(G25), .ZN(n944) );
  XNOR2_X1 U1046 ( .A(G27), .B(n942), .ZN(n943) );
  NOR2_X1 U1047 ( .A1(n944), .A2(n943), .ZN(n945) );
  NAND2_X1 U1048 ( .A1(n946), .A2(n945), .ZN(n947) );
  NOR2_X1 U1049 ( .A1(n948), .A2(n947), .ZN(n949) );
  XNOR2_X1 U1050 ( .A(KEYINPUT53), .B(n949), .ZN(n950) );
  NOR2_X1 U1051 ( .A1(n951), .A2(n950), .ZN(n952) );
  NAND2_X1 U1052 ( .A1(n953), .A2(n952), .ZN(n955) );
  INV_X1 U1053 ( .A(G29), .ZN(n954) );
  NAND2_X1 U1054 ( .A1(n955), .A2(n954), .ZN(n956) );
  XNOR2_X1 U1055 ( .A(n957), .B(n956), .ZN(n984) );
  XNOR2_X1 U1056 ( .A(KEYINPUT52), .B(KEYINPUT119), .ZN(n982) );
  XOR2_X1 U1057 ( .A(G2090), .B(G162), .Z(n958) );
  NOR2_X1 U1058 ( .A1(n959), .A2(n958), .ZN(n960) );
  XOR2_X1 U1059 ( .A(KEYINPUT118), .B(n960), .Z(n961) );
  XNOR2_X1 U1060 ( .A(KEYINPUT51), .B(n961), .ZN(n966) );
  NOR2_X1 U1061 ( .A1(n963), .A2(n962), .ZN(n964) );
  XOR2_X1 U1062 ( .A(KEYINPUT117), .B(n964), .Z(n965) );
  NAND2_X1 U1063 ( .A1(n966), .A2(n965), .ZN(n972) );
  XOR2_X1 U1064 ( .A(G2072), .B(n967), .Z(n969) );
  XOR2_X1 U1065 ( .A(G164), .B(G2078), .Z(n968) );
  NOR2_X1 U1066 ( .A1(n969), .A2(n968), .ZN(n970) );
  XOR2_X1 U1067 ( .A(KEYINPUT50), .B(n970), .Z(n971) );
  NOR2_X1 U1068 ( .A1(n972), .A2(n971), .ZN(n978) );
  NAND2_X1 U1069 ( .A1(n974), .A2(n973), .ZN(n976) );
  XOR2_X1 U1070 ( .A(G2084), .B(G160), .Z(n975) );
  NOR2_X1 U1071 ( .A1(n976), .A2(n975), .ZN(n977) );
  NAND2_X1 U1072 ( .A1(n978), .A2(n977), .ZN(n979) );
  NOR2_X1 U1073 ( .A1(n980), .A2(n979), .ZN(n981) );
  XNOR2_X1 U1074 ( .A(n982), .B(n981), .ZN(n983) );
  NAND2_X1 U1075 ( .A1(n984), .A2(n529), .ZN(n1041) );
  XNOR2_X1 U1076 ( .A(G16), .B(KEYINPUT56), .ZN(n1008) );
  XNOR2_X1 U1077 ( .A(G171), .B(G1961), .ZN(n989) );
  XNOR2_X1 U1078 ( .A(G1341), .B(n985), .ZN(n986) );
  NOR2_X1 U1079 ( .A1(n987), .A2(n986), .ZN(n988) );
  NAND2_X1 U1080 ( .A1(n989), .A2(n988), .ZN(n992) );
  XNOR2_X1 U1081 ( .A(G1348), .B(n990), .ZN(n991) );
  NOR2_X1 U1082 ( .A1(n992), .A2(n991), .ZN(n1006) );
  XNOR2_X1 U1083 ( .A(G1971), .B(G166), .ZN(n994) );
  NAND2_X1 U1084 ( .A1(n994), .A2(n993), .ZN(n996) );
  XNOR2_X1 U1085 ( .A(G1956), .B(G299), .ZN(n995) );
  NOR2_X1 U1086 ( .A1(n996), .A2(n995), .ZN(n998) );
  NAND2_X1 U1087 ( .A1(n998), .A2(n997), .ZN(n999) );
  XOR2_X1 U1088 ( .A(KEYINPUT121), .B(n999), .Z(n1004) );
  XNOR2_X1 U1089 ( .A(G168), .B(G1966), .ZN(n1001) );
  NAND2_X1 U1090 ( .A1(n1001), .A2(n1000), .ZN(n1002) );
  XOR2_X1 U1091 ( .A(KEYINPUT57), .B(n1002), .Z(n1003) );
  NOR2_X1 U1092 ( .A1(n1004), .A2(n1003), .ZN(n1005) );
  NAND2_X1 U1093 ( .A1(n1006), .A2(n1005), .ZN(n1007) );
  NAND2_X1 U1094 ( .A1(n1008), .A2(n1007), .ZN(n1038) );
  INV_X1 U1095 ( .A(G16), .ZN(n1036) );
  XOR2_X1 U1096 ( .A(G1966), .B(G21), .Z(n1022) );
  XNOR2_X1 U1097 ( .A(G1981), .B(G6), .ZN(n1010) );
  XNOR2_X1 U1098 ( .A(G1341), .B(G19), .ZN(n1009) );
  NOR2_X1 U1099 ( .A1(n1010), .A2(n1009), .ZN(n1011) );
  XOR2_X1 U1100 ( .A(KEYINPUT122), .B(n1011), .Z(n1014) );
  XOR2_X1 U1101 ( .A(n1012), .B(G20), .Z(n1013) );
  NOR2_X1 U1102 ( .A1(n1014), .A2(n1013), .ZN(n1018) );
  XOR2_X1 U1103 ( .A(KEYINPUT123), .B(G4), .Z(n1016) );
  XNOR2_X1 U1104 ( .A(G1348), .B(KEYINPUT59), .ZN(n1015) );
  XNOR2_X1 U1105 ( .A(n1016), .B(n1015), .ZN(n1017) );
  NAND2_X1 U1106 ( .A1(n1018), .A2(n1017), .ZN(n1019) );
  XOR2_X1 U1107 ( .A(KEYINPUT60), .B(n1019), .Z(n1020) );
  XNOR2_X1 U1108 ( .A(n1020), .B(KEYINPUT124), .ZN(n1021) );
  NAND2_X1 U1109 ( .A1(n1022), .A2(n1021), .ZN(n1023) );
  XNOR2_X1 U1110 ( .A(n1023), .B(KEYINPUT125), .ZN(n1031) );
  XOR2_X1 U1111 ( .A(G1971), .B(KEYINPUT126), .Z(n1024) );
  XNOR2_X1 U1112 ( .A(G22), .B(n1024), .ZN(n1028) );
  XNOR2_X1 U1113 ( .A(G1986), .B(G24), .ZN(n1026) );
  XNOR2_X1 U1114 ( .A(G23), .B(G1976), .ZN(n1025) );
  NOR2_X1 U1115 ( .A1(n1026), .A2(n1025), .ZN(n1027) );
  NAND2_X1 U1116 ( .A1(n1028), .A2(n1027), .ZN(n1029) );
  XOR2_X1 U1117 ( .A(KEYINPUT58), .B(n1029), .Z(n1030) );
  NAND2_X1 U1118 ( .A1(n1031), .A2(n1030), .ZN(n1033) );
  XNOR2_X1 U1119 ( .A(G5), .B(G1961), .ZN(n1032) );
  NOR2_X1 U1120 ( .A1(n1033), .A2(n1032), .ZN(n1034) );
  XNOR2_X1 U1121 ( .A(KEYINPUT61), .B(n1034), .ZN(n1035) );
  NAND2_X1 U1122 ( .A1(n1036), .A2(n1035), .ZN(n1037) );
  NAND2_X1 U1123 ( .A1(n1038), .A2(n1037), .ZN(n1039) );
  XOR2_X1 U1124 ( .A(KEYINPUT127), .B(n1039), .Z(n1040) );
  NOR2_X1 U1125 ( .A1(n1041), .A2(n1040), .ZN(n1042) );
  NAND2_X1 U1126 ( .A1(n1042), .A2(G11), .ZN(n1043) );
  XOR2_X1 U1127 ( .A(KEYINPUT62), .B(n1043), .Z(G311) );
  INV_X1 U1128 ( .A(G311), .ZN(G150) );
endmodule

