//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 1 0 0 1 1 1 1 1 0 1 1 0 1 0 1 1 1 1 0 0 1 0 0 1 0 1 1 0 1 0 1 0 1 1 0 1 0 0 0 0 1 0 0 1 0 1 0 0 1 1 1 1 1 1 1 0 1 0 0 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:17:12 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n724,
    new_n725, new_n726, new_n727, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n763, new_n764, new_n765, new_n767, new_n768, new_n769, new_n770,
    new_n772, new_n773, new_n774, new_n775, new_n776, new_n777, new_n778,
    new_n779, new_n780, new_n781, new_n782, new_n783, new_n784, new_n785,
    new_n786, new_n787, new_n788, new_n790, new_n791, new_n793, new_n794,
    new_n795, new_n796, new_n797, new_n798, new_n799, new_n800, new_n801,
    new_n802, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n818, new_n819, new_n820, new_n821, new_n822, new_n823, new_n824,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n878, new_n879, new_n880, new_n881, new_n883, new_n884,
    new_n886, new_n887, new_n888, new_n889, new_n890, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n949, new_n951,
    new_n952, new_n954, new_n955, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n973, new_n974, new_n975, new_n976,
    new_n978, new_n979, new_n980, new_n981, new_n982, new_n984, new_n985,
    new_n986, new_n987, new_n988, new_n989, new_n990, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1006, new_n1007;
  XOR2_X1   g000(.A(G1gat), .B(G29gat), .Z(new_n202));
  XNOR2_X1  g001(.A(G57gat), .B(G85gat), .ZN(new_n203));
  XNOR2_X1  g002(.A(new_n202), .B(new_n203), .ZN(new_n204));
  XNOR2_X1  g003(.A(KEYINPUT77), .B(KEYINPUT0), .ZN(new_n205));
  XOR2_X1   g004(.A(new_n204), .B(new_n205), .Z(new_n206));
  INV_X1    g005(.A(new_n206), .ZN(new_n207));
  XNOR2_X1  g006(.A(G127gat), .B(G134gat), .ZN(new_n208));
  INV_X1    g007(.A(KEYINPUT1), .ZN(new_n209));
  NAND2_X1  g008(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  INV_X1    g009(.A(G113gat), .ZN(new_n211));
  NOR2_X1   g010(.A1(new_n211), .A2(G120gat), .ZN(new_n212));
  XOR2_X1   g011(.A(KEYINPUT66), .B(G113gat), .Z(new_n213));
  AOI21_X1  g012(.A(new_n212), .B1(new_n213), .B2(G120gat), .ZN(new_n214));
  OR2_X1    g013(.A1(new_n214), .A2(KEYINPUT67), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n214), .A2(KEYINPUT67), .ZN(new_n216));
  AOI21_X1  g015(.A(new_n210), .B1(new_n215), .B2(new_n216), .ZN(new_n217));
  INV_X1    g016(.A(new_n217), .ZN(new_n218));
  INV_X1    g017(.A(new_n212), .ZN(new_n219));
  INV_X1    g018(.A(G120gat), .ZN(new_n220));
  NOR2_X1   g019(.A1(new_n220), .A2(G113gat), .ZN(new_n221));
  INV_X1    g020(.A(new_n221), .ZN(new_n222));
  AOI21_X1  g021(.A(KEYINPUT1), .B1(new_n219), .B2(new_n222), .ZN(new_n223));
  AND2_X1   g022(.A1(new_n208), .A2(KEYINPUT65), .ZN(new_n224));
  NOR2_X1   g023(.A1(new_n208), .A2(KEYINPUT65), .ZN(new_n225));
  NOR3_X1   g024(.A1(new_n223), .A2(new_n224), .A3(new_n225), .ZN(new_n226));
  INV_X1    g025(.A(new_n226), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n218), .A2(new_n227), .ZN(new_n228));
  XNOR2_X1  g027(.A(G155gat), .B(G162gat), .ZN(new_n229));
  OR2_X1    g028(.A1(new_n229), .A2(KEYINPUT74), .ZN(new_n230));
  INV_X1    g029(.A(KEYINPUT73), .ZN(new_n231));
  INV_X1    g030(.A(G148gat), .ZN(new_n232));
  OAI21_X1  g031(.A(new_n231), .B1(new_n232), .B2(G141gat), .ZN(new_n233));
  INV_X1    g032(.A(G141gat), .ZN(new_n234));
  NAND3_X1  g033(.A1(new_n234), .A2(KEYINPUT73), .A3(G148gat), .ZN(new_n235));
  OAI211_X1 g034(.A(new_n233), .B(new_n235), .C1(new_n234), .C2(G148gat), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n229), .A2(KEYINPUT74), .ZN(new_n237));
  INV_X1    g036(.A(G155gat), .ZN(new_n238));
  INV_X1    g037(.A(G162gat), .ZN(new_n239));
  OAI21_X1  g038(.A(KEYINPUT2), .B1(new_n238), .B2(new_n239), .ZN(new_n240));
  NAND4_X1  g039(.A1(new_n230), .A2(new_n236), .A3(new_n237), .A4(new_n240), .ZN(new_n241));
  INV_X1    g040(.A(new_n229), .ZN(new_n242));
  XNOR2_X1  g041(.A(G141gat), .B(G148gat), .ZN(new_n243));
  OAI21_X1  g042(.A(new_n242), .B1(KEYINPUT2), .B2(new_n243), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n241), .A2(new_n244), .ZN(new_n245));
  NAND2_X1  g044(.A1(new_n228), .A2(new_n245), .ZN(new_n246));
  INV_X1    g045(.A(new_n245), .ZN(new_n247));
  NAND3_X1  g046(.A1(new_n218), .A2(new_n247), .A3(new_n227), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n246), .A2(new_n248), .ZN(new_n249));
  NAND2_X1  g048(.A1(G225gat), .A2(G233gat), .ZN(new_n250));
  INV_X1    g049(.A(new_n250), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n249), .A2(new_n251), .ZN(new_n252));
  XOR2_X1   g051(.A(KEYINPUT76), .B(KEYINPUT5), .Z(new_n253));
  INV_X1    g052(.A(new_n253), .ZN(new_n254));
  NAND2_X1  g053(.A1(new_n252), .A2(new_n254), .ZN(new_n255));
  INV_X1    g054(.A(KEYINPUT4), .ZN(new_n256));
  NAND4_X1  g055(.A1(new_n218), .A2(new_n256), .A3(new_n247), .A4(new_n227), .ZN(new_n257));
  OR2_X1    g056(.A1(new_n257), .A2(KEYINPUT75), .ZN(new_n258));
  NAND2_X1  g057(.A1(new_n257), .A2(KEYINPUT75), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n248), .A2(KEYINPUT4), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  INV_X1    g061(.A(KEYINPUT3), .ZN(new_n263));
  NAND2_X1  g062(.A1(new_n247), .A2(new_n263), .ZN(new_n264));
  NAND2_X1  g063(.A1(new_n245), .A2(KEYINPUT3), .ZN(new_n265));
  NAND3_X1  g064(.A1(new_n228), .A2(new_n264), .A3(new_n265), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n266), .A2(new_n250), .ZN(new_n267));
  INV_X1    g066(.A(new_n267), .ZN(new_n268));
  AOI21_X1  g067(.A(new_n255), .B1(new_n262), .B2(new_n268), .ZN(new_n269));
  INV_X1    g068(.A(new_n266), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n257), .A2(KEYINPUT78), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n271), .A2(new_n261), .ZN(new_n272));
  NAND3_X1  g071(.A1(new_n248), .A2(KEYINPUT78), .A3(KEYINPUT4), .ZN(new_n273));
  AOI21_X1  g072(.A(new_n270), .B1(new_n272), .B2(new_n273), .ZN(new_n274));
  NOR2_X1   g073(.A1(new_n254), .A2(new_n251), .ZN(new_n275));
  AND2_X1   g074(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  OAI21_X1  g075(.A(new_n207), .B1(new_n269), .B2(new_n276), .ZN(new_n277));
  INV_X1    g076(.A(KEYINPUT6), .ZN(new_n278));
  AOI22_X1  g077(.A1(new_n258), .A2(new_n259), .B1(KEYINPUT4), .B2(new_n248), .ZN(new_n279));
  OAI211_X1 g078(.A(new_n252), .B(new_n254), .C1(new_n279), .C2(new_n267), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n274), .A2(new_n275), .ZN(new_n281));
  NAND3_X1  g080(.A1(new_n280), .A2(new_n206), .A3(new_n281), .ZN(new_n282));
  NAND3_X1  g081(.A1(new_n277), .A2(new_n278), .A3(new_n282), .ZN(new_n283));
  AOI21_X1  g082(.A(new_n206), .B1(new_n280), .B2(new_n281), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n284), .A2(KEYINPUT6), .ZN(new_n285));
  OAI21_X1  g084(.A(KEYINPUT64), .B1(G169gat), .B2(G176gat), .ZN(new_n286));
  XNOR2_X1  g085(.A(new_n286), .B(KEYINPUT23), .ZN(new_n287));
  INV_X1    g086(.A(KEYINPUT24), .ZN(new_n288));
  NAND3_X1  g087(.A1(new_n288), .A2(G183gat), .A3(G190gat), .ZN(new_n289));
  INV_X1    g088(.A(G169gat), .ZN(new_n290));
  INV_X1    g089(.A(G176gat), .ZN(new_n291));
  OAI21_X1  g090(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n292));
  AND2_X1   g091(.A1(G183gat), .A2(G190gat), .ZN(new_n293));
  OAI221_X1 g092(.A(new_n289), .B1(new_n290), .B2(new_n291), .C1(new_n292), .C2(new_n293), .ZN(new_n294));
  NOR2_X1   g093(.A1(new_n287), .A2(new_n294), .ZN(new_n295));
  XNOR2_X1  g094(.A(new_n295), .B(KEYINPUT25), .ZN(new_n296));
  XNOR2_X1  g095(.A(KEYINPUT27), .B(G183gat), .ZN(new_n297));
  INV_X1    g096(.A(G190gat), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n297), .A2(new_n298), .ZN(new_n299));
  XOR2_X1   g098(.A(new_n299), .B(KEYINPUT28), .Z(new_n300));
  NAND2_X1  g099(.A1(new_n290), .A2(new_n291), .ZN(new_n301));
  NOR2_X1   g100(.A1(new_n290), .A2(new_n291), .ZN(new_n302));
  OAI21_X1  g101(.A(new_n301), .B1(new_n302), .B2(KEYINPUT26), .ZN(new_n303));
  OR2_X1    g102(.A1(new_n301), .A2(KEYINPUT26), .ZN(new_n304));
  AOI21_X1  g103(.A(new_n293), .B1(new_n303), .B2(new_n304), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n300), .A2(new_n305), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n296), .A2(new_n306), .ZN(new_n307));
  NAND2_X1  g106(.A1(G226gat), .A2(G233gat), .ZN(new_n308));
  XOR2_X1   g107(.A(new_n308), .B(KEYINPUT71), .Z(new_n309));
  NOR2_X1   g108(.A1(new_n309), .A2(KEYINPUT29), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n307), .A2(new_n310), .ZN(new_n311));
  XNOR2_X1  g110(.A(new_n307), .B(KEYINPUT72), .ZN(new_n312));
  INV_X1    g111(.A(new_n309), .ZN(new_n313));
  OAI21_X1  g112(.A(new_n311), .B1(new_n312), .B2(new_n313), .ZN(new_n314));
  XNOR2_X1  g113(.A(G197gat), .B(G204gat), .ZN(new_n315));
  INV_X1    g114(.A(G211gat), .ZN(new_n316));
  INV_X1    g115(.A(G218gat), .ZN(new_n317));
  NOR2_X1   g116(.A1(new_n316), .A2(new_n317), .ZN(new_n318));
  OAI21_X1  g117(.A(new_n315), .B1(KEYINPUT22), .B2(new_n318), .ZN(new_n319));
  XOR2_X1   g118(.A(G211gat), .B(G218gat), .Z(new_n320));
  OR2_X1    g119(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  XNOR2_X1  g120(.A(new_n321), .B(KEYINPUT70), .ZN(new_n322));
  XNOR2_X1  g121(.A(new_n320), .B(KEYINPUT69), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n323), .A2(new_n319), .ZN(new_n324));
  AND2_X1   g123(.A1(new_n322), .A2(new_n324), .ZN(new_n325));
  INV_X1    g124(.A(new_n325), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n314), .A2(new_n326), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n312), .A2(new_n310), .ZN(new_n328));
  AND2_X1   g127(.A1(new_n296), .A2(new_n306), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n329), .A2(new_n309), .ZN(new_n330));
  NAND3_X1  g129(.A1(new_n328), .A2(new_n325), .A3(new_n330), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n327), .A2(new_n331), .ZN(new_n332));
  XNOR2_X1  g131(.A(G8gat), .B(G36gat), .ZN(new_n333));
  XNOR2_X1  g132(.A(G64gat), .B(G92gat), .ZN(new_n334));
  XNOR2_X1  g133(.A(new_n333), .B(new_n334), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n332), .A2(new_n335), .ZN(new_n336));
  INV_X1    g135(.A(new_n335), .ZN(new_n337));
  NAND3_X1  g136(.A1(new_n327), .A2(new_n331), .A3(new_n337), .ZN(new_n338));
  NAND3_X1  g137(.A1(new_n336), .A2(KEYINPUT30), .A3(new_n338), .ZN(new_n339));
  OR2_X1    g138(.A1(new_n338), .A2(KEYINPUT30), .ZN(new_n340));
  AOI22_X1  g139(.A1(new_n283), .A2(new_n285), .B1(new_n339), .B2(new_n340), .ZN(new_n341));
  INV_X1    g140(.A(G22gat), .ZN(new_n342));
  AND2_X1   g141(.A1(G228gat), .A2(G233gat), .ZN(new_n343));
  INV_X1    g142(.A(new_n343), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n319), .A2(new_n320), .ZN(new_n345));
  AOI21_X1  g144(.A(KEYINPUT29), .B1(new_n322), .B2(new_n345), .ZN(new_n346));
  OR2_X1    g145(.A1(new_n346), .A2(KEYINPUT80), .ZN(new_n347));
  AOI21_X1  g146(.A(KEYINPUT3), .B1(new_n346), .B2(KEYINPUT80), .ZN(new_n348));
  AOI21_X1  g147(.A(new_n247), .B1(new_n347), .B2(new_n348), .ZN(new_n349));
  INV_X1    g148(.A(KEYINPUT29), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n264), .A2(new_n350), .ZN(new_n351));
  AND2_X1   g150(.A1(new_n325), .A2(new_n351), .ZN(new_n352));
  OAI21_X1  g151(.A(new_n344), .B1(new_n349), .B2(new_n352), .ZN(new_n353));
  OAI21_X1  g152(.A(new_n263), .B1(new_n325), .B2(KEYINPUT29), .ZN(new_n354));
  AOI21_X1  g153(.A(new_n344), .B1(new_n354), .B2(new_n245), .ZN(new_n355));
  XOR2_X1   g154(.A(new_n351), .B(KEYINPUT81), .Z(new_n356));
  OAI21_X1  g155(.A(new_n355), .B1(new_n356), .B2(new_n326), .ZN(new_n357));
  AOI21_X1  g156(.A(new_n342), .B1(new_n353), .B2(new_n357), .ZN(new_n358));
  NAND3_X1  g157(.A1(new_n353), .A2(new_n357), .A3(new_n342), .ZN(new_n359));
  AOI21_X1  g158(.A(new_n358), .B1(KEYINPUT82), .B2(new_n359), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n353), .A2(new_n357), .ZN(new_n361));
  NAND3_X1  g160(.A1(new_n361), .A2(KEYINPUT82), .A3(G22gat), .ZN(new_n362));
  XNOR2_X1  g161(.A(G78gat), .B(G106gat), .ZN(new_n363));
  XNOR2_X1  g162(.A(KEYINPUT31), .B(G50gat), .ZN(new_n364));
  XNOR2_X1  g163(.A(new_n363), .B(new_n364), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n362), .A2(new_n365), .ZN(new_n366));
  INV_X1    g165(.A(new_n359), .ZN(new_n367));
  NOR2_X1   g166(.A1(new_n367), .A2(new_n358), .ZN(new_n368));
  XOR2_X1   g167(.A(new_n365), .B(KEYINPUT79), .Z(new_n369));
  OAI22_X1  g168(.A1(new_n360), .A2(new_n366), .B1(new_n368), .B2(new_n369), .ZN(new_n370));
  XNOR2_X1  g169(.A(G15gat), .B(G43gat), .ZN(new_n371));
  XNOR2_X1  g170(.A(G71gat), .B(G99gat), .ZN(new_n372));
  XNOR2_X1  g171(.A(new_n371), .B(new_n372), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n329), .A2(new_n228), .ZN(new_n374));
  NAND3_X1  g173(.A1(new_n307), .A2(new_n227), .A3(new_n218), .ZN(new_n375));
  NAND4_X1  g174(.A1(new_n374), .A2(G227gat), .A3(G233gat), .A4(new_n375), .ZN(new_n376));
  INV_X1    g175(.A(KEYINPUT33), .ZN(new_n377));
  AOI21_X1  g176(.A(new_n373), .B1(new_n376), .B2(new_n377), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n376), .A2(KEYINPUT32), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n378), .A2(new_n379), .ZN(new_n380));
  OAI211_X1 g179(.A(new_n376), .B(KEYINPUT32), .C1(new_n377), .C2(new_n373), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n380), .A2(new_n381), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n374), .A2(new_n375), .ZN(new_n383));
  NAND2_X1  g182(.A1(G227gat), .A2(G233gat), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  OR2_X1    g184(.A1(new_n385), .A2(KEYINPUT34), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n385), .A2(KEYINPUT34), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n382), .A2(new_n388), .ZN(new_n389));
  NAND4_X1  g188(.A1(new_n380), .A2(new_n386), .A3(new_n387), .A4(new_n381), .ZN(new_n390));
  AND2_X1   g189(.A1(new_n389), .A2(new_n390), .ZN(new_n391));
  NAND3_X1  g190(.A1(new_n341), .A2(new_n370), .A3(new_n391), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n392), .A2(KEYINPUT35), .ZN(new_n393));
  INV_X1    g192(.A(KEYINPUT87), .ZN(new_n394));
  INV_X1    g193(.A(KEYINPUT68), .ZN(new_n395));
  NAND3_X1  g194(.A1(new_n382), .A2(new_n388), .A3(new_n395), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n396), .A2(new_n390), .ZN(new_n397));
  AOI21_X1  g196(.A(new_n395), .B1(new_n382), .B2(new_n388), .ZN(new_n398));
  OAI21_X1  g197(.A(new_n394), .B1(new_n397), .B2(new_n398), .ZN(new_n399));
  INV_X1    g198(.A(new_n398), .ZN(new_n400));
  NAND4_X1  g199(.A1(new_n400), .A2(KEYINPUT87), .A3(new_n390), .A4(new_n396), .ZN(new_n401));
  NAND3_X1  g200(.A1(new_n370), .A2(new_n399), .A3(new_n401), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n285), .A2(KEYINPUT85), .ZN(new_n403));
  INV_X1    g202(.A(KEYINPUT85), .ZN(new_n404));
  NAND3_X1  g203(.A1(new_n284), .A2(new_n404), .A3(KEYINPUT6), .ZN(new_n405));
  NAND3_X1  g204(.A1(new_n403), .A2(new_n283), .A3(new_n405), .ZN(new_n406));
  INV_X1    g205(.A(KEYINPUT35), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n339), .A2(new_n340), .ZN(new_n408));
  NAND3_X1  g207(.A1(new_n406), .A2(new_n407), .A3(new_n408), .ZN(new_n409));
  OAI21_X1  g208(.A(new_n393), .B1(new_n402), .B2(new_n409), .ZN(new_n410));
  INV_X1    g209(.A(KEYINPUT38), .ZN(new_n411));
  INV_X1    g210(.A(KEYINPUT37), .ZN(new_n412));
  NAND3_X1  g211(.A1(new_n327), .A2(new_n412), .A3(new_n331), .ZN(new_n413));
  INV_X1    g212(.A(new_n413), .ZN(new_n414));
  AOI21_X1  g213(.A(new_n412), .B1(new_n327), .B2(new_n331), .ZN(new_n415));
  NOR2_X1   g214(.A1(new_n415), .A2(new_n337), .ZN(new_n416));
  INV_X1    g215(.A(KEYINPUT86), .ZN(new_n417));
  AOI21_X1  g216(.A(new_n414), .B1(new_n416), .B2(new_n417), .ZN(new_n418));
  OAI21_X1  g217(.A(KEYINPUT86), .B1(new_n415), .B2(new_n337), .ZN(new_n419));
  AOI21_X1  g218(.A(new_n411), .B1(new_n418), .B2(new_n419), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n314), .A2(new_n325), .ZN(new_n421));
  NAND3_X1  g220(.A1(new_n328), .A2(new_n326), .A3(new_n330), .ZN(new_n422));
  NAND3_X1  g221(.A1(new_n421), .A2(KEYINPUT37), .A3(new_n422), .ZN(new_n423));
  NAND4_X1  g222(.A1(new_n413), .A2(new_n423), .A3(new_n411), .A4(new_n335), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n424), .A2(new_n338), .ZN(new_n425));
  NOR3_X1   g224(.A1(new_n406), .A2(new_n420), .A3(new_n425), .ZN(new_n426));
  INV_X1    g225(.A(new_n408), .ZN(new_n427));
  INV_X1    g226(.A(KEYINPUT84), .ZN(new_n428));
  NAND3_X1  g227(.A1(new_n246), .A2(new_n248), .A3(new_n250), .ZN(new_n429));
  INV_X1    g228(.A(KEYINPUT83), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n429), .A2(new_n430), .ZN(new_n431));
  INV_X1    g230(.A(new_n431), .ZN(new_n432));
  OAI21_X1  g231(.A(KEYINPUT39), .B1(new_n429), .B2(new_n430), .ZN(new_n433));
  OAI21_X1  g232(.A(new_n428), .B1(new_n432), .B2(new_n433), .ZN(new_n434));
  OR2_X1    g233(.A1(new_n429), .A2(new_n430), .ZN(new_n435));
  NAND4_X1  g234(.A1(new_n435), .A2(KEYINPUT84), .A3(KEYINPUT39), .A4(new_n431), .ZN(new_n436));
  OAI211_X1 g235(.A(new_n434), .B(new_n436), .C1(new_n250), .C2(new_n274), .ZN(new_n437));
  NOR3_X1   g236(.A1(new_n274), .A2(KEYINPUT39), .A3(new_n250), .ZN(new_n438));
  NOR2_X1   g237(.A1(new_n438), .A2(new_n207), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n437), .A2(new_n439), .ZN(new_n440));
  INV_X1    g239(.A(KEYINPUT40), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n440), .A2(new_n441), .ZN(new_n442));
  NAND3_X1  g241(.A1(new_n437), .A2(KEYINPUT40), .A3(new_n439), .ZN(new_n443));
  NAND4_X1  g242(.A1(new_n427), .A2(new_n442), .A3(new_n277), .A4(new_n443), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n444), .A2(new_n370), .ZN(new_n445));
  NOR2_X1   g244(.A1(new_n426), .A2(new_n445), .ZN(new_n446));
  INV_X1    g245(.A(KEYINPUT36), .ZN(new_n447));
  OAI21_X1  g246(.A(new_n447), .B1(new_n397), .B2(new_n398), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n391), .A2(KEYINPUT36), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n448), .A2(new_n449), .ZN(new_n450));
  OAI21_X1  g249(.A(new_n450), .B1(new_n341), .B2(new_n370), .ZN(new_n451));
  OAI21_X1  g250(.A(new_n410), .B1(new_n446), .B2(new_n451), .ZN(new_n452));
  INV_X1    g251(.A(KEYINPUT90), .ZN(new_n453));
  XNOR2_X1  g252(.A(G15gat), .B(G22gat), .ZN(new_n454));
  INV_X1    g253(.A(G1gat), .ZN(new_n455));
  AND2_X1   g254(.A1(new_n455), .A2(KEYINPUT16), .ZN(new_n456));
  AND2_X1   g255(.A1(new_n454), .A2(new_n456), .ZN(new_n457));
  NOR2_X1   g256(.A1(new_n454), .A2(new_n455), .ZN(new_n458));
  OAI21_X1  g257(.A(G8gat), .B1(new_n457), .B2(new_n458), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n454), .A2(new_n456), .ZN(new_n460));
  INV_X1    g259(.A(G8gat), .ZN(new_n461));
  OAI211_X1 g260(.A(new_n460), .B(new_n461), .C1(new_n455), .C2(new_n454), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n459), .A2(new_n462), .ZN(new_n463));
  INV_X1    g262(.A(KEYINPUT15), .ZN(new_n464));
  INV_X1    g263(.A(G36gat), .ZN(new_n465));
  OR2_X1    g264(.A1(KEYINPUT89), .A2(G29gat), .ZN(new_n466));
  NAND2_X1  g265(.A1(KEYINPUT89), .A2(G29gat), .ZN(new_n467));
  AOI21_X1  g266(.A(new_n465), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  INV_X1    g267(.A(G29gat), .ZN(new_n469));
  NAND3_X1  g268(.A1(new_n469), .A2(new_n465), .A3(KEYINPUT14), .ZN(new_n470));
  INV_X1    g269(.A(KEYINPUT14), .ZN(new_n471));
  OAI21_X1  g270(.A(new_n471), .B1(G29gat), .B2(G36gat), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n470), .A2(new_n472), .ZN(new_n473));
  OAI21_X1  g272(.A(new_n464), .B1(new_n468), .B2(new_n473), .ZN(new_n474));
  XOR2_X1   g273(.A(G43gat), .B(G50gat), .Z(new_n475));
  INV_X1    g274(.A(new_n475), .ZN(new_n476));
  AND2_X1   g275(.A1(KEYINPUT89), .A2(G29gat), .ZN(new_n477));
  NOR2_X1   g276(.A1(KEYINPUT89), .A2(G29gat), .ZN(new_n478));
  OAI21_X1  g277(.A(G36gat), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  NAND4_X1  g278(.A1(new_n479), .A2(KEYINPUT15), .A3(new_n472), .A4(new_n470), .ZN(new_n480));
  NAND3_X1  g279(.A1(new_n474), .A2(new_n476), .A3(new_n480), .ZN(new_n481));
  INV_X1    g280(.A(KEYINPUT17), .ZN(new_n482));
  NOR2_X1   g281(.A1(new_n468), .A2(new_n473), .ZN(new_n483));
  NAND3_X1  g282(.A1(new_n483), .A2(KEYINPUT15), .A3(new_n475), .ZN(new_n484));
  AND3_X1   g283(.A1(new_n481), .A2(new_n482), .A3(new_n484), .ZN(new_n485));
  AOI21_X1  g284(.A(new_n482), .B1(new_n481), .B2(new_n484), .ZN(new_n486));
  OAI211_X1 g285(.A(new_n453), .B(new_n463), .C1(new_n485), .C2(new_n486), .ZN(new_n487));
  NAND2_X1  g286(.A1(G229gat), .A2(G233gat), .ZN(new_n488));
  AND2_X1   g287(.A1(new_n459), .A2(new_n462), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n481), .A2(new_n484), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n490), .A2(KEYINPUT17), .ZN(new_n491));
  NAND3_X1  g290(.A1(new_n481), .A2(new_n482), .A3(new_n484), .ZN(new_n492));
  AOI21_X1  g291(.A(new_n489), .B1(new_n491), .B2(new_n492), .ZN(new_n493));
  AOI21_X1  g292(.A(KEYINPUT90), .B1(new_n489), .B2(new_n490), .ZN(new_n494));
  OAI211_X1 g293(.A(new_n487), .B(new_n488), .C1(new_n493), .C2(new_n494), .ZN(new_n495));
  INV_X1    g294(.A(KEYINPUT18), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  INV_X1    g296(.A(KEYINPUT91), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  OAI21_X1  g298(.A(new_n463), .B1(new_n485), .B2(new_n486), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n489), .A2(new_n490), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n501), .A2(new_n453), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n500), .A2(new_n502), .ZN(new_n503));
  NAND4_X1  g302(.A1(new_n503), .A2(KEYINPUT18), .A3(new_n488), .A4(new_n487), .ZN(new_n504));
  NAND3_X1  g303(.A1(new_n495), .A2(KEYINPUT91), .A3(new_n496), .ZN(new_n505));
  INV_X1    g304(.A(new_n490), .ZN(new_n506));
  NAND2_X1  g305(.A1(new_n506), .A2(new_n463), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n507), .A2(new_n501), .ZN(new_n508));
  XOR2_X1   g307(.A(new_n488), .B(KEYINPUT13), .Z(new_n509));
  XOR2_X1   g308(.A(KEYINPUT88), .B(KEYINPUT12), .Z(new_n510));
  XNOR2_X1  g309(.A(G113gat), .B(G141gat), .ZN(new_n511));
  OR2_X1    g310(.A1(new_n511), .A2(KEYINPUT11), .ZN(new_n512));
  NAND2_X1  g311(.A1(new_n511), .A2(KEYINPUT11), .ZN(new_n513));
  NAND3_X1  g312(.A1(new_n512), .A2(new_n290), .A3(new_n513), .ZN(new_n514));
  INV_X1    g313(.A(new_n514), .ZN(new_n515));
  INV_X1    g314(.A(G197gat), .ZN(new_n516));
  AOI21_X1  g315(.A(new_n290), .B1(new_n512), .B2(new_n513), .ZN(new_n517));
  NOR3_X1   g316(.A1(new_n515), .A2(new_n516), .A3(new_n517), .ZN(new_n518));
  NAND2_X1  g317(.A1(new_n512), .A2(new_n513), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n519), .A2(G169gat), .ZN(new_n520));
  AOI21_X1  g319(.A(G197gat), .B1(new_n520), .B2(new_n514), .ZN(new_n521));
  OAI21_X1  g320(.A(new_n510), .B1(new_n518), .B2(new_n521), .ZN(new_n522));
  OAI21_X1  g321(.A(new_n516), .B1(new_n515), .B2(new_n517), .ZN(new_n523));
  NAND3_X1  g322(.A1(new_n520), .A2(G197gat), .A3(new_n514), .ZN(new_n524));
  INV_X1    g323(.A(new_n510), .ZN(new_n525));
  NAND3_X1  g324(.A1(new_n523), .A2(new_n524), .A3(new_n525), .ZN(new_n526));
  AOI22_X1  g325(.A1(new_n508), .A2(new_n509), .B1(new_n522), .B2(new_n526), .ZN(new_n527));
  NAND4_X1  g326(.A1(new_n499), .A2(new_n504), .A3(new_n505), .A4(new_n527), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n508), .A2(new_n509), .ZN(new_n529));
  NAND3_X1  g328(.A1(new_n497), .A2(new_n504), .A3(new_n529), .ZN(new_n530));
  NAND2_X1  g329(.A1(new_n522), .A2(new_n526), .ZN(new_n531));
  INV_X1    g330(.A(new_n531), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n530), .A2(new_n532), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n528), .A2(new_n533), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n452), .A2(new_n534), .ZN(new_n535));
  XNOR2_X1  g334(.A(G183gat), .B(G211gat), .ZN(new_n536));
  XNOR2_X1  g335(.A(new_n536), .B(KEYINPUT94), .ZN(new_n537));
  INV_X1    g336(.A(new_n537), .ZN(new_n538));
  XOR2_X1   g337(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n539));
  INV_X1    g338(.A(KEYINPUT93), .ZN(new_n540));
  AND2_X1   g339(.A1(G71gat), .A2(G78gat), .ZN(new_n541));
  NOR2_X1   g340(.A1(G71gat), .A2(G78gat), .ZN(new_n542));
  NOR2_X1   g341(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  INV_X1    g342(.A(new_n543), .ZN(new_n544));
  OR2_X1    g343(.A1(G57gat), .A2(G64gat), .ZN(new_n545));
  OR2_X1    g344(.A1(new_n541), .A2(KEYINPUT9), .ZN(new_n546));
  NAND2_X1  g345(.A1(G57gat), .A2(G64gat), .ZN(new_n547));
  NAND4_X1  g346(.A1(new_n544), .A2(new_n545), .A3(new_n546), .A4(new_n547), .ZN(new_n548));
  NAND3_X1  g347(.A1(new_n545), .A2(KEYINPUT9), .A3(new_n547), .ZN(new_n549));
  INV_X1    g348(.A(KEYINPUT92), .ZN(new_n550));
  AND3_X1   g349(.A1(new_n549), .A2(new_n550), .A3(new_n543), .ZN(new_n551));
  AOI21_X1  g350(.A(new_n550), .B1(new_n549), .B2(new_n543), .ZN(new_n552));
  OAI21_X1  g351(.A(new_n548), .B1(new_n551), .B2(new_n552), .ZN(new_n553));
  INV_X1    g352(.A(KEYINPUT21), .ZN(new_n554));
  AOI21_X1  g353(.A(new_n540), .B1(new_n553), .B2(new_n554), .ZN(new_n555));
  INV_X1    g354(.A(new_n555), .ZN(new_n556));
  NAND3_X1  g355(.A1(new_n553), .A2(new_n540), .A3(new_n554), .ZN(new_n557));
  NAND4_X1  g356(.A1(new_n556), .A2(G231gat), .A3(G233gat), .A4(new_n557), .ZN(new_n558));
  NAND2_X1  g357(.A1(G231gat), .A2(G233gat), .ZN(new_n559));
  INV_X1    g358(.A(new_n557), .ZN(new_n560));
  OAI21_X1  g359(.A(new_n559), .B1(new_n560), .B2(new_n555), .ZN(new_n561));
  XNOR2_X1  g360(.A(G127gat), .B(G155gat), .ZN(new_n562));
  NAND3_X1  g361(.A1(new_n558), .A2(new_n561), .A3(new_n562), .ZN(new_n563));
  INV_X1    g362(.A(new_n563), .ZN(new_n564));
  AOI21_X1  g363(.A(new_n562), .B1(new_n558), .B2(new_n561), .ZN(new_n565));
  OAI21_X1  g364(.A(new_n539), .B1(new_n564), .B2(new_n565), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n558), .A2(new_n561), .ZN(new_n567));
  INV_X1    g366(.A(new_n562), .ZN(new_n568));
  NAND2_X1  g367(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  INV_X1    g368(.A(new_n539), .ZN(new_n570));
  NAND3_X1  g369(.A1(new_n569), .A2(new_n563), .A3(new_n570), .ZN(new_n571));
  INV_X1    g370(.A(new_n553), .ZN(new_n572));
  NAND2_X1  g371(.A1(new_n572), .A2(KEYINPUT21), .ZN(new_n573));
  NAND2_X1  g372(.A1(new_n573), .A2(new_n463), .ZN(new_n574));
  AND3_X1   g373(.A1(new_n566), .A2(new_n571), .A3(new_n574), .ZN(new_n575));
  AOI21_X1  g374(.A(new_n574), .B1(new_n566), .B2(new_n571), .ZN(new_n576));
  OAI21_X1  g375(.A(new_n538), .B1(new_n575), .B2(new_n576), .ZN(new_n577));
  NAND2_X1  g376(.A1(new_n566), .A2(new_n571), .ZN(new_n578));
  INV_X1    g377(.A(new_n574), .ZN(new_n579));
  NAND2_X1  g378(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  NAND3_X1  g379(.A1(new_n566), .A2(new_n571), .A3(new_n574), .ZN(new_n581));
  NAND3_X1  g380(.A1(new_n580), .A2(new_n581), .A3(new_n537), .ZN(new_n582));
  NAND2_X1  g381(.A1(new_n577), .A2(new_n582), .ZN(new_n583));
  INV_X1    g382(.A(KEYINPUT98), .ZN(new_n584));
  XNOR2_X1  g383(.A(G190gat), .B(G218gat), .ZN(new_n585));
  INV_X1    g384(.A(new_n585), .ZN(new_n586));
  XOR2_X1   g385(.A(G99gat), .B(G106gat), .Z(new_n587));
  INV_X1    g386(.A(KEYINPUT7), .ZN(new_n588));
  NAND2_X1  g387(.A1(new_n588), .A2(KEYINPUT95), .ZN(new_n589));
  INV_X1    g388(.A(KEYINPUT95), .ZN(new_n590));
  NAND2_X1  g389(.A1(new_n590), .A2(KEYINPUT7), .ZN(new_n591));
  NAND2_X1  g390(.A1(G85gat), .A2(G92gat), .ZN(new_n592));
  NAND3_X1  g391(.A1(new_n589), .A2(new_n591), .A3(new_n592), .ZN(new_n593));
  NAND2_X1  g392(.A1(G99gat), .A2(G106gat), .ZN(new_n594));
  INV_X1    g393(.A(G85gat), .ZN(new_n595));
  INV_X1    g394(.A(G92gat), .ZN(new_n596));
  AOI22_X1  g395(.A1(KEYINPUT8), .A2(new_n594), .B1(new_n595), .B2(new_n596), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n593), .A2(new_n597), .ZN(new_n598));
  AOI21_X1  g397(.A(new_n592), .B1(new_n589), .B2(new_n591), .ZN(new_n599));
  OAI21_X1  g398(.A(new_n587), .B1(new_n598), .B2(new_n599), .ZN(new_n600));
  INV_X1    g399(.A(KEYINPUT96), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  OAI211_X1 g401(.A(KEYINPUT96), .B(new_n587), .C1(new_n598), .C2(new_n599), .ZN(new_n603));
  INV_X1    g402(.A(new_n599), .ZN(new_n604));
  INV_X1    g403(.A(new_n587), .ZN(new_n605));
  NAND4_X1  g404(.A1(new_n604), .A2(new_n605), .A3(new_n593), .A4(new_n597), .ZN(new_n606));
  NAND3_X1  g405(.A1(new_n602), .A2(new_n603), .A3(new_n606), .ZN(new_n607));
  OAI21_X1  g406(.A(new_n607), .B1(new_n485), .B2(new_n486), .ZN(new_n608));
  INV_X1    g407(.A(KEYINPUT97), .ZN(new_n609));
  NAND2_X1  g408(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  OAI211_X1 g409(.A(KEYINPUT97), .B(new_n607), .C1(new_n485), .C2(new_n486), .ZN(new_n611));
  NAND2_X1  g410(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  AND2_X1   g411(.A1(G232gat), .A2(G233gat), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n613), .A2(KEYINPUT41), .ZN(new_n614));
  OAI21_X1  g413(.A(new_n614), .B1(new_n506), .B2(new_n607), .ZN(new_n615));
  INV_X1    g414(.A(new_n615), .ZN(new_n616));
  AOI21_X1  g415(.A(new_n586), .B1(new_n612), .B2(new_n616), .ZN(new_n617));
  AOI211_X1 g416(.A(new_n615), .B(new_n585), .C1(new_n610), .C2(new_n611), .ZN(new_n618));
  OAI21_X1  g417(.A(new_n584), .B1(new_n617), .B2(new_n618), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n491), .A2(new_n492), .ZN(new_n620));
  AOI21_X1  g419(.A(KEYINPUT97), .B1(new_n620), .B2(new_n607), .ZN(new_n621));
  INV_X1    g420(.A(new_n611), .ZN(new_n622));
  OAI21_X1  g421(.A(new_n616), .B1(new_n621), .B2(new_n622), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n623), .A2(new_n585), .ZN(new_n624));
  NAND3_X1  g423(.A1(new_n612), .A2(new_n616), .A3(new_n586), .ZN(new_n625));
  NAND3_X1  g424(.A1(new_n624), .A2(KEYINPUT98), .A3(new_n625), .ZN(new_n626));
  NOR2_X1   g425(.A1(new_n613), .A2(KEYINPUT41), .ZN(new_n627));
  XNOR2_X1  g426(.A(G134gat), .B(G162gat), .ZN(new_n628));
  XOR2_X1   g427(.A(new_n627), .B(new_n628), .Z(new_n629));
  INV_X1    g428(.A(new_n629), .ZN(new_n630));
  NAND3_X1  g429(.A1(new_n619), .A2(new_n626), .A3(new_n630), .ZN(new_n631));
  NAND4_X1  g430(.A1(new_n624), .A2(KEYINPUT98), .A3(new_n629), .A4(new_n625), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  NAND2_X1  g432(.A1(new_n583), .A2(new_n633), .ZN(new_n634));
  NAND2_X1  g433(.A1(G230gat), .A2(G233gat), .ZN(new_n635));
  INV_X1    g434(.A(new_n635), .ZN(new_n636));
  NAND3_X1  g435(.A1(new_n604), .A2(new_n593), .A3(new_n597), .ZN(new_n637));
  AOI21_X1  g436(.A(KEYINPUT96), .B1(new_n637), .B2(new_n587), .ZN(new_n638));
  NAND2_X1  g437(.A1(new_n603), .A2(new_n606), .ZN(new_n639));
  OAI21_X1  g438(.A(new_n553), .B1(new_n638), .B2(new_n639), .ZN(new_n640));
  INV_X1    g439(.A(KEYINPUT10), .ZN(new_n641));
  AND2_X1   g440(.A1(new_n606), .A2(new_n600), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n642), .A2(new_n572), .ZN(new_n643));
  NAND3_X1  g442(.A1(new_n640), .A2(new_n641), .A3(new_n643), .ZN(new_n644));
  NOR2_X1   g443(.A1(new_n638), .A2(new_n639), .ZN(new_n645));
  NAND3_X1  g444(.A1(new_n645), .A2(KEYINPUT10), .A3(new_n572), .ZN(new_n646));
  AOI21_X1  g445(.A(new_n636), .B1(new_n644), .B2(new_n646), .ZN(new_n647));
  XNOR2_X1  g446(.A(G120gat), .B(G148gat), .ZN(new_n648));
  XNOR2_X1  g447(.A(G176gat), .B(G204gat), .ZN(new_n649));
  XNOR2_X1  g448(.A(new_n648), .B(new_n649), .ZN(new_n650));
  NOR2_X1   g449(.A1(new_n647), .A2(new_n650), .ZN(new_n651));
  AND2_X1   g450(.A1(new_n640), .A2(new_n643), .ZN(new_n652));
  NOR2_X1   g451(.A1(new_n652), .A2(new_n635), .ZN(new_n653));
  INV_X1    g452(.A(KEYINPUT99), .ZN(new_n654));
  NOR2_X1   g453(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  NOR3_X1   g454(.A1(new_n652), .A2(KEYINPUT99), .A3(new_n635), .ZN(new_n656));
  OAI21_X1  g455(.A(new_n651), .B1(new_n655), .B2(new_n656), .ZN(new_n657));
  OAI21_X1  g456(.A(new_n650), .B1(new_n653), .B2(new_n647), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  NOR3_X1   g458(.A1(new_n535), .A2(new_n634), .A3(new_n659), .ZN(new_n660));
  AND2_X1   g459(.A1(new_n283), .A2(new_n285), .ZN(new_n661));
  NAND2_X1  g460(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  XNOR2_X1  g461(.A(new_n662), .B(G1gat), .ZN(G1324gat));
  INV_X1    g462(.A(KEYINPUT100), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n660), .A2(new_n427), .ZN(new_n665));
  XNOR2_X1  g464(.A(KEYINPUT16), .B(G8gat), .ZN(new_n666));
  XNOR2_X1  g465(.A(new_n666), .B(KEYINPUT101), .ZN(new_n667));
  OAI21_X1  g466(.A(new_n664), .B1(new_n665), .B2(new_n667), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n668), .A2(KEYINPUT42), .ZN(new_n669));
  INV_X1    g468(.A(KEYINPUT42), .ZN(new_n670));
  OAI211_X1 g469(.A(new_n664), .B(new_n670), .C1(new_n665), .C2(new_n667), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n665), .A2(G8gat), .ZN(new_n672));
  NAND3_X1  g471(.A1(new_n669), .A2(new_n671), .A3(new_n672), .ZN(G1325gat));
  INV_X1    g472(.A(new_n660), .ZN(new_n674));
  XNOR2_X1  g473(.A(new_n450), .B(KEYINPUT102), .ZN(new_n675));
  INV_X1    g474(.A(new_n675), .ZN(new_n676));
  OAI21_X1  g475(.A(G15gat), .B1(new_n674), .B2(new_n676), .ZN(new_n677));
  NAND2_X1  g476(.A1(new_n399), .A2(new_n401), .ZN(new_n678));
  OR2_X1    g477(.A1(new_n678), .A2(G15gat), .ZN(new_n679));
  OAI21_X1  g478(.A(new_n677), .B1(new_n674), .B2(new_n679), .ZN(G1326gat));
  NAND2_X1  g479(.A1(new_n361), .A2(G22gat), .ZN(new_n681));
  AOI21_X1  g480(.A(new_n369), .B1(new_n681), .B2(new_n359), .ZN(new_n682));
  AND2_X1   g481(.A1(new_n362), .A2(new_n365), .ZN(new_n683));
  INV_X1    g482(.A(KEYINPUT82), .ZN(new_n684));
  OAI21_X1  g483(.A(new_n681), .B1(new_n367), .B2(new_n684), .ZN(new_n685));
  AOI21_X1  g484(.A(new_n682), .B1(new_n683), .B2(new_n685), .ZN(new_n686));
  NAND2_X1  g485(.A1(new_n660), .A2(new_n686), .ZN(new_n687));
  XNOR2_X1  g486(.A(KEYINPUT43), .B(G22gat), .ZN(new_n688));
  XNOR2_X1  g487(.A(new_n687), .B(new_n688), .ZN(G1327gat));
  INV_X1    g488(.A(new_n583), .ZN(new_n690));
  INV_X1    g489(.A(new_n659), .ZN(new_n691));
  NAND2_X1  g490(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  NOR3_X1   g491(.A1(new_n535), .A2(new_n633), .A3(new_n692), .ZN(new_n693));
  NAND4_X1  g492(.A1(new_n693), .A2(new_n661), .A3(new_n466), .A4(new_n467), .ZN(new_n694));
  XNOR2_X1  g493(.A(new_n694), .B(KEYINPUT45), .ZN(new_n695));
  AND2_X1   g494(.A1(new_n631), .A2(new_n632), .ZN(new_n696));
  INV_X1    g495(.A(new_n409), .ZN(new_n697));
  INV_X1    g496(.A(new_n402), .ZN(new_n698));
  AOI22_X1  g497(.A1(new_n697), .A2(new_n698), .B1(KEYINPUT35), .B2(new_n392), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n332), .A2(KEYINPUT37), .ZN(new_n700));
  NAND3_X1  g499(.A1(new_n700), .A2(new_n417), .A3(new_n335), .ZN(new_n701));
  NAND3_X1  g500(.A1(new_n701), .A2(new_n419), .A3(new_n413), .ZN(new_n702));
  AOI21_X1  g501(.A(new_n425), .B1(new_n702), .B2(KEYINPUT38), .ZN(new_n703));
  NAND4_X1  g502(.A1(new_n703), .A2(new_n283), .A3(new_n403), .A4(new_n405), .ZN(new_n704));
  NAND3_X1  g503(.A1(new_n339), .A2(new_n340), .A3(new_n277), .ZN(new_n705));
  AOI21_X1  g504(.A(KEYINPUT40), .B1(new_n437), .B2(new_n439), .ZN(new_n706));
  NOR2_X1   g505(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  AOI21_X1  g506(.A(new_n686), .B1(new_n707), .B2(new_n443), .ZN(new_n708));
  AOI21_X1  g507(.A(new_n451), .B1(new_n704), .B2(new_n708), .ZN(new_n709));
  OAI211_X1 g508(.A(KEYINPUT44), .B(new_n696), .C1(new_n699), .C2(new_n709), .ZN(new_n710));
  INV_X1    g509(.A(new_n534), .ZN(new_n711));
  NOR2_X1   g510(.A1(new_n692), .A2(new_n711), .ZN(new_n712));
  NAND2_X1  g511(.A1(new_n704), .A2(new_n708), .ZN(new_n713));
  OAI211_X1 g512(.A(new_n686), .B(KEYINPUT103), .C1(new_n661), .C2(new_n427), .ZN(new_n714));
  INV_X1    g513(.A(KEYINPUT103), .ZN(new_n715));
  OAI21_X1  g514(.A(new_n715), .B1(new_n341), .B2(new_n370), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n714), .A2(new_n716), .ZN(new_n717));
  NAND3_X1  g516(.A1(new_n713), .A2(new_n717), .A3(new_n450), .ZN(new_n718));
  AOI21_X1  g517(.A(new_n633), .B1(new_n718), .B2(new_n410), .ZN(new_n719));
  OAI211_X1 g518(.A(new_n710), .B(new_n712), .C1(new_n719), .C2(KEYINPUT44), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n283), .A2(new_n285), .ZN(new_n721));
  OAI22_X1  g520(.A1(new_n720), .A2(new_n721), .B1(new_n478), .B2(new_n477), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n695), .A2(new_n722), .ZN(G1328gat));
  NAND3_X1  g522(.A1(new_n693), .A2(new_n465), .A3(new_n427), .ZN(new_n724));
  INV_X1    g523(.A(KEYINPUT46), .ZN(new_n725));
  XNOR2_X1  g524(.A(new_n724), .B(new_n725), .ZN(new_n726));
  OAI21_X1  g525(.A(G36gat), .B1(new_n720), .B2(new_n408), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n726), .A2(new_n727), .ZN(G1329gat));
  OAI21_X1  g527(.A(G43gat), .B1(new_n720), .B2(new_n676), .ZN(new_n729));
  NOR2_X1   g528(.A1(new_n692), .A2(new_n633), .ZN(new_n730));
  NOR2_X1   g529(.A1(new_n678), .A2(G43gat), .ZN(new_n731));
  NAND4_X1  g530(.A1(new_n452), .A2(new_n534), .A3(new_n730), .A4(new_n731), .ZN(new_n732));
  INV_X1    g531(.A(KEYINPUT104), .ZN(new_n733));
  XNOR2_X1  g532(.A(new_n732), .B(new_n733), .ZN(new_n734));
  OAI21_X1  g533(.A(new_n729), .B1(new_n734), .B2(KEYINPUT105), .ZN(new_n735));
  INV_X1    g534(.A(KEYINPUT47), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  OAI21_X1  g536(.A(new_n450), .B1(new_n426), .B2(new_n445), .ZN(new_n738));
  AND2_X1   g537(.A1(new_n714), .A2(new_n716), .ZN(new_n739));
  OAI21_X1  g538(.A(new_n410), .B1(new_n738), .B2(new_n739), .ZN(new_n740));
  NAND2_X1  g539(.A1(new_n740), .A2(new_n696), .ZN(new_n741));
  INV_X1    g540(.A(KEYINPUT44), .ZN(new_n742));
  NAND2_X1  g541(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  INV_X1    g542(.A(new_n450), .ZN(new_n744));
  NAND4_X1  g543(.A1(new_n743), .A2(new_n744), .A3(new_n710), .A4(new_n712), .ZN(new_n745));
  AOI21_X1  g544(.A(new_n736), .B1(new_n745), .B2(G43gat), .ZN(new_n746));
  AND2_X1   g545(.A1(new_n736), .A2(KEYINPUT105), .ZN(new_n747));
  OAI21_X1  g546(.A(new_n734), .B1(new_n746), .B2(new_n747), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n737), .A2(new_n748), .ZN(G1330gat));
  INV_X1    g548(.A(KEYINPUT48), .ZN(new_n750));
  OAI21_X1  g549(.A(G50gat), .B1(new_n720), .B2(new_n370), .ZN(new_n751));
  INV_X1    g550(.A(KEYINPUT106), .ZN(new_n752));
  NOR2_X1   g551(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  OR2_X1    g552(.A1(new_n370), .A2(G50gat), .ZN(new_n754));
  XNOR2_X1  g553(.A(new_n754), .B(KEYINPUT107), .ZN(new_n755));
  NAND4_X1  g554(.A1(new_n452), .A2(new_n534), .A3(new_n730), .A4(new_n755), .ZN(new_n756));
  XNOR2_X1  g555(.A(new_n756), .B(KEYINPUT108), .ZN(new_n757));
  OAI21_X1  g556(.A(new_n750), .B1(new_n753), .B2(new_n757), .ZN(new_n758));
  NAND2_X1  g557(.A1(new_n756), .A2(KEYINPUT48), .ZN(new_n759));
  OAI21_X1  g558(.A(new_n759), .B1(KEYINPUT106), .B2(KEYINPUT48), .ZN(new_n760));
  NAND2_X1  g559(.A1(new_n751), .A2(new_n760), .ZN(new_n761));
  NAND2_X1  g560(.A1(new_n758), .A2(new_n761), .ZN(G1331gat));
  NOR3_X1   g561(.A1(new_n634), .A2(new_n534), .A3(new_n691), .ZN(new_n763));
  AND2_X1   g562(.A1(new_n740), .A2(new_n763), .ZN(new_n764));
  NAND2_X1  g563(.A1(new_n764), .A2(new_n661), .ZN(new_n765));
  XNOR2_X1  g564(.A(new_n765), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g565(.A1(new_n764), .A2(new_n427), .ZN(new_n767));
  NOR2_X1   g566(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n768));
  AND2_X1   g567(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n769));
  NOR3_X1   g568(.A1(new_n767), .A2(new_n768), .A3(new_n769), .ZN(new_n770));
  AOI21_X1  g569(.A(new_n770), .B1(new_n768), .B2(new_n767), .ZN(G1333gat));
  INV_X1    g570(.A(KEYINPUT50), .ZN(new_n772));
  INV_X1    g571(.A(KEYINPUT110), .ZN(new_n773));
  INV_X1    g572(.A(new_n678), .ZN(new_n774));
  AND2_X1   g573(.A1(new_n774), .A2(KEYINPUT109), .ZN(new_n775));
  NOR2_X1   g574(.A1(new_n774), .A2(KEYINPUT109), .ZN(new_n776));
  NOR2_X1   g575(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  INV_X1    g576(.A(new_n777), .ZN(new_n778));
  NAND3_X1  g577(.A1(new_n764), .A2(new_n773), .A3(new_n778), .ZN(new_n779));
  NAND2_X1  g578(.A1(new_n740), .A2(new_n763), .ZN(new_n780));
  OAI21_X1  g579(.A(KEYINPUT110), .B1(new_n780), .B2(new_n777), .ZN(new_n781));
  NAND2_X1  g580(.A1(new_n779), .A2(new_n781), .ZN(new_n782));
  INV_X1    g581(.A(G71gat), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n782), .A2(new_n783), .ZN(new_n784));
  AOI21_X1  g583(.A(new_n783), .B1(new_n764), .B2(new_n675), .ZN(new_n785));
  INV_X1    g584(.A(new_n785), .ZN(new_n786));
  AOI21_X1  g585(.A(new_n772), .B1(new_n784), .B2(new_n786), .ZN(new_n787));
  AOI211_X1 g586(.A(KEYINPUT50), .B(new_n785), .C1(new_n782), .C2(new_n783), .ZN(new_n788));
  NOR2_X1   g587(.A1(new_n787), .A2(new_n788), .ZN(G1334gat));
  NOR2_X1   g588(.A1(new_n780), .A2(new_n370), .ZN(new_n790));
  XOR2_X1   g589(.A(KEYINPUT111), .B(G78gat), .Z(new_n791));
  XNOR2_X1  g590(.A(new_n790), .B(new_n791), .ZN(G1335gat));
  NOR2_X1   g591(.A1(new_n583), .A2(new_n534), .ZN(new_n793));
  INV_X1    g592(.A(new_n793), .ZN(new_n794));
  NOR2_X1   g593(.A1(new_n794), .A2(new_n691), .ZN(new_n795));
  OAI211_X1 g594(.A(new_n710), .B(new_n795), .C1(new_n719), .C2(KEYINPUT44), .ZN(new_n796));
  OAI21_X1  g595(.A(G85gat), .B1(new_n796), .B2(new_n721), .ZN(new_n797));
  NAND3_X1  g596(.A1(new_n740), .A2(new_n696), .A3(new_n793), .ZN(new_n798));
  OR2_X1    g597(.A1(new_n798), .A2(KEYINPUT51), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n798), .A2(KEYINPUT51), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  NAND3_X1  g600(.A1(new_n661), .A2(new_n595), .A3(new_n659), .ZN(new_n802));
  OAI21_X1  g601(.A(new_n797), .B1(new_n801), .B2(new_n802), .ZN(G1336gat));
  OAI21_X1  g602(.A(G92gat), .B1(new_n796), .B2(new_n408), .ZN(new_n804));
  NAND3_X1  g603(.A1(new_n427), .A2(new_n596), .A3(new_n659), .ZN(new_n805));
  NOR2_X1   g604(.A1(KEYINPUT112), .A2(KEYINPUT51), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n798), .A2(new_n806), .ZN(new_n807));
  INV_X1    g606(.A(new_n806), .ZN(new_n808));
  NAND3_X1  g607(.A1(new_n719), .A2(new_n793), .A3(new_n808), .ZN(new_n809));
  AOI21_X1  g608(.A(new_n805), .B1(new_n807), .B2(new_n809), .ZN(new_n810));
  INV_X1    g609(.A(KEYINPUT113), .ZN(new_n811));
  OAI21_X1  g610(.A(new_n804), .B1(new_n810), .B2(new_n811), .ZN(new_n812));
  AOI211_X1 g611(.A(KEYINPUT113), .B(new_n805), .C1(new_n807), .C2(new_n809), .ZN(new_n813));
  OAI21_X1  g612(.A(KEYINPUT52), .B1(new_n812), .B2(new_n813), .ZN(new_n814));
  INV_X1    g613(.A(KEYINPUT52), .ZN(new_n815));
  OAI211_X1 g614(.A(new_n815), .B(new_n804), .C1(new_n801), .C2(new_n805), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n814), .A2(new_n816), .ZN(G1337gat));
  NOR3_X1   g616(.A1(new_n678), .A2(G99gat), .A3(new_n691), .ZN(new_n818));
  NAND3_X1  g617(.A1(new_n799), .A2(new_n800), .A3(new_n818), .ZN(new_n819));
  OAI21_X1  g618(.A(G99gat), .B1(new_n796), .B2(new_n676), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n821), .A2(KEYINPUT114), .ZN(new_n822));
  INV_X1    g621(.A(KEYINPUT114), .ZN(new_n823));
  NAND3_X1  g622(.A1(new_n819), .A2(new_n823), .A3(new_n820), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n822), .A2(new_n824), .ZN(G1338gat));
  INV_X1    g624(.A(G106gat), .ZN(new_n826));
  OR3_X1    g625(.A1(new_n796), .A2(KEYINPUT115), .A3(new_n370), .ZN(new_n827));
  NAND4_X1  g626(.A1(new_n743), .A2(new_n686), .A3(new_n710), .A4(new_n795), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n828), .A2(KEYINPUT115), .ZN(new_n829));
  AOI21_X1  g628(.A(new_n826), .B1(new_n827), .B2(new_n829), .ZN(new_n830));
  INV_X1    g629(.A(KEYINPUT53), .ZN(new_n831));
  NAND3_X1  g630(.A1(new_n686), .A2(new_n826), .A3(new_n659), .ZN(new_n832));
  OAI21_X1  g631(.A(new_n831), .B1(new_n801), .B2(new_n832), .ZN(new_n833));
  AOI21_X1  g632(.A(new_n832), .B1(new_n807), .B2(new_n809), .ZN(new_n834));
  AOI21_X1  g633(.A(new_n834), .B1(G106gat), .B2(new_n828), .ZN(new_n835));
  OAI22_X1  g634(.A1(new_n830), .A2(new_n833), .B1(new_n835), .B2(new_n831), .ZN(G1339gat));
  NAND2_X1  g635(.A1(new_n644), .A2(new_n646), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n837), .A2(new_n635), .ZN(new_n838));
  NAND3_X1  g637(.A1(new_n644), .A2(new_n646), .A3(new_n636), .ZN(new_n839));
  NAND3_X1  g638(.A1(new_n838), .A2(KEYINPUT54), .A3(new_n839), .ZN(new_n840));
  INV_X1    g639(.A(new_n650), .ZN(new_n841));
  INV_X1    g640(.A(KEYINPUT54), .ZN(new_n842));
  AOI21_X1  g641(.A(new_n841), .B1(new_n647), .B2(new_n842), .ZN(new_n843));
  AOI21_X1  g642(.A(KEYINPUT55), .B1(new_n840), .B2(new_n843), .ZN(new_n844));
  AOI21_X1  g643(.A(new_n844), .B1(new_n528), .B2(new_n533), .ZN(new_n845));
  NAND3_X1  g644(.A1(new_n840), .A2(KEYINPUT55), .A3(new_n843), .ZN(new_n846));
  AND3_X1   g645(.A1(new_n846), .A2(KEYINPUT116), .A3(new_n657), .ZN(new_n847));
  AOI21_X1  g646(.A(KEYINPUT116), .B1(new_n846), .B2(new_n657), .ZN(new_n848));
  OAI21_X1  g647(.A(new_n845), .B1(new_n847), .B2(new_n848), .ZN(new_n849));
  NAND2_X1  g648(.A1(new_n503), .A2(new_n487), .ZN(new_n850));
  INV_X1    g649(.A(new_n850), .ZN(new_n851));
  OAI22_X1  g650(.A1(new_n851), .A2(new_n488), .B1(new_n508), .B2(new_n509), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n523), .A2(new_n524), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  NAND3_X1  g653(.A1(new_n659), .A2(new_n528), .A3(new_n854), .ZN(new_n855));
  AOI21_X1  g654(.A(new_n696), .B1(new_n849), .B2(new_n855), .ZN(new_n856));
  AND3_X1   g655(.A1(new_n495), .A2(KEYINPUT91), .A3(new_n496), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n504), .A2(new_n527), .ZN(new_n858));
  NOR2_X1   g657(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  AOI22_X1  g658(.A1(new_n859), .A2(new_n499), .B1(new_n853), .B2(new_n852), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n840), .A2(new_n843), .ZN(new_n861));
  INV_X1    g660(.A(KEYINPUT55), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  NAND4_X1  g662(.A1(new_n860), .A2(new_n631), .A3(new_n632), .A4(new_n863), .ZN(new_n864));
  NOR2_X1   g663(.A1(new_n847), .A2(new_n848), .ZN(new_n865));
  NOR2_X1   g664(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  OAI21_X1  g665(.A(new_n690), .B1(new_n856), .B2(new_n866), .ZN(new_n867));
  NAND4_X1  g666(.A1(new_n583), .A2(new_n711), .A3(new_n633), .A4(new_n691), .ZN(new_n868));
  NAND2_X1  g667(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  NOR2_X1   g668(.A1(new_n721), .A2(new_n427), .ZN(new_n870));
  AND2_X1   g669(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  NAND3_X1  g670(.A1(new_n871), .A2(new_n370), .A3(new_n391), .ZN(new_n872));
  INV_X1    g671(.A(new_n213), .ZN(new_n873));
  NOR3_X1   g672(.A1(new_n872), .A2(new_n873), .A3(new_n711), .ZN(new_n874));
  NAND3_X1  g673(.A1(new_n871), .A2(new_n534), .A3(new_n698), .ZN(new_n875));
  AOI21_X1  g674(.A(new_n874), .B1(new_n875), .B2(G113gat), .ZN(new_n876));
  XOR2_X1   g675(.A(new_n876), .B(KEYINPUT117), .Z(G1340gat));
  NAND2_X1  g676(.A1(new_n871), .A2(new_n698), .ZN(new_n878));
  OAI21_X1  g677(.A(G120gat), .B1(new_n878), .B2(new_n691), .ZN(new_n879));
  NAND2_X1  g678(.A1(new_n659), .A2(new_n220), .ZN(new_n880));
  XNOR2_X1  g679(.A(new_n880), .B(KEYINPUT118), .ZN(new_n881));
  OAI21_X1  g680(.A(new_n879), .B1(new_n872), .B2(new_n881), .ZN(G1341gat));
  OAI21_X1  g681(.A(G127gat), .B1(new_n878), .B2(new_n690), .ZN(new_n883));
  OR2_X1    g682(.A1(new_n690), .A2(G127gat), .ZN(new_n884));
  OAI21_X1  g683(.A(new_n883), .B1(new_n872), .B2(new_n884), .ZN(G1342gat));
  NAND2_X1  g684(.A1(new_n370), .A2(new_n391), .ZN(new_n886));
  NOR3_X1   g685(.A1(new_n886), .A2(G134gat), .A3(new_n633), .ZN(new_n887));
  NAND2_X1  g686(.A1(new_n871), .A2(new_n887), .ZN(new_n888));
  XOR2_X1   g687(.A(new_n888), .B(KEYINPUT56), .Z(new_n889));
  OAI21_X1  g688(.A(G134gat), .B1(new_n878), .B2(new_n633), .ZN(new_n890));
  NAND2_X1  g689(.A1(new_n889), .A2(new_n890), .ZN(G1343gat));
  NOR2_X1   g690(.A1(new_n675), .A2(new_n370), .ZN(new_n892));
  AND2_X1   g691(.A1(new_n892), .A2(new_n871), .ZN(new_n893));
  NAND3_X1  g692(.A1(new_n893), .A2(new_n234), .A3(new_n534), .ZN(new_n894));
  NAND4_X1  g693(.A1(new_n534), .A2(new_n657), .A3(new_n863), .A4(new_n846), .ZN(new_n895));
  AOI22_X1  g694(.A1(new_n895), .A2(new_n855), .B1(new_n632), .B2(new_n631), .ZN(new_n896));
  OAI21_X1  g695(.A(new_n690), .B1(new_n896), .B2(new_n866), .ZN(new_n897));
  NAND2_X1  g696(.A1(new_n897), .A2(new_n868), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n898), .A2(new_n686), .ZN(new_n899));
  NAND2_X1  g698(.A1(new_n899), .A2(KEYINPUT57), .ZN(new_n900));
  NAND2_X1  g699(.A1(new_n870), .A2(new_n450), .ZN(new_n901));
  INV_X1    g700(.A(new_n901), .ZN(new_n902));
  INV_X1    g701(.A(KEYINPUT57), .ZN(new_n903));
  NAND3_X1  g702(.A1(new_n869), .A2(new_n903), .A3(new_n686), .ZN(new_n904));
  NAND3_X1  g703(.A1(new_n900), .A2(new_n902), .A3(new_n904), .ZN(new_n905));
  OAI21_X1  g704(.A(G141gat), .B1(new_n905), .B2(new_n711), .ZN(new_n906));
  NAND2_X1  g705(.A1(new_n894), .A2(new_n906), .ZN(new_n907));
  XNOR2_X1  g706(.A(new_n907), .B(KEYINPUT58), .ZN(G1344gat));
  NAND3_X1  g707(.A1(new_n893), .A2(new_n232), .A3(new_n659), .ZN(new_n909));
  INV_X1    g708(.A(KEYINPUT121), .ZN(new_n910));
  AOI211_X1 g709(.A(new_n903), .B(new_n370), .C1(new_n867), .C2(new_n868), .ZN(new_n911));
  INV_X1    g710(.A(KEYINPUT120), .ZN(new_n912));
  AOI21_X1  g711(.A(KEYINPUT91), .B1(new_n495), .B2(new_n496), .ZN(new_n913));
  NOR3_X1   g712(.A1(new_n857), .A2(new_n858), .A3(new_n913), .ZN(new_n914));
  AOI22_X1  g713(.A1(new_n495), .A2(new_n496), .B1(new_n508), .B2(new_n509), .ZN(new_n915));
  AOI21_X1  g714(.A(new_n531), .B1(new_n915), .B2(new_n504), .ZN(new_n916));
  OAI21_X1  g715(.A(new_n863), .B1(new_n914), .B2(new_n916), .ZN(new_n917));
  NAND2_X1  g716(.A1(new_n846), .A2(new_n657), .ZN(new_n918));
  OAI21_X1  g717(.A(new_n855), .B1(new_n917), .B2(new_n918), .ZN(new_n919));
  NAND2_X1  g718(.A1(new_n919), .A2(new_n633), .ZN(new_n920));
  INV_X1    g719(.A(KEYINPUT116), .ZN(new_n921));
  NAND2_X1  g720(.A1(new_n918), .A2(new_n921), .ZN(new_n922));
  NAND3_X1  g721(.A1(new_n846), .A2(KEYINPUT116), .A3(new_n657), .ZN(new_n923));
  NAND2_X1  g722(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  AND3_X1   g723(.A1(new_n863), .A2(new_n528), .A3(new_n854), .ZN(new_n925));
  NAND3_X1  g724(.A1(new_n696), .A2(new_n924), .A3(new_n925), .ZN(new_n926));
  AOI21_X1  g725(.A(new_n583), .B1(new_n920), .B2(new_n926), .ZN(new_n927));
  INV_X1    g726(.A(new_n868), .ZN(new_n928));
  OAI21_X1  g727(.A(new_n912), .B1(new_n927), .B2(new_n928), .ZN(new_n929));
  NAND3_X1  g728(.A1(new_n897), .A2(KEYINPUT120), .A3(new_n868), .ZN(new_n930));
  NAND3_X1  g729(.A1(new_n929), .A2(new_n930), .A3(new_n686), .ZN(new_n931));
  AOI21_X1  g730(.A(new_n911), .B1(new_n931), .B2(new_n903), .ZN(new_n932));
  NOR3_X1   g731(.A1(new_n932), .A2(new_n691), .A3(new_n901), .ZN(new_n933));
  OAI211_X1 g732(.A(new_n910), .B(KEYINPUT59), .C1(new_n933), .C2(new_n232), .ZN(new_n934));
  NAND4_X1  g733(.A1(new_n900), .A2(new_n659), .A3(new_n904), .A4(new_n902), .ZN(new_n935));
  NOR2_X1   g734(.A1(new_n232), .A2(KEYINPUT59), .ZN(new_n936));
  AND3_X1   g735(.A1(new_n935), .A2(KEYINPUT119), .A3(new_n936), .ZN(new_n937));
  AOI21_X1  g736(.A(KEYINPUT119), .B1(new_n935), .B2(new_n936), .ZN(new_n938));
  NOR2_X1   g737(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  NAND2_X1  g738(.A1(new_n934), .A2(new_n939), .ZN(new_n940));
  AOI21_X1  g739(.A(new_n370), .B1(new_n898), .B2(new_n912), .ZN(new_n941));
  AOI21_X1  g740(.A(KEYINPUT57), .B1(new_n941), .B2(new_n930), .ZN(new_n942));
  OAI211_X1 g741(.A(new_n659), .B(new_n902), .C1(new_n942), .C2(new_n911), .ZN(new_n943));
  NAND2_X1  g742(.A1(new_n943), .A2(G148gat), .ZN(new_n944));
  AOI21_X1  g743(.A(new_n910), .B1(new_n944), .B2(KEYINPUT59), .ZN(new_n945));
  OAI21_X1  g744(.A(new_n909), .B1(new_n940), .B2(new_n945), .ZN(new_n946));
  NAND2_X1  g745(.A1(new_n946), .A2(KEYINPUT122), .ZN(new_n947));
  INV_X1    g746(.A(KEYINPUT122), .ZN(new_n948));
  OAI211_X1 g747(.A(new_n948), .B(new_n909), .C1(new_n940), .C2(new_n945), .ZN(new_n949));
  NAND2_X1  g748(.A1(new_n947), .A2(new_n949), .ZN(G1345gat));
  NAND3_X1  g749(.A1(new_n893), .A2(new_n238), .A3(new_n583), .ZN(new_n951));
  OAI21_X1  g750(.A(G155gat), .B1(new_n905), .B2(new_n690), .ZN(new_n952));
  NAND2_X1  g751(.A1(new_n951), .A2(new_n952), .ZN(G1346gat));
  NAND3_X1  g752(.A1(new_n893), .A2(new_n239), .A3(new_n696), .ZN(new_n954));
  OAI21_X1  g753(.A(G162gat), .B1(new_n905), .B2(new_n633), .ZN(new_n955));
  NAND2_X1  g754(.A1(new_n954), .A2(new_n955), .ZN(G1347gat));
  NOR2_X1   g755(.A1(new_n661), .A2(new_n408), .ZN(new_n957));
  AND2_X1   g756(.A1(new_n869), .A2(new_n957), .ZN(new_n958));
  INV_X1    g757(.A(new_n958), .ZN(new_n959));
  NOR2_X1   g758(.A1(new_n959), .A2(new_n886), .ZN(new_n960));
  AOI21_X1  g759(.A(G169gat), .B1(new_n960), .B2(new_n534), .ZN(new_n961));
  NOR3_X1   g760(.A1(new_n777), .A2(new_n959), .A3(new_n686), .ZN(new_n962));
  NOR2_X1   g761(.A1(new_n711), .A2(new_n290), .ZN(new_n963));
  AOI21_X1  g762(.A(new_n961), .B1(new_n962), .B2(new_n963), .ZN(new_n964));
  XOR2_X1   g763(.A(new_n964), .B(KEYINPUT123), .Z(G1348gat));
  INV_X1    g764(.A(new_n962), .ZN(new_n966));
  NOR3_X1   g765(.A1(new_n966), .A2(new_n291), .A3(new_n691), .ZN(new_n967));
  AOI21_X1  g766(.A(G176gat), .B1(new_n960), .B2(new_n659), .ZN(new_n968));
  INV_X1    g767(.A(KEYINPUT124), .ZN(new_n969));
  AND2_X1   g768(.A1(new_n968), .A2(new_n969), .ZN(new_n970));
  NOR2_X1   g769(.A1(new_n968), .A2(new_n969), .ZN(new_n971));
  NOR3_X1   g770(.A1(new_n967), .A2(new_n970), .A3(new_n971), .ZN(G1349gat));
  OAI21_X1  g771(.A(G183gat), .B1(new_n966), .B2(new_n690), .ZN(new_n973));
  NAND3_X1  g772(.A1(new_n960), .A2(new_n297), .A3(new_n583), .ZN(new_n974));
  NAND2_X1  g773(.A1(new_n973), .A2(new_n974), .ZN(new_n975));
  XNOR2_X1  g774(.A(KEYINPUT125), .B(KEYINPUT60), .ZN(new_n976));
  XNOR2_X1  g775(.A(new_n975), .B(new_n976), .ZN(G1350gat));
  OAI21_X1  g776(.A(G190gat), .B1(new_n966), .B2(new_n633), .ZN(new_n978));
  XNOR2_X1  g777(.A(KEYINPUT126), .B(KEYINPUT61), .ZN(new_n979));
  OR2_X1    g778(.A1(new_n978), .A2(new_n979), .ZN(new_n980));
  NAND2_X1  g779(.A1(new_n978), .A2(new_n979), .ZN(new_n981));
  NAND3_X1  g780(.A1(new_n960), .A2(new_n298), .A3(new_n696), .ZN(new_n982));
  NAND3_X1  g781(.A1(new_n980), .A2(new_n981), .A3(new_n982), .ZN(G1351gat));
  NAND2_X1  g782(.A1(new_n892), .A2(new_n958), .ZN(new_n984));
  INV_X1    g783(.A(new_n984), .ZN(new_n985));
  AOI21_X1  g784(.A(G197gat), .B1(new_n985), .B2(new_n534), .ZN(new_n986));
  NOR3_X1   g785(.A1(new_n675), .A2(new_n661), .A3(new_n408), .ZN(new_n987));
  INV_X1    g786(.A(new_n987), .ZN(new_n988));
  NOR2_X1   g787(.A1(new_n988), .A2(new_n932), .ZN(new_n989));
  NOR2_X1   g788(.A1(new_n711), .A2(new_n516), .ZN(new_n990));
  AOI21_X1  g789(.A(new_n986), .B1(new_n989), .B2(new_n990), .ZN(G1352gat));
  INV_X1    g790(.A(G204gat), .ZN(new_n992));
  NAND3_X1  g791(.A1(new_n985), .A2(new_n992), .A3(new_n659), .ZN(new_n993));
  NAND2_X1  g792(.A1(new_n993), .A2(KEYINPUT62), .ZN(new_n994));
  INV_X1    g793(.A(KEYINPUT127), .ZN(new_n995));
  NAND2_X1  g794(.A1(new_n994), .A2(new_n995), .ZN(new_n996));
  NAND3_X1  g795(.A1(new_n993), .A2(KEYINPUT127), .A3(KEYINPUT62), .ZN(new_n997));
  NAND2_X1  g796(.A1(new_n996), .A2(new_n997), .ZN(new_n998));
  NOR3_X1   g797(.A1(new_n988), .A2(new_n691), .A3(new_n932), .ZN(new_n999));
  OAI221_X1 g798(.A(new_n998), .B1(KEYINPUT62), .B2(new_n993), .C1(new_n992), .C2(new_n999), .ZN(G1353gat));
  NAND3_X1  g799(.A1(new_n985), .A2(new_n316), .A3(new_n583), .ZN(new_n1001));
  NAND2_X1  g800(.A1(new_n989), .A2(new_n583), .ZN(new_n1002));
  AND3_X1   g801(.A1(new_n1002), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n1003));
  AOI21_X1  g802(.A(KEYINPUT63), .B1(new_n1002), .B2(G211gat), .ZN(new_n1004));
  OAI21_X1  g803(.A(new_n1001), .B1(new_n1003), .B2(new_n1004), .ZN(G1354gat));
  NAND3_X1  g804(.A1(new_n985), .A2(new_n317), .A3(new_n696), .ZN(new_n1006));
  NOR3_X1   g805(.A1(new_n988), .A2(new_n633), .A3(new_n932), .ZN(new_n1007));
  OAI21_X1  g806(.A(new_n1006), .B1(new_n1007), .B2(new_n317), .ZN(G1355gat));
endmodule


