//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 1 1 0 1 1 1 1 1 1 1 0 0 0 0 0 0 0 0 0 0 0 1 0 0 0 1 0 1 1 0 1 1 1 0 0 0 0 1 1 1 0 1 0 0 0 1 1 1 0 0 1 1 0 0 0 1 1 1 0 0 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:30:34 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n443, new_n448, new_n449, new_n451, new_n453, new_n455,
    new_n456, new_n457, new_n460, new_n461, new_n462, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n532, new_n533,
    new_n534, new_n535, new_n536, new_n537, new_n538, new_n539, new_n540,
    new_n541, new_n542, new_n543, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n552, new_n553, new_n554, new_n555, new_n556,
    new_n557, new_n559, new_n561, new_n562, new_n563, new_n565, new_n566,
    new_n567, new_n568, new_n569, new_n570, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n580, new_n581, new_n582, new_n583, new_n584,
    new_n585, new_n586, new_n587, new_n588, new_n589, new_n590, new_n591,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n623,
    new_n624, new_n627, new_n629, new_n630, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n827, new_n828, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1144, new_n1145;
  BUF_X1    g000(.A(G452), .Z(G350));
  XOR2_X1   g001(.A(KEYINPUT64), .B(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  XOR2_X1   g006(.A(KEYINPUT65), .B(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  XOR2_X1   g016(.A(KEYINPUT66), .B(G108), .Z(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(new_n443));
  XNOR2_X1  g018(.A(new_n443), .B(KEYINPUT67), .ZN(G158));
  NAND3_X1  g019(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g020(.A(G452), .Z(G391));
  AND2_X1   g021(.A1(G94), .A2(G452), .ZN(G173));
  XNOR2_X1  g022(.A(KEYINPUT68), .B(KEYINPUT1), .ZN(new_n448));
  NAND2_X1  g023(.A1(G7), .A2(G661), .ZN(new_n449));
  XNOR2_X1  g024(.A(new_n448), .B(new_n449), .ZN(G223));
  INV_X1    g025(.A(new_n449), .ZN(new_n451));
  NAND2_X1  g026(.A1(new_n451), .A2(G567), .ZN(G234));
  NAND2_X1  g027(.A1(new_n451), .A2(G2106), .ZN(new_n453));
  XNOR2_X1  g028(.A(new_n453), .B(KEYINPUT69), .ZN(G217));
  NAND4_X1  g029(.A1(new_n436), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n455));
  XOR2_X1   g030(.A(new_n455), .B(KEYINPUT2), .Z(new_n456));
  NOR4_X1   g031(.A1(G238), .A2(G237), .A3(G235), .A4(G236), .ZN(new_n457));
  NAND2_X1  g032(.A1(new_n456), .A2(new_n457), .ZN(G261));
  INV_X1    g033(.A(G261), .ZN(G325));
  INV_X1    g034(.A(G2106), .ZN(new_n460));
  INV_X1    g035(.A(G567), .ZN(new_n461));
  OAI22_X1  g036(.A1(new_n456), .A2(new_n460), .B1(new_n461), .B2(new_n457), .ZN(new_n462));
  XOR2_X1   g037(.A(new_n462), .B(KEYINPUT70), .Z(G319));
  NAND2_X1  g038(.A1(KEYINPUT71), .A2(KEYINPUT3), .ZN(new_n464));
  NAND3_X1  g039(.A1(new_n464), .A2(KEYINPUT72), .A3(G2104), .ZN(new_n465));
  NAND2_X1  g040(.A1(KEYINPUT72), .A2(G2104), .ZN(new_n466));
  NAND3_X1  g041(.A1(new_n466), .A2(KEYINPUT71), .A3(KEYINPUT3), .ZN(new_n467));
  INV_X1    g042(.A(KEYINPUT71), .ZN(new_n468));
  INV_X1    g043(.A(KEYINPUT3), .ZN(new_n469));
  OAI21_X1  g044(.A(new_n468), .B1(new_n469), .B2(G2104), .ZN(new_n470));
  INV_X1    g045(.A(G2105), .ZN(new_n471));
  NAND4_X1  g046(.A1(new_n465), .A2(new_n467), .A3(new_n470), .A4(new_n471), .ZN(new_n472));
  INV_X1    g047(.A(G137), .ZN(new_n473));
  INV_X1    g048(.A(G101), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n471), .A2(G2104), .ZN(new_n475));
  OAI22_X1  g050(.A1(new_n472), .A2(new_n473), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  INV_X1    g051(.A(KEYINPUT73), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  OAI221_X1 g053(.A(KEYINPUT73), .B1(new_n474), .B2(new_n475), .C1(new_n472), .C2(new_n473), .ZN(new_n479));
  NAND2_X1  g054(.A1(G113), .A2(G2104), .ZN(new_n480));
  XOR2_X1   g055(.A(KEYINPUT3), .B(G2104), .Z(new_n481));
  INV_X1    g056(.A(G125), .ZN(new_n482));
  OAI21_X1  g057(.A(new_n480), .B1(new_n481), .B2(new_n482), .ZN(new_n483));
  AOI22_X1  g058(.A1(new_n478), .A2(new_n479), .B1(G2105), .B2(new_n483), .ZN(G160));
  INV_X1    g059(.A(G136), .ZN(new_n485));
  OAI21_X1  g060(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n486));
  NOR2_X1   g061(.A1(new_n471), .A2(G112), .ZN(new_n487));
  OAI22_X1  g062(.A1(new_n472), .A2(new_n485), .B1(new_n486), .B2(new_n487), .ZN(new_n488));
  AND4_X1   g063(.A1(G2105), .A2(new_n465), .A3(new_n467), .A4(new_n470), .ZN(new_n489));
  AOI21_X1  g064(.A(new_n488), .B1(new_n489), .B2(G124), .ZN(G162));
  INV_X1    g065(.A(G138), .ZN(new_n491));
  OAI21_X1  g066(.A(KEYINPUT4), .B1(new_n472), .B2(new_n491), .ZN(new_n492));
  INV_X1    g067(.A(KEYINPUT74), .ZN(new_n493));
  NAND2_X1  g068(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  OAI211_X1 g069(.A(KEYINPUT74), .B(KEYINPUT4), .C1(new_n472), .C2(new_n491), .ZN(new_n495));
  NOR2_X1   g070(.A1(new_n481), .A2(KEYINPUT4), .ZN(new_n496));
  NAND3_X1  g071(.A1(new_n496), .A2(G138), .A3(new_n471), .ZN(new_n497));
  NAND3_X1  g072(.A1(new_n494), .A2(new_n495), .A3(new_n497), .ZN(new_n498));
  OAI21_X1  g073(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n499));
  INV_X1    g074(.A(G114), .ZN(new_n500));
  AOI21_X1  g075(.A(new_n499), .B1(new_n500), .B2(G2105), .ZN(new_n501));
  AOI21_X1  g076(.A(new_n501), .B1(new_n489), .B2(G126), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n498), .A2(new_n502), .ZN(new_n503));
  INV_X1    g078(.A(new_n503), .ZN(G164));
  INV_X1    g079(.A(G543), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n505), .A2(KEYINPUT5), .ZN(new_n506));
  INV_X1    g081(.A(KEYINPUT5), .ZN(new_n507));
  NAND2_X1  g082(.A1(new_n507), .A2(G543), .ZN(new_n508));
  AND2_X1   g083(.A1(new_n506), .A2(new_n508), .ZN(new_n509));
  XNOR2_X1  g084(.A(KEYINPUT6), .B(G651), .ZN(new_n510));
  INV_X1    g085(.A(KEYINPUT75), .ZN(new_n511));
  NAND3_X1  g086(.A1(new_n509), .A2(new_n510), .A3(new_n511), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n506), .A2(new_n508), .ZN(new_n513));
  INV_X1    g088(.A(G651), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n514), .A2(KEYINPUT6), .ZN(new_n515));
  INV_X1    g090(.A(KEYINPUT6), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n516), .A2(G651), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n515), .A2(new_n517), .ZN(new_n518));
  OAI21_X1  g093(.A(KEYINPUT75), .B1(new_n513), .B2(new_n518), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n512), .A2(new_n519), .ZN(new_n520));
  INV_X1    g095(.A(new_n520), .ZN(new_n521));
  XOR2_X1   g096(.A(KEYINPUT76), .B(G88), .Z(new_n522));
  NAND2_X1  g097(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  AND2_X1   g098(.A1(new_n509), .A2(G62), .ZN(new_n524));
  NAND2_X1  g099(.A1(G75), .A2(G543), .ZN(new_n525));
  XNOR2_X1  g100(.A(new_n525), .B(KEYINPUT77), .ZN(new_n526));
  OAI21_X1  g101(.A(G651), .B1(new_n524), .B2(new_n526), .ZN(new_n527));
  NOR2_X1   g102(.A1(new_n518), .A2(new_n505), .ZN(new_n528));
  NAND2_X1  g103(.A1(new_n528), .A2(G50), .ZN(new_n529));
  NAND3_X1  g104(.A1(new_n523), .A2(new_n527), .A3(new_n529), .ZN(G303));
  INV_X1    g105(.A(G303), .ZN(G166));
  NAND3_X1  g106(.A1(new_n509), .A2(G63), .A3(G651), .ZN(new_n532));
  INV_X1    g107(.A(KEYINPUT78), .ZN(new_n533));
  XNOR2_X1  g108(.A(new_n532), .B(new_n533), .ZN(new_n534));
  NAND3_X1  g109(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n535));
  XNOR2_X1  g110(.A(new_n535), .B(KEYINPUT7), .ZN(new_n536));
  INV_X1    g111(.A(KEYINPUT79), .ZN(new_n537));
  NAND2_X1  g112(.A1(new_n518), .A2(new_n537), .ZN(new_n538));
  NAND2_X1  g113(.A1(new_n510), .A2(KEYINPUT79), .ZN(new_n539));
  AND3_X1   g114(.A1(new_n538), .A2(new_n539), .A3(G543), .ZN(new_n540));
  NAND2_X1  g115(.A1(new_n540), .A2(G51), .ZN(new_n541));
  NAND3_X1  g116(.A1(new_n534), .A2(new_n536), .A3(new_n541), .ZN(new_n542));
  AND2_X1   g117(.A1(new_n521), .A2(G89), .ZN(new_n543));
  NOR2_X1   g118(.A1(new_n542), .A2(new_n543), .ZN(G168));
  AOI22_X1  g119(.A1(new_n509), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n545));
  OR2_X1    g120(.A1(new_n545), .A2(new_n514), .ZN(new_n546));
  NAND3_X1  g121(.A1(new_n538), .A2(new_n539), .A3(G543), .ZN(new_n547));
  INV_X1    g122(.A(G52), .ZN(new_n548));
  OAI21_X1  g123(.A(new_n546), .B1(new_n547), .B2(new_n548), .ZN(new_n549));
  AND2_X1   g124(.A1(new_n521), .A2(G90), .ZN(new_n550));
  NOR2_X1   g125(.A1(new_n549), .A2(new_n550), .ZN(G171));
  AOI22_X1  g126(.A1(new_n509), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n552));
  OR2_X1    g127(.A1(new_n552), .A2(new_n514), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n540), .A2(G43), .ZN(new_n554));
  INV_X1    g129(.A(G81), .ZN(new_n555));
  OAI211_X1 g130(.A(new_n553), .B(new_n554), .C1(new_n555), .C2(new_n520), .ZN(new_n556));
  INV_X1    g131(.A(new_n556), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n557), .A2(G860), .ZN(G153));
  AND3_X1   g133(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n559), .A2(G36), .ZN(G176));
  XOR2_X1   g135(.A(KEYINPUT80), .B(KEYINPUT8), .Z(new_n561));
  NAND2_X1  g136(.A1(G1), .A2(G3), .ZN(new_n562));
  XNOR2_X1  g137(.A(new_n561), .B(new_n562), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n559), .A2(new_n563), .ZN(G188));
  NAND2_X1  g139(.A1(new_n540), .A2(G53), .ZN(new_n565));
  XNOR2_X1  g140(.A(new_n565), .B(KEYINPUT9), .ZN(new_n566));
  AOI22_X1  g141(.A1(new_n509), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n567));
  XNOR2_X1  g142(.A(new_n567), .B(KEYINPUT81), .ZN(new_n568));
  NAND2_X1  g143(.A1(new_n568), .A2(G651), .ZN(new_n569));
  NAND2_X1  g144(.A1(new_n521), .A2(G91), .ZN(new_n570));
  NAND3_X1  g145(.A1(new_n566), .A2(new_n569), .A3(new_n570), .ZN(G299));
  OR2_X1    g146(.A1(new_n549), .A2(new_n550), .ZN(G301));
  INV_X1    g147(.A(G168), .ZN(G286));
  INV_X1    g148(.A(G87), .ZN(new_n574));
  OR3_X1    g149(.A1(new_n520), .A2(KEYINPUT82), .A3(new_n574), .ZN(new_n575));
  OR2_X1    g150(.A1(new_n509), .A2(G74), .ZN(new_n576));
  AOI22_X1  g151(.A1(new_n540), .A2(G49), .B1(G651), .B2(new_n576), .ZN(new_n577));
  OAI21_X1  g152(.A(KEYINPUT82), .B1(new_n520), .B2(new_n574), .ZN(new_n578));
  NAND3_X1  g153(.A1(new_n575), .A2(new_n577), .A3(new_n578), .ZN(G288));
  INV_X1    g154(.A(G61), .ZN(new_n580));
  OR3_X1    g155(.A1(new_n513), .A2(KEYINPUT83), .A3(new_n580), .ZN(new_n581));
  NAND2_X1  g156(.A1(G73), .A2(G543), .ZN(new_n582));
  XOR2_X1   g157(.A(new_n582), .B(KEYINPUT84), .Z(new_n583));
  OAI21_X1  g158(.A(KEYINPUT83), .B1(new_n513), .B2(new_n580), .ZN(new_n584));
  NAND3_X1  g159(.A1(new_n581), .A2(new_n583), .A3(new_n584), .ZN(new_n585));
  NAND2_X1  g160(.A1(new_n585), .A2(G651), .ZN(new_n586));
  XNOR2_X1  g161(.A(new_n586), .B(KEYINPUT85), .ZN(new_n587));
  NAND2_X1  g162(.A1(new_n528), .A2(G48), .ZN(new_n588));
  INV_X1    g163(.A(G86), .ZN(new_n589));
  OAI21_X1  g164(.A(new_n588), .B1(new_n520), .B2(new_n589), .ZN(new_n590));
  NOR2_X1   g165(.A1(new_n587), .A2(new_n590), .ZN(new_n591));
  INV_X1    g166(.A(new_n591), .ZN(G305));
  AOI22_X1  g167(.A1(new_n509), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n593));
  OR2_X1    g168(.A1(new_n593), .A2(new_n514), .ZN(new_n594));
  INV_X1    g169(.A(G85), .ZN(new_n595));
  INV_X1    g170(.A(G47), .ZN(new_n596));
  OAI22_X1  g171(.A1(new_n520), .A2(new_n595), .B1(new_n547), .B2(new_n596), .ZN(new_n597));
  AND2_X1   g172(.A1(new_n597), .A2(KEYINPUT86), .ZN(new_n598));
  NOR2_X1   g173(.A1(new_n597), .A2(KEYINPUT86), .ZN(new_n599));
  OAI21_X1  g174(.A(new_n594), .B1(new_n598), .B2(new_n599), .ZN(G290));
  NAND2_X1  g175(.A1(G301), .A2(G868), .ZN(new_n601));
  INV_X1    g176(.A(G92), .ZN(new_n602));
  OR3_X1    g177(.A1(new_n520), .A2(KEYINPUT88), .A3(new_n602), .ZN(new_n603));
  OAI21_X1  g178(.A(KEYINPUT88), .B1(new_n520), .B2(new_n602), .ZN(new_n604));
  NAND2_X1  g179(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  NAND2_X1  g180(.A1(new_n605), .A2(KEYINPUT87), .ZN(new_n606));
  INV_X1    g181(.A(KEYINPUT87), .ZN(new_n607));
  NAND3_X1  g182(.A1(new_n603), .A2(new_n607), .A3(new_n604), .ZN(new_n608));
  NAND2_X1  g183(.A1(new_n606), .A2(new_n608), .ZN(new_n609));
  INV_X1    g184(.A(KEYINPUT10), .ZN(new_n610));
  NAND2_X1  g185(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  OR2_X1    g186(.A1(KEYINPUT89), .A2(G66), .ZN(new_n612));
  NAND2_X1  g187(.A1(KEYINPUT89), .A2(G66), .ZN(new_n613));
  NAND3_X1  g188(.A1(new_n509), .A2(new_n612), .A3(new_n613), .ZN(new_n614));
  NAND2_X1  g189(.A1(G79), .A2(G543), .ZN(new_n615));
  AOI21_X1  g190(.A(new_n514), .B1(new_n614), .B2(new_n615), .ZN(new_n616));
  AOI21_X1  g191(.A(new_n616), .B1(G54), .B2(new_n540), .ZN(new_n617));
  NAND3_X1  g192(.A1(new_n606), .A2(KEYINPUT10), .A3(new_n608), .ZN(new_n618));
  NAND3_X1  g193(.A1(new_n611), .A2(new_n617), .A3(new_n618), .ZN(new_n619));
  XNOR2_X1  g194(.A(new_n619), .B(KEYINPUT90), .ZN(new_n620));
  OAI21_X1  g195(.A(new_n601), .B1(new_n620), .B2(G868), .ZN(G284));
  OAI21_X1  g196(.A(new_n601), .B1(new_n620), .B2(G868), .ZN(G321));
  NAND2_X1  g197(.A1(G286), .A2(G868), .ZN(new_n623));
  INV_X1    g198(.A(G299), .ZN(new_n624));
  OAI21_X1  g199(.A(new_n623), .B1(new_n624), .B2(G868), .ZN(G297));
  OAI21_X1  g200(.A(new_n623), .B1(new_n624), .B2(G868), .ZN(G280));
  INV_X1    g201(.A(G559), .ZN(new_n627));
  OAI21_X1  g202(.A(new_n620), .B1(new_n627), .B2(G860), .ZN(G148));
  NAND2_X1  g203(.A1(new_n620), .A2(new_n627), .ZN(new_n629));
  NAND2_X1  g204(.A1(new_n629), .A2(G868), .ZN(new_n630));
  OAI21_X1  g205(.A(new_n630), .B1(G868), .B2(new_n557), .ZN(G323));
  XNOR2_X1  g206(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NOR2_X1   g207(.A1(new_n481), .A2(new_n475), .ZN(new_n633));
  XOR2_X1   g208(.A(new_n633), .B(KEYINPUT12), .Z(new_n634));
  XOR2_X1   g209(.A(new_n634), .B(KEYINPUT13), .Z(new_n635));
  INV_X1    g210(.A(KEYINPUT91), .ZN(new_n636));
  NOR2_X1   g211(.A1(new_n636), .A2(G2100), .ZN(new_n637));
  XNOR2_X1  g212(.A(new_n635), .B(new_n637), .ZN(new_n638));
  INV_X1    g213(.A(G135), .ZN(new_n639));
  OAI21_X1  g214(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n640));
  NOR2_X1   g215(.A1(new_n471), .A2(G111), .ZN(new_n641));
  OAI22_X1  g216(.A1(new_n472), .A2(new_n639), .B1(new_n640), .B2(new_n641), .ZN(new_n642));
  AOI21_X1  g217(.A(new_n642), .B1(new_n489), .B2(G123), .ZN(new_n643));
  INV_X1    g218(.A(G2096), .ZN(new_n644));
  AOI22_X1  g219(.A1(new_n643), .A2(new_n644), .B1(new_n636), .B2(G2100), .ZN(new_n645));
  OAI211_X1 g220(.A(new_n638), .B(new_n645), .C1(new_n644), .C2(new_n643), .ZN(G156));
  XNOR2_X1  g221(.A(G2427), .B(G2438), .ZN(new_n647));
  XNOR2_X1  g222(.A(new_n647), .B(G2430), .ZN(new_n648));
  XNOR2_X1  g223(.A(new_n648), .B(KEYINPUT15), .ZN(new_n649));
  XOR2_X1   g224(.A(new_n649), .B(G2435), .Z(new_n650));
  NAND2_X1  g225(.A1(new_n650), .A2(KEYINPUT14), .ZN(new_n651));
  XOR2_X1   g226(.A(KEYINPUT92), .B(KEYINPUT16), .Z(new_n652));
  XNOR2_X1  g227(.A(new_n651), .B(new_n652), .ZN(new_n653));
  XNOR2_X1  g228(.A(G2443), .B(G2446), .ZN(new_n654));
  XNOR2_X1  g229(.A(G2451), .B(G2454), .ZN(new_n655));
  XNOR2_X1  g230(.A(new_n654), .B(new_n655), .ZN(new_n656));
  XNOR2_X1  g231(.A(new_n653), .B(new_n656), .ZN(new_n657));
  XNOR2_X1  g232(.A(G1341), .B(G1348), .ZN(new_n658));
  XOR2_X1   g233(.A(new_n657), .B(new_n658), .Z(new_n659));
  NAND2_X1  g234(.A1(new_n659), .A2(G14), .ZN(new_n660));
  INV_X1    g235(.A(new_n660), .ZN(G401));
  XOR2_X1   g236(.A(G2084), .B(G2090), .Z(new_n662));
  XNOR2_X1  g237(.A(G2072), .B(G2078), .ZN(new_n663));
  XOR2_X1   g238(.A(new_n663), .B(KEYINPUT93), .Z(new_n664));
  XOR2_X1   g239(.A(G2067), .B(G2678), .Z(new_n665));
  AOI21_X1  g240(.A(new_n662), .B1(new_n664), .B2(new_n665), .ZN(new_n666));
  XOR2_X1   g241(.A(new_n663), .B(KEYINPUT17), .Z(new_n667));
  OAI21_X1  g242(.A(new_n666), .B1(new_n665), .B2(new_n667), .ZN(new_n668));
  INV_X1    g243(.A(new_n665), .ZN(new_n669));
  NAND3_X1  g244(.A1(new_n669), .A2(new_n663), .A3(new_n662), .ZN(new_n670));
  XOR2_X1   g245(.A(new_n670), .B(KEYINPUT18), .Z(new_n671));
  NAND3_X1  g246(.A1(new_n667), .A2(new_n665), .A3(new_n662), .ZN(new_n672));
  NAND3_X1  g247(.A1(new_n668), .A2(new_n671), .A3(new_n672), .ZN(new_n673));
  XNOR2_X1  g248(.A(G2096), .B(G2100), .ZN(new_n674));
  XNOR2_X1  g249(.A(new_n673), .B(new_n674), .ZN(new_n675));
  INV_X1    g250(.A(new_n675), .ZN(G227));
  XOR2_X1   g251(.A(G1956), .B(G2474), .Z(new_n677));
  XOR2_X1   g252(.A(G1961), .B(G1966), .Z(new_n678));
  NOR2_X1   g253(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  INV_X1    g254(.A(new_n679), .ZN(new_n680));
  XNOR2_X1  g255(.A(G1971), .B(G1976), .ZN(new_n681));
  XNOR2_X1  g256(.A(new_n681), .B(KEYINPUT19), .ZN(new_n682));
  NOR2_X1   g257(.A1(new_n680), .A2(new_n682), .ZN(new_n683));
  NAND2_X1  g258(.A1(new_n677), .A2(new_n678), .ZN(new_n684));
  OR2_X1    g259(.A1(new_n682), .A2(new_n684), .ZN(new_n685));
  INV_X1    g260(.A(KEYINPUT20), .ZN(new_n686));
  AOI21_X1  g261(.A(new_n683), .B1(new_n685), .B2(new_n686), .ZN(new_n687));
  NAND3_X1  g262(.A1(new_n680), .A2(new_n682), .A3(new_n684), .ZN(new_n688));
  OAI211_X1 g263(.A(new_n687), .B(new_n688), .C1(new_n686), .C2(new_n685), .ZN(new_n689));
  XOR2_X1   g264(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n690));
  XNOR2_X1  g265(.A(new_n689), .B(new_n690), .ZN(new_n691));
  XNOR2_X1  g266(.A(G1991), .B(G1996), .ZN(new_n692));
  INV_X1    g267(.A(G1981), .ZN(new_n693));
  XNOR2_X1  g268(.A(new_n692), .B(new_n693), .ZN(new_n694));
  XNOR2_X1  g269(.A(new_n694), .B(G1986), .ZN(new_n695));
  XNOR2_X1  g270(.A(new_n691), .B(new_n695), .ZN(G229));
  NOR2_X1   g271(.A1(G4), .A2(G16), .ZN(new_n697));
  AOI21_X1  g272(.A(new_n697), .B1(new_n620), .B2(G16), .ZN(new_n698));
  INV_X1    g273(.A(G1348), .ZN(new_n699));
  OR2_X1    g274(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  NAND2_X1  g275(.A1(new_n698), .A2(new_n699), .ZN(new_n701));
  INV_X1    g276(.A(G29), .ZN(new_n702));
  NOR2_X1   g277(.A1(G164), .A2(new_n702), .ZN(new_n703));
  AOI21_X1  g278(.A(new_n703), .B1(G27), .B2(new_n702), .ZN(new_n704));
  INV_X1    g279(.A(new_n704), .ZN(new_n705));
  AOI22_X1  g280(.A1(new_n700), .A2(new_n701), .B1(G2078), .B2(new_n705), .ZN(new_n706));
  NAND2_X1  g281(.A1(new_n702), .A2(G35), .ZN(new_n707));
  OAI21_X1  g282(.A(new_n707), .B1(G162), .B2(new_n702), .ZN(new_n708));
  XOR2_X1   g283(.A(new_n708), .B(KEYINPUT29), .Z(new_n709));
  INV_X1    g284(.A(G2090), .ZN(new_n710));
  NAND2_X1  g285(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  OR2_X1    g286(.A1(KEYINPUT24), .A2(G34), .ZN(new_n712));
  NAND2_X1  g287(.A1(KEYINPUT24), .A2(G34), .ZN(new_n713));
  NAND3_X1  g288(.A1(new_n712), .A2(new_n702), .A3(new_n713), .ZN(new_n714));
  OAI21_X1  g289(.A(new_n714), .B1(G160), .B2(new_n702), .ZN(new_n715));
  XNOR2_X1  g290(.A(new_n715), .B(G2084), .ZN(new_n716));
  INV_X1    g291(.A(G16), .ZN(new_n717));
  NAND2_X1  g292(.A1(new_n717), .A2(G5), .ZN(new_n718));
  OAI21_X1  g293(.A(new_n718), .B1(G171), .B2(new_n717), .ZN(new_n719));
  XOR2_X1   g294(.A(new_n719), .B(KEYINPUT99), .Z(new_n720));
  INV_X1    g295(.A(new_n720), .ZN(new_n721));
  INV_X1    g296(.A(G1961), .ZN(new_n722));
  AOI21_X1  g297(.A(new_n716), .B1(new_n721), .B2(new_n722), .ZN(new_n723));
  OR2_X1    g298(.A1(G29), .A2(G33), .ZN(new_n724));
  NAND2_X1  g299(.A1(G115), .A2(G2104), .ZN(new_n725));
  INV_X1    g300(.A(G127), .ZN(new_n726));
  OAI21_X1  g301(.A(new_n725), .B1(new_n481), .B2(new_n726), .ZN(new_n727));
  NAND2_X1  g302(.A1(new_n727), .A2(G2105), .ZN(new_n728));
  NAND3_X1  g303(.A1(new_n471), .A2(G103), .A3(G2104), .ZN(new_n729));
  XOR2_X1   g304(.A(new_n729), .B(KEYINPUT25), .Z(new_n730));
  INV_X1    g305(.A(G139), .ZN(new_n731));
  OAI211_X1 g306(.A(new_n728), .B(new_n730), .C1(new_n731), .C2(new_n472), .ZN(new_n732));
  OAI21_X1  g307(.A(new_n724), .B1(new_n732), .B2(new_n702), .ZN(new_n733));
  INV_X1    g308(.A(G2072), .ZN(new_n734));
  NAND2_X1  g309(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  XNOR2_X1  g310(.A(new_n735), .B(KEYINPUT98), .ZN(new_n736));
  NAND4_X1  g311(.A1(new_n706), .A2(new_n711), .A3(new_n723), .A4(new_n736), .ZN(new_n737));
  INV_X1    g312(.A(KEYINPUT23), .ZN(new_n738));
  NAND2_X1  g313(.A1(new_n717), .A2(G20), .ZN(new_n739));
  AOI22_X1  g314(.A1(G299), .A2(G16), .B1(new_n738), .B2(new_n739), .ZN(new_n740));
  OAI21_X1  g315(.A(new_n740), .B1(new_n738), .B2(new_n739), .ZN(new_n741));
  INV_X1    g316(.A(G1956), .ZN(new_n742));
  XNOR2_X1  g317(.A(new_n741), .B(new_n742), .ZN(new_n743));
  OAI221_X1 g318(.A(new_n743), .B1(new_n722), .B2(new_n721), .C1(new_n710), .C2(new_n709), .ZN(new_n744));
  NAND2_X1  g319(.A1(new_n717), .A2(G19), .ZN(new_n745));
  OAI21_X1  g320(.A(new_n745), .B1(new_n557), .B2(new_n717), .ZN(new_n746));
  XNOR2_X1  g321(.A(new_n746), .B(G1341), .ZN(new_n747));
  NAND2_X1  g322(.A1(new_n702), .A2(G26), .ZN(new_n748));
  XNOR2_X1  g323(.A(new_n748), .B(KEYINPUT97), .ZN(new_n749));
  XNOR2_X1  g324(.A(new_n749), .B(KEYINPUT28), .ZN(new_n750));
  AND2_X1   g325(.A1(new_n489), .A2(G128), .ZN(new_n751));
  INV_X1    g326(.A(G140), .ZN(new_n752));
  OAI21_X1  g327(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n753));
  NOR2_X1   g328(.A1(new_n471), .A2(G116), .ZN(new_n754));
  OAI22_X1  g329(.A1(new_n472), .A2(new_n752), .B1(new_n753), .B2(new_n754), .ZN(new_n755));
  NOR2_X1   g330(.A1(new_n751), .A2(new_n755), .ZN(new_n756));
  OAI21_X1  g331(.A(new_n750), .B1(new_n756), .B2(new_n702), .ZN(new_n757));
  XNOR2_X1  g332(.A(new_n757), .B(G2067), .ZN(new_n758));
  NOR4_X1   g333(.A1(new_n737), .A2(new_n744), .A3(new_n747), .A4(new_n758), .ZN(new_n759));
  NAND2_X1  g334(.A1(new_n717), .A2(G23), .ZN(new_n760));
  INV_X1    g335(.A(G288), .ZN(new_n761));
  OAI21_X1  g336(.A(new_n760), .B1(new_n761), .B2(new_n717), .ZN(new_n762));
  XNOR2_X1  g337(.A(new_n762), .B(KEYINPUT33), .ZN(new_n763));
  XNOR2_X1  g338(.A(new_n763), .B(G1976), .ZN(new_n764));
  NAND2_X1  g339(.A1(new_n717), .A2(G6), .ZN(new_n765));
  OAI21_X1  g340(.A(new_n765), .B1(new_n591), .B2(new_n717), .ZN(new_n766));
  XOR2_X1   g341(.A(KEYINPUT32), .B(G1981), .Z(new_n767));
  XOR2_X1   g342(.A(new_n767), .B(KEYINPUT95), .Z(new_n768));
  XNOR2_X1  g343(.A(new_n766), .B(new_n768), .ZN(new_n769));
  NOR2_X1   g344(.A1(G16), .A2(G22), .ZN(new_n770));
  AOI21_X1  g345(.A(new_n770), .B1(G166), .B2(G16), .ZN(new_n771));
  INV_X1    g346(.A(G1971), .ZN(new_n772));
  XNOR2_X1  g347(.A(new_n771), .B(new_n772), .ZN(new_n773));
  NAND3_X1  g348(.A1(new_n764), .A2(new_n769), .A3(new_n773), .ZN(new_n774));
  XOR2_X1   g349(.A(new_n774), .B(KEYINPUT34), .Z(new_n775));
  NAND2_X1  g350(.A1(new_n717), .A2(G24), .ZN(new_n776));
  INV_X1    g351(.A(G290), .ZN(new_n777));
  OAI21_X1  g352(.A(new_n776), .B1(new_n777), .B2(new_n717), .ZN(new_n778));
  INV_X1    g353(.A(G1986), .ZN(new_n779));
  XNOR2_X1  g354(.A(new_n778), .B(new_n779), .ZN(new_n780));
  NAND2_X1  g355(.A1(new_n702), .A2(G25), .ZN(new_n781));
  OR2_X1    g356(.A1(G95), .A2(G2105), .ZN(new_n782));
  OAI211_X1 g357(.A(new_n782), .B(G2104), .C1(G107), .C2(new_n471), .ZN(new_n783));
  INV_X1    g358(.A(G131), .ZN(new_n784));
  OAI21_X1  g359(.A(new_n783), .B1(new_n472), .B2(new_n784), .ZN(new_n785));
  AOI21_X1  g360(.A(new_n785), .B1(new_n489), .B2(G119), .ZN(new_n786));
  OAI21_X1  g361(.A(new_n781), .B1(new_n786), .B2(new_n702), .ZN(new_n787));
  XNOR2_X1  g362(.A(KEYINPUT35), .B(G1991), .ZN(new_n788));
  XNOR2_X1  g363(.A(new_n788), .B(KEYINPUT94), .ZN(new_n789));
  XNOR2_X1  g364(.A(new_n787), .B(new_n789), .ZN(new_n790));
  INV_X1    g365(.A(KEYINPUT96), .ZN(new_n791));
  AOI21_X1  g366(.A(new_n790), .B1(new_n791), .B2(KEYINPUT36), .ZN(new_n792));
  NAND3_X1  g367(.A1(new_n775), .A2(new_n780), .A3(new_n792), .ZN(new_n793));
  NOR2_X1   g368(.A1(new_n791), .A2(KEYINPUT36), .ZN(new_n794));
  OR2_X1    g369(.A1(new_n793), .A2(new_n794), .ZN(new_n795));
  NAND2_X1  g370(.A1(new_n793), .A2(new_n794), .ZN(new_n796));
  OR2_X1    g371(.A1(new_n733), .A2(new_n734), .ZN(new_n797));
  INV_X1    g372(.A(G11), .ZN(new_n798));
  OR2_X1    g373(.A1(new_n798), .A2(KEYINPUT31), .ZN(new_n799));
  AOI22_X1  g374(.A1(new_n643), .A2(G29), .B1(KEYINPUT31), .B2(new_n798), .ZN(new_n800));
  INV_X1    g375(.A(KEYINPUT30), .ZN(new_n801));
  OR2_X1    g376(.A1(new_n801), .A2(G28), .ZN(new_n802));
  NAND2_X1  g377(.A1(new_n801), .A2(G28), .ZN(new_n803));
  NAND3_X1  g378(.A1(new_n802), .A2(new_n803), .A3(new_n702), .ZN(new_n804));
  NAND4_X1  g379(.A1(new_n797), .A2(new_n799), .A3(new_n800), .A4(new_n804), .ZN(new_n805));
  NOR2_X1   g380(.A1(G29), .A2(G32), .ZN(new_n806));
  NAND3_X1  g381(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n807));
  XOR2_X1   g382(.A(new_n807), .B(KEYINPUT26), .Z(new_n808));
  INV_X1    g383(.A(G105), .ZN(new_n809));
  INV_X1    g384(.A(G141), .ZN(new_n810));
  OAI221_X1 g385(.A(new_n808), .B1(new_n809), .B2(new_n475), .C1(new_n472), .C2(new_n810), .ZN(new_n811));
  AOI21_X1  g386(.A(new_n811), .B1(G129), .B2(new_n489), .ZN(new_n812));
  AOI21_X1  g387(.A(new_n806), .B1(new_n812), .B2(G29), .ZN(new_n813));
  INV_X1    g388(.A(new_n813), .ZN(new_n814));
  XOR2_X1   g389(.A(KEYINPUT27), .B(G1996), .Z(new_n815));
  INV_X1    g390(.A(new_n815), .ZN(new_n816));
  AOI21_X1  g391(.A(new_n805), .B1(new_n814), .B2(new_n816), .ZN(new_n817));
  NAND4_X1  g392(.A1(new_n759), .A2(new_n795), .A3(new_n796), .A4(new_n817), .ZN(new_n818));
  NOR2_X1   g393(.A1(new_n705), .A2(G2078), .ZN(new_n819));
  NOR2_X1   g394(.A1(new_n814), .A2(new_n816), .ZN(new_n820));
  NAND2_X1  g395(.A1(new_n717), .A2(G21), .ZN(new_n821));
  OAI21_X1  g396(.A(new_n821), .B1(G168), .B2(new_n717), .ZN(new_n822));
  INV_X1    g397(.A(G1966), .ZN(new_n823));
  XNOR2_X1  g398(.A(new_n822), .B(new_n823), .ZN(new_n824));
  INV_X1    g399(.A(new_n824), .ZN(new_n825));
  NOR4_X1   g400(.A1(new_n818), .A2(new_n819), .A3(new_n820), .A4(new_n825), .ZN(G311));
  NOR3_X1   g401(.A1(new_n818), .A2(new_n820), .A3(new_n825), .ZN(new_n827));
  INV_X1    g402(.A(new_n819), .ZN(new_n828));
  NAND2_X1  g403(.A1(new_n827), .A2(new_n828), .ZN(G150));
  NAND2_X1  g404(.A1(G80), .A2(G543), .ZN(new_n830));
  INV_X1    g405(.A(G67), .ZN(new_n831));
  OAI21_X1  g406(.A(new_n830), .B1(new_n513), .B2(new_n831), .ZN(new_n832));
  XNOR2_X1  g407(.A(new_n832), .B(KEYINPUT100), .ZN(new_n833));
  NOR2_X1   g408(.A1(new_n833), .A2(new_n514), .ZN(new_n834));
  INV_X1    g409(.A(G93), .ZN(new_n835));
  INV_X1    g410(.A(G55), .ZN(new_n836));
  OAI22_X1  g411(.A1(new_n520), .A2(new_n835), .B1(new_n547), .B2(new_n836), .ZN(new_n837));
  NOR2_X1   g412(.A1(new_n834), .A2(new_n837), .ZN(new_n838));
  INV_X1    g413(.A(new_n838), .ZN(new_n839));
  NAND2_X1  g414(.A1(new_n839), .A2(G860), .ZN(new_n840));
  XNOR2_X1  g415(.A(new_n840), .B(KEYINPUT101), .ZN(new_n841));
  XNOR2_X1  g416(.A(new_n841), .B(KEYINPUT37), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n620), .A2(G559), .ZN(new_n843));
  XNOR2_X1  g418(.A(new_n843), .B(KEYINPUT38), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n839), .A2(new_n557), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n838), .A2(new_n556), .ZN(new_n846));
  NAND2_X1  g421(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  XNOR2_X1  g422(.A(new_n847), .B(KEYINPUT39), .ZN(new_n848));
  XNOR2_X1  g423(.A(new_n844), .B(new_n848), .ZN(new_n849));
  OAI21_X1  g424(.A(new_n842), .B1(new_n849), .B2(G860), .ZN(G145));
  XOR2_X1   g425(.A(new_n732), .B(new_n786), .Z(new_n851));
  XNOR2_X1  g426(.A(new_n756), .B(KEYINPUT103), .ZN(new_n852));
  XNOR2_X1  g427(.A(new_n851), .B(new_n852), .ZN(new_n853));
  INV_X1    g428(.A(new_n812), .ZN(new_n854));
  XNOR2_X1  g429(.A(new_n854), .B(new_n503), .ZN(new_n855));
  XNOR2_X1  g430(.A(new_n853), .B(new_n855), .ZN(new_n856));
  XNOR2_X1  g431(.A(new_n634), .B(KEYINPUT104), .ZN(new_n857));
  INV_X1    g432(.A(G142), .ZN(new_n858));
  OAI21_X1  g433(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n859));
  NOR2_X1   g434(.A1(new_n471), .A2(G118), .ZN(new_n860));
  OAI22_X1  g435(.A1(new_n472), .A2(new_n858), .B1(new_n859), .B2(new_n860), .ZN(new_n861));
  AOI21_X1  g436(.A(new_n861), .B1(new_n489), .B2(G130), .ZN(new_n862));
  XNOR2_X1  g437(.A(new_n857), .B(new_n862), .ZN(new_n863));
  XNOR2_X1  g438(.A(new_n856), .B(new_n863), .ZN(new_n864));
  XNOR2_X1  g439(.A(G162), .B(KEYINPUT102), .ZN(new_n865));
  XNOR2_X1  g440(.A(new_n865), .B(G160), .ZN(new_n866));
  XNOR2_X1  g441(.A(new_n866), .B(new_n643), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n864), .A2(new_n867), .ZN(new_n868));
  XNOR2_X1  g443(.A(new_n868), .B(KEYINPUT105), .ZN(new_n869));
  INV_X1    g444(.A(G37), .ZN(new_n870));
  OAI211_X1 g445(.A(new_n869), .B(new_n870), .C1(new_n867), .C2(new_n864), .ZN(new_n871));
  XNOR2_X1  g446(.A(new_n871), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g447(.A1(new_n619), .A2(G299), .ZN(new_n873));
  NAND4_X1  g448(.A1(new_n611), .A2(new_n624), .A3(new_n617), .A4(new_n618), .ZN(new_n874));
  NAND2_X1  g449(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  INV_X1    g450(.A(new_n875), .ZN(new_n876));
  NAND3_X1  g451(.A1(new_n873), .A2(KEYINPUT41), .A3(new_n874), .ZN(new_n877));
  INV_X1    g452(.A(new_n877), .ZN(new_n878));
  AOI21_X1  g453(.A(KEYINPUT41), .B1(new_n873), .B2(new_n874), .ZN(new_n879));
  NOR2_X1   g454(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  XNOR2_X1  g455(.A(new_n629), .B(new_n847), .ZN(new_n881));
  MUX2_X1   g456(.A(new_n876), .B(new_n880), .S(new_n881), .Z(new_n882));
  NAND2_X1  g457(.A1(new_n777), .A2(new_n761), .ZN(new_n883));
  NAND2_X1  g458(.A1(G290), .A2(G288), .ZN(new_n884));
  AOI21_X1  g459(.A(G303), .B1(new_n883), .B2(new_n884), .ZN(new_n885));
  INV_X1    g460(.A(new_n885), .ZN(new_n886));
  NAND3_X1  g461(.A1(new_n883), .A2(G303), .A3(new_n884), .ZN(new_n887));
  AOI21_X1  g462(.A(new_n591), .B1(new_n886), .B2(new_n887), .ZN(new_n888));
  INV_X1    g463(.A(new_n887), .ZN(new_n889));
  NOR3_X1   g464(.A1(new_n889), .A2(new_n885), .A3(G305), .ZN(new_n890));
  NOR2_X1   g465(.A1(new_n888), .A2(new_n890), .ZN(new_n891));
  XOR2_X1   g466(.A(new_n891), .B(KEYINPUT42), .Z(new_n892));
  XNOR2_X1  g467(.A(new_n882), .B(new_n892), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n893), .A2(G868), .ZN(new_n894));
  OAI21_X1  g469(.A(new_n894), .B1(G868), .B2(new_n838), .ZN(G295));
  OAI21_X1  g470(.A(new_n894), .B1(G868), .B2(new_n838), .ZN(G331));
  INV_X1    g471(.A(KEYINPUT43), .ZN(new_n897));
  NAND2_X1  g472(.A1(G286), .A2(G171), .ZN(new_n898));
  NAND2_X1  g473(.A1(G301), .A2(G168), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n900), .A2(new_n847), .ZN(new_n901));
  NAND4_X1  g476(.A1(new_n898), .A2(new_n845), .A3(new_n846), .A4(new_n899), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  NOR2_X1   g478(.A1(new_n875), .A2(new_n903), .ZN(new_n904));
  INV_X1    g479(.A(KEYINPUT107), .ZN(new_n905));
  NAND3_X1  g480(.A1(new_n900), .A2(new_n905), .A3(new_n847), .ZN(new_n906));
  OAI21_X1  g481(.A(new_n906), .B1(new_n903), .B2(new_n905), .ZN(new_n907));
  INV_X1    g482(.A(new_n907), .ZN(new_n908));
  AOI21_X1  g483(.A(new_n904), .B1(new_n880), .B2(new_n908), .ZN(new_n909));
  AOI21_X1  g484(.A(G37), .B1(new_n909), .B2(new_n891), .ZN(new_n910));
  INV_X1    g485(.A(KEYINPUT108), .ZN(new_n911));
  INV_X1    g486(.A(new_n879), .ZN(new_n912));
  NAND3_X1  g487(.A1(new_n912), .A2(new_n877), .A3(new_n903), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n907), .A2(new_n876), .ZN(new_n914));
  AOI211_X1 g489(.A(new_n911), .B(new_n891), .C1(new_n913), .C2(new_n914), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n913), .A2(new_n914), .ZN(new_n916));
  INV_X1    g491(.A(new_n891), .ZN(new_n917));
  AOI21_X1  g492(.A(KEYINPUT108), .B1(new_n916), .B2(new_n917), .ZN(new_n918));
  OAI211_X1 g493(.A(new_n897), .B(new_n910), .C1(new_n915), .C2(new_n918), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n919), .A2(KEYINPUT109), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n916), .A2(new_n917), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n921), .A2(new_n911), .ZN(new_n922));
  NAND3_X1  g497(.A1(new_n916), .A2(KEYINPUT108), .A3(new_n917), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  INV_X1    g499(.A(KEYINPUT109), .ZN(new_n925));
  NAND4_X1  g500(.A1(new_n924), .A2(new_n925), .A3(new_n897), .A4(new_n910), .ZN(new_n926));
  INV_X1    g501(.A(new_n910), .ZN(new_n927));
  NOR2_X1   g502(.A1(new_n909), .A2(new_n891), .ZN(new_n928));
  OAI21_X1  g503(.A(KEYINPUT43), .B1(new_n927), .B2(new_n928), .ZN(new_n929));
  NAND3_X1  g504(.A1(new_n920), .A2(new_n926), .A3(new_n929), .ZN(new_n930));
  XNOR2_X1  g505(.A(KEYINPUT106), .B(KEYINPUT44), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  OAI211_X1 g507(.A(new_n910), .B(new_n897), .C1(new_n891), .C2(new_n909), .ZN(new_n933));
  AOI21_X1  g508(.A(new_n927), .B1(new_n922), .B2(new_n923), .ZN(new_n934));
  OAI211_X1 g509(.A(new_n933), .B(KEYINPUT44), .C1(new_n934), .C2(new_n897), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n932), .A2(new_n935), .ZN(new_n936));
  INV_X1    g511(.A(KEYINPUT110), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  NAND3_X1  g513(.A1(new_n932), .A2(KEYINPUT110), .A3(new_n935), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n938), .A2(new_n939), .ZN(G397));
  INV_X1    g515(.A(G1384), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n503), .A2(new_n941), .ZN(new_n942));
  INV_X1    g517(.A(KEYINPUT45), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  NAND2_X1  g519(.A1(G160), .A2(G40), .ZN(new_n945));
  NOR2_X1   g520(.A1(new_n944), .A2(new_n945), .ZN(new_n946));
  XNOR2_X1  g521(.A(new_n946), .B(KEYINPUT112), .ZN(new_n947));
  INV_X1    g522(.A(G1996), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n946), .A2(new_n948), .ZN(new_n949));
  XNOR2_X1  g524(.A(new_n949), .B(KEYINPUT111), .ZN(new_n950));
  INV_X1    g525(.A(new_n950), .ZN(new_n951));
  INV_X1    g526(.A(G2067), .ZN(new_n952));
  NOR2_X1   g527(.A1(new_n756), .A2(new_n952), .ZN(new_n953));
  NOR3_X1   g528(.A1(new_n751), .A2(G2067), .A3(new_n755), .ZN(new_n954));
  NOR2_X1   g529(.A1(new_n953), .A2(new_n954), .ZN(new_n955));
  OAI21_X1  g530(.A(new_n955), .B1(new_n948), .B2(new_n812), .ZN(new_n956));
  AOI22_X1  g531(.A1(new_n951), .A2(new_n812), .B1(new_n947), .B2(new_n956), .ZN(new_n957));
  INV_X1    g532(.A(new_n788), .ZN(new_n958));
  AND3_X1   g533(.A1(new_n957), .A2(new_n786), .A3(new_n958), .ZN(new_n959));
  OAI21_X1  g534(.A(new_n947), .B1(new_n959), .B2(new_n954), .ZN(new_n960));
  INV_X1    g535(.A(new_n955), .ZN(new_n961));
  OAI21_X1  g536(.A(new_n947), .B1(new_n854), .B2(new_n961), .ZN(new_n962));
  AND2_X1   g537(.A1(new_n950), .A2(KEYINPUT46), .ZN(new_n963));
  NOR2_X1   g538(.A1(new_n950), .A2(KEYINPUT46), .ZN(new_n964));
  OAI21_X1  g539(.A(new_n962), .B1(new_n963), .B2(new_n964), .ZN(new_n965));
  XNOR2_X1  g540(.A(new_n965), .B(KEYINPUT47), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n960), .A2(new_n966), .ZN(new_n967));
  INV_X1    g542(.A(new_n957), .ZN(new_n968));
  XNOR2_X1  g543(.A(new_n786), .B(new_n958), .ZN(new_n969));
  AOI21_X1  g544(.A(new_n968), .B1(new_n969), .B2(new_n947), .ZN(new_n970));
  NAND3_X1  g545(.A1(new_n946), .A2(new_n779), .A3(new_n777), .ZN(new_n971));
  XNOR2_X1  g546(.A(new_n971), .B(KEYINPUT48), .ZN(new_n972));
  AOI21_X1  g547(.A(new_n967), .B1(new_n970), .B2(new_n972), .ZN(new_n973));
  INV_X1    g548(.A(KEYINPUT127), .ZN(new_n974));
  INV_X1    g549(.A(KEYINPUT53), .ZN(new_n975));
  NAND3_X1  g550(.A1(new_n503), .A2(KEYINPUT45), .A3(new_n941), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n976), .A2(KEYINPUT113), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n977), .A2(new_n944), .ZN(new_n978));
  INV_X1    g553(.A(new_n945), .ZN(new_n979));
  AOI21_X1  g554(.A(G1384), .B1(new_n498), .B2(new_n502), .ZN(new_n980));
  INV_X1    g555(.A(KEYINPUT113), .ZN(new_n981));
  NOR3_X1   g556(.A1(new_n980), .A2(new_n981), .A3(KEYINPUT45), .ZN(new_n982));
  INV_X1    g557(.A(new_n982), .ZN(new_n983));
  NAND3_X1  g558(.A1(new_n978), .A2(new_n979), .A3(new_n983), .ZN(new_n984));
  OAI21_X1  g559(.A(new_n975), .B1(new_n984), .B2(G2078), .ZN(new_n985));
  NAND3_X1  g560(.A1(new_n944), .A2(new_n979), .A3(new_n976), .ZN(new_n986));
  OR3_X1    g561(.A1(new_n986), .A2(new_n975), .A3(G2078), .ZN(new_n987));
  INV_X1    g562(.A(KEYINPUT50), .ZN(new_n988));
  NOR2_X1   g563(.A1(new_n980), .A2(new_n988), .ZN(new_n989));
  AOI211_X1 g564(.A(KEYINPUT50), .B(G1384), .C1(new_n498), .C2(new_n502), .ZN(new_n990));
  NOR3_X1   g565(.A1(new_n989), .A2(new_n990), .A3(new_n945), .ZN(new_n991));
  OAI211_X1 g566(.A(new_n985), .B(new_n987), .C1(G1961), .C2(new_n991), .ZN(new_n992));
  NAND2_X1  g567(.A1(new_n992), .A2(G171), .ZN(new_n993));
  INV_X1    g568(.A(KEYINPUT51), .ZN(new_n994));
  INV_X1    g569(.A(KEYINPUT117), .ZN(new_n995));
  NOR2_X1   g570(.A1(new_n980), .A2(KEYINPUT45), .ZN(new_n996));
  AOI211_X1 g571(.A(new_n943), .B(G1384), .C1(new_n498), .C2(new_n502), .ZN(new_n997));
  NOR3_X1   g572(.A1(new_n996), .A2(new_n997), .A3(new_n945), .ZN(new_n998));
  OAI21_X1  g573(.A(new_n995), .B1(new_n998), .B2(G1966), .ZN(new_n999));
  INV_X1    g574(.A(G2084), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n991), .A2(new_n1000), .ZN(new_n1001));
  NAND3_X1  g576(.A1(new_n986), .A2(KEYINPUT117), .A3(new_n823), .ZN(new_n1002));
  NAND4_X1  g577(.A1(new_n999), .A2(G168), .A3(new_n1001), .A4(new_n1002), .ZN(new_n1003));
  AOI21_X1  g578(.A(new_n994), .B1(new_n1003), .B2(G8), .ZN(new_n1004));
  NAND3_X1  g579(.A1(new_n999), .A2(new_n1001), .A3(new_n1002), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n1005), .A2(G286), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n1006), .A2(KEYINPUT51), .ZN(new_n1007));
  AND2_X1   g582(.A1(new_n1003), .A2(G8), .ZN(new_n1008));
  AOI21_X1  g583(.A(new_n1004), .B1(new_n1007), .B2(new_n1008), .ZN(new_n1009));
  INV_X1    g584(.A(KEYINPUT62), .ZN(new_n1010));
  AOI21_X1  g585(.A(new_n993), .B1(new_n1009), .B2(new_n1010), .ZN(new_n1011));
  NOR4_X1   g586(.A1(new_n989), .A2(new_n990), .A3(G2090), .A4(new_n945), .ZN(new_n1012));
  AOI21_X1  g587(.A(new_n1012), .B1(new_n984), .B2(new_n772), .ZN(new_n1013));
  INV_X1    g588(.A(KEYINPUT114), .ZN(new_n1014));
  NOR2_X1   g589(.A1(new_n1013), .A2(new_n1014), .ZN(new_n1015));
  AOI211_X1 g590(.A(KEYINPUT114), .B(new_n1012), .C1(new_n984), .C2(new_n772), .ZN(new_n1016));
  NOR2_X1   g591(.A1(new_n1015), .A2(new_n1016), .ZN(new_n1017));
  NAND2_X1  g592(.A1(G303), .A2(G8), .ZN(new_n1018));
  XNOR2_X1  g593(.A(new_n1018), .B(KEYINPUT55), .ZN(new_n1019));
  INV_X1    g594(.A(new_n1019), .ZN(new_n1020));
  NAND4_X1  g595(.A1(new_n1017), .A2(KEYINPUT115), .A3(G8), .A4(new_n1020), .ZN(new_n1021));
  INV_X1    g596(.A(new_n1012), .ZN(new_n1022));
  AOI21_X1  g597(.A(new_n981), .B1(new_n980), .B2(KEYINPUT45), .ZN(new_n1023));
  NOR2_X1   g598(.A1(new_n1023), .A2(new_n996), .ZN(new_n1024));
  NOR3_X1   g599(.A1(new_n1024), .A2(new_n945), .A3(new_n982), .ZN(new_n1025));
  OAI21_X1  g600(.A(new_n1022), .B1(new_n1025), .B2(G1971), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n1026), .A2(KEYINPUT114), .ZN(new_n1027));
  NAND2_X1  g602(.A1(new_n1013), .A2(new_n1014), .ZN(new_n1028));
  NAND4_X1  g603(.A1(new_n1027), .A2(G8), .A3(new_n1020), .A4(new_n1028), .ZN(new_n1029));
  INV_X1    g604(.A(KEYINPUT115), .ZN(new_n1030));
  NAND2_X1  g605(.A1(new_n1029), .A2(new_n1030), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n1021), .A2(new_n1031), .ZN(new_n1032));
  INV_X1    g607(.A(G8), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n979), .A2(new_n980), .ZN(new_n1034));
  INV_X1    g609(.A(new_n1034), .ZN(new_n1035));
  AOI211_X1 g610(.A(new_n1033), .B(new_n1035), .C1(G1976), .C2(new_n761), .ZN(new_n1036));
  INV_X1    g611(.A(KEYINPUT52), .ZN(new_n1037));
  OR2_X1    g612(.A1(new_n1036), .A2(new_n1037), .ZN(new_n1038));
  OAI211_X1 g613(.A(new_n1036), .B(new_n1037), .C1(G1976), .C2(new_n761), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n591), .A2(new_n693), .ZN(new_n1040));
  INV_X1    g615(.A(new_n586), .ZN(new_n1041));
  OAI21_X1  g616(.A(G1981), .B1(new_n1041), .B2(new_n590), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n1040), .A2(new_n1042), .ZN(new_n1043));
  INV_X1    g618(.A(KEYINPUT49), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n1043), .A2(new_n1044), .ZN(new_n1045));
  NOR2_X1   g620(.A1(new_n1035), .A2(new_n1033), .ZN(new_n1046));
  NAND3_X1  g621(.A1(new_n1040), .A2(KEYINPUT49), .A3(new_n1042), .ZN(new_n1047));
  NAND3_X1  g622(.A1(new_n1045), .A2(new_n1046), .A3(new_n1047), .ZN(new_n1048));
  NAND3_X1  g623(.A1(new_n1038), .A2(new_n1039), .A3(new_n1048), .ZN(new_n1049));
  AOI21_X1  g624(.A(new_n1020), .B1(new_n1026), .B2(G8), .ZN(new_n1050));
  NOR2_X1   g625(.A1(new_n1049), .A2(new_n1050), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n1003), .A2(G8), .ZN(new_n1052));
  AOI21_X1  g627(.A(new_n1052), .B1(KEYINPUT51), .B2(new_n1006), .ZN(new_n1053));
  OAI21_X1  g628(.A(KEYINPUT62), .B1(new_n1053), .B2(new_n1004), .ZN(new_n1054));
  NAND4_X1  g629(.A1(new_n1011), .A2(new_n1032), .A3(new_n1051), .A4(new_n1054), .ZN(new_n1055));
  INV_X1    g630(.A(new_n1049), .ZN(new_n1056));
  NAND3_X1  g631(.A1(new_n1021), .A2(new_n1031), .A3(new_n1056), .ZN(new_n1057));
  INV_X1    g632(.A(G1976), .ZN(new_n1058));
  NAND3_X1  g633(.A1(new_n1048), .A2(new_n1058), .A3(new_n761), .ZN(new_n1059));
  AND2_X1   g634(.A1(new_n1059), .A2(new_n1040), .ZN(new_n1060));
  OR2_X1    g635(.A1(new_n1060), .A2(KEYINPUT116), .ZN(new_n1061));
  NAND2_X1  g636(.A1(new_n1060), .A2(KEYINPUT116), .ZN(new_n1062));
  NAND3_X1  g637(.A1(new_n1061), .A2(new_n1046), .A3(new_n1062), .ZN(new_n1063));
  NAND3_X1  g638(.A1(new_n1055), .A2(new_n1057), .A3(new_n1063), .ZN(new_n1064));
  XNOR2_X1  g639(.A(new_n992), .B(G301), .ZN(new_n1065));
  XNOR2_X1  g640(.A(new_n1065), .B(KEYINPUT54), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n1032), .A2(new_n1051), .ZN(new_n1067));
  NOR2_X1   g642(.A1(new_n1066), .A2(new_n1067), .ZN(new_n1068));
  INV_X1    g643(.A(KEYINPUT120), .ZN(new_n1069));
  NOR2_X1   g644(.A1(new_n1069), .A2(KEYINPUT57), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n1069), .A2(KEYINPUT57), .ZN(new_n1071));
  XOR2_X1   g646(.A(new_n1071), .B(KEYINPUT121), .Z(new_n1072));
  INV_X1    g647(.A(new_n1072), .ZN(new_n1073));
  OR3_X1    g648(.A1(G299), .A2(new_n1070), .A3(new_n1073), .ZN(new_n1074));
  OAI21_X1  g649(.A(new_n1073), .B1(G299), .B2(new_n1070), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n1074), .A2(new_n1075), .ZN(new_n1076));
  NOR2_X1   g651(.A1(new_n989), .A2(new_n990), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n1077), .A2(new_n979), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n1078), .A2(new_n742), .ZN(new_n1079));
  XNOR2_X1  g654(.A(KEYINPUT56), .B(G2072), .ZN(new_n1080));
  NAND4_X1  g655(.A1(new_n978), .A2(new_n983), .A3(new_n979), .A4(new_n1080), .ZN(new_n1081));
  NAND3_X1  g656(.A1(new_n1076), .A2(new_n1079), .A3(new_n1081), .ZN(new_n1082));
  INV_X1    g657(.A(KEYINPUT122), .ZN(new_n1083));
  OR2_X1    g658(.A1(new_n1082), .A2(new_n1083), .ZN(new_n1084));
  AOI21_X1  g659(.A(new_n1076), .B1(new_n1079), .B2(new_n1081), .ZN(new_n1085));
  INV_X1    g660(.A(new_n1085), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n1082), .A2(new_n1083), .ZN(new_n1087));
  NAND3_X1  g662(.A1(new_n1084), .A2(new_n1086), .A3(new_n1087), .ZN(new_n1088));
  INV_X1    g663(.A(KEYINPUT61), .ZN(new_n1089));
  NOR2_X1   g664(.A1(new_n1082), .A2(KEYINPUT124), .ZN(new_n1090));
  NOR2_X1   g665(.A1(new_n1090), .A2(new_n1089), .ZN(new_n1091));
  AOI21_X1  g666(.A(new_n1085), .B1(KEYINPUT124), .B2(new_n1082), .ZN(new_n1092));
  AOI22_X1  g667(.A1(new_n1088), .A2(new_n1089), .B1(new_n1091), .B2(new_n1092), .ZN(new_n1093));
  AOI22_X1  g668(.A1(new_n1078), .A2(new_n699), .B1(new_n952), .B2(new_n1035), .ZN(new_n1094));
  NAND3_X1  g669(.A1(new_n1094), .A2(KEYINPUT60), .A3(new_n619), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n1095), .A2(KEYINPUT125), .ZN(new_n1096));
  INV_X1    g671(.A(KEYINPUT126), .ZN(new_n1097));
  OAI22_X1  g672(.A1(new_n991), .A2(G1348), .B1(G2067), .B2(new_n1034), .ZN(new_n1098));
  INV_X1    g673(.A(KEYINPUT60), .ZN(new_n1099));
  NOR2_X1   g674(.A1(new_n1098), .A2(new_n1099), .ZN(new_n1100));
  OAI21_X1  g675(.A(new_n1097), .B1(new_n1100), .B2(new_n619), .ZN(new_n1101));
  INV_X1    g676(.A(KEYINPUT125), .ZN(new_n1102));
  NAND3_X1  g677(.A1(new_n1100), .A2(new_n1102), .A3(new_n619), .ZN(new_n1103));
  INV_X1    g678(.A(new_n619), .ZN(new_n1104));
  OAI211_X1 g679(.A(new_n1104), .B(KEYINPUT126), .C1(new_n1098), .C2(new_n1099), .ZN(new_n1105));
  NAND4_X1  g680(.A1(new_n1096), .A2(new_n1101), .A3(new_n1103), .A4(new_n1105), .ZN(new_n1106));
  OAI21_X1  g681(.A(new_n1106), .B1(KEYINPUT60), .B2(new_n1094), .ZN(new_n1107));
  XNOR2_X1  g682(.A(KEYINPUT58), .B(G1341), .ZN(new_n1108));
  OAI22_X1  g683(.A1(new_n984), .A2(G1996), .B1(new_n1035), .B2(new_n1108), .ZN(new_n1109));
  XNOR2_X1  g684(.A(new_n1109), .B(KEYINPUT123), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n1110), .A2(new_n557), .ZN(new_n1111));
  INV_X1    g686(.A(KEYINPUT59), .ZN(new_n1112));
  NAND2_X1  g687(.A1(new_n1111), .A2(new_n1112), .ZN(new_n1113));
  NAND3_X1  g688(.A1(new_n1110), .A2(KEYINPUT59), .A3(new_n557), .ZN(new_n1114));
  NAND4_X1  g689(.A1(new_n1093), .A2(new_n1107), .A3(new_n1113), .A4(new_n1114), .ZN(new_n1115));
  OAI21_X1  g690(.A(new_n1086), .B1(new_n619), .B2(new_n1094), .ZN(new_n1116));
  NAND3_X1  g691(.A1(new_n1116), .A2(new_n1084), .A3(new_n1087), .ZN(new_n1117));
  AOI21_X1  g692(.A(new_n1009), .B1(new_n1115), .B2(new_n1117), .ZN(new_n1118));
  AOI21_X1  g693(.A(new_n1064), .B1(new_n1068), .B2(new_n1118), .ZN(new_n1119));
  AND3_X1   g694(.A1(new_n1005), .A2(G8), .A3(G168), .ZN(new_n1120));
  AND2_X1   g695(.A1(new_n1029), .A2(new_n1030), .ZN(new_n1121));
  NOR2_X1   g696(.A1(new_n1029), .A2(new_n1030), .ZN(new_n1122));
  OAI211_X1 g697(.A(new_n1051), .B(new_n1120), .C1(new_n1121), .C2(new_n1122), .ZN(new_n1123));
  NAND2_X1  g698(.A1(new_n1123), .A2(KEYINPUT118), .ZN(new_n1124));
  INV_X1    g699(.A(KEYINPUT63), .ZN(new_n1125));
  INV_X1    g700(.A(KEYINPUT118), .ZN(new_n1126));
  NAND4_X1  g701(.A1(new_n1032), .A2(new_n1126), .A3(new_n1051), .A4(new_n1120), .ZN(new_n1127));
  NAND3_X1  g702(.A1(new_n1124), .A2(new_n1125), .A3(new_n1127), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n1017), .A2(G8), .ZN(new_n1129));
  AOI21_X1  g704(.A(new_n1049), .B1(new_n1129), .B2(new_n1019), .ZN(new_n1130));
  OR2_X1    g705(.A1(new_n1130), .A2(KEYINPUT119), .ZN(new_n1131));
  AOI21_X1  g706(.A(new_n1125), .B1(new_n1130), .B2(KEYINPUT119), .ZN(new_n1132));
  NAND4_X1  g707(.A1(new_n1131), .A2(new_n1132), .A3(new_n1032), .A4(new_n1120), .ZN(new_n1133));
  NAND2_X1  g708(.A1(new_n1128), .A2(new_n1133), .ZN(new_n1134));
  NAND2_X1  g709(.A1(new_n1119), .A2(new_n1134), .ZN(new_n1135));
  XNOR2_X1  g710(.A(G290), .B(G1986), .ZN(new_n1136));
  NAND2_X1  g711(.A1(new_n1136), .A2(new_n946), .ZN(new_n1137));
  NAND2_X1  g712(.A1(new_n970), .A2(new_n1137), .ZN(new_n1138));
  INV_X1    g713(.A(new_n1138), .ZN(new_n1139));
  AOI21_X1  g714(.A(new_n974), .B1(new_n1135), .B2(new_n1139), .ZN(new_n1140));
  AOI211_X1 g715(.A(KEYINPUT127), .B(new_n1138), .C1(new_n1119), .C2(new_n1134), .ZN(new_n1141));
  OAI21_X1  g716(.A(new_n973), .B1(new_n1140), .B2(new_n1141), .ZN(G329));
  assign    G231 = 1'b0;
  AND3_X1   g717(.A1(new_n871), .A2(new_n660), .A3(new_n675), .ZN(new_n1144));
  INV_X1    g718(.A(G229), .ZN(new_n1145));
  NAND4_X1  g719(.A1(new_n1144), .A2(G319), .A3(new_n1145), .A4(new_n930), .ZN(G225));
  INV_X1    g720(.A(G225), .ZN(G308));
endmodule


