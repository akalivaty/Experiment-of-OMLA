

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
         n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597,
         n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608,
         n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619,
         n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630,
         n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641,
         n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652,
         n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663,
         n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674,
         n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685,
         n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696,
         n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707,
         n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718,
         n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729,
         n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740,
         n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751,
         n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762,
         n763, n764, n765, n766, n767, n768;

  OR2_X1 U378 ( .A1(n571), .A2(n569), .ZN(n657) );
  NOR2_X1 U379 ( .A1(n768), .A2(n767), .ZN(n564) );
  AND2_X4 U380 ( .A1(n452), .A2(n451), .ZN(n734) );
  OR2_X1 U381 ( .A1(n635), .A2(n741), .ZN(n429) );
  XNOR2_X2 U382 ( .A(n408), .B(G119), .ZN(n491) );
  XNOR2_X2 U383 ( .A(G101), .B(KEYINPUT3), .ZN(n408) );
  OR2_X1 U384 ( .A1(n582), .A2(n465), .ZN(n464) );
  NAND2_X2 U385 ( .A1(n589), .A2(n590), .ZN(n436) );
  XOR2_X2 U386 ( .A(G137), .B(G140), .Z(n522) );
  INV_X2 U387 ( .A(G953), .ZN(n760) );
  AND2_X1 U388 ( .A1(n413), .A2(n411), .ZN(n410) );
  XNOR2_X1 U389 ( .A(n416), .B(n601), .ZN(n618) );
  NOR2_X1 U390 ( .A1(n554), .A2(n553), .ZN(n567) );
  XOR2_X1 U391 ( .A(KEYINPUT23), .B(KEYINPUT95), .Z(n526) );
  NOR2_X1 U392 ( .A1(n635), .A2(n428), .ZN(n450) );
  NAND2_X1 U393 ( .A1(n410), .A2(n409), .ZN(n412) );
  AND2_X1 U394 ( .A1(n437), .A2(KEYINPUT44), .ZN(n362) );
  XNOR2_X1 U395 ( .A(n577), .B(KEYINPUT83), .ZN(n409) );
  NOR2_X1 U396 ( .A1(n620), .A2(n399), .ZN(n643) );
  XNOR2_X1 U397 ( .A(n401), .B(n366), .ZN(n695) );
  XNOR2_X1 U398 ( .A(n532), .B(n531), .ZN(n675) );
  XNOR2_X1 U399 ( .A(n736), .B(n735), .ZN(n737) );
  XNOR2_X1 U400 ( .A(n727), .B(n726), .ZN(n728) );
  XNOR2_X1 U401 ( .A(n456), .B(n754), .ZN(n736) );
  OR2_X1 U402 ( .A1(n727), .A2(G902), .ZN(n396) );
  XNOR2_X1 U403 ( .A(n510), .B(n509), .ZN(n727) );
  XNOR2_X1 U404 ( .A(n503), .B(n454), .ZN(n521) );
  XNOR2_X1 U405 ( .A(n526), .B(n523), .ZN(n415) );
  XNOR2_X1 U406 ( .A(G128), .B(G119), .ZN(n523) );
  XNOR2_X1 U407 ( .A(G125), .B(G146), .ZN(n418) );
  XNOR2_X1 U408 ( .A(G116), .B(G107), .ZN(n490) );
  BUF_X1 U409 ( .A(n548), .Z(n673) );
  XOR2_X2 U410 ( .A(G143), .B(G128), .Z(n513) );
  XNOR2_X1 U411 ( .A(n548), .B(KEYINPUT106), .ZN(n621) );
  XNOR2_X2 U412 ( .A(n566), .B(KEYINPUT19), .ZN(n589) );
  NAND2_X2 U413 ( .A1(n382), .A2(n689), .ZN(n566) );
  XNOR2_X1 U414 ( .A(n718), .B(n717), .ZN(n719) );
  XNOR2_X2 U415 ( .A(n513), .B(n482), .ZN(n488) );
  AND2_X1 U416 ( .A1(n670), .A2(n557), .ZN(n558) );
  XOR2_X1 U417 ( .A(KEYINPUT15), .B(G902), .Z(n636) );
  XNOR2_X1 U418 ( .A(n378), .B(n358), .ZN(n548) );
  OR2_X1 U419 ( .A1(n500), .A2(G902), .ZN(n378) );
  XNOR2_X1 U420 ( .A(n379), .B(n753), .ZN(n500) );
  XNOR2_X1 U421 ( .A(n423), .B(n422), .ZN(n379) );
  XNOR2_X1 U422 ( .A(n480), .B(n487), .ZN(n423) );
  XNOR2_X1 U423 ( .A(n491), .B(n405), .ZN(n422) );
  XNOR2_X1 U424 ( .A(n521), .B(n522), .ZN(n754) );
  INV_X1 U425 ( .A(n643), .ZN(n398) );
  AND2_X1 U426 ( .A1(n665), .A2(n581), .ZN(n411) );
  NAND2_X1 U427 ( .A1(n469), .A2(n666), .ZN(n468) );
  NAND2_X1 U428 ( .A1(n468), .A2(KEYINPUT87), .ZN(n467) );
  XNOR2_X1 U429 ( .A(G113), .B(G104), .ZN(n441) );
  XNOR2_X1 U430 ( .A(n584), .B(KEYINPUT1), .ZN(n593) );
  AND2_X1 U431 ( .A1(n593), .A2(n414), .ZN(n603) );
  NOR2_X1 U432 ( .A1(n736), .A2(G902), .ZN(n532) );
  XNOR2_X1 U433 ( .A(n516), .B(n515), .ZN(n525) );
  INV_X1 U434 ( .A(KEYINPUT10), .ZN(n454) );
  INV_X1 U435 ( .A(n418), .ZN(n503) );
  XNOR2_X1 U436 ( .A(n483), .B(G131), .ZN(n430) );
  XOR2_X1 U437 ( .A(KEYINPUT68), .B(G134), .Z(n483) );
  NAND2_X1 U438 ( .A1(n475), .A2(n474), .ZN(n470) );
  INV_X1 U439 ( .A(KEYINPUT22), .ZN(n601) );
  NOR2_X1 U440 ( .A1(n718), .A2(n636), .ZN(n494) );
  BUF_X1 U441 ( .A(n675), .Z(n421) );
  INV_X1 U442 ( .A(KEYINPUT6), .ZN(n419) );
  INV_X1 U443 ( .A(n712), .ZN(n451) );
  XNOR2_X1 U444 ( .A(n402), .B(n753), .ZN(n724) );
  XNOR2_X1 U445 ( .A(n499), .B(n427), .ZN(n402) );
  XNOR2_X1 U446 ( .A(n498), .B(G146), .ZN(n427) );
  XNOR2_X1 U447 ( .A(n439), .B(n495), .ZN(n499) );
  XOR2_X1 U448 ( .A(KEYINPUT93), .B(n481), .Z(n740) );
  XNOR2_X1 U449 ( .A(n407), .B(n406), .ZN(n405) );
  XNOR2_X1 U450 ( .A(KEYINPUT98), .B(KEYINPUT99), .ZN(n407) );
  XNOR2_X1 U451 ( .A(G116), .B(KEYINPUT5), .ZN(n406) );
  XNOR2_X1 U452 ( .A(n484), .B(n455), .ZN(n480) );
  INV_X1 U453 ( .A(G146), .ZN(n455) );
  INV_X1 U454 ( .A(KEYINPUT97), .ZN(n485) );
  XNOR2_X1 U455 ( .A(G137), .B(G113), .ZN(n486) );
  NAND2_X1 U456 ( .A1(G234), .A2(G237), .ZN(n535) );
  NAND2_X1 U457 ( .A1(n400), .A2(n397), .ZN(n624) );
  AND2_X1 U458 ( .A1(n612), .A2(n398), .ZN(n397) );
  OR2_X1 U459 ( .A1(n764), .A2(KEYINPUT90), .ZN(n400) );
  NAND2_X1 U460 ( .A1(n675), .A2(n459), .ZN(n547) );
  NOR2_X1 U461 ( .A1(n674), .A2(n460), .ZN(n459) );
  XOR2_X1 U462 ( .A(KEYINPUT28), .B(KEYINPUT111), .Z(n551) );
  OR2_X1 U463 ( .A1(G237), .A2(G902), .ZN(n542) );
  NOR2_X1 U464 ( .A1(n675), .A2(n674), .ZN(n670) );
  INV_X1 U465 ( .A(KEYINPUT0), .ZN(n435) );
  NAND2_X2 U466 ( .A1(n466), .A2(n464), .ZN(n404) );
  AND2_X1 U467 ( .A1(n446), .A2(n467), .ZN(n466) );
  OR2_X1 U468 ( .A1(n468), .A2(KEYINPUT87), .ZN(n465) );
  XNOR2_X1 U469 ( .A(KEYINPUT104), .B(KEYINPUT7), .ZN(n433) );
  XOR2_X1 U470 ( .A(G134), .B(KEYINPUT9), .Z(n518) );
  INV_X1 U471 ( .A(KEYINPUT102), .ZN(n390) );
  XNOR2_X1 U472 ( .A(G143), .B(G122), .ZN(n505) );
  XOR2_X1 U473 ( .A(KEYINPUT11), .B(G140), .Z(n506) );
  NAND2_X1 U474 ( .A1(n638), .A2(n368), .ZN(n449) );
  XNOR2_X1 U475 ( .A(n522), .B(n364), .ZN(n439) );
  XNOR2_X1 U476 ( .A(n497), .B(n496), .ZN(n498) );
  INV_X1 U477 ( .A(G101), .ZN(n496) );
  XNOR2_X1 U478 ( .A(KEYINPUT4), .B(KEYINPUT64), .ZN(n482) );
  XNOR2_X1 U479 ( .A(n418), .B(n387), .ZN(n386) );
  XNOR2_X1 U480 ( .A(KEYINPUT18), .B(KEYINPUT75), .ZN(n387) );
  XNOR2_X1 U481 ( .A(n489), .B(KEYINPUT17), .ZN(n384) );
  XNOR2_X1 U482 ( .A(n417), .B(G110), .ZN(n495) );
  INV_X1 U483 ( .A(KEYINPUT69), .ZN(n417) );
  XNOR2_X1 U484 ( .A(n425), .B(n403), .ZN(n747) );
  XNOR2_X1 U485 ( .A(n441), .B(KEYINPUT16), .ZN(n425) );
  NAND2_X1 U486 ( .A1(n613), .A2(n603), .ZN(n401) );
  XNOR2_X1 U487 ( .A(n432), .B(n431), .ZN(n569) );
  INV_X1 U488 ( .A(G478), .ZN(n431) );
  OR2_X1 U489 ( .A1(n724), .A2(G902), .ZN(n426) );
  BUF_X1 U490 ( .A(n670), .Z(n414) );
  XNOR2_X1 U491 ( .A(n463), .B(n369), .ZN(n462) );
  NAND2_X1 U492 ( .A1(n734), .A2(G472), .ZN(n463) );
  INV_X1 U493 ( .A(n740), .ZN(n461) );
  XNOR2_X1 U494 ( .A(n458), .B(n457), .ZN(n456) );
  NAND2_X1 U495 ( .A1(n525), .A2(G221), .ZN(n457) );
  XNOR2_X1 U496 ( .A(n415), .B(n524), .ZN(n458) );
  XNOR2_X1 U497 ( .A(n376), .B(n747), .ZN(n718) );
  XNOR2_X1 U498 ( .A(n385), .B(n383), .ZN(n376) );
  XNOR2_X1 U499 ( .A(n384), .B(n495), .ZN(n383) );
  XNOR2_X1 U500 ( .A(n488), .B(n386), .ZN(n385) );
  XNOR2_X1 U501 ( .A(n424), .B(n367), .ZN(n543) );
  NAND2_X1 U502 ( .A1(n565), .A2(n356), .ZN(n424) );
  XNOR2_X1 U503 ( .A(n375), .B(n374), .ZN(n768) );
  INV_X1 U504 ( .A(KEYINPUT42), .ZN(n374) );
  XNOR2_X1 U505 ( .A(n479), .B(n478), .ZN(n767) );
  INV_X1 U506 ( .A(KEYINPUT40), .ZN(n478) );
  AND2_X1 U507 ( .A1(n477), .A2(n472), .ZN(n471) );
  XNOR2_X1 U508 ( .A(n393), .B(n392), .ZN(n391) );
  INV_X1 U509 ( .A(KEYINPUT36), .ZN(n392) );
  AND2_X1 U510 ( .A1(n475), .A2(n381), .ZN(n572) );
  INV_X1 U511 ( .A(n608), .ZN(n381) );
  NAND2_X1 U512 ( .A1(n389), .A2(n421), .ZN(n388) );
  INV_X1 U513 ( .A(n621), .ZN(n389) );
  OR2_X1 U514 ( .A1(n613), .A2(n421), .ZN(n399) );
  XNOR2_X1 U515 ( .A(n722), .B(n442), .ZN(n725) );
  XNOR2_X1 U516 ( .A(n724), .B(n723), .ZN(n442) );
  NOR2_X1 U517 ( .A1(n669), .A2(n544), .ZN(n356) );
  AND2_X1 U518 ( .A1(n638), .A2(KEYINPUT65), .ZN(n357) );
  XOR2_X1 U519 ( .A(G472), .B(KEYINPUT71), .Z(n358) );
  XOR2_X1 U520 ( .A(G131), .B(KEYINPUT12), .Z(n359) );
  AND2_X1 U521 ( .A1(G214), .A2(n507), .ZN(n360) );
  NOR2_X1 U522 ( .A1(n582), .A2(n667), .ZN(n361) );
  AND2_X1 U523 ( .A1(n477), .A2(n476), .ZN(n363) );
  XOR2_X1 U524 ( .A(G104), .B(G107), .Z(n364) );
  XOR2_X1 U525 ( .A(n563), .B(KEYINPUT39), .Z(n365) );
  XOR2_X1 U526 ( .A(KEYINPUT91), .B(KEYINPUT33), .Z(n366) );
  XOR2_X1 U527 ( .A(KEYINPUT43), .B(KEYINPUT108), .Z(n367) );
  OR2_X2 U528 ( .A1(n620), .A2(n388), .ZN(n649) );
  OR2_X1 U529 ( .A1(n636), .A2(n453), .ZN(n368) );
  XOR2_X1 U530 ( .A(n500), .B(KEYINPUT62), .Z(n369) );
  OR2_X1 U531 ( .A1(n638), .A2(n453), .ZN(n370) );
  INV_X1 U532 ( .A(KEYINPUT65), .ZN(n453) );
  NAND2_X1 U533 ( .A1(n636), .A2(n453), .ZN(n371) );
  AND2_X1 U534 ( .A1(n370), .A2(n449), .ZN(n372) );
  XOR2_X1 U535 ( .A(n642), .B(KEYINPUT92), .Z(n373) );
  NAND2_X1 U536 ( .A1(n391), .A2(n669), .ZN(n665) );
  NAND2_X1 U537 ( .A1(n668), .A2(n567), .ZN(n375) );
  XNOR2_X2 U538 ( .A(n494), .B(n493), .ZN(n382) );
  NAND2_X1 U539 ( .A1(n377), .A2(n689), .ZN(n545) );
  INV_X1 U540 ( .A(n688), .ZN(n377) );
  NAND2_X1 U541 ( .A1(n570), .A2(n571), .ZN(n688) );
  XNOR2_X2 U542 ( .A(n488), .B(n430), .ZN(n753) );
  NAND2_X1 U543 ( .A1(n380), .A2(n365), .ZN(n477) );
  NAND2_X1 U544 ( .A1(n562), .A2(n561), .ZN(n380) );
  INV_X1 U545 ( .A(n380), .ZN(n475) );
  XNOR2_X1 U546 ( .A(n382), .B(KEYINPUT38), .ZN(n686) );
  NAND2_X1 U547 ( .A1(n572), .A2(n382), .ZN(n653) );
  NOR2_X1 U548 ( .A1(n543), .A2(n382), .ZN(n667) );
  NAND2_X1 U549 ( .A1(n618), .A2(n602), .ZN(n620) );
  XNOR2_X1 U550 ( .A(n441), .B(n390), .ZN(n502) );
  NAND2_X1 U551 ( .A1(n395), .A2(n394), .ZN(n393) );
  INV_X1 U552 ( .A(n566), .ZN(n394) );
  XNOR2_X1 U553 ( .A(n565), .B(KEYINPUT112), .ZN(n395) );
  XNOR2_X2 U554 ( .A(n396), .B(n511), .ZN(n571) );
  XNOR2_X2 U555 ( .A(n611), .B(KEYINPUT35), .ZN(n764) );
  XNOR2_X1 U556 ( .A(n491), .B(n512), .ZN(n403) );
  NOR2_X1 U557 ( .A1(n404), .A2(n707), .ZN(n706) );
  XNOR2_X2 U558 ( .A(n404), .B(KEYINPUT73), .ZN(n635) );
  XNOR2_X1 U559 ( .A(n404), .B(KEYINPUT125), .ZN(n759) );
  XNOR2_X1 U560 ( .A(n564), .B(KEYINPUT46), .ZN(n413) );
  XNOR2_X2 U561 ( .A(n412), .B(KEYINPUT48), .ZN(n582) );
  XNOR2_X1 U562 ( .A(n434), .B(KEYINPUT78), .ZN(n654) );
  NAND2_X1 U563 ( .A1(n604), .A2(n600), .ZN(n416) );
  NAND2_X1 U564 ( .A1(n649), .A2(n765), .ZN(n628) );
  XNOR2_X2 U565 ( .A(n619), .B(KEYINPUT32), .ZN(n765) );
  XNOR2_X2 U566 ( .A(n673), .B(n419), .ZN(n613) );
  NOR2_X1 U567 ( .A1(n686), .A2(n545), .ZN(n546) );
  XNOR2_X1 U568 ( .A(n502), .B(n420), .ZN(n504) );
  XNOR2_X1 U569 ( .A(n501), .B(n359), .ZN(n420) );
  XNOR2_X1 U570 ( .A(n560), .B(n559), .ZN(n561) );
  XNOR2_X2 U571 ( .A(n541), .B(KEYINPUT107), .ZN(n565) );
  XNOR2_X2 U572 ( .A(n426), .B(G469), .ZN(n584) );
  OR2_X2 U573 ( .A1(n741), .A2(n371), .ZN(n428) );
  NAND2_X1 U574 ( .A1(n429), .A2(n357), .ZN(n447) );
  NOR2_X1 U575 ( .A1(n732), .A2(G902), .ZN(n432) );
  XNOR2_X1 U576 ( .A(n513), .B(n433), .ZN(n514) );
  NAND2_X1 U577 ( .A1(n567), .A2(n589), .ZN(n434) );
  XNOR2_X2 U578 ( .A(n436), .B(n435), .ZN(n604) );
  NAND2_X1 U579 ( .A1(n622), .A2(n623), .ZN(n437) );
  BUF_X1 U580 ( .A(n654), .Z(n438) );
  INV_X1 U581 ( .A(n669), .ZN(n602) );
  AND2_X2 U582 ( .A1(n631), .A2(n632), .ZN(n634) );
  XNOR2_X1 U583 ( .A(n440), .B(n373), .ZN(G57) );
  NAND2_X1 U584 ( .A1(n462), .A2(n461), .ZN(n440) );
  XNOR2_X1 U585 ( .A(n490), .B(G122), .ZN(n512) );
  XNOR2_X1 U586 ( .A(n443), .B(KEYINPUT122), .ZN(G66) );
  NOR2_X2 U587 ( .A1(n739), .A2(n740), .ZN(n443) );
  XNOR2_X1 U588 ( .A(n444), .B(KEYINPUT56), .ZN(G51) );
  NOR2_X2 U589 ( .A1(n721), .A2(n740), .ZN(n444) );
  XNOR2_X1 U590 ( .A(n445), .B(KEYINPUT60), .ZN(G60) );
  NOR2_X2 U591 ( .A1(n730), .A2(n740), .ZN(n445) );
  NAND2_X1 U592 ( .A1(n582), .A2(KEYINPUT87), .ZN(n446) );
  NAND2_X1 U593 ( .A1(n448), .A2(n447), .ZN(n452) );
  NOR2_X1 U594 ( .A1(n450), .A2(n372), .ZN(n448) );
  INV_X1 U595 ( .A(n421), .ZN(n614) );
  INV_X1 U596 ( .A(n547), .ZN(n549) );
  INV_X1 U597 ( .A(n557), .ZN(n460) );
  INV_X1 U598 ( .A(n667), .ZN(n469) );
  NAND2_X1 U599 ( .A1(n363), .A2(n470), .ZN(n583) );
  NAND2_X1 U600 ( .A1(n471), .A2(n470), .ZN(n479) );
  NOR2_X1 U601 ( .A1(n473), .A2(n657), .ZN(n472) );
  INV_X1 U602 ( .A(n476), .ZN(n473) );
  NOR2_X1 U603 ( .A1(n686), .A2(n365), .ZN(n474) );
  NAND2_X1 U604 ( .A1(n686), .A2(n365), .ZN(n476) );
  XNOR2_X1 U605 ( .A(n729), .B(n728), .ZN(n730) );
  XNOR2_X1 U606 ( .A(n720), .B(n719), .ZN(n721) );
  NOR2_X1 U607 ( .A1(n628), .A2(n764), .ZN(n626) );
  XNOR2_X1 U608 ( .A(n486), .B(n485), .ZN(n487) );
  INV_X1 U609 ( .A(KEYINPUT74), .ZN(n559) );
  XNOR2_X1 U610 ( .A(n508), .B(n360), .ZN(n509) );
  XNOR2_X1 U611 ( .A(n605), .B(KEYINPUT34), .ZN(n606) );
  XNOR2_X1 U612 ( .A(n492), .B(KEYINPUT79), .ZN(n493) );
  XNOR2_X1 U613 ( .A(n738), .B(n737), .ZN(n739) );
  BUF_X1 U614 ( .A(n593), .Z(n669) );
  NOR2_X1 U615 ( .A1(G952), .A2(n760), .ZN(n481) );
  NOR2_X2 U616 ( .A1(G953), .A2(G237), .ZN(n507) );
  NAND2_X1 U617 ( .A1(n507), .A2(G210), .ZN(n484) );
  NAND2_X1 U618 ( .A1(G224), .A2(n760), .ZN(n489) );
  AND2_X1 U619 ( .A1(G210), .A2(n542), .ZN(n492) );
  NAND2_X1 U620 ( .A1(G227), .A2(n760), .ZN(n497) );
  XNOR2_X1 U621 ( .A(KEYINPUT13), .B(G475), .ZN(n511) );
  XOR2_X1 U622 ( .A(KEYINPUT101), .B(KEYINPUT103), .Z(n501) );
  XNOR2_X1 U623 ( .A(n504), .B(n521), .ZN(n510) );
  XNOR2_X1 U624 ( .A(n506), .B(n505), .ZN(n508) );
  XNOR2_X1 U625 ( .A(n512), .B(n514), .ZN(n520) );
  NAND2_X1 U626 ( .A1(n760), .A2(G234), .ZN(n516) );
  XNOR2_X1 U627 ( .A(KEYINPUT67), .B(KEYINPUT8), .ZN(n515) );
  NAND2_X1 U628 ( .A1(G217), .A2(n525), .ZN(n517) );
  XNOR2_X1 U629 ( .A(n518), .B(n517), .ZN(n519) );
  XNOR2_X1 U630 ( .A(n520), .B(n519), .ZN(n732) );
  XOR2_X1 U631 ( .A(KEYINPUT24), .B(G110), .Z(n524) );
  XOR2_X1 U632 ( .A(KEYINPUT96), .B(KEYINPUT25), .Z(n530) );
  INV_X1 U633 ( .A(n636), .ZN(n527) );
  NAND2_X1 U634 ( .A1(n527), .A2(G234), .ZN(n528) );
  XNOR2_X1 U635 ( .A(n528), .B(KEYINPUT20), .ZN(n533) );
  NAND2_X1 U636 ( .A1(n533), .A2(G217), .ZN(n529) );
  XNOR2_X1 U637 ( .A(n530), .B(n529), .ZN(n531) );
  NAND2_X1 U638 ( .A1(G221), .A2(n533), .ZN(n534) );
  XNOR2_X1 U639 ( .A(KEYINPUT21), .B(n534), .ZN(n674) );
  XNOR2_X1 U640 ( .A(n535), .B(KEYINPUT14), .ZN(n537) );
  NAND2_X1 U641 ( .A1(G952), .A2(n537), .ZN(n536) );
  XOR2_X1 U642 ( .A(KEYINPUT94), .B(n536), .Z(n702) );
  NAND2_X1 U643 ( .A1(n760), .A2(n702), .ZN(n587) );
  NAND2_X1 U644 ( .A1(G902), .A2(n537), .ZN(n585) );
  NOR2_X1 U645 ( .A1(G900), .A2(n585), .ZN(n538) );
  NAND2_X1 U646 ( .A1(G953), .A2(n538), .ZN(n539) );
  NAND2_X1 U647 ( .A1(n587), .A2(n539), .ZN(n557) );
  NOR2_X1 U648 ( .A1(n657), .A2(n547), .ZN(n540) );
  NAND2_X1 U649 ( .A1(n613), .A2(n540), .ZN(n541) );
  NAND2_X1 U650 ( .A1(G214), .A2(n542), .ZN(n689) );
  INV_X1 U651 ( .A(n569), .ZN(n570) );
  INV_X1 U652 ( .A(n689), .ZN(n544) );
  XNOR2_X1 U653 ( .A(n546), .B(KEYINPUT41), .ZN(n683) );
  INV_X1 U654 ( .A(n683), .ZN(n668) );
  NAND2_X1 U655 ( .A1(n549), .A2(n621), .ZN(n550) );
  XNOR2_X1 U656 ( .A(n551), .B(n550), .ZN(n554) );
  INV_X1 U657 ( .A(n584), .ZN(n552) );
  XNOR2_X1 U658 ( .A(KEYINPUT110), .B(n552), .ZN(n553) );
  NAND2_X1 U659 ( .A1(n621), .A2(n689), .ZN(n556) );
  XNOR2_X1 U660 ( .A(KEYINPUT30), .B(KEYINPUT109), .ZN(n555) );
  XNOR2_X1 U661 ( .A(n556), .B(n555), .ZN(n562) );
  NAND2_X1 U662 ( .A1(n558), .A2(n584), .ZN(n560) );
  INV_X1 U663 ( .A(KEYINPUT89), .ZN(n563) );
  NAND2_X1 U664 ( .A1(n654), .A2(KEYINPUT47), .ZN(n568) );
  XNOR2_X1 U665 ( .A(n568), .B(KEYINPUT84), .ZN(n576) );
  NAND2_X1 U666 ( .A1(n569), .A2(n571), .ZN(n661) );
  NAND2_X1 U667 ( .A1(n657), .A2(n661), .ZN(n597) );
  INV_X1 U668 ( .A(n597), .ZN(n692) );
  NAND2_X1 U669 ( .A1(KEYINPUT47), .A2(n692), .ZN(n573) );
  OR2_X1 U670 ( .A1(n571), .A2(n570), .ZN(n608) );
  NAND2_X1 U671 ( .A1(n573), .A2(n653), .ZN(n574) );
  XNOR2_X1 U672 ( .A(KEYINPUT81), .B(n574), .ZN(n575) );
  NAND2_X1 U673 ( .A1(n576), .A2(n575), .ZN(n577) );
  NOR2_X1 U674 ( .A1(KEYINPUT47), .A2(n692), .ZN(n578) );
  XNOR2_X1 U675 ( .A(KEYINPUT72), .B(n578), .ZN(n580) );
  INV_X1 U676 ( .A(n438), .ZN(n579) );
  NAND2_X1 U677 ( .A1(n580), .A2(n579), .ZN(n581) );
  OR2_X1 U678 ( .A1(n583), .A2(n661), .ZN(n666) );
  AND2_X1 U679 ( .A1(n414), .A2(n584), .ZN(n592) );
  NOR2_X1 U680 ( .A1(G898), .A2(n760), .ZN(n749) );
  INV_X1 U681 ( .A(n585), .ZN(n586) );
  NAND2_X1 U682 ( .A1(n749), .A2(n586), .ZN(n588) );
  NAND2_X1 U683 ( .A1(n588), .A2(n587), .ZN(n590) );
  INV_X1 U684 ( .A(n604), .ZN(n594) );
  NOR2_X1 U685 ( .A1(n673), .A2(n594), .ZN(n591) );
  NAND2_X1 U686 ( .A1(n592), .A2(n591), .ZN(n645) );
  NAND2_X1 U687 ( .A1(n673), .A2(n603), .ZN(n679) );
  NOR2_X1 U688 ( .A1(n594), .A2(n679), .ZN(n596) );
  XNOR2_X1 U689 ( .A(KEYINPUT100), .B(KEYINPUT31), .ZN(n595) );
  XNOR2_X1 U690 ( .A(n596), .B(n595), .ZN(n662) );
  NAND2_X1 U691 ( .A1(n645), .A2(n662), .ZN(n598) );
  NAND2_X1 U692 ( .A1(n598), .A2(n597), .ZN(n612) );
  OR2_X1 U693 ( .A1(n688), .A2(n674), .ZN(n599) );
  XNOR2_X1 U694 ( .A(n599), .B(KEYINPUT105), .ZN(n600) );
  NAND2_X1 U695 ( .A1(n604), .A2(n695), .ZN(n607) );
  INV_X1 U696 ( .A(KEYINPUT70), .ZN(n605) );
  XNOR2_X1 U697 ( .A(n607), .B(n606), .ZN(n610) );
  XOR2_X1 U698 ( .A(n608), .B(KEYINPUT76), .Z(n609) );
  NAND2_X1 U699 ( .A1(n610), .A2(n609), .ZN(n611) );
  NAND2_X1 U700 ( .A1(n764), .A2(KEYINPUT90), .ZN(n623) );
  NOR2_X1 U701 ( .A1(n614), .A2(n613), .ZN(n615) );
  NAND2_X1 U702 ( .A1(n615), .A2(n669), .ZN(n616) );
  XNOR2_X1 U703 ( .A(n616), .B(KEYINPUT77), .ZN(n617) );
  NAND2_X1 U704 ( .A1(n618), .A2(n617), .ZN(n619) );
  NAND2_X1 U705 ( .A1(KEYINPUT66), .A2(n628), .ZN(n622) );
  NOR2_X1 U706 ( .A1(n624), .A2(n362), .ZN(n632) );
  NAND2_X1 U707 ( .A1(KEYINPUT90), .A2(KEYINPUT66), .ZN(n625) );
  NOR2_X1 U708 ( .A1(n626), .A2(n625), .ZN(n627) );
  NOR2_X1 U709 ( .A1(n627), .A2(KEYINPUT44), .ZN(n630) );
  NOR2_X1 U710 ( .A1(KEYINPUT66), .A2(n628), .ZN(n629) );
  NOR2_X1 U711 ( .A1(n630), .A2(n629), .ZN(n631) );
  XNOR2_X1 U712 ( .A(KEYINPUT88), .B(KEYINPUT45), .ZN(n633) );
  XNOR2_X2 U713 ( .A(n634), .B(n633), .ZN(n741) );
  XNOR2_X1 U714 ( .A(n636), .B(KEYINPUT86), .ZN(n637) );
  NAND2_X1 U715 ( .A1(n637), .A2(KEYINPUT2), .ZN(n638) );
  NAND2_X1 U716 ( .A1(KEYINPUT2), .A2(n666), .ZN(n639) );
  XOR2_X1 U717 ( .A(KEYINPUT80), .B(n639), .Z(n640) );
  NAND2_X1 U718 ( .A1(n361), .A2(n640), .ZN(n641) );
  NOR2_X1 U719 ( .A1(n741), .A2(n641), .ZN(n712) );
  INV_X1 U720 ( .A(KEYINPUT63), .ZN(n642) );
  XOR2_X1 U721 ( .A(G101), .B(n643), .Z(G3) );
  NOR2_X1 U722 ( .A1(n657), .A2(n645), .ZN(n644) );
  XOR2_X1 U723 ( .A(G104), .B(n644), .Z(G6) );
  NOR2_X1 U724 ( .A1(n661), .A2(n645), .ZN(n647) );
  XNOR2_X1 U725 ( .A(KEYINPUT27), .B(KEYINPUT26), .ZN(n646) );
  XNOR2_X1 U726 ( .A(n647), .B(n646), .ZN(n648) );
  XNOR2_X1 U727 ( .A(G107), .B(n648), .ZN(G9) );
  XNOR2_X1 U728 ( .A(G110), .B(n649), .ZN(G12) );
  XOR2_X1 U729 ( .A(G128), .B(KEYINPUT29), .Z(n651) );
  OR2_X1 U730 ( .A1(n661), .A2(n438), .ZN(n650) );
  XNOR2_X1 U731 ( .A(n651), .B(n650), .ZN(G30) );
  XOR2_X1 U732 ( .A(G143), .B(KEYINPUT113), .Z(n652) );
  XNOR2_X1 U733 ( .A(n653), .B(n652), .ZN(G45) );
  NOR2_X1 U734 ( .A1(n438), .A2(n657), .ZN(n655) );
  XOR2_X1 U735 ( .A(KEYINPUT114), .B(n655), .Z(n656) );
  XNOR2_X1 U736 ( .A(G146), .B(n656), .ZN(G48) );
  NOR2_X1 U737 ( .A1(n662), .A2(n657), .ZN(n659) );
  XNOR2_X1 U738 ( .A(KEYINPUT115), .B(KEYINPUT116), .ZN(n658) );
  XNOR2_X1 U739 ( .A(n659), .B(n658), .ZN(n660) );
  XNOR2_X1 U740 ( .A(G113), .B(n660), .ZN(G15) );
  NOR2_X1 U741 ( .A1(n662), .A2(n661), .ZN(n663) );
  XOR2_X1 U742 ( .A(G116), .B(n663), .Z(G18) );
  XOR2_X1 U743 ( .A(G125), .B(KEYINPUT37), .Z(n664) );
  XNOR2_X1 U744 ( .A(n665), .B(n664), .ZN(G27) );
  XNOR2_X1 U745 ( .A(G134), .B(n666), .ZN(G36) );
  XOR2_X1 U746 ( .A(G140), .B(n667), .Z(G42) );
  NAND2_X1 U747 ( .A1(n695), .A2(n668), .ZN(n705) );
  XOR2_X1 U748 ( .A(KEYINPUT51), .B(KEYINPUT117), .Z(n682) );
  NOR2_X1 U749 ( .A1(n414), .A2(n669), .ZN(n671) );
  XNOR2_X1 U750 ( .A(n671), .B(KEYINPUT50), .ZN(n672) );
  NOR2_X1 U751 ( .A1(n673), .A2(n672), .ZN(n678) );
  AND2_X1 U752 ( .A1(n421), .A2(n674), .ZN(n676) );
  XNOR2_X1 U753 ( .A(n676), .B(KEYINPUT49), .ZN(n677) );
  NAND2_X1 U754 ( .A1(n678), .A2(n677), .ZN(n680) );
  NAND2_X1 U755 ( .A1(n680), .A2(n679), .ZN(n681) );
  XNOR2_X1 U756 ( .A(n682), .B(n681), .ZN(n684) );
  NOR2_X1 U757 ( .A1(n684), .A2(n683), .ZN(n685) );
  XOR2_X1 U758 ( .A(KEYINPUT118), .B(n685), .Z(n700) );
  INV_X1 U759 ( .A(n686), .ZN(n690) );
  NOR2_X1 U760 ( .A1(n690), .A2(n689), .ZN(n687) );
  NOR2_X1 U761 ( .A1(n688), .A2(n687), .ZN(n694) );
  NAND2_X1 U762 ( .A1(n690), .A2(n689), .ZN(n691) );
  NOR2_X1 U763 ( .A1(n692), .A2(n691), .ZN(n693) );
  NOR2_X1 U764 ( .A1(n694), .A2(n693), .ZN(n697) );
  INV_X1 U765 ( .A(n695), .ZN(n696) );
  NOR2_X1 U766 ( .A1(n697), .A2(n696), .ZN(n698) );
  XNOR2_X1 U767 ( .A(KEYINPUT119), .B(n698), .ZN(n699) );
  NAND2_X1 U768 ( .A1(n700), .A2(n699), .ZN(n701) );
  XNOR2_X1 U769 ( .A(KEYINPUT52), .B(n701), .ZN(n703) );
  NAND2_X1 U770 ( .A1(n703), .A2(n702), .ZN(n704) );
  NAND2_X1 U771 ( .A1(n705), .A2(n704), .ZN(n714) );
  XNOR2_X1 U772 ( .A(KEYINPUT2), .B(KEYINPUT82), .ZN(n707) );
  XNOR2_X1 U773 ( .A(n706), .B(KEYINPUT85), .ZN(n710) );
  INV_X1 U774 ( .A(n707), .ZN(n708) );
  NAND2_X1 U775 ( .A1(n708), .A2(n741), .ZN(n709) );
  NAND2_X1 U776 ( .A1(n710), .A2(n709), .ZN(n711) );
  NOR2_X1 U777 ( .A1(n712), .A2(n711), .ZN(n713) );
  NOR2_X1 U778 ( .A1(n714), .A2(n713), .ZN(n715) );
  NAND2_X1 U779 ( .A1(n760), .A2(n715), .ZN(n716) );
  XOR2_X1 U780 ( .A(KEYINPUT53), .B(n716), .Z(G75) );
  NAND2_X1 U781 ( .A1(n734), .A2(G210), .ZN(n720) );
  XOR2_X1 U782 ( .A(KEYINPUT54), .B(KEYINPUT55), .Z(n717) );
  XOR2_X1 U783 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n723) );
  NAND2_X1 U784 ( .A1(n734), .A2(G469), .ZN(n722) );
  NOR2_X1 U785 ( .A1(n740), .A2(n725), .ZN(G54) );
  NAND2_X1 U786 ( .A1(n734), .A2(G475), .ZN(n729) );
  XOR2_X1 U787 ( .A(KEYINPUT120), .B(KEYINPUT59), .Z(n726) );
  NAND2_X1 U788 ( .A1(G478), .A2(n734), .ZN(n731) );
  XNOR2_X1 U789 ( .A(n732), .B(n731), .ZN(n733) );
  NOR2_X1 U790 ( .A1(n740), .A2(n733), .ZN(G63) );
  NAND2_X1 U791 ( .A1(n734), .A2(G217), .ZN(n738) );
  INV_X1 U792 ( .A(KEYINPUT121), .ZN(n735) );
  NOR2_X1 U793 ( .A1(G953), .A2(n741), .ZN(n742) );
  XNOR2_X1 U794 ( .A(KEYINPUT123), .B(n742), .ZN(n746) );
  NAND2_X1 U795 ( .A1(G953), .A2(G224), .ZN(n743) );
  XNOR2_X1 U796 ( .A(KEYINPUT61), .B(n743), .ZN(n744) );
  NAND2_X1 U797 ( .A1(n744), .A2(G898), .ZN(n745) );
  NAND2_X1 U798 ( .A1(n746), .A2(n745), .ZN(n751) );
  XNOR2_X1 U799 ( .A(n747), .B(G110), .ZN(n748) );
  NOR2_X1 U800 ( .A1(n749), .A2(n748), .ZN(n750) );
  XNOR2_X1 U801 ( .A(n751), .B(n750), .ZN(n752) );
  XNOR2_X1 U802 ( .A(KEYINPUT124), .B(n752), .ZN(G69) );
  XNOR2_X1 U803 ( .A(n753), .B(n754), .ZN(n758) );
  XNOR2_X1 U804 ( .A(G227), .B(n758), .ZN(n755) );
  NAND2_X1 U805 ( .A1(n755), .A2(G900), .ZN(n756) );
  NAND2_X1 U806 ( .A1(n756), .A2(G953), .ZN(n757) );
  XNOR2_X1 U807 ( .A(n757), .B(KEYINPUT126), .ZN(n763) );
  XNOR2_X1 U808 ( .A(n759), .B(n758), .ZN(n761) );
  NAND2_X1 U809 ( .A1(n761), .A2(n760), .ZN(n762) );
  NAND2_X1 U810 ( .A1(n763), .A2(n762), .ZN(G72) );
  XOR2_X1 U811 ( .A(n764), .B(G122), .Z(G24) );
  XOR2_X1 U812 ( .A(n765), .B(G119), .Z(n766) );
  XNOR2_X1 U813 ( .A(KEYINPUT127), .B(n766), .ZN(G21) );
  XOR2_X1 U814 ( .A(n767), .B(G131), .Z(G33) );
  XOR2_X1 U815 ( .A(n768), .B(G137), .Z(G39) );
endmodule

