

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589,
         n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600,
         n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611,
         n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622,
         n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633,
         n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644,
         n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655,
         n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666,
         n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677,
         n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688,
         n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699,
         n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710,
         n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721,
         n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732,
         n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743,
         n744, n745, n746, n747, n748, n749, n750, n751, n752, n753, n754,
         n755, n756, n757, n758, n759, n760, n761, n762, n763, n764, n765,
         n766, n767, n768, n769, n770, n771, n772, n773, n774, n775, n776,
         n777, n778, n779, n780, n781, n782, n783, n784, n785;

  NOR2_X1 U370 ( .A1(n424), .A2(n364), .ZN(n658) );
  AND2_X1 U371 ( .A1(n646), .A2(KEYINPUT44), .ZN(n364) );
  NOR2_X1 U372 ( .A1(n636), .A2(n647), .ZN(n714) );
  XNOR2_X1 U373 ( .A(n770), .B(n540), .ZN(n747) );
  NAND2_X1 U374 ( .A1(n715), .A2(n714), .ZN(n480) );
  INV_X1 U375 ( .A(G953), .ZN(n778) );
  OR2_X1 U376 ( .A1(n471), .A2(n467), .ZN(n348) );
  OR2_X2 U377 ( .A1(n499), .A2(n496), .ZN(n371) );
  OR2_X2 U378 ( .A1(n598), .A2(n445), .ZN(n439) );
  NOR2_X2 U379 ( .A1(n349), .A2(n378), .ZN(n656) );
  XNOR2_X2 U380 ( .A(n605), .B(KEYINPUT1), .ZN(n715) );
  XNOR2_X2 U381 ( .A(n666), .B(n665), .ZN(n668) );
  NOR2_X1 U382 ( .A1(n753), .A2(n757), .ZN(n754) );
  NOR2_X1 U383 ( .A1(n671), .A2(n757), .ZN(n673) );
  NOR2_X1 U384 ( .A1(n744), .A2(n757), .ZN(n436) );
  NAND2_X1 U385 ( .A1(n664), .A2(n663), .ZN(n666) );
  AND2_X1 U386 ( .A1(n629), .A2(n628), .ZN(n776) );
  NOR2_X1 U387 ( .A1(n785), .A2(n783), .ZN(n618) );
  AND2_X1 U388 ( .A1(n470), .A2(n348), .ZN(n469) );
  OR2_X1 U389 ( .A1(n695), .A2(n677), .ZN(n403) );
  XNOR2_X1 U390 ( .A(n406), .B(n405), .ZN(n782) );
  INV_X1 U391 ( .A(n474), .ZN(n473) );
  OR2_X1 U392 ( .A1(n712), .A2(n477), .ZN(n476) );
  AND2_X1 U393 ( .A1(n355), .A2(n426), .ZN(n615) );
  XNOR2_X1 U394 ( .A(n432), .B(n431), .ZN(n653) );
  NOR2_X1 U395 ( .A1(n633), .A2(n634), .ZN(n432) );
  XNOR2_X1 U396 ( .A(n603), .B(n358), .ZN(n633) );
  XNOR2_X1 U397 ( .A(n394), .B(n429), .ZN(n694) );
  XNOR2_X1 U398 ( .A(n741), .B(n740), .ZN(n742) );
  XNOR2_X1 U399 ( .A(n533), .B(G472), .ZN(n649) );
  XOR2_X1 U400 ( .A(n750), .B(KEYINPUT59), .Z(n752) );
  XNOR2_X1 U401 ( .A(n495), .B(n494), .ZN(n546) );
  XNOR2_X1 U402 ( .A(n536), .B(G110), .ZN(n759) );
  XNOR2_X1 U403 ( .A(n526), .B(G101), .ZN(n495) );
  INV_X1 U404 ( .A(G953), .ZN(n350) );
  XOR2_X1 U405 ( .A(G137), .B(G140), .Z(n535) );
  NOR2_X1 U406 ( .A1(n613), .A2(n732), .ZN(n614) );
  XNOR2_X1 U407 ( .A(n614), .B(KEYINPUT42), .ZN(n785) );
  NAND2_X1 U408 ( .A1(n470), .A2(n348), .ZN(n349) );
  AND2_X1 U409 ( .A1(n350), .A2(n351), .ZN(n738) );
  XNOR2_X1 U410 ( .A(KEYINPUT121), .B(n737), .ZN(n351) );
  NOR2_X1 U411 ( .A1(n668), .A2(n667), .ZN(n352) );
  NOR2_X2 U412 ( .A1(n668), .A2(n667), .ZN(n353) );
  XNOR2_X1 U413 ( .A(n480), .B(n391), .ZN(n354) );
  NOR2_X2 U414 ( .A1(n668), .A2(n667), .ZN(n755) );
  XNOR2_X1 U415 ( .A(G134), .B(G131), .ZN(n530) );
  XNOR2_X1 U416 ( .A(G113), .B(G119), .ZN(n494) );
  XNOR2_X1 U417 ( .A(G146), .B(G125), .ZN(n550) );
  XNOR2_X1 U418 ( .A(n611), .B(KEYINPUT108), .ZN(n707) );
  NAND2_X1 U419 ( .A1(n475), .A2(n635), .ZN(n474) );
  AND2_X1 U420 ( .A1(n452), .A2(n356), .ZN(n454) );
  NAND2_X1 U421 ( .A1(n613), .A2(n359), .ZN(n452) );
  NAND2_X1 U422 ( .A1(n487), .A2(n456), .ZN(n455) );
  NOR2_X1 U423 ( .A1(n687), .A2(n589), .ZN(n599) );
  NOR2_X1 U424 ( .A1(n595), .A2(n594), .ZN(n597) );
  NAND2_X1 U425 ( .A1(n542), .A2(n411), .ZN(n410) );
  INV_X1 U426 ( .A(G902), .ZN(n411) );
  NOR2_X1 U427 ( .A1(n691), .A2(n694), .ZN(n709) );
  XNOR2_X1 U428 ( .A(n527), .B(KEYINPUT5), .ZN(n399) );
  XNOR2_X1 U429 ( .A(G137), .B(G146), .ZN(n527) );
  XNOR2_X1 U430 ( .A(n437), .B(KEYINPUT110), .ZN(n424) );
  NAND2_X1 U431 ( .A1(n404), .A2(n401), .ZN(n437) );
  NAND2_X1 U432 ( .A1(n403), .A2(n402), .ZN(n401) );
  INV_X1 U433 ( .A(n782), .ZN(n404) );
  XNOR2_X1 U434 ( .A(n418), .B(n509), .ZN(n561) );
  XNOR2_X1 U435 ( .A(n508), .B(n419), .ZN(n418) );
  INV_X1 U436 ( .A(KEYINPUT83), .ZN(n419) );
  NOR2_X1 U437 ( .A1(G953), .A2(G237), .ZN(n531) );
  INV_X1 U438 ( .A(KEYINPUT4), .ZN(n529) );
  XNOR2_X1 U439 ( .A(n759), .B(KEYINPUT72), .ZN(n553) );
  XNOR2_X1 U440 ( .A(n551), .B(n550), .ZN(n422) );
  INV_X1 U441 ( .A(KEYINPUT115), .ZN(n434) );
  XOR2_X1 U442 ( .A(n586), .B(n585), .Z(n609) );
  NOR2_X1 U443 ( .A1(n750), .A2(G902), .ZN(n586) );
  XNOR2_X1 U444 ( .A(G122), .B(KEYINPUT16), .ZN(n545) );
  XNOR2_X1 U445 ( .A(n493), .B(n492), .ZN(n505) );
  XNOR2_X1 U446 ( .A(KEYINPUT94), .B(KEYINPUT93), .ZN(n493) );
  XNOR2_X1 U447 ( .A(G110), .B(KEYINPUT24), .ZN(n492) );
  XNOR2_X1 U448 ( .A(G143), .B(G122), .ZN(n579) );
  INV_X1 U449 ( .A(G131), .ZN(n578) );
  XNOR2_X1 U450 ( .A(G104), .B(KEYINPUT101), .ZN(n572) );
  XNOR2_X1 U451 ( .A(n550), .B(KEYINPUT10), .ZN(n771) );
  AND2_X1 U452 ( .A1(n654), .A2(n427), .ZN(n426) );
  INV_X1 U453 ( .A(n592), .ZN(n427) );
  XNOR2_X1 U454 ( .A(n513), .B(n512), .ZN(n514) );
  NOR2_X1 U455 ( .A1(n670), .A2(G902), .ZN(n515) );
  XNOR2_X1 U456 ( .A(n609), .B(n395), .ZN(n587) );
  INV_X1 U457 ( .A(KEYINPUT106), .ZN(n395) );
  XNOR2_X1 U458 ( .A(n425), .B(G478), .ZN(n610) );
  NOR2_X1 U459 ( .A1(n756), .A2(G902), .ZN(n425) );
  INV_X1 U460 ( .A(KEYINPUT6), .ZN(n396) );
  NAND2_X1 U461 ( .A1(n370), .A2(n473), .ZN(n372) );
  INV_X1 U462 ( .A(KEYINPUT47), .ZN(n456) );
  NAND2_X1 U463 ( .A1(n458), .A2(n359), .ZN(n457) );
  INV_X1 U464 ( .A(n488), .ZN(n458) );
  INV_X1 U465 ( .A(n698), .ZN(n442) );
  INV_X1 U466 ( .A(KEYINPUT44), .ZN(n379) );
  INV_X1 U467 ( .A(n709), .ZN(n402) );
  XNOR2_X1 U468 ( .A(G902), .B(KEYINPUT15), .ZN(n557) );
  OR2_X1 U469 ( .A1(G902), .A2(G237), .ZN(n560) );
  NAND2_X1 U470 ( .A1(n415), .A2(G902), .ZN(n413) );
  INV_X1 U471 ( .A(KEYINPUT73), .ZN(n462) );
  XNOR2_X1 U472 ( .A(G116), .B(G107), .ZN(n562) );
  XOR2_X1 U473 ( .A(KEYINPUT9), .B(KEYINPUT7), .Z(n563) );
  XOR2_X1 U474 ( .A(KEYINPUT11), .B(KEYINPUT102), .Z(n575) );
  XNOR2_X1 U475 ( .A(G140), .B(G113), .ZN(n574) );
  XOR2_X1 U476 ( .A(KEYINPUT12), .B(KEYINPUT103), .Z(n573) );
  XOR2_X1 U477 ( .A(G146), .B(G101), .Z(n538) );
  NAND2_X1 U478 ( .A1(G237), .A2(G234), .ZN(n516) );
  INV_X1 U479 ( .A(KEYINPUT38), .ZN(n433) );
  XNOR2_X1 U480 ( .A(n650), .B(KEYINPUT99), .ZN(n723) );
  INV_X1 U481 ( .A(KEYINPUT0), .ZN(n431) );
  XNOR2_X1 U482 ( .A(n399), .B(n528), .ZN(n398) );
  XNOR2_X1 U483 ( .A(n549), .B(n422), .ZN(n552) );
  INV_X1 U484 ( .A(KEYINPUT33), .ZN(n386) );
  OR2_X1 U485 ( .A1(n544), .A2(n543), .ZN(n613) );
  NOR2_X1 U486 ( .A1(n708), .A2(n707), .ZN(n612) );
  NAND2_X1 U487 ( .A1(n503), .A2(n498), .ZN(n497) );
  INV_X1 U488 ( .A(KEYINPUT32), .ZN(n498) );
  NAND2_X1 U489 ( .A1(n501), .A2(KEYINPUT32), .ZN(n500) );
  INV_X1 U490 ( .A(n503), .ZN(n501) );
  INV_X1 U491 ( .A(n633), .ZN(n488) );
  INV_X1 U492 ( .A(n613), .ZN(n459) );
  XNOR2_X1 U493 ( .A(n490), .B(n489), .ZN(n670) );
  XNOR2_X1 U494 ( .A(n491), .B(n506), .ZN(n490) );
  XNOR2_X1 U495 ( .A(n510), .B(n507), .ZN(n489) );
  XNOR2_X1 U496 ( .A(n392), .B(n393), .ZN(n750) );
  XNOR2_X1 U497 ( .A(n771), .B(n580), .ZN(n393) );
  XNOR2_X1 U498 ( .A(n579), .B(n578), .ZN(n580) );
  XNOR2_X1 U499 ( .A(KEYINPUT84), .B(KEYINPUT2), .ZN(n702) );
  NOR2_X1 U500 ( .A1(n625), .A2(n593), .ZN(n685) );
  INV_X1 U501 ( .A(KEYINPUT107), .ZN(n429) );
  NOR2_X1 U502 ( .A1(n587), .A2(n610), .ZN(n394) );
  INV_X1 U503 ( .A(KEYINPUT109), .ZN(n405) );
  INV_X1 U504 ( .A(KEYINPUT122), .ZN(n481) );
  XNOR2_X1 U505 ( .A(n485), .B(n484), .ZN(n483) );
  XNOR2_X1 U506 ( .A(n745), .B(n420), .ZN(n749) );
  XNOR2_X1 U507 ( .A(n748), .B(n746), .ZN(n420) );
  INV_X1 U508 ( .A(G122), .ZN(n380) );
  INV_X1 U509 ( .A(KEYINPUT89), .ZN(n657) );
  XNOR2_X1 U510 ( .A(n612), .B(KEYINPUT41), .ZN(n732) );
  XNOR2_X1 U511 ( .A(n608), .B(n434), .ZN(n708) );
  XOR2_X1 U512 ( .A(n428), .B(KEYINPUT30), .Z(n355) );
  AND2_X1 U513 ( .A1(n457), .A2(n455), .ZN(n356) );
  AND2_X1 U514 ( .A1(n488), .A2(n487), .ZN(n357) );
  INV_X1 U515 ( .A(KEYINPUT81), .ZN(n487) );
  XOR2_X1 U516 ( .A(KEYINPUT19), .B(KEYINPUT66), .Z(n358) );
  AND2_X1 U517 ( .A1(KEYINPUT81), .A2(KEYINPUT47), .ZN(n359) );
  XNOR2_X1 U518 ( .A(n546), .B(n545), .ZN(n758) );
  XOR2_X1 U519 ( .A(n674), .B(KEYINPUT62), .Z(n360) );
  XOR2_X1 U520 ( .A(n619), .B(KEYINPUT48), .Z(n361) );
  INV_X1 U521 ( .A(KEYINPUT74), .ZN(n448) );
  INV_X1 U522 ( .A(KEYINPUT35), .ZN(n467) );
  XOR2_X1 U523 ( .A(n675), .B(KEYINPUT116), .Z(n362) );
  NOR2_X1 U524 ( .A1(G952), .A2(n778), .ZN(n757) );
  INV_X1 U525 ( .A(n757), .ZN(n482) );
  AND2_X1 U526 ( .A1(n371), .A2(n681), .ZN(n363) );
  INV_X1 U527 ( .A(n605), .ZN(n365) );
  INV_X1 U528 ( .A(n365), .ZN(n366) );
  OR2_X1 U529 ( .A1(n499), .A2(n496), .ZN(n376) );
  OR2_X2 U530 ( .A1(n409), .A2(n412), .ZN(n605) );
  OR2_X1 U531 ( .A1(n712), .A2(n477), .ZN(n370) );
  NAND2_X1 U532 ( .A1(n367), .A2(n370), .ZN(n468) );
  NOR2_X1 U533 ( .A1(n474), .A2(n373), .ZN(n367) );
  AND2_X1 U534 ( .A1(n629), .A2(n368), .ZN(n660) );
  AND2_X1 U535 ( .A1(n628), .A2(n661), .ZN(n368) );
  OR2_X1 U536 ( .A1(n372), .A2(n373), .ZN(n369) );
  NAND2_X1 U537 ( .A1(n376), .A2(n681), .ZN(n382) );
  XNOR2_X1 U538 ( .A(n652), .B(n651), .ZN(n695) );
  NAND2_X1 U539 ( .A1(n414), .A2(n413), .ZN(n412) );
  NAND2_X1 U540 ( .A1(n471), .A2(n467), .ZN(n373) );
  XNOR2_X1 U541 ( .A(n400), .B(n398), .ZN(n397) );
  NAND2_X1 U542 ( .A1(n476), .A2(n473), .ZN(n472) );
  NAND2_X1 U543 ( .A1(n653), .A2(KEYINPUT34), .ZN(n475) );
  BUF_X1 U544 ( .A(n715), .Z(n435) );
  BUF_X1 U545 ( .A(n765), .Z(n374) );
  XNOR2_X1 U546 ( .A(n430), .B(n659), .ZN(n765) );
  NAND2_X1 U547 ( .A1(n353), .A2(G478), .ZN(n485) );
  AND2_X1 U548 ( .A1(n408), .A2(n641), .ZN(n503) );
  INV_X1 U549 ( .A(n408), .ZN(n389) );
  XNOR2_X1 U550 ( .A(n649), .B(n396), .ZN(n408) );
  OR2_X1 U551 ( .A1(n649), .A2(n423), .ZN(n428) );
  BUF_X1 U552 ( .A(n770), .Z(n375) );
  INV_X1 U553 ( .A(n704), .ZN(n423) );
  NAND2_X1 U554 ( .A1(n502), .A2(n500), .ZN(n499) );
  NAND2_X1 U555 ( .A1(n384), .A2(n371), .ZN(n383) );
  XNOR2_X1 U556 ( .A(n371), .B(G119), .ZN(G21) );
  NAND2_X1 U557 ( .A1(n377), .A2(n389), .ZN(n387) );
  AND2_X1 U558 ( .A1(n354), .A2(n390), .ZN(n650) );
  XNOR2_X1 U559 ( .A(n480), .B(n391), .ZN(n377) );
  NAND2_X1 U560 ( .A1(n469), .A2(n369), .ZN(n381) );
  NAND2_X1 U561 ( .A1(n468), .A2(n379), .ZN(n378) );
  INV_X1 U562 ( .A(n381), .ZN(n421) );
  XNOR2_X1 U563 ( .A(n381), .B(n380), .ZN(G24) );
  NAND2_X1 U564 ( .A1(n382), .A2(KEYINPUT89), .ZN(n385) );
  NAND2_X1 U565 ( .A1(n385), .A2(n383), .ZN(n464) );
  AND2_X1 U566 ( .A1(n681), .A2(n657), .ZN(n384) );
  XNOR2_X2 U567 ( .A(n387), .B(n386), .ZN(n712) );
  NAND2_X1 U568 ( .A1(n388), .A2(n444), .ZN(n446) );
  AND2_X1 U569 ( .A1(n447), .A2(n441), .ZN(n388) );
  INV_X1 U570 ( .A(n649), .ZN(n390) );
  INV_X1 U571 ( .A(KEYINPUT76), .ZN(n391) );
  XNOR2_X1 U572 ( .A(n581), .B(n582), .ZN(n392) );
  NAND2_X1 U573 ( .A1(n601), .A2(n389), .ZN(n602) );
  XNOR2_X1 U574 ( .A(n397), .B(n438), .ZN(n674) );
  XNOR2_X2 U575 ( .A(n554), .B(n530), .ZN(n438) );
  XNOR2_X2 U576 ( .A(n565), .B(n529), .ZN(n554) );
  XNOR2_X1 U577 ( .A(n546), .B(n532), .ZN(n400) );
  NOR2_X1 U578 ( .A1(n643), .A2(n407), .ZN(n406) );
  NAND2_X1 U579 ( .A1(n648), .A2(n408), .ZN(n407) );
  NOR2_X1 U580 ( .A1(n747), .A2(n410), .ZN(n409) );
  NAND2_X1 U581 ( .A1(n747), .A2(n415), .ZN(n414) );
  INV_X1 U582 ( .A(n542), .ZN(n415) );
  XNOR2_X1 U583 ( .A(n416), .B(n481), .ZN(G63) );
  NAND2_X1 U584 ( .A1(n483), .A2(n482), .ZN(n416) );
  XNOR2_X1 U585 ( .A(n751), .B(n752), .ZN(n753) );
  XNOR2_X1 U586 ( .A(n417), .B(KEYINPUT40), .ZN(n783) );
  NOR2_X1 U587 ( .A1(n620), .A2(n688), .ZN(n417) );
  NAND2_X1 U588 ( .A1(n363), .A2(n421), .ZN(n646) );
  XNOR2_X2 U589 ( .A(n438), .B(n535), .ZN(n770) );
  XNOR2_X1 U590 ( .A(n463), .B(n462), .ZN(n461) );
  NOR2_X1 U591 ( .A1(n443), .A2(n442), .ZN(n441) );
  NAND2_X1 U592 ( .A1(n461), .A2(n658), .ZN(n430) );
  XNOR2_X1 U593 ( .A(n446), .B(n361), .ZN(n629) );
  XNOR2_X2 U594 ( .A(n607), .B(n433), .ZN(n705) );
  NAND2_X1 U595 ( .A1(n765), .A2(n660), .ZN(n664) );
  XNOR2_X1 U596 ( .A(n436), .B(KEYINPUT56), .ZN(G51) );
  NAND2_X1 U597 ( .A1(n440), .A2(n439), .ZN(n444) );
  NAND2_X1 U598 ( .A1(n598), .A2(n448), .ZN(n440) );
  AND2_X1 U599 ( .A1(n599), .A2(KEYINPUT74), .ZN(n443) );
  NOR2_X1 U600 ( .A1(n599), .A2(KEYINPUT74), .ZN(n445) );
  XNOR2_X1 U601 ( .A(n618), .B(KEYINPUT46), .ZN(n447) );
  XNOR2_X1 U602 ( .A(n449), .B(n362), .ZN(G57) );
  NAND2_X1 U603 ( .A1(n450), .A2(n482), .ZN(n449) );
  XNOR2_X1 U604 ( .A(n451), .B(n360), .ZN(n450) );
  NAND2_X1 U605 ( .A1(n352), .A2(G472), .ZN(n451) );
  NAND2_X1 U606 ( .A1(n459), .A2(n488), .ZN(n687) );
  NAND2_X1 U607 ( .A1(n454), .A2(n453), .ZN(n486) );
  NAND2_X1 U608 ( .A1(n459), .A2(n357), .ZN(n453) );
  XNOR2_X2 U609 ( .A(n460), .B(G143), .ZN(n565) );
  XNOR2_X2 U610 ( .A(G128), .B(KEYINPUT79), .ZN(n460) );
  NAND2_X1 U611 ( .A1(n465), .A2(n464), .ZN(n463) );
  XNOR2_X1 U612 ( .A(n656), .B(n466), .ZN(n465) );
  INV_X1 U613 ( .A(KEYINPUT67), .ZN(n466) );
  NAND2_X1 U614 ( .A1(n712), .A2(KEYINPUT34), .ZN(n471) );
  NAND2_X1 U615 ( .A1(n472), .A2(KEYINPUT35), .ZN(n470) );
  NAND2_X1 U616 ( .A1(n478), .A2(n479), .ZN(n477) );
  INV_X1 U617 ( .A(n653), .ZN(n478) );
  INV_X1 U618 ( .A(KEYINPUT34), .ZN(n479) );
  INV_X1 U619 ( .A(n756), .ZN(n484) );
  NAND2_X1 U620 ( .A1(n705), .A2(n704), .ZN(n608) );
  BUF_X2 U621 ( .A(n591), .Z(n607) );
  NAND2_X1 U622 ( .A1(n590), .A2(n486), .ZN(n595) );
  NAND2_X1 U623 ( .A1(n561), .A2(G221), .ZN(n491) );
  NAND2_X1 U624 ( .A1(n643), .A2(KEYINPUT32), .ZN(n502) );
  XNOR2_X2 U625 ( .A(n640), .B(n639), .ZN(n643) );
  NOR2_X1 U626 ( .A1(n643), .A2(n497), .ZN(n496) );
  NAND2_X1 U627 ( .A1(n591), .A2(n704), .ZN(n603) );
  XNOR2_X1 U628 ( .A(n703), .B(n702), .ZN(n736) );
  AND2_X2 U629 ( .A1(KEYINPUT2), .A2(n703), .ZN(n667) );
  XNOR2_X1 U630 ( .A(n505), .B(KEYINPUT78), .ZN(n506) );
  XNOR2_X1 U631 ( .A(n743), .B(n742), .ZN(n744) );
  INV_X1 U632 ( .A(KEYINPUT80), .ZN(n596) );
  XNOR2_X1 U633 ( .A(n597), .B(n596), .ZN(n598) );
  XNOR2_X1 U634 ( .A(n541), .B(G469), .ZN(n542) );
  XNOR2_X1 U635 ( .A(n553), .B(n539), .ZN(n540) );
  INV_X1 U636 ( .A(KEYINPUT123), .ZN(n672) );
  XNOR2_X1 U637 ( .A(G128), .B(n535), .ZN(n504) );
  XNOR2_X1 U638 ( .A(n504), .B(G119), .ZN(n510) );
  XNOR2_X1 U639 ( .A(n771), .B(KEYINPUT23), .ZN(n507) );
  XOR2_X1 U640 ( .A(KEYINPUT8), .B(KEYINPUT68), .Z(n509) );
  NAND2_X1 U641 ( .A1(G234), .A2(n778), .ZN(n508) );
  NAND2_X1 U642 ( .A1(G234), .A2(n557), .ZN(n511) );
  XNOR2_X1 U643 ( .A(KEYINPUT20), .B(n511), .ZN(n522) );
  NAND2_X1 U644 ( .A1(G217), .A2(n522), .ZN(n513) );
  XNOR2_X1 U645 ( .A(KEYINPUT95), .B(KEYINPUT25), .ZN(n512) );
  XNOR2_X2 U646 ( .A(n515), .B(n514), .ZN(n647) );
  XNOR2_X1 U647 ( .A(n516), .B(KEYINPUT14), .ZN(n517) );
  NAND2_X1 U648 ( .A1(G952), .A2(n517), .ZN(n731) );
  NOR2_X1 U649 ( .A1(G953), .A2(n731), .ZN(n632) );
  NAND2_X1 U650 ( .A1(G902), .A2(n517), .ZN(n518) );
  XOR2_X1 U651 ( .A(KEYINPUT92), .B(n518), .Z(n519) );
  NAND2_X1 U652 ( .A1(G953), .A2(n519), .ZN(n630) );
  NOR2_X1 U653 ( .A1(G900), .A2(n630), .ZN(n520) );
  XOR2_X1 U654 ( .A(KEYINPUT111), .B(n520), .Z(n521) );
  NOR2_X1 U655 ( .A1(n632), .A2(n521), .ZN(n592) );
  NAND2_X1 U656 ( .A1(n522), .A2(G221), .ZN(n523) );
  XOR2_X1 U657 ( .A(KEYINPUT21), .B(n523), .Z(n524) );
  XOR2_X1 U658 ( .A(KEYINPUT96), .B(n524), .Z(n636) );
  NOR2_X1 U659 ( .A1(n592), .A2(n636), .ZN(n525) );
  NAND2_X1 U660 ( .A1(n647), .A2(n525), .ZN(n600) );
  XNOR2_X2 U661 ( .A(G116), .B(KEYINPUT3), .ZN(n526) );
  XOR2_X1 U662 ( .A(KEYINPUT98), .B(KEYINPUT97), .Z(n528) );
  XOR2_X1 U663 ( .A(KEYINPUT77), .B(n531), .Z(n571) );
  NAND2_X1 U664 ( .A1(n571), .A2(G210), .ZN(n532) );
  NOR2_X1 U665 ( .A1(G902), .A2(n674), .ZN(n533) );
  NOR2_X1 U666 ( .A1(n600), .A2(n649), .ZN(n534) );
  XOR2_X1 U667 ( .A(KEYINPUT28), .B(n534), .Z(n544) );
  XOR2_X1 U668 ( .A(G107), .B(G104), .Z(n536) );
  NAND2_X1 U669 ( .A1(G227), .A2(n778), .ZN(n537) );
  XNOR2_X1 U670 ( .A(n538), .B(n537), .ZN(n539) );
  XNOR2_X1 U671 ( .A(KEYINPUT70), .B(KEYINPUT71), .ZN(n541) );
  XOR2_X1 U672 ( .A(n366), .B(KEYINPUT114), .Z(n543) );
  XOR2_X1 U673 ( .A(KEYINPUT18), .B(KEYINPUT90), .Z(n548) );
  XNOR2_X1 U674 ( .A(KEYINPUT17), .B(KEYINPUT91), .ZN(n547) );
  XNOR2_X1 U675 ( .A(n548), .B(n547), .ZN(n549) );
  NAND2_X1 U676 ( .A1(G224), .A2(n778), .ZN(n551) );
  XNOR2_X1 U677 ( .A(n758), .B(n552), .ZN(n556) );
  XOR2_X1 U678 ( .A(n554), .B(n553), .Z(n555) );
  XNOR2_X1 U679 ( .A(n556), .B(n555), .ZN(n739) );
  INV_X1 U680 ( .A(n557), .ZN(n661) );
  NOR2_X2 U681 ( .A1(n739), .A2(n661), .ZN(n559) );
  NAND2_X1 U682 ( .A1(G210), .A2(n560), .ZN(n558) );
  XNOR2_X2 U683 ( .A(n559), .B(n558), .ZN(n591) );
  NAND2_X1 U684 ( .A1(G214), .A2(n560), .ZN(n704) );
  NAND2_X1 U685 ( .A1(n561), .A2(G217), .ZN(n570) );
  XNOR2_X1 U686 ( .A(n563), .B(n562), .ZN(n564) );
  XOR2_X1 U687 ( .A(n564), .B(G134), .Z(n568) );
  INV_X1 U688 ( .A(n565), .ZN(n566) );
  XOR2_X1 U689 ( .A(n566), .B(G122), .Z(n567) );
  XNOR2_X1 U690 ( .A(n567), .B(n568), .ZN(n569) );
  XOR2_X1 U691 ( .A(n570), .B(n569), .Z(n756) );
  NAND2_X1 U692 ( .A1(n571), .A2(G214), .ZN(n582) );
  XNOR2_X1 U693 ( .A(n573), .B(n572), .ZN(n577) );
  XNOR2_X1 U694 ( .A(n575), .B(n574), .ZN(n576) );
  XNOR2_X1 U695 ( .A(n577), .B(n576), .ZN(n581) );
  XOR2_X1 U696 ( .A(KEYINPUT105), .B(KEYINPUT104), .Z(n584) );
  XNOR2_X1 U697 ( .A(KEYINPUT13), .B(G475), .ZN(n583) );
  XNOR2_X1 U698 ( .A(n584), .B(n583), .ZN(n585) );
  NAND2_X1 U699 ( .A1(n610), .A2(n587), .ZN(n688) );
  INV_X1 U700 ( .A(n688), .ZN(n691) );
  NOR2_X1 U701 ( .A1(n709), .A2(KEYINPUT47), .ZN(n588) );
  XNOR2_X1 U702 ( .A(n588), .B(KEYINPUT75), .ZN(n589) );
  NAND2_X1 U703 ( .A1(n709), .A2(KEYINPUT47), .ZN(n590) );
  INV_X1 U704 ( .A(n607), .ZN(n625) );
  AND2_X1 U705 ( .A1(n366), .A2(n714), .ZN(n654) );
  NOR2_X1 U706 ( .A1(n609), .A2(n610), .ZN(n635) );
  NAND2_X1 U707 ( .A1(n615), .A2(n635), .ZN(n593) );
  XNOR2_X1 U708 ( .A(n685), .B(KEYINPUT82), .ZN(n594) );
  NOR2_X1 U709 ( .A1(n688), .A2(n600), .ZN(n601) );
  XNOR2_X1 U710 ( .A(KEYINPUT112), .B(n602), .ZN(n622) );
  NOR2_X1 U711 ( .A1(n622), .A2(n603), .ZN(n604) );
  XNOR2_X1 U712 ( .A(KEYINPUT36), .B(n604), .ZN(n606) );
  NAND2_X1 U713 ( .A1(n606), .A2(n435), .ZN(n698) );
  NAND2_X1 U714 ( .A1(n610), .A2(n609), .ZN(n611) );
  XOR2_X1 U715 ( .A(KEYINPUT88), .B(KEYINPUT39), .Z(n617) );
  NAND2_X1 U716 ( .A1(n615), .A2(n705), .ZN(n616) );
  XNOR2_X1 U717 ( .A(n616), .B(n617), .ZN(n620) );
  XNOR2_X1 U718 ( .A(KEYINPUT87), .B(KEYINPUT69), .ZN(n619) );
  INV_X1 U719 ( .A(n694), .ZN(n682) );
  NOR2_X1 U720 ( .A1(n620), .A2(n682), .ZN(n700) );
  INV_X1 U721 ( .A(n435), .ZN(n644) );
  NAND2_X1 U722 ( .A1(n644), .A2(n704), .ZN(n621) );
  NOR2_X1 U723 ( .A1(n622), .A2(n621), .ZN(n624) );
  XNOR2_X1 U724 ( .A(KEYINPUT113), .B(KEYINPUT43), .ZN(n623) );
  XNOR2_X1 U725 ( .A(n624), .B(n623), .ZN(n626) );
  NAND2_X1 U726 ( .A1(n626), .A2(n625), .ZN(n701) );
  INV_X1 U727 ( .A(n701), .ZN(n627) );
  NOR2_X1 U728 ( .A1(n700), .A2(n627), .ZN(n628) );
  NOR2_X1 U729 ( .A1(G898), .A2(n630), .ZN(n631) );
  NOR2_X1 U730 ( .A1(n632), .A2(n631), .ZN(n634) );
  INV_X1 U731 ( .A(n636), .ZN(n717) );
  INV_X1 U732 ( .A(n707), .ZN(n637) );
  NAND2_X1 U733 ( .A1(n717), .A2(n637), .ZN(n638) );
  NOR2_X1 U734 ( .A1(n653), .A2(n638), .ZN(n640) );
  XNOR2_X1 U735 ( .A(KEYINPUT65), .B(KEYINPUT22), .ZN(n639) );
  INV_X1 U736 ( .A(n647), .ZN(n718) );
  NOR2_X1 U737 ( .A1(n644), .A2(n718), .ZN(n641) );
  NAND2_X1 U738 ( .A1(n647), .A2(n649), .ZN(n642) );
  NOR2_X1 U739 ( .A1(n643), .A2(n642), .ZN(n645) );
  NAND2_X1 U740 ( .A1(n645), .A2(n644), .ZN(n681) );
  NOR2_X1 U741 ( .A1(n435), .A2(n647), .ZN(n648) );
  NOR2_X1 U742 ( .A1(n653), .A2(n723), .ZN(n652) );
  XOR2_X1 U743 ( .A(KEYINPUT100), .B(KEYINPUT31), .Z(n651) );
  NAND2_X1 U744 ( .A1(n654), .A2(n478), .ZN(n655) );
  NOR2_X1 U745 ( .A1(n390), .A2(n655), .ZN(n677) );
  XNOR2_X1 U746 ( .A(KEYINPUT86), .B(KEYINPUT45), .ZN(n659) );
  XOR2_X1 U747 ( .A(n661), .B(KEYINPUT85), .Z(n662) );
  NAND2_X1 U748 ( .A1(n662), .A2(KEYINPUT2), .ZN(n663) );
  INV_X1 U749 ( .A(KEYINPUT64), .ZN(n665) );
  AND2_X1 U750 ( .A1(n765), .A2(n776), .ZN(n703) );
  NAND2_X1 U751 ( .A1(n755), .A2(G217), .ZN(n669) );
  XNOR2_X1 U752 ( .A(n669), .B(n670), .ZN(n671) );
  XNOR2_X1 U753 ( .A(n673), .B(n672), .ZN(G66) );
  INV_X1 U754 ( .A(KEYINPUT63), .ZN(n675) );
  NAND2_X1 U755 ( .A1(n677), .A2(n691), .ZN(n676) );
  XNOR2_X1 U756 ( .A(n676), .B(G104), .ZN(G6) );
  XOR2_X1 U757 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n679) );
  NAND2_X1 U758 ( .A1(n677), .A2(n694), .ZN(n678) );
  XNOR2_X1 U759 ( .A(n679), .B(n678), .ZN(n680) );
  XNOR2_X1 U760 ( .A(G107), .B(n680), .ZN(G9) );
  XNOR2_X1 U761 ( .A(G110), .B(n681), .ZN(G12) );
  NOR2_X1 U762 ( .A1(n687), .A2(n682), .ZN(n684) );
  XNOR2_X1 U763 ( .A(G128), .B(KEYINPUT29), .ZN(n683) );
  XNOR2_X1 U764 ( .A(n684), .B(n683), .ZN(G30) );
  XNOR2_X1 U765 ( .A(G143), .B(n685), .ZN(n686) );
  XNOR2_X1 U766 ( .A(n686), .B(KEYINPUT117), .ZN(G45) );
  NOR2_X1 U767 ( .A1(n688), .A2(n687), .ZN(n689) );
  XOR2_X1 U768 ( .A(KEYINPUT118), .B(n689), .Z(n690) );
  XNOR2_X1 U769 ( .A(G146), .B(n690), .ZN(G48) );
  XOR2_X1 U770 ( .A(G113), .B(KEYINPUT119), .Z(n693) );
  NAND2_X1 U771 ( .A1(n691), .A2(n695), .ZN(n692) );
  XNOR2_X1 U772 ( .A(n693), .B(n692), .ZN(G15) );
  NAND2_X1 U773 ( .A1(n695), .A2(n694), .ZN(n696) );
  XNOR2_X1 U774 ( .A(n696), .B(G116), .ZN(G18) );
  XOR2_X1 U775 ( .A(KEYINPUT37), .B(KEYINPUT120), .Z(n697) );
  XNOR2_X1 U776 ( .A(n698), .B(n697), .ZN(n699) );
  XNOR2_X1 U777 ( .A(G125), .B(n699), .ZN(G27) );
  XOR2_X1 U778 ( .A(G134), .B(n700), .Z(G36) );
  XNOR2_X1 U779 ( .A(G140), .B(n701), .ZN(G42) );
  NOR2_X1 U780 ( .A1(n705), .A2(n704), .ZN(n706) );
  NOR2_X1 U781 ( .A1(n707), .A2(n706), .ZN(n711) );
  NOR2_X1 U782 ( .A1(n709), .A2(n708), .ZN(n710) );
  NOR2_X1 U783 ( .A1(n711), .A2(n710), .ZN(n713) );
  NOR2_X1 U784 ( .A1(n713), .A2(n712), .ZN(n728) );
  OR2_X1 U785 ( .A1(n435), .A2(n714), .ZN(n716) );
  XNOR2_X1 U786 ( .A(n716), .B(KEYINPUT50), .ZN(n722) );
  NOR2_X1 U787 ( .A1(n718), .A2(n717), .ZN(n719) );
  XOR2_X1 U788 ( .A(KEYINPUT49), .B(n719), .Z(n720) );
  NOR2_X1 U789 ( .A1(n390), .A2(n720), .ZN(n721) );
  NAND2_X1 U790 ( .A1(n722), .A2(n721), .ZN(n724) );
  NAND2_X1 U791 ( .A1(n724), .A2(n723), .ZN(n725) );
  XNOR2_X1 U792 ( .A(KEYINPUT51), .B(n725), .ZN(n726) );
  NOR2_X1 U793 ( .A1(n732), .A2(n726), .ZN(n727) );
  NOR2_X1 U794 ( .A1(n728), .A2(n727), .ZN(n729) );
  XNOR2_X1 U795 ( .A(n729), .B(KEYINPUT52), .ZN(n730) );
  NOR2_X1 U796 ( .A1(n731), .A2(n730), .ZN(n734) );
  NOR2_X1 U797 ( .A1(n712), .A2(n732), .ZN(n733) );
  NOR2_X1 U798 ( .A1(n734), .A2(n733), .ZN(n735) );
  NAND2_X1 U799 ( .A1(n736), .A2(n735), .ZN(n737) );
  XNOR2_X1 U800 ( .A(KEYINPUT53), .B(n738), .ZN(G75) );
  NAND2_X1 U801 ( .A1(n353), .A2(G210), .ZN(n743) );
  BUF_X1 U802 ( .A(n739), .Z(n741) );
  XOR2_X1 U803 ( .A(KEYINPUT54), .B(KEYINPUT55), .Z(n740) );
  XOR2_X1 U804 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n746) );
  NAND2_X1 U805 ( .A1(n352), .A2(G469), .ZN(n745) );
  BUF_X1 U806 ( .A(n747), .Z(n748) );
  NOR2_X1 U807 ( .A1(n757), .A2(n749), .ZN(G54) );
  NAND2_X1 U808 ( .A1(n755), .A2(G475), .ZN(n751) );
  XNOR2_X1 U809 ( .A(n754), .B(KEYINPUT60), .ZN(G60) );
  NOR2_X1 U810 ( .A1(G898), .A2(n778), .ZN(n761) );
  XOR2_X1 U811 ( .A(n759), .B(n758), .Z(n760) );
  NOR2_X1 U812 ( .A1(n761), .A2(n760), .ZN(n769) );
  NAND2_X1 U813 ( .A1(G953), .A2(G224), .ZN(n762) );
  XNOR2_X1 U814 ( .A(KEYINPUT61), .B(n762), .ZN(n763) );
  NAND2_X1 U815 ( .A1(n763), .A2(G898), .ZN(n764) );
  XNOR2_X1 U816 ( .A(n764), .B(KEYINPUT124), .ZN(n767) );
  NAND2_X1 U817 ( .A1(n374), .A2(n778), .ZN(n766) );
  NAND2_X1 U818 ( .A1(n767), .A2(n766), .ZN(n768) );
  XNOR2_X1 U819 ( .A(n769), .B(n768), .ZN(G69) );
  XNOR2_X1 U820 ( .A(n375), .B(n771), .ZN(n775) );
  XNOR2_X1 U821 ( .A(G227), .B(n775), .ZN(n772) );
  XNOR2_X1 U822 ( .A(n772), .B(KEYINPUT126), .ZN(n773) );
  NAND2_X1 U823 ( .A1(G900), .A2(n773), .ZN(n774) );
  NAND2_X1 U824 ( .A1(n774), .A2(G953), .ZN(n781) );
  XNOR2_X1 U825 ( .A(n776), .B(n775), .ZN(n777) );
  XNOR2_X1 U826 ( .A(n777), .B(KEYINPUT125), .ZN(n779) );
  NAND2_X1 U827 ( .A1(n779), .A2(n778), .ZN(n780) );
  NAND2_X1 U828 ( .A1(n781), .A2(n780), .ZN(G72) );
  XOR2_X1 U829 ( .A(G101), .B(n782), .Z(G3) );
  XNOR2_X1 U830 ( .A(G131), .B(KEYINPUT127), .ZN(n784) );
  XNOR2_X1 U831 ( .A(n784), .B(n783), .ZN(G33) );
  XOR2_X1 U832 ( .A(n785), .B(G137), .Z(G39) );
endmodule

