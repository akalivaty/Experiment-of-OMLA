

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
         n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706,
         n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717,
         n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
         n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739,
         n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750,
         n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761,
         n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772,
         n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783,
         n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n794,
         n795, n796, n797, n798, n799, n800, n801, n802, n803, n804, n805,
         n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n816,
         n817, n818, n819, n820, n821, n822, n823, n824, n825, n826, n827,
         n828, n829, n830, n831, n832, n833, n834, n835, n836, n837, n838,
         n839, n840, n841, n842, n843, n844, n845, n846, n847, n848, n849,
         n850, n851, n852, n853, n854, n855, n856, n857, n858, n859, n860,
         n861, n862, n863, n864, n865, n866, n867, n868, n869, n870, n871,
         n872, n873, n874, n875, n876, n877, n878, n879, n880, n881, n882,
         n883, n884, n885, n886, n887, n888, n889, n890, n891, n892, n893,
         n894, n895, n896, n897, n898, n899, n900, n901, n902, n903, n904,
         n905, n906, n907, n908, n909, n910, n911, n912, n913, n914, n915,
         n916, n917, n918, n919, n920, n921, n922, n923, n924, n925, n926,
         n927, n928, n929, n930, n931, n932, n933, n934, n935, n936, n937,
         n938, n939, n940, n941, n942, n943, n944, n945, n946, n947, n948,
         n949, n950, n951, n952, n953, n954, n955, n956, n957, n958, n959,
         n960, n961, n962, n963, n964, n965, n966, n967, n968, n969, n970,
         n971, n972, n973, n974, n975, n976, n977, n978, n979, n980, n981,
         n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, n992,
         n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003,
         n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013,
         n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023,
         n1024, n1025;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NAND2_X1 U551 ( .A1(G8), .A2(n727), .ZN(n799) );
  INV_X1 U552 ( .A(n705), .ZN(n727) );
  NOR2_X2 U553 ( .A1(n766), .A2(n680), .ZN(n705) );
  INV_X1 U554 ( .A(KEYINPUT28), .ZN(n685) );
  XNOR2_X1 U555 ( .A(n705), .B(n681), .ZN(n707) );
  INV_X1 U556 ( .A(KEYINPUT97), .ZN(n681) );
  XNOR2_X1 U557 ( .A(n704), .B(n703), .ZN(n712) );
  INV_X1 U558 ( .A(KEYINPUT29), .ZN(n703) );
  INV_X1 U559 ( .A(KEYINPUT17), .ZN(n516) );
  NAND2_X1 U560 ( .A1(n707), .A2(G2072), .ZN(n682) );
  INV_X1 U561 ( .A(KEYINPUT30), .ZN(n714) );
  INV_X1 U562 ( .A(KEYINPUT98), .ZN(n717) );
  XNOR2_X1 U563 ( .A(KEYINPUT99), .B(KEYINPUT31), .ZN(n722) );
  XNOR2_X1 U564 ( .A(n723), .B(n722), .ZN(n724) );
  INV_X1 U565 ( .A(KEYINPUT101), .ZN(n733) );
  XNOR2_X1 U566 ( .A(n734), .B(n733), .ZN(n735) );
  NOR2_X1 U567 ( .A1(G1384), .A2(G164), .ZN(n679) );
  NAND2_X1 U568 ( .A1(G160), .A2(G40), .ZN(n766) );
  NAND2_X1 U569 ( .A1(G114), .A2(n883), .ZN(n518) );
  AND2_X1 U570 ( .A1(n521), .A2(G2104), .ZN(n879) );
  NOR2_X2 U571 ( .A1(G2104), .A2(n521), .ZN(n884) );
  AND2_X2 U572 ( .A1(G2104), .A2(G2105), .ZN(n883) );
  NAND2_X1 U573 ( .A1(n880), .A2(G138), .ZN(n525) );
  AND2_X1 U574 ( .A1(n525), .A2(n524), .ZN(G164) );
  NOR2_X1 U575 ( .A1(G2104), .A2(G2105), .ZN(n517) );
  XNOR2_X2 U576 ( .A(n517), .B(n516), .ZN(n880) );
  INV_X1 U577 ( .A(G2105), .ZN(n521) );
  NAND2_X1 U578 ( .A1(n879), .A2(G102), .ZN(n520) );
  XOR2_X1 U579 ( .A(KEYINPUT91), .B(n518), .Z(n519) );
  NAND2_X1 U580 ( .A1(n520), .A2(n519), .ZN(n523) );
  AND2_X1 U581 ( .A1(G126), .A2(n884), .ZN(n522) );
  NOR2_X1 U582 ( .A1(n523), .A2(n522), .ZN(n524) );
  NAND2_X1 U583 ( .A1(G113), .A2(n883), .ZN(n526) );
  XNOR2_X1 U584 ( .A(n526), .B(KEYINPUT68), .ZN(n533) );
  NAND2_X1 U585 ( .A1(G137), .A2(n880), .ZN(n528) );
  NAND2_X1 U586 ( .A1(G125), .A2(n884), .ZN(n527) );
  NAND2_X1 U587 ( .A1(n528), .A2(n527), .ZN(n531) );
  NAND2_X1 U588 ( .A1(G101), .A2(n879), .ZN(n529) );
  XNOR2_X1 U589 ( .A(KEYINPUT23), .B(n529), .ZN(n530) );
  NOR2_X1 U590 ( .A1(n531), .A2(n530), .ZN(n532) );
  NAND2_X1 U591 ( .A1(n533), .A2(n532), .ZN(n534) );
  XNOR2_X2 U592 ( .A(KEYINPUT67), .B(n534), .ZN(G160) );
  XNOR2_X1 U593 ( .A(KEYINPUT74), .B(KEYINPUT6), .ZN(n541) );
  INV_X1 U594 ( .A(G651), .ZN(n544) );
  NOR2_X1 U595 ( .A1(G543), .A2(n544), .ZN(n535) );
  XOR2_X1 U596 ( .A(KEYINPUT1), .B(n535), .Z(n640) );
  NAND2_X1 U597 ( .A1(G63), .A2(n640), .ZN(n539) );
  XNOR2_X1 U598 ( .A(G543), .B(KEYINPUT0), .ZN(n536) );
  XNOR2_X1 U599 ( .A(n536), .B(KEYINPUT69), .ZN(n637) );
  NOR2_X1 U600 ( .A1(n637), .A2(G651), .ZN(n537) );
  XNOR2_X1 U601 ( .A(KEYINPUT66), .B(n537), .ZN(n647) );
  NAND2_X1 U602 ( .A1(G51), .A2(n647), .ZN(n538) );
  NAND2_X1 U603 ( .A1(n539), .A2(n538), .ZN(n540) );
  XNOR2_X1 U604 ( .A(n541), .B(n540), .ZN(n549) );
  NOR2_X1 U605 ( .A1(G543), .A2(G651), .ZN(n542) );
  XOR2_X1 U606 ( .A(KEYINPUT65), .B(n542), .Z(n642) );
  NAND2_X1 U607 ( .A1(n642), .A2(G89), .ZN(n543) );
  XNOR2_X1 U608 ( .A(n543), .B(KEYINPUT4), .ZN(n546) );
  NOR2_X1 U609 ( .A1(n637), .A2(n544), .ZN(n643) );
  NAND2_X1 U610 ( .A1(G76), .A2(n643), .ZN(n545) );
  NAND2_X1 U611 ( .A1(n546), .A2(n545), .ZN(n547) );
  XOR2_X1 U612 ( .A(KEYINPUT5), .B(n547), .Z(n548) );
  NOR2_X1 U613 ( .A1(n549), .A2(n548), .ZN(n551) );
  XNOR2_X1 U614 ( .A(KEYINPUT7), .B(KEYINPUT75), .ZN(n550) );
  XNOR2_X1 U615 ( .A(n551), .B(n550), .ZN(G168) );
  XOR2_X1 U616 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U617 ( .A1(G85), .A2(n642), .ZN(n553) );
  NAND2_X1 U618 ( .A1(G72), .A2(n643), .ZN(n552) );
  NAND2_X1 U619 ( .A1(n553), .A2(n552), .ZN(n557) );
  NAND2_X1 U620 ( .A1(G60), .A2(n640), .ZN(n555) );
  NAND2_X1 U621 ( .A1(G47), .A2(n647), .ZN(n554) );
  NAND2_X1 U622 ( .A1(n555), .A2(n554), .ZN(n556) );
  OR2_X1 U623 ( .A1(n557), .A2(n556), .ZN(G290) );
  AND2_X1 U624 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U625 ( .A(G132), .ZN(G219) );
  INV_X1 U626 ( .A(G82), .ZN(G220) );
  NAND2_X1 U627 ( .A1(G64), .A2(n640), .ZN(n559) );
  NAND2_X1 U628 ( .A1(G52), .A2(n647), .ZN(n558) );
  NAND2_X1 U629 ( .A1(n559), .A2(n558), .ZN(n564) );
  NAND2_X1 U630 ( .A1(G90), .A2(n642), .ZN(n561) );
  NAND2_X1 U631 ( .A1(G77), .A2(n643), .ZN(n560) );
  NAND2_X1 U632 ( .A1(n561), .A2(n560), .ZN(n562) );
  XOR2_X1 U633 ( .A(KEYINPUT9), .B(n562), .Z(n563) );
  NOR2_X1 U634 ( .A1(n564), .A2(n563), .ZN(G171) );
  NAND2_X1 U635 ( .A1(G7), .A2(G661), .ZN(n565) );
  XNOR2_X1 U636 ( .A(n565), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U637 ( .A(G223), .ZN(n822) );
  NAND2_X1 U638 ( .A1(n822), .A2(G567), .ZN(n566) );
  XOR2_X1 U639 ( .A(KEYINPUT11), .B(n566), .Z(G234) );
  NAND2_X1 U640 ( .A1(G56), .A2(n640), .ZN(n567) );
  XOR2_X1 U641 ( .A(KEYINPUT14), .B(n567), .Z(n574) );
  NAND2_X1 U642 ( .A1(G81), .A2(n642), .ZN(n568) );
  XOR2_X1 U643 ( .A(KEYINPUT71), .B(n568), .Z(n569) );
  XNOR2_X1 U644 ( .A(n569), .B(KEYINPUT12), .ZN(n571) );
  NAND2_X1 U645 ( .A1(G68), .A2(n643), .ZN(n570) );
  NAND2_X1 U646 ( .A1(n571), .A2(n570), .ZN(n572) );
  XOR2_X1 U647 ( .A(KEYINPUT13), .B(n572), .Z(n573) );
  NOR2_X1 U648 ( .A1(n574), .A2(n573), .ZN(n576) );
  NAND2_X1 U649 ( .A1(G43), .A2(n647), .ZN(n575) );
  NAND2_X1 U650 ( .A1(n576), .A2(n575), .ZN(n977) );
  INV_X1 U651 ( .A(G860), .ZN(n598) );
  OR2_X1 U652 ( .A1(n977), .A2(n598), .ZN(G153) );
  INV_X1 U653 ( .A(G171), .ZN(G301) );
  NAND2_X1 U654 ( .A1(n647), .A2(G54), .ZN(n583) );
  NAND2_X1 U655 ( .A1(G66), .A2(n640), .ZN(n578) );
  NAND2_X1 U656 ( .A1(G79), .A2(n643), .ZN(n577) );
  NAND2_X1 U657 ( .A1(n578), .A2(n577), .ZN(n581) );
  NAND2_X1 U658 ( .A1(n642), .A2(G92), .ZN(n579) );
  XOR2_X1 U659 ( .A(KEYINPUT72), .B(n579), .Z(n580) );
  NOR2_X1 U660 ( .A1(n581), .A2(n580), .ZN(n582) );
  NAND2_X1 U661 ( .A1(n583), .A2(n582), .ZN(n584) );
  XNOR2_X1 U662 ( .A(n584), .B(KEYINPUT15), .ZN(n966) );
  NOR2_X1 U663 ( .A1(n966), .A2(G868), .ZN(n585) );
  XNOR2_X1 U664 ( .A(n585), .B(KEYINPUT73), .ZN(n587) );
  NAND2_X1 U665 ( .A1(G868), .A2(G301), .ZN(n586) );
  NAND2_X1 U666 ( .A1(n587), .A2(n586), .ZN(G284) );
  NAND2_X1 U667 ( .A1(G65), .A2(n640), .ZN(n589) );
  NAND2_X1 U668 ( .A1(G53), .A2(n647), .ZN(n588) );
  NAND2_X1 U669 ( .A1(n589), .A2(n588), .ZN(n593) );
  NAND2_X1 U670 ( .A1(G91), .A2(n642), .ZN(n591) );
  NAND2_X1 U671 ( .A1(G78), .A2(n643), .ZN(n590) );
  NAND2_X1 U672 ( .A1(n591), .A2(n590), .ZN(n592) );
  NOR2_X1 U673 ( .A1(n593), .A2(n592), .ZN(n973) );
  INV_X1 U674 ( .A(n973), .ZN(G299) );
  INV_X1 U675 ( .A(G868), .ZN(n594) );
  NOR2_X1 U676 ( .A1(G286), .A2(n594), .ZN(n596) );
  NOR2_X1 U677 ( .A1(G868), .A2(G299), .ZN(n595) );
  NOR2_X1 U678 ( .A1(n596), .A2(n595), .ZN(n597) );
  XNOR2_X1 U679 ( .A(KEYINPUT76), .B(n597), .ZN(G297) );
  NAND2_X1 U680 ( .A1(n598), .A2(G559), .ZN(n599) );
  NAND2_X1 U681 ( .A1(n599), .A2(n966), .ZN(n600) );
  XNOR2_X1 U682 ( .A(n600), .B(KEYINPUT16), .ZN(G148) );
  AND2_X1 U683 ( .A1(n966), .A2(G868), .ZN(n601) );
  XNOR2_X1 U684 ( .A(n601), .B(KEYINPUT77), .ZN(n602) );
  NOR2_X1 U685 ( .A1(G559), .A2(n602), .ZN(n604) );
  NOR2_X1 U686 ( .A1(G868), .A2(n977), .ZN(n603) );
  NOR2_X1 U687 ( .A1(n604), .A2(n603), .ZN(n605) );
  XNOR2_X1 U688 ( .A(KEYINPUT78), .B(n605), .ZN(G282) );
  XOR2_X1 U689 ( .A(G2100), .B(KEYINPUT80), .Z(n615) );
  NAND2_X1 U690 ( .A1(G123), .A2(n884), .ZN(n606) );
  XNOR2_X1 U691 ( .A(n606), .B(KEYINPUT18), .ZN(n613) );
  NAND2_X1 U692 ( .A1(G111), .A2(n883), .ZN(n608) );
  NAND2_X1 U693 ( .A1(G99), .A2(n879), .ZN(n607) );
  NAND2_X1 U694 ( .A1(n608), .A2(n607), .ZN(n611) );
  NAND2_X1 U695 ( .A1(G135), .A2(n880), .ZN(n609) );
  XNOR2_X1 U696 ( .A(KEYINPUT79), .B(n609), .ZN(n610) );
  NOR2_X1 U697 ( .A1(n611), .A2(n610), .ZN(n612) );
  NAND2_X1 U698 ( .A1(n613), .A2(n612), .ZN(n997) );
  XOR2_X1 U699 ( .A(G2096), .B(n997), .Z(n614) );
  NAND2_X1 U700 ( .A1(n615), .A2(n614), .ZN(G156) );
  NAND2_X1 U701 ( .A1(G80), .A2(n643), .ZN(n616) );
  XNOR2_X1 U702 ( .A(n616), .B(KEYINPUT82), .ZN(n618) );
  NAND2_X1 U703 ( .A1(n640), .A2(G67), .ZN(n617) );
  NAND2_X1 U704 ( .A1(n618), .A2(n617), .ZN(n622) );
  NAND2_X1 U705 ( .A1(G93), .A2(n642), .ZN(n620) );
  NAND2_X1 U706 ( .A1(G55), .A2(n647), .ZN(n619) );
  NAND2_X1 U707 ( .A1(n620), .A2(n619), .ZN(n621) );
  NOR2_X1 U708 ( .A1(n622), .A2(n621), .ZN(n654) );
  NAND2_X1 U709 ( .A1(G559), .A2(n966), .ZN(n623) );
  XNOR2_X1 U710 ( .A(n623), .B(n977), .ZN(n662) );
  XOR2_X1 U711 ( .A(KEYINPUT81), .B(n662), .Z(n624) );
  NOR2_X1 U712 ( .A1(G860), .A2(n624), .ZN(n625) );
  XNOR2_X1 U713 ( .A(n654), .B(n625), .ZN(G145) );
  NAND2_X1 U714 ( .A1(G61), .A2(n640), .ZN(n627) );
  NAND2_X1 U715 ( .A1(G86), .A2(n642), .ZN(n626) );
  NAND2_X1 U716 ( .A1(n627), .A2(n626), .ZN(n630) );
  NAND2_X1 U717 ( .A1(n643), .A2(G73), .ZN(n628) );
  XOR2_X1 U718 ( .A(KEYINPUT2), .B(n628), .Z(n629) );
  NOR2_X1 U719 ( .A1(n630), .A2(n629), .ZN(n632) );
  NAND2_X1 U720 ( .A1(G48), .A2(n647), .ZN(n631) );
  NAND2_X1 U721 ( .A1(n632), .A2(n631), .ZN(G305) );
  NAND2_X1 U722 ( .A1(G651), .A2(G74), .ZN(n634) );
  NAND2_X1 U723 ( .A1(G49), .A2(n647), .ZN(n633) );
  NAND2_X1 U724 ( .A1(n634), .A2(n633), .ZN(n635) );
  NOR2_X1 U725 ( .A1(n640), .A2(n635), .ZN(n636) );
  XOR2_X1 U726 ( .A(KEYINPUT83), .B(n636), .Z(n639) );
  NAND2_X1 U727 ( .A1(n637), .A2(G87), .ZN(n638) );
  NAND2_X1 U728 ( .A1(n639), .A2(n638), .ZN(G288) );
  NAND2_X1 U729 ( .A1(G62), .A2(n640), .ZN(n641) );
  XNOR2_X1 U730 ( .A(n641), .B(KEYINPUT84), .ZN(n652) );
  NAND2_X1 U731 ( .A1(G88), .A2(n642), .ZN(n645) );
  NAND2_X1 U732 ( .A1(G75), .A2(n643), .ZN(n644) );
  NAND2_X1 U733 ( .A1(n645), .A2(n644), .ZN(n646) );
  XNOR2_X1 U734 ( .A(KEYINPUT86), .B(n646), .ZN(n650) );
  NAND2_X1 U735 ( .A1(G50), .A2(n647), .ZN(n648) );
  XNOR2_X1 U736 ( .A(KEYINPUT85), .B(n648), .ZN(n649) );
  NOR2_X1 U737 ( .A1(n650), .A2(n649), .ZN(n651) );
  NAND2_X1 U738 ( .A1(n652), .A2(n651), .ZN(G303) );
  INV_X1 U739 ( .A(G303), .ZN(G166) );
  NOR2_X1 U740 ( .A1(G868), .A2(n654), .ZN(n653) );
  XNOR2_X1 U741 ( .A(n653), .B(KEYINPUT89), .ZN(n665) );
  XOR2_X1 U742 ( .A(KEYINPUT87), .B(KEYINPUT19), .Z(n656) );
  XNOR2_X1 U743 ( .A(n654), .B(KEYINPUT88), .ZN(n655) );
  XNOR2_X1 U744 ( .A(n656), .B(n655), .ZN(n657) );
  XNOR2_X1 U745 ( .A(n657), .B(G290), .ZN(n658) );
  XNOR2_X1 U746 ( .A(n658), .B(G288), .ZN(n659) );
  XNOR2_X1 U747 ( .A(G305), .B(n659), .ZN(n661) );
  XNOR2_X1 U748 ( .A(n973), .B(G166), .ZN(n660) );
  XNOR2_X1 U749 ( .A(n661), .B(n660), .ZN(n894) );
  XNOR2_X1 U750 ( .A(n894), .B(n662), .ZN(n663) );
  NAND2_X1 U751 ( .A1(G868), .A2(n663), .ZN(n664) );
  NAND2_X1 U752 ( .A1(n665), .A2(n664), .ZN(G295) );
  NAND2_X1 U753 ( .A1(G2084), .A2(G2078), .ZN(n666) );
  XOR2_X1 U754 ( .A(KEYINPUT20), .B(n666), .Z(n667) );
  NAND2_X1 U755 ( .A1(G2090), .A2(n667), .ZN(n668) );
  XNOR2_X1 U756 ( .A(KEYINPUT21), .B(n668), .ZN(n669) );
  NAND2_X1 U757 ( .A1(n669), .A2(G2072), .ZN(G158) );
  XOR2_X1 U758 ( .A(KEYINPUT70), .B(G57), .Z(G237) );
  XNOR2_X1 U759 ( .A(KEYINPUT90), .B(G44), .ZN(n670) );
  XNOR2_X1 U760 ( .A(n670), .B(KEYINPUT3), .ZN(G218) );
  NAND2_X1 U761 ( .A1(G108), .A2(G120), .ZN(n671) );
  NOR2_X1 U762 ( .A1(G237), .A2(n671), .ZN(n672) );
  NAND2_X1 U763 ( .A1(G69), .A2(n672), .ZN(n826) );
  NAND2_X1 U764 ( .A1(n826), .A2(G567), .ZN(n677) );
  NOR2_X1 U765 ( .A1(G220), .A2(G219), .ZN(n673) );
  XOR2_X1 U766 ( .A(KEYINPUT22), .B(n673), .Z(n674) );
  NOR2_X1 U767 ( .A1(G218), .A2(n674), .ZN(n675) );
  NAND2_X1 U768 ( .A1(G96), .A2(n675), .ZN(n827) );
  NAND2_X1 U769 ( .A1(n827), .A2(G2106), .ZN(n676) );
  NAND2_X1 U770 ( .A1(n677), .A2(n676), .ZN(n828) );
  NAND2_X1 U771 ( .A1(G661), .A2(G483), .ZN(n678) );
  NOR2_X1 U772 ( .A1(n828), .A2(n678), .ZN(n825) );
  NAND2_X1 U773 ( .A1(n825), .A2(G36), .ZN(G176) );
  XNOR2_X1 U774 ( .A(n679), .B(KEYINPUT64), .ZN(n765) );
  INV_X1 U775 ( .A(n765), .ZN(n680) );
  XNOR2_X1 U776 ( .A(n682), .B(KEYINPUT27), .ZN(n684) );
  INV_X1 U777 ( .A(G1956), .ZN(n939) );
  NOR2_X1 U778 ( .A1(n939), .A2(n707), .ZN(n683) );
  NOR2_X1 U779 ( .A1(n684), .A2(n683), .ZN(n687) );
  NOR2_X1 U780 ( .A1(n973), .A2(n687), .ZN(n686) );
  XNOR2_X1 U781 ( .A(n686), .B(n685), .ZN(n702) );
  NAND2_X1 U782 ( .A1(n973), .A2(n687), .ZN(n700) );
  AND2_X1 U783 ( .A1(n705), .A2(G1996), .ZN(n688) );
  XOR2_X1 U784 ( .A(n688), .B(KEYINPUT26), .Z(n690) );
  NAND2_X1 U785 ( .A1(n727), .A2(G1341), .ZN(n689) );
  NAND2_X1 U786 ( .A1(n690), .A2(n689), .ZN(n691) );
  NOR2_X1 U787 ( .A1(n977), .A2(n691), .ZN(n692) );
  OR2_X1 U788 ( .A1(n966), .A2(n692), .ZN(n698) );
  NAND2_X1 U789 ( .A1(n966), .A2(n692), .ZN(n696) );
  NAND2_X1 U790 ( .A1(G2067), .A2(n707), .ZN(n694) );
  NAND2_X1 U791 ( .A1(G1348), .A2(n727), .ZN(n693) );
  NAND2_X1 U792 ( .A1(n694), .A2(n693), .ZN(n695) );
  NAND2_X1 U793 ( .A1(n696), .A2(n695), .ZN(n697) );
  NAND2_X1 U794 ( .A1(n698), .A2(n697), .ZN(n699) );
  NAND2_X1 U795 ( .A1(n700), .A2(n699), .ZN(n701) );
  NAND2_X1 U796 ( .A1(n702), .A2(n701), .ZN(n704) );
  XOR2_X1 U797 ( .A(KEYINPUT95), .B(G1961), .Z(n948) );
  NOR2_X1 U798 ( .A1(n705), .A2(n948), .ZN(n706) );
  XNOR2_X1 U799 ( .A(n706), .B(KEYINPUT96), .ZN(n710) );
  INV_X1 U800 ( .A(n707), .ZN(n708) );
  XOR2_X1 U801 ( .A(KEYINPUT25), .B(G2078), .Z(n917) );
  NOR2_X1 U802 ( .A1(n708), .A2(n917), .ZN(n709) );
  NOR2_X1 U803 ( .A1(n710), .A2(n709), .ZN(n719) );
  OR2_X1 U804 ( .A1(n719), .A2(G301), .ZN(n711) );
  NAND2_X1 U805 ( .A1(n712), .A2(n711), .ZN(n726) );
  NOR2_X1 U806 ( .A1(G2084), .A2(n727), .ZN(n741) );
  NOR2_X1 U807 ( .A1(G1966), .A2(n799), .ZN(n739) );
  NOR2_X1 U808 ( .A1(n741), .A2(n739), .ZN(n713) );
  AND2_X1 U809 ( .A1(n713), .A2(G8), .ZN(n715) );
  XNOR2_X1 U810 ( .A(n715), .B(n714), .ZN(n716) );
  NOR2_X1 U811 ( .A1(G168), .A2(n716), .ZN(n718) );
  XNOR2_X1 U812 ( .A(n718), .B(n717), .ZN(n721) );
  NAND2_X1 U813 ( .A1(G301), .A2(n719), .ZN(n720) );
  NAND2_X1 U814 ( .A1(n721), .A2(n720), .ZN(n723) );
  INV_X1 U815 ( .A(n724), .ZN(n725) );
  NAND2_X1 U816 ( .A1(n726), .A2(n725), .ZN(n737) );
  NAND2_X1 U817 ( .A1(n737), .A2(G286), .ZN(n732) );
  NOR2_X1 U818 ( .A1(G1971), .A2(n799), .ZN(n729) );
  NOR2_X1 U819 ( .A1(G2090), .A2(n727), .ZN(n728) );
  NOR2_X1 U820 ( .A1(n729), .A2(n728), .ZN(n730) );
  NAND2_X1 U821 ( .A1(n730), .A2(G303), .ZN(n731) );
  NAND2_X1 U822 ( .A1(n732), .A2(n731), .ZN(n734) );
  NAND2_X1 U823 ( .A1(n735), .A2(G8), .ZN(n736) );
  XNOR2_X1 U824 ( .A(n736), .B(KEYINPUT32), .ZN(n788) );
  INV_X1 U825 ( .A(n737), .ZN(n738) );
  NOR2_X1 U826 ( .A1(n739), .A2(n738), .ZN(n740) );
  XNOR2_X1 U827 ( .A(n740), .B(KEYINPUT100), .ZN(n743) );
  NAND2_X1 U828 ( .A1(n741), .A2(G8), .ZN(n742) );
  NAND2_X1 U829 ( .A1(n743), .A2(n742), .ZN(n786) );
  NAND2_X1 U830 ( .A1(n788), .A2(n786), .ZN(n746) );
  NOR2_X1 U831 ( .A1(G2090), .A2(G303), .ZN(n744) );
  NAND2_X1 U832 ( .A1(G8), .A2(n744), .ZN(n745) );
  NAND2_X1 U833 ( .A1(n746), .A2(n745), .ZN(n747) );
  XNOR2_X1 U834 ( .A(n747), .B(KEYINPUT102), .ZN(n779) );
  NAND2_X1 U835 ( .A1(G117), .A2(n883), .ZN(n749) );
  NAND2_X1 U836 ( .A1(G129), .A2(n884), .ZN(n748) );
  NAND2_X1 U837 ( .A1(n749), .A2(n748), .ZN(n752) );
  NAND2_X1 U838 ( .A1(n879), .A2(G105), .ZN(n750) );
  XOR2_X1 U839 ( .A(KEYINPUT38), .B(n750), .Z(n751) );
  NOR2_X1 U840 ( .A1(n752), .A2(n751), .ZN(n754) );
  NAND2_X1 U841 ( .A1(n880), .A2(G141), .ZN(n753) );
  NAND2_X1 U842 ( .A1(n754), .A2(n753), .ZN(n863) );
  NAND2_X1 U843 ( .A1(G1996), .A2(n863), .ZN(n755) );
  XNOR2_X1 U844 ( .A(n755), .B(KEYINPUT93), .ZN(n764) );
  NAND2_X1 U845 ( .A1(n883), .A2(G107), .ZN(n756) );
  XNOR2_X1 U846 ( .A(n756), .B(KEYINPUT92), .ZN(n758) );
  NAND2_X1 U847 ( .A1(G119), .A2(n884), .ZN(n757) );
  NAND2_X1 U848 ( .A1(n758), .A2(n757), .ZN(n762) );
  NAND2_X1 U849 ( .A1(G95), .A2(n879), .ZN(n760) );
  NAND2_X1 U850 ( .A1(G131), .A2(n880), .ZN(n759) );
  NAND2_X1 U851 ( .A1(n760), .A2(n759), .ZN(n761) );
  OR2_X1 U852 ( .A1(n762), .A2(n761), .ZN(n862) );
  AND2_X1 U853 ( .A1(G1991), .A2(n862), .ZN(n763) );
  NOR2_X1 U854 ( .A1(n764), .A2(n763), .ZN(n808) );
  XOR2_X1 U855 ( .A(G1986), .B(G290), .Z(n976) );
  NAND2_X1 U856 ( .A1(n808), .A2(n976), .ZN(n767) );
  NOR2_X1 U857 ( .A1(n766), .A2(n765), .ZN(n818) );
  NAND2_X1 U858 ( .A1(n767), .A2(n818), .ZN(n777) );
  NAND2_X1 U859 ( .A1(G104), .A2(n879), .ZN(n769) );
  NAND2_X1 U860 ( .A1(G140), .A2(n880), .ZN(n768) );
  NAND2_X1 U861 ( .A1(n769), .A2(n768), .ZN(n770) );
  XNOR2_X1 U862 ( .A(KEYINPUT34), .B(n770), .ZN(n775) );
  NAND2_X1 U863 ( .A1(G116), .A2(n883), .ZN(n772) );
  NAND2_X1 U864 ( .A1(G128), .A2(n884), .ZN(n771) );
  NAND2_X1 U865 ( .A1(n772), .A2(n771), .ZN(n773) );
  XOR2_X1 U866 ( .A(KEYINPUT35), .B(n773), .Z(n774) );
  NOR2_X1 U867 ( .A1(n775), .A2(n774), .ZN(n776) );
  XNOR2_X1 U868 ( .A(KEYINPUT36), .B(n776), .ZN(n890) );
  XNOR2_X1 U869 ( .A(G2067), .B(KEYINPUT37), .ZN(n815) );
  NOR2_X1 U870 ( .A1(n890), .A2(n815), .ZN(n1016) );
  NAND2_X1 U871 ( .A1(n818), .A2(n1016), .ZN(n813) );
  AND2_X1 U872 ( .A1(n777), .A2(n813), .ZN(n795) );
  AND2_X1 U873 ( .A1(n799), .A2(n795), .ZN(n778) );
  AND2_X1 U874 ( .A1(n779), .A2(n778), .ZN(n785) );
  NOR2_X1 U875 ( .A1(G1981), .A2(G305), .ZN(n780) );
  XOR2_X1 U876 ( .A(n780), .B(KEYINPUT24), .Z(n781) );
  XNOR2_X1 U877 ( .A(KEYINPUT94), .B(n781), .ZN(n782) );
  NOR2_X1 U878 ( .A1(n799), .A2(n782), .ZN(n783) );
  AND2_X1 U879 ( .A1(n795), .A2(n783), .ZN(n784) );
  NOR2_X1 U880 ( .A1(n785), .A2(n784), .ZN(n806) );
  NAND2_X1 U881 ( .A1(G1976), .A2(G288), .ZN(n967) );
  AND2_X1 U882 ( .A1(n786), .A2(n967), .ZN(n787) );
  AND2_X1 U883 ( .A1(n788), .A2(n787), .ZN(n792) );
  INV_X1 U884 ( .A(n967), .ZN(n790) );
  NOR2_X1 U885 ( .A1(G1976), .A2(G288), .ZN(n793) );
  NOR2_X1 U886 ( .A1(G1971), .A2(G303), .ZN(n789) );
  NOR2_X1 U887 ( .A1(n793), .A2(n789), .ZN(n991) );
  NOR2_X1 U888 ( .A1(n790), .A2(n991), .ZN(n791) );
  NOR2_X1 U889 ( .A1(n792), .A2(n791), .ZN(n801) );
  NAND2_X1 U890 ( .A1(n793), .A2(KEYINPUT33), .ZN(n794) );
  OR2_X1 U891 ( .A1(n794), .A2(n799), .ZN(n797) );
  XOR2_X1 U892 ( .A(G1981), .B(G305), .Z(n969) );
  AND2_X1 U893 ( .A1(n969), .A2(n795), .ZN(n796) );
  AND2_X1 U894 ( .A1(n797), .A2(n796), .ZN(n802) );
  INV_X1 U895 ( .A(n802), .ZN(n798) );
  OR2_X1 U896 ( .A1(n799), .A2(n798), .ZN(n800) );
  NOR2_X1 U897 ( .A1(n801), .A2(n800), .ZN(n804) );
  AND2_X1 U898 ( .A1(n802), .A2(KEYINPUT33), .ZN(n803) );
  NOR2_X1 U899 ( .A1(n804), .A2(n803), .ZN(n805) );
  NAND2_X1 U900 ( .A1(n806), .A2(n805), .ZN(n807) );
  XNOR2_X1 U901 ( .A(n807), .B(KEYINPUT103), .ZN(n820) );
  NOR2_X1 U902 ( .A1(G1996), .A2(n863), .ZN(n1007) );
  INV_X1 U903 ( .A(n808), .ZN(n1000) );
  NOR2_X1 U904 ( .A1(G1991), .A2(n862), .ZN(n996) );
  NOR2_X1 U905 ( .A1(G1986), .A2(G290), .ZN(n809) );
  NOR2_X1 U906 ( .A1(n996), .A2(n809), .ZN(n810) );
  NOR2_X1 U907 ( .A1(n1000), .A2(n810), .ZN(n811) );
  NOR2_X1 U908 ( .A1(n1007), .A2(n811), .ZN(n812) );
  XNOR2_X1 U909 ( .A(n812), .B(KEYINPUT39), .ZN(n814) );
  NAND2_X1 U910 ( .A1(n814), .A2(n813), .ZN(n816) );
  NAND2_X1 U911 ( .A1(n890), .A2(n815), .ZN(n1009) );
  NAND2_X1 U912 ( .A1(n816), .A2(n1009), .ZN(n817) );
  NAND2_X1 U913 ( .A1(n818), .A2(n817), .ZN(n819) );
  NAND2_X1 U914 ( .A1(n820), .A2(n819), .ZN(n821) );
  XNOR2_X1 U915 ( .A(n821), .B(KEYINPUT40), .ZN(G329) );
  NAND2_X1 U916 ( .A1(G2106), .A2(n822), .ZN(G217) );
  AND2_X1 U917 ( .A1(G15), .A2(G2), .ZN(n823) );
  NAND2_X1 U918 ( .A1(G661), .A2(n823), .ZN(G259) );
  NAND2_X1 U919 ( .A1(G3), .A2(G1), .ZN(n824) );
  NAND2_X1 U920 ( .A1(n825), .A2(n824), .ZN(G188) );
  NOR2_X1 U921 ( .A1(n827), .A2(n826), .ZN(G325) );
  XOR2_X1 U922 ( .A(KEYINPUT104), .B(G325), .Z(G261) );
  INV_X1 U924 ( .A(G120), .ZN(G236) );
  INV_X1 U925 ( .A(G108), .ZN(G238) );
  INV_X1 U926 ( .A(G96), .ZN(G221) );
  INV_X1 U927 ( .A(G69), .ZN(G235) );
  INV_X1 U928 ( .A(n828), .ZN(G319) );
  XOR2_X1 U929 ( .A(KEYINPUT42), .B(G2090), .Z(n830) );
  XNOR2_X1 U930 ( .A(G2084), .B(G2072), .ZN(n829) );
  XNOR2_X1 U931 ( .A(n830), .B(n829), .ZN(n831) );
  XOR2_X1 U932 ( .A(n831), .B(G2096), .Z(n833) );
  XNOR2_X1 U933 ( .A(G2067), .B(G2078), .ZN(n832) );
  XNOR2_X1 U934 ( .A(n833), .B(n832), .ZN(n837) );
  XOR2_X1 U935 ( .A(G2100), .B(KEYINPUT43), .Z(n835) );
  XNOR2_X1 U936 ( .A(G2678), .B(KEYINPUT105), .ZN(n834) );
  XNOR2_X1 U937 ( .A(n835), .B(n834), .ZN(n836) );
  XOR2_X1 U938 ( .A(n837), .B(n836), .Z(G227) );
  XOR2_X1 U939 ( .A(G1971), .B(G1986), .Z(n839) );
  XNOR2_X1 U940 ( .A(G1996), .B(G1991), .ZN(n838) );
  XNOR2_X1 U941 ( .A(n839), .B(n838), .ZN(n849) );
  XOR2_X1 U942 ( .A(KEYINPUT107), .B(KEYINPUT108), .Z(n841) );
  XNOR2_X1 U943 ( .A(G1956), .B(KEYINPUT41), .ZN(n840) );
  XNOR2_X1 U944 ( .A(n841), .B(n840), .ZN(n845) );
  XOR2_X1 U945 ( .A(G1976), .B(G1981), .Z(n843) );
  XNOR2_X1 U946 ( .A(G1966), .B(G1961), .ZN(n842) );
  XNOR2_X1 U947 ( .A(n843), .B(n842), .ZN(n844) );
  XOR2_X1 U948 ( .A(n845), .B(n844), .Z(n847) );
  XNOR2_X1 U949 ( .A(KEYINPUT106), .B(G2474), .ZN(n846) );
  XNOR2_X1 U950 ( .A(n847), .B(n846), .ZN(n848) );
  XNOR2_X1 U951 ( .A(n849), .B(n848), .ZN(G229) );
  NAND2_X1 U952 ( .A1(G124), .A2(n884), .ZN(n850) );
  XNOR2_X1 U953 ( .A(n850), .B(KEYINPUT44), .ZN(n853) );
  NAND2_X1 U954 ( .A1(G100), .A2(n879), .ZN(n851) );
  XOR2_X1 U955 ( .A(KEYINPUT109), .B(n851), .Z(n852) );
  NAND2_X1 U956 ( .A1(n853), .A2(n852), .ZN(n857) );
  NAND2_X1 U957 ( .A1(G112), .A2(n883), .ZN(n855) );
  NAND2_X1 U958 ( .A1(G136), .A2(n880), .ZN(n854) );
  NAND2_X1 U959 ( .A1(n855), .A2(n854), .ZN(n856) );
  NOR2_X1 U960 ( .A1(n857), .A2(n856), .ZN(G162) );
  XOR2_X1 U961 ( .A(G164), .B(G160), .Z(n858) );
  XNOR2_X1 U962 ( .A(n997), .B(n858), .ZN(n878) );
  XOR2_X1 U963 ( .A(KEYINPUT48), .B(KEYINPUT46), .Z(n860) );
  XNOR2_X1 U964 ( .A(KEYINPUT113), .B(KEYINPUT112), .ZN(n859) );
  XNOR2_X1 U965 ( .A(n860), .B(n859), .ZN(n861) );
  XNOR2_X1 U966 ( .A(G162), .B(n861), .ZN(n865) );
  XOR2_X1 U967 ( .A(n863), .B(n862), .Z(n864) );
  XNOR2_X1 U968 ( .A(n865), .B(n864), .ZN(n876) );
  NAND2_X1 U969 ( .A1(G118), .A2(n883), .ZN(n867) );
  NAND2_X1 U970 ( .A1(G130), .A2(n884), .ZN(n866) );
  NAND2_X1 U971 ( .A1(n867), .A2(n866), .ZN(n874) );
  NAND2_X1 U972 ( .A1(n879), .A2(G106), .ZN(n868) );
  XNOR2_X1 U973 ( .A(KEYINPUT110), .B(n868), .ZN(n871) );
  NAND2_X1 U974 ( .A1(n880), .A2(G142), .ZN(n869) );
  XOR2_X1 U975 ( .A(KEYINPUT111), .B(n869), .Z(n870) );
  NAND2_X1 U976 ( .A1(n871), .A2(n870), .ZN(n872) );
  XOR2_X1 U977 ( .A(n872), .B(KEYINPUT45), .Z(n873) );
  NOR2_X1 U978 ( .A1(n874), .A2(n873), .ZN(n875) );
  XOR2_X1 U979 ( .A(n876), .B(n875), .Z(n877) );
  XNOR2_X1 U980 ( .A(n878), .B(n877), .ZN(n892) );
  NAND2_X1 U981 ( .A1(G103), .A2(n879), .ZN(n882) );
  NAND2_X1 U982 ( .A1(G139), .A2(n880), .ZN(n881) );
  NAND2_X1 U983 ( .A1(n882), .A2(n881), .ZN(n889) );
  NAND2_X1 U984 ( .A1(G115), .A2(n883), .ZN(n886) );
  NAND2_X1 U985 ( .A1(G127), .A2(n884), .ZN(n885) );
  NAND2_X1 U986 ( .A1(n886), .A2(n885), .ZN(n887) );
  XOR2_X1 U987 ( .A(KEYINPUT47), .B(n887), .Z(n888) );
  NOR2_X1 U988 ( .A1(n889), .A2(n888), .ZN(n1001) );
  XNOR2_X1 U989 ( .A(n890), .B(n1001), .ZN(n891) );
  XNOR2_X1 U990 ( .A(n892), .B(n891), .ZN(n893) );
  NOR2_X1 U991 ( .A1(G37), .A2(n893), .ZN(G395) );
  XNOR2_X1 U992 ( .A(n977), .B(n894), .ZN(n896) );
  XNOR2_X1 U993 ( .A(G171), .B(n966), .ZN(n895) );
  XNOR2_X1 U994 ( .A(n896), .B(n895), .ZN(n897) );
  XOR2_X1 U995 ( .A(G286), .B(n897), .Z(n898) );
  NOR2_X1 U996 ( .A1(G37), .A2(n898), .ZN(G397) );
  XOR2_X1 U997 ( .A(G2451), .B(G2430), .Z(n900) );
  XNOR2_X1 U998 ( .A(G2438), .B(G2443), .ZN(n899) );
  XNOR2_X1 U999 ( .A(n900), .B(n899), .ZN(n906) );
  XOR2_X1 U1000 ( .A(G2435), .B(G2454), .Z(n902) );
  XNOR2_X1 U1001 ( .A(G1341), .B(G1348), .ZN(n901) );
  XNOR2_X1 U1002 ( .A(n902), .B(n901), .ZN(n904) );
  XOR2_X1 U1003 ( .A(G2446), .B(G2427), .Z(n903) );
  XNOR2_X1 U1004 ( .A(n904), .B(n903), .ZN(n905) );
  XOR2_X1 U1005 ( .A(n906), .B(n905), .Z(n907) );
  NAND2_X1 U1006 ( .A1(G14), .A2(n907), .ZN(n913) );
  NAND2_X1 U1007 ( .A1(G319), .A2(n913), .ZN(n910) );
  NOR2_X1 U1008 ( .A1(G227), .A2(G229), .ZN(n908) );
  XNOR2_X1 U1009 ( .A(KEYINPUT49), .B(n908), .ZN(n909) );
  NOR2_X1 U1010 ( .A1(n910), .A2(n909), .ZN(n912) );
  NOR2_X1 U1011 ( .A1(G395), .A2(G397), .ZN(n911) );
  NAND2_X1 U1012 ( .A1(n912), .A2(n911), .ZN(G225) );
  INV_X1 U1013 ( .A(G225), .ZN(G308) );
  INV_X1 U1014 ( .A(n913), .ZN(G401) );
  XNOR2_X1 U1015 ( .A(G32), .B(G1996), .ZN(n914) );
  XNOR2_X1 U1016 ( .A(n914), .B(KEYINPUT117), .ZN(n926) );
  XOR2_X1 U1017 ( .A(G1991), .B(G25), .Z(n915) );
  NAND2_X1 U1018 ( .A1(n915), .A2(G28), .ZN(n916) );
  XNOR2_X1 U1019 ( .A(n916), .B(KEYINPUT115), .ZN(n921) );
  XNOR2_X1 U1020 ( .A(G2067), .B(G26), .ZN(n919) );
  XNOR2_X1 U1021 ( .A(G27), .B(n917), .ZN(n918) );
  NOR2_X1 U1022 ( .A1(n919), .A2(n918), .ZN(n920) );
  NAND2_X1 U1023 ( .A1(n921), .A2(n920), .ZN(n924) );
  XNOR2_X1 U1024 ( .A(KEYINPUT116), .B(G2072), .ZN(n922) );
  XNOR2_X1 U1025 ( .A(G33), .B(n922), .ZN(n923) );
  NOR2_X1 U1026 ( .A1(n924), .A2(n923), .ZN(n925) );
  NAND2_X1 U1027 ( .A1(n926), .A2(n925), .ZN(n927) );
  XNOR2_X1 U1028 ( .A(KEYINPUT53), .B(n927), .ZN(n931) );
  XOR2_X1 U1029 ( .A(G34), .B(KEYINPUT118), .Z(n929) );
  XNOR2_X1 U1030 ( .A(G2084), .B(KEYINPUT54), .ZN(n928) );
  XNOR2_X1 U1031 ( .A(n929), .B(n928), .ZN(n930) );
  NAND2_X1 U1032 ( .A1(n931), .A2(n930), .ZN(n933) );
  XNOR2_X1 U1033 ( .A(G35), .B(G2090), .ZN(n932) );
  NOR2_X1 U1034 ( .A1(n933), .A2(n932), .ZN(n934) );
  XNOR2_X1 U1035 ( .A(n934), .B(KEYINPUT55), .ZN(n936) );
  INV_X1 U1036 ( .A(G29), .ZN(n935) );
  NAND2_X1 U1037 ( .A1(n936), .A2(n935), .ZN(n937) );
  NAND2_X1 U1038 ( .A1(n937), .A2(G11), .ZN(n938) );
  XNOR2_X1 U1039 ( .A(n938), .B(KEYINPUT119), .ZN(n965) );
  XNOR2_X1 U1040 ( .A(G20), .B(n939), .ZN(n943) );
  XNOR2_X1 U1041 ( .A(G1341), .B(G19), .ZN(n941) );
  XNOR2_X1 U1042 ( .A(G6), .B(G1981), .ZN(n940) );
  NOR2_X1 U1043 ( .A1(n941), .A2(n940), .ZN(n942) );
  NAND2_X1 U1044 ( .A1(n943), .A2(n942), .ZN(n946) );
  XOR2_X1 U1045 ( .A(KEYINPUT59), .B(G1348), .Z(n944) );
  XNOR2_X1 U1046 ( .A(G4), .B(n944), .ZN(n945) );
  NOR2_X1 U1047 ( .A1(n946), .A2(n945), .ZN(n947) );
  XNOR2_X1 U1048 ( .A(KEYINPUT60), .B(n947), .ZN(n952) );
  XNOR2_X1 U1049 ( .A(G1966), .B(G21), .ZN(n950) );
  XNOR2_X1 U1050 ( .A(n948), .B(G5), .ZN(n949) );
  NOR2_X1 U1051 ( .A1(n950), .A2(n949), .ZN(n951) );
  NAND2_X1 U1052 ( .A1(n952), .A2(n951), .ZN(n960) );
  XNOR2_X1 U1053 ( .A(G1986), .B(G24), .ZN(n954) );
  XNOR2_X1 U1054 ( .A(G23), .B(G1976), .ZN(n953) );
  NOR2_X1 U1055 ( .A1(n954), .A2(n953), .ZN(n957) );
  XNOR2_X1 U1056 ( .A(G1971), .B(KEYINPUT125), .ZN(n955) );
  XNOR2_X1 U1057 ( .A(n955), .B(G22), .ZN(n956) );
  NAND2_X1 U1058 ( .A1(n957), .A2(n956), .ZN(n958) );
  XNOR2_X1 U1059 ( .A(KEYINPUT58), .B(n958), .ZN(n959) );
  NOR2_X1 U1060 ( .A1(n960), .A2(n959), .ZN(n961) );
  XOR2_X1 U1061 ( .A(KEYINPUT61), .B(n961), .Z(n962) );
  NOR2_X1 U1062 ( .A1(G16), .A2(n962), .ZN(n963) );
  XOR2_X1 U1063 ( .A(KEYINPUT126), .B(n963), .Z(n964) );
  NAND2_X1 U1064 ( .A1(n965), .A2(n964), .ZN(n1024) );
  XNOR2_X1 U1065 ( .A(KEYINPUT56), .B(G16), .ZN(n994) );
  XNOR2_X1 U1066 ( .A(n966), .B(G1348), .ZN(n968) );
  NAND2_X1 U1067 ( .A1(n968), .A2(n967), .ZN(n989) );
  XNOR2_X1 U1068 ( .A(G1966), .B(G168), .ZN(n970) );
  NAND2_X1 U1069 ( .A1(n970), .A2(n969), .ZN(n971) );
  XNOR2_X1 U1070 ( .A(n971), .B(KEYINPUT120), .ZN(n972) );
  XNOR2_X1 U1071 ( .A(KEYINPUT57), .B(n972), .ZN(n987) );
  XNOR2_X1 U1072 ( .A(n973), .B(G1956), .ZN(n974) );
  XNOR2_X1 U1073 ( .A(n974), .B(KEYINPUT122), .ZN(n975) );
  NAND2_X1 U1074 ( .A1(n976), .A2(n975), .ZN(n980) );
  XOR2_X1 U1075 ( .A(G1341), .B(n977), .Z(n978) );
  XNOR2_X1 U1076 ( .A(KEYINPUT123), .B(n978), .ZN(n979) );
  NOR2_X1 U1077 ( .A1(n980), .A2(n979), .ZN(n982) );
  NAND2_X1 U1078 ( .A1(G1971), .A2(G303), .ZN(n981) );
  NAND2_X1 U1079 ( .A1(n982), .A2(n981), .ZN(n985) );
  XOR2_X1 U1080 ( .A(G1961), .B(G301), .Z(n983) );
  XNOR2_X1 U1081 ( .A(KEYINPUT121), .B(n983), .ZN(n984) );
  NOR2_X1 U1082 ( .A1(n985), .A2(n984), .ZN(n986) );
  NAND2_X1 U1083 ( .A1(n987), .A2(n986), .ZN(n988) );
  NOR2_X1 U1084 ( .A1(n989), .A2(n988), .ZN(n990) );
  NAND2_X1 U1085 ( .A1(n991), .A2(n990), .ZN(n992) );
  XNOR2_X1 U1086 ( .A(KEYINPUT124), .B(n992), .ZN(n993) );
  NAND2_X1 U1087 ( .A1(n994), .A2(n993), .ZN(n1022) );
  XOR2_X1 U1088 ( .A(G160), .B(G2084), .Z(n995) );
  NOR2_X1 U1089 ( .A1(n996), .A2(n995), .ZN(n998) );
  NAND2_X1 U1090 ( .A1(n998), .A2(n997), .ZN(n999) );
  NOR2_X1 U1091 ( .A1(n1000), .A2(n999), .ZN(n1014) );
  XNOR2_X1 U1092 ( .A(G2072), .B(n1001), .ZN(n1004) );
  XNOR2_X1 U1093 ( .A(G164), .B(G2078), .ZN(n1002) );
  XNOR2_X1 U1094 ( .A(n1002), .B(KEYINPUT114), .ZN(n1003) );
  NAND2_X1 U1095 ( .A1(n1004), .A2(n1003), .ZN(n1005) );
  XNOR2_X1 U1096 ( .A(n1005), .B(KEYINPUT50), .ZN(n1012) );
  XOR2_X1 U1097 ( .A(G2090), .B(G162), .Z(n1006) );
  NOR2_X1 U1098 ( .A1(n1007), .A2(n1006), .ZN(n1008) );
  XOR2_X1 U1099 ( .A(KEYINPUT51), .B(n1008), .Z(n1010) );
  NAND2_X1 U1100 ( .A1(n1010), .A2(n1009), .ZN(n1011) );
  NOR2_X1 U1101 ( .A1(n1012), .A2(n1011), .ZN(n1013) );
  NAND2_X1 U1102 ( .A1(n1014), .A2(n1013), .ZN(n1015) );
  NOR2_X1 U1103 ( .A1(n1016), .A2(n1015), .ZN(n1017) );
  XNOR2_X1 U1104 ( .A(KEYINPUT52), .B(n1017), .ZN(n1019) );
  INV_X1 U1105 ( .A(KEYINPUT55), .ZN(n1018) );
  NAND2_X1 U1106 ( .A1(n1019), .A2(n1018), .ZN(n1020) );
  NAND2_X1 U1107 ( .A1(n1020), .A2(G29), .ZN(n1021) );
  NAND2_X1 U1108 ( .A1(n1022), .A2(n1021), .ZN(n1023) );
  NOR2_X1 U1109 ( .A1(n1024), .A2(n1023), .ZN(n1025) );
  XNOR2_X1 U1110 ( .A(n1025), .B(KEYINPUT62), .ZN(G311) );
  INV_X1 U1111 ( .A(G311), .ZN(G150) );
endmodule

