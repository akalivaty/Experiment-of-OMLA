//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 0 1 0 0 0 1 1 1 0 0 1 1 0 1 0 0 1 1 0 0 0 0 1 0 0 1 0 1 1 1 0 1 0 0 0 1 1 0 1 1 0 0 1 0 0 1 1 0 0 0 1 1 0 0 1 0 0 1 0 0 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:24:06 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n590, new_n591, new_n592, new_n593, new_n594,
    new_n595, new_n596, new_n597, new_n598, new_n599, new_n600, new_n602,
    new_n603, new_n604, new_n605, new_n606, new_n607, new_n608, new_n609,
    new_n611, new_n612, new_n613, new_n614, new_n615, new_n616, new_n617,
    new_n618, new_n619, new_n620, new_n621, new_n622, new_n623, new_n624,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n643, new_n644, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n654, new_n655, new_n657,
    new_n658, new_n659, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n672, new_n673,
    new_n674, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n686, new_n687, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n863,
    new_n864, new_n865, new_n866, new_n867, new_n868, new_n869, new_n870,
    new_n871, new_n872, new_n873, new_n875, new_n876, new_n877, new_n878,
    new_n879, new_n880, new_n881, new_n882, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n933, new_n934, new_n935, new_n936, new_n937, new_n938,
    new_n939, new_n940, new_n941, new_n942, new_n943, new_n944, new_n945,
    new_n946;
  XNOR2_X1  g000(.A(KEYINPUT22), .B(G137), .ZN(new_n187));
  INV_X1    g001(.A(G953), .ZN(new_n188));
  NAND3_X1  g002(.A1(new_n188), .A2(G221), .A3(G234), .ZN(new_n189));
  XNOR2_X1  g003(.A(new_n187), .B(new_n189), .ZN(new_n190));
  INV_X1    g004(.A(new_n190), .ZN(new_n191));
  INV_X1    g005(.A(G125), .ZN(new_n192));
  NOR3_X1   g006(.A1(new_n192), .A2(KEYINPUT16), .A3(G140), .ZN(new_n193));
  XNOR2_X1  g007(.A(G125), .B(G140), .ZN(new_n194));
  AOI21_X1  g008(.A(new_n193), .B1(new_n194), .B2(KEYINPUT16), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n195), .A2(G146), .ZN(new_n196));
  INV_X1    g010(.A(KEYINPUT78), .ZN(new_n197));
  XNOR2_X1  g011(.A(new_n196), .B(new_n197), .ZN(new_n198));
  INV_X1    g012(.A(KEYINPUT77), .ZN(new_n199));
  INV_X1    g013(.A(G128), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n200), .A2(G119), .ZN(new_n201));
  INV_X1    g015(.A(new_n201), .ZN(new_n202));
  INV_X1    g016(.A(G119), .ZN(new_n203));
  AOI21_X1  g017(.A(KEYINPUT75), .B1(new_n203), .B2(G128), .ZN(new_n204));
  NOR2_X1   g018(.A1(new_n202), .A2(new_n204), .ZN(new_n205));
  NOR2_X1   g019(.A1(new_n201), .A2(KEYINPUT75), .ZN(new_n206));
  NOR2_X1   g020(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  XOR2_X1   g021(.A(KEYINPUT24), .B(G110), .Z(new_n208));
  OAI21_X1  g022(.A(new_n199), .B1(new_n207), .B2(new_n208), .ZN(new_n209));
  NOR2_X1   g023(.A1(new_n202), .A2(KEYINPUT23), .ZN(new_n210));
  NOR2_X1   g024(.A1(new_n200), .A2(G119), .ZN(new_n211));
  INV_X1    g025(.A(KEYINPUT23), .ZN(new_n212));
  NOR2_X1   g026(.A1(new_n201), .A2(new_n212), .ZN(new_n213));
  NOR3_X1   g027(.A1(new_n210), .A2(new_n211), .A3(new_n213), .ZN(new_n214));
  INV_X1    g028(.A(G110), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n214), .A2(new_n215), .ZN(new_n216));
  INV_X1    g030(.A(new_n208), .ZN(new_n217));
  OAI211_X1 g031(.A(new_n217), .B(KEYINPUT77), .C1(new_n205), .C2(new_n206), .ZN(new_n218));
  NAND3_X1  g032(.A1(new_n209), .A2(new_n216), .A3(new_n218), .ZN(new_n219));
  INV_X1    g033(.A(G146), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n194), .A2(new_n220), .ZN(new_n221));
  NAND3_X1  g035(.A1(new_n198), .A2(new_n219), .A3(new_n221), .ZN(new_n222));
  INV_X1    g036(.A(KEYINPUT76), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n196), .A2(new_n223), .ZN(new_n224));
  OR2_X1    g038(.A1(new_n195), .A2(G146), .ZN(new_n225));
  NAND3_X1  g039(.A1(new_n195), .A2(KEYINPUT76), .A3(G146), .ZN(new_n226));
  NAND3_X1  g040(.A1(new_n224), .A2(new_n225), .A3(new_n226), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n207), .A2(new_n208), .ZN(new_n228));
  OAI211_X1 g042(.A(new_n227), .B(new_n228), .C1(new_n215), .C2(new_n214), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n222), .A2(new_n229), .ZN(new_n230));
  OAI21_X1  g044(.A(new_n191), .B1(new_n230), .B2(KEYINPUT79), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n230), .A2(KEYINPUT79), .ZN(new_n232));
  XNOR2_X1  g046(.A(new_n231), .B(new_n232), .ZN(new_n233));
  OAI21_X1  g047(.A(KEYINPUT25), .B1(new_n233), .B2(G902), .ZN(new_n234));
  INV_X1    g048(.A(G217), .ZN(new_n235));
  INV_X1    g049(.A(G902), .ZN(new_n236));
  AOI21_X1  g050(.A(new_n235), .B1(G234), .B2(new_n236), .ZN(new_n237));
  OR2_X1    g051(.A1(new_n230), .A2(KEYINPUT79), .ZN(new_n238));
  NAND3_X1  g052(.A1(new_n238), .A2(new_n232), .A3(new_n191), .ZN(new_n239));
  NAND3_X1  g053(.A1(new_n230), .A2(KEYINPUT79), .A3(new_n190), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n239), .A2(new_n240), .ZN(new_n241));
  INV_X1    g055(.A(KEYINPUT25), .ZN(new_n242));
  NAND3_X1  g056(.A1(new_n241), .A2(new_n242), .A3(new_n236), .ZN(new_n243));
  NAND3_X1  g057(.A1(new_n234), .A2(new_n237), .A3(new_n243), .ZN(new_n244));
  NOR2_X1   g058(.A1(new_n237), .A2(G902), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n241), .A2(new_n245), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n244), .A2(new_n246), .ZN(new_n247));
  INV_X1    g061(.A(new_n247), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n188), .A2(G227), .ZN(new_n249));
  XNOR2_X1  g063(.A(new_n249), .B(G140), .ZN(new_n250));
  XNOR2_X1  g064(.A(KEYINPUT80), .B(G110), .ZN(new_n251));
  XNOR2_X1  g065(.A(new_n250), .B(new_n251), .ZN(new_n252));
  INV_X1    g066(.A(KEYINPUT84), .ZN(new_n253));
  INV_X1    g067(.A(G104), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n254), .A2(G107), .ZN(new_n255));
  INV_X1    g069(.A(new_n255), .ZN(new_n256));
  NOR2_X1   g070(.A1(new_n254), .A2(G107), .ZN(new_n257));
  OAI21_X1  g071(.A(G101), .B1(new_n256), .B2(new_n257), .ZN(new_n258));
  OAI21_X1  g072(.A(KEYINPUT3), .B1(new_n254), .B2(G107), .ZN(new_n259));
  INV_X1    g073(.A(KEYINPUT3), .ZN(new_n260));
  INV_X1    g074(.A(G107), .ZN(new_n261));
  NAND3_X1  g075(.A1(new_n260), .A2(new_n261), .A3(G104), .ZN(new_n262));
  INV_X1    g076(.A(G101), .ZN(new_n263));
  NAND4_X1  g077(.A1(new_n259), .A2(new_n262), .A3(new_n263), .A4(new_n255), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n258), .A2(new_n264), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n220), .A2(G143), .ZN(new_n266));
  INV_X1    g080(.A(G143), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n267), .A2(G146), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n266), .A2(new_n268), .ZN(new_n269));
  OAI21_X1  g083(.A(KEYINPUT1), .B1(new_n267), .B2(G146), .ZN(new_n270));
  INV_X1    g084(.A(KEYINPUT83), .ZN(new_n271));
  OAI21_X1  g085(.A(G128), .B1(new_n270), .B2(new_n271), .ZN(new_n272));
  INV_X1    g086(.A(KEYINPUT1), .ZN(new_n273));
  AOI21_X1  g087(.A(new_n273), .B1(G143), .B2(new_n220), .ZN(new_n274));
  NOR2_X1   g088(.A1(new_n274), .A2(KEYINPUT83), .ZN(new_n275));
  OAI21_X1  g089(.A(new_n269), .B1(new_n272), .B2(new_n275), .ZN(new_n276));
  AND4_X1   g090(.A1(new_n273), .A2(new_n266), .A3(new_n268), .A4(G128), .ZN(new_n277));
  INV_X1    g091(.A(new_n277), .ZN(new_n278));
  AOI21_X1  g092(.A(new_n265), .B1(new_n276), .B2(new_n278), .ZN(new_n279));
  OAI21_X1  g093(.A(new_n253), .B1(new_n279), .B2(KEYINPUT10), .ZN(new_n280));
  INV_X1    g094(.A(new_n265), .ZN(new_n281));
  XNOR2_X1  g095(.A(G143), .B(G146), .ZN(new_n282));
  AOI21_X1  g096(.A(new_n200), .B1(new_n274), .B2(KEYINPUT83), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n270), .A2(new_n271), .ZN(new_n284));
  AOI21_X1  g098(.A(new_n282), .B1(new_n283), .B2(new_n284), .ZN(new_n285));
  OAI21_X1  g099(.A(new_n281), .B1(new_n285), .B2(new_n277), .ZN(new_n286));
  INV_X1    g100(.A(KEYINPUT10), .ZN(new_n287));
  NAND3_X1  g101(.A1(new_n286), .A2(KEYINPUT84), .A3(new_n287), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n280), .A2(new_n288), .ZN(new_n289));
  NAND3_X1  g103(.A1(new_n259), .A2(new_n262), .A3(new_n255), .ZN(new_n290));
  INV_X1    g104(.A(KEYINPUT82), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  NAND4_X1  g106(.A1(new_n259), .A2(new_n262), .A3(KEYINPUT82), .A4(new_n255), .ZN(new_n293));
  NAND3_X1  g107(.A1(new_n292), .A2(G101), .A3(new_n293), .ZN(new_n294));
  NAND3_X1  g108(.A1(new_n294), .A2(KEYINPUT4), .A3(new_n264), .ZN(new_n295));
  INV_X1    g109(.A(KEYINPUT0), .ZN(new_n296));
  NOR2_X1   g110(.A1(new_n296), .A2(new_n200), .ZN(new_n297));
  NOR2_X1   g111(.A1(KEYINPUT0), .A2(G128), .ZN(new_n298));
  OAI21_X1  g112(.A(new_n269), .B1(new_n297), .B2(new_n298), .ZN(new_n299));
  OAI21_X1  g113(.A(new_n282), .B1(new_n296), .B2(new_n200), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n299), .A2(new_n300), .ZN(new_n301));
  OAI211_X1 g115(.A(new_n295), .B(new_n301), .C1(KEYINPUT4), .C2(new_n294), .ZN(new_n302));
  INV_X1    g116(.A(KEYINPUT65), .ZN(new_n303));
  OAI211_X1 g117(.A(new_n303), .B(KEYINPUT1), .C1(new_n267), .C2(G146), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n304), .A2(G128), .ZN(new_n305));
  AOI21_X1  g119(.A(new_n303), .B1(new_n266), .B2(KEYINPUT1), .ZN(new_n306));
  OAI21_X1  g120(.A(new_n269), .B1(new_n305), .B2(new_n306), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n307), .A2(new_n278), .ZN(new_n308));
  NAND3_X1  g122(.A1(new_n308), .A2(KEYINPUT10), .A3(new_n281), .ZN(new_n309));
  NAND3_X1  g123(.A1(new_n289), .A2(new_n302), .A3(new_n309), .ZN(new_n310));
  INV_X1    g124(.A(KEYINPUT11), .ZN(new_n311));
  INV_X1    g125(.A(G134), .ZN(new_n312));
  OAI21_X1  g126(.A(new_n311), .B1(new_n312), .B2(G137), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n312), .A2(G137), .ZN(new_n314));
  INV_X1    g128(.A(G137), .ZN(new_n315));
  NAND3_X1  g129(.A1(new_n315), .A2(KEYINPUT11), .A3(G134), .ZN(new_n316));
  NAND3_X1  g130(.A1(new_n313), .A2(new_n314), .A3(new_n316), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n317), .A2(G131), .ZN(new_n318));
  INV_X1    g132(.A(G131), .ZN(new_n319));
  NAND4_X1  g133(.A1(new_n313), .A2(new_n316), .A3(new_n319), .A4(new_n314), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n318), .A2(new_n320), .ZN(new_n321));
  AND2_X1   g135(.A1(new_n310), .A2(new_n321), .ZN(new_n322));
  INV_X1    g136(.A(new_n321), .ZN(new_n323));
  NAND4_X1  g137(.A1(new_n289), .A2(new_n302), .A3(new_n323), .A4(new_n309), .ZN(new_n324));
  INV_X1    g138(.A(new_n324), .ZN(new_n325));
  OAI21_X1  g139(.A(new_n252), .B1(new_n322), .B2(new_n325), .ZN(new_n326));
  NOR2_X1   g140(.A1(new_n308), .A2(new_n281), .ZN(new_n327));
  OAI21_X1  g141(.A(new_n321), .B1(new_n327), .B2(new_n279), .ZN(new_n328));
  INV_X1    g142(.A(KEYINPUT12), .ZN(new_n329));
  XNOR2_X1  g143(.A(new_n328), .B(new_n329), .ZN(new_n330));
  INV_X1    g144(.A(new_n252), .ZN(new_n331));
  NAND3_X1  g145(.A1(new_n330), .A2(new_n324), .A3(new_n331), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n326), .A2(new_n332), .ZN(new_n333));
  INV_X1    g147(.A(G469), .ZN(new_n334));
  NAND3_X1  g148(.A1(new_n333), .A2(new_n334), .A3(new_n236), .ZN(new_n335));
  XOR2_X1   g149(.A(new_n252), .B(KEYINPUT81), .Z(new_n336));
  AND3_X1   g150(.A1(new_n330), .A2(KEYINPUT85), .A3(new_n324), .ZN(new_n337));
  AOI21_X1  g151(.A(KEYINPUT85), .B1(new_n330), .B2(new_n324), .ZN(new_n338));
  OAI21_X1  g152(.A(new_n336), .B1(new_n337), .B2(new_n338), .ZN(new_n339));
  OR3_X1    g153(.A1(new_n322), .A2(new_n325), .A3(new_n252), .ZN(new_n340));
  NAND3_X1  g154(.A1(new_n339), .A2(new_n340), .A3(G469), .ZN(new_n341));
  NAND2_X1  g155(.A1(G469), .A2(G902), .ZN(new_n342));
  NAND3_X1  g156(.A1(new_n335), .A2(new_n341), .A3(new_n342), .ZN(new_n343));
  XNOR2_X1  g157(.A(KEYINPUT9), .B(G234), .ZN(new_n344));
  OAI21_X1  g158(.A(G221), .B1(new_n344), .B2(G902), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n343), .A2(new_n345), .ZN(new_n346));
  NOR2_X1   g160(.A1(G237), .A2(G953), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n347), .A2(G214), .ZN(new_n348));
  NAND3_X1  g162(.A1(new_n348), .A2(KEYINPUT88), .A3(G143), .ZN(new_n349));
  OR2_X1    g163(.A1(KEYINPUT88), .A2(G143), .ZN(new_n350));
  NAND2_X1  g164(.A1(KEYINPUT88), .A2(G143), .ZN(new_n351));
  NAND4_X1  g165(.A1(new_n350), .A2(G214), .A3(new_n347), .A4(new_n351), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n349), .A2(new_n352), .ZN(new_n353));
  NOR2_X1   g167(.A1(new_n353), .A2(new_n319), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n354), .A2(KEYINPUT18), .ZN(new_n355));
  INV_X1    g169(.A(KEYINPUT89), .ZN(new_n356));
  XNOR2_X1  g170(.A(new_n194), .B(new_n356), .ZN(new_n357));
  OAI21_X1  g171(.A(new_n221), .B1(new_n357), .B2(new_n220), .ZN(new_n358));
  INV_X1    g172(.A(KEYINPUT18), .ZN(new_n359));
  OAI21_X1  g173(.A(new_n353), .B1(new_n359), .B2(new_n319), .ZN(new_n360));
  NAND3_X1  g174(.A1(new_n355), .A2(new_n358), .A3(new_n360), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n354), .A2(KEYINPUT17), .ZN(new_n362));
  XNOR2_X1  g176(.A(new_n353), .B(new_n319), .ZN(new_n363));
  OAI21_X1  g177(.A(new_n362), .B1(new_n363), .B2(KEYINPUT17), .ZN(new_n364));
  OAI21_X1  g178(.A(new_n361), .B1(new_n364), .B2(new_n227), .ZN(new_n365));
  XNOR2_X1  g179(.A(G113), .B(G122), .ZN(new_n366));
  XNOR2_X1  g180(.A(new_n366), .B(new_n254), .ZN(new_n367));
  INV_X1    g181(.A(new_n367), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n365), .A2(new_n368), .ZN(new_n369));
  OAI211_X1 g183(.A(new_n367), .B(new_n361), .C1(new_n364), .C2(new_n227), .ZN(new_n370));
  AOI21_X1  g184(.A(G902), .B1(new_n369), .B2(new_n370), .ZN(new_n371));
  XOR2_X1   g185(.A(KEYINPUT91), .B(G475), .Z(new_n372));
  NOR2_X1   g186(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  INV_X1    g187(.A(KEYINPUT19), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n194), .A2(new_n374), .ZN(new_n375));
  OAI211_X1 g189(.A(new_n220), .B(new_n375), .C1(new_n357), .C2(new_n374), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n363), .A2(new_n376), .ZN(new_n377));
  XNOR2_X1  g191(.A(new_n196), .B(KEYINPUT78), .ZN(new_n378));
  OAI21_X1  g192(.A(new_n361), .B1(new_n377), .B2(new_n378), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n379), .A2(new_n368), .ZN(new_n380));
  AOI21_X1  g194(.A(G475), .B1(new_n380), .B2(new_n370), .ZN(new_n381));
  INV_X1    g195(.A(KEYINPUT20), .ZN(new_n382));
  NAND3_X1  g196(.A1(new_n381), .A2(new_n382), .A3(new_n236), .ZN(new_n383));
  AOI21_X1  g197(.A(new_n382), .B1(new_n381), .B2(new_n236), .ZN(new_n384));
  OAI21_X1  g198(.A(new_n383), .B1(new_n384), .B2(KEYINPUT90), .ZN(new_n385));
  INV_X1    g199(.A(KEYINPUT90), .ZN(new_n386));
  NAND4_X1  g200(.A1(new_n381), .A2(new_n386), .A3(new_n382), .A4(new_n236), .ZN(new_n387));
  AOI21_X1  g201(.A(new_n373), .B1(new_n385), .B2(new_n387), .ZN(new_n388));
  NAND2_X1  g202(.A1(G234), .A2(G237), .ZN(new_n389));
  NAND3_X1  g203(.A1(new_n389), .A2(G952), .A3(new_n188), .ZN(new_n390));
  INV_X1    g204(.A(new_n390), .ZN(new_n391));
  XOR2_X1   g205(.A(KEYINPUT21), .B(G898), .Z(new_n392));
  INV_X1    g206(.A(new_n392), .ZN(new_n393));
  NAND3_X1  g207(.A1(new_n389), .A2(G902), .A3(G953), .ZN(new_n394));
  INV_X1    g208(.A(new_n394), .ZN(new_n395));
  AOI21_X1  g209(.A(new_n391), .B1(new_n393), .B2(new_n395), .ZN(new_n396));
  INV_X1    g210(.A(new_n396), .ZN(new_n397));
  INV_X1    g211(.A(G478), .ZN(new_n398));
  NOR2_X1   g212(.A1(new_n398), .A2(KEYINPUT15), .ZN(new_n399));
  XNOR2_X1  g213(.A(G128), .B(G143), .ZN(new_n400));
  XNOR2_X1  g214(.A(new_n400), .B(new_n312), .ZN(new_n401));
  XNOR2_X1  g215(.A(G116), .B(G122), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n402), .A2(new_n261), .ZN(new_n403));
  INV_X1    g217(.A(G116), .ZN(new_n404));
  NAND3_X1  g218(.A1(new_n404), .A2(KEYINPUT14), .A3(G122), .ZN(new_n405));
  XOR2_X1   g219(.A(G116), .B(G122), .Z(new_n406));
  OAI211_X1 g220(.A(G107), .B(new_n405), .C1(new_n406), .C2(KEYINPUT14), .ZN(new_n407));
  NAND3_X1  g221(.A1(new_n401), .A2(new_n403), .A3(new_n407), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n406), .A2(G107), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n409), .A2(new_n403), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n400), .A2(new_n312), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n400), .A2(KEYINPUT13), .ZN(new_n412));
  OR3_X1    g226(.A1(new_n200), .A2(KEYINPUT13), .A3(G143), .ZN(new_n413));
  NAND3_X1  g227(.A1(new_n412), .A2(G134), .A3(new_n413), .ZN(new_n414));
  NAND3_X1  g228(.A1(new_n410), .A2(new_n411), .A3(new_n414), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n408), .A2(new_n415), .ZN(new_n416));
  NOR3_X1   g230(.A1(new_n344), .A2(new_n235), .A3(G953), .ZN(new_n417));
  XOR2_X1   g231(.A(new_n416), .B(new_n417), .Z(new_n418));
  NAND2_X1  g232(.A1(new_n418), .A2(new_n236), .ZN(new_n419));
  INV_X1    g233(.A(KEYINPUT92), .ZN(new_n420));
  AOI21_X1  g234(.A(new_n399), .B1(new_n419), .B2(new_n420), .ZN(new_n421));
  XNOR2_X1  g235(.A(new_n419), .B(new_n420), .ZN(new_n422));
  AOI21_X1  g236(.A(new_n421), .B1(new_n422), .B2(new_n399), .ZN(new_n423));
  NAND3_X1  g237(.A1(new_n388), .A2(new_n397), .A3(new_n423), .ZN(new_n424));
  INV_X1    g238(.A(G113), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n425), .A2(KEYINPUT2), .ZN(new_n426));
  INV_X1    g240(.A(KEYINPUT2), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n427), .A2(G113), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n426), .A2(new_n428), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n404), .A2(G119), .ZN(new_n430));
  INV_X1    g244(.A(KEYINPUT67), .ZN(new_n431));
  OAI21_X1  g245(.A(new_n431), .B1(new_n404), .B2(G119), .ZN(new_n432));
  NAND3_X1  g246(.A1(new_n203), .A2(KEYINPUT67), .A3(G116), .ZN(new_n433));
  NAND4_X1  g247(.A1(new_n429), .A2(new_n430), .A3(new_n432), .A4(new_n433), .ZN(new_n434));
  INV_X1    g248(.A(KEYINPUT5), .ZN(new_n435));
  NAND3_X1  g249(.A1(new_n435), .A2(new_n203), .A3(G116), .ZN(new_n436));
  NAND3_X1  g250(.A1(new_n432), .A2(new_n430), .A3(new_n433), .ZN(new_n437));
  OAI21_X1  g251(.A(new_n436), .B1(new_n437), .B2(new_n435), .ZN(new_n438));
  OAI21_X1  g252(.A(new_n434), .B1(new_n438), .B2(new_n425), .ZN(new_n439));
  OR2_X1    g253(.A1(new_n439), .A2(new_n265), .ZN(new_n440));
  OAI21_X1  g254(.A(new_n295), .B1(KEYINPUT4), .B2(new_n294), .ZN(new_n441));
  AND2_X1   g255(.A1(new_n426), .A2(new_n428), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n437), .A2(new_n442), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n443), .A2(new_n434), .ZN(new_n444));
  INV_X1    g258(.A(KEYINPUT68), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n444), .A2(new_n445), .ZN(new_n446));
  NAND3_X1  g260(.A1(new_n443), .A2(new_n434), .A3(KEYINPUT68), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n446), .A2(new_n447), .ZN(new_n448));
  INV_X1    g262(.A(new_n448), .ZN(new_n449));
  OAI21_X1  g263(.A(new_n440), .B1(new_n441), .B2(new_n449), .ZN(new_n450));
  XNOR2_X1  g264(.A(G110), .B(G122), .ZN(new_n451));
  XNOR2_X1  g265(.A(new_n451), .B(KEYINPUT86), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n450), .A2(new_n452), .ZN(new_n453));
  INV_X1    g267(.A(new_n452), .ZN(new_n454));
  OAI211_X1 g268(.A(new_n454), .B(new_n440), .C1(new_n441), .C2(new_n449), .ZN(new_n455));
  NAND3_X1  g269(.A1(new_n453), .A2(KEYINPUT6), .A3(new_n455), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n301), .A2(G125), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n270), .A2(KEYINPUT65), .ZN(new_n458));
  NAND3_X1  g272(.A1(new_n458), .A2(G128), .A3(new_n304), .ZN(new_n459));
  AOI21_X1  g273(.A(new_n277), .B1(new_n459), .B2(new_n269), .ZN(new_n460));
  OAI21_X1  g274(.A(new_n457), .B1(new_n460), .B2(G125), .ZN(new_n461));
  INV_X1    g275(.A(G224), .ZN(new_n462));
  NOR2_X1   g276(.A1(new_n462), .A2(G953), .ZN(new_n463));
  XOR2_X1   g277(.A(new_n461), .B(new_n463), .Z(new_n464));
  INV_X1    g278(.A(KEYINPUT6), .ZN(new_n465));
  NAND3_X1  g279(.A1(new_n450), .A2(new_n465), .A3(new_n452), .ZN(new_n466));
  NAND3_X1  g280(.A1(new_n456), .A2(new_n464), .A3(new_n466), .ZN(new_n467));
  INV_X1    g281(.A(KEYINPUT7), .ZN(new_n468));
  NOR2_X1   g282(.A1(new_n463), .A2(new_n468), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n461), .A2(new_n469), .ZN(new_n470));
  XOR2_X1   g284(.A(new_n470), .B(KEYINPUT87), .Z(new_n471));
  OR2_X1    g285(.A1(new_n461), .A2(new_n469), .ZN(new_n472));
  XNOR2_X1  g286(.A(new_n439), .B(new_n265), .ZN(new_n473));
  XOR2_X1   g287(.A(new_n452), .B(KEYINPUT8), .Z(new_n474));
  NAND2_X1  g288(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  NAND4_X1  g289(.A1(new_n471), .A2(new_n472), .A3(new_n455), .A4(new_n475), .ZN(new_n476));
  NAND3_X1  g290(.A1(new_n467), .A2(new_n236), .A3(new_n476), .ZN(new_n477));
  OAI21_X1  g291(.A(G210), .B1(G237), .B2(G902), .ZN(new_n478));
  INV_X1    g292(.A(new_n478), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n477), .A2(new_n479), .ZN(new_n480));
  NAND4_X1  g294(.A1(new_n467), .A2(new_n476), .A3(new_n236), .A4(new_n478), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  OAI21_X1  g296(.A(G214), .B1(G237), .B2(G902), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  NOR3_X1   g298(.A1(new_n346), .A2(new_n424), .A3(new_n484), .ZN(new_n485));
  NOR2_X1   g299(.A1(G472), .A2(G902), .ZN(new_n486));
  INV_X1    g300(.A(new_n486), .ZN(new_n487));
  INV_X1    g301(.A(KEYINPUT28), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n321), .A2(new_n301), .ZN(new_n489));
  INV_X1    g303(.A(KEYINPUT64), .ZN(new_n490));
  XNOR2_X1  g304(.A(G134), .B(G137), .ZN(new_n491));
  OAI21_X1  g305(.A(new_n490), .B1(new_n491), .B2(new_n319), .ZN(new_n492));
  NOR2_X1   g306(.A1(new_n315), .A2(G134), .ZN(new_n493));
  NOR2_X1   g307(.A1(new_n312), .A2(G137), .ZN(new_n494));
  OAI211_X1 g308(.A(KEYINPUT64), .B(G131), .C1(new_n493), .C2(new_n494), .ZN(new_n495));
  NAND3_X1  g309(.A1(new_n492), .A2(new_n320), .A3(new_n495), .ZN(new_n496));
  OAI21_X1  g310(.A(new_n489), .B1(new_n460), .B2(new_n496), .ZN(new_n497));
  OAI21_X1  g311(.A(new_n488), .B1(new_n497), .B2(new_n448), .ZN(new_n498));
  XNOR2_X1  g312(.A(new_n498), .B(KEYINPUT72), .ZN(new_n499));
  AND3_X1   g313(.A1(new_n492), .A2(new_n320), .A3(new_n495), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n500), .A2(new_n308), .ZN(new_n501));
  NAND4_X1  g315(.A1(new_n501), .A2(new_n446), .A3(new_n447), .A4(new_n489), .ZN(new_n502));
  INV_X1    g316(.A(new_n489), .ZN(new_n503));
  INV_X1    g317(.A(KEYINPUT66), .ZN(new_n504));
  OAI21_X1  g318(.A(new_n504), .B1(new_n460), .B2(new_n496), .ZN(new_n505));
  NAND3_X1  g319(.A1(new_n500), .A2(new_n308), .A3(KEYINPUT66), .ZN(new_n506));
  AOI21_X1  g320(.A(new_n503), .B1(new_n505), .B2(new_n506), .ZN(new_n507));
  OAI21_X1  g321(.A(new_n502), .B1(new_n507), .B2(new_n449), .ZN(new_n508));
  INV_X1    g322(.A(KEYINPUT71), .ZN(new_n509));
  AND3_X1   g323(.A1(new_n508), .A2(new_n509), .A3(KEYINPUT28), .ZN(new_n510));
  AOI21_X1  g324(.A(new_n509), .B1(new_n508), .B2(KEYINPUT28), .ZN(new_n511));
  OAI21_X1  g325(.A(new_n499), .B1(new_n510), .B2(new_n511), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n347), .A2(G210), .ZN(new_n513));
  XNOR2_X1  g327(.A(new_n513), .B(new_n263), .ZN(new_n514));
  XNOR2_X1  g328(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n515));
  XNOR2_X1  g329(.A(new_n514), .B(new_n515), .ZN(new_n516));
  NAND3_X1  g330(.A1(new_n501), .A2(KEYINPUT30), .A3(new_n489), .ZN(new_n517));
  OAI211_X1 g331(.A(new_n448), .B(new_n517), .C1(new_n507), .C2(KEYINPUT30), .ZN(new_n518));
  INV_X1    g332(.A(KEYINPUT31), .ZN(new_n519));
  NOR2_X1   g333(.A1(new_n497), .A2(new_n448), .ZN(new_n520));
  NOR2_X1   g334(.A1(new_n520), .A2(new_n516), .ZN(new_n521));
  NAND3_X1  g335(.A1(new_n518), .A2(new_n519), .A3(new_n521), .ZN(new_n522));
  INV_X1    g336(.A(KEYINPUT70), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  NAND4_X1  g338(.A1(new_n518), .A2(KEYINPUT70), .A3(new_n519), .A4(new_n521), .ZN(new_n525));
  AOI22_X1  g339(.A1(new_n512), .A2(new_n516), .B1(new_n524), .B2(new_n525), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n518), .A2(new_n521), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n527), .A2(KEYINPUT31), .ZN(new_n528));
  INV_X1    g342(.A(KEYINPUT69), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  AOI21_X1  g344(.A(new_n519), .B1(new_n518), .B2(new_n521), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n531), .A2(KEYINPUT69), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n530), .A2(new_n532), .ZN(new_n533));
  AOI21_X1  g347(.A(new_n487), .B1(new_n526), .B2(new_n533), .ZN(new_n534));
  NOR3_X1   g348(.A1(new_n534), .A2(KEYINPUT73), .A3(KEYINPUT32), .ZN(new_n535));
  INV_X1    g349(.A(KEYINPUT32), .ZN(new_n536));
  AOI211_X1 g350(.A(new_n536), .B(new_n487), .C1(new_n526), .C2(new_n533), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n512), .A2(new_n516), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n524), .A2(new_n525), .ZN(new_n539));
  NAND3_X1  g353(.A1(new_n538), .A2(new_n533), .A3(new_n539), .ZN(new_n540));
  AOI21_X1  g354(.A(KEYINPUT32), .B1(new_n540), .B2(new_n486), .ZN(new_n541));
  NOR2_X1   g355(.A1(new_n537), .A2(new_n541), .ZN(new_n542));
  AOI21_X1  g356(.A(new_n535), .B1(new_n542), .B2(KEYINPUT73), .ZN(new_n543));
  INV_X1    g357(.A(G472), .ZN(new_n544));
  INV_X1    g358(.A(KEYINPUT29), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n518), .A2(new_n502), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n546), .A2(new_n516), .ZN(new_n547));
  OAI211_X1 g361(.A(new_n545), .B(new_n547), .C1(new_n512), .C2(new_n516), .ZN(new_n548));
  INV_X1    g362(.A(KEYINPUT72), .ZN(new_n549));
  XNOR2_X1  g363(.A(new_n498), .B(new_n549), .ZN(new_n550));
  INV_X1    g364(.A(new_n497), .ZN(new_n551));
  OR3_X1    g365(.A1(new_n551), .A2(new_n449), .A3(KEYINPUT74), .ZN(new_n552));
  OAI21_X1  g366(.A(KEYINPUT74), .B1(new_n551), .B2(new_n449), .ZN(new_n553));
  NAND3_X1  g367(.A1(new_n552), .A2(new_n502), .A3(new_n553), .ZN(new_n554));
  AOI21_X1  g368(.A(new_n550), .B1(new_n554), .B2(KEYINPUT28), .ZN(new_n555));
  NOR2_X1   g369(.A1(new_n516), .A2(new_n545), .ZN(new_n556));
  AOI21_X1  g370(.A(G902), .B1(new_n555), .B2(new_n556), .ZN(new_n557));
  AOI21_X1  g371(.A(new_n544), .B1(new_n548), .B2(new_n557), .ZN(new_n558));
  OAI211_X1 g372(.A(new_n248), .B(new_n485), .C1(new_n543), .C2(new_n558), .ZN(new_n559));
  XNOR2_X1  g373(.A(new_n559), .B(G101), .ZN(G3));
  NOR3_X1   g374(.A1(new_n460), .A2(new_n496), .A3(new_n504), .ZN(new_n561));
  AOI21_X1  g375(.A(KEYINPUT66), .B1(new_n500), .B2(new_n308), .ZN(new_n562));
  OAI21_X1  g376(.A(new_n489), .B1(new_n561), .B2(new_n562), .ZN(new_n563));
  AOI21_X1  g377(.A(new_n520), .B1(new_n563), .B2(new_n448), .ZN(new_n564));
  OAI21_X1  g378(.A(KEYINPUT71), .B1(new_n564), .B2(new_n488), .ZN(new_n565));
  NAND3_X1  g379(.A1(new_n508), .A2(new_n509), .A3(KEYINPUT28), .ZN(new_n566));
  AOI21_X1  g380(.A(new_n550), .B1(new_n565), .B2(new_n566), .ZN(new_n567));
  INV_X1    g381(.A(new_n516), .ZN(new_n568));
  OAI21_X1  g382(.A(new_n539), .B1(new_n567), .B2(new_n568), .ZN(new_n569));
  XNOR2_X1  g383(.A(new_n531), .B(new_n529), .ZN(new_n570));
  OAI21_X1  g384(.A(new_n486), .B1(new_n569), .B2(new_n570), .ZN(new_n571));
  AOI21_X1  g385(.A(G902), .B1(new_n526), .B2(new_n533), .ZN(new_n572));
  OAI21_X1  g386(.A(new_n571), .B1(new_n572), .B2(new_n544), .ZN(new_n573));
  NOR3_X1   g387(.A1(new_n573), .A2(new_n346), .A3(new_n247), .ZN(new_n574));
  INV_X1    g388(.A(new_n388), .ZN(new_n575));
  NOR2_X1   g389(.A1(new_n398), .A2(new_n236), .ZN(new_n576));
  INV_X1    g390(.A(new_n576), .ZN(new_n577));
  INV_X1    g391(.A(new_n419), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n578), .A2(new_n398), .ZN(new_n579));
  XOR2_X1   g393(.A(new_n418), .B(KEYINPUT33), .Z(new_n580));
  INV_X1    g394(.A(new_n580), .ZN(new_n581));
  OAI211_X1 g395(.A(new_n577), .B(new_n579), .C1(new_n581), .C2(new_n398), .ZN(new_n582));
  INV_X1    g396(.A(new_n582), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n575), .A2(new_n583), .ZN(new_n584));
  NAND3_X1  g398(.A1(new_n482), .A2(new_n483), .A3(new_n397), .ZN(new_n585));
  NOR2_X1   g399(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n574), .A2(new_n586), .ZN(new_n587));
  XOR2_X1   g401(.A(KEYINPUT34), .B(G104), .Z(new_n588));
  XNOR2_X1  g402(.A(new_n587), .B(new_n588), .ZN(G6));
  INV_X1    g403(.A(new_n421), .ZN(new_n590));
  XNOR2_X1  g404(.A(new_n419), .B(KEYINPUT92), .ZN(new_n591));
  INV_X1    g405(.A(new_n399), .ZN(new_n592));
  OAI21_X1  g406(.A(new_n590), .B1(new_n591), .B2(new_n592), .ZN(new_n593));
  INV_X1    g407(.A(new_n373), .ZN(new_n594));
  INV_X1    g408(.A(new_n384), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n595), .A2(new_n383), .ZN(new_n596));
  NAND3_X1  g410(.A1(new_n593), .A2(new_n594), .A3(new_n596), .ZN(new_n597));
  NOR2_X1   g411(.A1(new_n585), .A2(new_n597), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n574), .A2(new_n598), .ZN(new_n599));
  XOR2_X1   g413(.A(KEYINPUT35), .B(G107), .Z(new_n600));
  XNOR2_X1  g414(.A(new_n599), .B(new_n600), .ZN(G9));
  INV_X1    g415(.A(new_n573), .ZN(new_n602));
  NOR2_X1   g416(.A1(new_n191), .A2(KEYINPUT36), .ZN(new_n603));
  XNOR2_X1  g417(.A(new_n230), .B(new_n603), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n604), .A2(new_n245), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n244), .A2(new_n605), .ZN(new_n606));
  NAND3_X1  g420(.A1(new_n485), .A2(new_n602), .A3(new_n606), .ZN(new_n607));
  XNOR2_X1  g421(.A(new_n607), .B(G110), .ZN(new_n608));
  XOR2_X1   g422(.A(KEYINPUT93), .B(KEYINPUT37), .Z(new_n609));
  XNOR2_X1  g423(.A(new_n608), .B(new_n609), .ZN(G12));
  NAND2_X1  g424(.A1(new_n571), .A2(new_n536), .ZN(new_n611));
  NAND3_X1  g425(.A1(new_n540), .A2(KEYINPUT32), .A3(new_n486), .ZN(new_n612));
  NAND3_X1  g426(.A1(new_n611), .A2(KEYINPUT73), .A3(new_n612), .ZN(new_n613));
  INV_X1    g427(.A(KEYINPUT73), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n541), .A2(new_n614), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n613), .A2(new_n615), .ZN(new_n616));
  INV_X1    g430(.A(new_n558), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  XOR2_X1   g432(.A(KEYINPUT94), .B(G900), .Z(new_n619));
  AOI21_X1  g433(.A(new_n391), .B1(new_n619), .B2(new_n395), .ZN(new_n620));
  NOR2_X1   g434(.A1(new_n597), .A2(new_n620), .ZN(new_n621));
  XNOR2_X1  g435(.A(new_n621), .B(KEYINPUT95), .ZN(new_n622));
  NOR2_X1   g436(.A1(new_n346), .A2(new_n484), .ZN(new_n623));
  NAND4_X1  g437(.A1(new_n618), .A2(new_n622), .A3(new_n623), .A4(new_n606), .ZN(new_n624));
  XNOR2_X1  g438(.A(new_n624), .B(G128), .ZN(G30));
  AND2_X1   g439(.A1(new_n343), .A2(new_n345), .ZN(new_n626));
  XOR2_X1   g440(.A(new_n620), .B(KEYINPUT39), .Z(new_n627));
  NAND2_X1  g441(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  XNOR2_X1  g442(.A(new_n628), .B(KEYINPUT97), .ZN(new_n629));
  XOR2_X1   g443(.A(new_n629), .B(KEYINPUT40), .Z(new_n630));
  INV_X1    g444(.A(new_n483), .ZN(new_n631));
  NOR2_X1   g445(.A1(new_n606), .A2(new_n631), .ZN(new_n632));
  OAI21_X1  g446(.A(new_n236), .B1(new_n554), .B2(new_n568), .ZN(new_n633));
  AOI21_X1  g447(.A(new_n516), .B1(new_n518), .B2(new_n502), .ZN(new_n634));
  OAI21_X1  g448(.A(G472), .B1(new_n633), .B2(new_n634), .ZN(new_n635));
  NAND2_X1  g449(.A1(new_n616), .A2(new_n635), .ZN(new_n636));
  XNOR2_X1  g450(.A(KEYINPUT96), .B(KEYINPUT38), .ZN(new_n637));
  XNOR2_X1  g451(.A(new_n482), .B(new_n637), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n575), .A2(new_n593), .ZN(new_n639));
  NOR2_X1   g453(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  NAND4_X1  g454(.A1(new_n630), .A2(new_n632), .A3(new_n636), .A4(new_n640), .ZN(new_n641));
  XNOR2_X1  g455(.A(new_n641), .B(G143), .ZN(G45));
  NOR3_X1   g456(.A1(new_n388), .A2(new_n582), .A3(new_n620), .ZN(new_n643));
  NAND4_X1  g457(.A1(new_n618), .A2(new_n623), .A3(new_n606), .A4(new_n643), .ZN(new_n644));
  XNOR2_X1  g458(.A(new_n644), .B(G146), .ZN(G48));
  AOI21_X1  g459(.A(new_n247), .B1(new_n616), .B2(new_n617), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n333), .A2(new_n236), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n647), .A2(G469), .ZN(new_n648));
  NAND3_X1  g462(.A1(new_n648), .A2(new_n345), .A3(new_n335), .ZN(new_n649));
  XNOR2_X1  g463(.A(new_n649), .B(KEYINPUT98), .ZN(new_n650));
  NAND3_X1  g464(.A1(new_n646), .A2(new_n586), .A3(new_n650), .ZN(new_n651));
  XNOR2_X1  g465(.A(KEYINPUT41), .B(G113), .ZN(new_n652));
  XNOR2_X1  g466(.A(new_n651), .B(new_n652), .ZN(G15));
  NAND3_X1  g467(.A1(new_n646), .A2(new_n598), .A3(new_n650), .ZN(new_n654));
  XOR2_X1   g468(.A(KEYINPUT99), .B(G116), .Z(new_n655));
  XNOR2_X1  g469(.A(new_n654), .B(new_n655), .ZN(G18));
  INV_X1    g470(.A(new_n424), .ZN(new_n657));
  NOR2_X1   g471(.A1(new_n649), .A2(new_n484), .ZN(new_n658));
  NAND4_X1  g472(.A1(new_n618), .A2(new_n657), .A3(new_n606), .A4(new_n658), .ZN(new_n659));
  XNOR2_X1  g473(.A(new_n659), .B(G119), .ZN(G21));
  OAI21_X1  g474(.A(new_n539), .B1(new_n555), .B2(new_n568), .ZN(new_n661));
  OAI21_X1  g475(.A(new_n486), .B1(new_n661), .B2(new_n531), .ZN(new_n662));
  NAND2_X1  g476(.A1(new_n540), .A2(new_n236), .ZN(new_n663));
  XOR2_X1   g477(.A(KEYINPUT100), .B(G472), .Z(new_n664));
  NAND2_X1  g478(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  AND3_X1   g479(.A1(new_n248), .A2(new_n662), .A3(new_n665), .ZN(new_n666));
  INV_X1    g480(.A(new_n585), .ZN(new_n667));
  INV_X1    g481(.A(new_n639), .ZN(new_n668));
  NAND4_X1  g482(.A1(new_n666), .A2(new_n650), .A3(new_n667), .A4(new_n668), .ZN(new_n669));
  XNOR2_X1  g483(.A(KEYINPUT101), .B(G122), .ZN(new_n670));
  XNOR2_X1  g484(.A(new_n669), .B(new_n670), .ZN(G24));
  AND3_X1   g485(.A1(new_n665), .A2(new_n606), .A3(new_n662), .ZN(new_n672));
  NAND3_X1  g486(.A1(new_n672), .A2(new_n643), .A3(new_n658), .ZN(new_n673));
  XNOR2_X1  g487(.A(KEYINPUT102), .B(G125), .ZN(new_n674));
  XNOR2_X1  g488(.A(new_n673), .B(new_n674), .ZN(G27));
  NAND3_X1  g489(.A1(new_n480), .A2(new_n483), .A3(new_n481), .ZN(new_n676));
  NOR2_X1   g490(.A1(new_n346), .A2(new_n676), .ZN(new_n677));
  AND2_X1   g491(.A1(new_n677), .A2(new_n643), .ZN(new_n678));
  NAND2_X1  g492(.A1(new_n646), .A2(new_n678), .ZN(new_n679));
  INV_X1    g493(.A(KEYINPUT42), .ZN(new_n680));
  NAND2_X1  g494(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  AOI21_X1  g495(.A(new_n247), .B1(new_n542), .B2(new_n617), .ZN(new_n682));
  NAND3_X1  g496(.A1(new_n678), .A2(new_n682), .A3(KEYINPUT42), .ZN(new_n683));
  NAND2_X1  g497(.A1(new_n681), .A2(new_n683), .ZN(new_n684));
  XNOR2_X1  g498(.A(new_n684), .B(G131), .ZN(G33));
  NAND4_X1  g499(.A1(new_n618), .A2(new_n622), .A3(new_n248), .A4(new_n677), .ZN(new_n686));
  XOR2_X1   g500(.A(KEYINPUT103), .B(G134), .Z(new_n687));
  XNOR2_X1  g501(.A(new_n686), .B(new_n687), .ZN(G36));
  NAND2_X1  g502(.A1(new_n339), .A2(new_n340), .ZN(new_n689));
  XNOR2_X1  g503(.A(new_n689), .B(KEYINPUT45), .ZN(new_n690));
  NAND2_X1  g504(.A1(new_n690), .A2(G469), .ZN(new_n691));
  NAND2_X1  g505(.A1(new_n691), .A2(new_n342), .ZN(new_n692));
  INV_X1    g506(.A(KEYINPUT46), .ZN(new_n693));
  NAND2_X1  g507(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  INV_X1    g508(.A(KEYINPUT104), .ZN(new_n695));
  NAND2_X1  g509(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  NAND3_X1  g510(.A1(new_n691), .A2(KEYINPUT46), .A3(new_n342), .ZN(new_n697));
  NAND3_X1  g511(.A1(new_n692), .A2(KEYINPUT104), .A3(new_n693), .ZN(new_n698));
  NAND4_X1  g512(.A1(new_n696), .A2(new_n335), .A3(new_n697), .A4(new_n698), .ZN(new_n699));
  AND3_X1   g513(.A1(new_n699), .A2(new_n345), .A3(new_n627), .ZN(new_n700));
  INV_X1    g514(.A(new_n676), .ZN(new_n701));
  NAND2_X1  g515(.A1(new_n573), .A2(new_n606), .ZN(new_n702));
  XOR2_X1   g516(.A(new_n702), .B(KEYINPUT105), .Z(new_n703));
  NAND2_X1  g517(.A1(new_n583), .A2(new_n388), .ZN(new_n704));
  XOR2_X1   g518(.A(new_n704), .B(KEYINPUT43), .Z(new_n705));
  NAND2_X1  g519(.A1(new_n703), .A2(new_n705), .ZN(new_n706));
  INV_X1    g520(.A(KEYINPUT44), .ZN(new_n707));
  NAND2_X1  g521(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  NAND3_X1  g522(.A1(new_n703), .A2(KEYINPUT44), .A3(new_n705), .ZN(new_n709));
  NAND4_X1  g523(.A1(new_n700), .A2(new_n701), .A3(new_n708), .A4(new_n709), .ZN(new_n710));
  XNOR2_X1  g524(.A(new_n710), .B(G137), .ZN(G39));
  NAND2_X1  g525(.A1(new_n699), .A2(new_n345), .ZN(new_n712));
  INV_X1    g526(.A(KEYINPUT47), .ZN(new_n713));
  XNOR2_X1  g527(.A(new_n712), .B(new_n713), .ZN(new_n714));
  NOR3_X1   g528(.A1(new_n618), .A2(new_n248), .A3(new_n676), .ZN(new_n715));
  NAND3_X1  g529(.A1(new_n714), .A2(new_n643), .A3(new_n715), .ZN(new_n716));
  XNOR2_X1  g530(.A(new_n716), .B(G140), .ZN(G42));
  AND2_X1   g531(.A1(new_n648), .A2(new_n335), .ZN(new_n718));
  INV_X1    g532(.A(new_n718), .ZN(new_n719));
  NAND2_X1  g533(.A1(new_n719), .A2(KEYINPUT49), .ZN(new_n720));
  INV_X1    g534(.A(new_n704), .ZN(new_n721));
  NOR2_X1   g535(.A1(new_n247), .A2(new_n631), .ZN(new_n722));
  NAND4_X1  g536(.A1(new_n720), .A2(new_n345), .A3(new_n721), .A4(new_n722), .ZN(new_n723));
  XNOR2_X1  g537(.A(new_n723), .B(KEYINPUT106), .ZN(new_n724));
  INV_X1    g538(.A(new_n636), .ZN(new_n725));
  OR2_X1    g539(.A1(new_n719), .A2(KEYINPUT49), .ZN(new_n726));
  NAND4_X1  g540(.A1(new_n724), .A2(new_n725), .A3(new_n638), .A4(new_n726), .ZN(new_n727));
  INV_X1    g541(.A(KEYINPUT110), .ZN(new_n728));
  NOR2_X1   g542(.A1(new_n606), .A2(new_n620), .ZN(new_n729));
  NOR2_X1   g543(.A1(new_n639), .A2(new_n484), .ZN(new_n730));
  NAND4_X1  g544(.A1(new_n636), .A2(new_n626), .A3(new_n729), .A4(new_n730), .ZN(new_n731));
  NAND4_X1  g545(.A1(new_n624), .A2(new_n644), .A3(new_n731), .A4(new_n673), .ZN(new_n732));
  INV_X1    g546(.A(KEYINPUT52), .ZN(new_n733));
  OAI21_X1  g547(.A(new_n728), .B1(new_n732), .B2(new_n733), .ZN(new_n734));
  INV_X1    g548(.A(KEYINPUT111), .ZN(new_n735));
  NAND3_X1  g549(.A1(new_n732), .A2(new_n735), .A3(new_n733), .ZN(new_n736));
  INV_X1    g550(.A(new_n736), .ZN(new_n737));
  AOI21_X1  g551(.A(new_n735), .B1(new_n732), .B2(new_n733), .ZN(new_n738));
  OAI21_X1  g552(.A(new_n734), .B1(new_n737), .B2(new_n738), .ZN(new_n739));
  NAND2_X1  g553(.A1(new_n732), .A2(new_n733), .ZN(new_n740));
  NAND2_X1  g554(.A1(new_n740), .A2(KEYINPUT111), .ZN(new_n741));
  AND2_X1   g555(.A1(new_n624), .A2(new_n644), .ZN(new_n742));
  NAND4_X1  g556(.A1(new_n742), .A2(KEYINPUT52), .A3(new_n673), .A4(new_n731), .ZN(new_n743));
  NAND4_X1  g557(.A1(new_n741), .A2(new_n728), .A3(new_n743), .A4(new_n736), .ZN(new_n744));
  NAND2_X1  g558(.A1(new_n739), .A2(new_n744), .ZN(new_n745));
  INV_X1    g559(.A(KEYINPUT53), .ZN(new_n746));
  INV_X1    g560(.A(KEYINPUT108), .ZN(new_n747));
  NAND2_X1  g561(.A1(new_n596), .A2(new_n594), .ZN(new_n748));
  OR2_X1    g562(.A1(new_n748), .A2(new_n620), .ZN(new_n749));
  NAND4_X1  g563(.A1(new_n423), .A2(new_n480), .A3(new_n483), .A4(new_n481), .ZN(new_n750));
  OAI21_X1  g564(.A(new_n747), .B1(new_n749), .B2(new_n750), .ZN(new_n751));
  NOR2_X1   g565(.A1(new_n748), .A2(new_n620), .ZN(new_n752));
  NAND4_X1  g566(.A1(new_n701), .A2(new_n752), .A3(KEYINPUT108), .A4(new_n423), .ZN(new_n753));
  NAND2_X1  g567(.A1(new_n751), .A2(new_n753), .ZN(new_n754));
  NAND4_X1  g568(.A1(new_n618), .A2(new_n626), .A3(new_n606), .A4(new_n754), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n686), .A2(new_n755), .ZN(new_n756));
  OAI21_X1  g570(.A(new_n584), .B1(new_n575), .B2(new_n423), .ZN(new_n757));
  NAND3_X1  g571(.A1(new_n574), .A2(new_n667), .A3(new_n757), .ZN(new_n758));
  NAND3_X1  g572(.A1(new_n559), .A2(new_n607), .A3(new_n758), .ZN(new_n759));
  INV_X1    g573(.A(KEYINPUT109), .ZN(new_n760));
  NAND4_X1  g574(.A1(new_n643), .A2(new_n665), .A3(new_n606), .A4(new_n662), .ZN(new_n761));
  NAND2_X1  g575(.A1(new_n626), .A2(new_n701), .ZN(new_n762));
  OAI21_X1  g576(.A(new_n760), .B1(new_n761), .B2(new_n762), .ZN(new_n763));
  NAND4_X1  g577(.A1(new_n672), .A2(KEYINPUT109), .A3(new_n643), .A4(new_n677), .ZN(new_n764));
  AND2_X1   g578(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  NOR3_X1   g579(.A1(new_n756), .A2(new_n759), .A3(new_n765), .ZN(new_n766));
  INV_X1    g580(.A(new_n684), .ZN(new_n767));
  NAND4_X1  g581(.A1(new_n651), .A2(new_n654), .A3(new_n669), .A4(new_n659), .ZN(new_n768));
  OR2_X1    g582(.A1(new_n768), .A2(KEYINPUT107), .ZN(new_n769));
  NAND2_X1  g583(.A1(new_n768), .A2(KEYINPUT107), .ZN(new_n770));
  AOI21_X1  g584(.A(new_n767), .B1(new_n769), .B2(new_n770), .ZN(new_n771));
  NAND4_X1  g585(.A1(new_n745), .A2(new_n746), .A3(new_n766), .A4(new_n771), .ZN(new_n772));
  NAND2_X1  g586(.A1(new_n771), .A2(new_n766), .ZN(new_n773));
  NAND2_X1  g587(.A1(new_n743), .A2(new_n740), .ZN(new_n774));
  INV_X1    g588(.A(new_n774), .ZN(new_n775));
  OAI21_X1  g589(.A(KEYINPUT53), .B1(new_n773), .B2(new_n775), .ZN(new_n776));
  AND2_X1   g590(.A1(new_n772), .A2(new_n776), .ZN(new_n777));
  NAND2_X1  g591(.A1(new_n777), .A2(KEYINPUT54), .ZN(new_n778));
  INV_X1    g592(.A(KEYINPUT54), .ZN(new_n779));
  AND2_X1   g593(.A1(new_n651), .A2(new_n669), .ZN(new_n780));
  NAND4_X1  g594(.A1(new_n684), .A2(new_n780), .A3(new_n654), .A4(new_n659), .ZN(new_n781));
  INV_X1    g595(.A(KEYINPUT112), .ZN(new_n782));
  AND3_X1   g596(.A1(new_n559), .A2(new_n607), .A3(new_n758), .ZN(new_n783));
  NAND3_X1  g597(.A1(new_n783), .A2(new_n686), .A3(new_n755), .ZN(new_n784));
  OAI21_X1  g598(.A(new_n782), .B1(new_n784), .B2(new_n765), .ZN(new_n785));
  NAND2_X1  g599(.A1(new_n766), .A2(KEYINPUT112), .ZN(new_n786));
  AOI21_X1  g600(.A(new_n781), .B1(new_n785), .B2(new_n786), .ZN(new_n787));
  AOI21_X1  g601(.A(new_n746), .B1(new_n745), .B2(new_n787), .ZN(new_n788));
  NAND4_X1  g602(.A1(new_n771), .A2(new_n746), .A3(new_n774), .A4(new_n766), .ZN(new_n789));
  INV_X1    g603(.A(new_n789), .ZN(new_n790));
  OAI21_X1  g604(.A(new_n779), .B1(new_n788), .B2(new_n790), .ZN(new_n791));
  NAND2_X1  g605(.A1(new_n778), .A2(new_n791), .ZN(new_n792));
  AND2_X1   g606(.A1(new_n705), .A2(new_n391), .ZN(new_n793));
  NAND2_X1  g607(.A1(new_n793), .A2(new_n666), .ZN(new_n794));
  INV_X1    g608(.A(new_n794), .ZN(new_n795));
  NOR2_X1   g609(.A1(new_n719), .A2(new_n345), .ZN(new_n796));
  OAI211_X1 g610(.A(new_n701), .B(new_n795), .C1(new_n714), .C2(new_n796), .ZN(new_n797));
  NAND4_X1  g611(.A1(new_n638), .A2(new_n631), .A3(new_n345), .A4(new_n718), .ZN(new_n798));
  XOR2_X1   g612(.A(new_n798), .B(KEYINPUT113), .Z(new_n799));
  NOR2_X1   g613(.A1(new_n799), .A2(new_n794), .ZN(new_n800));
  XNOR2_X1  g614(.A(new_n800), .B(KEYINPUT50), .ZN(new_n801));
  NOR2_X1   g615(.A1(new_n649), .A2(new_n676), .ZN(new_n802));
  NAND3_X1  g616(.A1(new_n793), .A2(new_n672), .A3(new_n802), .ZN(new_n803));
  XOR2_X1   g617(.A(new_n803), .B(KEYINPUT114), .Z(new_n804));
  AND3_X1   g618(.A1(new_n797), .A2(new_n801), .A3(new_n804), .ZN(new_n805));
  NAND4_X1  g619(.A1(new_n725), .A2(new_n248), .A3(new_n391), .A4(new_n802), .ZN(new_n806));
  OR3_X1    g620(.A1(new_n806), .A2(new_n575), .A3(new_n583), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n805), .A2(new_n807), .ZN(new_n808));
  NAND3_X1  g622(.A1(new_n797), .A2(KEYINPUT115), .A3(new_n801), .ZN(new_n809));
  NAND2_X1  g623(.A1(new_n809), .A2(KEYINPUT51), .ZN(new_n810));
  NAND2_X1  g624(.A1(new_n808), .A2(new_n810), .ZN(new_n811));
  NAND3_X1  g625(.A1(new_n793), .A2(new_n682), .A3(new_n802), .ZN(new_n812));
  INV_X1    g626(.A(KEYINPUT48), .ZN(new_n813));
  NAND2_X1  g627(.A1(new_n812), .A2(new_n813), .ZN(new_n814));
  NAND3_X1  g628(.A1(new_n814), .A2(G952), .A3(new_n188), .ZN(new_n815));
  NOR2_X1   g629(.A1(new_n806), .A2(new_n584), .ZN(new_n816));
  NOR2_X1   g630(.A1(new_n812), .A2(new_n813), .ZN(new_n817));
  NOR3_X1   g631(.A1(new_n815), .A2(new_n816), .A3(new_n817), .ZN(new_n818));
  NAND2_X1  g632(.A1(new_n811), .A2(new_n818), .ZN(new_n819));
  NOR3_X1   g633(.A1(new_n794), .A2(new_n484), .A3(new_n649), .ZN(new_n820));
  NOR2_X1   g634(.A1(new_n808), .A2(new_n810), .ZN(new_n821));
  NOR4_X1   g635(.A1(new_n792), .A2(new_n819), .A3(new_n820), .A4(new_n821), .ZN(new_n822));
  NOR2_X1   g636(.A1(G952), .A2(G953), .ZN(new_n823));
  OAI21_X1  g637(.A(new_n727), .B1(new_n822), .B2(new_n823), .ZN(G75));
  NOR2_X1   g638(.A1(new_n767), .A2(new_n768), .ZN(new_n825));
  NOR2_X1   g639(.A1(new_n756), .A2(new_n759), .ZN(new_n826));
  INV_X1    g640(.A(new_n765), .ZN(new_n827));
  AOI21_X1  g641(.A(KEYINPUT112), .B1(new_n826), .B2(new_n827), .ZN(new_n828));
  NOR4_X1   g642(.A1(new_n756), .A2(new_n759), .A3(new_n765), .A4(new_n782), .ZN(new_n829));
  OAI21_X1  g643(.A(new_n825), .B1(new_n828), .B2(new_n829), .ZN(new_n830));
  AOI21_X1  g644(.A(new_n830), .B1(new_n744), .B2(new_n739), .ZN(new_n831));
  OAI211_X1 g645(.A(G902), .B(new_n789), .C1(new_n831), .C2(new_n746), .ZN(new_n832));
  NAND2_X1  g646(.A1(new_n832), .A2(KEYINPUT116), .ZN(new_n833));
  NOR3_X1   g647(.A1(new_n737), .A2(new_n734), .A3(new_n738), .ZN(new_n834));
  AOI22_X1  g648(.A1(new_n741), .A2(new_n736), .B1(new_n728), .B2(new_n743), .ZN(new_n835));
  OAI21_X1  g649(.A(new_n787), .B1(new_n834), .B2(new_n835), .ZN(new_n836));
  NAND2_X1  g650(.A1(new_n836), .A2(KEYINPUT53), .ZN(new_n837));
  INV_X1    g651(.A(KEYINPUT116), .ZN(new_n838));
  NAND4_X1  g652(.A1(new_n837), .A2(new_n838), .A3(G902), .A4(new_n789), .ZN(new_n839));
  NAND3_X1  g653(.A1(new_n833), .A2(new_n479), .A3(new_n839), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n456), .A2(new_n466), .ZN(new_n841));
  XOR2_X1   g655(.A(new_n841), .B(new_n464), .Z(new_n842));
  XNOR2_X1  g656(.A(new_n842), .B(KEYINPUT55), .ZN(new_n843));
  INV_X1    g657(.A(new_n843), .ZN(new_n844));
  XOR2_X1   g658(.A(KEYINPUT117), .B(KEYINPUT56), .Z(new_n845));
  NAND3_X1  g659(.A1(new_n840), .A2(new_n844), .A3(new_n845), .ZN(new_n846));
  NOR2_X1   g660(.A1(new_n188), .A2(G952), .ZN(new_n847));
  INV_X1    g661(.A(KEYINPUT56), .ZN(new_n848));
  INV_X1    g662(.A(G210), .ZN(new_n849));
  OAI21_X1  g663(.A(new_n848), .B1(new_n832), .B2(new_n849), .ZN(new_n850));
  AOI21_X1  g664(.A(new_n847), .B1(new_n850), .B2(new_n843), .ZN(new_n851));
  AND2_X1   g665(.A1(new_n846), .A2(new_n851), .ZN(G51));
  OAI211_X1 g666(.A(KEYINPUT54), .B(new_n789), .C1(new_n831), .C2(new_n746), .ZN(new_n853));
  NAND2_X1  g667(.A1(new_n853), .A2(KEYINPUT118), .ZN(new_n854));
  INV_X1    g668(.A(KEYINPUT118), .ZN(new_n855));
  NAND4_X1  g669(.A1(new_n837), .A2(new_n855), .A3(KEYINPUT54), .A4(new_n789), .ZN(new_n856));
  NAND3_X1  g670(.A1(new_n854), .A2(new_n791), .A3(new_n856), .ZN(new_n857));
  XOR2_X1   g671(.A(new_n342), .B(KEYINPUT57), .Z(new_n858));
  NAND2_X1  g672(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  NAND2_X1  g673(.A1(new_n859), .A2(new_n333), .ZN(new_n860));
  NAND4_X1  g674(.A1(new_n833), .A2(new_n839), .A3(G469), .A4(new_n690), .ZN(new_n861));
  AOI21_X1  g675(.A(new_n847), .B1(new_n860), .B2(new_n861), .ZN(G54));
  AND2_X1   g676(.A1(KEYINPUT58), .A2(G475), .ZN(new_n863));
  NAND3_X1  g677(.A1(new_n833), .A2(new_n839), .A3(new_n863), .ZN(new_n864));
  NAND2_X1  g678(.A1(new_n380), .A2(new_n370), .ZN(new_n865));
  INV_X1    g679(.A(new_n865), .ZN(new_n866));
  NAND2_X1  g680(.A1(new_n864), .A2(new_n866), .ZN(new_n867));
  INV_X1    g681(.A(new_n847), .ZN(new_n868));
  NAND4_X1  g682(.A1(new_n833), .A2(new_n839), .A3(new_n865), .A4(new_n863), .ZN(new_n869));
  NAND3_X1  g683(.A1(new_n867), .A2(new_n868), .A3(new_n869), .ZN(new_n870));
  NAND2_X1  g684(.A1(new_n870), .A2(KEYINPUT119), .ZN(new_n871));
  INV_X1    g685(.A(KEYINPUT119), .ZN(new_n872));
  NAND4_X1  g686(.A1(new_n867), .A2(new_n872), .A3(new_n868), .A4(new_n869), .ZN(new_n873));
  NAND2_X1  g687(.A1(new_n871), .A2(new_n873), .ZN(G60));
  INV_X1    g688(.A(KEYINPUT120), .ZN(new_n875));
  XNOR2_X1  g689(.A(new_n576), .B(KEYINPUT59), .ZN(new_n876));
  NOR2_X1   g690(.A1(new_n580), .A2(new_n876), .ZN(new_n877));
  NAND2_X1  g691(.A1(new_n857), .A2(new_n877), .ZN(new_n878));
  AOI21_X1  g692(.A(new_n875), .B1(new_n878), .B2(new_n868), .ZN(new_n879));
  AOI211_X1 g693(.A(KEYINPUT120), .B(new_n847), .C1(new_n857), .C2(new_n877), .ZN(new_n880));
  INV_X1    g694(.A(new_n876), .ZN(new_n881));
  AOI21_X1  g695(.A(new_n581), .B1(new_n792), .B2(new_n881), .ZN(new_n882));
  NOR3_X1   g696(.A1(new_n879), .A2(new_n880), .A3(new_n882), .ZN(G63));
  NOR2_X1   g697(.A1(new_n788), .A2(new_n790), .ZN(new_n884));
  NAND2_X1  g698(.A1(G217), .A2(G902), .ZN(new_n885));
  XOR2_X1   g699(.A(new_n885), .B(KEYINPUT60), .Z(new_n886));
  NAND3_X1  g700(.A1(new_n884), .A2(new_n604), .A3(new_n886), .ZN(new_n887));
  AND2_X1   g701(.A1(new_n884), .A2(new_n886), .ZN(new_n888));
  OAI211_X1 g702(.A(new_n868), .B(new_n887), .C1(new_n888), .C2(new_n241), .ZN(new_n889));
  INV_X1    g703(.A(KEYINPUT61), .ZN(new_n890));
  XNOR2_X1  g704(.A(new_n889), .B(new_n890), .ZN(G66));
  OAI21_X1  g705(.A(G953), .B1(new_n393), .B2(new_n462), .ZN(new_n892));
  NAND2_X1  g706(.A1(new_n769), .A2(new_n770), .ZN(new_n893));
  NAND2_X1  g707(.A1(new_n893), .A2(new_n783), .ZN(new_n894));
  XOR2_X1   g708(.A(new_n894), .B(KEYINPUT121), .Z(new_n895));
  INV_X1    g709(.A(new_n895), .ZN(new_n896));
  OAI21_X1  g710(.A(new_n892), .B1(new_n896), .B2(G953), .ZN(new_n897));
  OAI21_X1  g711(.A(new_n841), .B1(G898), .B2(new_n188), .ZN(new_n898));
  XNOR2_X1  g712(.A(new_n897), .B(new_n898), .ZN(G69));
  AOI21_X1  g713(.A(new_n188), .B1(G227), .B2(G900), .ZN(new_n900));
  INV_X1    g714(.A(KEYINPUT124), .ZN(new_n901));
  NAND2_X1  g715(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  XOR2_X1   g716(.A(new_n902), .B(KEYINPUT125), .Z(new_n903));
  INV_X1    g717(.A(new_n629), .ZN(new_n904));
  NAND4_X1  g718(.A1(new_n904), .A2(new_n646), .A3(new_n701), .A4(new_n757), .ZN(new_n905));
  NAND2_X1  g719(.A1(new_n710), .A2(new_n905), .ZN(new_n906));
  INV_X1    g720(.A(KEYINPUT123), .ZN(new_n907));
  XNOR2_X1  g721(.A(new_n906), .B(new_n907), .ZN(new_n908));
  NAND2_X1  g722(.A1(new_n908), .A2(new_n716), .ZN(new_n909));
  AND2_X1   g723(.A1(new_n742), .A2(new_n673), .ZN(new_n910));
  NAND2_X1  g724(.A1(KEYINPUT122), .A2(KEYINPUT62), .ZN(new_n911));
  NAND3_X1  g725(.A1(new_n641), .A2(new_n910), .A3(new_n911), .ZN(new_n912));
  NOR2_X1   g726(.A1(KEYINPUT122), .A2(KEYINPUT62), .ZN(new_n913));
  XOR2_X1   g727(.A(new_n912), .B(new_n913), .Z(new_n914));
  OAI21_X1  g728(.A(new_n188), .B1(new_n909), .B2(new_n914), .ZN(new_n915));
  MUX2_X1   g729(.A(new_n507), .B(new_n497), .S(KEYINPUT30), .Z(new_n916));
  OAI21_X1  g730(.A(new_n375), .B1(new_n357), .B2(new_n374), .ZN(new_n917));
  XOR2_X1   g731(.A(new_n916), .B(new_n917), .Z(new_n918));
  INV_X1    g732(.A(new_n918), .ZN(new_n919));
  NAND2_X1  g733(.A1(new_n915), .A2(new_n919), .ZN(new_n920));
  NAND2_X1  g734(.A1(G900), .A2(G953), .ZN(new_n921));
  NAND3_X1  g735(.A1(new_n700), .A2(new_n682), .A3(new_n730), .ZN(new_n922));
  AND3_X1   g736(.A1(new_n716), .A2(new_n710), .A3(new_n922), .ZN(new_n923));
  NAND4_X1  g737(.A1(new_n923), .A2(new_n684), .A3(new_n686), .A4(new_n910), .ZN(new_n924));
  OAI211_X1 g738(.A(new_n918), .B(new_n921), .C1(new_n924), .C2(G953), .ZN(new_n925));
  NAND2_X1  g739(.A1(new_n920), .A2(new_n925), .ZN(new_n926));
  NOR2_X1   g740(.A1(new_n900), .A2(new_n901), .ZN(new_n927));
  INV_X1    g741(.A(new_n927), .ZN(new_n928));
  AOI21_X1  g742(.A(new_n903), .B1(new_n926), .B2(new_n928), .ZN(new_n929));
  INV_X1    g743(.A(new_n903), .ZN(new_n930));
  AOI211_X1 g744(.A(new_n927), .B(new_n930), .C1(new_n920), .C2(new_n925), .ZN(new_n931));
  NOR2_X1   g745(.A1(new_n929), .A2(new_n931), .ZN(G72));
  NAND2_X1  g746(.A1(new_n546), .A2(new_n568), .ZN(new_n933));
  XNOR2_X1  g747(.A(KEYINPUT126), .B(KEYINPUT63), .ZN(new_n934));
  NOR2_X1   g748(.A1(new_n544), .A2(new_n236), .ZN(new_n935));
  XOR2_X1   g749(.A(new_n934), .B(new_n935), .Z(new_n936));
  NOR2_X1   g750(.A1(new_n546), .A2(new_n568), .ZN(new_n937));
  INV_X1    g751(.A(new_n937), .ZN(new_n938));
  NAND4_X1  g752(.A1(new_n777), .A2(new_n933), .A3(new_n936), .A4(new_n938), .ZN(new_n939));
  INV_X1    g753(.A(KEYINPUT127), .ZN(new_n940));
  XNOR2_X1  g754(.A(new_n939), .B(new_n940), .ZN(new_n941));
  OR2_X1    g755(.A1(new_n909), .A2(new_n914), .ZN(new_n942));
  OAI21_X1  g756(.A(new_n936), .B1(new_n942), .B2(new_n895), .ZN(new_n943));
  NAND2_X1  g757(.A1(new_n943), .A2(new_n634), .ZN(new_n944));
  OAI21_X1  g758(.A(new_n936), .B1(new_n924), .B2(new_n895), .ZN(new_n945));
  AOI21_X1  g759(.A(new_n847), .B1(new_n945), .B2(new_n937), .ZN(new_n946));
  AND3_X1   g760(.A1(new_n941), .A2(new_n944), .A3(new_n946), .ZN(G57));
endmodule


