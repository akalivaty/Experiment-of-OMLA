//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 1 1 0 1 1 0 1 0 0 1 0 0 1 1 1 1 1 0 0 0 1 1 0 1 1 0 0 0 1 0 1 0 0 0 1 1 0 1 1 0 1 0 0 1 0 1 1 0 1 0 0 0 1 1 1 1 1 1 0 1 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:30:00 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n447, new_n451, new_n452, new_n453, new_n454, new_n455,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n531, new_n532,
    new_n533, new_n534, new_n535, new_n536, new_n537, new_n538, new_n540,
    new_n541, new_n542, new_n543, new_n544, new_n545, new_n546, new_n547,
    new_n548, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n558, new_n559, new_n560, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n570, new_n574, new_n575, new_n577,
    new_n578, new_n579, new_n580, new_n581, new_n582, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n603, new_n604, new_n607, new_n608, new_n610, new_n611, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1163, new_n1164, new_n1165, new_n1166,
    new_n1167, new_n1168, new_n1169, new_n1170;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(new_n442));
  XOR2_X1   g017(.A(new_n442), .B(KEYINPUT64), .Z(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n451));
  XNOR2_X1  g026(.A(new_n451), .B(KEYINPUT2), .ZN(new_n452));
  INV_X1    g027(.A(new_n452), .ZN(new_n453));
  NOR4_X1   g028(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n453), .A2(new_n455), .ZN(G325));
  INV_X1    g031(.A(G325), .ZN(G261));
  AOI22_X1  g032(.A1(new_n453), .A2(G2106), .B1(G567), .B2(new_n455), .ZN(G319));
  INV_X1    g033(.A(KEYINPUT65), .ZN(new_n459));
  INV_X1    g034(.A(G2105), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  NAND2_X1  g036(.A1(KEYINPUT65), .A2(G2105), .ZN(new_n462));
  AND2_X1   g037(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n463));
  NOR2_X1   g038(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n464));
  OAI211_X1 g039(.A(new_n461), .B(new_n462), .C1(new_n463), .C2(new_n464), .ZN(new_n465));
  INV_X1    g040(.A(G137), .ZN(new_n466));
  INV_X1    g041(.A(G101), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n460), .A2(G2104), .ZN(new_n468));
  OAI22_X1  g043(.A1(new_n465), .A2(new_n466), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  AND2_X1   g044(.A1(KEYINPUT65), .A2(G2105), .ZN(new_n470));
  NOR2_X1   g045(.A1(KEYINPUT65), .A2(G2105), .ZN(new_n471));
  NOR2_X1   g046(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  OAI21_X1  g047(.A(G125), .B1(new_n463), .B2(new_n464), .ZN(new_n473));
  NAND2_X1  g048(.A1(G113), .A2(G2104), .ZN(new_n474));
  AOI21_X1  g049(.A(new_n472), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  NOR2_X1   g050(.A1(new_n469), .A2(new_n475), .ZN(G160));
  NOR2_X1   g051(.A1(new_n472), .A2(G112), .ZN(new_n477));
  OAI21_X1  g052(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n478));
  XNOR2_X1  g053(.A(KEYINPUT3), .B(G2104), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n479), .A2(new_n460), .ZN(new_n480));
  INV_X1    g055(.A(G136), .ZN(new_n481));
  OAI22_X1  g056(.A1(new_n477), .A2(new_n478), .B1(new_n480), .B2(new_n481), .ZN(new_n482));
  OAI22_X1  g057(.A1(new_n464), .A2(new_n463), .B1(new_n470), .B2(new_n471), .ZN(new_n483));
  INV_X1    g058(.A(KEYINPUT66), .ZN(new_n484));
  XNOR2_X1  g059(.A(new_n483), .B(new_n484), .ZN(new_n485));
  AOI21_X1  g060(.A(new_n482), .B1(new_n485), .B2(G124), .ZN(G162));
  INV_X1    g061(.A(KEYINPUT69), .ZN(new_n487));
  NOR2_X1   g062(.A1(new_n487), .A2(KEYINPUT4), .ZN(new_n488));
  INV_X1    g063(.A(G138), .ZN(new_n489));
  AOI21_X1  g064(.A(new_n489), .B1(new_n487), .B2(KEYINPUT4), .ZN(new_n490));
  INV_X1    g065(.A(new_n490), .ZN(new_n491));
  OAI21_X1  g066(.A(new_n488), .B1(new_n465), .B2(new_n491), .ZN(new_n492));
  INV_X1    g067(.A(new_n488), .ZN(new_n493));
  NAND4_X1  g068(.A1(new_n472), .A2(new_n479), .A3(new_n493), .A4(new_n490), .ZN(new_n494));
  NAND2_X1  g069(.A1(new_n492), .A2(new_n494), .ZN(new_n495));
  OAI21_X1  g070(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n496));
  INV_X1    g071(.A(G114), .ZN(new_n497));
  AOI21_X1  g072(.A(new_n496), .B1(new_n497), .B2(G2105), .ZN(new_n498));
  INV_X1    g073(.A(new_n498), .ZN(new_n499));
  INV_X1    g074(.A(KEYINPUT67), .ZN(new_n500));
  AND2_X1   g075(.A1(G126), .A2(G2105), .ZN(new_n501));
  AOI21_X1  g076(.A(new_n500), .B1(new_n479), .B2(new_n501), .ZN(new_n502));
  OAI211_X1 g077(.A(new_n500), .B(new_n501), .C1(new_n463), .C2(new_n464), .ZN(new_n503));
  INV_X1    g078(.A(new_n503), .ZN(new_n504));
  OAI21_X1  g079(.A(new_n499), .B1(new_n502), .B2(new_n504), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n505), .A2(KEYINPUT68), .ZN(new_n506));
  OAI21_X1  g081(.A(new_n501), .B1(new_n463), .B2(new_n464), .ZN(new_n507));
  NAND2_X1  g082(.A1(new_n507), .A2(KEYINPUT67), .ZN(new_n508));
  AOI21_X1  g083(.A(new_n498), .B1(new_n508), .B2(new_n503), .ZN(new_n509));
  INV_X1    g084(.A(KEYINPUT68), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  AOI21_X1  g086(.A(new_n495), .B1(new_n506), .B2(new_n511), .ZN(G164));
  INV_X1    g087(.A(G543), .ZN(new_n513));
  OR2_X1    g088(.A1(KEYINPUT6), .A2(G651), .ZN(new_n514));
  NAND2_X1  g089(.A1(KEYINPUT6), .A2(G651), .ZN(new_n515));
  AOI21_X1  g090(.A(new_n513), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n516), .A2(G50), .ZN(new_n517));
  NAND2_X1  g092(.A1(KEYINPUT70), .A2(G543), .ZN(new_n518));
  INV_X1    g093(.A(KEYINPUT5), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  NAND3_X1  g095(.A1(KEYINPUT70), .A2(KEYINPUT5), .A3(G543), .ZN(new_n521));
  AOI22_X1  g096(.A1(new_n520), .A2(new_n521), .B1(new_n514), .B2(new_n515), .ZN(new_n522));
  INV_X1    g097(.A(new_n522), .ZN(new_n523));
  XNOR2_X1  g098(.A(KEYINPUT71), .B(G88), .ZN(new_n524));
  OAI21_X1  g099(.A(new_n517), .B1(new_n523), .B2(new_n524), .ZN(new_n525));
  NAND2_X1  g100(.A1(new_n520), .A2(new_n521), .ZN(new_n526));
  AOI22_X1  g101(.A1(new_n526), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n527));
  INV_X1    g102(.A(G651), .ZN(new_n528));
  NOR2_X1   g103(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  NOR2_X1   g104(.A1(new_n525), .A2(new_n529), .ZN(G166));
  NAND3_X1  g105(.A1(new_n526), .A2(G63), .A3(G651), .ZN(new_n531));
  NAND2_X1  g106(.A1(new_n516), .A2(G51), .ZN(new_n532));
  NAND3_X1  g107(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n533));
  XNOR2_X1  g108(.A(new_n533), .B(KEYINPUT7), .ZN(new_n534));
  INV_X1    g109(.A(G89), .ZN(new_n535));
  OAI21_X1  g110(.A(new_n534), .B1(new_n523), .B2(new_n535), .ZN(new_n536));
  OAI211_X1 g111(.A(new_n531), .B(new_n532), .C1(new_n536), .C2(KEYINPUT72), .ZN(new_n537));
  AND2_X1   g112(.A1(new_n536), .A2(KEYINPUT72), .ZN(new_n538));
  NOR2_X1   g113(.A1(new_n537), .A2(new_n538), .ZN(G168));
  NAND2_X1  g114(.A1(G77), .A2(G543), .ZN(new_n540));
  AND2_X1   g115(.A1(new_n520), .A2(new_n521), .ZN(new_n541));
  INV_X1    g116(.A(G64), .ZN(new_n542));
  OAI21_X1  g117(.A(new_n540), .B1(new_n541), .B2(new_n542), .ZN(new_n543));
  AOI21_X1  g118(.A(new_n528), .B1(new_n543), .B2(KEYINPUT73), .ZN(new_n544));
  OAI21_X1  g119(.A(new_n544), .B1(KEYINPUT73), .B2(new_n543), .ZN(new_n545));
  XOR2_X1   g120(.A(KEYINPUT74), .B(G52), .Z(new_n546));
  AOI22_X1  g121(.A1(new_n522), .A2(G90), .B1(new_n516), .B2(new_n546), .ZN(new_n547));
  NAND2_X1  g122(.A1(new_n545), .A2(new_n547), .ZN(new_n548));
  INV_X1    g123(.A(new_n548), .ZN(G171));
  NAND2_X1  g124(.A1(new_n516), .A2(G43), .ZN(new_n550));
  INV_X1    g125(.A(G81), .ZN(new_n551));
  OAI21_X1  g126(.A(new_n550), .B1(new_n523), .B2(new_n551), .ZN(new_n552));
  AOI22_X1  g127(.A1(new_n526), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n553));
  NOR2_X1   g128(.A1(new_n553), .A2(new_n528), .ZN(new_n554));
  NOR2_X1   g129(.A1(new_n552), .A2(new_n554), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n555), .A2(G860), .ZN(G153));
  NAND4_X1  g131(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g132(.A1(G1), .A2(G3), .ZN(new_n558));
  XNOR2_X1  g133(.A(new_n558), .B(KEYINPUT75), .ZN(new_n559));
  XNOR2_X1  g134(.A(new_n559), .B(KEYINPUT8), .ZN(new_n560));
  NAND4_X1  g135(.A1(G319), .A2(G483), .A3(G661), .A4(new_n560), .ZN(G188));
  NAND2_X1  g136(.A1(new_n516), .A2(G53), .ZN(new_n562));
  XNOR2_X1  g137(.A(new_n562), .B(KEYINPUT9), .ZN(new_n563));
  AOI22_X1  g138(.A1(new_n526), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n564));
  OR2_X1    g139(.A1(new_n564), .A2(new_n528), .ZN(new_n565));
  AND2_X1   g140(.A1(new_n563), .A2(new_n565), .ZN(new_n566));
  AND2_X1   g141(.A1(new_n522), .A2(G91), .ZN(new_n567));
  XNOR2_X1  g142(.A(new_n567), .B(KEYINPUT76), .ZN(new_n568));
  NAND2_X1  g143(.A1(new_n566), .A2(new_n568), .ZN(G299));
  XNOR2_X1  g144(.A(new_n548), .B(KEYINPUT77), .ZN(new_n570));
  INV_X1    g145(.A(new_n570), .ZN(G301));
  INV_X1    g146(.A(G168), .ZN(G286));
  INV_X1    g147(.A(G166), .ZN(G303));
  AOI22_X1  g148(.A1(new_n522), .A2(G87), .B1(new_n516), .B2(G49), .ZN(new_n574));
  OAI21_X1  g149(.A(G651), .B1(new_n526), .B2(G74), .ZN(new_n575));
  NAND2_X1  g150(.A1(new_n574), .A2(new_n575), .ZN(G288));
  AOI22_X1  g151(.A1(new_n522), .A2(G86), .B1(new_n516), .B2(G48), .ZN(new_n577));
  INV_X1    g152(.A(G61), .ZN(new_n578));
  AOI21_X1  g153(.A(new_n578), .B1(new_n520), .B2(new_n521), .ZN(new_n579));
  AND2_X1   g154(.A1(G73), .A2(G543), .ZN(new_n580));
  OAI21_X1  g155(.A(G651), .B1(new_n579), .B2(new_n580), .ZN(new_n581));
  NAND2_X1  g156(.A1(new_n577), .A2(new_n581), .ZN(new_n582));
  XNOR2_X1  g157(.A(new_n582), .B(KEYINPUT78), .ZN(G305));
  NAND2_X1  g158(.A1(new_n516), .A2(G47), .ZN(new_n584));
  INV_X1    g159(.A(G85), .ZN(new_n585));
  OAI21_X1  g160(.A(new_n584), .B1(new_n523), .B2(new_n585), .ZN(new_n586));
  AOI22_X1  g161(.A1(new_n526), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n587));
  NOR2_X1   g162(.A1(new_n587), .A2(new_n528), .ZN(new_n588));
  NOR2_X1   g163(.A1(new_n586), .A2(new_n588), .ZN(new_n589));
  INV_X1    g164(.A(new_n589), .ZN(G290));
  NAND2_X1  g165(.A1(new_n522), .A2(G92), .ZN(new_n591));
  INV_X1    g166(.A(KEYINPUT10), .ZN(new_n592));
  XNOR2_X1  g167(.A(new_n591), .B(new_n592), .ZN(new_n593));
  NAND2_X1  g168(.A1(G79), .A2(G543), .ZN(new_n594));
  XNOR2_X1  g169(.A(new_n594), .B(KEYINPUT79), .ZN(new_n595));
  INV_X1    g170(.A(G66), .ZN(new_n596));
  OAI21_X1  g171(.A(new_n595), .B1(new_n541), .B2(new_n596), .ZN(new_n597));
  AOI22_X1  g172(.A1(new_n597), .A2(G651), .B1(G54), .B2(new_n516), .ZN(new_n598));
  NAND2_X1  g173(.A1(new_n593), .A2(new_n598), .ZN(new_n599));
  NOR2_X1   g174(.A1(new_n599), .A2(G868), .ZN(new_n600));
  AOI21_X1  g175(.A(new_n600), .B1(new_n570), .B2(G868), .ZN(G284));
  AOI21_X1  g176(.A(new_n600), .B1(new_n570), .B2(G868), .ZN(G321));
  INV_X1    g177(.A(G868), .ZN(new_n603));
  NAND2_X1  g178(.A1(G299), .A2(new_n603), .ZN(new_n604));
  OAI21_X1  g179(.A(new_n604), .B1(new_n603), .B2(G168), .ZN(G297));
  OAI21_X1  g180(.A(new_n604), .B1(new_n603), .B2(G168), .ZN(G280));
  INV_X1    g181(.A(new_n599), .ZN(new_n607));
  INV_X1    g182(.A(G559), .ZN(new_n608));
  OAI21_X1  g183(.A(new_n607), .B1(new_n608), .B2(G860), .ZN(G148));
  NAND2_X1  g184(.A1(new_n607), .A2(new_n608), .ZN(new_n610));
  NAND2_X1  g185(.A1(new_n610), .A2(G868), .ZN(new_n611));
  OAI21_X1  g186(.A(new_n611), .B1(G868), .B2(new_n555), .ZN(G323));
  XNOR2_X1  g187(.A(G323), .B(KEYINPUT11), .ZN(G282));
  INV_X1    g188(.A(new_n480), .ZN(new_n614));
  NAND2_X1  g189(.A1(new_n614), .A2(G135), .ZN(new_n615));
  NOR2_X1   g190(.A1(new_n472), .A2(G111), .ZN(new_n616));
  OAI21_X1  g191(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n617));
  XNOR2_X1  g192(.A(new_n483), .B(KEYINPUT66), .ZN(new_n618));
  INV_X1    g193(.A(G123), .ZN(new_n619));
  OAI221_X1 g194(.A(new_n615), .B1(new_n616), .B2(new_n617), .C1(new_n618), .C2(new_n619), .ZN(new_n620));
  OR2_X1    g195(.A1(new_n620), .A2(G2096), .ZN(new_n621));
  NAND3_X1  g196(.A1(new_n460), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n622));
  XNOR2_X1  g197(.A(new_n622), .B(KEYINPUT12), .ZN(new_n623));
  XNOR2_X1  g198(.A(new_n623), .B(KEYINPUT13), .ZN(new_n624));
  INV_X1    g199(.A(new_n624), .ZN(new_n625));
  OR2_X1    g200(.A1(new_n625), .A2(G2100), .ZN(new_n626));
  NAND2_X1  g201(.A1(new_n625), .A2(G2100), .ZN(new_n627));
  NAND2_X1  g202(.A1(new_n620), .A2(G2096), .ZN(new_n628));
  NAND4_X1  g203(.A1(new_n621), .A2(new_n626), .A3(new_n627), .A4(new_n628), .ZN(G156));
  XOR2_X1   g204(.A(KEYINPUT15), .B(G2435), .Z(new_n630));
  XNOR2_X1  g205(.A(new_n630), .B(G2438), .ZN(new_n631));
  XOR2_X1   g206(.A(G2427), .B(G2430), .Z(new_n632));
  OR2_X1    g207(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  XNOR2_X1  g208(.A(KEYINPUT81), .B(KEYINPUT14), .ZN(new_n634));
  NAND2_X1  g209(.A1(new_n631), .A2(new_n632), .ZN(new_n635));
  NAND3_X1  g210(.A1(new_n633), .A2(new_n634), .A3(new_n635), .ZN(new_n636));
  XOR2_X1   g211(.A(G1341), .B(G1348), .Z(new_n637));
  XNOR2_X1  g212(.A(KEYINPUT80), .B(KEYINPUT16), .ZN(new_n638));
  XNOR2_X1  g213(.A(new_n637), .B(new_n638), .ZN(new_n639));
  XNOR2_X1  g214(.A(new_n636), .B(new_n639), .ZN(new_n640));
  INV_X1    g215(.A(new_n640), .ZN(new_n641));
  XOR2_X1   g216(.A(G2443), .B(G2446), .Z(new_n642));
  XNOR2_X1  g217(.A(G2451), .B(G2454), .ZN(new_n643));
  XNOR2_X1  g218(.A(new_n642), .B(new_n643), .ZN(new_n644));
  INV_X1    g219(.A(new_n644), .ZN(new_n645));
  OAI21_X1  g220(.A(G14), .B1(new_n641), .B2(new_n645), .ZN(new_n646));
  AOI21_X1  g221(.A(new_n646), .B1(new_n645), .B2(new_n641), .ZN(G401));
  XOR2_X1   g222(.A(G2084), .B(G2090), .Z(new_n648));
  XNOR2_X1  g223(.A(new_n648), .B(KEYINPUT82), .ZN(new_n649));
  XNOR2_X1  g224(.A(G2067), .B(G2678), .ZN(new_n650));
  NAND2_X1  g225(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  NAND2_X1  g226(.A1(new_n651), .A2(KEYINPUT18), .ZN(new_n652));
  XNOR2_X1  g227(.A(G2072), .B(G2078), .ZN(new_n653));
  NAND2_X1  g228(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  XOR2_X1   g229(.A(G2096), .B(G2100), .Z(new_n655));
  XNOR2_X1  g230(.A(new_n655), .B(KEYINPUT83), .ZN(new_n656));
  XNOR2_X1  g231(.A(new_n654), .B(new_n656), .ZN(new_n657));
  AND2_X1   g232(.A1(new_n651), .A2(KEYINPUT17), .ZN(new_n658));
  OR2_X1    g233(.A1(new_n649), .A2(new_n650), .ZN(new_n659));
  AOI21_X1  g234(.A(KEYINPUT18), .B1(new_n658), .B2(new_n659), .ZN(new_n660));
  XNOR2_X1  g235(.A(new_n657), .B(new_n660), .ZN(G227));
  XOR2_X1   g236(.A(G1971), .B(G1976), .Z(new_n662));
  XNOR2_X1  g237(.A(new_n662), .B(KEYINPUT19), .ZN(new_n663));
  XNOR2_X1  g238(.A(G1956), .B(G2474), .ZN(new_n664));
  XNOR2_X1  g239(.A(G1961), .B(G1966), .ZN(new_n665));
  NOR2_X1   g240(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  AND2_X1   g241(.A1(new_n664), .A2(new_n665), .ZN(new_n667));
  NOR3_X1   g242(.A1(new_n663), .A2(new_n666), .A3(new_n667), .ZN(new_n668));
  NAND2_X1  g243(.A1(new_n663), .A2(new_n666), .ZN(new_n669));
  XNOR2_X1  g244(.A(KEYINPUT84), .B(KEYINPUT20), .ZN(new_n670));
  XNOR2_X1  g245(.A(new_n669), .B(new_n670), .ZN(new_n671));
  AOI211_X1 g246(.A(new_n668), .B(new_n671), .C1(new_n663), .C2(new_n667), .ZN(new_n672));
  XOR2_X1   g247(.A(new_n672), .B(KEYINPUT85), .Z(new_n673));
  XNOR2_X1  g248(.A(new_n673), .B(KEYINPUT86), .ZN(new_n674));
  XOR2_X1   g249(.A(G1981), .B(G1986), .Z(new_n675));
  XNOR2_X1  g250(.A(G1991), .B(G1996), .ZN(new_n676));
  XNOR2_X1  g251(.A(new_n675), .B(new_n676), .ZN(new_n677));
  XOR2_X1   g252(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n678));
  XNOR2_X1  g253(.A(new_n677), .B(new_n678), .ZN(new_n679));
  XNOR2_X1  g254(.A(new_n674), .B(new_n679), .ZN(new_n680));
  INV_X1    g255(.A(new_n680), .ZN(G229));
  OAI221_X1 g256(.A(G2104), .B1(G95), .B2(G2105), .C1(new_n472), .C2(G107), .ZN(new_n682));
  XOR2_X1   g257(.A(new_n682), .B(KEYINPUT87), .Z(new_n683));
  AOI21_X1  g258(.A(new_n683), .B1(G131), .B2(new_n614), .ZN(new_n684));
  INV_X1    g259(.A(G119), .ZN(new_n685));
  OAI21_X1  g260(.A(new_n684), .B1(new_n685), .B2(new_n618), .ZN(new_n686));
  MUX2_X1   g261(.A(G25), .B(new_n686), .S(G29), .Z(new_n687));
  XOR2_X1   g262(.A(KEYINPUT35), .B(G1991), .Z(new_n688));
  INV_X1    g263(.A(new_n688), .ZN(new_n689));
  XNOR2_X1  g264(.A(new_n687), .B(new_n689), .ZN(new_n690));
  INV_X1    g265(.A(KEYINPUT88), .ZN(new_n691));
  NOR2_X1   g266(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  XOR2_X1   g267(.A(KEYINPUT89), .B(G16), .Z(new_n693));
  NOR2_X1   g268(.A1(new_n589), .A2(new_n693), .ZN(new_n694));
  AOI21_X1  g269(.A(new_n694), .B1(G24), .B2(new_n693), .ZN(new_n695));
  INV_X1    g270(.A(new_n695), .ZN(new_n696));
  AOI21_X1  g271(.A(KEYINPUT93), .B1(new_n696), .B2(G1986), .ZN(new_n697));
  OAI21_X1  g272(.A(new_n697), .B1(G1986), .B2(new_n696), .ZN(new_n698));
  NOR2_X1   g273(.A1(new_n692), .A2(new_n698), .ZN(new_n699));
  INV_X1    g274(.A(G16), .ZN(new_n700));
  NAND2_X1  g275(.A1(new_n700), .A2(G6), .ZN(new_n701));
  INV_X1    g276(.A(G305), .ZN(new_n702));
  OAI21_X1  g277(.A(new_n701), .B1(new_n702), .B2(new_n700), .ZN(new_n703));
  XOR2_X1   g278(.A(KEYINPUT32), .B(G1981), .Z(new_n704));
  XNOR2_X1  g279(.A(new_n703), .B(new_n704), .ZN(new_n705));
  NAND2_X1  g280(.A1(new_n693), .A2(G22), .ZN(new_n706));
  XOR2_X1   g281(.A(new_n706), .B(KEYINPUT92), .Z(new_n707));
  OAI21_X1  g282(.A(new_n707), .B1(G166), .B2(new_n693), .ZN(new_n708));
  XNOR2_X1  g283(.A(new_n708), .B(G1971), .ZN(new_n709));
  INV_X1    g284(.A(KEYINPUT91), .ZN(new_n710));
  NAND2_X1  g285(.A1(new_n700), .A2(G23), .ZN(new_n711));
  AND2_X1   g286(.A1(new_n574), .A2(new_n575), .ZN(new_n712));
  OAI21_X1  g287(.A(new_n711), .B1(new_n712), .B2(new_n700), .ZN(new_n713));
  XOR2_X1   g288(.A(KEYINPUT33), .B(G1976), .Z(new_n714));
  XNOR2_X1  g289(.A(new_n714), .B(KEYINPUT90), .ZN(new_n715));
  XNOR2_X1  g290(.A(new_n713), .B(new_n715), .ZN(new_n716));
  AOI21_X1  g291(.A(new_n709), .B1(new_n710), .B2(new_n716), .ZN(new_n717));
  OAI211_X1 g292(.A(new_n705), .B(new_n717), .C1(new_n710), .C2(new_n716), .ZN(new_n718));
  OR2_X1    g293(.A1(new_n718), .A2(KEYINPUT34), .ZN(new_n719));
  NAND2_X1  g294(.A1(new_n718), .A2(KEYINPUT34), .ZN(new_n720));
  NAND2_X1  g295(.A1(new_n690), .A2(new_n691), .ZN(new_n721));
  NAND4_X1  g296(.A1(new_n699), .A2(new_n719), .A3(new_n720), .A4(new_n721), .ZN(new_n722));
  INV_X1    g297(.A(KEYINPUT36), .ZN(new_n723));
  OR2_X1    g298(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  NAND2_X1  g299(.A1(new_n722), .A2(new_n723), .ZN(new_n725));
  XNOR2_X1  g300(.A(KEYINPUT31), .B(G11), .ZN(new_n726));
  XNOR2_X1  g301(.A(KEYINPUT30), .B(G28), .ZN(new_n727));
  INV_X1    g302(.A(G29), .ZN(new_n728));
  NAND2_X1  g303(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  OAI211_X1 g304(.A(new_n726), .B(new_n729), .C1(new_n620), .C2(new_n728), .ZN(new_n730));
  NAND2_X1  g305(.A1(new_n700), .A2(G21), .ZN(new_n731));
  OAI21_X1  g306(.A(new_n731), .B1(G168), .B2(new_n700), .ZN(new_n732));
  NOR2_X1   g307(.A1(G5), .A2(G16), .ZN(new_n733));
  XNOR2_X1  g308(.A(new_n733), .B(KEYINPUT99), .ZN(new_n734));
  OAI21_X1  g309(.A(new_n734), .B1(new_n548), .B2(new_n700), .ZN(new_n735));
  INV_X1    g310(.A(G1961), .ZN(new_n736));
  OAI22_X1  g311(.A1(new_n732), .A2(G1966), .B1(new_n735), .B2(new_n736), .ZN(new_n737));
  AOI211_X1 g312(.A(new_n730), .B(new_n737), .C1(G1966), .C2(new_n732), .ZN(new_n738));
  INV_X1    g313(.A(new_n738), .ZN(new_n739));
  OR2_X1    g314(.A1(new_n739), .A2(KEYINPUT100), .ZN(new_n740));
  NAND2_X1  g315(.A1(new_n739), .A2(KEYINPUT100), .ZN(new_n741));
  NAND2_X1  g316(.A1(new_n728), .A2(G33), .ZN(new_n742));
  NAND3_X1  g317(.A1(new_n472), .A2(G103), .A3(G2104), .ZN(new_n743));
  XOR2_X1   g318(.A(new_n743), .B(KEYINPUT25), .Z(new_n744));
  AOI22_X1  g319(.A1(new_n479), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n745));
  OR2_X1    g320(.A1(new_n745), .A2(new_n472), .ZN(new_n746));
  NAND2_X1  g321(.A1(new_n614), .A2(G139), .ZN(new_n747));
  NAND3_X1  g322(.A1(new_n744), .A2(new_n746), .A3(new_n747), .ZN(new_n748));
  INV_X1    g323(.A(new_n748), .ZN(new_n749));
  OAI21_X1  g324(.A(new_n742), .B1(new_n749), .B2(new_n728), .ZN(new_n750));
  OR2_X1    g325(.A1(new_n750), .A2(G2072), .ZN(new_n751));
  NAND2_X1  g326(.A1(new_n750), .A2(G2072), .ZN(new_n752));
  INV_X1    g327(.A(KEYINPUT24), .ZN(new_n753));
  INV_X1    g328(.A(G34), .ZN(new_n754));
  AOI21_X1  g329(.A(G29), .B1(new_n753), .B2(new_n754), .ZN(new_n755));
  OAI21_X1  g330(.A(new_n755), .B1(new_n753), .B2(new_n754), .ZN(new_n756));
  OAI21_X1  g331(.A(new_n756), .B1(G160), .B2(new_n728), .ZN(new_n757));
  INV_X1    g332(.A(G2084), .ZN(new_n758));
  XNOR2_X1  g333(.A(new_n757), .B(new_n758), .ZN(new_n759));
  NAND3_X1  g334(.A1(new_n751), .A2(new_n752), .A3(new_n759), .ZN(new_n760));
  NAND2_X1  g335(.A1(new_n700), .A2(G4), .ZN(new_n761));
  OAI21_X1  g336(.A(new_n761), .B1(new_n607), .B2(new_n700), .ZN(new_n762));
  INV_X1    g337(.A(G1348), .ZN(new_n763));
  XNOR2_X1  g338(.A(new_n762), .B(new_n763), .ZN(new_n764));
  NAND2_X1  g339(.A1(new_n735), .A2(new_n736), .ZN(new_n765));
  NAND2_X1  g340(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  NAND2_X1  g341(.A1(new_n728), .A2(G35), .ZN(new_n767));
  OAI21_X1  g342(.A(new_n767), .B1(G162), .B2(new_n728), .ZN(new_n768));
  XOR2_X1   g343(.A(new_n768), .B(KEYINPUT29), .Z(new_n769));
  INV_X1    g344(.A(new_n769), .ZN(new_n770));
  AOI211_X1 g345(.A(new_n760), .B(new_n766), .C1(G2090), .C2(new_n770), .ZN(new_n771));
  NAND2_X1  g346(.A1(new_n693), .A2(G19), .ZN(new_n772));
  XNOR2_X1  g347(.A(new_n772), .B(KEYINPUT94), .ZN(new_n773));
  OAI21_X1  g348(.A(new_n773), .B1(new_n555), .B2(new_n693), .ZN(new_n774));
  XOR2_X1   g349(.A(new_n774), .B(KEYINPUT95), .Z(new_n775));
  XNOR2_X1  g350(.A(new_n775), .B(G1341), .ZN(new_n776));
  NAND2_X1  g351(.A1(new_n728), .A2(G26), .ZN(new_n777));
  XOR2_X1   g352(.A(new_n777), .B(KEYINPUT28), .Z(new_n778));
  OAI221_X1 g353(.A(G2104), .B1(G104), .B2(G2105), .C1(new_n472), .C2(G116), .ZN(new_n779));
  INV_X1    g354(.A(G140), .ZN(new_n780));
  OAI21_X1  g355(.A(new_n779), .B1(new_n780), .B2(new_n480), .ZN(new_n781));
  AOI21_X1  g356(.A(new_n781), .B1(G128), .B2(new_n485), .ZN(new_n782));
  INV_X1    g357(.A(KEYINPUT96), .ZN(new_n783));
  NAND2_X1  g358(.A1(new_n782), .A2(new_n783), .ZN(new_n784));
  AND2_X1   g359(.A1(new_n485), .A2(G128), .ZN(new_n785));
  OAI21_X1  g360(.A(KEYINPUT96), .B1(new_n785), .B2(new_n781), .ZN(new_n786));
  NAND2_X1  g361(.A1(new_n784), .A2(new_n786), .ZN(new_n787));
  AOI21_X1  g362(.A(new_n778), .B1(new_n787), .B2(G29), .ZN(new_n788));
  INV_X1    g363(.A(G2067), .ZN(new_n789));
  XNOR2_X1  g364(.A(new_n788), .B(new_n789), .ZN(new_n790));
  NOR2_X1   g365(.A1(new_n776), .A2(new_n790), .ZN(new_n791));
  NAND4_X1  g366(.A1(new_n740), .A2(new_n741), .A3(new_n771), .A4(new_n791), .ZN(new_n792));
  NAND2_X1  g367(.A1(new_n728), .A2(G32), .ZN(new_n793));
  NAND3_X1  g368(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n794));
  INV_X1    g369(.A(KEYINPUT26), .ZN(new_n795));
  XNOR2_X1  g370(.A(new_n794), .B(new_n795), .ZN(new_n796));
  INV_X1    g371(.A(G105), .ZN(new_n797));
  INV_X1    g372(.A(G141), .ZN(new_n798));
  OAI221_X1 g373(.A(new_n796), .B1(new_n797), .B2(new_n468), .C1(new_n480), .C2(new_n798), .ZN(new_n799));
  AOI21_X1  g374(.A(new_n799), .B1(new_n485), .B2(G129), .ZN(new_n800));
  OR2_X1    g375(.A1(new_n800), .A2(KEYINPUT97), .ZN(new_n801));
  NAND2_X1  g376(.A1(new_n800), .A2(KEYINPUT97), .ZN(new_n802));
  NAND2_X1  g377(.A1(new_n801), .A2(new_n802), .ZN(new_n803));
  XNOR2_X1  g378(.A(new_n803), .B(KEYINPUT98), .ZN(new_n804));
  OAI21_X1  g379(.A(new_n793), .B1(new_n804), .B2(new_n728), .ZN(new_n805));
  INV_X1    g380(.A(new_n805), .ZN(new_n806));
  XNOR2_X1  g381(.A(KEYINPUT27), .B(G1996), .ZN(new_n807));
  AND2_X1   g382(.A1(new_n806), .A2(new_n807), .ZN(new_n808));
  NOR2_X1   g383(.A1(new_n806), .A2(new_n807), .ZN(new_n809));
  NAND2_X1  g384(.A1(new_n693), .A2(G20), .ZN(new_n810));
  XOR2_X1   g385(.A(new_n810), .B(KEYINPUT23), .Z(new_n811));
  AOI21_X1  g386(.A(new_n811), .B1(G299), .B2(G16), .ZN(new_n812));
  XNOR2_X1  g387(.A(KEYINPUT101), .B(G1956), .ZN(new_n813));
  XNOR2_X1  g388(.A(new_n812), .B(new_n813), .ZN(new_n814));
  NAND2_X1  g389(.A1(new_n728), .A2(G27), .ZN(new_n815));
  OAI21_X1  g390(.A(new_n815), .B1(G164), .B2(new_n728), .ZN(new_n816));
  INV_X1    g391(.A(G2078), .ZN(new_n817));
  XNOR2_X1  g392(.A(new_n816), .B(new_n817), .ZN(new_n818));
  OAI211_X1 g393(.A(new_n814), .B(new_n818), .C1(new_n770), .C2(G2090), .ZN(new_n819));
  NOR4_X1   g394(.A1(new_n792), .A2(new_n808), .A3(new_n809), .A4(new_n819), .ZN(new_n820));
  NAND3_X1  g395(.A1(new_n724), .A2(new_n725), .A3(new_n820), .ZN(G150));
  INV_X1    g396(.A(G150), .ZN(G311));
  NAND2_X1  g397(.A1(new_n607), .A2(G559), .ZN(new_n823));
  XNOR2_X1  g398(.A(new_n823), .B(KEYINPUT38), .ZN(new_n824));
  INV_X1    g399(.A(new_n555), .ZN(new_n825));
  NAND2_X1  g400(.A1(new_n516), .A2(G55), .ZN(new_n826));
  XNOR2_X1  g401(.A(KEYINPUT102), .B(G93), .ZN(new_n827));
  OAI21_X1  g402(.A(new_n826), .B1(new_n523), .B2(new_n827), .ZN(new_n828));
  AOI22_X1  g403(.A1(new_n526), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n829));
  NOR2_X1   g404(.A1(new_n829), .A2(new_n528), .ZN(new_n830));
  NOR2_X1   g405(.A1(new_n828), .A2(new_n830), .ZN(new_n831));
  INV_X1    g406(.A(new_n831), .ZN(new_n832));
  NAND2_X1  g407(.A1(new_n825), .A2(new_n832), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n555), .A2(new_n831), .ZN(new_n834));
  NAND2_X1  g409(.A1(new_n833), .A2(new_n834), .ZN(new_n835));
  INV_X1    g410(.A(new_n835), .ZN(new_n836));
  XNOR2_X1  g411(.A(new_n824), .B(new_n836), .ZN(new_n837));
  OR2_X1    g412(.A1(new_n837), .A2(KEYINPUT39), .ZN(new_n838));
  INV_X1    g413(.A(G860), .ZN(new_n839));
  NAND2_X1  g414(.A1(new_n837), .A2(KEYINPUT39), .ZN(new_n840));
  NAND3_X1  g415(.A1(new_n838), .A2(new_n839), .A3(new_n840), .ZN(new_n841));
  NOR2_X1   g416(.A1(new_n831), .A2(new_n839), .ZN(new_n842));
  XNOR2_X1  g417(.A(new_n842), .B(KEYINPUT37), .ZN(new_n843));
  NAND2_X1  g418(.A1(new_n841), .A2(new_n843), .ZN(new_n844));
  XNOR2_X1  g419(.A(new_n844), .B(KEYINPUT103), .ZN(G145));
  XNOR2_X1  g420(.A(G160), .B(KEYINPUT104), .ZN(new_n846));
  XNOR2_X1  g421(.A(new_n846), .B(G162), .ZN(new_n847));
  XOR2_X1   g422(.A(new_n847), .B(new_n620), .Z(new_n848));
  XNOR2_X1  g423(.A(new_n803), .B(new_n787), .ZN(new_n849));
  NAND2_X1  g424(.A1(new_n508), .A2(new_n503), .ZN(new_n850));
  NAND4_X1  g425(.A1(new_n850), .A2(new_n492), .A3(new_n494), .A4(new_n499), .ZN(new_n851));
  INV_X1    g426(.A(new_n851), .ZN(new_n852));
  OR2_X1    g427(.A1(new_n849), .A2(new_n852), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n849), .A2(new_n852), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n749), .A2(KEYINPUT105), .ZN(new_n855));
  NAND3_X1  g430(.A1(new_n853), .A2(new_n854), .A3(new_n855), .ZN(new_n856));
  INV_X1    g431(.A(KEYINPUT98), .ZN(new_n857));
  AOI21_X1  g432(.A(KEYINPUT105), .B1(new_n749), .B2(new_n857), .ZN(new_n858));
  NAND2_X1  g433(.A1(new_n856), .A2(new_n858), .ZN(new_n859));
  XNOR2_X1  g434(.A(new_n686), .B(new_n623), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n614), .A2(G142), .ZN(new_n861));
  OAI221_X1 g436(.A(G2104), .B1(G106), .B2(G2105), .C1(new_n472), .C2(G118), .ZN(new_n862));
  INV_X1    g437(.A(G130), .ZN(new_n863));
  OAI211_X1 g438(.A(new_n861), .B(new_n862), .C1(new_n618), .C2(new_n863), .ZN(new_n864));
  XOR2_X1   g439(.A(new_n860), .B(new_n864), .Z(new_n865));
  INV_X1    g440(.A(new_n858), .ZN(new_n866));
  NAND4_X1  g441(.A1(new_n853), .A2(new_n866), .A3(new_n854), .A4(new_n855), .ZN(new_n867));
  NAND3_X1  g442(.A1(new_n859), .A2(new_n865), .A3(new_n867), .ZN(new_n868));
  INV_X1    g443(.A(new_n868), .ZN(new_n869));
  AOI21_X1  g444(.A(new_n865), .B1(new_n859), .B2(new_n867), .ZN(new_n870));
  OAI21_X1  g445(.A(new_n848), .B1(new_n869), .B2(new_n870), .ZN(new_n871));
  INV_X1    g446(.A(G37), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n859), .A2(new_n867), .ZN(new_n873));
  INV_X1    g448(.A(new_n865), .ZN(new_n874));
  NAND2_X1  g449(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  INV_X1    g450(.A(new_n848), .ZN(new_n876));
  NAND3_X1  g451(.A1(new_n875), .A2(new_n876), .A3(new_n868), .ZN(new_n877));
  NAND3_X1  g452(.A1(new_n871), .A2(new_n872), .A3(new_n877), .ZN(new_n878));
  XNOR2_X1  g453(.A(new_n878), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g454(.A1(new_n832), .A2(new_n603), .ZN(new_n880));
  XNOR2_X1  g455(.A(G305), .B(new_n589), .ZN(new_n881));
  XNOR2_X1  g456(.A(G166), .B(new_n712), .ZN(new_n882));
  XOR2_X1   g457(.A(new_n881), .B(new_n882), .Z(new_n883));
  NOR2_X1   g458(.A1(new_n883), .A2(KEYINPUT108), .ZN(new_n884));
  XNOR2_X1  g459(.A(new_n884), .B(KEYINPUT42), .ZN(new_n885));
  NAND2_X1  g460(.A1(G299), .A2(new_n607), .ZN(new_n886));
  INV_X1    g461(.A(KEYINPUT106), .ZN(new_n887));
  XNOR2_X1  g462(.A(new_n886), .B(new_n887), .ZN(new_n888));
  OR3_X1    g463(.A1(G299), .A2(new_n607), .A3(KEYINPUT107), .ZN(new_n889));
  OAI21_X1  g464(.A(KEYINPUT107), .B1(G299), .B2(new_n607), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  NOR2_X1   g466(.A1(new_n888), .A2(new_n891), .ZN(new_n892));
  OAI21_X1  g467(.A(KEYINPUT41), .B1(new_n888), .B2(new_n891), .ZN(new_n893));
  XNOR2_X1  g468(.A(new_n886), .B(KEYINPUT106), .ZN(new_n894));
  INV_X1    g469(.A(KEYINPUT41), .ZN(new_n895));
  NAND4_X1  g470(.A1(new_n894), .A2(new_n895), .A3(new_n890), .A4(new_n889), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n893), .A2(new_n896), .ZN(new_n897));
  XOR2_X1   g472(.A(new_n835), .B(new_n610), .Z(new_n898));
  MUX2_X1   g473(.A(new_n892), .B(new_n897), .S(new_n898), .Z(new_n899));
  XNOR2_X1  g474(.A(new_n885), .B(new_n899), .ZN(new_n900));
  OAI21_X1  g475(.A(new_n880), .B1(new_n900), .B2(new_n603), .ZN(G295));
  OAI21_X1  g476(.A(new_n880), .B1(new_n900), .B2(new_n603), .ZN(G331));
  NAND2_X1  g477(.A1(new_n570), .A2(G168), .ZN(new_n903));
  NAND2_X1  g478(.A1(G286), .A2(new_n548), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n905), .A2(new_n836), .ZN(new_n906));
  NAND3_X1  g481(.A1(new_n903), .A2(new_n835), .A3(new_n904), .ZN(new_n907));
  NAND4_X1  g482(.A1(new_n893), .A2(new_n896), .A3(new_n906), .A4(new_n907), .ZN(new_n908));
  AND2_X1   g483(.A1(new_n906), .A2(new_n907), .ZN(new_n909));
  OAI21_X1  g484(.A(new_n908), .B1(new_n909), .B2(new_n892), .ZN(new_n910));
  INV_X1    g485(.A(new_n883), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  OAI211_X1 g487(.A(new_n908), .B(new_n883), .C1(new_n909), .C2(new_n892), .ZN(new_n913));
  NAND3_X1  g488(.A1(new_n912), .A2(new_n872), .A3(new_n913), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n914), .A2(KEYINPUT43), .ZN(new_n915));
  INV_X1    g490(.A(KEYINPUT43), .ZN(new_n916));
  NAND4_X1  g491(.A1(new_n912), .A2(new_n916), .A3(new_n872), .A4(new_n913), .ZN(new_n917));
  OR2_X1    g492(.A1(KEYINPUT109), .A2(KEYINPUT44), .ZN(new_n918));
  NAND3_X1  g493(.A1(new_n915), .A2(new_n917), .A3(new_n918), .ZN(new_n919));
  NAND2_X1  g494(.A1(KEYINPUT109), .A2(KEYINPUT44), .ZN(new_n920));
  XOR2_X1   g495(.A(new_n920), .B(KEYINPUT110), .Z(new_n921));
  XNOR2_X1  g496(.A(new_n919), .B(new_n921), .ZN(G397));
  INV_X1    g497(.A(G1384), .ZN(new_n923));
  AOI21_X1  g498(.A(KEYINPUT45), .B1(new_n851), .B2(new_n923), .ZN(new_n924));
  INV_X1    g499(.A(new_n924), .ZN(new_n925));
  NAND2_X1  g500(.A1(G160), .A2(G40), .ZN(new_n926));
  NOR2_X1   g501(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  NAND3_X1  g502(.A1(new_n803), .A2(G1996), .A3(new_n927), .ZN(new_n928));
  XOR2_X1   g503(.A(new_n928), .B(KEYINPUT111), .Z(new_n929));
  INV_X1    g504(.A(G1996), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n804), .A2(new_n930), .ZN(new_n931));
  XNOR2_X1  g506(.A(new_n787), .B(new_n789), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n931), .A2(new_n932), .ZN(new_n933));
  AOI21_X1  g508(.A(new_n929), .B1(new_n933), .B2(new_n927), .ZN(new_n934));
  INV_X1    g509(.A(KEYINPUT112), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  INV_X1    g511(.A(new_n927), .ZN(new_n937));
  AOI21_X1  g512(.A(new_n937), .B1(new_n931), .B2(new_n932), .ZN(new_n938));
  OAI21_X1  g513(.A(KEYINPUT112), .B1(new_n938), .B2(new_n929), .ZN(new_n939));
  XNOR2_X1  g514(.A(new_n686), .B(new_n688), .ZN(new_n940));
  INV_X1    g515(.A(KEYINPUT113), .ZN(new_n941));
  AOI21_X1  g516(.A(new_n937), .B1(new_n940), .B2(new_n941), .ZN(new_n942));
  OAI21_X1  g517(.A(new_n942), .B1(new_n941), .B2(new_n940), .ZN(new_n943));
  NOR2_X1   g518(.A1(G290), .A2(G1986), .ZN(new_n944));
  AND2_X1   g519(.A1(G290), .A2(G1986), .ZN(new_n945));
  OAI21_X1  g520(.A(new_n927), .B1(new_n944), .B2(new_n945), .ZN(new_n946));
  NAND4_X1  g521(.A1(new_n936), .A2(new_n939), .A3(new_n943), .A4(new_n946), .ZN(new_n947));
  XOR2_X1   g522(.A(new_n947), .B(KEYINPUT114), .Z(new_n948));
  INV_X1    g523(.A(KEYINPUT62), .ZN(new_n949));
  INV_X1    g524(.A(KEYINPUT119), .ZN(new_n950));
  INV_X1    g525(.A(G40), .ZN(new_n951));
  NOR3_X1   g526(.A1(new_n469), .A2(new_n475), .A3(new_n951), .ZN(new_n952));
  AND2_X1   g527(.A1(new_n492), .A2(new_n494), .ZN(new_n953));
  AOI21_X1  g528(.A(G1384), .B1(new_n953), .B2(new_n509), .ZN(new_n954));
  OAI211_X1 g529(.A(new_n950), .B(new_n952), .C1(new_n954), .C2(KEYINPUT45), .ZN(new_n955));
  OAI21_X1  g530(.A(KEYINPUT119), .B1(new_n924), .B2(new_n926), .ZN(new_n956));
  AOI21_X1  g531(.A(new_n510), .B1(new_n850), .B2(new_n499), .ZN(new_n957));
  AOI211_X1 g532(.A(KEYINPUT68), .B(new_n498), .C1(new_n508), .C2(new_n503), .ZN(new_n958));
  OAI21_X1  g533(.A(new_n953), .B1(new_n957), .B2(new_n958), .ZN(new_n959));
  NAND3_X1  g534(.A1(new_n959), .A2(KEYINPUT45), .A3(new_n923), .ZN(new_n960));
  NAND3_X1  g535(.A1(new_n955), .A2(new_n956), .A3(new_n960), .ZN(new_n961));
  INV_X1    g536(.A(G1966), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n961), .A2(new_n962), .ZN(new_n963));
  INV_X1    g538(.A(KEYINPUT120), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n963), .A2(new_n964), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n851), .A2(new_n923), .ZN(new_n966));
  OAI21_X1  g541(.A(new_n952), .B1(new_n966), .B2(KEYINPUT50), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n959), .A2(new_n923), .ZN(new_n968));
  AOI21_X1  g543(.A(new_n967), .B1(KEYINPUT50), .B2(new_n968), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n969), .A2(new_n758), .ZN(new_n970));
  NAND3_X1  g545(.A1(new_n961), .A2(KEYINPUT120), .A3(new_n962), .ZN(new_n971));
  NAND4_X1  g546(.A1(new_n965), .A2(G168), .A3(new_n970), .A4(new_n971), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n972), .A2(G8), .ZN(new_n973));
  INV_X1    g548(.A(KEYINPUT51), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n973), .A2(new_n974), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n971), .A2(new_n970), .ZN(new_n976));
  AOI21_X1  g551(.A(KEYINPUT120), .B1(new_n961), .B2(new_n962), .ZN(new_n977));
  OAI21_X1  g552(.A(G286), .B1(new_n976), .B2(new_n977), .ZN(new_n978));
  NAND4_X1  g553(.A1(new_n978), .A2(new_n972), .A3(KEYINPUT51), .A4(G8), .ZN(new_n979));
  INV_X1    g554(.A(KEYINPUT123), .ZN(new_n980));
  NAND3_X1  g555(.A1(new_n975), .A2(new_n979), .A3(new_n980), .ZN(new_n981));
  INV_X1    g556(.A(new_n981), .ZN(new_n982));
  AOI21_X1  g557(.A(new_n980), .B1(new_n975), .B2(new_n979), .ZN(new_n983));
  OAI21_X1  g558(.A(new_n949), .B1(new_n982), .B2(new_n983), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n975), .A2(new_n979), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n985), .A2(KEYINPUT123), .ZN(new_n986));
  NAND3_X1  g561(.A1(new_n986), .A2(new_n981), .A3(KEYINPUT62), .ZN(new_n987));
  INV_X1    g562(.A(G8), .ZN(new_n988));
  NOR2_X1   g563(.A1(G166), .A2(new_n988), .ZN(new_n989));
  XOR2_X1   g564(.A(KEYINPUT116), .B(KEYINPUT55), .Z(new_n990));
  NAND2_X1  g565(.A1(new_n989), .A2(new_n990), .ZN(new_n991));
  INV_X1    g566(.A(KEYINPUT55), .ZN(new_n992));
  OAI22_X1  g567(.A1(G166), .A2(new_n988), .B1(KEYINPUT116), .B2(new_n992), .ZN(new_n993));
  NAND2_X1  g568(.A1(new_n991), .A2(new_n993), .ZN(new_n994));
  INV_X1    g569(.A(KEYINPUT45), .ZN(new_n995));
  OAI211_X1 g570(.A(KEYINPUT45), .B(new_n923), .C1(new_n495), .C2(new_n505), .ZN(new_n996));
  INV_X1    g571(.A(KEYINPUT115), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n996), .A2(new_n997), .ZN(new_n998));
  NAND4_X1  g573(.A1(new_n851), .A2(KEYINPUT115), .A3(KEYINPUT45), .A4(new_n923), .ZN(new_n999));
  AOI22_X1  g574(.A1(new_n968), .A2(new_n995), .B1(new_n998), .B2(new_n999), .ZN(new_n1000));
  AOI21_X1  g575(.A(G1971), .B1(new_n1000), .B2(new_n952), .ZN(new_n1001));
  OAI21_X1  g576(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n1002));
  INV_X1    g577(.A(KEYINPUT50), .ZN(new_n1003));
  AOI21_X1  g578(.A(new_n926), .B1(new_n954), .B2(new_n1003), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n1002), .A2(new_n1004), .ZN(new_n1005));
  NOR2_X1   g580(.A1(new_n1005), .A2(G2090), .ZN(new_n1006));
  OAI211_X1 g581(.A(G8), .B(new_n994), .C1(new_n1001), .C2(new_n1006), .ZN(new_n1007));
  INV_X1    g582(.A(KEYINPUT118), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n712), .A2(G1976), .ZN(new_n1009));
  NAND3_X1  g584(.A1(new_n952), .A2(new_n851), .A3(new_n923), .ZN(new_n1010));
  NAND3_X1  g585(.A1(new_n1009), .A2(new_n1010), .A3(G8), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n1011), .A2(KEYINPUT52), .ZN(new_n1012));
  INV_X1    g587(.A(G1976), .ZN(new_n1013));
  AOI21_X1  g588(.A(KEYINPUT52), .B1(G288), .B2(new_n1013), .ZN(new_n1014));
  NAND4_X1  g589(.A1(new_n1010), .A2(new_n1009), .A3(new_n1014), .A4(G8), .ZN(new_n1015));
  NAND2_X1  g590(.A1(new_n1012), .A2(new_n1015), .ZN(new_n1016));
  INV_X1    g591(.A(G1981), .ZN(new_n1017));
  AOI21_X1  g592(.A(new_n1017), .B1(new_n581), .B2(KEYINPUT117), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n1018), .A2(new_n582), .ZN(new_n1019));
  OAI211_X1 g594(.A(new_n577), .B(new_n581), .C1(KEYINPUT117), .C2(new_n1017), .ZN(new_n1020));
  AND3_X1   g595(.A1(new_n1019), .A2(KEYINPUT49), .A3(new_n1020), .ZN(new_n1021));
  AOI21_X1  g596(.A(KEYINPUT49), .B1(new_n1019), .B2(new_n1020), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n1010), .A2(G8), .ZN(new_n1023));
  NOR3_X1   g598(.A1(new_n1021), .A2(new_n1022), .A3(new_n1023), .ZN(new_n1024));
  OAI21_X1  g599(.A(new_n1008), .B1(new_n1016), .B2(new_n1024), .ZN(new_n1025));
  INV_X1    g600(.A(new_n1022), .ZN(new_n1026));
  INV_X1    g601(.A(new_n1023), .ZN(new_n1027));
  NAND3_X1  g602(.A1(new_n1019), .A2(KEYINPUT49), .A3(new_n1020), .ZN(new_n1028));
  NAND3_X1  g603(.A1(new_n1026), .A2(new_n1027), .A3(new_n1028), .ZN(new_n1029));
  NAND4_X1  g604(.A1(new_n1029), .A2(KEYINPUT118), .A3(new_n1012), .A4(new_n1015), .ZN(new_n1030));
  NAND2_X1  g605(.A1(new_n1025), .A2(new_n1030), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n1007), .A2(new_n1031), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n998), .A2(new_n999), .ZN(new_n1033));
  OAI21_X1  g608(.A(new_n995), .B1(G164), .B2(G1384), .ZN(new_n1034));
  NAND3_X1  g609(.A1(new_n1033), .A2(new_n1034), .A3(new_n952), .ZN(new_n1035));
  INV_X1    g610(.A(G1971), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n1035), .A2(new_n1036), .ZN(new_n1037));
  NAND3_X1  g612(.A1(new_n959), .A2(new_n1003), .A3(new_n923), .ZN(new_n1038));
  INV_X1    g613(.A(G2090), .ZN(new_n1039));
  AOI21_X1  g614(.A(new_n926), .B1(new_n966), .B2(KEYINPUT50), .ZN(new_n1040));
  NAND3_X1  g615(.A1(new_n1038), .A2(new_n1039), .A3(new_n1040), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n1037), .A2(new_n1041), .ZN(new_n1042));
  AOI21_X1  g617(.A(new_n994), .B1(new_n1042), .B2(G8), .ZN(new_n1043));
  OAI21_X1  g618(.A(KEYINPUT125), .B1(new_n1032), .B2(new_n1043), .ZN(new_n1044));
  INV_X1    g619(.A(new_n1041), .ZN(new_n1045));
  AOI21_X1  g620(.A(new_n1045), .B1(new_n1036), .B2(new_n1035), .ZN(new_n1046));
  OAI211_X1 g621(.A(new_n991), .B(new_n993), .C1(new_n1046), .C2(new_n988), .ZN(new_n1047));
  INV_X1    g622(.A(KEYINPUT125), .ZN(new_n1048));
  NAND4_X1  g623(.A1(new_n1047), .A2(new_n1048), .A3(new_n1031), .A4(new_n1007), .ZN(new_n1049));
  AOI21_X1  g624(.A(G1961), .B1(new_n1002), .B2(new_n1004), .ZN(new_n1050));
  NAND4_X1  g625(.A1(new_n1033), .A2(new_n1034), .A3(new_n817), .A4(new_n952), .ZN(new_n1051));
  INV_X1    g626(.A(KEYINPUT53), .ZN(new_n1052));
  AOI21_X1  g627(.A(new_n1050), .B1(new_n1051), .B2(new_n1052), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n817), .A2(KEYINPUT53), .ZN(new_n1054));
  OR2_X1    g629(.A1(new_n961), .A2(new_n1054), .ZN(new_n1055));
  AOI21_X1  g630(.A(G301), .B1(new_n1053), .B2(new_n1055), .ZN(new_n1056));
  AND3_X1   g631(.A1(new_n1044), .A2(new_n1049), .A3(new_n1056), .ZN(new_n1057));
  NAND3_X1  g632(.A1(new_n984), .A2(new_n987), .A3(new_n1057), .ZN(new_n1058));
  NOR3_X1   g633(.A1(new_n1024), .A2(G1976), .A3(G288), .ZN(new_n1059));
  NOR2_X1   g634(.A1(new_n582), .A2(G1981), .ZN(new_n1060));
  OAI21_X1  g635(.A(new_n1027), .B1(new_n1059), .B2(new_n1060), .ZN(new_n1061));
  NAND3_X1  g636(.A1(new_n1029), .A2(new_n1012), .A3(new_n1015), .ZN(new_n1062));
  OAI21_X1  g637(.A(new_n1061), .B1(new_n1007), .B2(new_n1062), .ZN(new_n1063));
  INV_X1    g638(.A(KEYINPUT63), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n969), .A2(new_n1039), .ZN(new_n1065));
  AOI21_X1  g640(.A(new_n988), .B1(new_n1037), .B2(new_n1065), .ZN(new_n1066));
  AOI211_X1 g641(.A(new_n1064), .B(new_n1062), .C1(new_n1066), .C2(new_n994), .ZN(new_n1067));
  OAI21_X1  g642(.A(new_n1067), .B1(new_n994), .B2(new_n1066), .ZN(new_n1068));
  OAI211_X1 g643(.A(G8), .B(G168), .C1(new_n976), .C2(new_n977), .ZN(new_n1069));
  OR2_X1    g644(.A1(new_n1068), .A2(new_n1069), .ZN(new_n1070));
  NAND3_X1  g645(.A1(new_n1047), .A2(new_n1031), .A3(new_n1007), .ZN(new_n1071));
  OAI21_X1  g646(.A(new_n1064), .B1(new_n1071), .B2(new_n1069), .ZN(new_n1072));
  AOI21_X1  g647(.A(new_n1063), .B1(new_n1070), .B2(new_n1072), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n1058), .A2(new_n1073), .ZN(new_n1074));
  INV_X1    g649(.A(KEYINPUT57), .ZN(new_n1075));
  AOI21_X1  g650(.A(new_n1075), .B1(new_n566), .B2(new_n568), .ZN(new_n1076));
  INV_X1    g651(.A(KEYINPUT76), .ZN(new_n1077));
  XNOR2_X1  g652(.A(new_n567), .B(new_n1077), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n563), .A2(new_n565), .ZN(new_n1079));
  NOR3_X1   g654(.A1(new_n1078), .A2(new_n1079), .A3(KEYINPUT57), .ZN(new_n1080));
  NOR2_X1   g655(.A1(new_n1076), .A2(new_n1080), .ZN(new_n1081));
  XNOR2_X1  g656(.A(KEYINPUT56), .B(G2072), .ZN(new_n1082));
  NAND4_X1  g657(.A1(new_n1033), .A2(new_n1034), .A3(new_n952), .A4(new_n1082), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n1038), .A2(new_n1040), .ZN(new_n1084));
  INV_X1    g659(.A(G1956), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n1084), .A2(new_n1085), .ZN(new_n1086));
  AOI21_X1  g661(.A(new_n1081), .B1(new_n1083), .B2(new_n1086), .ZN(new_n1087));
  NAND3_X1  g662(.A1(new_n1083), .A2(new_n1086), .A3(new_n1081), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n1088), .A2(KEYINPUT61), .ZN(new_n1089));
  INV_X1    g664(.A(KEYINPUT59), .ZN(new_n1090));
  NOR2_X1   g665(.A1(new_n926), .A2(G1996), .ZN(new_n1091));
  NAND3_X1  g666(.A1(new_n1033), .A2(new_n1034), .A3(new_n1091), .ZN(new_n1092));
  XOR2_X1   g667(.A(KEYINPUT58), .B(G1341), .Z(new_n1093));
  NAND2_X1  g668(.A1(new_n1010), .A2(new_n1093), .ZN(new_n1094));
  NAND2_X1  g669(.A1(new_n1092), .A2(new_n1094), .ZN(new_n1095));
  AOI21_X1  g670(.A(new_n1090), .B1(new_n1095), .B2(new_n555), .ZN(new_n1096));
  AOI211_X1 g671(.A(KEYINPUT59), .B(new_n825), .C1(new_n1092), .C2(new_n1094), .ZN(new_n1097));
  OAI22_X1  g672(.A1(new_n1087), .A2(new_n1089), .B1(new_n1096), .B2(new_n1097), .ZN(new_n1098));
  INV_X1    g673(.A(new_n1087), .ZN(new_n1099));
  AOI21_X1  g674(.A(KEYINPUT61), .B1(new_n1099), .B2(new_n1088), .ZN(new_n1100));
  OAI21_X1  g675(.A(KEYINPUT121), .B1(new_n1098), .B2(new_n1100), .ZN(new_n1101));
  OR2_X1    g676(.A1(new_n1096), .A2(new_n1097), .ZN(new_n1102));
  INV_X1    g677(.A(KEYINPUT121), .ZN(new_n1103));
  INV_X1    g678(.A(KEYINPUT61), .ZN(new_n1104));
  INV_X1    g679(.A(new_n1088), .ZN(new_n1105));
  OAI21_X1  g680(.A(new_n1104), .B1(new_n1105), .B2(new_n1087), .ZN(new_n1106));
  NAND3_X1  g681(.A1(new_n1099), .A2(KEYINPUT61), .A3(new_n1088), .ZN(new_n1107));
  NAND4_X1  g682(.A1(new_n1102), .A2(new_n1103), .A3(new_n1106), .A4(new_n1107), .ZN(new_n1108));
  NAND2_X1  g683(.A1(new_n1005), .A2(new_n763), .ZN(new_n1109));
  INV_X1    g684(.A(new_n1010), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n1110), .A2(new_n789), .ZN(new_n1111));
  NAND2_X1  g686(.A1(new_n1109), .A2(new_n1111), .ZN(new_n1112));
  INV_X1    g687(.A(KEYINPUT60), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n1112), .A2(new_n1113), .ZN(new_n1114));
  NOR2_X1   g689(.A1(new_n1112), .A2(new_n1113), .ZN(new_n1115));
  NOR2_X1   g690(.A1(new_n1115), .A2(new_n599), .ZN(new_n1116));
  NOR3_X1   g691(.A1(new_n1112), .A2(new_n1113), .A3(new_n607), .ZN(new_n1117));
  OAI21_X1  g692(.A(new_n1114), .B1(new_n1116), .B2(new_n1117), .ZN(new_n1118));
  NAND3_X1  g693(.A1(new_n1101), .A2(new_n1108), .A3(new_n1118), .ZN(new_n1119));
  NAND2_X1  g694(.A1(new_n1112), .A2(new_n607), .ZN(new_n1120));
  AOI21_X1  g695(.A(new_n1105), .B1(new_n1099), .B2(new_n1120), .ZN(new_n1121));
  INV_X1    g696(.A(new_n1121), .ZN(new_n1122));
  AND3_X1   g697(.A1(new_n1119), .A2(KEYINPUT122), .A3(new_n1122), .ZN(new_n1123));
  AOI21_X1  g698(.A(KEYINPUT122), .B1(new_n1119), .B2(new_n1122), .ZN(new_n1124));
  INV_X1    g699(.A(KEYINPUT124), .ZN(new_n1125));
  OR2_X1    g700(.A1(new_n469), .A2(new_n1125), .ZN(new_n1126));
  NOR3_X1   g701(.A1(new_n475), .A2(new_n951), .A3(new_n1054), .ZN(new_n1127));
  NAND2_X1  g702(.A1(new_n469), .A2(new_n1125), .ZN(new_n1128));
  AND3_X1   g703(.A1(new_n1126), .A2(new_n1127), .A3(new_n1128), .ZN(new_n1129));
  NAND3_X1  g704(.A1(new_n1033), .A2(new_n925), .A3(new_n1129), .ZN(new_n1130));
  NAND2_X1  g705(.A1(new_n1053), .A2(new_n1130), .ZN(new_n1131));
  NAND2_X1  g706(.A1(new_n1131), .A2(G171), .ZN(new_n1132));
  NAND3_X1  g707(.A1(new_n1053), .A2(G301), .A3(new_n1055), .ZN(new_n1133));
  NAND3_X1  g708(.A1(new_n1132), .A2(KEYINPUT54), .A3(new_n1133), .ZN(new_n1134));
  INV_X1    g709(.A(KEYINPUT54), .ZN(new_n1135));
  NAND2_X1  g710(.A1(new_n1051), .A2(new_n1052), .ZN(new_n1136));
  INV_X1    g711(.A(new_n1050), .ZN(new_n1137));
  AND4_X1   g712(.A1(G301), .A2(new_n1136), .A3(new_n1137), .A4(new_n1130), .ZN(new_n1138));
  OAI21_X1  g713(.A(new_n1135), .B1(new_n1138), .B2(new_n1056), .ZN(new_n1139));
  AND4_X1   g714(.A1(new_n1044), .A2(new_n1049), .A3(new_n1134), .A4(new_n1139), .ZN(new_n1140));
  NAND3_X1  g715(.A1(new_n1140), .A2(new_n986), .A3(new_n981), .ZN(new_n1141));
  NOR3_X1   g716(.A1(new_n1123), .A2(new_n1124), .A3(new_n1141), .ZN(new_n1142));
  OAI21_X1  g717(.A(new_n948), .B1(new_n1074), .B2(new_n1142), .ZN(new_n1143));
  INV_X1    g718(.A(new_n803), .ZN(new_n1144));
  AOI21_X1  g719(.A(new_n937), .B1(new_n932), .B2(new_n1144), .ZN(new_n1145));
  NAND2_X1  g720(.A1(new_n927), .A2(new_n930), .ZN(new_n1146));
  XOR2_X1   g721(.A(new_n1146), .B(KEYINPUT46), .Z(new_n1147));
  NOR2_X1   g722(.A1(new_n1145), .A2(new_n1147), .ZN(new_n1148));
  XOR2_X1   g723(.A(new_n1148), .B(KEYINPUT47), .Z(new_n1149));
  AND2_X1   g724(.A1(new_n936), .A2(new_n939), .ZN(new_n1150));
  NAND2_X1  g725(.A1(new_n1150), .A2(new_n943), .ZN(new_n1151));
  NAND2_X1  g726(.A1(new_n927), .A2(new_n944), .ZN(new_n1152));
  XOR2_X1   g727(.A(new_n1152), .B(KEYINPUT126), .Z(new_n1153));
  XNOR2_X1  g728(.A(new_n1153), .B(KEYINPUT48), .ZN(new_n1154));
  OAI21_X1  g729(.A(new_n1149), .B1(new_n1151), .B2(new_n1154), .ZN(new_n1155));
  NOR2_X1   g730(.A1(new_n686), .A2(new_n689), .ZN(new_n1156));
  NAND2_X1  g731(.A1(new_n1150), .A2(new_n1156), .ZN(new_n1157));
  NAND3_X1  g732(.A1(new_n784), .A2(new_n786), .A3(new_n789), .ZN(new_n1158));
  AOI21_X1  g733(.A(new_n937), .B1(new_n1157), .B2(new_n1158), .ZN(new_n1159));
  NOR2_X1   g734(.A1(new_n1155), .A2(new_n1159), .ZN(new_n1160));
  NAND2_X1  g735(.A1(new_n1143), .A2(new_n1160), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g736(.A(G319), .ZN(new_n1163));
  OR3_X1    g737(.A1(G401), .A2(new_n1163), .A3(G227), .ZN(new_n1164));
  INV_X1    g738(.A(KEYINPUT127), .ZN(new_n1165));
  NAND2_X1  g739(.A1(new_n1164), .A2(new_n1165), .ZN(new_n1166));
  OR2_X1    g740(.A1(new_n1164), .A2(new_n1165), .ZN(new_n1167));
  NAND3_X1  g741(.A1(new_n680), .A2(new_n1166), .A3(new_n1167), .ZN(new_n1168));
  INV_X1    g742(.A(new_n1168), .ZN(new_n1169));
  NAND2_X1  g743(.A1(new_n915), .A2(new_n917), .ZN(new_n1170));
  NAND3_X1  g744(.A1(new_n1169), .A2(new_n878), .A3(new_n1170), .ZN(G225));
  INV_X1    g745(.A(G225), .ZN(G308));
endmodule


