//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 0 1 0 0 0 0 1 0 1 0 0 1 1 1 1 0 1 1 0 1 1 0 1 0 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 1 1 1 1 1 1 0 0 1 0 0 0 0 0 1 1 0 1 0 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:18:00 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n671, new_n672,
    new_n673, new_n674, new_n676, new_n677, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n715, new_n716, new_n717,
    new_n718, new_n720, new_n721, new_n722, new_n723, new_n724, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n732, new_n733, new_n734,
    new_n735, new_n737, new_n738, new_n739, new_n740, new_n741, new_n743,
    new_n744, new_n745, new_n746, new_n747, new_n748, new_n749, new_n750,
    new_n751, new_n753, new_n755, new_n756, new_n757, new_n758, new_n759,
    new_n760, new_n761, new_n762, new_n763, new_n764, new_n765, new_n766,
    new_n767, new_n768, new_n769, new_n770, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n782,
    new_n783, new_n784, new_n785, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n830, new_n831, new_n833, new_n834, new_n836,
    new_n837, new_n838, new_n839, new_n840, new_n841, new_n842, new_n843,
    new_n844, new_n845, new_n846, new_n847, new_n848, new_n849, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n898, new_n899, new_n900, new_n901, new_n902, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n921, new_n922, new_n923, new_n924, new_n925, new_n926, new_n927,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n949, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n963, new_n964, new_n965, new_n966,
    new_n967, new_n968, new_n969, new_n971, new_n972, new_n973, new_n974;
  INV_X1    g000(.A(KEYINPUT97), .ZN(new_n202));
  XNOR2_X1  g001(.A(G190gat), .B(G218gat), .ZN(new_n203));
  NAND2_X1  g002(.A1(G232gat), .A2(G233gat), .ZN(new_n204));
  INV_X1    g003(.A(KEYINPUT41), .ZN(new_n205));
  NOR2_X1   g004(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  INV_X1    g005(.A(G29gat), .ZN(new_n207));
  INV_X1    g006(.A(G36gat), .ZN(new_n208));
  NAND3_X1  g007(.A1(new_n207), .A2(new_n208), .A3(KEYINPUT14), .ZN(new_n209));
  INV_X1    g008(.A(KEYINPUT14), .ZN(new_n210));
  OAI21_X1  g009(.A(new_n210), .B1(G29gat), .B2(G36gat), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n209), .A2(new_n211), .ZN(new_n212));
  INV_X1    g011(.A(KEYINPUT85), .ZN(new_n213));
  XNOR2_X1  g012(.A(new_n212), .B(new_n213), .ZN(new_n214));
  XOR2_X1   g013(.A(G43gat), .B(G50gat), .Z(new_n215));
  INV_X1    g014(.A(KEYINPUT15), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  XNOR2_X1  g016(.A(G43gat), .B(G50gat), .ZN(new_n218));
  INV_X1    g017(.A(KEYINPUT87), .ZN(new_n219));
  NAND3_X1  g018(.A1(new_n218), .A2(new_n219), .A3(KEYINPUT15), .ZN(new_n220));
  INV_X1    g019(.A(new_n212), .ZN(new_n221));
  XNOR2_X1  g020(.A(KEYINPUT86), .B(G29gat), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n222), .A2(G36gat), .ZN(new_n223));
  NAND4_X1  g022(.A1(new_n217), .A2(new_n220), .A3(new_n221), .A4(new_n223), .ZN(new_n224));
  NAND3_X1  g023(.A1(new_n214), .A2(new_n224), .A3(new_n223), .ZN(new_n225));
  NOR2_X1   g024(.A1(new_n215), .A2(new_n216), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  INV_X1    g026(.A(KEYINPUT88), .ZN(new_n228));
  OR2_X1    g027(.A1(new_n224), .A2(KEYINPUT87), .ZN(new_n229));
  AND3_X1   g028(.A1(new_n227), .A2(new_n228), .A3(new_n229), .ZN(new_n230));
  AOI21_X1  g029(.A(new_n228), .B1(new_n227), .B2(new_n229), .ZN(new_n231));
  NOR2_X1   g030(.A1(new_n230), .A2(new_n231), .ZN(new_n232));
  INV_X1    g031(.A(KEYINPUT17), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n232), .A2(new_n233), .ZN(new_n234));
  AOI21_X1  g033(.A(new_n233), .B1(new_n227), .B2(new_n229), .ZN(new_n235));
  INV_X1    g034(.A(new_n235), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n234), .A2(new_n236), .ZN(new_n237));
  INV_X1    g036(.A(G85gat), .ZN(new_n238));
  INV_X1    g037(.A(G92gat), .ZN(new_n239));
  OAI21_X1  g038(.A(KEYINPUT7), .B1(new_n238), .B2(new_n239), .ZN(new_n240));
  INV_X1    g039(.A(KEYINPUT7), .ZN(new_n241));
  NAND3_X1  g040(.A1(new_n241), .A2(G85gat), .A3(G92gat), .ZN(new_n242));
  NAND2_X1  g041(.A1(G99gat), .A2(G106gat), .ZN(new_n243));
  AOI22_X1  g042(.A1(new_n240), .A2(new_n242), .B1(KEYINPUT8), .B2(new_n243), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n238), .A2(new_n239), .ZN(new_n245));
  NAND2_X1  g044(.A1(new_n244), .A2(new_n245), .ZN(new_n246));
  XOR2_X1   g045(.A(G99gat), .B(G106gat), .Z(new_n247));
  NAND2_X1  g046(.A1(new_n246), .A2(new_n247), .ZN(new_n248));
  INV_X1    g047(.A(new_n247), .ZN(new_n249));
  NAND3_X1  g048(.A1(new_n244), .A2(new_n249), .A3(new_n245), .ZN(new_n250));
  NAND3_X1  g049(.A1(new_n248), .A2(KEYINPUT95), .A3(new_n250), .ZN(new_n251));
  OR3_X1    g050(.A1(new_n246), .A2(KEYINPUT95), .A3(new_n247), .ZN(new_n252));
  AND3_X1   g051(.A1(new_n251), .A2(new_n252), .A3(KEYINPUT96), .ZN(new_n253));
  AOI21_X1  g052(.A(KEYINPUT96), .B1(new_n251), .B2(new_n252), .ZN(new_n254));
  NOR2_X1   g053(.A1(new_n253), .A2(new_n254), .ZN(new_n255));
  AOI21_X1  g054(.A(new_n206), .B1(new_n237), .B2(new_n255), .ZN(new_n256));
  OR2_X1    g055(.A1(new_n230), .A2(new_n231), .ZN(new_n257));
  INV_X1    g056(.A(new_n255), .ZN(new_n258));
  NAND2_X1  g057(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  AOI21_X1  g058(.A(new_n203), .B1(new_n256), .B2(new_n259), .ZN(new_n260));
  AOI21_X1  g059(.A(new_n258), .B1(new_n234), .B2(new_n236), .ZN(new_n261));
  NOR2_X1   g060(.A1(new_n232), .A2(new_n255), .ZN(new_n262));
  INV_X1    g061(.A(new_n203), .ZN(new_n263));
  NOR4_X1   g062(.A1(new_n261), .A2(new_n262), .A3(new_n206), .A4(new_n263), .ZN(new_n264));
  OAI21_X1  g063(.A(new_n202), .B1(new_n260), .B2(new_n264), .ZN(new_n265));
  NOR3_X1   g064(.A1(new_n230), .A2(new_n231), .A3(KEYINPUT17), .ZN(new_n266));
  NOR2_X1   g065(.A1(new_n266), .A2(new_n235), .ZN(new_n267));
  OAI221_X1 g066(.A(new_n259), .B1(new_n205), .B2(new_n204), .C1(new_n267), .C2(new_n258), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n268), .A2(new_n263), .ZN(new_n269));
  NAND3_X1  g068(.A1(new_n256), .A2(new_n259), .A3(new_n203), .ZN(new_n270));
  NAND3_X1  g069(.A1(new_n269), .A2(new_n270), .A3(KEYINPUT97), .ZN(new_n271));
  XNOR2_X1  g070(.A(KEYINPUT94), .B(G134gat), .ZN(new_n272));
  XNOR2_X1  g071(.A(new_n272), .B(G162gat), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n204), .A2(new_n205), .ZN(new_n274));
  XOR2_X1   g073(.A(new_n273), .B(new_n274), .Z(new_n275));
  INV_X1    g074(.A(new_n275), .ZN(new_n276));
  NAND3_X1  g075(.A1(new_n265), .A2(new_n271), .A3(new_n276), .ZN(new_n277));
  OAI211_X1 g076(.A(new_n202), .B(new_n275), .C1(new_n260), .C2(new_n264), .ZN(new_n278));
  AND2_X1   g077(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  XOR2_X1   g078(.A(G57gat), .B(G64gat), .Z(new_n280));
  NOR2_X1   g079(.A1(new_n280), .A2(KEYINPUT92), .ZN(new_n281));
  INV_X1    g080(.A(KEYINPUT9), .ZN(new_n282));
  XNOR2_X1  g081(.A(G57gat), .B(G64gat), .ZN(new_n283));
  INV_X1    g082(.A(KEYINPUT92), .ZN(new_n284));
  NOR2_X1   g083(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  OR3_X1    g084(.A1(new_n281), .A2(new_n282), .A3(new_n285), .ZN(new_n286));
  OR2_X1    g085(.A1(G71gat), .A2(G78gat), .ZN(new_n287));
  NAND2_X1  g086(.A1(G71gat), .A2(G78gat), .ZN(new_n288));
  AND2_X1   g087(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  OAI21_X1  g088(.A(new_n288), .B1(new_n287), .B2(new_n282), .ZN(new_n290));
  AOI22_X1  g089(.A1(new_n286), .A2(new_n289), .B1(new_n290), .B2(new_n280), .ZN(new_n291));
  NOR2_X1   g090(.A1(new_n291), .A2(KEYINPUT21), .ZN(new_n292));
  NAND2_X1  g091(.A1(G231gat), .A2(G233gat), .ZN(new_n293));
  XNOR2_X1  g092(.A(new_n292), .B(new_n293), .ZN(new_n294));
  XNOR2_X1  g093(.A(new_n294), .B(G211gat), .ZN(new_n295));
  XNOR2_X1  g094(.A(G15gat), .B(G22gat), .ZN(new_n296));
  INV_X1    g095(.A(KEYINPUT16), .ZN(new_n297));
  OAI21_X1  g096(.A(new_n296), .B1(new_n297), .B2(G1gat), .ZN(new_n298));
  OAI21_X1  g097(.A(new_n298), .B1(G1gat), .B2(new_n296), .ZN(new_n299));
  INV_X1    g098(.A(G8gat), .ZN(new_n300));
  XNOR2_X1  g099(.A(new_n299), .B(new_n300), .ZN(new_n301));
  INV_X1    g100(.A(new_n301), .ZN(new_n302));
  AOI21_X1  g101(.A(new_n302), .B1(KEYINPUT21), .B2(new_n291), .ZN(new_n303));
  XNOR2_X1  g102(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n304));
  XNOR2_X1  g103(.A(new_n303), .B(new_n304), .ZN(new_n305));
  XNOR2_X1  g104(.A(new_n295), .B(new_n305), .ZN(new_n306));
  XNOR2_X1  g105(.A(KEYINPUT93), .B(G183gat), .ZN(new_n307));
  XNOR2_X1  g106(.A(G127gat), .B(G155gat), .ZN(new_n308));
  XNOR2_X1  g107(.A(new_n307), .B(new_n308), .ZN(new_n309));
  XNOR2_X1  g108(.A(new_n306), .B(new_n309), .ZN(new_n310));
  NOR2_X1   g109(.A1(new_n279), .A2(new_n310), .ZN(new_n311));
  NAND2_X1  g110(.A1(G230gat), .A2(G233gat), .ZN(new_n312));
  INV_X1    g111(.A(new_n312), .ZN(new_n313));
  OAI211_X1 g112(.A(KEYINPUT10), .B(new_n291), .C1(new_n253), .C2(new_n254), .ZN(new_n314));
  AOI21_X1  g113(.A(new_n249), .B1(new_n244), .B2(new_n245), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n315), .A2(KEYINPUT98), .ZN(new_n316));
  INV_X1    g115(.A(KEYINPUT98), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n250), .A2(new_n317), .ZN(new_n318));
  OAI21_X1  g117(.A(new_n316), .B1(new_n318), .B2(new_n315), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n291), .A2(new_n319), .ZN(new_n320));
  INV_X1    g119(.A(KEYINPUT10), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n290), .A2(new_n280), .ZN(new_n322));
  NOR3_X1   g121(.A1(new_n281), .A2(new_n282), .A3(new_n285), .ZN(new_n323));
  INV_X1    g122(.A(new_n289), .ZN(new_n324));
  OAI21_X1  g123(.A(new_n322), .B1(new_n323), .B2(new_n324), .ZN(new_n325));
  NAND3_X1  g124(.A1(new_n325), .A2(new_n252), .A3(new_n251), .ZN(new_n326));
  NAND3_X1  g125(.A1(new_n320), .A2(new_n321), .A3(new_n326), .ZN(new_n327));
  AOI21_X1  g126(.A(new_n313), .B1(new_n314), .B2(new_n327), .ZN(new_n328));
  XNOR2_X1  g127(.A(new_n328), .B(KEYINPUT99), .ZN(new_n329));
  INV_X1    g128(.A(KEYINPUT101), .ZN(new_n330));
  XNOR2_X1  g129(.A(G120gat), .B(G148gat), .ZN(new_n331));
  INV_X1    g130(.A(G204gat), .ZN(new_n332));
  XNOR2_X1  g131(.A(new_n331), .B(new_n332), .ZN(new_n333));
  XNOR2_X1  g132(.A(KEYINPUT100), .B(G176gat), .ZN(new_n334));
  XOR2_X1   g133(.A(new_n333), .B(new_n334), .Z(new_n335));
  INV_X1    g134(.A(new_n335), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n320), .A2(new_n326), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n337), .A2(new_n313), .ZN(new_n338));
  NAND4_X1  g137(.A1(new_n329), .A2(new_n330), .A3(new_n336), .A4(new_n338), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n314), .A2(new_n327), .ZN(new_n340));
  AOI21_X1  g139(.A(KEYINPUT99), .B1(new_n340), .B2(new_n312), .ZN(new_n341));
  INV_X1    g140(.A(KEYINPUT99), .ZN(new_n342));
  AOI211_X1 g141(.A(new_n342), .B(new_n313), .C1(new_n314), .C2(new_n327), .ZN(new_n343));
  OAI211_X1 g142(.A(new_n336), .B(new_n338), .C1(new_n341), .C2(new_n343), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n344), .A2(KEYINPUT101), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n339), .A2(new_n345), .ZN(new_n346));
  INV_X1    g145(.A(new_n338), .ZN(new_n347));
  OAI21_X1  g146(.A(new_n335), .B1(new_n328), .B2(new_n347), .ZN(new_n348));
  AOI21_X1  g147(.A(KEYINPUT102), .B1(new_n346), .B2(new_n348), .ZN(new_n349));
  INV_X1    g148(.A(KEYINPUT102), .ZN(new_n350));
  INV_X1    g149(.A(new_n348), .ZN(new_n351));
  AOI211_X1 g150(.A(new_n350), .B(new_n351), .C1(new_n339), .C2(new_n345), .ZN(new_n352));
  NOR2_X1   g151(.A1(new_n349), .A2(new_n352), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n311), .A2(new_n353), .ZN(new_n354));
  XNOR2_X1  g153(.A(new_n354), .B(KEYINPUT103), .ZN(new_n355));
  INV_X1    g154(.A(G120gat), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n356), .A2(G113gat), .ZN(new_n357));
  INV_X1    g156(.A(G113gat), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n358), .A2(G120gat), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n357), .A2(new_n359), .ZN(new_n360));
  XNOR2_X1  g159(.A(G127gat), .B(G134gat), .ZN(new_n361));
  INV_X1    g160(.A(KEYINPUT1), .ZN(new_n362));
  AND3_X1   g161(.A1(new_n360), .A2(new_n361), .A3(new_n362), .ZN(new_n363));
  INV_X1    g162(.A(G134gat), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n364), .A2(G127gat), .ZN(new_n365));
  INV_X1    g164(.A(G127gat), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n366), .A2(G134gat), .ZN(new_n367));
  AOI22_X1  g166(.A1(new_n360), .A2(new_n362), .B1(new_n365), .B2(new_n367), .ZN(new_n368));
  NOR2_X1   g167(.A1(new_n363), .A2(new_n368), .ZN(new_n369));
  INV_X1    g168(.A(new_n369), .ZN(new_n370));
  OAI21_X1  g169(.A(KEYINPUT76), .B1(G155gat), .B2(G162gat), .ZN(new_n371));
  XNOR2_X1  g170(.A(G141gat), .B(G148gat), .ZN(new_n372));
  INV_X1    g171(.A(KEYINPUT2), .ZN(new_n373));
  AOI21_X1  g172(.A(new_n373), .B1(G155gat), .B2(G162gat), .ZN(new_n374));
  OAI21_X1  g173(.A(new_n371), .B1(new_n372), .B2(new_n374), .ZN(new_n375));
  XNOR2_X1  g174(.A(G155gat), .B(G162gat), .ZN(new_n376));
  INV_X1    g175(.A(new_n376), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n375), .A2(new_n377), .ZN(new_n378));
  OAI211_X1 g177(.A(new_n376), .B(new_n371), .C1(new_n372), .C2(new_n374), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n378), .A2(new_n379), .ZN(new_n380));
  XNOR2_X1  g179(.A(new_n370), .B(new_n380), .ZN(new_n381));
  NAND2_X1  g180(.A1(G225gat), .A2(G233gat), .ZN(new_n382));
  INV_X1    g181(.A(new_n382), .ZN(new_n383));
  NAND3_X1  g182(.A1(new_n381), .A2(KEYINPUT5), .A3(new_n383), .ZN(new_n384));
  INV_X1    g183(.A(new_n384), .ZN(new_n385));
  INV_X1    g184(.A(KEYINPUT77), .ZN(new_n386));
  INV_X1    g185(.A(KEYINPUT67), .ZN(new_n387));
  OAI21_X1  g186(.A(new_n387), .B1(new_n363), .B2(new_n368), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n365), .A2(new_n367), .ZN(new_n389));
  XNOR2_X1  g188(.A(G113gat), .B(G120gat), .ZN(new_n390));
  OAI21_X1  g189(.A(new_n389), .B1(new_n390), .B2(KEYINPUT1), .ZN(new_n391));
  NAND3_X1  g190(.A1(new_n360), .A2(new_n361), .A3(new_n362), .ZN(new_n392));
  NAND3_X1  g191(.A1(new_n391), .A2(new_n392), .A3(KEYINPUT67), .ZN(new_n393));
  AOI22_X1  g192(.A1(new_n388), .A2(new_n393), .B1(new_n378), .B2(new_n379), .ZN(new_n394));
  INV_X1    g193(.A(KEYINPUT4), .ZN(new_n395));
  OAI21_X1  g194(.A(new_n386), .B1(new_n394), .B2(new_n395), .ZN(new_n396));
  NAND3_X1  g195(.A1(new_n380), .A2(new_n395), .A3(new_n369), .ZN(new_n397));
  AND3_X1   g196(.A1(new_n391), .A2(new_n392), .A3(KEYINPUT67), .ZN(new_n398));
  AOI21_X1  g197(.A(KEYINPUT67), .B1(new_n391), .B2(new_n392), .ZN(new_n399));
  NOR2_X1   g198(.A1(new_n398), .A2(new_n399), .ZN(new_n400));
  INV_X1    g199(.A(new_n380), .ZN(new_n401));
  OAI211_X1 g200(.A(KEYINPUT77), .B(KEYINPUT4), .C1(new_n400), .C2(new_n401), .ZN(new_n402));
  NAND3_X1  g201(.A1(new_n396), .A2(new_n397), .A3(new_n402), .ZN(new_n403));
  INV_X1    g202(.A(KEYINPUT3), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n380), .A2(new_n404), .ZN(new_n405));
  NAND3_X1  g204(.A1(new_n378), .A2(KEYINPUT3), .A3(new_n379), .ZN(new_n406));
  NAND3_X1  g205(.A1(new_n405), .A2(new_n370), .A3(new_n406), .ZN(new_n407));
  NAND3_X1  g206(.A1(new_n403), .A2(KEYINPUT5), .A3(new_n407), .ZN(new_n408));
  NAND3_X1  g207(.A1(new_n380), .A2(KEYINPUT4), .A3(new_n369), .ZN(new_n409));
  OAI211_X1 g208(.A(new_n407), .B(new_n409), .C1(KEYINPUT4), .C2(new_n394), .ZN(new_n410));
  INV_X1    g209(.A(KEYINPUT5), .ZN(new_n411));
  AOI21_X1  g210(.A(new_n383), .B1(new_n410), .B2(new_n411), .ZN(new_n412));
  AOI21_X1  g211(.A(new_n385), .B1(new_n408), .B2(new_n412), .ZN(new_n413));
  XNOR2_X1  g212(.A(G1gat), .B(G29gat), .ZN(new_n414));
  XNOR2_X1  g213(.A(new_n414), .B(KEYINPUT79), .ZN(new_n415));
  XOR2_X1   g214(.A(G57gat), .B(G85gat), .Z(new_n416));
  XNOR2_X1  g215(.A(new_n415), .B(new_n416), .ZN(new_n417));
  XNOR2_X1  g216(.A(KEYINPUT78), .B(KEYINPUT0), .ZN(new_n418));
  XNOR2_X1  g217(.A(new_n417), .B(new_n418), .ZN(new_n419));
  AOI21_X1  g218(.A(KEYINPUT6), .B1(new_n413), .B2(new_n419), .ZN(new_n420));
  NOR2_X1   g219(.A1(new_n413), .A2(new_n419), .ZN(new_n421));
  XNOR2_X1  g220(.A(new_n420), .B(new_n421), .ZN(new_n422));
  INV_X1    g221(.A(KEYINPUT83), .ZN(new_n423));
  XNOR2_X1  g222(.A(KEYINPUT69), .B(G204gat), .ZN(new_n424));
  INV_X1    g223(.A(G197gat), .ZN(new_n425));
  AND2_X1   g224(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  NOR2_X1   g225(.A1(new_n424), .A2(new_n425), .ZN(new_n427));
  INV_X1    g226(.A(G211gat), .ZN(new_n428));
  INV_X1    g227(.A(G218gat), .ZN(new_n429));
  NOR2_X1   g228(.A1(new_n428), .A2(new_n429), .ZN(new_n430));
  OAI22_X1  g229(.A1(new_n426), .A2(new_n427), .B1(KEYINPUT22), .B2(new_n430), .ZN(new_n431));
  XOR2_X1   g230(.A(G211gat), .B(G218gat), .Z(new_n432));
  XOR2_X1   g231(.A(new_n431), .B(new_n432), .Z(new_n433));
  INV_X1    g232(.A(KEYINPUT70), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n433), .A2(new_n434), .ZN(new_n435));
  NAND3_X1  g234(.A1(new_n431), .A2(KEYINPUT70), .A3(new_n432), .ZN(new_n436));
  AND2_X1   g235(.A1(new_n435), .A2(new_n436), .ZN(new_n437));
  AND2_X1   g236(.A1(G183gat), .A2(G190gat), .ZN(new_n438));
  OAI21_X1  g237(.A(KEYINPUT24), .B1(new_n438), .B2(KEYINPUT64), .ZN(new_n439));
  OR2_X1    g238(.A1(G183gat), .A2(G190gat), .ZN(new_n440));
  AOI21_X1  g239(.A(KEYINPUT64), .B1(G183gat), .B2(G190gat), .ZN(new_n441));
  INV_X1    g240(.A(KEYINPUT24), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n441), .A2(new_n442), .ZN(new_n443));
  NAND3_X1  g242(.A1(new_n439), .A2(new_n440), .A3(new_n443), .ZN(new_n444));
  INV_X1    g243(.A(G169gat), .ZN(new_n445));
  INV_X1    g244(.A(G176gat), .ZN(new_n446));
  NAND3_X1  g245(.A1(new_n445), .A2(new_n446), .A3(KEYINPUT23), .ZN(new_n447));
  INV_X1    g246(.A(KEYINPUT23), .ZN(new_n448));
  OAI21_X1  g247(.A(new_n448), .B1(G169gat), .B2(G176gat), .ZN(new_n449));
  NAND2_X1  g248(.A1(G169gat), .A2(G176gat), .ZN(new_n450));
  AND3_X1   g249(.A1(new_n447), .A2(new_n449), .A3(new_n450), .ZN(new_n451));
  NAND3_X1  g250(.A1(new_n444), .A2(KEYINPUT25), .A3(new_n451), .ZN(new_n452));
  INV_X1    g251(.A(KEYINPUT25), .ZN(new_n453));
  NAND2_X1  g252(.A1(G183gat), .A2(G190gat), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n454), .A2(new_n442), .ZN(new_n455));
  NAND3_X1  g254(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n456));
  AND3_X1   g255(.A1(new_n455), .A2(new_n456), .A3(new_n440), .ZN(new_n457));
  NAND3_X1  g256(.A1(new_n447), .A2(new_n449), .A3(new_n450), .ZN(new_n458));
  OAI21_X1  g257(.A(new_n453), .B1(new_n457), .B2(new_n458), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n452), .A2(new_n459), .ZN(new_n460));
  INV_X1    g259(.A(KEYINPUT27), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n461), .A2(G183gat), .ZN(new_n462));
  AOI21_X1  g261(.A(KEYINPUT28), .B1(new_n462), .B2(KEYINPUT66), .ZN(new_n463));
  INV_X1    g262(.A(G190gat), .ZN(new_n464));
  XNOR2_X1  g263(.A(KEYINPUT27), .B(G183gat), .ZN(new_n465));
  OAI211_X1 g264(.A(new_n463), .B(new_n464), .C1(KEYINPUT66), .C2(new_n465), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n465), .A2(new_n464), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n467), .A2(KEYINPUT28), .ZN(new_n468));
  OR3_X1    g267(.A1(KEYINPUT26), .A2(G169gat), .A3(G176gat), .ZN(new_n469));
  OAI21_X1  g268(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n470));
  NAND3_X1  g269(.A1(new_n469), .A2(new_n450), .A3(new_n470), .ZN(new_n471));
  NAND4_X1  g270(.A1(new_n466), .A2(new_n468), .A3(new_n454), .A4(new_n471), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n460), .A2(new_n472), .ZN(new_n473));
  INV_X1    g272(.A(KEYINPUT72), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  NAND3_X1  g274(.A1(new_n460), .A2(new_n472), .A3(KEYINPUT72), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  NAND2_X1  g276(.A1(G226gat), .A2(G233gat), .ZN(new_n478));
  INV_X1    g277(.A(KEYINPUT29), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  NAND4_X1  g279(.A1(new_n447), .A2(new_n449), .A3(KEYINPUT25), .A4(new_n450), .ZN(new_n481));
  XNOR2_X1  g280(.A(new_n441), .B(KEYINPUT24), .ZN(new_n482));
  AOI21_X1  g281(.A(new_n481), .B1(new_n482), .B2(new_n440), .ZN(new_n483));
  NAND3_X1  g282(.A1(new_n455), .A2(new_n440), .A3(new_n456), .ZN(new_n484));
  AOI21_X1  g283(.A(KEYINPUT25), .B1(new_n451), .B2(new_n484), .ZN(new_n485));
  OAI21_X1  g284(.A(KEYINPUT65), .B1(new_n483), .B2(new_n485), .ZN(new_n486));
  INV_X1    g285(.A(KEYINPUT65), .ZN(new_n487));
  NAND3_X1  g286(.A1(new_n452), .A2(new_n459), .A3(new_n487), .ZN(new_n488));
  NAND2_X1  g287(.A1(new_n486), .A2(new_n488), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n489), .A2(new_n472), .ZN(new_n490));
  OAI22_X1  g289(.A1(new_n477), .A2(new_n480), .B1(new_n490), .B2(new_n478), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n437), .A2(new_n491), .ZN(new_n492));
  XNOR2_X1  g291(.A(G8gat), .B(G36gat), .ZN(new_n493));
  XNOR2_X1  g292(.A(G64gat), .B(G92gat), .ZN(new_n494));
  XNOR2_X1  g293(.A(new_n493), .B(new_n494), .ZN(new_n495));
  INV_X1    g294(.A(new_n495), .ZN(new_n496));
  INV_X1    g295(.A(KEYINPUT71), .ZN(new_n497));
  AOI21_X1  g296(.A(KEYINPUT29), .B1(new_n489), .B2(new_n472), .ZN(new_n498));
  INV_X1    g297(.A(new_n478), .ZN(new_n499));
  OAI21_X1  g298(.A(new_n497), .B1(new_n498), .B2(new_n499), .ZN(new_n500));
  AND4_X1   g299(.A1(new_n468), .A2(new_n466), .A3(new_n454), .A4(new_n471), .ZN(new_n501));
  AOI21_X1  g300(.A(new_n501), .B1(new_n486), .B2(new_n488), .ZN(new_n502));
  OAI211_X1 g301(.A(KEYINPUT71), .B(new_n478), .C1(new_n502), .C2(KEYINPUT29), .ZN(new_n503));
  NAND3_X1  g302(.A1(new_n475), .A2(new_n499), .A3(new_n476), .ZN(new_n504));
  INV_X1    g303(.A(KEYINPUT73), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  NAND4_X1  g305(.A1(new_n475), .A2(KEYINPUT73), .A3(new_n499), .A4(new_n476), .ZN(new_n507));
  AOI22_X1  g306(.A1(new_n500), .A2(new_n503), .B1(new_n506), .B2(new_n507), .ZN(new_n508));
  OAI211_X1 g307(.A(new_n492), .B(new_n496), .C1(new_n508), .C2(new_n437), .ZN(new_n509));
  INV_X1    g308(.A(KEYINPUT37), .ZN(new_n510));
  OAI211_X1 g309(.A(new_n510), .B(new_n492), .C1(new_n508), .C2(new_n437), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n435), .A2(new_n436), .ZN(new_n512));
  NAND2_X1  g311(.A1(new_n491), .A2(new_n512), .ZN(new_n513));
  OAI211_X1 g312(.A(KEYINPUT37), .B(new_n513), .C1(new_n508), .C2(new_n512), .ZN(new_n514));
  XNOR2_X1  g313(.A(KEYINPUT82), .B(KEYINPUT38), .ZN(new_n515));
  INV_X1    g314(.A(new_n515), .ZN(new_n516));
  NAND4_X1  g315(.A1(new_n511), .A2(new_n514), .A3(new_n495), .A4(new_n516), .ZN(new_n517));
  NAND4_X1  g316(.A1(new_n422), .A2(new_n423), .A3(new_n509), .A4(new_n517), .ZN(new_n518));
  NAND2_X1  g317(.A1(new_n408), .A2(new_n412), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n519), .A2(new_n384), .ZN(new_n520));
  INV_X1    g319(.A(new_n419), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n522), .A2(new_n420), .ZN(new_n523));
  NAND3_X1  g322(.A1(new_n520), .A2(KEYINPUT6), .A3(new_n521), .ZN(new_n524));
  NAND3_X1  g323(.A1(new_n523), .A2(new_n524), .A3(new_n509), .ZN(new_n525));
  AND4_X1   g324(.A1(new_n495), .A2(new_n511), .A3(new_n514), .A4(new_n516), .ZN(new_n526));
  OAI21_X1  g325(.A(KEYINPUT83), .B1(new_n525), .B2(new_n526), .ZN(new_n527));
  NOR2_X1   g326(.A1(new_n508), .A2(new_n437), .ZN(new_n528));
  INV_X1    g327(.A(new_n528), .ZN(new_n529));
  AOI21_X1  g328(.A(new_n510), .B1(new_n529), .B2(new_n492), .ZN(new_n530));
  NAND2_X1  g329(.A1(new_n511), .A2(new_n495), .ZN(new_n531));
  OAI21_X1  g330(.A(new_n515), .B1(new_n530), .B2(new_n531), .ZN(new_n532));
  NAND3_X1  g331(.A1(new_n518), .A2(new_n527), .A3(new_n532), .ZN(new_n533));
  INV_X1    g332(.A(new_n405), .ZN(new_n534));
  OAI21_X1  g333(.A(new_n512), .B1(KEYINPUT29), .B2(new_n534), .ZN(new_n535));
  NAND2_X1  g334(.A1(G228gat), .A2(G233gat), .ZN(new_n536));
  OAI21_X1  g335(.A(new_n404), .B1(new_n433), .B2(KEYINPUT29), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n537), .A2(new_n401), .ZN(new_n538));
  NAND3_X1  g337(.A1(new_n535), .A2(new_n536), .A3(new_n538), .ZN(new_n539));
  INV_X1    g338(.A(new_n535), .ZN(new_n540));
  NAND3_X1  g339(.A1(new_n435), .A2(new_n479), .A3(new_n436), .ZN(new_n541));
  AOI21_X1  g340(.A(new_n380), .B1(new_n541), .B2(new_n404), .ZN(new_n542));
  NOR2_X1   g341(.A1(new_n540), .A2(new_n542), .ZN(new_n543));
  OAI21_X1  g342(.A(new_n539), .B1(new_n543), .B2(new_n536), .ZN(new_n544));
  XOR2_X1   g343(.A(KEYINPUT31), .B(G50gat), .Z(new_n545));
  XNOR2_X1  g344(.A(new_n545), .B(KEYINPUT80), .ZN(new_n546));
  XOR2_X1   g345(.A(G78gat), .B(G106gat), .Z(new_n547));
  XNOR2_X1  g346(.A(new_n547), .B(G22gat), .ZN(new_n548));
  XNOR2_X1  g347(.A(new_n546), .B(new_n548), .ZN(new_n549));
  INV_X1    g348(.A(new_n549), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n544), .A2(new_n550), .ZN(new_n551));
  OAI211_X1 g350(.A(new_n539), .B(new_n549), .C1(new_n543), .C2(new_n536), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  INV_X1    g352(.A(KEYINPUT39), .ZN(new_n554));
  INV_X1    g353(.A(KEYINPUT81), .ZN(new_n555));
  NAND3_X1  g354(.A1(new_n410), .A2(new_n555), .A3(new_n383), .ZN(new_n556));
  INV_X1    g355(.A(new_n556), .ZN(new_n557));
  AOI21_X1  g356(.A(new_n555), .B1(new_n410), .B2(new_n383), .ZN(new_n558));
  OAI21_X1  g357(.A(new_n554), .B1(new_n557), .B2(new_n558), .ZN(new_n559));
  INV_X1    g358(.A(new_n558), .ZN(new_n560));
  AOI21_X1  g359(.A(new_n554), .B1(new_n381), .B2(new_n382), .ZN(new_n561));
  NAND3_X1  g360(.A1(new_n560), .A2(new_n556), .A3(new_n561), .ZN(new_n562));
  NAND3_X1  g361(.A1(new_n559), .A2(new_n562), .A3(new_n419), .ZN(new_n563));
  INV_X1    g362(.A(KEYINPUT40), .ZN(new_n564));
  OAI21_X1  g363(.A(new_n522), .B1(new_n563), .B2(new_n564), .ZN(new_n565));
  AOI21_X1  g364(.A(new_n565), .B1(new_n564), .B2(new_n563), .ZN(new_n566));
  NAND4_X1  g365(.A1(new_n529), .A2(KEYINPUT30), .A3(new_n492), .A4(new_n496), .ZN(new_n567));
  INV_X1    g366(.A(new_n492), .ZN(new_n568));
  OAI21_X1  g367(.A(new_n495), .B1(new_n528), .B2(new_n568), .ZN(new_n569));
  XOR2_X1   g368(.A(KEYINPUT74), .B(KEYINPUT30), .Z(new_n570));
  AND3_X1   g369(.A1(new_n509), .A2(KEYINPUT75), .A3(new_n570), .ZN(new_n571));
  AOI21_X1  g370(.A(KEYINPUT75), .B1(new_n509), .B2(new_n570), .ZN(new_n572));
  OAI211_X1 g371(.A(new_n567), .B(new_n569), .C1(new_n571), .C2(new_n572), .ZN(new_n573));
  AOI21_X1  g372(.A(new_n553), .B1(new_n566), .B2(new_n573), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n533), .A2(new_n574), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n575), .A2(KEYINPUT84), .ZN(new_n576));
  INV_X1    g375(.A(new_n573), .ZN(new_n577));
  INV_X1    g376(.A(new_n422), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  NAND2_X1  g378(.A1(new_n579), .A2(new_n553), .ZN(new_n580));
  INV_X1    g379(.A(KEYINPUT68), .ZN(new_n581));
  NAND3_X1  g380(.A1(new_n490), .A2(new_n581), .A3(new_n400), .ZN(new_n582));
  INV_X1    g381(.A(new_n400), .ZN(new_n583));
  OAI21_X1  g382(.A(KEYINPUT68), .B1(new_n502), .B2(new_n583), .ZN(new_n584));
  NAND2_X1  g383(.A1(new_n502), .A2(new_n583), .ZN(new_n585));
  NAND3_X1  g384(.A1(new_n582), .A2(new_n584), .A3(new_n585), .ZN(new_n586));
  AND2_X1   g385(.A1(G227gat), .A2(G233gat), .ZN(new_n587));
  NAND2_X1  g386(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  NAND2_X1  g387(.A1(new_n588), .A2(KEYINPUT32), .ZN(new_n589));
  NAND2_X1  g388(.A1(new_n589), .A2(KEYINPUT34), .ZN(new_n590));
  INV_X1    g389(.A(KEYINPUT34), .ZN(new_n591));
  NAND3_X1  g390(.A1(new_n588), .A2(KEYINPUT32), .A3(new_n591), .ZN(new_n592));
  NOR2_X1   g391(.A1(new_n586), .A2(new_n587), .ZN(new_n593));
  INV_X1    g392(.A(new_n593), .ZN(new_n594));
  NAND3_X1  g393(.A1(new_n590), .A2(new_n592), .A3(new_n594), .ZN(new_n595));
  AOI21_X1  g394(.A(new_n591), .B1(new_n588), .B2(KEYINPUT32), .ZN(new_n596));
  INV_X1    g395(.A(KEYINPUT32), .ZN(new_n597));
  AOI211_X1 g396(.A(new_n597), .B(KEYINPUT34), .C1(new_n586), .C2(new_n587), .ZN(new_n598));
  OAI21_X1  g397(.A(new_n593), .B1(new_n596), .B2(new_n598), .ZN(new_n599));
  INV_X1    g398(.A(KEYINPUT33), .ZN(new_n600));
  NAND2_X1  g399(.A1(new_n588), .A2(new_n600), .ZN(new_n601));
  XNOR2_X1  g400(.A(G15gat), .B(G43gat), .ZN(new_n602));
  XNOR2_X1  g401(.A(G71gat), .B(G99gat), .ZN(new_n603));
  XOR2_X1   g402(.A(new_n602), .B(new_n603), .Z(new_n604));
  NAND2_X1  g403(.A1(new_n601), .A2(new_n604), .ZN(new_n605));
  INV_X1    g404(.A(new_n605), .ZN(new_n606));
  AND3_X1   g405(.A1(new_n595), .A2(new_n599), .A3(new_n606), .ZN(new_n607));
  AOI21_X1  g406(.A(new_n606), .B1(new_n595), .B2(new_n599), .ZN(new_n608));
  NOR2_X1   g407(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  NAND2_X1  g408(.A1(new_n609), .A2(KEYINPUT36), .ZN(new_n610));
  INV_X1    g409(.A(KEYINPUT36), .ZN(new_n611));
  OAI21_X1  g410(.A(new_n611), .B1(new_n607), .B2(new_n608), .ZN(new_n612));
  NAND2_X1  g411(.A1(new_n610), .A2(new_n612), .ZN(new_n613));
  INV_X1    g412(.A(KEYINPUT84), .ZN(new_n614));
  NAND3_X1  g413(.A1(new_n533), .A2(new_n614), .A3(new_n574), .ZN(new_n615));
  NAND4_X1  g414(.A1(new_n576), .A2(new_n580), .A3(new_n613), .A4(new_n615), .ZN(new_n616));
  INV_X1    g415(.A(new_n553), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n609), .A2(new_n617), .ZN(new_n618));
  OAI21_X1  g417(.A(KEYINPUT35), .B1(new_n618), .B2(new_n579), .ZN(new_n619));
  NOR3_X1   g418(.A1(new_n553), .A2(new_n607), .A3(new_n608), .ZN(new_n620));
  INV_X1    g419(.A(KEYINPUT35), .ZN(new_n621));
  NOR2_X1   g420(.A1(new_n573), .A2(new_n422), .ZN(new_n622));
  NAND3_X1  g421(.A1(new_n620), .A2(new_n621), .A3(new_n622), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n619), .A2(new_n623), .ZN(new_n624));
  NAND2_X1  g423(.A1(new_n616), .A2(new_n624), .ZN(new_n625));
  OAI21_X1  g424(.A(new_n301), .B1(new_n266), .B2(new_n235), .ZN(new_n626));
  NAND2_X1  g425(.A1(G229gat), .A2(G233gat), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n257), .A2(new_n302), .ZN(new_n628));
  NAND4_X1  g427(.A1(new_n626), .A2(KEYINPUT18), .A3(new_n627), .A4(new_n628), .ZN(new_n629));
  XNOR2_X1  g428(.A(new_n627), .B(KEYINPUT13), .ZN(new_n630));
  INV_X1    g429(.A(new_n630), .ZN(new_n631));
  NOR2_X1   g430(.A1(new_n257), .A2(new_n302), .ZN(new_n632));
  NOR2_X1   g431(.A1(new_n232), .A2(new_n301), .ZN(new_n633));
  OAI21_X1  g432(.A(new_n631), .B1(new_n632), .B2(new_n633), .ZN(new_n634));
  NAND2_X1  g433(.A1(new_n629), .A2(new_n634), .ZN(new_n635));
  NAND3_X1  g434(.A1(new_n626), .A2(new_n627), .A3(new_n628), .ZN(new_n636));
  AOI21_X1  g435(.A(KEYINPUT18), .B1(new_n636), .B2(KEYINPUT89), .ZN(new_n637));
  INV_X1    g436(.A(KEYINPUT89), .ZN(new_n638));
  NAND4_X1  g437(.A1(new_n626), .A2(new_n638), .A3(new_n627), .A4(new_n628), .ZN(new_n639));
  AOI21_X1  g438(.A(new_n635), .B1(new_n637), .B2(new_n639), .ZN(new_n640));
  XNOR2_X1  g439(.A(G113gat), .B(G141gat), .ZN(new_n641));
  XNOR2_X1  g440(.A(new_n641), .B(G197gat), .ZN(new_n642));
  XNOR2_X1  g441(.A(KEYINPUT11), .B(G169gat), .ZN(new_n643));
  XNOR2_X1  g442(.A(new_n642), .B(new_n643), .ZN(new_n644));
  XOR2_X1   g443(.A(new_n644), .B(KEYINPUT12), .Z(new_n645));
  INV_X1    g444(.A(new_n645), .ZN(new_n646));
  OAI21_X1  g445(.A(new_n646), .B1(new_n635), .B2(KEYINPUT90), .ZN(new_n647));
  AND2_X1   g446(.A1(new_n640), .A2(new_n647), .ZN(new_n648));
  NOR2_X1   g447(.A1(new_n640), .A2(new_n647), .ZN(new_n649));
  OR2_X1    g448(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  AOI21_X1  g449(.A(KEYINPUT91), .B1(new_n625), .B2(new_n650), .ZN(new_n651));
  INV_X1    g450(.A(KEYINPUT91), .ZN(new_n652));
  INV_X1    g451(.A(new_n650), .ZN(new_n653));
  AOI211_X1 g452(.A(new_n652), .B(new_n653), .C1(new_n616), .C2(new_n624), .ZN(new_n654));
  OAI21_X1  g453(.A(new_n355), .B1(new_n651), .B2(new_n654), .ZN(new_n655));
  INV_X1    g454(.A(KEYINPUT104), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  OAI211_X1 g456(.A(KEYINPUT104), .B(new_n355), .C1(new_n651), .C2(new_n654), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n659), .A2(new_n422), .ZN(new_n660));
  XNOR2_X1  g459(.A(new_n660), .B(G1gat), .ZN(G1324gat));
  NAND2_X1  g460(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n297), .A2(new_n300), .ZN(new_n663));
  NAND4_X1  g462(.A1(new_n659), .A2(new_n573), .A3(new_n662), .A4(new_n663), .ZN(new_n664));
  INV_X1    g463(.A(KEYINPUT42), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  AOI21_X1  g465(.A(new_n577), .B1(new_n657), .B2(new_n658), .ZN(new_n667));
  OR2_X1    g466(.A1(new_n667), .A2(new_n300), .ZN(new_n668));
  NAND4_X1  g467(.A1(new_n667), .A2(KEYINPUT42), .A3(new_n662), .A4(new_n663), .ZN(new_n669));
  NAND3_X1  g468(.A1(new_n666), .A2(new_n668), .A3(new_n669), .ZN(G1325gat));
  AOI21_X1  g469(.A(G15gat), .B1(new_n659), .B2(new_n609), .ZN(new_n671));
  INV_X1    g470(.A(new_n613), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n672), .A2(G15gat), .ZN(new_n673));
  XNOR2_X1  g472(.A(new_n673), .B(KEYINPUT105), .ZN(new_n674));
  AOI21_X1  g473(.A(new_n671), .B1(new_n659), .B2(new_n674), .ZN(G1326gat));
  NAND2_X1  g474(.A1(new_n659), .A2(new_n553), .ZN(new_n676));
  XNOR2_X1  g475(.A(KEYINPUT43), .B(G22gat), .ZN(new_n677));
  XNOR2_X1  g476(.A(new_n676), .B(new_n677), .ZN(G1327gat));
  AND3_X1   g477(.A1(new_n533), .A2(new_n614), .A3(new_n574), .ZN(new_n679));
  AOI21_X1  g478(.A(new_n614), .B1(new_n533), .B2(new_n574), .ZN(new_n680));
  NOR3_X1   g479(.A1(new_n607), .A2(new_n608), .A3(new_n611), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n595), .A2(new_n599), .ZN(new_n682));
  NAND2_X1  g481(.A1(new_n682), .A2(new_n605), .ZN(new_n683));
  NAND3_X1  g482(.A1(new_n595), .A2(new_n599), .A3(new_n606), .ZN(new_n684));
  AOI21_X1  g483(.A(KEYINPUT36), .B1(new_n683), .B2(new_n684), .ZN(new_n685));
  OAI22_X1  g484(.A1(new_n681), .A2(new_n685), .B1(new_n622), .B2(new_n617), .ZN(new_n686));
  NOR3_X1   g485(.A1(new_n679), .A2(new_n680), .A3(new_n686), .ZN(new_n687));
  AND2_X1   g486(.A1(new_n619), .A2(new_n623), .ZN(new_n688));
  OAI21_X1  g487(.A(new_n279), .B1(new_n687), .B2(new_n688), .ZN(new_n689));
  INV_X1    g488(.A(KEYINPUT44), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  INV_X1    g490(.A(new_n279), .ZN(new_n692));
  AOI21_X1  g491(.A(new_n692), .B1(new_n616), .B2(new_n624), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n693), .A2(KEYINPUT44), .ZN(new_n694));
  INV_X1    g493(.A(new_n353), .ZN(new_n695));
  INV_X1    g494(.A(new_n310), .ZN(new_n696));
  NOR2_X1   g495(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  NAND4_X1  g496(.A1(new_n691), .A2(new_n694), .A3(new_n650), .A4(new_n697), .ZN(new_n698));
  OAI21_X1  g497(.A(new_n222), .B1(new_n698), .B2(new_n578), .ZN(new_n699));
  INV_X1    g498(.A(new_n697), .ZN(new_n700));
  OAI21_X1  g499(.A(new_n650), .B1(new_n687), .B2(new_n688), .ZN(new_n701));
  NAND2_X1  g500(.A1(new_n701), .A2(new_n652), .ZN(new_n702));
  NAND3_X1  g501(.A1(new_n625), .A2(KEYINPUT91), .A3(new_n650), .ZN(new_n703));
  AOI21_X1  g502(.A(new_n700), .B1(new_n702), .B2(new_n703), .ZN(new_n704));
  INV_X1    g503(.A(new_n222), .ZN(new_n705));
  NAND4_X1  g504(.A1(new_n704), .A2(new_n422), .A3(new_n705), .A4(new_n279), .ZN(new_n706));
  NAND3_X1  g505(.A1(new_n699), .A2(new_n706), .A3(KEYINPUT45), .ZN(new_n707));
  INV_X1    g506(.A(KEYINPUT106), .ZN(new_n708));
  AOI211_X1 g507(.A(new_n692), .B(new_n700), .C1(new_n702), .C2(new_n703), .ZN(new_n709));
  INV_X1    g508(.A(KEYINPUT45), .ZN(new_n710));
  NAND4_X1  g509(.A1(new_n709), .A2(new_n710), .A3(new_n422), .A4(new_n705), .ZN(new_n711));
  AND3_X1   g510(.A1(new_n707), .A2(new_n708), .A3(new_n711), .ZN(new_n712));
  AOI21_X1  g511(.A(new_n708), .B1(new_n707), .B2(new_n711), .ZN(new_n713));
  NOR2_X1   g512(.A1(new_n712), .A2(new_n713), .ZN(G1328gat));
  NAND3_X1  g513(.A1(new_n709), .A2(new_n208), .A3(new_n573), .ZN(new_n715));
  OR2_X1    g514(.A1(new_n715), .A2(KEYINPUT46), .ZN(new_n716));
  OAI21_X1  g515(.A(G36gat), .B1(new_n698), .B2(new_n577), .ZN(new_n717));
  NAND2_X1  g516(.A1(new_n715), .A2(KEYINPUT46), .ZN(new_n718));
  NAND3_X1  g517(.A1(new_n716), .A2(new_n717), .A3(new_n718), .ZN(G1329gat));
  INV_X1    g518(.A(G43gat), .ZN(new_n720));
  NAND3_X1  g519(.A1(new_n709), .A2(new_n720), .A3(new_n609), .ZN(new_n721));
  OAI21_X1  g520(.A(G43gat), .B1(new_n698), .B2(new_n613), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  INV_X1    g522(.A(KEYINPUT47), .ZN(new_n724));
  XNOR2_X1  g523(.A(new_n723), .B(new_n724), .ZN(G1330gat));
  INV_X1    g524(.A(G50gat), .ZN(new_n726));
  NAND3_X1  g525(.A1(new_n709), .A2(new_n726), .A3(new_n553), .ZN(new_n727));
  OAI21_X1  g526(.A(G50gat), .B1(new_n698), .B2(new_n617), .ZN(new_n728));
  NAND2_X1  g527(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  INV_X1    g528(.A(KEYINPUT48), .ZN(new_n730));
  XNOR2_X1  g529(.A(new_n729), .B(new_n730), .ZN(G1331gat));
  AOI21_X1  g530(.A(new_n650), .B1(new_n616), .B2(new_n624), .ZN(new_n732));
  NOR3_X1   g531(.A1(new_n279), .A2(new_n353), .A3(new_n310), .ZN(new_n733));
  AND2_X1   g532(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n734), .A2(new_n422), .ZN(new_n735));
  XNOR2_X1  g534(.A(new_n735), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g535(.A1(new_n732), .A2(new_n733), .ZN(new_n737));
  NOR2_X1   g536(.A1(new_n737), .A2(new_n577), .ZN(new_n738));
  NOR2_X1   g537(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n739));
  AND2_X1   g538(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n740));
  OAI21_X1  g539(.A(new_n738), .B1(new_n739), .B2(new_n740), .ZN(new_n741));
  OAI21_X1  g540(.A(new_n741), .B1(new_n738), .B2(new_n739), .ZN(G1333gat));
  INV_X1    g541(.A(G71gat), .ZN(new_n743));
  NAND3_X1  g542(.A1(new_n734), .A2(new_n743), .A3(new_n609), .ZN(new_n744));
  OAI21_X1  g543(.A(G71gat), .B1(new_n737), .B2(new_n613), .ZN(new_n745));
  NAND2_X1  g544(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  NAND2_X1  g545(.A1(new_n746), .A2(KEYINPUT107), .ZN(new_n747));
  INV_X1    g546(.A(KEYINPUT107), .ZN(new_n748));
  NAND3_X1  g547(.A1(new_n744), .A2(new_n748), .A3(new_n745), .ZN(new_n749));
  NAND2_X1  g548(.A1(new_n747), .A2(new_n749), .ZN(new_n750));
  INV_X1    g549(.A(KEYINPUT50), .ZN(new_n751));
  XNOR2_X1  g550(.A(new_n750), .B(new_n751), .ZN(G1334gat));
  NAND2_X1  g551(.A1(new_n734), .A2(new_n553), .ZN(new_n753));
  XNOR2_X1  g552(.A(new_n753), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g553(.A1(new_n650), .A2(new_n696), .ZN(new_n755));
  AND4_X1   g554(.A1(new_n695), .A2(new_n691), .A3(new_n694), .A4(new_n755), .ZN(new_n756));
  INV_X1    g555(.A(new_n756), .ZN(new_n757));
  OAI21_X1  g556(.A(G85gat), .B1(new_n757), .B2(new_n578), .ZN(new_n758));
  NAND4_X1  g557(.A1(new_n625), .A2(KEYINPUT51), .A3(new_n279), .A4(new_n755), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n759), .A2(KEYINPUT108), .ZN(new_n760));
  INV_X1    g559(.A(KEYINPUT108), .ZN(new_n761));
  NAND4_X1  g560(.A1(new_n693), .A2(new_n761), .A3(KEYINPUT51), .A4(new_n755), .ZN(new_n762));
  NAND3_X1  g561(.A1(new_n760), .A2(KEYINPUT109), .A3(new_n762), .ZN(new_n763));
  INV_X1    g562(.A(KEYINPUT51), .ZN(new_n764));
  INV_X1    g563(.A(new_n755), .ZN(new_n765));
  OAI21_X1  g564(.A(new_n764), .B1(new_n689), .B2(new_n765), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n763), .A2(new_n766), .ZN(new_n767));
  AOI21_X1  g566(.A(KEYINPUT109), .B1(new_n760), .B2(new_n762), .ZN(new_n768));
  OAI21_X1  g567(.A(new_n695), .B1(new_n767), .B2(new_n768), .ZN(new_n769));
  NAND2_X1  g568(.A1(new_n422), .A2(new_n238), .ZN(new_n770));
  OAI21_X1  g569(.A(new_n758), .B1(new_n769), .B2(new_n770), .ZN(G1336gat));
  AOI21_X1  g570(.A(new_n239), .B1(new_n756), .B2(new_n573), .ZN(new_n772));
  NOR2_X1   g571(.A1(new_n772), .A2(KEYINPUT52), .ZN(new_n773));
  NOR2_X1   g572(.A1(new_n767), .A2(new_n768), .ZN(new_n774));
  NAND3_X1  g573(.A1(new_n695), .A2(new_n239), .A3(new_n573), .ZN(new_n775));
  XNOR2_X1  g574(.A(new_n775), .B(KEYINPUT110), .ZN(new_n776));
  OAI21_X1  g575(.A(new_n773), .B1(new_n774), .B2(new_n776), .ZN(new_n777));
  NAND2_X1  g576(.A1(new_n760), .A2(new_n762), .ZN(new_n778));
  AOI21_X1  g577(.A(new_n776), .B1(new_n778), .B2(new_n766), .ZN(new_n779));
  OAI21_X1  g578(.A(KEYINPUT52), .B1(new_n772), .B2(new_n779), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n777), .A2(new_n780), .ZN(G1337gat));
  OAI21_X1  g580(.A(G99gat), .B1(new_n757), .B2(new_n613), .ZN(new_n782));
  INV_X1    g581(.A(G99gat), .ZN(new_n783));
  NAND3_X1  g582(.A1(new_n695), .A2(new_n783), .A3(new_n609), .ZN(new_n784));
  XNOR2_X1  g583(.A(new_n784), .B(KEYINPUT111), .ZN(new_n785));
  OAI21_X1  g584(.A(new_n782), .B1(new_n774), .B2(new_n785), .ZN(G1338gat));
  INV_X1    g585(.A(G106gat), .ZN(new_n787));
  AOI21_X1  g586(.A(new_n787), .B1(new_n756), .B2(new_n553), .ZN(new_n788));
  NOR2_X1   g587(.A1(new_n788), .A2(KEYINPUT53), .ZN(new_n789));
  NOR2_X1   g588(.A1(new_n617), .A2(G106gat), .ZN(new_n790));
  INV_X1    g589(.A(new_n790), .ZN(new_n791));
  OAI21_X1  g590(.A(new_n789), .B1(new_n769), .B2(new_n791), .ZN(new_n792));
  AOI211_X1 g591(.A(new_n353), .B(new_n791), .C1(new_n778), .C2(new_n766), .ZN(new_n793));
  OAI21_X1  g592(.A(KEYINPUT53), .B1(new_n793), .B2(new_n788), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n792), .A2(new_n794), .ZN(G1339gat));
  INV_X1    g594(.A(KEYINPUT112), .ZN(new_n796));
  NAND3_X1  g595(.A1(new_n314), .A2(new_n313), .A3(new_n327), .ZN(new_n797));
  OAI211_X1 g596(.A(new_n797), .B(KEYINPUT54), .C1(new_n341), .C2(new_n343), .ZN(new_n798));
  INV_X1    g597(.A(KEYINPUT54), .ZN(new_n799));
  AOI21_X1  g598(.A(new_n336), .B1(new_n328), .B2(new_n799), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n798), .A2(new_n800), .ZN(new_n801));
  INV_X1    g600(.A(KEYINPUT55), .ZN(new_n802));
  AOI21_X1  g601(.A(new_n796), .B1(new_n801), .B2(new_n802), .ZN(new_n803));
  AOI211_X1 g602(.A(KEYINPUT112), .B(KEYINPUT55), .C1(new_n798), .C2(new_n800), .ZN(new_n804));
  NOR2_X1   g603(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  NAND3_X1  g604(.A1(new_n798), .A2(KEYINPUT55), .A3(new_n800), .ZN(new_n806));
  AND2_X1   g605(.A1(new_n346), .A2(new_n806), .ZN(new_n807));
  OAI211_X1 g606(.A(new_n805), .B(new_n807), .C1(new_n648), .C2(new_n649), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n626), .A2(new_n628), .ZN(new_n809));
  NAND3_X1  g608(.A1(new_n809), .A2(G229gat), .A3(G233gat), .ZN(new_n810));
  OR3_X1    g609(.A1(new_n632), .A2(new_n633), .A3(new_n631), .ZN(new_n811));
  AOI21_X1  g610(.A(new_n644), .B1(new_n810), .B2(new_n811), .ZN(new_n812));
  AOI21_X1  g611(.A(new_n812), .B1(new_n640), .B2(new_n645), .ZN(new_n813));
  OAI21_X1  g612(.A(new_n813), .B1(new_n349), .B2(new_n352), .ZN(new_n814));
  AOI21_X1  g613(.A(new_n279), .B1(new_n808), .B2(new_n814), .ZN(new_n815));
  NAND3_X1  g614(.A1(new_n277), .A2(new_n813), .A3(new_n278), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n805), .A2(new_n807), .ZN(new_n817));
  NOR2_X1   g616(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  OAI21_X1  g617(.A(new_n310), .B1(new_n815), .B2(new_n818), .ZN(new_n819));
  NAND3_X1  g618(.A1(new_n311), .A2(new_n653), .A3(new_n353), .ZN(new_n820));
  AOI21_X1  g619(.A(new_n618), .B1(new_n819), .B2(new_n820), .ZN(new_n821));
  NAND3_X1  g620(.A1(new_n821), .A2(new_n422), .A3(new_n577), .ZN(new_n822));
  OAI21_X1  g621(.A(G113gat), .B1(new_n822), .B2(new_n653), .ZN(new_n823));
  AND3_X1   g622(.A1(new_n821), .A2(KEYINPUT113), .A3(new_n422), .ZN(new_n824));
  AOI21_X1  g623(.A(KEYINPUT113), .B1(new_n821), .B2(new_n422), .ZN(new_n825));
  NOR3_X1   g624(.A1(new_n824), .A2(new_n825), .A3(new_n573), .ZN(new_n826));
  INV_X1    g625(.A(new_n826), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n650), .A2(new_n358), .ZN(new_n828));
  OAI21_X1  g627(.A(new_n823), .B1(new_n827), .B2(new_n828), .ZN(G1340gat));
  OAI21_X1  g628(.A(G120gat), .B1(new_n822), .B2(new_n353), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n695), .A2(new_n356), .ZN(new_n831));
  OAI21_X1  g630(.A(new_n830), .B1(new_n827), .B2(new_n831), .ZN(G1341gat));
  NOR3_X1   g631(.A1(new_n822), .A2(new_n366), .A3(new_n310), .ZN(new_n833));
  NAND2_X1  g632(.A1(new_n826), .A2(new_n696), .ZN(new_n834));
  AOI21_X1  g633(.A(new_n833), .B1(new_n834), .B2(new_n366), .ZN(G1342gat));
  INV_X1    g634(.A(KEYINPUT56), .ZN(new_n836));
  NAND4_X1  g635(.A1(new_n826), .A2(new_n836), .A3(new_n364), .A4(new_n279), .ZN(new_n837));
  OAI21_X1  g636(.A(G134gat), .B1(new_n822), .B2(new_n692), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n819), .A2(new_n820), .ZN(new_n839));
  NAND3_X1  g638(.A1(new_n839), .A2(new_n422), .A3(new_n620), .ZN(new_n840));
  INV_X1    g639(.A(KEYINPUT113), .ZN(new_n841));
  NAND2_X1  g640(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  NAND3_X1  g641(.A1(new_n821), .A2(KEYINPUT113), .A3(new_n422), .ZN(new_n843));
  NAND4_X1  g642(.A1(new_n842), .A2(new_n577), .A3(new_n279), .A4(new_n843), .ZN(new_n844));
  OAI21_X1  g643(.A(KEYINPUT56), .B1(new_n844), .B2(G134gat), .ZN(new_n845));
  NAND3_X1  g644(.A1(new_n837), .A2(new_n838), .A3(new_n845), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n846), .A2(KEYINPUT114), .ZN(new_n847));
  INV_X1    g646(.A(KEYINPUT114), .ZN(new_n848));
  NAND4_X1  g647(.A1(new_n837), .A2(new_n845), .A3(new_n848), .A4(new_n838), .ZN(new_n849));
  NAND2_X1  g648(.A1(new_n847), .A2(new_n849), .ZN(G1343gat));
  INV_X1    g649(.A(new_n820), .ZN(new_n851));
  NAND2_X1  g650(.A1(new_n801), .A2(new_n802), .ZN(new_n852));
  NAND3_X1  g651(.A1(new_n650), .A2(new_n852), .A3(new_n807), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n853), .A2(new_n814), .ZN(new_n854));
  NAND2_X1  g653(.A1(new_n854), .A2(new_n692), .ZN(new_n855));
  INV_X1    g654(.A(new_n818), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n855), .A2(new_n856), .ZN(new_n857));
  AOI21_X1  g656(.A(new_n851), .B1(new_n857), .B2(new_n310), .ZN(new_n858));
  OAI21_X1  g657(.A(KEYINPUT57), .B1(new_n858), .B2(new_n617), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n839), .A2(new_n553), .ZN(new_n860));
  NOR2_X1   g659(.A1(new_n860), .A2(KEYINPUT57), .ZN(new_n861));
  INV_X1    g660(.A(new_n861), .ZN(new_n862));
  NOR3_X1   g661(.A1(new_n672), .A2(new_n578), .A3(new_n573), .ZN(new_n863));
  NAND3_X1  g662(.A1(new_n859), .A2(new_n862), .A3(new_n863), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n650), .A2(G141gat), .ZN(new_n865));
  INV_X1    g664(.A(new_n860), .ZN(new_n866));
  NAND2_X1  g665(.A1(new_n866), .A2(new_n863), .ZN(new_n867));
  NOR2_X1   g666(.A1(new_n867), .A2(new_n653), .ZN(new_n868));
  OAI22_X1  g667(.A1(new_n864), .A2(new_n865), .B1(G141gat), .B2(new_n868), .ZN(new_n869));
  XNOR2_X1  g668(.A(KEYINPUT115), .B(KEYINPUT58), .ZN(new_n870));
  XNOR2_X1  g669(.A(new_n869), .B(new_n870), .ZN(G1344gat));
  OR3_X1    g670(.A1(new_n867), .A2(G148gat), .A3(new_n353), .ZN(new_n872));
  INV_X1    g671(.A(KEYINPUT59), .ZN(new_n873));
  NOR2_X1   g672(.A1(new_n617), .A2(KEYINPUT57), .ZN(new_n874));
  INV_X1    g673(.A(KEYINPUT116), .ZN(new_n875));
  NAND3_X1  g674(.A1(new_n855), .A2(new_n875), .A3(new_n856), .ZN(new_n876));
  AOI21_X1  g675(.A(new_n279), .B1(new_n853), .B2(new_n814), .ZN(new_n877));
  OAI21_X1  g676(.A(KEYINPUT116), .B1(new_n877), .B2(new_n818), .ZN(new_n878));
  AND3_X1   g677(.A1(new_n876), .A2(new_n310), .A3(new_n878), .ZN(new_n879));
  AND2_X1   g678(.A1(new_n355), .A2(new_n653), .ZN(new_n880));
  OAI21_X1  g679(.A(new_n874), .B1(new_n879), .B2(new_n880), .ZN(new_n881));
  NAND2_X1  g680(.A1(new_n860), .A2(KEYINPUT57), .ZN(new_n882));
  NAND4_X1  g681(.A1(new_n881), .A2(new_n695), .A3(new_n863), .A4(new_n882), .ZN(new_n883));
  AOI21_X1  g682(.A(new_n873), .B1(new_n883), .B2(G148gat), .ZN(new_n884));
  NAND4_X1  g683(.A1(new_n859), .A2(new_n862), .A3(new_n695), .A4(new_n863), .ZN(new_n885));
  AND3_X1   g684(.A1(new_n885), .A2(new_n873), .A3(G148gat), .ZN(new_n886));
  OAI21_X1  g685(.A(new_n872), .B1(new_n884), .B2(new_n886), .ZN(G1345gat));
  INV_X1    g686(.A(G155gat), .ZN(new_n888));
  NOR3_X1   g687(.A1(new_n864), .A2(new_n888), .A3(new_n310), .ZN(new_n889));
  OAI21_X1  g688(.A(new_n888), .B1(new_n867), .B2(new_n310), .ZN(new_n890));
  INV_X1    g689(.A(new_n890), .ZN(new_n891));
  OAI21_X1  g690(.A(KEYINPUT117), .B1(new_n889), .B2(new_n891), .ZN(new_n892));
  INV_X1    g691(.A(KEYINPUT117), .ZN(new_n893));
  NOR2_X1   g692(.A1(new_n310), .A2(new_n888), .ZN(new_n894));
  INV_X1    g693(.A(new_n894), .ZN(new_n895));
  OAI211_X1 g694(.A(new_n893), .B(new_n890), .C1(new_n864), .C2(new_n895), .ZN(new_n896));
  NAND2_X1  g695(.A1(new_n892), .A2(new_n896), .ZN(G1346gat));
  INV_X1    g696(.A(new_n867), .ZN(new_n898));
  AOI21_X1  g697(.A(G162gat), .B1(new_n898), .B2(new_n279), .ZN(new_n899));
  NAND2_X1  g698(.A1(new_n859), .A2(new_n863), .ZN(new_n900));
  NOR2_X1   g699(.A1(new_n900), .A2(new_n861), .ZN(new_n901));
  AND2_X1   g700(.A1(new_n279), .A2(G162gat), .ZN(new_n902));
  AOI21_X1  g701(.A(new_n899), .B1(new_n901), .B2(new_n902), .ZN(G1347gat));
  NAND3_X1  g702(.A1(new_n821), .A2(new_n578), .A3(new_n573), .ZN(new_n904));
  NOR3_X1   g703(.A1(new_n904), .A2(G169gat), .A3(new_n653), .ZN(new_n905));
  XNOR2_X1  g704(.A(new_n905), .B(KEYINPUT118), .ZN(new_n906));
  AND3_X1   g705(.A1(new_n821), .A2(new_n578), .A3(new_n573), .ZN(new_n907));
  NAND2_X1  g706(.A1(new_n907), .A2(KEYINPUT119), .ZN(new_n908));
  INV_X1    g707(.A(KEYINPUT119), .ZN(new_n909));
  NAND2_X1  g708(.A1(new_n904), .A2(new_n909), .ZN(new_n910));
  AND2_X1   g709(.A1(new_n908), .A2(new_n910), .ZN(new_n911));
  AND2_X1   g710(.A1(new_n911), .A2(new_n650), .ZN(new_n912));
  OAI21_X1  g711(.A(new_n906), .B1(new_n912), .B2(new_n445), .ZN(G1348gat));
  AOI21_X1  g712(.A(G176gat), .B1(new_n907), .B2(new_n695), .ZN(new_n914));
  XNOR2_X1  g713(.A(new_n914), .B(KEYINPUT120), .ZN(new_n915));
  NAND3_X1  g714(.A1(new_n911), .A2(G176gat), .A3(new_n695), .ZN(new_n916));
  NAND2_X1  g715(.A1(new_n916), .A2(KEYINPUT121), .ZN(new_n917));
  INV_X1    g716(.A(KEYINPUT121), .ZN(new_n918));
  NAND4_X1  g717(.A1(new_n911), .A2(new_n918), .A3(G176gat), .A4(new_n695), .ZN(new_n919));
  AOI21_X1  g718(.A(new_n915), .B1(new_n917), .B2(new_n919), .ZN(G1349gat));
  NAND3_X1  g719(.A1(new_n908), .A2(new_n696), .A3(new_n910), .ZN(new_n921));
  NAND2_X1  g720(.A1(new_n921), .A2(G183gat), .ZN(new_n922));
  NAND3_X1  g721(.A1(new_n907), .A2(new_n465), .A3(new_n696), .ZN(new_n923));
  NAND2_X1  g722(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  NAND2_X1  g723(.A1(new_n924), .A2(KEYINPUT60), .ZN(new_n925));
  INV_X1    g724(.A(KEYINPUT60), .ZN(new_n926));
  NAND3_X1  g725(.A1(new_n922), .A2(new_n926), .A3(new_n923), .ZN(new_n927));
  NAND2_X1  g726(.A1(new_n925), .A2(new_n927), .ZN(G1350gat));
  NAND3_X1  g727(.A1(new_n907), .A2(new_n464), .A3(new_n279), .ZN(new_n929));
  NAND3_X1  g728(.A1(new_n908), .A2(new_n279), .A3(new_n910), .ZN(new_n930));
  INV_X1    g729(.A(KEYINPUT61), .ZN(new_n931));
  AND3_X1   g730(.A1(new_n930), .A2(new_n931), .A3(G190gat), .ZN(new_n932));
  AOI21_X1  g731(.A(new_n931), .B1(new_n930), .B2(G190gat), .ZN(new_n933));
  OAI21_X1  g732(.A(new_n929), .B1(new_n932), .B2(new_n933), .ZN(G1351gat));
  AOI21_X1  g733(.A(new_n577), .B1(new_n610), .B2(new_n612), .ZN(new_n935));
  NAND2_X1  g734(.A1(new_n935), .A2(new_n578), .ZN(new_n936));
  INV_X1    g735(.A(new_n936), .ZN(new_n937));
  NOR2_X1   g736(.A1(new_n653), .A2(new_n425), .ZN(new_n938));
  NAND4_X1  g737(.A1(new_n881), .A2(new_n882), .A3(new_n937), .A4(new_n938), .ZN(new_n939));
  AOI21_X1  g738(.A(new_n422), .B1(new_n819), .B2(new_n820), .ZN(new_n940));
  NAND2_X1  g739(.A1(new_n935), .A2(new_n553), .ZN(new_n941));
  XNOR2_X1  g740(.A(new_n941), .B(KEYINPUT122), .ZN(new_n942));
  AND2_X1   g741(.A1(new_n940), .A2(new_n942), .ZN(new_n943));
  NAND2_X1  g742(.A1(new_n943), .A2(new_n650), .ZN(new_n944));
  INV_X1    g743(.A(new_n944), .ZN(new_n945));
  OAI21_X1  g744(.A(new_n939), .B1(G197gat), .B2(new_n945), .ZN(new_n946));
  INV_X1    g745(.A(KEYINPUT123), .ZN(new_n947));
  NAND2_X1  g746(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  OAI211_X1 g747(.A(new_n939), .B(KEYINPUT123), .C1(G197gat), .C2(new_n945), .ZN(new_n949));
  NAND2_X1  g748(.A1(new_n948), .A2(new_n949), .ZN(G1352gat));
  NAND4_X1  g749(.A1(new_n940), .A2(new_n942), .A3(new_n332), .A4(new_n695), .ZN(new_n951));
  INV_X1    g750(.A(KEYINPUT124), .ZN(new_n952));
  OR2_X1    g751(.A1(new_n951), .A2(new_n952), .ZN(new_n953));
  NAND2_X1  g752(.A1(new_n951), .A2(new_n952), .ZN(new_n954));
  AND2_X1   g753(.A1(new_n953), .A2(new_n954), .ZN(new_n955));
  INV_X1    g754(.A(KEYINPUT62), .ZN(new_n956));
  OR2_X1    g755(.A1(new_n955), .A2(new_n956), .ZN(new_n957));
  NAND3_X1  g756(.A1(new_n881), .A2(new_n695), .A3(new_n882), .ZN(new_n958));
  OAI21_X1  g757(.A(G204gat), .B1(new_n958), .B2(new_n936), .ZN(new_n959));
  AOI21_X1  g758(.A(KEYINPUT125), .B1(new_n955), .B2(new_n956), .ZN(new_n960));
  AND4_X1   g759(.A1(KEYINPUT125), .A2(new_n953), .A3(new_n956), .A4(new_n954), .ZN(new_n961));
  OAI211_X1 g760(.A(new_n957), .B(new_n959), .C1(new_n960), .C2(new_n961), .ZN(G1353gat));
  NAND4_X1  g761(.A1(new_n881), .A2(new_n696), .A3(new_n882), .A4(new_n937), .ZN(new_n963));
  NAND2_X1  g762(.A1(new_n963), .A2(G211gat), .ZN(new_n964));
  NAND2_X1  g763(.A1(new_n964), .A2(KEYINPUT63), .ZN(new_n965));
  INV_X1    g764(.A(KEYINPUT63), .ZN(new_n966));
  NAND3_X1  g765(.A1(new_n963), .A2(new_n966), .A3(G211gat), .ZN(new_n967));
  NAND3_X1  g766(.A1(new_n943), .A2(new_n428), .A3(new_n696), .ZN(new_n968));
  XNOR2_X1  g767(.A(new_n968), .B(KEYINPUT126), .ZN(new_n969));
  NAND3_X1  g768(.A1(new_n965), .A2(new_n967), .A3(new_n969), .ZN(G1354gat));
  NAND3_X1  g769(.A1(new_n881), .A2(new_n882), .A3(new_n937), .ZN(new_n971));
  NOR3_X1   g770(.A1(new_n971), .A2(new_n429), .A3(new_n692), .ZN(new_n972));
  AOI21_X1  g771(.A(G218gat), .B1(new_n943), .B2(new_n279), .ZN(new_n973));
  XOR2_X1   g772(.A(new_n973), .B(KEYINPUT127), .Z(new_n974));
  NOR2_X1   g773(.A1(new_n972), .A2(new_n974), .ZN(G1355gat));
endmodule


