//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 0 0 1 0 1 0 0 1 1 0 1 0 1 0 1 0 1 0 1 1 0 0 0 1 0 0 0 0 0 0 0 0 0 0 0 1 0 0 0 0 0 1 1 0 1 0 0 1 1 0 0 0 1 1 1 1 1 1 0 1 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:28:59 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n454, new_n458,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n527, new_n528, new_n529, new_n530, new_n531, new_n532,
    new_n533, new_n535, new_n536, new_n537, new_n538, new_n539, new_n542,
    new_n543, new_n544, new_n545, new_n546, new_n547, new_n550, new_n551,
    new_n553, new_n554, new_n555, new_n556, new_n557, new_n558, new_n559,
    new_n560, new_n562, new_n565, new_n566, new_n567, new_n569, new_n570,
    new_n571, new_n572, new_n573, new_n574, new_n576, new_n577, new_n578,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n594, new_n597,
    new_n599, new_n600, new_n601, new_n602, new_n603, new_n604, new_n605,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1123, new_n1124,
    new_n1125;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n450), .B(KEYINPUT2), .ZN(new_n451));
  INV_X1    g026(.A(new_n451), .ZN(new_n452));
  NOR4_X1   g027(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NOR2_X1   g029(.A1(new_n452), .A2(new_n454), .ZN(G325));
  INV_X1    g030(.A(G325), .ZN(G261));
  AOI22_X1  g031(.A1(new_n452), .A2(G2106), .B1(G567), .B2(new_n454), .ZN(G319));
  INV_X1    g032(.A(G2105), .ZN(new_n458));
  AND2_X1   g033(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n459));
  NOR2_X1   g034(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n460));
  OAI21_X1  g035(.A(G125), .B1(new_n459), .B2(new_n460), .ZN(new_n461));
  NAND2_X1  g036(.A1(G113), .A2(G2104), .ZN(new_n462));
  AOI21_X1  g037(.A(new_n458), .B1(new_n461), .B2(new_n462), .ZN(new_n463));
  OAI211_X1 g038(.A(G137), .B(new_n458), .C1(new_n459), .C2(new_n460), .ZN(new_n464));
  INV_X1    g039(.A(G2104), .ZN(new_n465));
  NOR2_X1   g040(.A1(new_n465), .A2(G2105), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n466), .A2(G101), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n464), .A2(new_n467), .ZN(new_n468));
  NOR2_X1   g043(.A1(new_n463), .A2(new_n468), .ZN(G160));
  NOR2_X1   g044(.A1(new_n459), .A2(new_n460), .ZN(new_n470));
  INV_X1    g045(.A(KEYINPUT64), .ZN(new_n471));
  NOR2_X1   g046(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  NOR3_X1   g047(.A1(new_n459), .A2(new_n460), .A3(KEYINPUT64), .ZN(new_n473));
  NOR2_X1   g048(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  NOR2_X1   g049(.A1(new_n474), .A2(new_n458), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n475), .A2(G124), .ZN(new_n476));
  OAI21_X1  g051(.A(new_n458), .B1(new_n472), .B2(new_n473), .ZN(new_n477));
  INV_X1    g052(.A(new_n477), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n478), .A2(G136), .ZN(new_n479));
  NOR2_X1   g054(.A1(new_n458), .A2(G112), .ZN(new_n480));
  OAI21_X1  g055(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n481));
  OAI211_X1 g056(.A(new_n476), .B(new_n479), .C1(new_n480), .C2(new_n481), .ZN(new_n482));
  XOR2_X1   g057(.A(new_n482), .B(KEYINPUT65), .Z(G162));
  NAND2_X1  g058(.A1(KEYINPUT4), .A2(G138), .ZN(new_n484));
  INV_X1    g059(.A(new_n484), .ZN(new_n485));
  OAI21_X1  g060(.A(new_n485), .B1(new_n459), .B2(new_n460), .ZN(new_n486));
  NAND2_X1  g061(.A1(G102), .A2(G2104), .ZN(new_n487));
  AOI21_X1  g062(.A(G2105), .B1(new_n486), .B2(new_n487), .ZN(new_n488));
  OAI21_X1  g063(.A(G126), .B1(new_n459), .B2(new_n460), .ZN(new_n489));
  NAND2_X1  g064(.A1(G114), .A2(G2104), .ZN(new_n490));
  AOI21_X1  g065(.A(new_n458), .B1(new_n489), .B2(new_n490), .ZN(new_n491));
  NOR2_X1   g066(.A1(new_n488), .A2(new_n491), .ZN(new_n492));
  OAI211_X1 g067(.A(G138), .B(new_n458), .C1(new_n459), .C2(new_n460), .ZN(new_n493));
  INV_X1    g068(.A(KEYINPUT4), .ZN(new_n494));
  NAND2_X1  g069(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  AOI21_X1  g070(.A(KEYINPUT66), .B1(new_n492), .B2(new_n495), .ZN(new_n496));
  INV_X1    g071(.A(KEYINPUT3), .ZN(new_n497));
  NAND2_X1  g072(.A1(new_n497), .A2(new_n465), .ZN(new_n498));
  NAND2_X1  g073(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n499));
  AOI21_X1  g074(.A(new_n484), .B1(new_n498), .B2(new_n499), .ZN(new_n500));
  INV_X1    g075(.A(new_n487), .ZN(new_n501));
  OAI21_X1  g076(.A(new_n458), .B1(new_n500), .B2(new_n501), .ZN(new_n502));
  INV_X1    g077(.A(G126), .ZN(new_n503));
  AOI21_X1  g078(.A(new_n503), .B1(new_n498), .B2(new_n499), .ZN(new_n504));
  INV_X1    g079(.A(new_n490), .ZN(new_n505));
  OAI21_X1  g080(.A(G2105), .B1(new_n504), .B2(new_n505), .ZN(new_n506));
  NAND4_X1  g081(.A1(new_n502), .A2(new_n506), .A3(KEYINPUT66), .A4(new_n495), .ZN(new_n507));
  INV_X1    g082(.A(new_n507), .ZN(new_n508));
  NOR2_X1   g083(.A1(new_n496), .A2(new_n508), .ZN(G164));
  INV_X1    g084(.A(G651), .ZN(new_n510));
  XNOR2_X1  g085(.A(KEYINPUT5), .B(G543), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n511), .A2(G62), .ZN(new_n512));
  NAND2_X1  g087(.A1(G75), .A2(G543), .ZN(new_n513));
  XNOR2_X1  g088(.A(new_n513), .B(KEYINPUT68), .ZN(new_n514));
  AOI21_X1  g089(.A(new_n510), .B1(new_n512), .B2(new_n514), .ZN(new_n515));
  INV_X1    g090(.A(G50), .ZN(new_n516));
  AND2_X1   g091(.A1(KEYINPUT6), .A2(G651), .ZN(new_n517));
  NOR2_X1   g092(.A1(KEYINPUT6), .A2(G651), .ZN(new_n518));
  OR2_X1    g093(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n519), .A2(G543), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n519), .A2(new_n511), .ZN(new_n521));
  INV_X1    g096(.A(G88), .ZN(new_n522));
  OAI22_X1  g097(.A1(new_n516), .A2(new_n520), .B1(new_n521), .B2(new_n522), .ZN(new_n523));
  OR2_X1    g098(.A1(new_n523), .A2(KEYINPUT67), .ZN(new_n524));
  NAND2_X1  g099(.A1(new_n523), .A2(KEYINPUT67), .ZN(new_n525));
  AOI21_X1  g100(.A(new_n515), .B1(new_n524), .B2(new_n525), .ZN(G166));
  NAND3_X1  g101(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n527));
  XNOR2_X1  g102(.A(new_n527), .B(KEYINPUT7), .ZN(new_n528));
  XNOR2_X1  g103(.A(KEYINPUT69), .B(G51), .ZN(new_n529));
  OAI21_X1  g104(.A(new_n528), .B1(new_n520), .B2(new_n529), .ZN(new_n530));
  NAND2_X1  g105(.A1(new_n519), .A2(G89), .ZN(new_n531));
  NAND2_X1  g106(.A1(G63), .A2(G651), .ZN(new_n532));
  NAND2_X1  g107(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  AOI21_X1  g108(.A(new_n530), .B1(new_n511), .B2(new_n533), .ZN(G168));
  INV_X1    g109(.A(G52), .ZN(new_n535));
  INV_X1    g110(.A(G90), .ZN(new_n536));
  OAI22_X1  g111(.A1(new_n535), .A2(new_n520), .B1(new_n521), .B2(new_n536), .ZN(new_n537));
  AOI22_X1  g112(.A1(new_n511), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n538));
  NOR2_X1   g113(.A1(new_n538), .A2(new_n510), .ZN(new_n539));
  OR2_X1    g114(.A1(new_n537), .A2(new_n539), .ZN(G301));
  INV_X1    g115(.A(G301), .ZN(G171));
  INV_X1    g116(.A(G43), .ZN(new_n542));
  INV_X1    g117(.A(G81), .ZN(new_n543));
  OAI22_X1  g118(.A1(new_n542), .A2(new_n520), .B1(new_n521), .B2(new_n543), .ZN(new_n544));
  AOI22_X1  g119(.A1(new_n511), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n545));
  NOR2_X1   g120(.A1(new_n545), .A2(new_n510), .ZN(new_n546));
  NOR2_X1   g121(.A1(new_n544), .A2(new_n546), .ZN(new_n547));
  NAND2_X1  g122(.A1(new_n547), .A2(G860), .ZN(G153));
  NAND4_X1  g123(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g124(.A1(G1), .A2(G3), .ZN(new_n550));
  XNOR2_X1  g125(.A(new_n550), .B(KEYINPUT8), .ZN(new_n551));
  NAND4_X1  g126(.A1(G319), .A2(G483), .A3(G661), .A4(new_n551), .ZN(G188));
  NOR2_X1   g127(.A1(new_n517), .A2(new_n518), .ZN(new_n553));
  INV_X1    g128(.A(G543), .ZN(new_n554));
  NOR2_X1   g129(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n555), .A2(G53), .ZN(new_n556));
  XNOR2_X1  g131(.A(new_n556), .B(KEYINPUT9), .ZN(new_n557));
  INV_X1    g132(.A(new_n521), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n558), .A2(G91), .ZN(new_n559));
  AOI22_X1  g134(.A1(new_n511), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n560));
  OAI211_X1 g135(.A(new_n557), .B(new_n559), .C1(new_n510), .C2(new_n560), .ZN(G299));
  XNOR2_X1  g136(.A(G168), .B(KEYINPUT70), .ZN(new_n562));
  INV_X1    g137(.A(new_n562), .ZN(G286));
  INV_X1    g138(.A(G166), .ZN(G303));
  NAND2_X1  g139(.A1(new_n558), .A2(G87), .ZN(new_n565));
  OAI21_X1  g140(.A(G651), .B1(new_n511), .B2(G74), .ZN(new_n566));
  INV_X1    g141(.A(G49), .ZN(new_n567));
  OAI211_X1 g142(.A(new_n565), .B(new_n566), .C1(new_n567), .C2(new_n520), .ZN(G288));
  INV_X1    g143(.A(G48), .ZN(new_n569));
  INV_X1    g144(.A(G86), .ZN(new_n570));
  OAI22_X1  g145(.A1(new_n569), .A2(new_n520), .B1(new_n521), .B2(new_n570), .ZN(new_n571));
  AOI22_X1  g146(.A1(new_n511), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n572));
  NOR2_X1   g147(.A1(new_n572), .A2(new_n510), .ZN(new_n573));
  NOR2_X1   g148(.A1(new_n571), .A2(new_n573), .ZN(new_n574));
  INV_X1    g149(.A(new_n574), .ZN(G305));
  AOI22_X1  g150(.A1(new_n558), .A2(G85), .B1(new_n555), .B2(G47), .ZN(new_n576));
  AOI22_X1  g151(.A1(new_n511), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n577));
  OR2_X1    g152(.A1(new_n577), .A2(new_n510), .ZN(new_n578));
  NAND2_X1  g153(.A1(new_n576), .A2(new_n578), .ZN(G290));
  NAND2_X1  g154(.A1(G301), .A2(G868), .ZN(new_n580));
  XOR2_X1   g155(.A(new_n580), .B(KEYINPUT71), .Z(new_n581));
  NAND2_X1  g156(.A1(new_n555), .A2(G54), .ZN(new_n582));
  XOR2_X1   g157(.A(KEYINPUT72), .B(G66), .Z(new_n583));
  AOI22_X1  g158(.A1(new_n583), .A2(new_n511), .B1(G79), .B2(G543), .ZN(new_n584));
  OAI21_X1  g159(.A(new_n582), .B1(new_n584), .B2(new_n510), .ZN(new_n585));
  INV_X1    g160(.A(KEYINPUT73), .ZN(new_n586));
  XNOR2_X1  g161(.A(new_n585), .B(new_n586), .ZN(new_n587));
  INV_X1    g162(.A(G92), .ZN(new_n588));
  NOR2_X1   g163(.A1(new_n521), .A2(new_n588), .ZN(new_n589));
  XNOR2_X1  g164(.A(new_n589), .B(KEYINPUT10), .ZN(new_n590));
  AND2_X1   g165(.A1(new_n587), .A2(new_n590), .ZN(new_n591));
  OAI21_X1  g166(.A(new_n581), .B1(G868), .B2(new_n591), .ZN(G284));
  OAI21_X1  g167(.A(new_n581), .B1(G868), .B2(new_n591), .ZN(G321));
  NOR2_X1   g168(.A1(G299), .A2(G868), .ZN(new_n594));
  AOI21_X1  g169(.A(new_n594), .B1(G868), .B2(new_n562), .ZN(G297));
  AOI21_X1  g170(.A(new_n594), .B1(G868), .B2(new_n562), .ZN(G280));
  INV_X1    g171(.A(G559), .ZN(new_n597));
  OAI21_X1  g172(.A(new_n591), .B1(new_n597), .B2(G860), .ZN(G148));
  INV_X1    g173(.A(new_n547), .ZN(new_n599));
  INV_X1    g174(.A(G868), .ZN(new_n600));
  NAND2_X1  g175(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  NAND2_X1  g176(.A1(new_n587), .A2(new_n590), .ZN(new_n602));
  NOR2_X1   g177(.A1(new_n602), .A2(G559), .ZN(new_n603));
  XNOR2_X1  g178(.A(new_n603), .B(KEYINPUT74), .ZN(new_n604));
  OAI21_X1  g179(.A(new_n601), .B1(new_n604), .B2(new_n600), .ZN(new_n605));
  XOR2_X1   g180(.A(new_n605), .B(KEYINPUT75), .Z(G323));
  XNOR2_X1  g181(.A(G323), .B(KEYINPUT11), .ZN(G282));
  INV_X1    g182(.A(new_n466), .ZN(new_n608));
  NOR2_X1   g183(.A1(new_n470), .A2(new_n608), .ZN(new_n609));
  XOR2_X1   g184(.A(new_n609), .B(KEYINPUT12), .Z(new_n610));
  XOR2_X1   g185(.A(new_n610), .B(KEYINPUT13), .Z(new_n611));
  NAND2_X1  g186(.A1(new_n611), .A2(G2100), .ZN(new_n612));
  XNOR2_X1  g187(.A(new_n612), .B(KEYINPUT76), .ZN(new_n613));
  NAND2_X1  g188(.A1(new_n475), .A2(G123), .ZN(new_n614));
  NAND2_X1  g189(.A1(new_n478), .A2(G135), .ZN(new_n615));
  OR2_X1    g190(.A1(G99), .A2(G2105), .ZN(new_n616));
  OAI211_X1 g191(.A(new_n616), .B(G2104), .C1(G111), .C2(new_n458), .ZN(new_n617));
  NAND3_X1  g192(.A1(new_n614), .A2(new_n615), .A3(new_n617), .ZN(new_n618));
  XOR2_X1   g193(.A(new_n618), .B(G2096), .Z(new_n619));
  OAI211_X1 g194(.A(new_n613), .B(new_n619), .C1(G2100), .C2(new_n611), .ZN(G156));
  XNOR2_X1  g195(.A(G2427), .B(G2438), .ZN(new_n621));
  XNOR2_X1  g196(.A(new_n621), .B(G2430), .ZN(new_n622));
  XNOR2_X1  g197(.A(KEYINPUT15), .B(G2435), .ZN(new_n623));
  OR2_X1    g198(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  NAND2_X1  g199(.A1(new_n622), .A2(new_n623), .ZN(new_n625));
  NAND3_X1  g200(.A1(new_n624), .A2(KEYINPUT14), .A3(new_n625), .ZN(new_n626));
  XOR2_X1   g201(.A(KEYINPUT77), .B(KEYINPUT16), .Z(new_n627));
  XNOR2_X1  g202(.A(new_n626), .B(new_n627), .ZN(new_n628));
  XOR2_X1   g203(.A(G2451), .B(G2454), .Z(new_n629));
  XNOR2_X1  g204(.A(G2443), .B(G2446), .ZN(new_n630));
  XOR2_X1   g205(.A(new_n629), .B(new_n630), .Z(new_n631));
  XNOR2_X1  g206(.A(new_n628), .B(new_n631), .ZN(new_n632));
  XNOR2_X1  g207(.A(G1341), .B(G1348), .ZN(new_n633));
  NAND2_X1  g208(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  XOR2_X1   g209(.A(new_n634), .B(KEYINPUT78), .Z(new_n635));
  OAI21_X1  g210(.A(G14), .B1(new_n632), .B2(new_n633), .ZN(new_n636));
  NOR2_X1   g211(.A1(new_n635), .A2(new_n636), .ZN(G401));
  XOR2_X1   g212(.A(G2084), .B(G2090), .Z(new_n638));
  XNOR2_X1  g213(.A(G2067), .B(G2678), .ZN(new_n639));
  NAND2_X1  g214(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  XOR2_X1   g215(.A(G2072), .B(G2078), .Z(new_n641));
  NOR2_X1   g216(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  XNOR2_X1  g217(.A(new_n642), .B(KEYINPUT18), .ZN(new_n643));
  XNOR2_X1  g218(.A(new_n641), .B(KEYINPUT17), .ZN(new_n644));
  INV_X1    g219(.A(new_n638), .ZN(new_n645));
  INV_X1    g220(.A(new_n639), .ZN(new_n646));
  AOI21_X1  g221(.A(new_n644), .B1(new_n645), .B2(new_n646), .ZN(new_n647));
  NAND3_X1  g222(.A1(new_n645), .A2(new_n641), .A3(new_n646), .ZN(new_n648));
  NAND2_X1  g223(.A1(new_n648), .A2(new_n640), .ZN(new_n649));
  OAI21_X1  g224(.A(new_n643), .B1(new_n647), .B2(new_n649), .ZN(new_n650));
  XNOR2_X1  g225(.A(G2096), .B(G2100), .ZN(new_n651));
  XNOR2_X1  g226(.A(new_n651), .B(KEYINPUT79), .ZN(new_n652));
  XNOR2_X1  g227(.A(new_n650), .B(new_n652), .ZN(G227));
  XNOR2_X1  g228(.A(G1971), .B(G1976), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n654), .B(KEYINPUT81), .ZN(new_n655));
  XNOR2_X1  g230(.A(KEYINPUT80), .B(KEYINPUT19), .ZN(new_n656));
  XNOR2_X1  g231(.A(new_n655), .B(new_n656), .ZN(new_n657));
  XNOR2_X1  g232(.A(G1956), .B(G2474), .ZN(new_n658));
  XNOR2_X1  g233(.A(G1961), .B(G1966), .ZN(new_n659));
  NOR2_X1   g234(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  NAND2_X1  g235(.A1(new_n657), .A2(new_n660), .ZN(new_n661));
  XNOR2_X1  g236(.A(new_n661), .B(KEYINPUT20), .ZN(new_n662));
  AND2_X1   g237(.A1(new_n658), .A2(new_n659), .ZN(new_n663));
  NOR3_X1   g238(.A1(new_n657), .A2(new_n660), .A3(new_n663), .ZN(new_n664));
  AOI21_X1  g239(.A(new_n664), .B1(new_n657), .B2(new_n663), .ZN(new_n665));
  NAND2_X1  g240(.A1(new_n662), .A2(new_n665), .ZN(new_n666));
  XNOR2_X1  g241(.A(G1981), .B(G1986), .ZN(new_n667));
  XNOR2_X1  g242(.A(new_n666), .B(new_n667), .ZN(new_n668));
  XNOR2_X1  g243(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n669));
  XNOR2_X1  g244(.A(new_n668), .B(new_n669), .ZN(new_n670));
  XOR2_X1   g245(.A(G1991), .B(G1996), .Z(new_n671));
  XNOR2_X1  g246(.A(new_n671), .B(KEYINPUT83), .ZN(new_n672));
  XNOR2_X1  g247(.A(new_n672), .B(KEYINPUT82), .ZN(new_n673));
  XNOR2_X1  g248(.A(new_n670), .B(new_n673), .ZN(G229));
  XNOR2_X1  g249(.A(KEYINPUT90), .B(KEYINPUT28), .ZN(new_n675));
  INV_X1    g250(.A(G29), .ZN(new_n676));
  NAND2_X1  g251(.A1(new_n676), .A2(G26), .ZN(new_n677));
  XNOR2_X1  g252(.A(new_n675), .B(new_n677), .ZN(new_n678));
  NAND2_X1  g253(.A1(new_n478), .A2(G140), .ZN(new_n679));
  XNOR2_X1  g254(.A(new_n679), .B(KEYINPUT89), .ZN(new_n680));
  OAI21_X1  g255(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n681));
  INV_X1    g256(.A(G116), .ZN(new_n682));
  AOI21_X1  g257(.A(new_n681), .B1(new_n682), .B2(G2105), .ZN(new_n683));
  AOI21_X1  g258(.A(new_n683), .B1(new_n475), .B2(G128), .ZN(new_n684));
  NAND2_X1  g259(.A1(new_n680), .A2(new_n684), .ZN(new_n685));
  AOI21_X1  g260(.A(new_n678), .B1(new_n685), .B2(G29), .ZN(new_n686));
  XNOR2_X1  g261(.A(new_n686), .B(G2067), .ZN(new_n687));
  NAND2_X1  g262(.A1(new_n676), .A2(G27), .ZN(new_n688));
  OAI21_X1  g263(.A(new_n688), .B1(G164), .B2(new_n676), .ZN(new_n689));
  INV_X1    g264(.A(G2078), .ZN(new_n690));
  XNOR2_X1  g265(.A(new_n689), .B(new_n690), .ZN(new_n691));
  INV_X1    g266(.A(G2072), .ZN(new_n692));
  AND2_X1   g267(.A1(new_n676), .A2(G33), .ZN(new_n693));
  NAND3_X1  g268(.A1(new_n458), .A2(G103), .A3(G2104), .ZN(new_n694));
  XOR2_X1   g269(.A(new_n694), .B(KEYINPUT25), .Z(new_n695));
  INV_X1    g270(.A(G139), .ZN(new_n696));
  OAI21_X1  g271(.A(new_n695), .B1(new_n477), .B2(new_n696), .ZN(new_n697));
  XNOR2_X1  g272(.A(new_n697), .B(KEYINPUT91), .ZN(new_n698));
  NAND2_X1  g273(.A1(new_n498), .A2(new_n499), .ZN(new_n699));
  AOI22_X1  g274(.A1(new_n699), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n700));
  OAI21_X1  g275(.A(new_n698), .B1(new_n458), .B2(new_n700), .ZN(new_n701));
  AOI21_X1  g276(.A(new_n693), .B1(new_n701), .B2(G29), .ZN(new_n702));
  OAI211_X1 g277(.A(new_n687), .B(new_n691), .C1(new_n692), .C2(new_n702), .ZN(new_n703));
  NAND2_X1  g278(.A1(new_n475), .A2(G129), .ZN(new_n704));
  INV_X1    g279(.A(KEYINPUT94), .ZN(new_n705));
  XNOR2_X1  g280(.A(new_n704), .B(new_n705), .ZN(new_n706));
  NAND3_X1  g281(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n707));
  XOR2_X1   g282(.A(new_n707), .B(KEYINPUT26), .Z(new_n708));
  INV_X1    g283(.A(G105), .ZN(new_n709));
  OAI21_X1  g284(.A(new_n708), .B1(new_n709), .B2(new_n608), .ZN(new_n710));
  AOI21_X1  g285(.A(new_n710), .B1(new_n478), .B2(G141), .ZN(new_n711));
  NAND2_X1  g286(.A1(new_n706), .A2(new_n711), .ZN(new_n712));
  INV_X1    g287(.A(new_n712), .ZN(new_n713));
  NAND2_X1  g288(.A1(new_n713), .A2(G29), .ZN(new_n714));
  INV_X1    g289(.A(KEYINPUT95), .ZN(new_n715));
  OAI21_X1  g290(.A(new_n715), .B1(G29), .B2(G32), .ZN(new_n716));
  NAND2_X1  g291(.A1(new_n714), .A2(new_n716), .ZN(new_n717));
  OAI21_X1  g292(.A(new_n717), .B1(KEYINPUT95), .B2(new_n714), .ZN(new_n718));
  XOR2_X1   g293(.A(KEYINPUT27), .B(G1996), .Z(new_n719));
  XOR2_X1   g294(.A(new_n719), .B(KEYINPUT96), .Z(new_n720));
  XNOR2_X1  g295(.A(new_n718), .B(new_n720), .ZN(new_n721));
  INV_X1    g296(.A(G16), .ZN(new_n722));
  NAND2_X1  g297(.A1(new_n722), .A2(G20), .ZN(new_n723));
  XOR2_X1   g298(.A(new_n723), .B(KEYINPUT23), .Z(new_n724));
  AOI21_X1  g299(.A(new_n724), .B1(G299), .B2(G16), .ZN(new_n725));
  XNOR2_X1  g300(.A(new_n725), .B(KEYINPUT98), .ZN(new_n726));
  INV_X1    g301(.A(G1956), .ZN(new_n727));
  XNOR2_X1  g302(.A(new_n726), .B(new_n727), .ZN(new_n728));
  NOR2_X1   g303(.A1(G171), .A2(new_n722), .ZN(new_n729));
  AOI21_X1  g304(.A(new_n729), .B1(G5), .B2(new_n722), .ZN(new_n730));
  INV_X1    g305(.A(G1961), .ZN(new_n731));
  NAND2_X1  g306(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  XOR2_X1   g307(.A(KEYINPUT30), .B(G28), .Z(new_n733));
  NOR2_X1   g308(.A1(KEYINPUT31), .A2(G11), .ZN(new_n734));
  AND2_X1   g309(.A1(KEYINPUT31), .A2(G11), .ZN(new_n735));
  OAI221_X1 g310(.A(new_n732), .B1(G29), .B2(new_n733), .C1(new_n734), .C2(new_n735), .ZN(new_n736));
  XOR2_X1   g311(.A(KEYINPUT92), .B(KEYINPUT24), .Z(new_n737));
  INV_X1    g312(.A(G34), .ZN(new_n738));
  OAI21_X1  g313(.A(new_n676), .B1(new_n737), .B2(new_n738), .ZN(new_n739));
  AOI21_X1  g314(.A(new_n739), .B1(new_n738), .B2(new_n737), .ZN(new_n740));
  XOR2_X1   g315(.A(new_n740), .B(KEYINPUT93), .Z(new_n741));
  AOI21_X1  g316(.A(new_n741), .B1(G29), .B2(G160), .ZN(new_n742));
  OR2_X1    g317(.A1(new_n742), .A2(G2084), .ZN(new_n743));
  NOR2_X1   g318(.A1(G168), .A2(new_n722), .ZN(new_n744));
  AOI21_X1  g319(.A(new_n744), .B1(new_n722), .B2(G21), .ZN(new_n745));
  INV_X1    g320(.A(G1966), .ZN(new_n746));
  NAND2_X1  g321(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  NAND2_X1  g322(.A1(new_n742), .A2(G2084), .ZN(new_n748));
  OR2_X1    g323(.A1(new_n618), .A2(new_n676), .ZN(new_n749));
  NAND4_X1  g324(.A1(new_n743), .A2(new_n747), .A3(new_n748), .A4(new_n749), .ZN(new_n750));
  XNOR2_X1  g325(.A(KEYINPUT88), .B(G1341), .ZN(new_n751));
  NAND2_X1  g326(.A1(new_n722), .A2(G19), .ZN(new_n752));
  XNOR2_X1  g327(.A(new_n752), .B(KEYINPUT87), .ZN(new_n753));
  AOI21_X1  g328(.A(new_n753), .B1(new_n599), .B2(G16), .ZN(new_n754));
  OAI22_X1  g329(.A1(new_n730), .A2(new_n731), .B1(new_n751), .B2(new_n754), .ZN(new_n755));
  NAND2_X1  g330(.A1(new_n754), .A2(new_n751), .ZN(new_n756));
  OAI21_X1  g331(.A(new_n756), .B1(new_n745), .B2(new_n746), .ZN(new_n757));
  NOR4_X1   g332(.A1(new_n736), .A2(new_n750), .A3(new_n755), .A4(new_n757), .ZN(new_n758));
  NOR2_X1   g333(.A1(G4), .A2(G16), .ZN(new_n759));
  XNOR2_X1  g334(.A(new_n759), .B(KEYINPUT86), .ZN(new_n760));
  OAI21_X1  g335(.A(new_n760), .B1(new_n602), .B2(new_n722), .ZN(new_n761));
  INV_X1    g336(.A(G1348), .ZN(new_n762));
  XNOR2_X1  g337(.A(new_n761), .B(new_n762), .ZN(new_n763));
  AOI21_X1  g338(.A(new_n763), .B1(new_n692), .B2(new_n702), .ZN(new_n764));
  NAND4_X1  g339(.A1(new_n721), .A2(new_n728), .A3(new_n758), .A4(new_n764), .ZN(new_n765));
  INV_X1    g340(.A(G2090), .ZN(new_n766));
  NAND2_X1  g341(.A1(new_n676), .A2(G35), .ZN(new_n767));
  OAI21_X1  g342(.A(new_n767), .B1(G162), .B2(new_n676), .ZN(new_n768));
  XOR2_X1   g343(.A(new_n768), .B(KEYINPUT29), .Z(new_n769));
  AOI211_X1 g344(.A(new_n703), .B(new_n765), .C1(new_n766), .C2(new_n769), .ZN(new_n770));
  NOR2_X1   g345(.A1(G6), .A2(G16), .ZN(new_n771));
  AOI21_X1  g346(.A(new_n771), .B1(new_n574), .B2(G16), .ZN(new_n772));
  XOR2_X1   g347(.A(new_n772), .B(KEYINPUT85), .Z(new_n773));
  XNOR2_X1  g348(.A(KEYINPUT32), .B(G1981), .ZN(new_n774));
  INV_X1    g349(.A(new_n774), .ZN(new_n775));
  NOR2_X1   g350(.A1(new_n773), .A2(new_n775), .ZN(new_n776));
  NAND2_X1  g351(.A1(new_n722), .A2(G23), .ZN(new_n777));
  INV_X1    g352(.A(G288), .ZN(new_n778));
  OAI21_X1  g353(.A(new_n777), .B1(new_n778), .B2(new_n722), .ZN(new_n779));
  XOR2_X1   g354(.A(KEYINPUT33), .B(G1976), .Z(new_n780));
  XNOR2_X1  g355(.A(new_n779), .B(new_n780), .ZN(new_n781));
  NOR2_X1   g356(.A1(new_n776), .A2(new_n781), .ZN(new_n782));
  NAND2_X1  g357(.A1(G166), .A2(G16), .ZN(new_n783));
  OAI21_X1  g358(.A(new_n783), .B1(G16), .B2(G22), .ZN(new_n784));
  INV_X1    g359(.A(G1971), .ZN(new_n785));
  AOI22_X1  g360(.A1(new_n773), .A2(new_n775), .B1(new_n784), .B2(new_n785), .ZN(new_n786));
  OAI211_X1 g361(.A(new_n782), .B(new_n786), .C1(new_n785), .C2(new_n784), .ZN(new_n787));
  OR2_X1    g362(.A1(new_n787), .A2(KEYINPUT34), .ZN(new_n788));
  NAND2_X1  g363(.A1(new_n787), .A2(KEYINPUT34), .ZN(new_n789));
  NAND2_X1  g364(.A1(new_n475), .A2(G119), .ZN(new_n790));
  NAND2_X1  g365(.A1(new_n478), .A2(G131), .ZN(new_n791));
  OAI21_X1  g366(.A(KEYINPUT84), .B1(G95), .B2(G2105), .ZN(new_n792));
  INV_X1    g367(.A(new_n792), .ZN(new_n793));
  NOR3_X1   g368(.A1(KEYINPUT84), .A2(G95), .A3(G2105), .ZN(new_n794));
  OAI221_X1 g369(.A(G2104), .B1(G107), .B2(new_n458), .C1(new_n793), .C2(new_n794), .ZN(new_n795));
  NAND3_X1  g370(.A1(new_n790), .A2(new_n791), .A3(new_n795), .ZN(new_n796));
  INV_X1    g371(.A(new_n796), .ZN(new_n797));
  NAND2_X1  g372(.A1(new_n797), .A2(G29), .ZN(new_n798));
  OAI21_X1  g373(.A(new_n798), .B1(G25), .B2(G29), .ZN(new_n799));
  XOR2_X1   g374(.A(KEYINPUT35), .B(G1991), .Z(new_n800));
  AND2_X1   g375(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  NOR2_X1   g376(.A1(new_n799), .A2(new_n800), .ZN(new_n802));
  NAND2_X1  g377(.A1(new_n722), .A2(G24), .ZN(new_n803));
  INV_X1    g378(.A(G290), .ZN(new_n804));
  OAI21_X1  g379(.A(new_n803), .B1(new_n804), .B2(new_n722), .ZN(new_n805));
  XNOR2_X1  g380(.A(new_n805), .B(G1986), .ZN(new_n806));
  NOR3_X1   g381(.A1(new_n801), .A2(new_n802), .A3(new_n806), .ZN(new_n807));
  NAND3_X1  g382(.A1(new_n788), .A2(new_n789), .A3(new_n807), .ZN(new_n808));
  XNOR2_X1  g383(.A(new_n808), .B(KEYINPUT36), .ZN(new_n809));
  NOR2_X1   g384(.A1(new_n769), .A2(new_n766), .ZN(new_n810));
  XNOR2_X1  g385(.A(new_n810), .B(KEYINPUT97), .ZN(new_n811));
  NAND3_X1  g386(.A1(new_n770), .A2(new_n809), .A3(new_n811), .ZN(G150));
  INV_X1    g387(.A(G150), .ZN(G311));
  INV_X1    g388(.A(G55), .ZN(new_n814));
  INV_X1    g389(.A(G93), .ZN(new_n815));
  OAI22_X1  g390(.A1(new_n814), .A2(new_n520), .B1(new_n521), .B2(new_n815), .ZN(new_n816));
  AOI22_X1  g391(.A1(new_n511), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n817));
  NOR2_X1   g392(.A1(new_n817), .A2(new_n510), .ZN(new_n818));
  NOR2_X1   g393(.A1(new_n816), .A2(new_n818), .ZN(new_n819));
  XNOR2_X1  g394(.A(KEYINPUT100), .B(G860), .ZN(new_n820));
  NOR2_X1   g395(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  XNOR2_X1  g396(.A(new_n821), .B(KEYINPUT37), .ZN(new_n822));
  NOR2_X1   g397(.A1(new_n602), .A2(new_n597), .ZN(new_n823));
  XNOR2_X1  g398(.A(new_n823), .B(KEYINPUT99), .ZN(new_n824));
  XNOR2_X1  g399(.A(new_n824), .B(KEYINPUT38), .ZN(new_n825));
  XOR2_X1   g400(.A(new_n547), .B(new_n819), .Z(new_n826));
  XNOR2_X1  g401(.A(new_n825), .B(new_n826), .ZN(new_n827));
  NAND2_X1  g402(.A1(new_n827), .A2(KEYINPUT39), .ZN(new_n828));
  XOR2_X1   g403(.A(new_n828), .B(KEYINPUT101), .Z(new_n829));
  OAI21_X1  g404(.A(new_n820), .B1(new_n827), .B2(KEYINPUT39), .ZN(new_n830));
  OAI21_X1  g405(.A(new_n822), .B1(new_n829), .B2(new_n830), .ZN(G145));
  INV_X1    g406(.A(KEYINPUT40), .ZN(new_n832));
  XNOR2_X1  g407(.A(new_n712), .B(new_n701), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n475), .A2(G130), .ZN(new_n834));
  NAND2_X1  g409(.A1(new_n478), .A2(G142), .ZN(new_n835));
  NOR3_X1   g410(.A1(new_n458), .A2(KEYINPUT104), .A3(G118), .ZN(new_n836));
  OAI21_X1  g411(.A(KEYINPUT104), .B1(new_n458), .B2(G118), .ZN(new_n837));
  OR2_X1    g412(.A1(G106), .A2(G2105), .ZN(new_n838));
  NAND3_X1  g413(.A1(new_n837), .A2(G2104), .A3(new_n838), .ZN(new_n839));
  OAI211_X1 g414(.A(new_n834), .B(new_n835), .C1(new_n836), .C2(new_n839), .ZN(new_n840));
  XOR2_X1   g415(.A(new_n840), .B(new_n610), .Z(new_n841));
  XNOR2_X1  g416(.A(new_n833), .B(new_n841), .ZN(new_n842));
  NAND3_X1  g417(.A1(new_n502), .A2(new_n506), .A3(new_n495), .ZN(new_n843));
  XNOR2_X1  g418(.A(new_n685), .B(new_n843), .ZN(new_n844));
  XNOR2_X1  g419(.A(new_n844), .B(new_n796), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n842), .A2(new_n845), .ZN(new_n846));
  OR2_X1    g421(.A1(new_n842), .A2(new_n845), .ZN(new_n847));
  XNOR2_X1  g422(.A(G162), .B(new_n618), .ZN(new_n848));
  INV_X1    g423(.A(G160), .ZN(new_n849));
  OR2_X1    g424(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  XNOR2_X1  g425(.A(KEYINPUT102), .B(KEYINPUT103), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n848), .A2(new_n849), .ZN(new_n852));
  NAND3_X1  g427(.A1(new_n850), .A2(new_n851), .A3(new_n852), .ZN(new_n853));
  INV_X1    g428(.A(new_n853), .ZN(new_n854));
  AOI21_X1  g429(.A(new_n851), .B1(new_n850), .B2(new_n852), .ZN(new_n855));
  OAI211_X1 g430(.A(new_n846), .B(new_n847), .C1(new_n854), .C2(new_n855), .ZN(new_n856));
  INV_X1    g431(.A(G37), .ZN(new_n857));
  NAND2_X1  g432(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  INV_X1    g433(.A(new_n855), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n859), .A2(new_n853), .ZN(new_n860));
  AND2_X1   g435(.A1(new_n847), .A2(new_n846), .ZN(new_n861));
  NOR2_X1   g436(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  OAI21_X1  g437(.A(new_n832), .B1(new_n858), .B2(new_n862), .ZN(new_n863));
  OR2_X1    g438(.A1(new_n860), .A2(new_n861), .ZN(new_n864));
  AOI21_X1  g439(.A(G37), .B1(new_n860), .B2(new_n861), .ZN(new_n865));
  NAND3_X1  g440(.A1(new_n864), .A2(new_n865), .A3(KEYINPUT40), .ZN(new_n866));
  AND2_X1   g441(.A1(new_n863), .A2(new_n866), .ZN(G395));
  OAI21_X1  g442(.A(new_n600), .B1(new_n816), .B2(new_n818), .ZN(new_n868));
  INV_X1    g443(.A(new_n826), .ZN(new_n869));
  XNOR2_X1  g444(.A(new_n604), .B(new_n869), .ZN(new_n870));
  XNOR2_X1  g445(.A(new_n591), .B(G299), .ZN(new_n871));
  XNOR2_X1  g446(.A(new_n871), .B(KEYINPUT41), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n870), .A2(new_n872), .ZN(new_n873));
  OAI21_X1  g448(.A(new_n873), .B1(new_n871), .B2(new_n870), .ZN(new_n874));
  XNOR2_X1  g449(.A(G288), .B(G290), .ZN(new_n875));
  INV_X1    g450(.A(KEYINPUT105), .ZN(new_n876));
  AND2_X1   g451(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  XNOR2_X1  g452(.A(G166), .B(G305), .ZN(new_n878));
  NOR2_X1   g453(.A1(new_n875), .A2(new_n876), .ZN(new_n879));
  OR3_X1    g454(.A1(new_n877), .A2(new_n878), .A3(new_n879), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n877), .A2(new_n878), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  XNOR2_X1  g457(.A(new_n882), .B(KEYINPUT42), .ZN(new_n883));
  XNOR2_X1  g458(.A(new_n874), .B(new_n883), .ZN(new_n884));
  OAI21_X1  g459(.A(new_n868), .B1(new_n884), .B2(new_n600), .ZN(G295));
  OAI21_X1  g460(.A(new_n868), .B1(new_n884), .B2(new_n600), .ZN(G331));
  NOR2_X1   g461(.A1(G171), .A2(G168), .ZN(new_n887));
  AOI21_X1  g462(.A(new_n887), .B1(new_n562), .B2(G171), .ZN(new_n888));
  XNOR2_X1  g463(.A(new_n888), .B(new_n869), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n889), .A2(new_n871), .ZN(new_n890));
  OAI21_X1  g465(.A(new_n890), .B1(new_n872), .B2(new_n889), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n891), .A2(new_n882), .ZN(new_n892));
  INV_X1    g467(.A(new_n882), .ZN(new_n893));
  OAI211_X1 g468(.A(new_n893), .B(new_n890), .C1(new_n872), .C2(new_n889), .ZN(new_n894));
  XNOR2_X1  g469(.A(KEYINPUT106), .B(KEYINPUT43), .ZN(new_n895));
  NAND4_X1  g470(.A1(new_n892), .A2(new_n894), .A3(new_n857), .A4(new_n895), .ZN(new_n896));
  INV_X1    g471(.A(KEYINPUT108), .ZN(new_n897));
  OR2_X1    g472(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n896), .A2(new_n897), .ZN(new_n899));
  INV_X1    g474(.A(KEYINPUT44), .ZN(new_n900));
  NAND3_X1  g475(.A1(new_n892), .A2(new_n894), .A3(new_n857), .ZN(new_n901));
  AOI21_X1  g476(.A(new_n900), .B1(new_n901), .B2(KEYINPUT43), .ZN(new_n902));
  NAND3_X1  g477(.A1(new_n898), .A2(new_n899), .A3(new_n902), .ZN(new_n903));
  INV_X1    g478(.A(KEYINPUT107), .ZN(new_n904));
  INV_X1    g479(.A(new_n895), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n901), .A2(new_n905), .ZN(new_n906));
  NAND2_X1  g481(.A1(new_n906), .A2(new_n896), .ZN(new_n907));
  AOI21_X1  g482(.A(new_n904), .B1(new_n907), .B2(new_n900), .ZN(new_n908));
  AOI211_X1 g483(.A(KEYINPUT107), .B(KEYINPUT44), .C1(new_n906), .C2(new_n896), .ZN(new_n909));
  OAI21_X1  g484(.A(new_n903), .B1(new_n908), .B2(new_n909), .ZN(G397));
  INV_X1    g485(.A(G1384), .ZN(new_n911));
  AOI21_X1  g486(.A(KEYINPUT45), .B1(new_n843), .B2(new_n911), .ZN(new_n912));
  INV_X1    g487(.A(new_n912), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n461), .A2(new_n462), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n914), .A2(G2105), .ZN(new_n915));
  AND2_X1   g490(.A1(new_n464), .A2(new_n467), .ZN(new_n916));
  NAND3_X1  g491(.A1(new_n915), .A2(new_n916), .A3(G40), .ZN(new_n917));
  INV_X1    g492(.A(KEYINPUT109), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  NAND3_X1  g494(.A1(G160), .A2(KEYINPUT109), .A3(G40), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  NOR2_X1   g496(.A1(new_n913), .A2(new_n921), .ZN(new_n922));
  INV_X1    g497(.A(G1996), .ZN(new_n923));
  XNOR2_X1  g498(.A(new_n712), .B(new_n923), .ZN(new_n924));
  INV_X1    g499(.A(G2067), .ZN(new_n925));
  XNOR2_X1  g500(.A(new_n685), .B(new_n925), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n797), .A2(new_n800), .ZN(new_n927));
  OR2_X1    g502(.A1(new_n797), .A2(new_n800), .ZN(new_n928));
  NAND4_X1  g503(.A1(new_n924), .A2(new_n926), .A3(new_n927), .A4(new_n928), .ZN(new_n929));
  INV_X1    g504(.A(G1986), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n804), .A2(new_n930), .ZN(new_n931));
  XOR2_X1   g506(.A(new_n931), .B(KEYINPUT110), .Z(new_n932));
  INV_X1    g507(.A(new_n932), .ZN(new_n933));
  OAI21_X1  g508(.A(new_n933), .B1(new_n930), .B2(new_n804), .ZN(new_n934));
  OAI21_X1  g509(.A(new_n922), .B1(new_n929), .B2(new_n934), .ZN(new_n935));
  INV_X1    g510(.A(KEYINPUT54), .ZN(new_n936));
  INV_X1    g511(.A(new_n921), .ZN(new_n937));
  NAND3_X1  g512(.A1(new_n843), .A2(KEYINPUT45), .A3(new_n911), .ZN(new_n938));
  INV_X1    g513(.A(KEYINPUT111), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  OAI21_X1  g515(.A(new_n911), .B1(new_n496), .B2(new_n508), .ZN(new_n941));
  INV_X1    g516(.A(KEYINPUT45), .ZN(new_n942));
  AOI21_X1  g517(.A(new_n940), .B1(new_n941), .B2(new_n942), .ZN(new_n943));
  INV_X1    g518(.A(KEYINPUT66), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n843), .A2(new_n944), .ZN(new_n945));
  AOI21_X1  g520(.A(G1384), .B1(new_n945), .B2(new_n507), .ZN(new_n946));
  NOR3_X1   g521(.A1(new_n946), .A2(new_n939), .A3(KEYINPUT45), .ZN(new_n947));
  OAI21_X1  g522(.A(new_n937), .B1(new_n943), .B2(new_n947), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n948), .A2(KEYINPUT112), .ZN(new_n949));
  OAI211_X1 g524(.A(new_n939), .B(new_n938), .C1(new_n946), .C2(KEYINPUT45), .ZN(new_n950));
  NAND3_X1  g525(.A1(new_n941), .A2(KEYINPUT111), .A3(new_n942), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n950), .A2(new_n951), .ZN(new_n952));
  INV_X1    g527(.A(KEYINPUT112), .ZN(new_n953));
  NAND3_X1  g528(.A1(new_n952), .A2(new_n953), .A3(new_n937), .ZN(new_n954));
  AOI21_X1  g529(.A(G2078), .B1(new_n949), .B2(new_n954), .ZN(new_n955));
  OAI21_X1  g530(.A(KEYINPUT125), .B1(new_n955), .B2(KEYINPUT53), .ZN(new_n956));
  AOI21_X1  g531(.A(new_n953), .B1(new_n952), .B2(new_n937), .ZN(new_n957));
  AOI211_X1 g532(.A(KEYINPUT112), .B(new_n921), .C1(new_n950), .C2(new_n951), .ZN(new_n958));
  OAI21_X1  g533(.A(new_n690), .B1(new_n957), .B2(new_n958), .ZN(new_n959));
  INV_X1    g534(.A(KEYINPUT125), .ZN(new_n960));
  INV_X1    g535(.A(KEYINPUT53), .ZN(new_n961));
  NAND3_X1  g536(.A1(new_n959), .A2(new_n960), .A3(new_n961), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n956), .A2(new_n962), .ZN(new_n963));
  NAND3_X1  g538(.A1(new_n937), .A2(KEYINPUT116), .A3(new_n913), .ZN(new_n964));
  INV_X1    g539(.A(KEYINPUT116), .ZN(new_n965));
  OAI21_X1  g540(.A(new_n965), .B1(new_n921), .B2(new_n912), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n946), .A2(KEYINPUT45), .ZN(new_n967));
  NAND3_X1  g542(.A1(new_n964), .A2(new_n966), .A3(new_n967), .ZN(new_n968));
  NOR3_X1   g543(.A1(new_n968), .A2(new_n961), .A3(G2078), .ZN(new_n969));
  INV_X1    g544(.A(KEYINPUT50), .ZN(new_n970));
  NAND3_X1  g545(.A1(new_n843), .A2(new_n970), .A3(new_n911), .ZN(new_n971));
  OAI211_X1 g546(.A(new_n937), .B(new_n971), .C1(new_n946), .C2(new_n970), .ZN(new_n972));
  AOI21_X1  g547(.A(new_n969), .B1(new_n731), .B2(new_n972), .ZN(new_n973));
  AOI21_X1  g548(.A(G301), .B1(new_n963), .B2(new_n973), .ZN(new_n974));
  NOR3_X1   g549(.A1(new_n917), .A2(new_n961), .A3(G2078), .ZN(new_n975));
  NAND3_X1  g550(.A1(new_n913), .A2(new_n938), .A3(new_n975), .ZN(new_n976));
  NAND3_X1  g551(.A1(new_n971), .A2(new_n919), .A3(new_n920), .ZN(new_n977));
  AOI21_X1  g552(.A(new_n977), .B1(new_n941), .B2(KEYINPUT50), .ZN(new_n978));
  OAI21_X1  g553(.A(new_n976), .B1(new_n978), .B2(G1961), .ZN(new_n979));
  AOI211_X1 g554(.A(G171), .B(new_n979), .C1(new_n956), .C2(new_n962), .ZN(new_n980));
  OAI21_X1  g555(.A(new_n936), .B1(new_n974), .B2(new_n980), .ZN(new_n981));
  XNOR2_X1  g556(.A(KEYINPUT56), .B(G2072), .ZN(new_n982));
  OAI211_X1 g557(.A(new_n937), .B(new_n982), .C1(new_n943), .C2(new_n947), .ZN(new_n983));
  AOI21_X1  g558(.A(KEYINPUT57), .B1(new_n557), .B2(KEYINPUT117), .ZN(new_n984));
  XNOR2_X1  g559(.A(G299), .B(new_n984), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n843), .A2(new_n911), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n986), .A2(KEYINPUT50), .ZN(new_n987));
  OAI211_X1 g562(.A(new_n937), .B(new_n987), .C1(new_n941), .C2(KEYINPUT50), .ZN(new_n988));
  NAND2_X1  g563(.A1(new_n988), .A2(new_n727), .ZN(new_n989));
  NAND3_X1  g564(.A1(new_n983), .A2(new_n985), .A3(new_n989), .ZN(new_n990));
  INV_X1    g565(.A(KEYINPUT118), .ZN(new_n991));
  NOR3_X1   g566(.A1(new_n921), .A2(G2067), .A3(new_n986), .ZN(new_n992));
  AOI211_X1 g567(.A(new_n991), .B(new_n992), .C1(new_n972), .C2(new_n762), .ZN(new_n993));
  NOR2_X1   g568(.A1(new_n946), .A2(new_n970), .ZN(new_n994));
  OAI21_X1  g569(.A(new_n762), .B1(new_n994), .B2(new_n977), .ZN(new_n995));
  INV_X1    g570(.A(new_n992), .ZN(new_n996));
  AOI21_X1  g571(.A(KEYINPUT118), .B1(new_n995), .B2(new_n996), .ZN(new_n997));
  NOR3_X1   g572(.A1(new_n993), .A2(new_n997), .A3(new_n602), .ZN(new_n998));
  AOI21_X1  g573(.A(new_n985), .B1(new_n983), .B2(new_n989), .ZN(new_n999));
  OAI21_X1  g574(.A(new_n990), .B1(new_n998), .B2(new_n999), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n983), .A2(new_n989), .ZN(new_n1001));
  INV_X1    g576(.A(new_n985), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n1001), .A2(new_n1002), .ZN(new_n1003));
  NAND3_X1  g578(.A1(new_n1003), .A2(KEYINPUT121), .A3(new_n990), .ZN(new_n1004));
  INV_X1    g579(.A(KEYINPUT121), .ZN(new_n1005));
  AOI21_X1  g580(.A(KEYINPUT61), .B1(new_n999), .B2(new_n1005), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n1004), .A2(new_n1006), .ZN(new_n1007));
  XNOR2_X1  g582(.A(new_n591), .B(KEYINPUT123), .ZN(new_n1008));
  OAI211_X1 g583(.A(KEYINPUT60), .B(new_n1008), .C1(new_n993), .C2(new_n997), .ZN(new_n1009));
  OAI21_X1  g584(.A(new_n996), .B1(new_n978), .B2(G1348), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n1010), .A2(new_n991), .ZN(new_n1011));
  INV_X1    g586(.A(KEYINPUT60), .ZN(new_n1012));
  NAND3_X1  g587(.A1(new_n995), .A2(KEYINPUT118), .A3(new_n996), .ZN(new_n1013));
  NAND3_X1  g588(.A1(new_n1011), .A2(new_n1012), .A3(new_n1013), .ZN(new_n1014));
  AOI21_X1  g589(.A(new_n1012), .B1(new_n1011), .B2(new_n1013), .ZN(new_n1015));
  NAND2_X1  g590(.A1(new_n602), .A2(KEYINPUT123), .ZN(new_n1016));
  OAI211_X1 g591(.A(new_n1009), .B(new_n1014), .C1(new_n1015), .C2(new_n1016), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n937), .A2(new_n923), .ZN(new_n1018));
  AOI21_X1  g593(.A(new_n1018), .B1(new_n950), .B2(new_n951), .ZN(new_n1019));
  INV_X1    g594(.A(KEYINPUT119), .ZN(new_n1020));
  NOR2_X1   g595(.A1(new_n921), .A2(new_n986), .ZN(new_n1021));
  XNOR2_X1  g596(.A(KEYINPUT58), .B(G1341), .ZN(new_n1022));
  NOR2_X1   g597(.A1(new_n1021), .A2(new_n1022), .ZN(new_n1023));
  OR3_X1    g598(.A1(new_n1019), .A2(new_n1020), .A3(new_n1023), .ZN(new_n1024));
  OAI21_X1  g599(.A(new_n1020), .B1(new_n1019), .B2(new_n1023), .ZN(new_n1025));
  AND2_X1   g600(.A1(KEYINPUT120), .A2(KEYINPUT59), .ZN(new_n1026));
  NAND4_X1  g601(.A1(new_n1024), .A2(new_n547), .A3(new_n1025), .A4(new_n1026), .ZN(new_n1027));
  NAND3_X1  g602(.A1(new_n1024), .A2(new_n547), .A3(new_n1025), .ZN(new_n1028));
  NOR2_X1   g603(.A1(KEYINPUT120), .A2(KEYINPUT59), .ZN(new_n1029));
  NOR2_X1   g604(.A1(new_n1026), .A2(new_n1029), .ZN(new_n1030));
  NAND2_X1  g605(.A1(new_n1028), .A2(new_n1030), .ZN(new_n1031));
  NAND4_X1  g606(.A1(new_n1007), .A2(new_n1017), .A3(new_n1027), .A4(new_n1031), .ZN(new_n1032));
  NAND3_X1  g607(.A1(new_n1003), .A2(KEYINPUT61), .A3(new_n990), .ZN(new_n1033));
  INV_X1    g608(.A(KEYINPUT122), .ZN(new_n1034));
  XNOR2_X1  g609(.A(new_n1033), .B(new_n1034), .ZN(new_n1035));
  OAI21_X1  g610(.A(new_n1000), .B1(new_n1032), .B2(new_n1035), .ZN(new_n1036));
  AND2_X1   g611(.A1(new_n973), .A2(G301), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n963), .A2(new_n1037), .ZN(new_n1038));
  AOI21_X1  g613(.A(new_n979), .B1(new_n956), .B2(new_n962), .ZN(new_n1039));
  OAI211_X1 g614(.A(new_n1038), .B(KEYINPUT54), .C1(G301), .C2(new_n1039), .ZN(new_n1040));
  NAND2_X1  g615(.A1(G305), .A2(G1981), .ZN(new_n1041));
  OR3_X1    g616(.A1(new_n571), .A2(G1981), .A3(new_n573), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n1041), .A2(new_n1042), .ZN(new_n1043));
  XNOR2_X1  g618(.A(new_n1043), .B(KEYINPUT49), .ZN(new_n1044));
  INV_X1    g619(.A(G8), .ZN(new_n1045));
  NOR2_X1   g620(.A1(new_n1021), .A2(new_n1045), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n1044), .A2(new_n1046), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n778), .A2(G1976), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n1046), .A2(new_n1048), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n1049), .A2(KEYINPUT52), .ZN(new_n1050));
  INV_X1    g625(.A(G1976), .ZN(new_n1051));
  AOI21_X1  g626(.A(KEYINPUT52), .B1(G288), .B2(new_n1051), .ZN(new_n1052));
  NAND3_X1  g627(.A1(new_n1046), .A2(new_n1048), .A3(new_n1052), .ZN(new_n1053));
  AND2_X1   g628(.A1(new_n1053), .A2(KEYINPUT114), .ZN(new_n1054));
  NOR2_X1   g629(.A1(new_n1053), .A2(KEYINPUT114), .ZN(new_n1055));
  OAI211_X1 g630(.A(new_n1047), .B(new_n1050), .C1(new_n1054), .C2(new_n1055), .ZN(new_n1056));
  NAND3_X1  g631(.A1(new_n949), .A2(new_n785), .A3(new_n954), .ZN(new_n1057));
  NAND2_X1  g632(.A1(new_n978), .A2(new_n766), .ZN(new_n1058));
  AOI21_X1  g633(.A(new_n1045), .B1(new_n1057), .B2(new_n1058), .ZN(new_n1059));
  NOR2_X1   g634(.A1(G166), .A2(new_n1045), .ZN(new_n1060));
  NAND3_X1  g635(.A1(new_n1060), .A2(KEYINPUT113), .A3(KEYINPUT55), .ZN(new_n1061));
  OAI21_X1  g636(.A(new_n1061), .B1(KEYINPUT55), .B2(new_n1060), .ZN(new_n1062));
  AOI21_X1  g637(.A(KEYINPUT113), .B1(new_n1060), .B2(KEYINPUT55), .ZN(new_n1063));
  NOR2_X1   g638(.A1(new_n1062), .A2(new_n1063), .ZN(new_n1064));
  INV_X1    g639(.A(new_n1064), .ZN(new_n1065));
  AOI21_X1  g640(.A(new_n1056), .B1(new_n1059), .B2(new_n1065), .ZN(new_n1066));
  INV_X1    g641(.A(G2084), .ZN(new_n1067));
  AOI22_X1  g642(.A1(new_n968), .A2(new_n746), .B1(new_n1067), .B2(new_n978), .ZN(new_n1068));
  OR3_X1    g643(.A1(new_n1068), .A2(new_n1045), .A3(G168), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n1068), .A2(G168), .ZN(new_n1070));
  NOR2_X1   g645(.A1(new_n1045), .A2(KEYINPUT124), .ZN(new_n1071));
  AOI21_X1  g646(.A(KEYINPUT51), .B1(new_n1070), .B2(new_n1071), .ZN(new_n1072));
  INV_X1    g647(.A(KEYINPUT51), .ZN(new_n1073));
  INV_X1    g648(.A(new_n1071), .ZN(new_n1074));
  AOI211_X1 g649(.A(new_n1073), .B(new_n1074), .C1(new_n1068), .C2(G168), .ZN(new_n1075));
  OAI21_X1  g650(.A(new_n1069), .B1(new_n1072), .B2(new_n1075), .ZN(new_n1076));
  NOR2_X1   g651(.A1(new_n988), .A2(G2090), .ZN(new_n1077));
  NOR2_X1   g652(.A1(new_n957), .A2(new_n958), .ZN(new_n1078));
  AOI21_X1  g653(.A(new_n1077), .B1(new_n1078), .B2(new_n785), .ZN(new_n1079));
  OAI21_X1  g654(.A(new_n1064), .B1(new_n1079), .B2(new_n1045), .ZN(new_n1080));
  AND3_X1   g655(.A1(new_n1066), .A2(new_n1076), .A3(new_n1080), .ZN(new_n1081));
  AND4_X1   g656(.A1(new_n981), .A2(new_n1036), .A3(new_n1040), .A4(new_n1081), .ZN(new_n1082));
  NOR3_X1   g657(.A1(new_n1068), .A2(new_n1045), .A3(G286), .ZN(new_n1083));
  NAND3_X1  g658(.A1(new_n1066), .A2(new_n1080), .A3(new_n1083), .ZN(new_n1084));
  INV_X1    g659(.A(KEYINPUT63), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n1084), .A2(new_n1085), .ZN(new_n1086));
  AND2_X1   g661(.A1(new_n1083), .A2(KEYINPUT63), .ZN(new_n1087));
  OAI211_X1 g662(.A(new_n1066), .B(new_n1087), .C1(new_n1065), .C2(new_n1059), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n1086), .A2(new_n1088), .ZN(new_n1089));
  INV_X1    g664(.A(KEYINPUT62), .ZN(new_n1090));
  NAND2_X1  g665(.A1(new_n1076), .A2(new_n1090), .ZN(new_n1091));
  OAI211_X1 g666(.A(KEYINPUT62), .B(new_n1069), .C1(new_n1072), .C2(new_n1075), .ZN(new_n1092));
  NAND2_X1  g667(.A1(new_n1091), .A2(new_n1092), .ZN(new_n1093));
  AND2_X1   g668(.A1(new_n1066), .A2(new_n1080), .ZN(new_n1094));
  NAND3_X1  g669(.A1(new_n1093), .A2(new_n1094), .A3(new_n974), .ZN(new_n1095));
  XNOR2_X1  g670(.A(new_n1046), .B(KEYINPUT115), .ZN(new_n1096));
  NAND3_X1  g671(.A1(new_n1047), .A2(new_n1051), .A3(new_n778), .ZN(new_n1097));
  AOI21_X1  g672(.A(new_n1096), .B1(new_n1097), .B2(new_n1042), .ZN(new_n1098));
  AND2_X1   g673(.A1(new_n1059), .A2(new_n1065), .ZN(new_n1099));
  INV_X1    g674(.A(new_n1056), .ZN(new_n1100));
  AOI21_X1  g675(.A(new_n1098), .B1(new_n1099), .B2(new_n1100), .ZN(new_n1101));
  NAND3_X1  g676(.A1(new_n1089), .A2(new_n1095), .A3(new_n1101), .ZN(new_n1102));
  OAI21_X1  g677(.A(new_n935), .B1(new_n1082), .B2(new_n1102), .ZN(new_n1103));
  NAND2_X1  g678(.A1(new_n926), .A2(new_n713), .ZN(new_n1104));
  INV_X1    g679(.A(KEYINPUT46), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n922), .A2(new_n923), .ZN(new_n1106));
  AOI22_X1  g681(.A1(new_n1104), .A2(new_n922), .B1(new_n1105), .B2(new_n1106), .ZN(new_n1107));
  NOR2_X1   g682(.A1(new_n1106), .A2(new_n1105), .ZN(new_n1108));
  XNOR2_X1  g683(.A(new_n1108), .B(KEYINPUT126), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n1107), .A2(new_n1109), .ZN(new_n1110));
  XNOR2_X1  g685(.A(new_n1110), .B(KEYINPUT127), .ZN(new_n1111));
  OR2_X1    g686(.A1(new_n1111), .A2(KEYINPUT47), .ZN(new_n1112));
  NAND2_X1  g687(.A1(new_n1111), .A2(KEYINPUT47), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n929), .A2(new_n922), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n932), .A2(new_n922), .ZN(new_n1115));
  XNOR2_X1  g690(.A(new_n1115), .B(KEYINPUT48), .ZN(new_n1116));
  NAND2_X1  g691(.A1(new_n924), .A2(new_n926), .ZN(new_n1117));
  OAI22_X1  g692(.A1(new_n1117), .A2(new_n927), .B1(G2067), .B2(new_n685), .ZN(new_n1118));
  AOI22_X1  g693(.A1(new_n1114), .A2(new_n1116), .B1(new_n1118), .B2(new_n922), .ZN(new_n1119));
  AND3_X1   g694(.A1(new_n1112), .A2(new_n1113), .A3(new_n1119), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n1103), .A2(new_n1120), .ZN(G329));
  assign    G231 = 1'b0;
  NAND2_X1  g696(.A1(new_n864), .A2(new_n865), .ZN(new_n1123));
  INV_X1    g697(.A(G319), .ZN(new_n1124));
  NOR4_X1   g698(.A1(G229), .A2(G401), .A3(new_n1124), .A4(G227), .ZN(new_n1125));
  NAND3_X1  g699(.A1(new_n1123), .A2(new_n907), .A3(new_n1125), .ZN(G225));
  INV_X1    g700(.A(G225), .ZN(G308));
endmodule


