//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 0 1 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 0 1 0 1 0 0 0 0 1 0 0 0 0 0 1 0 0 0 0 0 0 1 0 0 1 0 1 0 0 0 0 1 0 0 1 0 0 1 1 1 1 1 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:21:35 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n615,
    new_n616, new_n617, new_n618, new_n619, new_n620, new_n621, new_n622,
    new_n624, new_n625, new_n626, new_n627, new_n628, new_n629, new_n630,
    new_n631, new_n632, new_n633, new_n634, new_n635, new_n637, new_n638,
    new_n639, new_n640, new_n641, new_n642, new_n643, new_n644, new_n645,
    new_n646, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n666, new_n667, new_n668,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n686, new_n687, new_n689, new_n690, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n697, new_n698, new_n699, new_n700,
    new_n702, new_n703, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n727, new_n728, new_n729, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n885, new_n886, new_n887, new_n888, new_n890, new_n891, new_n892,
    new_n893, new_n894, new_n895, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n945,
    new_n946, new_n947, new_n948, new_n949, new_n950, new_n951, new_n952,
    new_n953, new_n954, new_n955, new_n956, new_n957, new_n958;
  INV_X1    g000(.A(G125), .ZN(new_n187));
  NOR3_X1   g001(.A1(new_n187), .A2(KEYINPUT16), .A3(G140), .ZN(new_n188));
  XNOR2_X1  g002(.A(G125), .B(G140), .ZN(new_n189));
  AOI21_X1  g003(.A(new_n188), .B1(new_n189), .B2(KEYINPUT16), .ZN(new_n190));
  OR2_X1    g004(.A1(new_n190), .A2(G146), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n190), .A2(G146), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n191), .A2(new_n192), .ZN(new_n193));
  INV_X1    g007(.A(G237), .ZN(new_n194));
  INV_X1    g008(.A(G953), .ZN(new_n195));
  NAND3_X1  g009(.A1(new_n194), .A2(new_n195), .A3(G214), .ZN(new_n196));
  INV_X1    g010(.A(KEYINPUT88), .ZN(new_n197));
  INV_X1    g011(.A(G143), .ZN(new_n198));
  NAND3_X1  g012(.A1(new_n196), .A2(new_n197), .A3(new_n198), .ZN(new_n199));
  NOR2_X1   g013(.A1(G237), .A2(G953), .ZN(new_n200));
  OAI211_X1 g014(.A(new_n200), .B(G214), .C1(KEYINPUT88), .C2(G143), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n199), .A2(new_n201), .ZN(new_n202));
  NAND3_X1  g016(.A1(new_n202), .A2(KEYINPUT17), .A3(G131), .ZN(new_n203));
  INV_X1    g017(.A(new_n203), .ZN(new_n204));
  OAI21_X1  g018(.A(KEYINPUT92), .B1(new_n193), .B2(new_n204), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n202), .A2(G131), .ZN(new_n206));
  INV_X1    g020(.A(KEYINPUT17), .ZN(new_n207));
  INV_X1    g021(.A(G131), .ZN(new_n208));
  NAND3_X1  g022(.A1(new_n199), .A2(new_n208), .A3(new_n201), .ZN(new_n209));
  NAND3_X1  g023(.A1(new_n206), .A2(new_n207), .A3(new_n209), .ZN(new_n210));
  INV_X1    g024(.A(KEYINPUT92), .ZN(new_n211));
  NAND4_X1  g025(.A1(new_n191), .A2(new_n203), .A3(new_n211), .A4(new_n192), .ZN(new_n212));
  NAND3_X1  g026(.A1(new_n205), .A2(new_n210), .A3(new_n212), .ZN(new_n213));
  INV_X1    g027(.A(G146), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n214), .A2(KEYINPUT64), .ZN(new_n215));
  INV_X1    g029(.A(KEYINPUT64), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n216), .A2(G146), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n215), .A2(new_n217), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n218), .A2(new_n189), .ZN(new_n219));
  OAI21_X1  g033(.A(new_n219), .B1(new_n214), .B2(new_n189), .ZN(new_n220));
  NOR2_X1   g034(.A1(new_n202), .A2(KEYINPUT89), .ZN(new_n221));
  AOI21_X1  g035(.A(new_n221), .B1(KEYINPUT18), .B2(G131), .ZN(new_n222));
  NAND2_X1  g036(.A1(KEYINPUT18), .A2(G131), .ZN(new_n223));
  NOR3_X1   g037(.A1(new_n202), .A2(KEYINPUT89), .A3(new_n223), .ZN(new_n224));
  OAI21_X1  g038(.A(new_n220), .B1(new_n222), .B2(new_n224), .ZN(new_n225));
  XOR2_X1   g039(.A(G113), .B(G122), .Z(new_n226));
  XNOR2_X1  g040(.A(new_n226), .B(KEYINPUT91), .ZN(new_n227));
  INV_X1    g041(.A(G104), .ZN(new_n228));
  XNOR2_X1  g042(.A(new_n227), .B(new_n228), .ZN(new_n229));
  NAND3_X1  g043(.A1(new_n213), .A2(new_n225), .A3(new_n229), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n206), .A2(new_n209), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n231), .A2(KEYINPUT90), .ZN(new_n232));
  INV_X1    g046(.A(KEYINPUT90), .ZN(new_n233));
  NAND3_X1  g047(.A1(new_n206), .A2(new_n233), .A3(new_n209), .ZN(new_n234));
  XNOR2_X1  g048(.A(new_n189), .B(KEYINPUT19), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n235), .A2(new_n218), .ZN(new_n236));
  NAND4_X1  g050(.A1(new_n232), .A2(new_n234), .A3(new_n192), .A4(new_n236), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n225), .A2(new_n237), .ZN(new_n238));
  INV_X1    g052(.A(new_n229), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n238), .A2(new_n239), .ZN(new_n240));
  AOI21_X1  g054(.A(G475), .B1(new_n230), .B2(new_n240), .ZN(new_n241));
  INV_X1    g055(.A(KEYINPUT20), .ZN(new_n242));
  INV_X1    g056(.A(G902), .ZN(new_n243));
  NAND3_X1  g057(.A1(new_n241), .A2(new_n242), .A3(new_n243), .ZN(new_n244));
  AOI21_X1  g058(.A(new_n242), .B1(new_n241), .B2(new_n243), .ZN(new_n245));
  OAI21_X1  g059(.A(new_n244), .B1(new_n245), .B2(KEYINPUT93), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n230), .A2(new_n240), .ZN(new_n247));
  INV_X1    g061(.A(G475), .ZN(new_n248));
  NAND3_X1  g062(.A1(new_n247), .A2(new_n248), .A3(new_n243), .ZN(new_n249));
  OR3_X1    g063(.A1(new_n249), .A2(KEYINPUT93), .A3(KEYINPUT20), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n246), .A2(new_n250), .ZN(new_n251));
  INV_X1    g065(.A(new_n230), .ZN(new_n252));
  AOI21_X1  g066(.A(new_n229), .B1(new_n213), .B2(new_n225), .ZN(new_n253));
  OAI21_X1  g067(.A(new_n243), .B1(new_n252), .B2(new_n253), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n254), .A2(G475), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n251), .A2(new_n255), .ZN(new_n256));
  XNOR2_X1  g070(.A(G116), .B(G122), .ZN(new_n257));
  XNOR2_X1  g071(.A(new_n257), .B(G107), .ZN(new_n258));
  INV_X1    g072(.A(KEYINPUT94), .ZN(new_n259));
  INV_X1    g073(.A(G128), .ZN(new_n260));
  NOR2_X1   g074(.A1(new_n260), .A2(G143), .ZN(new_n261));
  NOR2_X1   g075(.A1(new_n261), .A2(KEYINPUT13), .ZN(new_n262));
  NOR2_X1   g076(.A1(new_n198), .A2(G128), .ZN(new_n263));
  OAI21_X1  g077(.A(new_n259), .B1(new_n262), .B2(new_n263), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n261), .A2(KEYINPUT13), .ZN(new_n265));
  INV_X1    g079(.A(new_n263), .ZN(new_n266));
  OAI211_X1 g080(.A(new_n266), .B(KEYINPUT94), .C1(KEYINPUT13), .C2(new_n261), .ZN(new_n267));
  NAND3_X1  g081(.A1(new_n264), .A2(new_n265), .A3(new_n267), .ZN(new_n268));
  AOI21_X1  g082(.A(new_n258), .B1(new_n268), .B2(G134), .ZN(new_n269));
  NOR3_X1   g083(.A1(new_n261), .A2(new_n263), .A3(G134), .ZN(new_n270));
  INV_X1    g084(.A(new_n270), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n269), .A2(new_n271), .ZN(new_n272));
  OAI21_X1  g086(.A(G134), .B1(new_n261), .B2(new_n263), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n271), .A2(new_n273), .ZN(new_n274));
  INV_X1    g088(.A(G107), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n257), .A2(new_n275), .ZN(new_n276));
  INV_X1    g090(.A(G116), .ZN(new_n277));
  NAND3_X1  g091(.A1(new_n277), .A2(KEYINPUT14), .A3(G122), .ZN(new_n278));
  INV_X1    g092(.A(new_n257), .ZN(new_n279));
  OAI211_X1 g093(.A(G107), .B(new_n278), .C1(new_n279), .C2(KEYINPUT14), .ZN(new_n280));
  NAND3_X1  g094(.A1(new_n274), .A2(new_n276), .A3(new_n280), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n272), .A2(new_n281), .ZN(new_n282));
  XOR2_X1   g096(.A(KEYINPUT9), .B(G234), .Z(new_n283));
  INV_X1    g097(.A(new_n283), .ZN(new_n284));
  INV_X1    g098(.A(G217), .ZN(new_n285));
  NOR3_X1   g099(.A1(new_n284), .A2(new_n285), .A3(G953), .ZN(new_n286));
  INV_X1    g100(.A(new_n286), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n282), .A2(new_n287), .ZN(new_n288));
  NAND3_X1  g102(.A1(new_n272), .A2(new_n281), .A3(new_n286), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  AOI21_X1  g104(.A(KEYINPUT95), .B1(new_n290), .B2(new_n243), .ZN(new_n291));
  INV_X1    g105(.A(G478), .ZN(new_n292));
  NOR2_X1   g106(.A1(new_n292), .A2(KEYINPUT15), .ZN(new_n293));
  OR2_X1    g107(.A1(new_n291), .A2(new_n293), .ZN(new_n294));
  INV_X1    g108(.A(KEYINPUT95), .ZN(new_n295));
  AOI211_X1 g109(.A(new_n295), .B(G902), .C1(new_n288), .C2(new_n289), .ZN(new_n296));
  OAI21_X1  g110(.A(new_n293), .B1(new_n291), .B2(new_n296), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n294), .A2(new_n297), .ZN(new_n298));
  INV_X1    g112(.A(G952), .ZN(new_n299));
  NOR2_X1   g113(.A1(new_n299), .A2(G953), .ZN(new_n300));
  NAND2_X1  g114(.A1(G234), .A2(G237), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  INV_X1    g116(.A(new_n302), .ZN(new_n303));
  XOR2_X1   g117(.A(KEYINPUT21), .B(G898), .Z(new_n304));
  INV_X1    g118(.A(new_n304), .ZN(new_n305));
  NAND3_X1  g119(.A1(new_n301), .A2(G902), .A3(G953), .ZN(new_n306));
  INV_X1    g120(.A(new_n306), .ZN(new_n307));
  AOI21_X1  g121(.A(new_n303), .B1(new_n305), .B2(new_n307), .ZN(new_n308));
  NOR3_X1   g122(.A1(new_n256), .A2(new_n298), .A3(new_n308), .ZN(new_n309));
  NAND3_X1  g123(.A1(new_n215), .A2(new_n217), .A3(new_n198), .ZN(new_n310));
  NOR2_X1   g124(.A1(new_n198), .A2(G146), .ZN(new_n311));
  INV_X1    g125(.A(new_n311), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n310), .A2(new_n312), .ZN(new_n313));
  AND2_X1   g127(.A1(KEYINPUT0), .A2(G128), .ZN(new_n314));
  NOR2_X1   g128(.A1(KEYINPUT0), .A2(G128), .ZN(new_n315));
  NOR2_X1   g129(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n313), .A2(new_n316), .ZN(new_n317));
  OAI21_X1  g131(.A(KEYINPUT65), .B1(new_n214), .B2(G143), .ZN(new_n318));
  INV_X1    g132(.A(KEYINPUT65), .ZN(new_n319));
  NAND3_X1  g133(.A1(new_n319), .A2(new_n198), .A3(G146), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n318), .A2(new_n320), .ZN(new_n321));
  XNOR2_X1  g135(.A(KEYINPUT64), .B(G146), .ZN(new_n322));
  OAI211_X1 g136(.A(new_n321), .B(new_n314), .C1(new_n198), .C2(new_n322), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n317), .A2(new_n323), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n324), .A2(G125), .ZN(new_n325));
  INV_X1    g139(.A(KEYINPUT1), .ZN(new_n326));
  AOI21_X1  g140(.A(new_n326), .B1(new_n218), .B2(G143), .ZN(new_n327));
  OAI21_X1  g141(.A(new_n313), .B1(new_n327), .B2(new_n260), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n218), .A2(G143), .ZN(new_n329));
  NAND4_X1  g143(.A1(new_n329), .A2(new_n326), .A3(G128), .A4(new_n321), .ZN(new_n330));
  NAND3_X1  g144(.A1(new_n328), .A2(new_n187), .A3(new_n330), .ZN(new_n331));
  INV_X1    g145(.A(G224), .ZN(new_n332));
  NOR2_X1   g146(.A1(new_n332), .A2(G953), .ZN(new_n333));
  INV_X1    g147(.A(new_n333), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n334), .A2(KEYINPUT7), .ZN(new_n335));
  NAND3_X1  g149(.A1(new_n325), .A2(new_n331), .A3(new_n335), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n325), .A2(new_n331), .ZN(new_n337));
  NAND3_X1  g151(.A1(new_n337), .A2(KEYINPUT7), .A3(new_n334), .ZN(new_n338));
  INV_X1    g152(.A(KEYINPUT5), .ZN(new_n339));
  INV_X1    g153(.A(G119), .ZN(new_n340));
  NAND3_X1  g154(.A1(new_n339), .A2(new_n340), .A3(G116), .ZN(new_n341));
  INV_X1    g155(.A(KEYINPUT86), .ZN(new_n342));
  XNOR2_X1  g156(.A(new_n341), .B(new_n342), .ZN(new_n343));
  INV_X1    g157(.A(KEYINPUT69), .ZN(new_n344));
  OAI21_X1  g158(.A(new_n344), .B1(new_n277), .B2(G119), .ZN(new_n345));
  NAND3_X1  g159(.A1(new_n340), .A2(KEYINPUT69), .A3(G116), .ZN(new_n346));
  OAI211_X1 g160(.A(new_n345), .B(new_n346), .C1(G116), .C2(new_n340), .ZN(new_n347));
  OAI211_X1 g161(.A(new_n343), .B(G113), .C1(new_n339), .C2(new_n347), .ZN(new_n348));
  XNOR2_X1  g162(.A(KEYINPUT2), .B(G113), .ZN(new_n349));
  OR2_X1    g163(.A1(new_n347), .A2(new_n349), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n348), .A2(new_n350), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n228), .A2(G107), .ZN(new_n352));
  INV_X1    g166(.A(new_n352), .ZN(new_n353));
  NOR2_X1   g167(.A1(new_n228), .A2(G107), .ZN(new_n354));
  OAI21_X1  g168(.A(G101), .B1(new_n353), .B2(new_n354), .ZN(new_n355));
  OAI21_X1  g169(.A(KEYINPUT3), .B1(new_n228), .B2(G107), .ZN(new_n356));
  INV_X1    g170(.A(KEYINPUT3), .ZN(new_n357));
  NAND3_X1  g171(.A1(new_n357), .A2(new_n275), .A3(G104), .ZN(new_n358));
  INV_X1    g172(.A(G101), .ZN(new_n359));
  NAND4_X1  g173(.A1(new_n356), .A2(new_n358), .A3(new_n359), .A4(new_n352), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n355), .A2(new_n360), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n351), .A2(new_n361), .ZN(new_n362));
  INV_X1    g176(.A(new_n361), .ZN(new_n363));
  NAND3_X1  g177(.A1(new_n348), .A2(new_n350), .A3(new_n363), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n362), .A2(new_n364), .ZN(new_n365));
  XNOR2_X1  g179(.A(G110), .B(G122), .ZN(new_n366));
  XOR2_X1   g180(.A(new_n366), .B(KEYINPUT8), .Z(new_n367));
  INV_X1    g181(.A(new_n367), .ZN(new_n368));
  AOI22_X1  g182(.A1(new_n336), .A2(new_n338), .B1(new_n365), .B2(new_n368), .ZN(new_n369));
  XNOR2_X1  g183(.A(new_n347), .B(new_n349), .ZN(new_n370));
  NAND3_X1  g184(.A1(new_n356), .A2(new_n358), .A3(new_n352), .ZN(new_n371));
  NAND2_X1  g185(.A1(KEYINPUT83), .A2(KEYINPUT4), .ZN(new_n372));
  NAND3_X1  g186(.A1(new_n371), .A2(G101), .A3(new_n372), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n371), .A2(G101), .ZN(new_n374));
  NAND4_X1  g188(.A1(new_n374), .A2(KEYINPUT83), .A3(KEYINPUT4), .A4(new_n360), .ZN(new_n375));
  NAND3_X1  g189(.A1(new_n370), .A2(new_n373), .A3(new_n375), .ZN(new_n376));
  NAND3_X1  g190(.A1(new_n376), .A2(new_n364), .A3(new_n366), .ZN(new_n377));
  AOI21_X1  g191(.A(G902), .B1(new_n369), .B2(new_n377), .ZN(new_n378));
  XNOR2_X1  g192(.A(new_n337), .B(new_n333), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n376), .A2(new_n364), .ZN(new_n380));
  INV_X1    g194(.A(KEYINPUT6), .ZN(new_n381));
  INV_X1    g195(.A(new_n366), .ZN(new_n382));
  NAND4_X1  g196(.A1(new_n380), .A2(KEYINPUT87), .A3(new_n381), .A4(new_n382), .ZN(new_n383));
  AND3_X1   g197(.A1(new_n380), .A2(KEYINPUT87), .A3(new_n382), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n377), .A2(KEYINPUT6), .ZN(new_n385));
  OAI211_X1 g199(.A(new_n379), .B(new_n383), .C1(new_n384), .C2(new_n385), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n378), .A2(new_n386), .ZN(new_n387));
  OAI21_X1  g201(.A(G210), .B1(G237), .B2(G902), .ZN(new_n388));
  INV_X1    g202(.A(new_n388), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n387), .A2(new_n389), .ZN(new_n390));
  NAND3_X1  g204(.A1(new_n378), .A2(new_n388), .A3(new_n386), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n390), .A2(new_n391), .ZN(new_n392));
  INV_X1    g206(.A(new_n392), .ZN(new_n393));
  OAI21_X1  g207(.A(G214), .B1(G237), .B2(G902), .ZN(new_n394));
  INV_X1    g208(.A(new_n394), .ZN(new_n395));
  NOR2_X1   g209(.A1(new_n393), .A2(new_n395), .ZN(new_n396));
  OAI21_X1  g210(.A(G221), .B1(new_n284), .B2(G902), .ZN(new_n397));
  XNOR2_X1  g211(.A(new_n397), .B(KEYINPUT81), .ZN(new_n398));
  INV_X1    g212(.A(new_n398), .ZN(new_n399));
  INV_X1    g213(.A(G469), .ZN(new_n400));
  INV_X1    g214(.A(KEYINPUT85), .ZN(new_n401));
  INV_X1    g215(.A(G137), .ZN(new_n402));
  AND2_X1   g216(.A1(new_n402), .A2(KEYINPUT68), .ZN(new_n403));
  NOR2_X1   g217(.A1(new_n402), .A2(KEYINPUT68), .ZN(new_n404));
  OAI211_X1 g218(.A(KEYINPUT11), .B(G134), .C1(new_n403), .C2(new_n404), .ZN(new_n405));
  INV_X1    g219(.A(G134), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n406), .A2(G137), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n405), .A2(new_n407), .ZN(new_n408));
  AOI21_X1  g222(.A(KEYINPUT11), .B1(new_n402), .B2(G134), .ZN(new_n409));
  XNOR2_X1  g223(.A(new_n409), .B(KEYINPUT67), .ZN(new_n410));
  OAI21_X1  g224(.A(G131), .B1(new_n408), .B2(new_n410), .ZN(new_n411));
  INV_X1    g225(.A(KEYINPUT67), .ZN(new_n412));
  XNOR2_X1  g226(.A(new_n409), .B(new_n412), .ZN(new_n413));
  NAND4_X1  g227(.A1(new_n413), .A2(new_n208), .A3(new_n407), .A4(new_n405), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n411), .A2(new_n414), .ZN(new_n415));
  INV_X1    g229(.A(new_n415), .ZN(new_n416));
  AOI22_X1  g230(.A1(new_n218), .A2(G143), .B1(new_n318), .B2(new_n320), .ZN(new_n417));
  AOI22_X1  g231(.A1(new_n417), .A2(new_n314), .B1(new_n313), .B2(new_n316), .ZN(new_n418));
  AND3_X1   g232(.A1(new_n418), .A2(new_n375), .A3(new_n373), .ZN(new_n419));
  OAI21_X1  g233(.A(G128), .B1(new_n311), .B2(new_n326), .ZN(new_n420));
  AND2_X1   g234(.A1(new_n318), .A2(new_n320), .ZN(new_n421));
  AOI21_X1  g235(.A(new_n198), .B1(new_n215), .B2(new_n217), .ZN(new_n422));
  OAI21_X1  g236(.A(new_n420), .B1(new_n421), .B2(new_n422), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n330), .A2(new_n423), .ZN(new_n424));
  AOI21_X1  g238(.A(KEYINPUT10), .B1(new_n424), .B2(new_n363), .ZN(new_n425));
  NOR2_X1   g239(.A1(new_n419), .A2(new_n425), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n328), .A2(new_n330), .ZN(new_n427));
  NAND3_X1  g241(.A1(new_n427), .A2(KEYINPUT10), .A3(new_n363), .ZN(new_n428));
  INV_X1    g242(.A(KEYINPUT84), .ZN(new_n429));
  NOR2_X1   g243(.A1(new_n428), .A2(new_n429), .ZN(new_n430));
  INV_X1    g244(.A(KEYINPUT10), .ZN(new_n431));
  AOI21_X1  g245(.A(new_n431), .B1(new_n328), .B2(new_n330), .ZN(new_n432));
  AOI21_X1  g246(.A(KEYINPUT84), .B1(new_n432), .B2(new_n363), .ZN(new_n433));
  OAI211_X1 g247(.A(new_n416), .B(new_n426), .C1(new_n430), .C2(new_n433), .ZN(new_n434));
  XNOR2_X1  g248(.A(G110), .B(G140), .ZN(new_n435));
  XNOR2_X1  g249(.A(new_n435), .B(KEYINPUT82), .ZN(new_n436));
  AND2_X1   g250(.A1(new_n195), .A2(G227), .ZN(new_n437));
  XNOR2_X1  g251(.A(new_n436), .B(new_n437), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n434), .A2(new_n438), .ZN(new_n439));
  NAND3_X1  g253(.A1(new_n418), .A2(new_n375), .A3(new_n373), .ZN(new_n440));
  AOI21_X1  g254(.A(new_n361), .B1(new_n330), .B2(new_n423), .ZN(new_n441));
  OAI21_X1  g255(.A(new_n440), .B1(KEYINPUT10), .B2(new_n441), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n428), .A2(new_n429), .ZN(new_n443));
  NAND3_X1  g257(.A1(new_n432), .A2(KEYINPUT84), .A3(new_n363), .ZN(new_n444));
  AOI21_X1  g258(.A(new_n442), .B1(new_n443), .B2(new_n444), .ZN(new_n445));
  NOR2_X1   g259(.A1(new_n445), .A2(new_n416), .ZN(new_n446));
  NOR2_X1   g260(.A1(new_n439), .A2(new_n446), .ZN(new_n447));
  AND3_X1   g261(.A1(new_n328), .A2(new_n330), .A3(new_n361), .ZN(new_n448));
  OAI21_X1  g262(.A(new_n415), .B1(new_n448), .B2(new_n441), .ZN(new_n449));
  INV_X1    g263(.A(KEYINPUT12), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n449), .A2(new_n450), .ZN(new_n451));
  OAI211_X1 g265(.A(KEYINPUT12), .B(new_n415), .C1(new_n448), .C2(new_n441), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n451), .A2(new_n452), .ZN(new_n453));
  AOI21_X1  g267(.A(new_n438), .B1(new_n453), .B2(new_n434), .ZN(new_n454));
  OAI21_X1  g268(.A(new_n401), .B1(new_n447), .B2(new_n454), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n453), .A2(new_n434), .ZN(new_n456));
  INV_X1    g270(.A(new_n438), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  AOI21_X1  g272(.A(new_n457), .B1(new_n445), .B2(new_n416), .ZN(new_n459));
  OAI21_X1  g273(.A(new_n426), .B1(new_n430), .B2(new_n433), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n460), .A2(new_n415), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n459), .A2(new_n461), .ZN(new_n462));
  NAND3_X1  g276(.A1(new_n458), .A2(new_n462), .A3(KEYINPUT85), .ZN(new_n463));
  AOI21_X1  g277(.A(new_n400), .B1(new_n455), .B2(new_n463), .ZN(new_n464));
  AOI21_X1  g278(.A(new_n438), .B1(new_n461), .B2(new_n434), .ZN(new_n465));
  AND3_X1   g279(.A1(new_n453), .A2(new_n434), .A3(new_n438), .ZN(new_n466));
  OAI211_X1 g280(.A(new_n400), .B(new_n243), .C1(new_n465), .C2(new_n466), .ZN(new_n467));
  NOR2_X1   g281(.A1(new_n400), .A2(new_n243), .ZN(new_n468));
  INV_X1    g282(.A(new_n468), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n467), .A2(new_n469), .ZN(new_n470));
  OAI21_X1  g284(.A(new_n399), .B1(new_n464), .B2(new_n470), .ZN(new_n471));
  INV_X1    g285(.A(new_n471), .ZN(new_n472));
  AND3_X1   g286(.A1(new_n309), .A2(new_n396), .A3(new_n472), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n415), .A2(new_n418), .ZN(new_n474));
  XNOR2_X1  g288(.A(KEYINPUT68), .B(G137), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n475), .A2(new_n406), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n402), .A2(G134), .ZN(new_n477));
  AOI21_X1  g291(.A(new_n208), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  AOI21_X1  g292(.A(new_n478), .B1(new_n328), .B2(new_n330), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n479), .A2(new_n414), .ZN(new_n480));
  NAND3_X1  g294(.A1(new_n474), .A2(new_n480), .A3(KEYINPUT30), .ZN(new_n481));
  AND3_X1   g295(.A1(new_n317), .A2(KEYINPUT66), .A3(new_n323), .ZN(new_n482));
  AOI21_X1  g296(.A(KEYINPUT66), .B1(new_n317), .B2(new_n323), .ZN(new_n483));
  NOR2_X1   g297(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  AOI22_X1  g298(.A1(new_n484), .A2(new_n415), .B1(new_n414), .B2(new_n479), .ZN(new_n485));
  OAI211_X1 g299(.A(new_n370), .B(new_n481), .C1(new_n485), .C2(KEYINPUT30), .ZN(new_n486));
  INV_X1    g300(.A(new_n370), .ZN(new_n487));
  NAND3_X1  g301(.A1(new_n474), .A2(new_n480), .A3(new_n487), .ZN(new_n488));
  XNOR2_X1  g302(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n489));
  XNOR2_X1  g303(.A(new_n489), .B(G101), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n200), .A2(G210), .ZN(new_n491));
  XNOR2_X1  g305(.A(new_n490), .B(new_n491), .ZN(new_n492));
  NAND3_X1  g306(.A1(new_n486), .A2(new_n488), .A3(new_n492), .ZN(new_n493));
  INV_X1    g307(.A(KEYINPUT31), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  NAND4_X1  g309(.A1(new_n486), .A2(KEYINPUT31), .A3(new_n488), .A4(new_n492), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n488), .A2(KEYINPUT28), .ZN(new_n498));
  AOI22_X1  g312(.A1(new_n415), .A2(new_n418), .B1(new_n479), .B2(new_n414), .ZN(new_n499));
  INV_X1    g313(.A(KEYINPUT28), .ZN(new_n500));
  NAND3_X1  g314(.A1(new_n499), .A2(new_n500), .A3(new_n487), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n498), .A2(new_n501), .ZN(new_n502));
  OR2_X1    g316(.A1(new_n485), .A2(new_n487), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  INV_X1    g318(.A(new_n492), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n497), .A2(new_n506), .ZN(new_n507));
  NOR2_X1   g321(.A1(G472), .A2(G902), .ZN(new_n508));
  NAND3_X1  g322(.A1(new_n507), .A2(KEYINPUT32), .A3(new_n508), .ZN(new_n509));
  INV_X1    g323(.A(KEYINPUT73), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  INV_X1    g325(.A(KEYINPUT32), .ZN(new_n512));
  NOR2_X1   g326(.A1(new_n510), .A2(new_n512), .ZN(new_n513));
  INV_X1    g327(.A(new_n508), .ZN(new_n514));
  AOI21_X1  g328(.A(new_n514), .B1(new_n497), .B2(new_n506), .ZN(new_n515));
  OAI21_X1  g329(.A(new_n513), .B1(new_n515), .B2(KEYINPUT70), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n486), .A2(new_n488), .ZN(new_n517));
  AOI21_X1  g331(.A(KEYINPUT29), .B1(new_n517), .B2(new_n505), .ZN(new_n518));
  NAND3_X1  g332(.A1(new_n502), .A2(new_n503), .A3(new_n492), .ZN(new_n519));
  AOI21_X1  g333(.A(G902), .B1(new_n518), .B2(new_n519), .ZN(new_n520));
  INV_X1    g334(.A(KEYINPUT71), .ZN(new_n521));
  OAI21_X1  g335(.A(new_n521), .B1(new_n499), .B2(new_n487), .ZN(new_n522));
  AOI21_X1  g336(.A(new_n522), .B1(new_n498), .B2(new_n501), .ZN(new_n523));
  NOR2_X1   g337(.A1(new_n488), .A2(new_n521), .ZN(new_n524));
  OAI211_X1 g338(.A(KEYINPUT29), .B(new_n492), .C1(new_n523), .C2(new_n524), .ZN(new_n525));
  INV_X1    g339(.A(KEYINPUT72), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  INV_X1    g341(.A(new_n522), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n502), .A2(new_n528), .ZN(new_n529));
  INV_X1    g343(.A(new_n524), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  NAND4_X1  g345(.A1(new_n531), .A2(KEYINPUT72), .A3(KEYINPUT29), .A4(new_n492), .ZN(new_n532));
  NAND3_X1  g346(.A1(new_n520), .A2(new_n527), .A3(new_n532), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n533), .A2(G472), .ZN(new_n534));
  INV_X1    g348(.A(KEYINPUT70), .ZN(new_n535));
  INV_X1    g349(.A(new_n513), .ZN(new_n536));
  AOI22_X1  g350(.A1(new_n495), .A2(new_n496), .B1(new_n504), .B2(new_n505), .ZN(new_n537));
  OAI211_X1 g351(.A(new_n535), .B(new_n536), .C1(new_n537), .C2(new_n514), .ZN(new_n538));
  NAND4_X1  g352(.A1(new_n511), .A2(new_n516), .A3(new_n534), .A4(new_n538), .ZN(new_n539));
  INV_X1    g353(.A(KEYINPUT80), .ZN(new_n540));
  XOR2_X1   g354(.A(KEYINPUT22), .B(G137), .Z(new_n541));
  XNOR2_X1  g355(.A(new_n541), .B(KEYINPUT79), .ZN(new_n542));
  AND3_X1   g356(.A1(new_n195), .A2(G221), .A3(G234), .ZN(new_n543));
  XNOR2_X1  g357(.A(new_n542), .B(new_n543), .ZN(new_n544));
  XOR2_X1   g358(.A(KEYINPUT24), .B(G110), .Z(new_n545));
  INV_X1    g359(.A(new_n545), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n340), .A2(G128), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n260), .A2(G119), .ZN(new_n548));
  NAND3_X1  g362(.A1(new_n547), .A2(new_n548), .A3(KEYINPUT74), .ZN(new_n549));
  INV_X1    g363(.A(new_n549), .ZN(new_n550));
  AOI21_X1  g364(.A(KEYINPUT74), .B1(new_n547), .B2(new_n548), .ZN(new_n551));
  OAI21_X1  g365(.A(new_n546), .B1(new_n550), .B2(new_n551), .ZN(new_n552));
  INV_X1    g366(.A(KEYINPUT77), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  OAI211_X1 g368(.A(new_n546), .B(KEYINPUT77), .C1(new_n550), .C2(new_n551), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  INV_X1    g370(.A(KEYINPUT23), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n548), .A2(new_n557), .ZN(new_n558));
  NAND3_X1  g372(.A1(new_n260), .A2(KEYINPUT23), .A3(G119), .ZN(new_n559));
  NAND3_X1  g373(.A1(new_n558), .A2(new_n547), .A3(new_n559), .ZN(new_n560));
  XOR2_X1   g374(.A(KEYINPUT76), .B(G110), .Z(new_n561));
  NOR2_X1   g375(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  OAI211_X1 g376(.A(new_n219), .B(new_n192), .C1(new_n556), .C2(new_n562), .ZN(new_n563));
  INV_X1    g377(.A(KEYINPUT78), .ZN(new_n564));
  INV_X1    g378(.A(new_n551), .ZN(new_n565));
  NAND3_X1  g379(.A1(new_n565), .A2(new_n549), .A3(new_n545), .ZN(new_n566));
  INV_X1    g380(.A(KEYINPUT75), .ZN(new_n567));
  OR2_X1    g381(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n560), .A2(G110), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n566), .A2(new_n567), .ZN(new_n570));
  NAND4_X1  g384(.A1(new_n568), .A2(new_n193), .A3(new_n569), .A4(new_n570), .ZN(new_n571));
  AND3_X1   g385(.A1(new_n563), .A2(new_n564), .A3(new_n571), .ZN(new_n572));
  AOI21_X1  g386(.A(new_n564), .B1(new_n563), .B2(new_n571), .ZN(new_n573));
  OAI21_X1  g387(.A(new_n544), .B1(new_n572), .B2(new_n573), .ZN(new_n574));
  INV_X1    g388(.A(new_n544), .ZN(new_n575));
  NAND3_X1  g389(.A1(new_n575), .A2(new_n563), .A3(new_n571), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n574), .A2(new_n576), .ZN(new_n577));
  OAI21_X1  g391(.A(KEYINPUT25), .B1(new_n577), .B2(G902), .ZN(new_n578));
  AOI21_X1  g392(.A(new_n285), .B1(G234), .B2(new_n243), .ZN(new_n579));
  INV_X1    g393(.A(KEYINPUT25), .ZN(new_n580));
  NAND4_X1  g394(.A1(new_n574), .A2(new_n580), .A3(new_n243), .A4(new_n576), .ZN(new_n581));
  NAND3_X1  g395(.A1(new_n578), .A2(new_n579), .A3(new_n581), .ZN(new_n582));
  NOR2_X1   g396(.A1(new_n579), .A2(G902), .ZN(new_n583));
  NAND3_X1  g397(.A1(new_n574), .A2(new_n576), .A3(new_n583), .ZN(new_n584));
  AND2_X1   g398(.A1(new_n582), .A2(new_n584), .ZN(new_n585));
  AND3_X1   g399(.A1(new_n539), .A2(new_n540), .A3(new_n585), .ZN(new_n586));
  AOI21_X1  g400(.A(new_n540), .B1(new_n539), .B2(new_n585), .ZN(new_n587));
  OAI21_X1  g401(.A(new_n473), .B1(new_n586), .B2(new_n587), .ZN(new_n588));
  XNOR2_X1  g402(.A(new_n588), .B(G101), .ZN(G3));
  AND2_X1   g403(.A1(new_n585), .A2(new_n399), .ZN(new_n590));
  OR2_X1    g404(.A1(new_n464), .A2(new_n470), .ZN(new_n591));
  OAI21_X1  g405(.A(G472), .B1(new_n537), .B2(G902), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n507), .A2(new_n508), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  INV_X1    g408(.A(new_n594), .ZN(new_n595));
  AND3_X1   g409(.A1(new_n590), .A2(new_n591), .A3(new_n595), .ZN(new_n596));
  INV_X1    g410(.A(new_n308), .ZN(new_n597));
  AOI21_X1  g411(.A(new_n388), .B1(new_n378), .B2(new_n386), .ZN(new_n598));
  AOI21_X1  g412(.A(new_n395), .B1(new_n598), .B2(KEYINPUT96), .ZN(new_n599));
  OAI21_X1  g413(.A(new_n599), .B1(new_n392), .B2(KEYINPUT96), .ZN(new_n600));
  AOI22_X1  g414(.A1(new_n246), .A2(new_n250), .B1(G475), .B2(new_n254), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n290), .A2(new_n243), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n602), .A2(new_n292), .ZN(new_n603));
  OR2_X1    g417(.A1(new_n603), .A2(KEYINPUT98), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n603), .A2(KEYINPUT98), .ZN(new_n605));
  AOI21_X1  g419(.A(KEYINPUT97), .B1(new_n288), .B2(new_n289), .ZN(new_n606));
  OR2_X1    g420(.A1(new_n606), .A2(KEYINPUT33), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n606), .A2(KEYINPUT33), .ZN(new_n608));
  AOI21_X1  g422(.A(G902), .B1(new_n607), .B2(new_n608), .ZN(new_n609));
  AOI22_X1  g423(.A1(new_n604), .A2(new_n605), .B1(new_n609), .B2(G478), .ZN(new_n610));
  NOR3_X1   g424(.A1(new_n600), .A2(new_n601), .A3(new_n610), .ZN(new_n611));
  NAND3_X1  g425(.A1(new_n596), .A2(new_n597), .A3(new_n611), .ZN(new_n612));
  XNOR2_X1  g426(.A(new_n612), .B(KEYINPUT34), .ZN(new_n613));
  XNOR2_X1  g427(.A(new_n613), .B(new_n228), .ZN(G6));
  INV_X1    g428(.A(new_n298), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n249), .A2(KEYINPUT20), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n616), .A2(new_n244), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n617), .A2(new_n255), .ZN(new_n618));
  NOR3_X1   g432(.A1(new_n600), .A2(new_n615), .A3(new_n618), .ZN(new_n619));
  NAND3_X1  g433(.A1(new_n596), .A2(new_n597), .A3(new_n619), .ZN(new_n620));
  XNOR2_X1  g434(.A(new_n620), .B(KEYINPUT99), .ZN(new_n621));
  XNOR2_X1  g435(.A(KEYINPUT35), .B(G107), .ZN(new_n622));
  XNOR2_X1  g436(.A(new_n621), .B(new_n622), .ZN(G9));
  NOR2_X1   g437(.A1(new_n572), .A2(new_n573), .ZN(new_n624));
  NOR2_X1   g438(.A1(new_n544), .A2(KEYINPUT36), .ZN(new_n625));
  XOR2_X1   g439(.A(new_n624), .B(new_n625), .Z(new_n626));
  NAND2_X1  g440(.A1(new_n626), .A2(new_n583), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n627), .A2(new_n582), .ZN(new_n628));
  INV_X1    g442(.A(KEYINPUT100), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  NAND3_X1  g444(.A1(new_n627), .A2(new_n582), .A3(KEYINPUT100), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  NAND3_X1  g446(.A1(new_n473), .A2(new_n595), .A3(new_n632), .ZN(new_n633));
  XNOR2_X1  g447(.A(KEYINPUT101), .B(KEYINPUT37), .ZN(new_n634));
  XNOR2_X1  g448(.A(new_n634), .B(G110), .ZN(new_n635));
  XNOR2_X1  g449(.A(new_n633), .B(new_n635), .ZN(G12));
  INV_X1    g450(.A(G900), .ZN(new_n637));
  AOI21_X1  g451(.A(new_n303), .B1(new_n307), .B2(new_n637), .ZN(new_n638));
  INV_X1    g452(.A(new_n638), .ZN(new_n639));
  NAND4_X1  g453(.A1(new_n298), .A2(new_n617), .A3(new_n255), .A4(new_n639), .ZN(new_n640));
  NOR3_X1   g454(.A1(new_n471), .A2(new_n600), .A3(new_n640), .ZN(new_n641));
  NAND3_X1  g455(.A1(new_n539), .A2(new_n641), .A3(new_n632), .ZN(new_n642));
  INV_X1    g456(.A(KEYINPUT102), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  NAND4_X1  g458(.A1(new_n539), .A2(new_n641), .A3(new_n632), .A4(KEYINPUT102), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  XNOR2_X1  g460(.A(new_n646), .B(G128), .ZN(G30));
  XNOR2_X1  g461(.A(new_n638), .B(KEYINPUT39), .ZN(new_n648));
  INV_X1    g462(.A(new_n648), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n472), .A2(new_n649), .ZN(new_n650));
  XOR2_X1   g464(.A(new_n650), .B(KEYINPUT40), .Z(new_n651));
  XNOR2_X1  g465(.A(new_n392), .B(KEYINPUT38), .ZN(new_n652));
  INV_X1    g466(.A(new_n628), .ZN(new_n653));
  NAND4_X1  g467(.A1(new_n653), .A2(new_n394), .A3(new_n256), .A4(new_n298), .ZN(new_n654));
  XNOR2_X1  g468(.A(new_n654), .B(KEYINPUT104), .ZN(new_n655));
  AND3_X1   g469(.A1(new_n511), .A2(new_n516), .A3(new_n538), .ZN(new_n656));
  AOI211_X1 g470(.A(new_n492), .B(new_n524), .C1(new_n488), .C2(new_n528), .ZN(new_n657));
  INV_X1    g471(.A(new_n493), .ZN(new_n658));
  OR2_X1    g472(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  AND2_X1   g473(.A1(new_n659), .A2(KEYINPUT103), .ZN(new_n660));
  OAI21_X1  g474(.A(new_n243), .B1(new_n659), .B2(KEYINPUT103), .ZN(new_n661));
  OAI21_X1  g475(.A(G472), .B1(new_n660), .B2(new_n661), .ZN(new_n662));
  NAND2_X1  g476(.A1(new_n656), .A2(new_n662), .ZN(new_n663));
  NAND4_X1  g477(.A1(new_n651), .A2(new_n652), .A3(new_n655), .A4(new_n663), .ZN(new_n664));
  XNOR2_X1  g478(.A(new_n664), .B(G143), .ZN(G45));
  NOR3_X1   g479(.A1(new_n601), .A2(new_n610), .A3(new_n638), .ZN(new_n666));
  NOR2_X1   g480(.A1(new_n471), .A2(new_n600), .ZN(new_n667));
  NAND4_X1  g481(.A1(new_n539), .A2(new_n632), .A3(new_n666), .A4(new_n667), .ZN(new_n668));
  XNOR2_X1  g482(.A(new_n668), .B(G146), .ZN(G48));
  AND2_X1   g483(.A1(new_n539), .A2(new_n585), .ZN(new_n670));
  NAND2_X1  g484(.A1(new_n461), .A2(new_n434), .ZN(new_n671));
  AOI22_X1  g485(.A1(new_n671), .A2(new_n457), .B1(new_n453), .B2(new_n459), .ZN(new_n672));
  OAI21_X1  g486(.A(G469), .B1(new_n672), .B2(G902), .ZN(new_n673));
  NAND3_X1  g487(.A1(new_n673), .A2(new_n399), .A3(new_n467), .ZN(new_n674));
  INV_X1    g488(.A(KEYINPUT105), .ZN(new_n675));
  NAND2_X1  g489(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  NAND4_X1  g490(.A1(new_n673), .A2(KEYINPUT105), .A3(new_n399), .A4(new_n467), .ZN(new_n677));
  AOI21_X1  g491(.A(new_n308), .B1(new_n676), .B2(new_n677), .ZN(new_n678));
  NAND4_X1  g492(.A1(new_n670), .A2(KEYINPUT106), .A3(new_n611), .A4(new_n678), .ZN(new_n679));
  NAND4_X1  g493(.A1(new_n678), .A2(new_n539), .A3(new_n611), .A4(new_n585), .ZN(new_n680));
  INV_X1    g494(.A(KEYINPUT106), .ZN(new_n681));
  NAND2_X1  g495(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  NAND2_X1  g496(.A1(new_n679), .A2(new_n682), .ZN(new_n683));
  XNOR2_X1  g497(.A(new_n683), .B(KEYINPUT41), .ZN(new_n684));
  XNOR2_X1  g498(.A(new_n684), .B(G113), .ZN(G15));
  AND4_X1   g499(.A1(new_n539), .A2(new_n678), .A3(new_n585), .A4(new_n619), .ZN(new_n686));
  XNOR2_X1  g500(.A(KEYINPUT107), .B(G116), .ZN(new_n687));
  XNOR2_X1  g501(.A(new_n686), .B(new_n687), .ZN(G18));
  NOR2_X1   g502(.A1(new_n600), .A2(new_n674), .ZN(new_n689));
  NAND4_X1  g503(.A1(new_n539), .A2(new_n309), .A3(new_n632), .A4(new_n689), .ZN(new_n690));
  XNOR2_X1  g504(.A(new_n690), .B(G119), .ZN(G21));
  OAI21_X1  g505(.A(new_n497), .B1(new_n492), .B2(new_n531), .ZN(new_n692));
  NAND2_X1  g506(.A1(new_n692), .A2(new_n508), .ZN(new_n693));
  AND3_X1   g507(.A1(new_n585), .A2(new_n693), .A3(new_n592), .ZN(new_n694));
  NOR3_X1   g508(.A1(new_n600), .A2(new_n601), .A3(new_n615), .ZN(new_n695));
  NAND3_X1  g509(.A1(new_n678), .A2(new_n694), .A3(new_n695), .ZN(new_n696));
  NAND2_X1  g510(.A1(new_n696), .A2(KEYINPUT108), .ZN(new_n697));
  INV_X1    g511(.A(KEYINPUT108), .ZN(new_n698));
  NAND4_X1  g512(.A1(new_n678), .A2(new_n694), .A3(new_n698), .A4(new_n695), .ZN(new_n699));
  NAND2_X1  g513(.A1(new_n697), .A2(new_n699), .ZN(new_n700));
  XNOR2_X1  g514(.A(new_n700), .B(G122), .ZN(G24));
  AND2_X1   g515(.A1(new_n693), .A2(new_n592), .ZN(new_n702));
  NAND4_X1  g516(.A1(new_n666), .A2(new_n702), .A3(new_n689), .A4(new_n628), .ZN(new_n703));
  XNOR2_X1  g517(.A(new_n703), .B(G125), .ZN(G27));
  NOR2_X1   g518(.A1(new_n392), .A2(new_n395), .ZN(new_n705));
  NAND2_X1  g519(.A1(new_n705), .A2(new_n399), .ZN(new_n706));
  INV_X1    g520(.A(new_n706), .ZN(new_n707));
  INV_X1    g521(.A(new_n470), .ZN(new_n708));
  NOR2_X1   g522(.A1(new_n447), .A2(new_n454), .ZN(new_n709));
  NAND2_X1  g523(.A1(new_n709), .A2(G469), .ZN(new_n710));
  NAND2_X1  g524(.A1(new_n708), .A2(new_n710), .ZN(new_n711));
  NAND4_X1  g525(.A1(new_n539), .A2(new_n585), .A3(new_n707), .A4(new_n711), .ZN(new_n712));
  INV_X1    g526(.A(new_n666), .ZN(new_n713));
  NOR2_X1   g527(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  NAND2_X1  g528(.A1(new_n593), .A2(new_n512), .ZN(new_n715));
  NAND3_X1  g529(.A1(new_n715), .A2(KEYINPUT109), .A3(new_n509), .ZN(new_n716));
  INV_X1    g530(.A(KEYINPUT109), .ZN(new_n717));
  NOR2_X1   g531(.A1(new_n515), .A2(KEYINPUT32), .ZN(new_n718));
  NOR3_X1   g532(.A1(new_n537), .A2(new_n512), .A3(new_n514), .ZN(new_n719));
  OAI21_X1  g533(.A(new_n717), .B1(new_n718), .B2(new_n719), .ZN(new_n720));
  NAND3_X1  g534(.A1(new_n716), .A2(new_n720), .A3(new_n534), .ZN(new_n721));
  AOI21_X1  g535(.A(new_n398), .B1(new_n708), .B2(new_n710), .ZN(new_n722));
  NAND4_X1  g536(.A1(new_n721), .A2(KEYINPUT42), .A3(new_n585), .A4(new_n722), .ZN(new_n723));
  NAND2_X1  g537(.A1(new_n666), .A2(new_n705), .ZN(new_n724));
  OAI22_X1  g538(.A1(new_n714), .A2(KEYINPUT42), .B1(new_n723), .B2(new_n724), .ZN(new_n725));
  XNOR2_X1  g539(.A(new_n725), .B(G131), .ZN(G33));
  XNOR2_X1  g540(.A(new_n640), .B(KEYINPUT110), .ZN(new_n727));
  OR2_X1    g541(.A1(new_n712), .A2(new_n727), .ZN(new_n728));
  XNOR2_X1  g542(.A(new_n728), .B(KEYINPUT111), .ZN(new_n729));
  XNOR2_X1  g543(.A(new_n729), .B(new_n406), .ZN(G36));
  INV_X1    g544(.A(KEYINPUT112), .ZN(new_n731));
  INV_X1    g545(.A(KEYINPUT45), .ZN(new_n732));
  NAND3_X1  g546(.A1(new_n455), .A2(new_n463), .A3(new_n732), .ZN(new_n733));
  NAND2_X1  g547(.A1(new_n709), .A2(KEYINPUT45), .ZN(new_n734));
  NAND3_X1  g548(.A1(new_n733), .A2(new_n734), .A3(G469), .ZN(new_n735));
  NAND2_X1  g549(.A1(new_n735), .A2(new_n469), .ZN(new_n736));
  INV_X1    g550(.A(KEYINPUT46), .ZN(new_n737));
  AOI21_X1  g551(.A(new_n731), .B1(new_n736), .B2(new_n737), .ZN(new_n738));
  AOI211_X1 g552(.A(KEYINPUT112), .B(KEYINPUT46), .C1(new_n735), .C2(new_n469), .ZN(new_n739));
  NAND3_X1  g553(.A1(new_n735), .A2(KEYINPUT46), .A3(new_n469), .ZN(new_n740));
  NAND2_X1  g554(.A1(new_n740), .A2(new_n467), .ZN(new_n741));
  NOR3_X1   g555(.A1(new_n738), .A2(new_n739), .A3(new_n741), .ZN(new_n742));
  NOR2_X1   g556(.A1(new_n742), .A2(new_n398), .ZN(new_n743));
  NAND2_X1  g557(.A1(new_n594), .A2(new_n628), .ZN(new_n744));
  XNOR2_X1  g558(.A(new_n744), .B(KEYINPUT113), .ZN(new_n745));
  NAND2_X1  g559(.A1(new_n604), .A2(new_n605), .ZN(new_n746));
  NAND2_X1  g560(.A1(new_n609), .A2(G478), .ZN(new_n747));
  NAND2_X1  g561(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  NAND2_X1  g562(.A1(new_n601), .A2(new_n748), .ZN(new_n749));
  INV_X1    g563(.A(KEYINPUT43), .ZN(new_n750));
  XNOR2_X1  g564(.A(new_n749), .B(new_n750), .ZN(new_n751));
  NAND3_X1  g565(.A1(new_n745), .A2(KEYINPUT44), .A3(new_n751), .ZN(new_n752));
  AND3_X1   g566(.A1(new_n743), .A2(new_n649), .A3(new_n752), .ZN(new_n753));
  AOI21_X1  g567(.A(KEYINPUT44), .B1(new_n745), .B2(new_n751), .ZN(new_n754));
  NOR3_X1   g568(.A1(new_n754), .A2(new_n392), .A3(new_n395), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n753), .A2(new_n755), .ZN(new_n756));
  XNOR2_X1  g570(.A(new_n756), .B(G137), .ZN(G39));
  NOR3_X1   g571(.A1(new_n724), .A2(new_n539), .A3(new_n585), .ZN(new_n758));
  XOR2_X1   g572(.A(new_n758), .B(KEYINPUT114), .Z(new_n759));
  NAND2_X1  g573(.A1(new_n743), .A2(KEYINPUT47), .ZN(new_n760));
  INV_X1    g574(.A(KEYINPUT47), .ZN(new_n761));
  OAI21_X1  g575(.A(new_n761), .B1(new_n742), .B2(new_n398), .ZN(new_n762));
  NAND2_X1  g576(.A1(new_n760), .A2(new_n762), .ZN(new_n763));
  NAND2_X1  g577(.A1(new_n759), .A2(new_n763), .ZN(new_n764));
  XNOR2_X1  g578(.A(new_n764), .B(G140), .ZN(G42));
  INV_X1    g579(.A(KEYINPUT54), .ZN(new_n766));
  AND2_X1   g580(.A1(new_n668), .A2(new_n703), .ZN(new_n767));
  AND2_X1   g581(.A1(new_n722), .A2(new_n639), .ZN(new_n768));
  NAND4_X1  g582(.A1(new_n663), .A2(new_n653), .A3(new_n695), .A4(new_n768), .ZN(new_n769));
  NAND3_X1  g583(.A1(new_n646), .A2(new_n767), .A3(new_n769), .ZN(new_n770));
  INV_X1    g584(.A(KEYINPUT52), .ZN(new_n771));
  NAND2_X1  g585(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  NAND4_X1  g586(.A1(new_n646), .A2(new_n767), .A3(KEYINPUT52), .A4(new_n769), .ZN(new_n773));
  NAND2_X1  g587(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  INV_X1    g588(.A(new_n690), .ZN(new_n775));
  AOI21_X1  g589(.A(new_n775), .B1(new_n679), .B2(new_n682), .ZN(new_n776));
  AOI21_X1  g590(.A(new_n686), .B1(new_n699), .B2(new_n697), .ZN(new_n777));
  AND3_X1   g591(.A1(new_n776), .A2(new_n725), .A3(new_n777), .ZN(new_n778));
  OR3_X1    g592(.A1(new_n601), .A2(new_n610), .A3(KEYINPUT116), .ZN(new_n779));
  NAND2_X1  g593(.A1(new_n256), .A2(new_n748), .ZN(new_n780));
  NAND2_X1  g594(.A1(new_n780), .A2(KEYINPUT116), .ZN(new_n781));
  OAI211_X1 g595(.A(new_n779), .B(new_n781), .C1(new_n615), .C2(new_n256), .ZN(new_n782));
  NAND4_X1  g596(.A1(new_n782), .A2(new_n596), .A3(new_n396), .A4(new_n597), .ZN(new_n783));
  NAND4_X1  g597(.A1(new_n588), .A2(new_n783), .A3(new_n728), .A4(new_n633), .ZN(new_n784));
  AND3_X1   g598(.A1(new_n539), .A2(new_n591), .A3(new_n632), .ZN(new_n785));
  INV_X1    g599(.A(new_n618), .ZN(new_n786));
  NAND4_X1  g600(.A1(new_n785), .A2(new_n615), .A3(new_n786), .A4(new_n639), .ZN(new_n787));
  AND2_X1   g601(.A1(new_n702), .A2(new_n628), .ZN(new_n788));
  NAND3_X1  g602(.A1(new_n788), .A2(new_n666), .A3(new_n711), .ZN(new_n789));
  AOI21_X1  g603(.A(new_n706), .B1(new_n787), .B2(new_n789), .ZN(new_n790));
  NOR2_X1   g604(.A1(new_n784), .A2(new_n790), .ZN(new_n791));
  AND3_X1   g605(.A1(new_n774), .A2(new_n778), .A3(new_n791), .ZN(new_n792));
  AND2_X1   g606(.A1(new_n774), .A2(KEYINPUT117), .ZN(new_n793));
  OAI21_X1  g607(.A(new_n792), .B1(new_n793), .B2(KEYINPUT53), .ZN(new_n794));
  AOI21_X1  g608(.A(KEYINPUT53), .B1(new_n774), .B2(KEYINPUT117), .ZN(new_n795));
  NAND3_X1  g609(.A1(new_n774), .A2(new_n778), .A3(new_n791), .ZN(new_n796));
  NAND2_X1  g610(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  AOI21_X1  g611(.A(new_n766), .B1(new_n794), .B2(new_n797), .ZN(new_n798));
  INV_X1    g612(.A(KEYINPUT118), .ZN(new_n799));
  NAND4_X1  g613(.A1(new_n776), .A2(new_n725), .A3(new_n799), .A4(new_n777), .ZN(new_n800));
  AND2_X1   g614(.A1(new_n800), .A2(KEYINPUT53), .ZN(new_n801));
  NAND3_X1  g615(.A1(new_n776), .A2(new_n725), .A3(new_n777), .ZN(new_n802));
  NAND2_X1  g616(.A1(new_n802), .A2(KEYINPUT118), .ZN(new_n803));
  NAND4_X1  g617(.A1(new_n801), .A2(new_n774), .A3(new_n791), .A4(new_n803), .ZN(new_n804));
  INV_X1    g618(.A(KEYINPUT53), .ZN(new_n805));
  NAND2_X1  g619(.A1(new_n796), .A2(new_n805), .ZN(new_n806));
  AND3_X1   g620(.A1(new_n804), .A2(new_n766), .A3(new_n806), .ZN(new_n807));
  NOR2_X1   g621(.A1(new_n798), .A2(new_n807), .ZN(new_n808));
  INV_X1    g622(.A(KEYINPUT120), .ZN(new_n809));
  NAND2_X1  g623(.A1(new_n673), .A2(new_n467), .ZN(new_n810));
  NOR3_X1   g624(.A1(new_n706), .A2(new_n302), .A3(new_n810), .ZN(new_n811));
  AND2_X1   g625(.A1(new_n751), .A2(new_n811), .ZN(new_n812));
  AND2_X1   g626(.A1(new_n721), .A2(new_n585), .ZN(new_n813));
  NAND2_X1  g627(.A1(new_n812), .A2(new_n813), .ZN(new_n814));
  XNOR2_X1  g628(.A(new_n814), .B(KEYINPUT48), .ZN(new_n815));
  AND3_X1   g629(.A1(new_n656), .A2(new_n585), .A3(new_n662), .ZN(new_n816));
  NAND2_X1  g630(.A1(new_n816), .A2(new_n811), .ZN(new_n817));
  OAI211_X1 g631(.A(new_n815), .B(new_n300), .C1(new_n780), .C2(new_n817), .ZN(new_n818));
  OAI211_X1 g632(.A(new_n760), .B(new_n762), .C1(new_n399), .C2(new_n810), .ZN(new_n819));
  AND2_X1   g633(.A1(new_n694), .A2(new_n303), .ZN(new_n820));
  AND2_X1   g634(.A1(new_n820), .A2(new_n751), .ZN(new_n821));
  AND2_X1   g635(.A1(new_n821), .A2(new_n705), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n819), .A2(new_n822), .ZN(new_n823));
  NAND4_X1  g637(.A1(new_n816), .A2(new_n601), .A3(new_n610), .A4(new_n811), .ZN(new_n824));
  NAND2_X1  g638(.A1(new_n812), .A2(new_n788), .ZN(new_n825));
  INV_X1    g639(.A(KEYINPUT119), .ZN(new_n826));
  XNOR2_X1  g640(.A(new_n825), .B(new_n826), .ZN(new_n827));
  INV_X1    g641(.A(new_n674), .ZN(new_n828));
  NOR2_X1   g642(.A1(new_n652), .A2(new_n394), .ZN(new_n829));
  NAND4_X1  g643(.A1(new_n820), .A2(new_n751), .A3(new_n828), .A4(new_n829), .ZN(new_n830));
  XNOR2_X1  g644(.A(new_n830), .B(KEYINPUT50), .ZN(new_n831));
  INV_X1    g645(.A(new_n831), .ZN(new_n832));
  NAND4_X1  g646(.A1(new_n823), .A2(new_n824), .A3(new_n827), .A4(new_n832), .ZN(new_n833));
  NAND2_X1  g647(.A1(new_n833), .A2(KEYINPUT51), .ZN(new_n834));
  AOI21_X1  g648(.A(new_n831), .B1(new_n819), .B2(new_n822), .ZN(new_n835));
  INV_X1    g649(.A(KEYINPUT51), .ZN(new_n836));
  NAND4_X1  g650(.A1(new_n835), .A2(new_n836), .A3(new_n824), .A4(new_n827), .ZN(new_n837));
  AOI21_X1  g651(.A(new_n818), .B1(new_n834), .B2(new_n837), .ZN(new_n838));
  NAND2_X1  g652(.A1(new_n821), .A2(new_n689), .ZN(new_n839));
  NAND4_X1  g653(.A1(new_n808), .A2(new_n809), .A3(new_n838), .A4(new_n839), .ZN(new_n840));
  AND2_X1   g654(.A1(new_n795), .A2(new_n796), .ZN(new_n841));
  NOR2_X1   g655(.A1(new_n795), .A2(new_n796), .ZN(new_n842));
  OAI21_X1  g656(.A(KEYINPUT54), .B1(new_n841), .B2(new_n842), .ZN(new_n843));
  NAND3_X1  g657(.A1(new_n804), .A2(new_n766), .A3(new_n806), .ZN(new_n844));
  NAND4_X1  g658(.A1(new_n843), .A2(new_n838), .A3(new_n844), .A4(new_n839), .ZN(new_n845));
  NAND2_X1  g659(.A1(new_n845), .A2(KEYINPUT120), .ZN(new_n846));
  NAND2_X1  g660(.A1(new_n299), .A2(new_n195), .ZN(new_n847));
  NAND3_X1  g661(.A1(new_n840), .A2(new_n846), .A3(new_n847), .ZN(new_n848));
  NOR2_X1   g662(.A1(new_n810), .A2(KEYINPUT49), .ZN(new_n849));
  NAND2_X1  g663(.A1(new_n810), .A2(KEYINPUT49), .ZN(new_n850));
  NAND3_X1  g664(.A1(new_n590), .A2(new_n394), .A3(new_n850), .ZN(new_n851));
  NOR2_X1   g665(.A1(new_n851), .A2(new_n749), .ZN(new_n852));
  INV_X1    g666(.A(KEYINPUT115), .ZN(new_n853));
  AOI21_X1  g667(.A(new_n849), .B1(new_n852), .B2(new_n853), .ZN(new_n854));
  NOR2_X1   g668(.A1(new_n663), .A2(new_n652), .ZN(new_n855));
  OAI211_X1 g669(.A(new_n854), .B(new_n855), .C1(new_n853), .C2(new_n852), .ZN(new_n856));
  NAND2_X1  g670(.A1(new_n848), .A2(new_n856), .ZN(G75));
  OAI21_X1  g671(.A(new_n383), .B1(new_n384), .B2(new_n385), .ZN(new_n858));
  XOR2_X1   g672(.A(new_n858), .B(new_n379), .Z(new_n859));
  XNOR2_X1  g673(.A(new_n859), .B(KEYINPUT55), .ZN(new_n860));
  INV_X1    g674(.A(G210), .ZN(new_n861));
  AOI211_X1 g675(.A(new_n861), .B(new_n243), .C1(new_n804), .C2(new_n806), .ZN(new_n862));
  OAI21_X1  g676(.A(new_n860), .B1(new_n862), .B2(KEYINPUT56), .ZN(new_n863));
  NOR2_X1   g677(.A1(new_n195), .A2(G952), .ZN(new_n864));
  INV_X1    g678(.A(new_n864), .ZN(new_n865));
  NAND2_X1  g679(.A1(new_n804), .A2(new_n806), .ZN(new_n866));
  NAND3_X1  g680(.A1(new_n866), .A2(G210), .A3(G902), .ZN(new_n867));
  INV_X1    g681(.A(KEYINPUT56), .ZN(new_n868));
  INV_X1    g682(.A(new_n860), .ZN(new_n869));
  NAND3_X1  g683(.A1(new_n867), .A2(new_n868), .A3(new_n869), .ZN(new_n870));
  NAND3_X1  g684(.A1(new_n863), .A2(new_n865), .A3(new_n870), .ZN(new_n871));
  INV_X1    g685(.A(KEYINPUT121), .ZN(new_n872));
  NAND2_X1  g686(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  NAND4_X1  g687(.A1(new_n863), .A2(KEYINPUT121), .A3(new_n870), .A4(new_n865), .ZN(new_n874));
  NAND2_X1  g688(.A1(new_n873), .A2(new_n874), .ZN(G51));
  XNOR2_X1  g689(.A(new_n468), .B(KEYINPUT57), .ZN(new_n876));
  AOI21_X1  g690(.A(new_n766), .B1(new_n804), .B2(new_n806), .ZN(new_n877));
  OAI21_X1  g691(.A(new_n876), .B1(new_n807), .B2(new_n877), .ZN(new_n878));
  XOR2_X1   g692(.A(new_n672), .B(KEYINPUT122), .Z(new_n879));
  NAND2_X1  g693(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  AOI21_X1  g694(.A(new_n243), .B1(new_n804), .B2(new_n806), .ZN(new_n881));
  INV_X1    g695(.A(new_n735), .ZN(new_n882));
  NAND2_X1  g696(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  AOI21_X1  g697(.A(new_n864), .B1(new_n880), .B2(new_n883), .ZN(G54));
  NAND3_X1  g698(.A1(new_n881), .A2(KEYINPUT58), .A3(G475), .ZN(new_n885));
  INV_X1    g699(.A(new_n247), .ZN(new_n886));
  AND2_X1   g700(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  NOR2_X1   g701(.A1(new_n885), .A2(new_n886), .ZN(new_n888));
  NOR3_X1   g702(.A1(new_n887), .A2(new_n888), .A3(new_n864), .ZN(G60));
  NAND2_X1  g703(.A1(new_n607), .A2(new_n608), .ZN(new_n890));
  OAI21_X1  g704(.A(new_n890), .B1(new_n807), .B2(new_n877), .ZN(new_n891));
  NAND2_X1  g705(.A1(G478), .A2(G902), .ZN(new_n892));
  XOR2_X1   g706(.A(new_n892), .B(KEYINPUT59), .Z(new_n893));
  AOI21_X1  g707(.A(new_n893), .B1(new_n843), .B2(new_n844), .ZN(new_n894));
  OAI221_X1 g708(.A(new_n865), .B1(new_n891), .B2(new_n893), .C1(new_n890), .C2(new_n894), .ZN(new_n895));
  INV_X1    g709(.A(new_n895), .ZN(G63));
  INV_X1    g710(.A(KEYINPUT61), .ZN(new_n897));
  NAND2_X1  g711(.A1(G217), .A2(G902), .ZN(new_n898));
  XNOR2_X1  g712(.A(new_n898), .B(KEYINPUT60), .ZN(new_n899));
  AOI21_X1  g713(.A(new_n899), .B1(new_n804), .B2(new_n806), .ZN(new_n900));
  AOI21_X1  g714(.A(new_n864), .B1(new_n900), .B2(new_n626), .ZN(new_n901));
  INV_X1    g715(.A(KEYINPUT123), .ZN(new_n902));
  AOI21_X1  g716(.A(new_n897), .B1(new_n901), .B2(new_n902), .ZN(new_n903));
  INV_X1    g717(.A(new_n900), .ZN(new_n904));
  NAND2_X1  g718(.A1(new_n904), .A2(new_n577), .ZN(new_n905));
  NAND2_X1  g719(.A1(new_n905), .A2(new_n901), .ZN(new_n906));
  NAND2_X1  g720(.A1(new_n903), .A2(new_n906), .ZN(new_n907));
  OAI211_X1 g721(.A(new_n905), .B(new_n901), .C1(new_n902), .C2(new_n897), .ZN(new_n908));
  AND2_X1   g722(.A1(new_n907), .A2(new_n908), .ZN(G66));
  OAI21_X1  g723(.A(G953), .B1(new_n305), .B2(new_n332), .ZN(new_n910));
  AND3_X1   g724(.A1(new_n783), .A2(new_n588), .A3(new_n633), .ZN(new_n911));
  NAND3_X1  g725(.A1(new_n911), .A2(new_n776), .A3(new_n777), .ZN(new_n912));
  INV_X1    g726(.A(new_n912), .ZN(new_n913));
  OAI21_X1  g727(.A(new_n910), .B1(new_n913), .B2(G953), .ZN(new_n914));
  OAI21_X1  g728(.A(new_n858), .B1(G898), .B2(new_n195), .ZN(new_n915));
  XNOR2_X1  g729(.A(new_n914), .B(new_n915), .ZN(G69));
  NAND3_X1  g730(.A1(new_n664), .A2(new_n646), .A3(new_n767), .ZN(new_n917));
  XNOR2_X1  g731(.A(new_n917), .B(KEYINPUT62), .ZN(new_n918));
  AOI22_X1  g732(.A1(new_n763), .A2(new_n759), .B1(new_n753), .B2(new_n755), .ZN(new_n919));
  INV_X1    g733(.A(KEYINPUT124), .ZN(new_n920));
  OAI211_X1 g734(.A(new_n472), .B(new_n649), .C1(new_n782), .C2(new_n920), .ZN(new_n921));
  AOI21_X1  g735(.A(new_n921), .B1(new_n920), .B2(new_n782), .ZN(new_n922));
  OR2_X1    g736(.A1(new_n586), .A2(new_n587), .ZN(new_n923));
  NAND3_X1  g737(.A1(new_n922), .A2(new_n923), .A3(new_n705), .ZN(new_n924));
  NAND2_X1  g738(.A1(new_n919), .A2(new_n924), .ZN(new_n925));
  OAI21_X1  g739(.A(new_n195), .B1(new_n918), .B2(new_n925), .ZN(new_n926));
  INV_X1    g740(.A(new_n499), .ZN(new_n927));
  MUX2_X1   g741(.A(new_n485), .B(new_n927), .S(KEYINPUT30), .Z(new_n928));
  XOR2_X1   g742(.A(new_n928), .B(new_n235), .Z(new_n929));
  NAND2_X1  g743(.A1(new_n926), .A2(new_n929), .ZN(new_n930));
  INV_X1    g744(.A(new_n929), .ZN(new_n931));
  NAND2_X1  g745(.A1(G900), .A2(G953), .ZN(new_n932));
  NAND4_X1  g746(.A1(new_n743), .A2(new_n649), .A3(new_n695), .A4(new_n813), .ZN(new_n933));
  AND3_X1   g747(.A1(new_n933), .A2(new_n646), .A3(new_n767), .ZN(new_n934));
  NAND4_X1  g748(.A1(new_n919), .A2(new_n725), .A3(new_n728), .A4(new_n934), .ZN(new_n935));
  OAI211_X1 g749(.A(new_n931), .B(new_n932), .C1(new_n935), .C2(G953), .ZN(new_n936));
  NAND2_X1  g750(.A1(new_n930), .A2(new_n936), .ZN(new_n937));
  NAND2_X1  g751(.A1(new_n937), .A2(KEYINPUT125), .ZN(new_n938));
  AOI21_X1  g752(.A(new_n195), .B1(G227), .B2(G900), .ZN(new_n939));
  INV_X1    g753(.A(KEYINPUT125), .ZN(new_n940));
  NAND3_X1  g754(.A1(new_n930), .A2(new_n936), .A3(new_n940), .ZN(new_n941));
  AND3_X1   g755(.A1(new_n938), .A2(new_n939), .A3(new_n941), .ZN(new_n942));
  AOI21_X1  g756(.A(new_n939), .B1(new_n938), .B2(new_n941), .ZN(new_n943));
  NOR2_X1   g757(.A1(new_n942), .A2(new_n943), .ZN(G72));
  XNOR2_X1  g758(.A(KEYINPUT126), .B(KEYINPUT63), .ZN(new_n945));
  NAND2_X1  g759(.A1(G472), .A2(G902), .ZN(new_n946));
  XNOR2_X1  g760(.A(new_n945), .B(new_n946), .ZN(new_n947));
  INV_X1    g761(.A(new_n517), .ZN(new_n948));
  NOR2_X1   g762(.A1(new_n948), .A2(new_n492), .ZN(new_n949));
  OAI221_X1 g763(.A(new_n947), .B1(new_n949), .B2(new_n658), .C1(new_n841), .C2(new_n842), .ZN(new_n950));
  OR2_X1    g764(.A1(new_n918), .A2(new_n925), .ZN(new_n951));
  OAI21_X1  g765(.A(new_n947), .B1(new_n951), .B2(new_n912), .ZN(new_n952));
  NAND3_X1  g766(.A1(new_n952), .A2(new_n492), .A3(new_n517), .ZN(new_n953));
  OAI21_X1  g767(.A(new_n947), .B1(new_n935), .B2(new_n912), .ZN(new_n954));
  NAND3_X1  g768(.A1(new_n954), .A2(new_n505), .A3(new_n948), .ZN(new_n955));
  AND3_X1   g769(.A1(new_n955), .A2(KEYINPUT127), .A3(new_n865), .ZN(new_n956));
  AOI21_X1  g770(.A(KEYINPUT127), .B1(new_n955), .B2(new_n865), .ZN(new_n957));
  OAI211_X1 g771(.A(new_n950), .B(new_n953), .C1(new_n956), .C2(new_n957), .ZN(new_n958));
  INV_X1    g772(.A(new_n958), .ZN(G57));
endmodule


