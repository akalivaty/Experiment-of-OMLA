//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 1 1 1 1 1 0 0 0 1 1 1 1 0 1 1 0 1 0 1 1 1 0 0 0 1 0 1 1 1 1 0 0 1 0 0 1 1 0 0 0 1 0 1 1 0 0 1 0 1 1 1 0 1 1 0 1 0 0 0 1 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:31:07 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n443, new_n444, new_n445, new_n450, new_n454, new_n455,
    new_n456, new_n457, new_n460, new_n461, new_n462, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n525,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n531, new_n532,
    new_n533, new_n534, new_n535, new_n536, new_n537, new_n538, new_n539,
    new_n541, new_n542, new_n543, new_n544, new_n545, new_n546, new_n547,
    new_n548, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n558, new_n560, new_n561, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n580, new_n581, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n597, new_n598,
    new_n599, new_n600, new_n601, new_n602, new_n603, new_n604, new_n605,
    new_n606, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n637,
    new_n640, new_n642, new_n643, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n692, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n845, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1187, new_n1188, new_n1189, new_n1190,
    new_n1191;
  BUF_X1    g000(.A(G452), .Z(G350));
  XNOR2_X1  g001(.A(KEYINPUT64), .B(G452), .ZN(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  XNOR2_X1  g007(.A(KEYINPUT65), .B(G2066), .ZN(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  XOR2_X1   g009(.A(KEYINPUT66), .B(G132), .Z(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  INV_X1    g016(.A(G2072), .ZN(new_n442));
  INV_X1    g017(.A(G2078), .ZN(new_n443));
  NOR2_X1   g018(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  NAND3_X1  g019(.A1(new_n444), .A2(G2084), .A3(G2090), .ZN(new_n445));
  XNOR2_X1  g020(.A(new_n445), .B(KEYINPUT67), .ZN(G158));
  NAND3_X1  g021(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g022(.A(G452), .Z(G391));
  AND2_X1   g023(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g024(.A1(G7), .A2(G661), .ZN(new_n450));
  XOR2_X1   g025(.A(new_n450), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g026(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g027(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g028(.A1(G219), .A2(G220), .A3(G218), .A4(G221), .ZN(new_n454));
  XOR2_X1   g029(.A(new_n454), .B(KEYINPUT2), .Z(new_n455));
  NOR4_X1   g030(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n456));
  INV_X1    g031(.A(new_n456), .ZN(new_n457));
  NOR2_X1   g032(.A1(new_n455), .A2(new_n457), .ZN(G325));
  INV_X1    g033(.A(G325), .ZN(G261));
  NAND2_X1  g034(.A1(new_n455), .A2(G2106), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n457), .A2(G567), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  INV_X1    g037(.A(new_n462), .ZN(G319));
  XNOR2_X1  g038(.A(KEYINPUT3), .B(G2104), .ZN(new_n464));
  INV_X1    g039(.A(G2105), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  INV_X1    g041(.A(new_n466), .ZN(new_n467));
  INV_X1    g042(.A(G2104), .ZN(new_n468));
  NOR2_X1   g043(.A1(new_n468), .A2(G2105), .ZN(new_n469));
  AOI22_X1  g044(.A1(new_n467), .A2(G137), .B1(G101), .B2(new_n469), .ZN(new_n470));
  INV_X1    g045(.A(new_n470), .ZN(new_n471));
  AOI22_X1  g046(.A1(new_n464), .A2(G125), .B1(G113), .B2(G2104), .ZN(new_n472));
  OAI21_X1  g047(.A(KEYINPUT68), .B1(new_n472), .B2(new_n465), .ZN(new_n473));
  NAND2_X1  g048(.A1(G113), .A2(G2104), .ZN(new_n474));
  AND2_X1   g049(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n475));
  NOR2_X1   g050(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n476));
  NOR2_X1   g051(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  INV_X1    g052(.A(G125), .ZN(new_n478));
  OAI21_X1  g053(.A(new_n474), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  INV_X1    g054(.A(KEYINPUT68), .ZN(new_n480));
  NAND3_X1  g055(.A1(new_n479), .A2(new_n480), .A3(G2105), .ZN(new_n481));
  AOI21_X1  g056(.A(new_n471), .B1(new_n473), .B2(new_n481), .ZN(G160));
  OR2_X1    g057(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n483));
  NAND2_X1  g058(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n484));
  AOI21_X1  g059(.A(new_n465), .B1(new_n483), .B2(new_n484), .ZN(new_n485));
  NAND2_X1  g060(.A1(new_n485), .A2(G124), .ZN(new_n486));
  XNOR2_X1  g061(.A(new_n486), .B(KEYINPUT69), .ZN(new_n487));
  NAND2_X1  g062(.A1(new_n467), .A2(G136), .ZN(new_n488));
  NOR2_X1   g063(.A1(G100), .A2(G2105), .ZN(new_n489));
  XNOR2_X1  g064(.A(new_n489), .B(KEYINPUT70), .ZN(new_n490));
  OAI21_X1  g065(.A(G2104), .B1(new_n465), .B2(G112), .ZN(new_n491));
  OAI211_X1 g066(.A(new_n487), .B(new_n488), .C1(new_n490), .C2(new_n491), .ZN(new_n492));
  XNOR2_X1  g067(.A(new_n492), .B(KEYINPUT71), .ZN(G162));
  OAI211_X1 g068(.A(G126), .B(G2105), .C1(new_n475), .C2(new_n476), .ZN(new_n494));
  OR2_X1    g069(.A1(G102), .A2(G2105), .ZN(new_n495));
  INV_X1    g070(.A(G114), .ZN(new_n496));
  NAND2_X1  g071(.A1(new_n496), .A2(G2105), .ZN(new_n497));
  NAND3_X1  g072(.A1(new_n495), .A2(new_n497), .A3(G2104), .ZN(new_n498));
  NAND2_X1  g073(.A1(new_n494), .A2(new_n498), .ZN(new_n499));
  INV_X1    g074(.A(G138), .ZN(new_n500));
  NOR2_X1   g075(.A1(new_n500), .A2(G2105), .ZN(new_n501));
  OAI21_X1  g076(.A(new_n501), .B1(new_n475), .B2(new_n476), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n502), .A2(KEYINPUT4), .ZN(new_n503));
  INV_X1    g078(.A(KEYINPUT4), .ZN(new_n504));
  OAI211_X1 g079(.A(new_n501), .B(new_n504), .C1(new_n476), .C2(new_n475), .ZN(new_n505));
  AOI21_X1  g080(.A(new_n499), .B1(new_n503), .B2(new_n505), .ZN(G164));
  XNOR2_X1  g081(.A(KEYINPUT5), .B(G543), .ZN(new_n507));
  XNOR2_X1  g082(.A(KEYINPUT6), .B(G651), .ZN(new_n508));
  AND2_X1   g083(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  XOR2_X1   g084(.A(KEYINPUT72), .B(G88), .Z(new_n510));
  INV_X1    g085(.A(G543), .ZN(new_n511));
  OR2_X1    g086(.A1(KEYINPUT6), .A2(G651), .ZN(new_n512));
  NAND2_X1  g087(.A1(KEYINPUT6), .A2(G651), .ZN(new_n513));
  AOI21_X1  g088(.A(new_n511), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  AOI22_X1  g089(.A1(new_n509), .A2(new_n510), .B1(G50), .B2(new_n514), .ZN(new_n515));
  INV_X1    g090(.A(new_n515), .ZN(new_n516));
  AOI22_X1  g091(.A1(new_n507), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n517));
  INV_X1    g092(.A(G651), .ZN(new_n518));
  OR2_X1    g093(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  INV_X1    g094(.A(KEYINPUT73), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  NOR2_X1   g096(.A1(new_n517), .A2(new_n518), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n522), .A2(KEYINPUT73), .ZN(new_n523));
  AOI21_X1  g098(.A(new_n516), .B1(new_n521), .B2(new_n523), .ZN(G166));
  NAND3_X1  g099(.A1(new_n507), .A2(G63), .A3(G651), .ZN(new_n525));
  NAND2_X1  g100(.A1(new_n508), .A2(G543), .ZN(new_n526));
  INV_X1    g101(.A(G51), .ZN(new_n527));
  OAI21_X1  g102(.A(new_n525), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  NAND2_X1  g103(.A1(new_n528), .A2(KEYINPUT74), .ZN(new_n529));
  INV_X1    g104(.A(KEYINPUT74), .ZN(new_n530));
  OAI211_X1 g105(.A(new_n525), .B(new_n530), .C1(new_n526), .C2(new_n527), .ZN(new_n531));
  NAND3_X1  g106(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n532));
  NAND2_X1  g107(.A1(new_n532), .A2(KEYINPUT7), .ZN(new_n533));
  OR2_X1    g108(.A1(new_n532), .A2(KEYINPUT7), .ZN(new_n534));
  AOI22_X1  g109(.A1(new_n509), .A2(G89), .B1(new_n533), .B2(new_n534), .ZN(new_n535));
  NAND3_X1  g110(.A1(new_n529), .A2(new_n531), .A3(new_n535), .ZN(new_n536));
  INV_X1    g111(.A(KEYINPUT75), .ZN(new_n537));
  NAND2_X1  g112(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  NAND4_X1  g113(.A1(new_n529), .A2(new_n535), .A3(KEYINPUT75), .A4(new_n531), .ZN(new_n539));
  NAND2_X1  g114(.A1(new_n538), .A2(new_n539), .ZN(G168));
  AOI22_X1  g115(.A1(new_n507), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n541));
  NOR2_X1   g116(.A1(new_n541), .A2(new_n518), .ZN(new_n542));
  NAND2_X1  g117(.A1(new_n514), .A2(G52), .ZN(new_n543));
  NAND3_X1  g118(.A1(new_n507), .A2(new_n508), .A3(G90), .ZN(new_n544));
  NAND2_X1  g119(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  INV_X1    g120(.A(KEYINPUT76), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  NAND3_X1  g122(.A1(new_n543), .A2(new_n544), .A3(KEYINPUT76), .ZN(new_n548));
  AOI21_X1  g123(.A(new_n542), .B1(new_n547), .B2(new_n548), .ZN(G171));
  NAND2_X1  g124(.A1(new_n507), .A2(new_n508), .ZN(new_n550));
  INV_X1    g125(.A(G81), .ZN(new_n551));
  INV_X1    g126(.A(G43), .ZN(new_n552));
  OAI22_X1  g127(.A1(new_n550), .A2(new_n551), .B1(new_n526), .B2(new_n552), .ZN(new_n553));
  AOI22_X1  g128(.A1(new_n507), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n554));
  NOR2_X1   g129(.A1(new_n554), .A2(new_n518), .ZN(new_n555));
  NOR2_X1   g130(.A1(new_n553), .A2(new_n555), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n556), .A2(G860), .ZN(G153));
  NAND4_X1  g132(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(new_n558));
  XNOR2_X1  g133(.A(new_n558), .B(KEYINPUT77), .ZN(G176));
  NAND2_X1  g134(.A1(G1), .A2(G3), .ZN(new_n560));
  XNOR2_X1  g135(.A(new_n560), .B(KEYINPUT8), .ZN(new_n561));
  NAND4_X1  g136(.A1(G319), .A2(G483), .A3(G661), .A4(new_n561), .ZN(G188));
  INV_X1    g137(.A(new_n513), .ZN(new_n563));
  NOR2_X1   g138(.A1(KEYINPUT6), .A2(G651), .ZN(new_n564));
  OAI211_X1 g139(.A(G53), .B(G543), .C1(new_n563), .C2(new_n564), .ZN(new_n565));
  NAND2_X1  g140(.A1(new_n565), .A2(KEYINPUT78), .ZN(new_n566));
  NAND3_X1  g141(.A1(new_n507), .A2(new_n508), .A3(G91), .ZN(new_n567));
  AOI22_X1  g142(.A1(new_n507), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n568));
  OAI211_X1 g143(.A(new_n566), .B(new_n567), .C1(new_n568), .C2(new_n518), .ZN(new_n569));
  INV_X1    g144(.A(new_n569), .ZN(new_n570));
  INV_X1    g145(.A(KEYINPUT9), .ZN(new_n571));
  INV_X1    g146(.A(KEYINPUT79), .ZN(new_n572));
  OAI21_X1  g147(.A(new_n571), .B1(new_n565), .B2(new_n572), .ZN(new_n573));
  NOR2_X1   g148(.A1(new_n571), .A2(KEYINPUT78), .ZN(new_n574));
  NAND4_X1  g149(.A1(new_n514), .A2(KEYINPUT79), .A3(G53), .A4(new_n574), .ZN(new_n575));
  AND2_X1   g150(.A1(new_n573), .A2(new_n575), .ZN(new_n576));
  NAND2_X1  g151(.A1(new_n570), .A2(new_n576), .ZN(G299));
  INV_X1    g152(.A(G171), .ZN(G301));
  INV_X1    g153(.A(G168), .ZN(G286));
  INV_X1    g154(.A(new_n523), .ZN(new_n580));
  NOR2_X1   g155(.A1(new_n522), .A2(KEYINPUT73), .ZN(new_n581));
  OAI21_X1  g156(.A(new_n515), .B1(new_n580), .B2(new_n581), .ZN(G303));
  OR2_X1    g157(.A1(new_n507), .A2(G74), .ZN(new_n583));
  AOI22_X1  g158(.A1(G651), .A2(new_n583), .B1(new_n509), .B2(G87), .ZN(new_n584));
  NAND3_X1  g159(.A1(new_n514), .A2(KEYINPUT80), .A3(G49), .ZN(new_n585));
  INV_X1    g160(.A(KEYINPUT80), .ZN(new_n586));
  INV_X1    g161(.A(G49), .ZN(new_n587));
  OAI21_X1  g162(.A(new_n586), .B1(new_n526), .B2(new_n587), .ZN(new_n588));
  NAND3_X1  g163(.A1(new_n584), .A2(new_n585), .A3(new_n588), .ZN(G288));
  INV_X1    g164(.A(G86), .ZN(new_n590));
  INV_X1    g165(.A(G48), .ZN(new_n591));
  OAI22_X1  g166(.A1(new_n550), .A2(new_n590), .B1(new_n526), .B2(new_n591), .ZN(new_n592));
  NAND2_X1  g167(.A1(new_n507), .A2(G61), .ZN(new_n593));
  NAND2_X1  g168(.A1(G73), .A2(G543), .ZN(new_n594));
  AOI21_X1  g169(.A(new_n518), .B1(new_n593), .B2(new_n594), .ZN(new_n595));
  OR2_X1    g170(.A1(new_n595), .A2(KEYINPUT81), .ZN(new_n596));
  NAND2_X1  g171(.A1(new_n595), .A2(KEYINPUT81), .ZN(new_n597));
  AOI21_X1  g172(.A(new_n592), .B1(new_n596), .B2(new_n597), .ZN(new_n598));
  NOR2_X1   g173(.A1(new_n598), .A2(KEYINPUT82), .ZN(new_n599));
  INV_X1    g174(.A(new_n592), .ZN(new_n600));
  NOR2_X1   g175(.A1(new_n595), .A2(KEYINPUT81), .ZN(new_n601));
  INV_X1    g176(.A(KEYINPUT81), .ZN(new_n602));
  AOI211_X1 g177(.A(new_n602), .B(new_n518), .C1(new_n593), .C2(new_n594), .ZN(new_n603));
  OAI21_X1  g178(.A(new_n600), .B1(new_n601), .B2(new_n603), .ZN(new_n604));
  INV_X1    g179(.A(KEYINPUT82), .ZN(new_n605));
  NOR2_X1   g180(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  NOR2_X1   g181(.A1(new_n599), .A2(new_n606), .ZN(G305));
  INV_X1    g182(.A(G85), .ZN(new_n608));
  INV_X1    g183(.A(G47), .ZN(new_n609));
  OAI22_X1  g184(.A1(new_n550), .A2(new_n608), .B1(new_n526), .B2(new_n609), .ZN(new_n610));
  AOI22_X1  g185(.A1(new_n507), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n611));
  NOR2_X1   g186(.A1(new_n611), .A2(new_n518), .ZN(new_n612));
  NOR2_X1   g187(.A1(new_n610), .A2(new_n612), .ZN(new_n613));
  INV_X1    g188(.A(new_n613), .ZN(G290));
  INV_X1    g189(.A(G868), .ZN(new_n615));
  NOR2_X1   g190(.A1(G171), .A2(new_n615), .ZN(new_n616));
  XNOR2_X1  g191(.A(new_n616), .B(KEYINPUT83), .ZN(new_n617));
  INV_X1    g192(.A(G92), .ZN(new_n618));
  XOR2_X1   g193(.A(KEYINPUT84), .B(KEYINPUT10), .Z(new_n619));
  OR3_X1    g194(.A1(new_n550), .A2(new_n618), .A3(new_n619), .ZN(new_n620));
  OAI21_X1  g195(.A(new_n619), .B1(new_n550), .B2(new_n618), .ZN(new_n621));
  AOI22_X1  g196(.A1(new_n620), .A2(new_n621), .B1(G54), .B2(new_n514), .ZN(new_n622));
  INV_X1    g197(.A(KEYINPUT85), .ZN(new_n623));
  OR2_X1    g198(.A1(new_n623), .A2(G66), .ZN(new_n624));
  NAND2_X1  g199(.A1(new_n623), .A2(G66), .ZN(new_n625));
  NAND3_X1  g200(.A1(new_n507), .A2(new_n624), .A3(new_n625), .ZN(new_n626));
  INV_X1    g201(.A(G79), .ZN(new_n627));
  OAI21_X1  g202(.A(new_n626), .B1(new_n627), .B2(new_n511), .ZN(new_n628));
  INV_X1    g203(.A(KEYINPUT86), .ZN(new_n629));
  NAND2_X1  g204(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  OAI211_X1 g205(.A(new_n626), .B(KEYINPUT86), .C1(new_n627), .C2(new_n511), .ZN(new_n631));
  NAND3_X1  g206(.A1(new_n630), .A2(G651), .A3(new_n631), .ZN(new_n632));
  NAND2_X1  g207(.A1(new_n622), .A2(new_n632), .ZN(new_n633));
  XNOR2_X1  g208(.A(new_n633), .B(KEYINPUT87), .ZN(new_n634));
  OAI21_X1  g209(.A(new_n617), .B1(new_n634), .B2(G868), .ZN(G284));
  OAI21_X1  g210(.A(new_n617), .B1(new_n634), .B2(G868), .ZN(G321));
  NOR2_X1   g211(.A1(G299), .A2(G868), .ZN(new_n637));
  AOI21_X1  g212(.A(new_n637), .B1(G168), .B2(G868), .ZN(G297));
  AOI21_X1  g213(.A(new_n637), .B1(G168), .B2(G868), .ZN(G280));
  XNOR2_X1  g214(.A(KEYINPUT88), .B(G559), .ZN(new_n640));
  OAI21_X1  g215(.A(new_n634), .B1(G860), .B2(new_n640), .ZN(G148));
  NAND2_X1  g216(.A1(new_n634), .A2(new_n640), .ZN(new_n642));
  NAND2_X1  g217(.A1(new_n642), .A2(G868), .ZN(new_n643));
  OAI21_X1  g218(.A(new_n643), .B1(G868), .B2(new_n556), .ZN(G323));
  XNOR2_X1  g219(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g220(.A1(new_n464), .A2(new_n469), .ZN(new_n646));
  XOR2_X1   g221(.A(KEYINPUT89), .B(KEYINPUT12), .Z(new_n647));
  XNOR2_X1  g222(.A(new_n646), .B(new_n647), .ZN(new_n648));
  XNOR2_X1  g223(.A(new_n648), .B(KEYINPUT13), .ZN(new_n649));
  INV_X1    g224(.A(G2100), .ZN(new_n650));
  OR2_X1    g225(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  NAND2_X1  g226(.A1(new_n649), .A2(new_n650), .ZN(new_n652));
  NAND2_X1  g227(.A1(new_n485), .A2(G123), .ZN(new_n653));
  OR2_X1    g228(.A1(G99), .A2(G2105), .ZN(new_n654));
  OAI211_X1 g229(.A(new_n654), .B(G2104), .C1(G111), .C2(new_n465), .ZN(new_n655));
  INV_X1    g230(.A(G135), .ZN(new_n656));
  OAI211_X1 g231(.A(new_n653), .B(new_n655), .C1(new_n656), .C2(new_n466), .ZN(new_n657));
  XOR2_X1   g232(.A(new_n657), .B(G2096), .Z(new_n658));
  NAND3_X1  g233(.A1(new_n651), .A2(new_n652), .A3(new_n658), .ZN(G156));
  XNOR2_X1  g234(.A(G2427), .B(G2438), .ZN(new_n660));
  XNOR2_X1  g235(.A(new_n660), .B(G2430), .ZN(new_n661));
  XNOR2_X1  g236(.A(KEYINPUT15), .B(G2435), .ZN(new_n662));
  OR2_X1    g237(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  NAND2_X1  g238(.A1(new_n661), .A2(new_n662), .ZN(new_n664));
  NAND3_X1  g239(.A1(new_n663), .A2(KEYINPUT14), .A3(new_n664), .ZN(new_n665));
  XOR2_X1   g240(.A(KEYINPUT90), .B(KEYINPUT16), .Z(new_n666));
  XNOR2_X1  g241(.A(new_n665), .B(new_n666), .ZN(new_n667));
  XOR2_X1   g242(.A(G2451), .B(G2454), .Z(new_n668));
  XNOR2_X1  g243(.A(G2443), .B(G2446), .ZN(new_n669));
  XNOR2_X1  g244(.A(new_n668), .B(new_n669), .ZN(new_n670));
  XNOR2_X1  g245(.A(new_n667), .B(new_n670), .ZN(new_n671));
  XNOR2_X1  g246(.A(G1341), .B(G1348), .ZN(new_n672));
  NAND2_X1  g247(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  INV_X1    g248(.A(KEYINPUT91), .ZN(new_n674));
  XNOR2_X1  g249(.A(new_n673), .B(new_n674), .ZN(new_n675));
  OR2_X1    g250(.A1(new_n671), .A2(new_n672), .ZN(new_n676));
  AND2_X1   g251(.A1(new_n676), .A2(G14), .ZN(new_n677));
  AND2_X1   g252(.A1(new_n675), .A2(new_n677), .ZN(G401));
  XOR2_X1   g253(.A(G2084), .B(G2090), .Z(new_n679));
  XNOR2_X1  g254(.A(G2067), .B(G2678), .ZN(new_n680));
  XOR2_X1   g255(.A(new_n680), .B(KEYINPUT92), .Z(new_n681));
  NOR2_X1   g256(.A1(G2072), .A2(G2078), .ZN(new_n682));
  NOR2_X1   g257(.A1(new_n444), .A2(new_n682), .ZN(new_n683));
  AOI21_X1  g258(.A(new_n679), .B1(new_n681), .B2(new_n683), .ZN(new_n684));
  XNOR2_X1  g259(.A(new_n683), .B(KEYINPUT17), .ZN(new_n685));
  OAI21_X1  g260(.A(new_n684), .B1(new_n681), .B2(new_n685), .ZN(new_n686));
  OAI211_X1 g261(.A(new_n679), .B(new_n680), .C1(new_n444), .C2(new_n682), .ZN(new_n687));
  XOR2_X1   g262(.A(new_n687), .B(KEYINPUT18), .Z(new_n688));
  NAND3_X1  g263(.A1(new_n685), .A2(new_n681), .A3(new_n679), .ZN(new_n689));
  NAND3_X1  g264(.A1(new_n686), .A2(new_n688), .A3(new_n689), .ZN(new_n690));
  XNOR2_X1  g265(.A(new_n690), .B(new_n650), .ZN(new_n691));
  XNOR2_X1  g266(.A(KEYINPUT93), .B(G2096), .ZN(new_n692));
  XNOR2_X1  g267(.A(new_n691), .B(new_n692), .ZN(G227));
  XNOR2_X1  g268(.A(G1971), .B(G1976), .ZN(new_n694));
  INV_X1    g269(.A(KEYINPUT19), .ZN(new_n695));
  XNOR2_X1  g270(.A(new_n694), .B(new_n695), .ZN(new_n696));
  XOR2_X1   g271(.A(G1956), .B(G2474), .Z(new_n697));
  XOR2_X1   g272(.A(G1961), .B(G1966), .Z(new_n698));
  NOR2_X1   g273(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  AND2_X1   g274(.A1(new_n696), .A2(new_n699), .ZN(new_n700));
  AND2_X1   g275(.A1(new_n697), .A2(new_n698), .ZN(new_n701));
  NOR3_X1   g276(.A1(new_n696), .A2(new_n701), .A3(new_n699), .ZN(new_n702));
  NAND2_X1  g277(.A1(new_n696), .A2(new_n701), .ZN(new_n703));
  XOR2_X1   g278(.A(KEYINPUT94), .B(KEYINPUT20), .Z(new_n704));
  AOI211_X1 g279(.A(new_n700), .B(new_n702), .C1(new_n703), .C2(new_n704), .ZN(new_n705));
  OAI21_X1  g280(.A(new_n705), .B1(new_n703), .B2(new_n704), .ZN(new_n706));
  XNOR2_X1  g281(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n707));
  XNOR2_X1  g282(.A(new_n706), .B(new_n707), .ZN(new_n708));
  XNOR2_X1  g283(.A(G1991), .B(G1996), .ZN(new_n709));
  AND2_X1   g284(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  NOR2_X1   g285(.A1(new_n708), .A2(new_n709), .ZN(new_n711));
  XNOR2_X1  g286(.A(G1981), .B(G1986), .ZN(new_n712));
  INV_X1    g287(.A(new_n712), .ZN(new_n713));
  OR3_X1    g288(.A1(new_n710), .A2(new_n711), .A3(new_n713), .ZN(new_n714));
  OAI21_X1  g289(.A(new_n713), .B1(new_n710), .B2(new_n711), .ZN(new_n715));
  AND2_X1   g290(.A1(new_n714), .A2(new_n715), .ZN(G229));
  NOR2_X1   g291(.A1(G29), .A2(G35), .ZN(new_n717));
  AOI21_X1  g292(.A(new_n717), .B1(G162), .B2(G29), .ZN(new_n718));
  XNOR2_X1  g293(.A(new_n718), .B(KEYINPUT29), .ZN(new_n719));
  XNOR2_X1  g294(.A(new_n719), .B(G2090), .ZN(new_n720));
  INV_X1    g295(.A(G16), .ZN(new_n721));
  NAND2_X1  g296(.A1(new_n721), .A2(G21), .ZN(new_n722));
  OAI21_X1  g297(.A(new_n722), .B1(G168), .B2(new_n721), .ZN(new_n723));
  NAND2_X1  g298(.A1(new_n723), .A2(G1966), .ZN(new_n724));
  XNOR2_X1  g299(.A(new_n724), .B(KEYINPUT100), .ZN(new_n725));
  NOR2_X1   g300(.A1(new_n720), .A2(new_n725), .ZN(new_n726));
  XNOR2_X1  g301(.A(KEYINPUT30), .B(G28), .ZN(new_n727));
  INV_X1    g302(.A(G29), .ZN(new_n728));
  OR2_X1    g303(.A1(KEYINPUT31), .A2(G11), .ZN(new_n729));
  NAND2_X1  g304(.A1(KEYINPUT31), .A2(G11), .ZN(new_n730));
  AOI22_X1  g305(.A1(new_n727), .A2(new_n728), .B1(new_n729), .B2(new_n730), .ZN(new_n731));
  NAND2_X1  g306(.A1(G164), .A2(G29), .ZN(new_n732));
  OAI21_X1  g307(.A(new_n732), .B1(G27), .B2(G29), .ZN(new_n733));
  OAI221_X1 g308(.A(new_n731), .B1(new_n728), .B2(new_n657), .C1(new_n733), .C2(new_n443), .ZN(new_n734));
  AND2_X1   g309(.A1(new_n728), .A2(G33), .ZN(new_n735));
  NAND3_X1  g310(.A1(new_n465), .A2(G103), .A3(G2104), .ZN(new_n736));
  INV_X1    g311(.A(KEYINPUT25), .ZN(new_n737));
  XNOR2_X1  g312(.A(new_n736), .B(new_n737), .ZN(new_n738));
  INV_X1    g313(.A(G139), .ZN(new_n739));
  OAI21_X1  g314(.A(new_n738), .B1(new_n739), .B2(new_n466), .ZN(new_n740));
  NAND2_X1  g315(.A1(new_n464), .A2(G127), .ZN(new_n741));
  NAND2_X1  g316(.A1(G115), .A2(G2104), .ZN(new_n742));
  AOI21_X1  g317(.A(new_n465), .B1(new_n741), .B2(new_n742), .ZN(new_n743));
  NOR2_X1   g318(.A1(new_n740), .A2(new_n743), .ZN(new_n744));
  XNOR2_X1  g319(.A(new_n744), .B(KEYINPUT97), .ZN(new_n745));
  AOI21_X1  g320(.A(new_n735), .B1(new_n745), .B2(G29), .ZN(new_n746));
  NOR2_X1   g321(.A1(new_n746), .A2(new_n442), .ZN(new_n747));
  AOI211_X1 g322(.A(new_n734), .B(new_n747), .C1(new_n443), .C2(new_n733), .ZN(new_n748));
  NAND2_X1  g323(.A1(G160), .A2(G29), .ZN(new_n749));
  INV_X1    g324(.A(KEYINPUT24), .ZN(new_n750));
  OAI21_X1  g325(.A(new_n728), .B1(new_n750), .B2(G34), .ZN(new_n751));
  AND2_X1   g326(.A1(new_n751), .A2(KEYINPUT98), .ZN(new_n752));
  NAND2_X1  g327(.A1(new_n750), .A2(G34), .ZN(new_n753));
  OAI21_X1  g328(.A(new_n753), .B1(new_n751), .B2(KEYINPUT98), .ZN(new_n754));
  OAI21_X1  g329(.A(new_n749), .B1(new_n752), .B2(new_n754), .ZN(new_n755));
  INV_X1    g330(.A(G2084), .ZN(new_n756));
  AOI22_X1  g331(.A1(new_n442), .A2(new_n746), .B1(new_n755), .B2(new_n756), .ZN(new_n757));
  NAND2_X1  g332(.A1(new_n721), .A2(G20), .ZN(new_n758));
  XOR2_X1   g333(.A(new_n758), .B(KEYINPUT23), .Z(new_n759));
  AOI21_X1  g334(.A(new_n759), .B1(G299), .B2(G16), .ZN(new_n760));
  XNOR2_X1  g335(.A(new_n760), .B(G1956), .ZN(new_n761));
  NAND2_X1  g336(.A1(new_n728), .A2(G32), .ZN(new_n762));
  AOI22_X1  g337(.A1(new_n467), .A2(G141), .B1(G105), .B2(new_n469), .ZN(new_n763));
  NAND2_X1  g338(.A1(new_n485), .A2(G129), .ZN(new_n764));
  NAND3_X1  g339(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n765));
  XOR2_X1   g340(.A(new_n765), .B(KEYINPUT26), .Z(new_n766));
  AND3_X1   g341(.A1(new_n763), .A2(new_n764), .A3(new_n766), .ZN(new_n767));
  OAI21_X1  g342(.A(new_n762), .B1(new_n767), .B2(new_n728), .ZN(new_n768));
  XNOR2_X1  g343(.A(new_n768), .B(KEYINPUT27), .ZN(new_n769));
  XNOR2_X1  g344(.A(new_n769), .B(G1996), .ZN(new_n770));
  NAND4_X1  g345(.A1(new_n748), .A2(new_n757), .A3(new_n761), .A4(new_n770), .ZN(new_n771));
  NOR2_X1   g346(.A1(new_n755), .A2(new_n756), .ZN(new_n772));
  XOR2_X1   g347(.A(new_n772), .B(KEYINPUT99), .Z(new_n773));
  NAND2_X1  g348(.A1(new_n721), .A2(G5), .ZN(new_n774));
  OAI21_X1  g349(.A(new_n774), .B1(G171), .B2(new_n721), .ZN(new_n775));
  XOR2_X1   g350(.A(new_n775), .B(KEYINPUT101), .Z(new_n776));
  INV_X1    g351(.A(G1961), .ZN(new_n777));
  AND2_X1   g352(.A1(new_n776), .A2(new_n777), .ZN(new_n778));
  OAI22_X1  g353(.A1(new_n776), .A2(new_n777), .B1(G1966), .B2(new_n723), .ZN(new_n779));
  NOR4_X1   g354(.A1(new_n771), .A2(new_n773), .A3(new_n778), .A4(new_n779), .ZN(new_n780));
  NOR2_X1   g355(.A1(new_n634), .A2(new_n721), .ZN(new_n781));
  AND2_X1   g356(.A1(new_n721), .A2(G4), .ZN(new_n782));
  OR3_X1    g357(.A1(new_n781), .A2(G1348), .A3(new_n782), .ZN(new_n783));
  OAI21_X1  g358(.A(G1348), .B1(new_n781), .B2(new_n782), .ZN(new_n784));
  NAND2_X1  g359(.A1(new_n721), .A2(G19), .ZN(new_n785));
  OAI21_X1  g360(.A(new_n785), .B1(new_n556), .B2(new_n721), .ZN(new_n786));
  XOR2_X1   g361(.A(new_n786), .B(G1341), .Z(new_n787));
  NAND2_X1  g362(.A1(new_n728), .A2(G26), .ZN(new_n788));
  XNOR2_X1  g363(.A(new_n788), .B(KEYINPUT28), .ZN(new_n789));
  NAND2_X1  g364(.A1(new_n467), .A2(G140), .ZN(new_n790));
  NAND2_X1  g365(.A1(new_n485), .A2(G128), .ZN(new_n791));
  OR2_X1    g366(.A1(G104), .A2(G2105), .ZN(new_n792));
  OAI211_X1 g367(.A(new_n792), .B(G2104), .C1(G116), .C2(new_n465), .ZN(new_n793));
  NAND3_X1  g368(.A1(new_n790), .A2(new_n791), .A3(new_n793), .ZN(new_n794));
  INV_X1    g369(.A(new_n794), .ZN(new_n795));
  OAI21_X1  g370(.A(new_n789), .B1(new_n795), .B2(new_n728), .ZN(new_n796));
  INV_X1    g371(.A(G2067), .ZN(new_n797));
  XNOR2_X1  g372(.A(new_n796), .B(new_n797), .ZN(new_n798));
  NAND4_X1  g373(.A1(new_n783), .A2(new_n784), .A3(new_n787), .A4(new_n798), .ZN(new_n799));
  XNOR2_X1  g374(.A(new_n799), .B(KEYINPUT96), .ZN(new_n800));
  NAND3_X1  g375(.A1(new_n726), .A2(new_n780), .A3(new_n800), .ZN(new_n801));
  NOR2_X1   g376(.A1(G16), .A2(G22), .ZN(new_n802));
  AOI21_X1  g377(.A(new_n802), .B1(G166), .B2(G16), .ZN(new_n803));
  XNOR2_X1  g378(.A(new_n803), .B(G1971), .ZN(new_n804));
  NAND2_X1  g379(.A1(new_n721), .A2(G23), .ZN(new_n805));
  INV_X1    g380(.A(G288), .ZN(new_n806));
  OAI21_X1  g381(.A(new_n805), .B1(new_n806), .B2(new_n721), .ZN(new_n807));
  XOR2_X1   g382(.A(KEYINPUT33), .B(G1976), .Z(new_n808));
  XNOR2_X1  g383(.A(new_n807), .B(new_n808), .ZN(new_n809));
  NOR2_X1   g384(.A1(new_n804), .A2(new_n809), .ZN(new_n810));
  MUX2_X1   g385(.A(G6), .B(G305), .S(G16), .Z(new_n811));
  XOR2_X1   g386(.A(KEYINPUT32), .B(G1981), .Z(new_n812));
  AND2_X1   g387(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  NOR2_X1   g388(.A1(new_n811), .A2(new_n812), .ZN(new_n814));
  OAI21_X1  g389(.A(new_n810), .B1(new_n813), .B2(new_n814), .ZN(new_n815));
  INV_X1    g390(.A(KEYINPUT34), .ZN(new_n816));
  NAND2_X1  g391(.A1(new_n815), .A2(new_n816), .ZN(new_n817));
  OAI211_X1 g392(.A(new_n810), .B(KEYINPUT34), .C1(new_n813), .C2(new_n814), .ZN(new_n818));
  NAND2_X1  g393(.A1(new_n817), .A2(new_n818), .ZN(new_n819));
  NAND2_X1  g394(.A1(new_n485), .A2(G119), .ZN(new_n820));
  XNOR2_X1  g395(.A(new_n820), .B(KEYINPUT95), .ZN(new_n821));
  OAI21_X1  g396(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n822));
  INV_X1    g397(.A(G107), .ZN(new_n823));
  AOI21_X1  g398(.A(new_n822), .B1(new_n823), .B2(G2105), .ZN(new_n824));
  AOI21_X1  g399(.A(new_n824), .B1(new_n467), .B2(G131), .ZN(new_n825));
  NAND2_X1  g400(.A1(new_n821), .A2(new_n825), .ZN(new_n826));
  INV_X1    g401(.A(new_n826), .ZN(new_n827));
  NAND2_X1  g402(.A1(new_n827), .A2(G29), .ZN(new_n828));
  OAI21_X1  g403(.A(new_n828), .B1(G25), .B2(G29), .ZN(new_n829));
  XOR2_X1   g404(.A(KEYINPUT35), .B(G1991), .Z(new_n830));
  OR2_X1    g405(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  NOR2_X1   g406(.A1(new_n613), .A2(new_n721), .ZN(new_n832));
  AOI21_X1  g407(.A(new_n832), .B1(new_n721), .B2(G24), .ZN(new_n833));
  INV_X1    g408(.A(G1986), .ZN(new_n834));
  OR2_X1    g409(.A1(new_n833), .A2(new_n834), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n829), .A2(new_n830), .ZN(new_n836));
  NAND2_X1  g411(.A1(new_n833), .A2(new_n834), .ZN(new_n837));
  NAND4_X1  g412(.A1(new_n831), .A2(new_n835), .A3(new_n836), .A4(new_n837), .ZN(new_n838));
  INV_X1    g413(.A(new_n838), .ZN(new_n839));
  NAND2_X1  g414(.A1(new_n819), .A2(new_n839), .ZN(new_n840));
  NAND2_X1  g415(.A1(new_n840), .A2(KEYINPUT36), .ZN(new_n841));
  INV_X1    g416(.A(KEYINPUT36), .ZN(new_n842));
  NAND3_X1  g417(.A1(new_n819), .A2(new_n842), .A3(new_n839), .ZN(new_n843));
  AOI21_X1  g418(.A(new_n801), .B1(new_n841), .B2(new_n843), .ZN(G311));
  NAND2_X1  g419(.A1(new_n841), .A2(new_n843), .ZN(new_n845));
  NAND4_X1  g420(.A1(new_n845), .A2(new_n800), .A3(new_n780), .A4(new_n726), .ZN(G150));
  AOI22_X1  g421(.A1(new_n507), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n847));
  OR2_X1    g422(.A1(new_n847), .A2(new_n518), .ZN(new_n848));
  AOI22_X1  g423(.A1(new_n509), .A2(G93), .B1(G55), .B2(new_n514), .ZN(new_n849));
  NAND3_X1  g424(.A1(new_n556), .A2(new_n848), .A3(new_n849), .ZN(new_n850));
  INV_X1    g425(.A(KEYINPUT102), .ZN(new_n851));
  NAND3_X1  g426(.A1(new_n848), .A2(new_n849), .A3(new_n851), .ZN(new_n852));
  INV_X1    g427(.A(G93), .ZN(new_n853));
  INV_X1    g428(.A(G55), .ZN(new_n854));
  OAI22_X1  g429(.A1(new_n550), .A2(new_n853), .B1(new_n526), .B2(new_n854), .ZN(new_n855));
  NOR2_X1   g430(.A1(new_n847), .A2(new_n518), .ZN(new_n856));
  OAI21_X1  g431(.A(KEYINPUT102), .B1(new_n855), .B2(new_n856), .ZN(new_n857));
  NAND2_X1  g432(.A1(new_n852), .A2(new_n857), .ZN(new_n858));
  INV_X1    g433(.A(new_n858), .ZN(new_n859));
  OAI21_X1  g434(.A(new_n850), .B1(new_n859), .B2(new_n556), .ZN(new_n860));
  XNOR2_X1  g435(.A(new_n860), .B(KEYINPUT38), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n634), .A2(G559), .ZN(new_n862));
  XNOR2_X1  g437(.A(new_n861), .B(new_n862), .ZN(new_n863));
  INV_X1    g438(.A(KEYINPUT39), .ZN(new_n864));
  AOI21_X1  g439(.A(G860), .B1(new_n863), .B2(new_n864), .ZN(new_n865));
  OAI21_X1  g440(.A(new_n865), .B1(new_n864), .B2(new_n863), .ZN(new_n866));
  XOR2_X1   g441(.A(new_n866), .B(KEYINPUT103), .Z(new_n867));
  NAND2_X1  g442(.A1(new_n858), .A2(G860), .ZN(new_n868));
  XOR2_X1   g443(.A(new_n868), .B(KEYINPUT37), .Z(new_n869));
  NAND2_X1  g444(.A1(new_n867), .A2(new_n869), .ZN(G145));
  XOR2_X1   g445(.A(G160), .B(new_n657), .Z(new_n871));
  XNOR2_X1  g446(.A(new_n871), .B(G162), .ZN(new_n872));
  INV_X1    g447(.A(new_n872), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n485), .A2(G130), .ZN(new_n874));
  NOR2_X1   g449(.A1(new_n465), .A2(G118), .ZN(new_n875));
  OAI21_X1  g450(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n876));
  INV_X1    g451(.A(G142), .ZN(new_n877));
  OAI221_X1 g452(.A(new_n874), .B1(new_n875), .B2(new_n876), .C1(new_n877), .C2(new_n466), .ZN(new_n878));
  XNOR2_X1  g453(.A(new_n878), .B(KEYINPUT104), .ZN(new_n879));
  XOR2_X1   g454(.A(new_n879), .B(new_n648), .Z(new_n880));
  XNOR2_X1  g455(.A(new_n745), .B(new_n767), .ZN(new_n881));
  XNOR2_X1  g456(.A(new_n880), .B(new_n881), .ZN(new_n882));
  XNOR2_X1  g457(.A(new_n794), .B(G164), .ZN(new_n883));
  XNOR2_X1  g458(.A(new_n883), .B(new_n826), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n882), .A2(new_n884), .ZN(new_n885));
  INV_X1    g460(.A(new_n885), .ZN(new_n886));
  NOR2_X1   g461(.A1(new_n882), .A2(new_n884), .ZN(new_n887));
  OAI21_X1  g462(.A(new_n873), .B1(new_n886), .B2(new_n887), .ZN(new_n888));
  OR2_X1    g463(.A1(new_n882), .A2(new_n884), .ZN(new_n889));
  NAND3_X1  g464(.A1(new_n889), .A2(new_n872), .A3(new_n885), .ZN(new_n890));
  INV_X1    g465(.A(G37), .ZN(new_n891));
  NAND3_X1  g466(.A1(new_n888), .A2(new_n890), .A3(new_n891), .ZN(new_n892));
  XNOR2_X1  g467(.A(new_n892), .B(KEYINPUT40), .ZN(G395));
  NOR4_X1   g468(.A1(new_n555), .A2(new_n553), .A3(new_n855), .A4(new_n856), .ZN(new_n894));
  INV_X1    g469(.A(new_n556), .ZN(new_n895));
  AOI21_X1  g470(.A(new_n894), .B1(new_n895), .B2(new_n858), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n642), .A2(new_n896), .ZN(new_n897));
  NAND3_X1  g472(.A1(new_n634), .A2(new_n640), .A3(new_n860), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  INV_X1    g474(.A(KEYINPUT105), .ZN(new_n900));
  NAND3_X1  g475(.A1(new_n633), .A2(new_n900), .A3(G299), .ZN(new_n901));
  NAND3_X1  g476(.A1(new_n570), .A2(KEYINPUT105), .A3(new_n576), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n573), .A2(new_n575), .ZN(new_n903));
  OAI21_X1  g478(.A(new_n900), .B1(new_n569), .B2(new_n903), .ZN(new_n904));
  NAND4_X1  g479(.A1(new_n902), .A2(new_n632), .A3(new_n622), .A4(new_n904), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n901), .A2(new_n905), .ZN(new_n906));
  INV_X1    g481(.A(KEYINPUT106), .ZN(new_n907));
  NAND3_X1  g482(.A1(new_n906), .A2(new_n907), .A3(KEYINPUT41), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n906), .A2(KEYINPUT41), .ZN(new_n909));
  INV_X1    g484(.A(KEYINPUT41), .ZN(new_n910));
  NAND3_X1  g485(.A1(new_n901), .A2(new_n905), .A3(new_n910), .ZN(new_n911));
  NAND3_X1  g486(.A1(new_n909), .A2(KEYINPUT106), .A3(new_n911), .ZN(new_n912));
  NAND3_X1  g487(.A1(new_n899), .A2(new_n908), .A3(new_n912), .ZN(new_n913));
  INV_X1    g488(.A(new_n906), .ZN(new_n914));
  NAND3_X1  g489(.A1(new_n897), .A2(new_n914), .A3(new_n898), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n913), .A2(new_n915), .ZN(new_n916));
  XNOR2_X1  g491(.A(G166), .B(G288), .ZN(new_n917));
  NOR3_X1   g492(.A1(new_n599), .A2(new_n606), .A3(new_n613), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n598), .A2(KEYINPUT82), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n604), .A2(new_n605), .ZN(new_n920));
  AOI21_X1  g495(.A(G290), .B1(new_n919), .B2(new_n920), .ZN(new_n921));
  OAI21_X1  g496(.A(new_n917), .B1(new_n918), .B2(new_n921), .ZN(new_n922));
  XNOR2_X1  g497(.A(G166), .B(new_n806), .ZN(new_n923));
  OAI21_X1  g498(.A(new_n613), .B1(new_n599), .B2(new_n606), .ZN(new_n924));
  NAND3_X1  g499(.A1(new_n919), .A2(new_n920), .A3(G290), .ZN(new_n925));
  NAND3_X1  g500(.A1(new_n923), .A2(new_n924), .A3(new_n925), .ZN(new_n926));
  AND2_X1   g501(.A1(new_n922), .A2(new_n926), .ZN(new_n927));
  INV_X1    g502(.A(KEYINPUT42), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n922), .A2(new_n926), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n930), .A2(KEYINPUT42), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n929), .A2(new_n931), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n916), .A2(new_n932), .ZN(new_n933));
  NAND4_X1  g508(.A1(new_n913), .A2(new_n929), .A3(new_n915), .A4(new_n931), .ZN(new_n934));
  AOI21_X1  g509(.A(new_n615), .B1(new_n933), .B2(new_n934), .ZN(new_n935));
  NOR2_X1   g510(.A1(new_n859), .A2(G868), .ZN(new_n936));
  NOR2_X1   g511(.A1(new_n935), .A2(new_n936), .ZN(new_n937));
  XNOR2_X1  g512(.A(new_n937), .B(KEYINPUT107), .ZN(G295));
  INV_X1    g513(.A(new_n937), .ZN(G331));
  INV_X1    g514(.A(KEYINPUT108), .ZN(new_n940));
  AND3_X1   g515(.A1(new_n538), .A2(G301), .A3(new_n539), .ZN(new_n941));
  AOI21_X1  g516(.A(G301), .B1(new_n538), .B2(new_n539), .ZN(new_n942));
  OAI21_X1  g517(.A(new_n860), .B1(new_n941), .B2(new_n942), .ZN(new_n943));
  NAND2_X1  g518(.A1(G168), .A2(G171), .ZN(new_n944));
  NAND3_X1  g519(.A1(new_n538), .A2(G301), .A3(new_n539), .ZN(new_n945));
  NAND3_X1  g520(.A1(new_n944), .A2(new_n896), .A3(new_n945), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n943), .A2(new_n946), .ZN(new_n947));
  NAND3_X1  g522(.A1(new_n912), .A2(new_n947), .A3(new_n908), .ZN(new_n948));
  NAND3_X1  g523(.A1(new_n943), .A2(new_n946), .A3(new_n914), .ZN(new_n949));
  NAND3_X1  g524(.A1(new_n948), .A2(new_n927), .A3(new_n949), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n950), .A2(new_n891), .ZN(new_n951));
  AOI21_X1  g526(.A(new_n927), .B1(new_n948), .B2(new_n949), .ZN(new_n952));
  OAI21_X1  g527(.A(KEYINPUT43), .B1(new_n951), .B2(new_n952), .ZN(new_n953));
  AOI22_X1  g528(.A1(new_n946), .A2(new_n943), .B1(new_n909), .B2(new_n911), .ZN(new_n954));
  AND3_X1   g529(.A1(new_n943), .A2(new_n946), .A3(new_n914), .ZN(new_n955));
  OAI21_X1  g530(.A(new_n930), .B1(new_n954), .B2(new_n955), .ZN(new_n956));
  INV_X1    g531(.A(KEYINPUT43), .ZN(new_n957));
  NAND4_X1  g532(.A1(new_n950), .A2(new_n956), .A3(new_n957), .A4(new_n891), .ZN(new_n958));
  AOI21_X1  g533(.A(new_n940), .B1(new_n953), .B2(new_n958), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n948), .A2(new_n949), .ZN(new_n960));
  NAND2_X1  g535(.A1(new_n960), .A2(new_n930), .ZN(new_n961));
  NAND3_X1  g536(.A1(new_n961), .A2(new_n891), .A3(new_n950), .ZN(new_n962));
  AOI21_X1  g537(.A(KEYINPUT108), .B1(new_n962), .B2(KEYINPUT43), .ZN(new_n963));
  NOR3_X1   g538(.A1(new_n959), .A2(KEYINPUT44), .A3(new_n963), .ZN(new_n964));
  INV_X1    g539(.A(KEYINPUT44), .ZN(new_n965));
  NAND3_X1  g540(.A1(new_n950), .A2(new_n956), .A3(new_n891), .ZN(new_n966));
  AOI21_X1  g541(.A(KEYINPUT109), .B1(new_n966), .B2(KEYINPUT43), .ZN(new_n967));
  NOR3_X1   g542(.A1(new_n951), .A2(KEYINPUT43), .A3(new_n952), .ZN(new_n968));
  NOR2_X1   g543(.A1(new_n967), .A2(new_n968), .ZN(new_n969));
  NAND3_X1  g544(.A1(new_n966), .A2(KEYINPUT109), .A3(KEYINPUT43), .ZN(new_n970));
  AOI21_X1  g545(.A(new_n965), .B1(new_n969), .B2(new_n970), .ZN(new_n971));
  NOR2_X1   g546(.A1(new_n964), .A2(new_n971), .ZN(G397));
  NAND2_X1  g547(.A1(new_n469), .A2(G101), .ZN(new_n973));
  INV_X1    g548(.A(G137), .ZN(new_n974));
  OAI211_X1 g549(.A(G40), .B(new_n973), .C1(new_n466), .C2(new_n974), .ZN(new_n975));
  INV_X1    g550(.A(KEYINPUT45), .ZN(new_n976));
  OAI21_X1  g551(.A(new_n976), .B1(G164), .B2(G1384), .ZN(new_n977));
  AOI211_X1 g552(.A(new_n975), .B(new_n977), .C1(new_n473), .C2(new_n481), .ZN(new_n978));
  INV_X1    g553(.A(G1996), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n978), .A2(new_n979), .ZN(new_n980));
  XNOR2_X1  g555(.A(new_n980), .B(KEYINPUT46), .ZN(new_n981));
  XNOR2_X1  g556(.A(new_n794), .B(new_n797), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n982), .A2(new_n767), .ZN(new_n983));
  NAND2_X1  g558(.A1(new_n978), .A2(new_n983), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n981), .A2(new_n984), .ZN(new_n985));
  XNOR2_X1  g560(.A(new_n985), .B(KEYINPUT125), .ZN(new_n986));
  INV_X1    g561(.A(KEYINPUT47), .ZN(new_n987));
  OR2_X1    g562(.A1(new_n986), .A2(new_n987), .ZN(new_n988));
  NAND2_X1  g563(.A1(new_n986), .A2(new_n987), .ZN(new_n989));
  NAND3_X1  g564(.A1(new_n978), .A2(new_n834), .A3(new_n613), .ZN(new_n990));
  XOR2_X1   g565(.A(KEYINPUT126), .B(KEYINPUT48), .Z(new_n991));
  XNOR2_X1  g566(.A(new_n990), .B(new_n991), .ZN(new_n992));
  XNOR2_X1  g567(.A(new_n767), .B(G1996), .ZN(new_n993));
  OR2_X1    g568(.A1(new_n827), .A2(new_n830), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n827), .A2(new_n830), .ZN(new_n995));
  NAND4_X1  g570(.A1(new_n993), .A2(new_n994), .A3(new_n982), .A4(new_n995), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n996), .A2(new_n978), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n993), .A2(new_n982), .ZN(new_n998));
  OAI22_X1  g573(.A1(new_n998), .A2(new_n995), .B1(G2067), .B2(new_n794), .ZN(new_n999));
  AOI22_X1  g574(.A1(new_n992), .A2(new_n997), .B1(new_n978), .B2(new_n999), .ZN(new_n1000));
  AND3_X1   g575(.A1(new_n988), .A2(new_n989), .A3(new_n1000), .ZN(new_n1001));
  INV_X1    g576(.A(G1384), .ZN(new_n1002));
  INV_X1    g577(.A(new_n505), .ZN(new_n1003));
  AOI21_X1  g578(.A(new_n504), .B1(new_n464), .B2(new_n501), .ZN(new_n1004));
  NOR2_X1   g579(.A1(new_n1003), .A2(new_n1004), .ZN(new_n1005));
  OAI211_X1 g580(.A(KEYINPUT45), .B(new_n1002), .C1(new_n1005), .C2(new_n499), .ZN(new_n1006));
  AOI21_X1  g581(.A(new_n975), .B1(new_n473), .B2(new_n481), .ZN(new_n1007));
  NAND3_X1  g582(.A1(new_n977), .A2(new_n1006), .A3(new_n1007), .ZN(new_n1008));
  INV_X1    g583(.A(G1966), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n1008), .A2(new_n1009), .ZN(new_n1010));
  OAI21_X1  g585(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n1011));
  INV_X1    g586(.A(KEYINPUT50), .ZN(new_n1012));
  OAI211_X1 g587(.A(new_n1012), .B(new_n1002), .C1(new_n1005), .C2(new_n499), .ZN(new_n1013));
  NAND4_X1  g588(.A1(new_n1011), .A2(new_n1013), .A3(new_n1007), .A4(new_n756), .ZN(new_n1014));
  NAND3_X1  g589(.A1(new_n1010), .A2(G168), .A3(new_n1014), .ZN(new_n1015));
  AND2_X1   g590(.A1(KEYINPUT121), .A2(G8), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n1015), .A2(new_n1016), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n1017), .A2(KEYINPUT51), .ZN(new_n1018));
  INV_X1    g593(.A(G8), .ZN(new_n1019));
  AOI21_X1  g594(.A(new_n1019), .B1(new_n1010), .B2(new_n1014), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n1020), .A2(G286), .ZN(new_n1021));
  INV_X1    g596(.A(KEYINPUT51), .ZN(new_n1022));
  NAND3_X1  g597(.A1(new_n1015), .A2(new_n1022), .A3(new_n1016), .ZN(new_n1023));
  NAND3_X1  g598(.A1(new_n1018), .A2(new_n1021), .A3(new_n1023), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n1024), .A2(KEYINPUT62), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n1025), .A2(KEYINPUT123), .ZN(new_n1026));
  INV_X1    g601(.A(KEYINPUT123), .ZN(new_n1027));
  NAND3_X1  g602(.A1(new_n1024), .A2(new_n1027), .A3(KEYINPUT62), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n503), .A2(new_n505), .ZN(new_n1029));
  AND2_X1   g604(.A1(new_n494), .A2(new_n498), .ZN(new_n1030));
  AOI21_X1  g605(.A(G1384), .B1(new_n1029), .B2(new_n1030), .ZN(new_n1031));
  OAI21_X1  g606(.A(KEYINPUT110), .B1(new_n1031), .B2(KEYINPUT45), .ZN(new_n1032));
  INV_X1    g607(.A(KEYINPUT110), .ZN(new_n1033));
  OAI211_X1 g608(.A(new_n1033), .B(new_n976), .C1(G164), .C2(G1384), .ZN(new_n1034));
  NAND4_X1  g609(.A1(new_n1032), .A2(new_n1007), .A3(new_n1006), .A4(new_n1034), .ZN(new_n1035));
  XNOR2_X1  g610(.A(KEYINPUT111), .B(G1971), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n1035), .A2(new_n1036), .ZN(new_n1037));
  AND3_X1   g612(.A1(new_n1011), .A2(new_n1007), .A3(new_n1013), .ZN(new_n1038));
  INV_X1    g613(.A(G2090), .ZN(new_n1039));
  NAND3_X1  g614(.A1(new_n1038), .A2(KEYINPUT112), .A3(new_n1039), .ZN(new_n1040));
  NAND4_X1  g615(.A1(new_n1011), .A2(new_n1013), .A3(new_n1007), .A4(new_n1039), .ZN(new_n1041));
  INV_X1    g616(.A(KEYINPUT112), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n1041), .A2(new_n1042), .ZN(new_n1043));
  NAND3_X1  g618(.A1(new_n1037), .A2(new_n1040), .A3(new_n1043), .ZN(new_n1044));
  NAND3_X1  g619(.A1(G303), .A2(KEYINPUT55), .A3(G8), .ZN(new_n1045));
  INV_X1    g620(.A(KEYINPUT55), .ZN(new_n1046));
  OAI21_X1  g621(.A(new_n1046), .B1(G166), .B2(new_n1019), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n1045), .A2(new_n1047), .ZN(new_n1048));
  NAND3_X1  g623(.A1(new_n1044), .A2(G8), .A3(new_n1048), .ZN(new_n1049));
  AOI22_X1  g624(.A1(new_n1035), .A2(new_n1036), .B1(new_n1038), .B2(new_n1039), .ZN(new_n1050));
  OAI211_X1 g625(.A(new_n1047), .B(new_n1045), .C1(new_n1050), .C2(new_n1019), .ZN(new_n1051));
  AOI21_X1  g626(.A(new_n1019), .B1(new_n1007), .B2(new_n1031), .ZN(new_n1052));
  NAND4_X1  g627(.A1(new_n584), .A2(G1976), .A3(new_n585), .A4(new_n588), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n1052), .A2(new_n1053), .ZN(new_n1054));
  NAND2_X1  g629(.A1(new_n1054), .A2(KEYINPUT52), .ZN(new_n1055));
  INV_X1    g630(.A(G1976), .ZN(new_n1056));
  AOI21_X1  g631(.A(KEYINPUT52), .B1(G288), .B2(new_n1056), .ZN(new_n1057));
  NAND3_X1  g632(.A1(new_n1057), .A2(new_n1052), .A3(new_n1053), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n1055), .A2(new_n1058), .ZN(new_n1059));
  INV_X1    g634(.A(G1981), .ZN(new_n1060));
  OAI211_X1 g635(.A(new_n1060), .B(new_n600), .C1(new_n601), .C2(new_n603), .ZN(new_n1061));
  OAI21_X1  g636(.A(G1981), .B1(new_n592), .B2(new_n595), .ZN(new_n1062));
  AND3_X1   g637(.A1(new_n1061), .A2(KEYINPUT49), .A3(new_n1062), .ZN(new_n1063));
  AOI21_X1  g638(.A(KEYINPUT49), .B1(new_n1061), .B2(new_n1062), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n1007), .A2(new_n1031), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n1065), .A2(G8), .ZN(new_n1066));
  NOR3_X1   g641(.A1(new_n1063), .A2(new_n1064), .A3(new_n1066), .ZN(new_n1067));
  NOR2_X1   g642(.A1(new_n1059), .A2(new_n1067), .ZN(new_n1068));
  NAND3_X1  g643(.A1(new_n1049), .A2(new_n1051), .A3(new_n1068), .ZN(new_n1069));
  INV_X1    g644(.A(KEYINPUT53), .ZN(new_n1070));
  OAI21_X1  g645(.A(new_n1070), .B1(new_n1035), .B2(G2078), .ZN(new_n1071));
  NAND3_X1  g646(.A1(new_n1011), .A2(new_n1007), .A3(new_n1013), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n1072), .A2(new_n777), .ZN(new_n1073));
  AND2_X1   g648(.A1(new_n1006), .A2(new_n1007), .ZN(new_n1074));
  NOR2_X1   g649(.A1(new_n1070), .A2(G2078), .ZN(new_n1075));
  NAND3_X1  g650(.A1(new_n1074), .A2(new_n977), .A3(new_n1075), .ZN(new_n1076));
  NAND3_X1  g651(.A1(new_n1071), .A2(new_n1073), .A3(new_n1076), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n1077), .A2(G171), .ZN(new_n1078));
  NOR2_X1   g653(.A1(new_n1069), .A2(new_n1078), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n1023), .A2(new_n1021), .ZN(new_n1080));
  AOI21_X1  g655(.A(new_n1022), .B1(new_n1015), .B2(new_n1016), .ZN(new_n1081));
  OR3_X1    g656(.A1(new_n1080), .A2(KEYINPUT62), .A3(new_n1081), .ZN(new_n1082));
  NAND4_X1  g657(.A1(new_n1026), .A2(new_n1028), .A3(new_n1079), .A4(new_n1082), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n1061), .A2(new_n1062), .ZN(new_n1084));
  INV_X1    g659(.A(KEYINPUT49), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n1084), .A2(new_n1085), .ZN(new_n1086));
  NAND3_X1  g661(.A1(new_n1061), .A2(KEYINPUT49), .A3(new_n1062), .ZN(new_n1087));
  NAND3_X1  g662(.A1(new_n1086), .A2(new_n1052), .A3(new_n1087), .ZN(new_n1088));
  AND3_X1   g663(.A1(new_n1088), .A2(new_n1056), .A3(new_n806), .ZN(new_n1089));
  INV_X1    g664(.A(new_n1061), .ZN(new_n1090));
  OAI21_X1  g665(.A(new_n1052), .B1(new_n1089), .B2(new_n1090), .ZN(new_n1091));
  NAND3_X1  g666(.A1(new_n1088), .A2(new_n1055), .A3(new_n1058), .ZN(new_n1092));
  OAI21_X1  g667(.A(new_n1091), .B1(new_n1049), .B2(new_n1092), .ZN(new_n1093));
  XOR2_X1   g668(.A(KEYINPUT114), .B(KEYINPUT63), .Z(new_n1094));
  INV_X1    g669(.A(KEYINPUT113), .ZN(new_n1095));
  NAND3_X1  g670(.A1(new_n1020), .A2(new_n1095), .A3(G168), .ZN(new_n1096));
  INV_X1    g671(.A(new_n1096), .ZN(new_n1097));
  AOI21_X1  g672(.A(new_n1095), .B1(new_n1020), .B2(G168), .ZN(new_n1098));
  NOR2_X1   g673(.A1(new_n1097), .A2(new_n1098), .ZN(new_n1099));
  OAI21_X1  g674(.A(new_n1094), .B1(new_n1069), .B2(new_n1099), .ZN(new_n1100));
  AOI22_X1  g675(.A1(new_n1035), .A2(new_n1036), .B1(new_n1042), .B2(new_n1041), .ZN(new_n1101));
  AOI21_X1  g676(.A(new_n1019), .B1(new_n1101), .B2(new_n1040), .ZN(new_n1102));
  OR2_X1    g677(.A1(new_n1102), .A2(new_n1048), .ZN(new_n1103));
  AOI21_X1  g678(.A(new_n1092), .B1(new_n1102), .B2(new_n1048), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n1020), .A2(G168), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n1105), .A2(KEYINPUT113), .ZN(new_n1106));
  NAND2_X1  g681(.A1(new_n1106), .A2(new_n1096), .ZN(new_n1107));
  NAND4_X1  g682(.A1(new_n1103), .A2(new_n1104), .A3(new_n1107), .A4(KEYINPUT63), .ZN(new_n1108));
  AOI21_X1  g683(.A(new_n1093), .B1(new_n1100), .B2(new_n1108), .ZN(new_n1109));
  INV_X1    g684(.A(KEYINPUT122), .ZN(new_n1110));
  OR2_X1    g685(.A1(G171), .A2(KEYINPUT54), .ZN(new_n1111));
  NAND2_X1  g686(.A1(G171), .A2(KEYINPUT54), .ZN(new_n1112));
  OAI21_X1  g687(.A(new_n1075), .B1(new_n472), .B2(new_n465), .ZN(new_n1113));
  AOI211_X1 g688(.A(new_n975), .B(new_n1113), .C1(new_n1031), .C2(KEYINPUT45), .ZN(new_n1114));
  AOI22_X1  g689(.A1(new_n1111), .A2(new_n1112), .B1(new_n1114), .B2(new_n977), .ZN(new_n1115));
  NAND3_X1  g690(.A1(new_n1071), .A2(new_n1115), .A3(new_n1073), .ZN(new_n1116));
  AND2_X1   g691(.A1(new_n1111), .A2(new_n1112), .ZN(new_n1117));
  NAND2_X1  g692(.A1(new_n1077), .A2(new_n1117), .ZN(new_n1118));
  OAI211_X1 g693(.A(new_n1116), .B(new_n1118), .C1(new_n1080), .C2(new_n1081), .ZN(new_n1119));
  OAI21_X1  g694(.A(new_n1110), .B1(new_n1119), .B2(new_n1069), .ZN(new_n1120));
  AND3_X1   g695(.A1(new_n1049), .A2(new_n1051), .A3(new_n1068), .ZN(new_n1121));
  AND2_X1   g696(.A1(new_n1071), .A2(new_n1073), .ZN(new_n1122));
  AOI22_X1  g697(.A1(new_n1122), .A2(new_n1115), .B1(new_n1077), .B2(new_n1117), .ZN(new_n1123));
  NAND4_X1  g698(.A1(new_n1121), .A2(KEYINPUT122), .A3(new_n1024), .A4(new_n1123), .ZN(new_n1124));
  NAND2_X1  g699(.A1(new_n1120), .A2(new_n1124), .ZN(new_n1125));
  XOR2_X1   g700(.A(KEYINPUT115), .B(G1956), .Z(new_n1126));
  NAND2_X1  g701(.A1(new_n1072), .A2(new_n1126), .ZN(new_n1127));
  INV_X1    g702(.A(KEYINPUT57), .ZN(new_n1128));
  NAND3_X1  g703(.A1(new_n570), .A2(new_n1128), .A3(new_n576), .ZN(new_n1129));
  OAI21_X1  g704(.A(KEYINPUT57), .B1(new_n569), .B2(new_n903), .ZN(new_n1130));
  AND2_X1   g705(.A1(new_n1129), .A2(new_n1130), .ZN(new_n1131));
  XNOR2_X1  g706(.A(KEYINPUT56), .B(G2072), .ZN(new_n1132));
  INV_X1    g707(.A(new_n1132), .ZN(new_n1133));
  OAI211_X1 g708(.A(new_n1127), .B(new_n1131), .C1(new_n1035), .C2(new_n1133), .ZN(new_n1134));
  INV_X1    g709(.A(G1348), .ZN(new_n1135));
  NAND2_X1  g710(.A1(new_n1072), .A2(new_n1135), .ZN(new_n1136));
  INV_X1    g711(.A(KEYINPUT116), .ZN(new_n1137));
  OAI21_X1  g712(.A(new_n1137), .B1(new_n1065), .B2(G2067), .ZN(new_n1138));
  NAND4_X1  g713(.A1(new_n1007), .A2(KEYINPUT116), .A3(new_n797), .A4(new_n1031), .ZN(new_n1139));
  NAND3_X1  g714(.A1(new_n1136), .A2(new_n1138), .A3(new_n1139), .ZN(new_n1140));
  NAND3_X1  g715(.A1(new_n1134), .A2(new_n634), .A3(new_n1140), .ZN(new_n1141));
  INV_X1    g716(.A(KEYINPUT117), .ZN(new_n1142));
  AND3_X1   g717(.A1(new_n1129), .A2(new_n1142), .A3(new_n1130), .ZN(new_n1143));
  AOI21_X1  g718(.A(new_n1142), .B1(new_n1129), .B2(new_n1130), .ZN(new_n1144));
  NOR2_X1   g719(.A1(new_n1143), .A2(new_n1144), .ZN(new_n1145));
  OAI21_X1  g720(.A(new_n1127), .B1(new_n1035), .B2(new_n1133), .ZN(new_n1146));
  NAND2_X1  g721(.A1(new_n1145), .A2(new_n1146), .ZN(new_n1147));
  NAND2_X1  g722(.A1(new_n1141), .A2(new_n1147), .ZN(new_n1148));
  NAND2_X1  g723(.A1(new_n1148), .A2(KEYINPUT118), .ZN(new_n1149));
  INV_X1    g724(.A(KEYINPUT118), .ZN(new_n1150));
  NAND3_X1  g725(.A1(new_n1141), .A2(new_n1150), .A3(new_n1147), .ZN(new_n1151));
  NAND2_X1  g726(.A1(new_n1149), .A2(new_n1151), .ZN(new_n1152));
  XOR2_X1   g727(.A(KEYINPUT58), .B(G1341), .Z(new_n1153));
  NAND2_X1  g728(.A1(new_n1065), .A2(new_n1153), .ZN(new_n1154));
  OAI21_X1  g729(.A(new_n1154), .B1(new_n1035), .B2(G1996), .ZN(new_n1155));
  NAND2_X1  g730(.A1(new_n1155), .A2(new_n556), .ZN(new_n1156));
  NAND2_X1  g731(.A1(new_n1156), .A2(KEYINPUT59), .ZN(new_n1157));
  INV_X1    g732(.A(KEYINPUT59), .ZN(new_n1158));
  NAND3_X1  g733(.A1(new_n1155), .A2(new_n1158), .A3(new_n556), .ZN(new_n1159));
  NAND2_X1  g734(.A1(new_n1157), .A2(new_n1159), .ZN(new_n1160));
  INV_X1    g735(.A(KEYINPUT119), .ZN(new_n1161));
  NAND2_X1  g736(.A1(new_n1134), .A2(new_n1161), .ZN(new_n1162));
  NAND4_X1  g737(.A1(new_n1074), .A2(new_n1032), .A3(new_n1034), .A4(new_n1132), .ZN(new_n1163));
  NAND4_X1  g738(.A1(new_n1163), .A2(KEYINPUT119), .A3(new_n1131), .A4(new_n1127), .ZN(new_n1164));
  NAND4_X1  g739(.A1(new_n1162), .A2(new_n1147), .A3(KEYINPUT61), .A4(new_n1164), .ZN(new_n1165));
  INV_X1    g740(.A(KEYINPUT61), .ZN(new_n1166));
  INV_X1    g741(.A(new_n1134), .ZN(new_n1167));
  AOI21_X1  g742(.A(new_n1131), .B1(new_n1163), .B2(new_n1127), .ZN(new_n1168));
  OAI21_X1  g743(.A(new_n1166), .B1(new_n1167), .B2(new_n1168), .ZN(new_n1169));
  AND3_X1   g744(.A1(new_n1160), .A2(new_n1165), .A3(new_n1169), .ZN(new_n1170));
  AND2_X1   g745(.A1(new_n1136), .A2(new_n1139), .ZN(new_n1171));
  NAND4_X1  g746(.A1(new_n1171), .A2(KEYINPUT120), .A3(KEYINPUT60), .A4(new_n1138), .ZN(new_n1172));
  INV_X1    g747(.A(KEYINPUT120), .ZN(new_n1173));
  INV_X1    g748(.A(KEYINPUT60), .ZN(new_n1174));
  OAI21_X1  g749(.A(new_n1173), .B1(new_n1140), .B2(new_n1174), .ZN(new_n1175));
  NAND3_X1  g750(.A1(new_n1172), .A2(new_n1175), .A3(new_n634), .ZN(new_n1176));
  NAND2_X1  g751(.A1(new_n1140), .A2(new_n1174), .ZN(new_n1177));
  OAI211_X1 g752(.A(new_n1176), .B(new_n1177), .C1(new_n634), .C2(new_n1175), .ZN(new_n1178));
  AOI21_X1  g753(.A(new_n1152), .B1(new_n1170), .B2(new_n1178), .ZN(new_n1179));
  OAI211_X1 g754(.A(new_n1083), .B(new_n1109), .C1(new_n1125), .C2(new_n1179), .ZN(new_n1180));
  XNOR2_X1  g755(.A(new_n613), .B(new_n834), .ZN(new_n1181));
  OAI21_X1  g756(.A(new_n978), .B1(new_n996), .B2(new_n1181), .ZN(new_n1182));
  AND3_X1   g757(.A1(new_n1180), .A2(KEYINPUT124), .A3(new_n1182), .ZN(new_n1183));
  AOI21_X1  g758(.A(KEYINPUT124), .B1(new_n1180), .B2(new_n1182), .ZN(new_n1184));
  OAI21_X1  g759(.A(new_n1001), .B1(new_n1183), .B2(new_n1184), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g760(.A1(new_n959), .A2(new_n963), .ZN(new_n1187));
  AOI22_X1  g761(.A1(new_n714), .A2(new_n715), .B1(new_n675), .B2(new_n677), .ZN(new_n1188));
  NOR2_X1   g762(.A1(G227), .A2(new_n462), .ZN(new_n1189));
  XNOR2_X1  g763(.A(new_n1189), .B(KEYINPUT127), .ZN(new_n1190));
  NAND3_X1  g764(.A1(new_n892), .A2(new_n1188), .A3(new_n1190), .ZN(new_n1191));
  NOR2_X1   g765(.A1(new_n1187), .A2(new_n1191), .ZN(G308));
  OR2_X1    g766(.A1(new_n1187), .A2(new_n1191), .ZN(G225));
endmodule


