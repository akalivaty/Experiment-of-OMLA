

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
         n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706,
         n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717,
         n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
         n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739,
         n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750,
         n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761,
         n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772,
         n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783,
         n784, n785, n786, n787, n788, n789, n790, n791, n792, n793;

  XNOR2_X1 U375 ( .A(n485), .B(n583), .ZN(n452) );
  XNOR2_X1 U376 ( .A(n571), .B(G134), .ZN(n485) );
  XNOR2_X1 U377 ( .A(n417), .B(n606), .ZN(n768) );
  XNOR2_X2 U378 ( .A(G128), .B(KEYINPUT64), .ZN(n535) );
  XNOR2_X2 U379 ( .A(n425), .B(n424), .ZN(n785) );
  XNOR2_X2 U380 ( .A(n423), .B(KEYINPUT31), .ZN(n743) );
  NOR2_X2 U381 ( .A1(n373), .A2(n681), .ZN(n682) );
  NOR2_X2 U382 ( .A1(n503), .A2(n692), .ZN(n641) );
  XNOR2_X2 U383 ( .A(n503), .B(n490), .ZN(n681) );
  XNOR2_X2 U384 ( .A(n497), .B(n361), .ZN(n503) );
  XNOR2_X1 U385 ( .A(n506), .B(n505), .ZN(n791) );
  NOR2_X1 U386 ( .A1(n664), .A2(n653), .ZN(n733) );
  NOR2_X1 U387 ( .A1(n791), .A2(n733), .ZN(n658) );
  INV_X1 U388 ( .A(KEYINPUT84), .ZN(n420) );
  NOR2_X1 U389 ( .A1(n723), .A2(n762), .ZN(n507) );
  NOR2_X1 U390 ( .A1(n752), .A2(n762), .ZN(n753) );
  XNOR2_X1 U391 ( .A(n421), .B(n420), .ZN(n704) );
  NOR2_X1 U392 ( .A1(n775), .A2(n600), .ZN(n529) );
  NAND2_X1 U393 ( .A1(n658), .A2(n785), .ZN(n384) );
  XNOR2_X1 U394 ( .A(n464), .B(n684), .ZN(n455) );
  XNOR2_X1 U395 ( .A(n427), .B(n426), .ZN(n792) );
  NOR2_X2 U396 ( .A1(n372), .A2(n686), .ZN(n737) );
  XNOR2_X1 U397 ( .A(n676), .B(n536), .ZN(n372) );
  OR2_X1 U398 ( .A1(n695), .A2(n693), .ZN(n429) );
  NAND2_X2 U399 ( .A1(n442), .A2(n441), .ZN(n675) );
  XNOR2_X1 U400 ( .A(n615), .B(n502), .ZN(n677) );
  AND2_X1 U401 ( .A1(n720), .A2(n476), .ZN(n615) );
  XNOR2_X1 U402 ( .A(n450), .B(n577), .ZN(n657) );
  XNOR2_X1 U403 ( .A(n451), .B(n569), .ZN(n579) );
  XNOR2_X1 U404 ( .A(n773), .B(n517), .ZN(n375) );
  XNOR2_X1 U405 ( .A(n452), .B(n516), .ZN(n773) );
  XNOR2_X1 U406 ( .A(n683), .B(KEYINPUT86), .ZN(n684) );
  NAND2_X1 U407 ( .A1(n702), .A2(n745), .ZN(n775) );
  XNOR2_X2 U408 ( .A(n514), .B(n513), .ZN(n793) );
  XNOR2_X1 U409 ( .A(n698), .B(KEYINPUT105), .ZN(n439) );
  NOR2_X1 U410 ( .A1(n706), .A2(n461), .ZN(n487) );
  NOR2_X1 U411 ( .A1(n666), .A2(n665), .ZN(n667) );
  INV_X1 U412 ( .A(n687), .ZN(n661) );
  AND2_X1 U413 ( .A1(n675), .A2(n473), .ZN(n512) );
  NAND2_X1 U414 ( .A1(n472), .A2(n474), .ZN(n471) );
  XNOR2_X1 U415 ( .A(n377), .B(n508), .ZN(n376) );
  INV_X1 U416 ( .A(n591), .ZN(n516) );
  AND2_X1 U417 ( .A1(n659), .A2(n663), .ZN(n628) );
  NOR2_X1 U418 ( .A1(n430), .A2(n429), .ZN(n696) );
  OR2_X1 U419 ( .A1(n755), .A2(G902), .ZN(n450) );
  INV_X1 U420 ( .A(KEYINPUT0), .ZN(n462) );
  NAND2_X1 U421 ( .A1(n468), .A2(n786), .ZN(n374) );
  NAND2_X1 U422 ( .A1(n469), .A2(KEYINPUT81), .ZN(n468) );
  NAND2_X1 U423 ( .A1(n470), .A2(n737), .ZN(n469) );
  NOR2_X1 U424 ( .A1(n687), .A2(n690), .ZN(n470) );
  INV_X1 U425 ( .A(KEYINPUT48), .ZN(n409) );
  XOR2_X1 U426 ( .A(KEYINPUT4), .B(G146), .Z(n582) );
  AND2_X1 U427 ( .A1(n428), .A2(n668), .ZN(n382) );
  XNOR2_X1 U428 ( .A(n499), .B(G119), .ZN(n498) );
  INV_X1 U429 ( .A(KEYINPUT70), .ZN(n499) );
  XNOR2_X1 U430 ( .A(n535), .B(n534), .ZN(n571) );
  INV_X1 U431 ( .A(G143), .ZN(n534) );
  XNOR2_X1 U432 ( .A(G101), .B(KEYINPUT75), .ZN(n459) );
  NAND2_X1 U433 ( .A1(n478), .A2(G902), .ZN(n477) );
  OR2_X1 U434 ( .A1(n760), .A2(G902), .ZN(n369) );
  XNOR2_X1 U435 ( .A(n479), .B(n613), .ZN(n720) );
  XNOR2_X1 U436 ( .A(n452), .B(n606), .ZN(n479) );
  XNOR2_X1 U437 ( .A(n496), .B(n573), .ZN(n592) );
  XNOR2_X1 U438 ( .A(n572), .B(KEYINPUT83), .ZN(n496) );
  XNOR2_X1 U439 ( .A(n447), .B(n446), .ZN(n574) );
  XNOR2_X1 U440 ( .A(G107), .B(KEYINPUT99), .ZN(n446) );
  XNOR2_X1 U441 ( .A(n448), .B(KEYINPUT98), .ZN(n447) );
  INV_X1 U442 ( .A(KEYINPUT7), .ZN(n448) );
  XNOR2_X1 U443 ( .A(n575), .B(n527), .ZN(n526) );
  INV_X1 U444 ( .A(KEYINPUT9), .ZN(n527) );
  XNOR2_X1 U445 ( .A(G116), .B(G122), .ZN(n575) );
  XNOR2_X1 U446 ( .A(n387), .B(KEYINPUT80), .ZN(n386) );
  INV_X1 U447 ( .A(n775), .ZN(n531) );
  NOR2_X1 U448 ( .A1(n484), .A2(n438), .ZN(n437) );
  NOR2_X1 U449 ( .A1(n435), .A2(n467), .ZN(n434) );
  NOR2_X1 U450 ( .A1(n699), .A2(KEYINPUT43), .ZN(n435) );
  INV_X1 U451 ( .A(KEYINPUT43), .ZN(n438) );
  INV_X1 U452 ( .A(KEYINPUT39), .ZN(n515) );
  NOR2_X1 U453 ( .A1(n483), .A2(n480), .ZN(n399) );
  AND2_X1 U454 ( .A1(n696), .A2(n363), .ZN(n483) );
  NAND2_X1 U455 ( .A1(n481), .A2(n484), .ZN(n480) );
  INV_X1 U456 ( .A(n489), .ZN(n467) );
  INV_X1 U457 ( .A(KEYINPUT109), .ZN(n536) );
  XNOR2_X1 U458 ( .A(n568), .B(G475), .ZN(n569) );
  INV_X1 U459 ( .A(KEYINPUT22), .ZN(n445) );
  AND2_X1 U460 ( .A1(n649), .A2(n472), .ZN(n650) );
  INV_X2 U461 ( .A(G953), .ZN(n776) );
  XNOR2_X1 U462 ( .A(n586), .B(G104), .ZN(n587) );
  NOR2_X1 U463 ( .A1(G952), .A2(n776), .ZN(n762) );
  XNOR2_X1 U464 ( .A(n394), .B(n620), .ZN(n707) );
  NAND2_X1 U465 ( .A1(n393), .A2(n391), .ZN(n394) );
  AND2_X1 U466 ( .A1(n649), .A2(n392), .ZN(n391) );
  XNOR2_X1 U467 ( .A(n617), .B(n488), .ZN(n706) );
  INV_X1 U468 ( .A(KEYINPUT33), .ZN(n488) );
  NAND2_X1 U469 ( .A1(n521), .A2(n691), .ZN(n520) );
  NAND2_X1 U470 ( .A1(n458), .A2(n523), .ZN(n457) );
  INV_X1 U471 ( .A(n520), .ZN(n402) );
  XOR2_X1 U472 ( .A(KEYINPUT90), .B(KEYINPUT18), .Z(n550) );
  NOR2_X1 U473 ( .A1(n455), .A2(KEYINPUT48), .ZN(n454) );
  OR2_X1 U474 ( .A1(G237), .A2(G902), .ZN(n557) );
  OR2_X1 U475 ( .A1(n701), .A2(n739), .ZN(n687) );
  XNOR2_X1 U476 ( .A(KEYINPUT96), .B(G137), .ZN(n607) );
  NAND2_X1 U477 ( .A1(n379), .A2(n378), .ZN(n377) );
  INV_X1 U478 ( .A(KEYINPUT44), .ZN(n378) );
  INV_X1 U479 ( .A(n384), .ZN(n379) );
  INV_X1 U480 ( .A(KEYINPUT88), .ZN(n396) );
  XNOR2_X1 U481 ( .A(n539), .B(n538), .ZN(n772) );
  XNOR2_X1 U482 ( .A(G125), .B(G140), .ZN(n538) );
  XNOR2_X1 U483 ( .A(n540), .B(KEYINPUT66), .ZN(n539) );
  INV_X1 U484 ( .A(KEYINPUT10), .ZN(n540) );
  INV_X1 U485 ( .A(KEYINPUT2), .ZN(n533) );
  XNOR2_X1 U486 ( .A(n371), .B(KEYINPUT68), .ZN(n370) );
  NOR2_X1 U487 ( .A1(n671), .A2(n679), .ZN(n371) );
  OR2_X1 U488 ( .A1(n692), .A2(n407), .ZN(n406) );
  NAND2_X1 U489 ( .A1(n482), .A2(n407), .ZN(n481) );
  NAND2_X1 U490 ( .A1(n467), .A2(n392), .ZN(n482) );
  XNOR2_X1 U491 ( .A(n614), .B(G472), .ZN(n502) );
  NAND2_X1 U492 ( .A1(n493), .A2(n492), .ZN(n606) );
  NAND2_X1 U493 ( .A1(n495), .A2(KEYINPUT3), .ZN(n493) );
  INV_X1 U494 ( .A(KEYINPUT3), .ZN(n544) );
  XOR2_X1 U495 ( .A(G137), .B(KEYINPUT67), .Z(n591) );
  XNOR2_X1 U496 ( .A(n772), .B(n537), .ZN(n590) );
  INV_X1 U497 ( .A(G146), .ZN(n537) );
  NOR2_X1 U498 ( .A1(G237), .A2(G953), .ZN(n563) );
  XNOR2_X1 U499 ( .A(G113), .B(G131), .ZN(n560) );
  XOR2_X1 U500 ( .A(KEYINPUT12), .B(G143), .Z(n561) );
  XOR2_X1 U501 ( .A(G122), .B(G104), .Z(n559) );
  XOR2_X1 U502 ( .A(n585), .B(KEYINPUT93), .Z(n586) );
  XNOR2_X1 U503 ( .A(n584), .B(G140), .ZN(n585) );
  XNOR2_X1 U504 ( .A(n415), .B(n541), .ZN(n418) );
  XNOR2_X1 U505 ( .A(n459), .B(n416), .ZN(n415) );
  INV_X1 U506 ( .A(G110), .ZN(n416) );
  AND2_X1 U507 ( .A1(n715), .A2(G210), .ZN(n528) );
  NOR2_X1 U508 ( .A1(n656), .A2(n657), .ZN(n649) );
  XNOR2_X1 U509 ( .A(n742), .B(KEYINPUT102), .ZN(n701) );
  AND2_X1 U510 ( .A1(n443), .A2(n477), .ZN(n442) );
  NAND2_X1 U511 ( .A1(n589), .A2(n476), .ZN(n475) );
  XOR2_X1 U512 ( .A(n720), .B(KEYINPUT62), .Z(n722) );
  AND2_X1 U513 ( .A1(n715), .A2(G472), .ZN(n389) );
  XNOR2_X1 U514 ( .A(n418), .B(n419), .ZN(n417) );
  XNOR2_X1 U515 ( .A(n559), .B(KEYINPUT16), .ZN(n419) );
  XNOR2_X1 U516 ( .A(n576), .B(n524), .ZN(n755) );
  XNOR2_X1 U517 ( .A(n574), .B(n526), .ZN(n525) );
  NAND2_X1 U518 ( .A1(n715), .A2(n386), .ZN(n385) );
  AND2_X1 U519 ( .A1(n436), .A2(n434), .ZN(n433) );
  INV_X1 U520 ( .A(KEYINPUT42), .ZN(n426) );
  INV_X1 U521 ( .A(KEYINPUT40), .ZN(n513) );
  XNOR2_X1 U522 ( .A(n398), .B(n397), .ZN(n789) );
  INV_X1 U523 ( .A(KEYINPUT111), .ZN(n397) );
  NAND2_X1 U524 ( .A1(n399), .A2(n360), .ZN(n398) );
  INV_X1 U525 ( .A(KEYINPUT35), .ZN(n424) );
  INV_X1 U526 ( .A(KEYINPUT32), .ZN(n505) );
  INV_X1 U527 ( .A(n662), .ZN(n460) );
  XNOR2_X1 U528 ( .A(n465), .B(KEYINPUT107), .ZN(n786) );
  NAND2_X1 U529 ( .A1(n467), .A2(n359), .ZN(n466) );
  NAND2_X1 U530 ( .A1(n494), .A2(n358), .ZN(n668) );
  XNOR2_X1 U531 ( .A(n491), .B(KEYINPUT87), .ZN(n494) );
  XOR2_X1 U532 ( .A(n749), .B(KEYINPUT59), .Z(n751) );
  XNOR2_X1 U533 ( .A(n746), .B(n504), .ZN(n748) );
  XOR2_X1 U534 ( .A(KEYINPUT92), .B(n558), .Z(n692) );
  INV_X1 U535 ( .A(n692), .ZN(n392) );
  INV_X1 U536 ( .A(n699), .ZN(n484) );
  BUF_X1 U537 ( .A(n503), .Z(n489) );
  AND2_X1 U538 ( .A1(n372), .A2(n690), .ZN(n355) );
  XNOR2_X1 U539 ( .A(KEYINPUT25), .B(n602), .ZN(n356) );
  XNOR2_X1 U540 ( .A(n677), .B(n616), .ZN(n694) );
  INV_X1 U541 ( .A(n694), .ZN(n430) );
  XNOR2_X1 U542 ( .A(n675), .B(KEYINPUT1), .ZN(n659) );
  XNOR2_X1 U543 ( .A(n605), .B(KEYINPUT21), .ZN(n671) );
  XNOR2_X1 U544 ( .A(KEYINPUT79), .B(n703), .ZN(n357) );
  AND2_X1 U545 ( .A1(n699), .A2(n660), .ZN(n358) );
  AND2_X1 U546 ( .A1(n657), .A2(n656), .ZN(n359) );
  OR2_X1 U547 ( .A1(n696), .A2(n697), .ZN(n360) );
  INV_X1 U548 ( .A(G902), .ZN(n476) );
  NAND2_X1 U549 ( .A1(n557), .A2(G210), .ZN(n361) );
  NOR2_X1 U550 ( .A1(n680), .A2(n664), .ZN(n362) );
  NOR2_X1 U551 ( .A1(n489), .A2(n406), .ZN(n363) );
  AND2_X1 U552 ( .A1(n655), .A2(n430), .ZN(n364) );
  AND2_X1 U553 ( .A1(n699), .A2(n654), .ZN(n365) );
  INV_X1 U554 ( .A(n697), .ZN(n407) );
  INV_X1 U555 ( .A(KEYINPUT71), .ZN(n508) );
  XNOR2_X1 U556 ( .A(G902), .B(KEYINPUT15), .ZN(n600) );
  XNOR2_X1 U557 ( .A(KEYINPUT72), .B(KEYINPUT34), .ZN(n366) );
  OR2_X1 U558 ( .A1(n600), .A2(n533), .ZN(n367) );
  INV_X1 U559 ( .A(KEYINPUT74), .ZN(n522) );
  XOR2_X1 U560 ( .A(KEYINPUT56), .B(KEYINPUT122), .Z(n368) );
  NAND2_X1 U561 ( .A1(n370), .A2(n672), .ZN(n693) );
  XNOR2_X2 U562 ( .A(n369), .B(n356), .ZN(n672) );
  XNOR2_X1 U563 ( .A(n598), .B(n599), .ZN(n760) );
  OR2_X1 U564 ( .A1(n707), .A2(n372), .ZN(n427) );
  NOR2_X1 U565 ( .A1(n466), .A2(n373), .ZN(n465) );
  NAND2_X1 U566 ( .A1(n422), .A2(n510), .ZN(n373) );
  INV_X1 U567 ( .A(n374), .ZN(n519) );
  NAND2_X1 U568 ( .A1(n374), .A2(KEYINPUT74), .ZN(n404) );
  NAND2_X1 U569 ( .A1(n375), .A2(n478), .ZN(n443) );
  OR2_X1 U570 ( .A1(n375), .A2(n475), .ZN(n441) );
  XNOR2_X1 U571 ( .A(n375), .B(n747), .ZN(n504) );
  NAND2_X1 U572 ( .A1(n380), .A2(n376), .ZN(n395) );
  XNOR2_X1 U573 ( .A(n381), .B(n396), .ZN(n380) );
  NAND2_X1 U574 ( .A1(n383), .A2(n382), .ZN(n381) );
  NAND2_X1 U575 ( .A1(n384), .A2(KEYINPUT44), .ZN(n383) );
  NAND2_X1 U576 ( .A1(n385), .A2(n705), .ZN(n709) );
  NAND2_X1 U577 ( .A1(n530), .A2(n533), .ZN(n387) );
  NAND2_X1 U578 ( .A1(n388), .A2(n509), .ZN(n750) );
  AND2_X1 U579 ( .A1(n715), .A2(G475), .ZN(n388) );
  AND2_X1 U580 ( .A1(n509), .A2(n715), .ZN(n390) );
  NAND2_X1 U581 ( .A1(n389), .A2(n509), .ZN(n721) );
  NAND2_X1 U582 ( .A1(n390), .A2(G217), .ZN(n759) );
  NAND2_X1 U583 ( .A1(n390), .A2(G469), .ZN(n746) );
  NAND2_X1 U584 ( .A1(n390), .A2(G478), .ZN(n757) );
  INV_X1 U585 ( .A(n681), .ZN(n393) );
  NOR2_X1 U586 ( .A1(n681), .A2(n692), .ZN(n619) );
  XNOR2_X2 U587 ( .A(n395), .B(KEYINPUT45), .ZN(n532) );
  NAND2_X1 U588 ( .A1(n400), .A2(n789), .ZN(n456) );
  NAND2_X1 U589 ( .A1(n403), .A2(n401), .ZN(n400) );
  NAND2_X1 U590 ( .A1(n402), .A2(n522), .ZN(n401) );
  NAND2_X1 U591 ( .A1(n405), .A2(n404), .ZN(n403) );
  NAND2_X1 U592 ( .A1(n519), .A2(n518), .ZN(n405) );
  NAND2_X1 U593 ( .A1(n454), .A2(n453), .ZN(n414) );
  NAND2_X1 U594 ( .A1(n410), .A2(n408), .ZN(n412) );
  NAND2_X1 U595 ( .A1(n787), .A2(n409), .ZN(n408) );
  NAND2_X1 U596 ( .A1(n411), .A2(n787), .ZN(n410) );
  NOR2_X1 U597 ( .A1(n456), .A2(n455), .ZN(n411) );
  NAND2_X1 U598 ( .A1(n412), .A2(n414), .ZN(n413) );
  XNOR2_X2 U599 ( .A(n413), .B(KEYINPUT85), .ZN(n702) );
  INV_X1 U600 ( .A(n418), .ZN(n588) );
  NAND2_X1 U601 ( .A1(n702), .A2(n357), .ZN(n421) );
  XNOR2_X1 U602 ( .A(n678), .B(KEYINPUT30), .ZN(n422) );
  NAND2_X2 U603 ( .A1(n463), .A2(n367), .ZN(n509) );
  NAND2_X1 U604 ( .A1(n460), .A2(n651), .ZN(n423) );
  NAND2_X1 U605 ( .A1(n486), .A2(n359), .ZN(n425) );
  XNOR2_X1 U606 ( .A(n667), .B(KEYINPUT103), .ZN(n428) );
  NAND2_X1 U607 ( .A1(n439), .A2(n437), .ZN(n436) );
  NAND2_X1 U608 ( .A1(n433), .A2(n431), .ZN(n700) );
  NAND2_X1 U609 ( .A1(n432), .A2(n438), .ZN(n431) );
  INV_X1 U610 ( .A(n439), .ZN(n432) );
  NAND2_X1 U611 ( .A1(n440), .A2(n739), .ZN(n514) );
  XNOR2_X1 U612 ( .A(n682), .B(n515), .ZN(n440) );
  NAND2_X1 U613 ( .A1(n440), .A2(n701), .ZN(n745) );
  NAND2_X1 U614 ( .A1(n444), .A2(n364), .ZN(n506) );
  NAND2_X1 U615 ( .A1(n444), .A2(n365), .ZN(n653) );
  NAND2_X1 U616 ( .A1(n444), .A2(n430), .ZN(n491) );
  XNOR2_X2 U617 ( .A(n652), .B(n445), .ZN(n444) );
  XNOR2_X2 U618 ( .A(n449), .B(KEYINPUT101), .ZN(n742) );
  NAND2_X1 U619 ( .A1(n579), .A2(n657), .ZN(n449) );
  NOR2_X1 U620 ( .A1(n749), .A2(G902), .ZN(n451) );
  INV_X1 U621 ( .A(n456), .ZN(n453) );
  NOR2_X1 U622 ( .A1(n457), .A2(n355), .ZN(n521) );
  NAND2_X1 U623 ( .A1(n686), .A2(n690), .ZN(n458) );
  INV_X1 U624 ( .A(n651), .ZN(n461) );
  AND2_X1 U625 ( .A1(n651), .A2(n362), .ZN(n728) );
  XNOR2_X2 U626 ( .A(n648), .B(n462), .ZN(n651) );
  NAND2_X1 U627 ( .A1(n529), .A2(n532), .ZN(n463) );
  NOR2_X2 U628 ( .A1(n792), .A2(n793), .ZN(n464) );
  NOR2_X1 U629 ( .A1(n672), .A2(n471), .ZN(n473) );
  INV_X1 U630 ( .A(n671), .ZN(n472) );
  NOR2_X1 U631 ( .A1(n672), .A2(n671), .ZN(n663) );
  NAND2_X1 U632 ( .A1(n675), .A2(n663), .ZN(n680) );
  INV_X1 U633 ( .A(n679), .ZN(n474) );
  INV_X1 U634 ( .A(n589), .ZN(n478) );
  NAND2_X1 U635 ( .A1(n696), .A2(n392), .ZN(n698) );
  XNOR2_X1 U636 ( .A(n485), .B(n525), .ZN(n524) );
  XNOR2_X1 U637 ( .A(n487), .B(n366), .ZN(n486) );
  INV_X1 U638 ( .A(KEYINPUT38), .ZN(n490) );
  NAND2_X1 U639 ( .A1(n543), .A2(n544), .ZN(n492) );
  XNOR2_X1 U640 ( .A(n641), .B(n640), .ZN(n685) );
  NAND2_X1 U641 ( .A1(n685), .A2(n647), .ZN(n648) );
  INV_X1 U642 ( .A(n668), .ZN(n726) );
  XNOR2_X1 U643 ( .A(n750), .B(n751), .ZN(n752) );
  XNOR2_X1 U644 ( .A(n721), .B(n722), .ZN(n723) );
  XNOR2_X1 U645 ( .A(n597), .B(n596), .ZN(n598) );
  INV_X1 U646 ( .A(n543), .ZN(n495) );
  XNOR2_X1 U647 ( .A(n498), .B(n542), .ZN(n543) );
  NAND2_X1 U648 ( .A1(n712), .A2(n600), .ZN(n497) );
  NOR2_X1 U649 ( .A1(n709), .A2(n708), .ZN(n711) );
  NAND2_X1 U650 ( .A1(n603), .A2(G221), .ZN(n604) );
  XNOR2_X1 U651 ( .A(n601), .B(KEYINPUT20), .ZN(n603) );
  XNOR2_X2 U652 ( .A(n556), .B(n555), .ZN(n712) );
  XNOR2_X1 U653 ( .A(n500), .B(n368), .ZN(G51) );
  NAND2_X1 U654 ( .A1(n718), .A2(n719), .ZN(n500) );
  NAND2_X1 U655 ( .A1(n501), .A2(n675), .ZN(n676) );
  XNOR2_X1 U656 ( .A(n674), .B(n673), .ZN(n501) );
  XNOR2_X1 U657 ( .A(n507), .B(n725), .ZN(G57) );
  NAND2_X1 U658 ( .A1(n528), .A2(n509), .ZN(n716) );
  XNOR2_X1 U659 ( .A(n512), .B(n511), .ZN(n510) );
  INV_X1 U660 ( .A(KEYINPUT77), .ZN(n511) );
  XNOR2_X1 U661 ( .A(n588), .B(n587), .ZN(n517) );
  NAND2_X1 U662 ( .A1(n520), .A2(KEYINPUT74), .ZN(n518) );
  INV_X1 U663 ( .A(KEYINPUT81), .ZN(n523) );
  NAND2_X2 U664 ( .A1(n704), .A2(n532), .ZN(n715) );
  NAND2_X1 U665 ( .A1(n532), .A2(n531), .ZN(n530) );
  INV_X1 U666 ( .A(n571), .ZN(n570) );
  XNOR2_X1 U667 ( .A(n755), .B(n754), .ZN(n756) );
  XNOR2_X1 U668 ( .A(n554), .B(n553), .ZN(n555) );
  INV_X1 U669 ( .A(KEYINPUT19), .ZN(n640) );
  XNOR2_X1 U670 ( .A(n612), .B(n611), .ZN(n613) );
  XNOR2_X1 U671 ( .A(n565), .B(n564), .ZN(n566) );
  INV_X1 U672 ( .A(KEYINPUT13), .ZN(n568) );
  XNOR2_X1 U673 ( .A(n567), .B(n566), .ZN(n749) );
  INV_X1 U674 ( .A(KEYINPUT63), .ZN(n724) );
  XNOR2_X1 U675 ( .A(n724), .B(KEYINPUT112), .ZN(n725) );
  XNOR2_X1 U676 ( .A(n757), .B(n756), .ZN(n758) );
  XNOR2_X1 U677 ( .A(n711), .B(n710), .ZN(G75) );
  XNOR2_X1 U678 ( .A(KEYINPUT91), .B(G107), .ZN(n541) );
  XNOR2_X1 U679 ( .A(G116), .B(G113), .ZN(n542) );
  INV_X1 U680 ( .A(n768), .ZN(n546) );
  INV_X1 U681 ( .A(n582), .ZN(n545) );
  NAND2_X1 U682 ( .A1(n546), .A2(n545), .ZN(n548) );
  NAND2_X1 U683 ( .A1(n768), .A2(n582), .ZN(n547) );
  NAND2_X1 U684 ( .A1(n548), .A2(n547), .ZN(n556) );
  NAND2_X1 U685 ( .A1(G224), .A2(n776), .ZN(n549) );
  XNOR2_X1 U686 ( .A(n550), .B(n549), .ZN(n551) );
  XNOR2_X1 U687 ( .A(KEYINPUT78), .B(n551), .ZN(n552) );
  XNOR2_X1 U688 ( .A(n552), .B(n570), .ZN(n554) );
  XOR2_X1 U689 ( .A(G125), .B(KEYINPUT17), .Z(n553) );
  NAND2_X1 U690 ( .A1(G214), .A2(n557), .ZN(n558) );
  NAND2_X1 U691 ( .A1(n681), .A2(n692), .ZN(n578) );
  XNOR2_X1 U692 ( .A(n559), .B(n590), .ZN(n567) );
  XNOR2_X1 U693 ( .A(n561), .B(n560), .ZN(n562) );
  XOR2_X1 U694 ( .A(n562), .B(KEYINPUT11), .Z(n565) );
  XNOR2_X1 U695 ( .A(n563), .B(KEYINPUT76), .ZN(n610) );
  NAND2_X1 U696 ( .A1(n610), .A2(G214), .ZN(n564) );
  INV_X1 U697 ( .A(n579), .ZN(n656) );
  XOR2_X1 U698 ( .A(KEYINPUT8), .B(KEYINPUT65), .Z(n573) );
  NAND2_X1 U699 ( .A1(G234), .A2(n776), .ZN(n572) );
  NAND2_X1 U700 ( .A1(n592), .A2(G217), .ZN(n576) );
  XNOR2_X1 U701 ( .A(KEYINPUT100), .B(G478), .ZN(n577) );
  NAND2_X1 U702 ( .A1(n578), .A2(n649), .ZN(n581) );
  NOR2_X1 U703 ( .A1(n579), .A2(n657), .ZN(n739) );
  NAND2_X1 U704 ( .A1(n687), .A2(n619), .ZN(n580) );
  AND2_X1 U705 ( .A1(n581), .A2(n580), .ZN(n618) );
  XNOR2_X1 U706 ( .A(G131), .B(n582), .ZN(n583) );
  NAND2_X1 U707 ( .A1(n776), .A2(G227), .ZN(n584) );
  XNOR2_X1 U708 ( .A(KEYINPUT69), .B(G469), .ZN(n589) );
  XNOR2_X1 U709 ( .A(n591), .B(n590), .ZN(n599) );
  NAND2_X1 U710 ( .A1(n592), .A2(G221), .ZN(n597) );
  XOR2_X1 U711 ( .A(KEYINPUT24), .B(G110), .Z(n594) );
  XNOR2_X1 U712 ( .A(G119), .B(G128), .ZN(n593) );
  XNOR2_X1 U713 ( .A(n594), .B(n593), .ZN(n595) );
  XOR2_X1 U714 ( .A(n595), .B(KEYINPUT23), .Z(n596) );
  NAND2_X1 U715 ( .A1(G234), .A2(n600), .ZN(n601) );
  NAND2_X1 U716 ( .A1(G217), .A2(n603), .ZN(n602) );
  XNOR2_X1 U717 ( .A(n604), .B(KEYINPUT94), .ZN(n605) );
  XNOR2_X1 U718 ( .A(KEYINPUT6), .B(KEYINPUT104), .ZN(n616) );
  XOR2_X1 U719 ( .A(KEYINPUT95), .B(G101), .Z(n608) );
  XNOR2_X1 U720 ( .A(n608), .B(n607), .ZN(n609) );
  XOR2_X1 U721 ( .A(n609), .B(KEYINPUT5), .Z(n612) );
  NAND2_X1 U722 ( .A1(n610), .A2(G210), .ZN(n611) );
  XNOR2_X1 U723 ( .A(KEYINPUT97), .B(KEYINPUT73), .ZN(n614) );
  NAND2_X1 U724 ( .A1(n628), .A2(n694), .ZN(n617) );
  NOR2_X1 U725 ( .A1(n618), .A2(n706), .ZN(n633) );
  XOR2_X1 U726 ( .A(KEYINPUT110), .B(KEYINPUT41), .Z(n620) );
  XOR2_X1 U727 ( .A(KEYINPUT49), .B(KEYINPUT117), .Z(n622) );
  NAND2_X1 U728 ( .A1(n654), .A2(n671), .ZN(n621) );
  XNOR2_X1 U729 ( .A(n622), .B(n621), .ZN(n625) );
  NOR2_X1 U730 ( .A1(n663), .A2(n659), .ZN(n623) );
  XNOR2_X1 U731 ( .A(n623), .B(KEYINPUT50), .ZN(n624) );
  NOR2_X1 U732 ( .A1(n625), .A2(n624), .ZN(n626) );
  NAND2_X1 U733 ( .A1(n626), .A2(n677), .ZN(n627) );
  XNOR2_X1 U734 ( .A(n627), .B(KEYINPUT118), .ZN(n629) );
  INV_X1 U735 ( .A(n677), .ZN(n664) );
  NAND2_X1 U736 ( .A1(n664), .A2(n628), .ZN(n662) );
  NAND2_X1 U737 ( .A1(n629), .A2(n662), .ZN(n630) );
  XNOR2_X1 U738 ( .A(KEYINPUT51), .B(n630), .ZN(n631) );
  NOR2_X1 U739 ( .A1(n707), .A2(n631), .ZN(n632) );
  NOR2_X1 U740 ( .A1(n633), .A2(n632), .ZN(n634) );
  XOR2_X1 U741 ( .A(n634), .B(KEYINPUT119), .Z(n635) );
  XNOR2_X1 U742 ( .A(KEYINPUT52), .B(n635), .ZN(n638) );
  NAND2_X1 U743 ( .A1(G234), .A2(G237), .ZN(n636) );
  XNOR2_X1 U744 ( .A(n636), .B(KEYINPUT14), .ZN(n643) );
  NAND2_X1 U745 ( .A1(G952), .A2(n643), .ZN(n637) );
  NOR2_X1 U746 ( .A1(n638), .A2(n637), .ZN(n639) );
  NOR2_X1 U747 ( .A1(G953), .A2(n639), .ZN(n705) );
  INV_X1 U748 ( .A(n672), .ZN(n660) );
  INV_X1 U749 ( .A(n660), .ZN(n654) );
  NAND2_X1 U750 ( .A1(G953), .A2(n476), .ZN(n642) );
  NAND2_X1 U751 ( .A1(n643), .A2(n642), .ZN(n645) );
  NOR2_X1 U752 ( .A1(G953), .A2(G952), .ZN(n644) );
  NOR2_X1 U753 ( .A1(n645), .A2(n644), .ZN(n670) );
  NAND2_X1 U754 ( .A1(G898), .A2(G953), .ZN(n646) );
  AND2_X1 U755 ( .A1(n670), .A2(n646), .ZN(n647) );
  NAND2_X1 U756 ( .A1(n651), .A2(n650), .ZN(n652) );
  AND2_X1 U757 ( .A1(n659), .A2(n654), .ZN(n655) );
  INV_X1 U758 ( .A(n659), .ZN(n699) );
  XNOR2_X1 U759 ( .A(n661), .B(KEYINPUT82), .ZN(n666) );
  NOR2_X1 U760 ( .A1(n743), .A2(n728), .ZN(n665) );
  NAND2_X1 U761 ( .A1(G953), .A2(G900), .ZN(n669) );
  NAND2_X1 U762 ( .A1(n670), .A2(n669), .ZN(n679) );
  NOR2_X1 U763 ( .A1(n677), .A2(n693), .ZN(n674) );
  XNOR2_X1 U764 ( .A(KEYINPUT28), .B(KEYINPUT108), .ZN(n673) );
  NOR2_X1 U765 ( .A1(n692), .A2(n677), .ZN(n678) );
  INV_X1 U766 ( .A(KEYINPUT46), .ZN(n683) );
  INV_X1 U767 ( .A(n685), .ZN(n686) );
  INV_X1 U768 ( .A(KEYINPUT47), .ZN(n690) );
  NAND2_X1 U769 ( .A1(n690), .A2(KEYINPUT82), .ZN(n688) );
  XNOR2_X1 U770 ( .A(n688), .B(n687), .ZN(n689) );
  NAND2_X1 U771 ( .A1(n689), .A2(n737), .ZN(n691) );
  INV_X1 U772 ( .A(n739), .ZN(n695) );
  XNOR2_X1 U773 ( .A(KEYINPUT36), .B(KEYINPUT89), .ZN(n697) );
  XNOR2_X1 U774 ( .A(KEYINPUT106), .B(n700), .ZN(n787) );
  NAND2_X1 U775 ( .A1(KEYINPUT2), .A2(n745), .ZN(n703) );
  NOR2_X1 U776 ( .A1(n707), .A2(n706), .ZN(n708) );
  XNOR2_X1 U777 ( .A(KEYINPUT120), .B(KEYINPUT53), .ZN(n710) );
  INV_X1 U778 ( .A(n762), .ZN(n719) );
  XNOR2_X1 U779 ( .A(KEYINPUT54), .B(KEYINPUT121), .ZN(n714) );
  XNOR2_X1 U780 ( .A(n712), .B(KEYINPUT55), .ZN(n713) );
  XNOR2_X1 U781 ( .A(n714), .B(n713), .ZN(n717) );
  XNOR2_X1 U782 ( .A(n717), .B(n716), .ZN(n718) );
  XOR2_X1 U783 ( .A(G101), .B(n726), .Z(G3) );
  NAND2_X1 U784 ( .A1(n728), .A2(n739), .ZN(n727) );
  XNOR2_X1 U785 ( .A(n727), .B(G104), .ZN(G6) );
  XOR2_X1 U786 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n730) );
  NAND2_X1 U787 ( .A1(n728), .A2(n742), .ZN(n729) );
  XNOR2_X1 U788 ( .A(n730), .B(n729), .ZN(n732) );
  XOR2_X1 U789 ( .A(G107), .B(KEYINPUT113), .Z(n731) );
  XNOR2_X1 U790 ( .A(n732), .B(n731), .ZN(G9) );
  XOR2_X1 U791 ( .A(G110), .B(n733), .Z(G12) );
  XOR2_X1 U792 ( .A(KEYINPUT114), .B(KEYINPUT29), .Z(n735) );
  NAND2_X1 U793 ( .A1(n737), .A2(n742), .ZN(n734) );
  XNOR2_X1 U794 ( .A(n735), .B(n734), .ZN(n736) );
  XNOR2_X1 U795 ( .A(G128), .B(n736), .ZN(G30) );
  NAND2_X1 U796 ( .A1(n737), .A2(n739), .ZN(n738) );
  XNOR2_X1 U797 ( .A(n738), .B(G146), .ZN(G48) );
  XOR2_X1 U798 ( .A(G113), .B(KEYINPUT115), .Z(n741) );
  NAND2_X1 U799 ( .A1(n743), .A2(n739), .ZN(n740) );
  XNOR2_X1 U800 ( .A(n741), .B(n740), .ZN(G15) );
  NAND2_X1 U801 ( .A1(n743), .A2(n742), .ZN(n744) );
  XNOR2_X1 U802 ( .A(n744), .B(G116), .ZN(G18) );
  XNOR2_X1 U803 ( .A(G134), .B(n745), .ZN(G36) );
  XOR2_X1 U804 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n747) );
  NOR2_X1 U805 ( .A1(n762), .A2(n748), .ZN(G54) );
  XNOR2_X1 U806 ( .A(n753), .B(KEYINPUT60), .ZN(G60) );
  INV_X1 U807 ( .A(KEYINPUT123), .ZN(n754) );
  NOR2_X1 U808 ( .A1(n762), .A2(n758), .ZN(G63) );
  XNOR2_X1 U809 ( .A(n760), .B(n759), .ZN(n761) );
  NOR2_X1 U810 ( .A1(n762), .A2(n761), .ZN(G66) );
  NAND2_X1 U811 ( .A1(n532), .A2(n776), .ZN(n766) );
  NAND2_X1 U812 ( .A1(G953), .A2(G224), .ZN(n763) );
  XNOR2_X1 U813 ( .A(KEYINPUT61), .B(n763), .ZN(n764) );
  NAND2_X1 U814 ( .A1(n764), .A2(G898), .ZN(n765) );
  NAND2_X1 U815 ( .A1(n766), .A2(n765), .ZN(n770) );
  NOR2_X1 U816 ( .A1(G898), .A2(n776), .ZN(n767) );
  NOR2_X1 U817 ( .A1(n768), .A2(n767), .ZN(n769) );
  XNOR2_X1 U818 ( .A(n770), .B(n769), .ZN(n771) );
  XNOR2_X1 U819 ( .A(KEYINPUT124), .B(n771), .ZN(G69) );
  XNOR2_X1 U820 ( .A(n773), .B(n772), .ZN(n774) );
  XNOR2_X1 U821 ( .A(n774), .B(KEYINPUT125), .ZN(n778) );
  XNOR2_X1 U822 ( .A(n775), .B(n778), .ZN(n777) );
  NAND2_X1 U823 ( .A1(n777), .A2(n776), .ZN(n784) );
  XNOR2_X1 U824 ( .A(n778), .B(KEYINPUT126), .ZN(n779) );
  XNOR2_X1 U825 ( .A(G227), .B(n779), .ZN(n780) );
  NAND2_X1 U826 ( .A1(G900), .A2(n780), .ZN(n781) );
  NAND2_X1 U827 ( .A1(G953), .A2(n781), .ZN(n782) );
  XOR2_X1 U828 ( .A(KEYINPUT127), .B(n782), .Z(n783) );
  NAND2_X1 U829 ( .A1(n784), .A2(n783), .ZN(G72) );
  XNOR2_X1 U830 ( .A(n785), .B(G122), .ZN(G24) );
  XNOR2_X1 U831 ( .A(G143), .B(n786), .ZN(G45) );
  XNOR2_X1 U832 ( .A(G140), .B(n787), .ZN(G42) );
  XOR2_X1 U833 ( .A(KEYINPUT37), .B(KEYINPUT116), .Z(n788) );
  XNOR2_X1 U834 ( .A(n789), .B(n788), .ZN(n790) );
  XNOR2_X1 U835 ( .A(G125), .B(n790), .ZN(G27) );
  XOR2_X1 U836 ( .A(n791), .B(G119), .Z(G21) );
  XOR2_X1 U837 ( .A(n792), .B(G137), .Z(G39) );
  XOR2_X1 U838 ( .A(n793), .B(G131), .Z(G33) );
endmodule

