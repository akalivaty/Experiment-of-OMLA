

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598,
         n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609,
         n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620,
         n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631,
         n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642,
         n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653,
         n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664,
         n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675,
         n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686,
         n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697,
         n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708,
         n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719,
         n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730,
         n731, n732;

  NAND2_X1 U379 ( .A1(n382), .A2(n383), .ZN(n381) );
  XNOR2_X1 U380 ( .A(n572), .B(n420), .ZN(n419) );
  NOR2_X1 U381 ( .A1(n500), .A2(n523), .ZN(n615) );
  XNOR2_X1 U382 ( .A(n714), .B(G146), .ZN(n452) );
  XNOR2_X1 U383 ( .A(n379), .B(KEYINPUT22), .ZN(n556) );
  XNOR2_X1 U384 ( .A(n397), .B(G953), .ZN(n722) );
  XNOR2_X2 U385 ( .A(n393), .B(KEYINPUT19), .ZN(n550) );
  XNOR2_X2 U386 ( .A(KEYINPUT65), .B(G128), .ZN(n410) );
  XNOR2_X2 U387 ( .A(n386), .B(n448), .ZN(n714) );
  XNOR2_X2 U388 ( .A(n460), .B(n459), .ZN(n506) );
  NOR2_X1 U389 ( .A1(n702), .A2(n681), .ZN(n682) );
  AND2_X1 U390 ( .A1(n635), .A2(n571), .ZN(n572) );
  INV_X1 U391 ( .A(n555), .ZN(n634) );
  NOR2_X1 U392 ( .A1(n702), .A2(n596), .ZN(n599) );
  NOR2_X1 U393 ( .A1(n702), .A2(n693), .ZN(n694) );
  NAND2_X1 U394 ( .A1(n591), .A2(n367), .ZN(n382) );
  NAND2_X1 U395 ( .A1(n705), .A2(n367), .ZN(n383) );
  NOR2_X1 U396 ( .A1(n566), .A2(n729), .ZN(n567) );
  XNOR2_X1 U397 ( .A(n414), .B(KEYINPUT35), .ZN(n729) );
  XNOR2_X1 U398 ( .A(n412), .B(n411), .ZN(n652) );
  XNOR2_X1 U399 ( .A(n398), .B(G146), .ZN(n465) );
  XNOR2_X2 U400 ( .A(n535), .B(n534), .ZN(n387) );
  XNOR2_X1 U401 ( .A(n468), .B(n469), .ZN(n399) );
  AND2_X1 U402 ( .A1(n585), .A2(n401), .ZN(n515) );
  NOR2_X1 U403 ( .A1(n440), .A2(n659), .ZN(n401) );
  XNOR2_X1 U404 ( .A(n384), .B(n358), .ZN(n499) );
  NAND2_X1 U405 ( .A1(n676), .A2(n543), .ZN(n384) );
  XNOR2_X1 U406 ( .A(n458), .B(KEYINPUT73), .ZN(n459) );
  XNOR2_X1 U407 ( .A(n494), .B(n403), .ZN(n715) );
  INV_X1 U408 ( .A(n454), .ZN(n403) );
  XNOR2_X1 U409 ( .A(G137), .B(G113), .ZN(n445) );
  XNOR2_X1 U410 ( .A(n444), .B(n409), .ZN(n408) );
  XOR2_X1 U411 ( .A(KEYINPUT78), .B(KEYINPUT95), .Z(n444) );
  AND2_X1 U412 ( .A1(n488), .A2(G210), .ZN(n409) );
  XOR2_X1 U413 ( .A(KEYINPUT11), .B(G122), .Z(n485) );
  NOR2_X1 U414 ( .A1(G953), .A2(G237), .ZN(n488) );
  XNOR2_X1 U415 ( .A(n493), .B(G134), .ZN(n448) );
  NAND2_X1 U416 ( .A1(n499), .A2(n643), .ZN(n393) );
  XOR2_X1 U417 ( .A(KEYINPUT76), .B(KEYINPUT16), .Z(n462) );
  XNOR2_X1 U418 ( .A(G101), .B(G116), .ZN(n441) );
  XNOR2_X1 U419 ( .A(G119), .B(KEYINPUT93), .ZN(n426) );
  XOR2_X1 U420 ( .A(KEYINPUT23), .B(KEYINPUT92), .Z(n427) );
  XOR2_X1 U421 ( .A(G113), .B(G104), .Z(n492) );
  XNOR2_X1 U422 ( .A(n465), .B(n423), .ZN(n494) );
  XOR2_X1 U423 ( .A(G104), .B(G107), .Z(n451) );
  XNOR2_X1 U424 ( .A(n385), .B(n703), .ZN(n676) );
  XNOR2_X1 U425 ( .A(n394), .B(n386), .ZN(n385) );
  XNOR2_X1 U426 ( .A(n399), .B(n467), .ZN(n394) );
  INV_X1 U427 ( .A(n624), .ZN(n541) );
  XNOR2_X1 U428 ( .A(KEYINPUT71), .B(KEYINPUT48), .ZN(n534) );
  AND2_X1 U429 ( .A1(n589), .A2(n588), .ZN(n590) );
  INV_X1 U430 ( .A(n506), .ZN(n517) );
  INV_X1 U431 ( .A(n514), .ZN(n539) );
  XNOR2_X1 U432 ( .A(n406), .B(KEYINPUT109), .ZN(n405) );
  AND2_X1 U433 ( .A1(n515), .A2(n615), .ZN(n370) );
  INV_X1 U434 ( .A(KEYINPUT1), .ZN(n413) );
  XNOR2_X1 U435 ( .A(n435), .B(n434), .ZN(n585) );
  XNOR2_X1 U436 ( .A(n433), .B(n360), .ZN(n434) );
  NOR2_X1 U437 ( .A1(n700), .A2(G902), .ZN(n435) );
  BUF_X1 U438 ( .A(n722), .Z(n369) );
  INV_X1 U439 ( .A(KEYINPUT4), .ZN(n447) );
  INV_X1 U440 ( .A(G125), .ZN(n398) );
  XNOR2_X1 U441 ( .A(KEYINPUT38), .B(n539), .ZN(n644) );
  XNOR2_X1 U442 ( .A(n452), .B(n357), .ZN(n593) );
  XNOR2_X1 U443 ( .A(n408), .B(n407), .ZN(n446) );
  XNOR2_X1 U444 ( .A(n445), .B(KEYINPUT5), .ZN(n407) );
  INV_X1 U445 ( .A(KEYINPUT64), .ZN(n397) );
  XOR2_X1 U446 ( .A(KEYINPUT105), .B(KEYINPUT7), .Z(n474) );
  XOR2_X1 U447 ( .A(KEYINPUT70), .B(G131), .Z(n493) );
  XNOR2_X1 U448 ( .A(n495), .B(n491), .ZN(n378) );
  XNOR2_X1 U449 ( .A(n489), .B(n490), .ZN(n377) );
  NAND2_X1 U450 ( .A1(G234), .A2(G237), .ZN(n422) );
  INV_X1 U451 ( .A(KEYINPUT33), .ZN(n411) );
  NAND2_X1 U452 ( .A1(n562), .A2(n570), .ZN(n412) );
  AND2_X1 U453 ( .A1(n570), .A2(n569), .ZN(n635) );
  AND2_X1 U454 ( .A1(n507), .A2(n391), .ZN(n528) );
  AND2_X1 U455 ( .A1(n573), .A2(n366), .ZN(n391) );
  NOR2_X1 U456 ( .A1(n526), .A2(n471), .ZN(n472) );
  NAND2_X1 U457 ( .A1(n380), .A2(n363), .ZN(n379) );
  INV_X1 U458 ( .A(n576), .ZN(n380) );
  XNOR2_X1 U459 ( .A(n483), .B(n371), .ZN(n500) );
  INV_X1 U460 ( .A(G478), .ZN(n371) );
  XNOR2_X1 U461 ( .A(n498), .B(n361), .ZN(n523) );
  BUF_X1 U462 ( .A(n555), .Z(n574) );
  XNOR2_X1 U463 ( .A(n464), .B(n418), .ZN(n417) );
  XNOR2_X1 U464 ( .A(n475), .B(n462), .ZN(n418) );
  XNOR2_X1 U465 ( .A(n431), .B(n402), .ZN(n700) );
  XNOR2_X1 U466 ( .A(n404), .B(n715), .ZN(n402) );
  XNOR2_X1 U467 ( .A(n376), .B(n374), .ZN(n690) );
  XNOR2_X1 U468 ( .A(n494), .B(n375), .ZN(n374) );
  XNOR2_X1 U469 ( .A(n378), .B(n377), .ZN(n376) );
  XNOR2_X1 U470 ( .A(n492), .B(n493), .ZN(n375) );
  BUF_X1 U471 ( .A(n688), .Z(n698) );
  XNOR2_X1 U472 ( .A(n452), .B(n416), .ZN(n684) );
  XNOR2_X1 U473 ( .A(n457), .B(n453), .ZN(n416) );
  NOR2_X1 U474 ( .A1(n369), .A2(G952), .ZN(n702) );
  INV_X1 U475 ( .A(G953), .ZN(n664) );
  XNOR2_X1 U476 ( .A(n388), .B(KEYINPUT86), .ZN(n592) );
  NAND2_X1 U477 ( .A1(n372), .A2(n539), .ZN(n624) );
  XNOR2_X1 U478 ( .A(n538), .B(n373), .ZN(n372) );
  XNOR2_X1 U479 ( .A(KEYINPUT43), .B(KEYINPUT111), .ZN(n373) );
  XOR2_X1 U480 ( .A(n464), .B(n446), .Z(n357) );
  AND2_X1 U481 ( .A1(G210), .A2(n470), .ZN(n358) );
  XOR2_X1 U482 ( .A(n437), .B(KEYINPUT21), .Z(n359) );
  XOR2_X1 U483 ( .A(KEYINPUT25), .B(KEYINPUT94), .Z(n360) );
  XOR2_X1 U484 ( .A(n497), .B(n496), .Z(n361) );
  AND2_X1 U485 ( .A1(n542), .A2(KEYINPUT2), .ZN(n362) );
  AND2_X1 U486 ( .A1(n551), .A2(n359), .ZN(n363) );
  XOR2_X1 U487 ( .A(G472), .B(KEYINPUT96), .Z(n364) );
  XOR2_X1 U488 ( .A(KEYINPUT67), .B(KEYINPUT0), .Z(n365) );
  AND2_X1 U489 ( .A1(n503), .A2(n502), .ZN(n366) );
  OR2_X1 U490 ( .A1(n668), .A2(n421), .ZN(n367) );
  NAND2_X1 U491 ( .A1(n368), .A2(n533), .ZN(n535) );
  XNOR2_X1 U492 ( .A(n532), .B(KEYINPUT46), .ZN(n368) );
  AND2_X2 U493 ( .A1(n387), .A2(n542), .ZN(n720) );
  NAND2_X1 U494 ( .A1(n561), .A2(n370), .ZN(n406) );
  NOR2_X2 U495 ( .A1(n556), .A2(n561), .ZN(n582) );
  NOR2_X4 U496 ( .A1(n672), .A2(n381), .ZN(n688) );
  NOR2_X2 U497 ( .A1(n705), .A2(n592), .ZN(n672) );
  XNOR2_X2 U498 ( .A(n590), .B(KEYINPUT45), .ZN(n705) );
  XNOR2_X2 U499 ( .A(n477), .B(n447), .ZN(n386) );
  NAND2_X1 U500 ( .A1(n387), .A2(n362), .ZN(n388) );
  XNOR2_X2 U501 ( .A(n389), .B(n364), .ZN(n555) );
  OR2_X2 U502 ( .A1(n593), .A2(G902), .ZN(n389) );
  XNOR2_X1 U503 ( .A(n390), .B(n529), .ZN(n540) );
  NAND2_X1 U504 ( .A1(n528), .A2(n644), .ZN(n390) );
  XNOR2_X2 U505 ( .A(n392), .B(n365), .ZN(n576) );
  NAND2_X1 U506 ( .A1(n550), .A2(n549), .ZN(n392) );
  XNOR2_X2 U507 ( .A(n410), .B(G143), .ZN(n477) );
  NAND2_X1 U508 ( .A1(n395), .A2(n612), .ZN(n509) );
  NAND2_X1 U509 ( .A1(n396), .A2(KEYINPUT47), .ZN(n395) );
  NAND2_X1 U510 ( .A1(n512), .A2(n647), .ZN(n396) );
  XNOR2_X1 U511 ( .A(n472), .B(KEYINPUT80), .ZN(n512) );
  XNOR2_X1 U512 ( .A(n400), .B(n449), .ZN(n461) );
  NAND2_X1 U513 ( .A1(n634), .A2(n515), .ZN(n400) );
  NAND2_X1 U514 ( .A1(n480), .A2(G221), .ZN(n404) );
  NAND2_X1 U515 ( .A1(n405), .A2(n643), .ZN(n536) );
  XNOR2_X2 U516 ( .A(n506), .B(n413), .ZN(n570) );
  NAND2_X1 U517 ( .A1(n415), .A2(n565), .ZN(n414) );
  XNOR2_X1 U518 ( .A(n564), .B(n563), .ZN(n415) );
  XNOR2_X1 U519 ( .A(n417), .B(n463), .ZN(n703) );
  NOR2_X1 U520 ( .A1(n419), .A2(n604), .ZN(n577) );
  NAND2_X1 U521 ( .A1(n419), .A2(n615), .ZN(n616) );
  NAND2_X1 U522 ( .A1(n419), .A2(n618), .ZN(n619) );
  INV_X1 U523 ( .A(KEYINPUT31), .ZN(n420) );
  INV_X1 U524 ( .A(n600), .ZN(n586) );
  INV_X1 U525 ( .A(KEYINPUT88), .ZN(n559) );
  INV_X1 U526 ( .A(KEYINPUT106), .ZN(n580) );
  NAND2_X1 U527 ( .A1(n720), .A2(n544), .ZN(n591) );
  INV_X1 U528 ( .A(KEYINPUT10), .ZN(n423) );
  AND2_X1 U529 ( .A1(n587), .A2(n586), .ZN(n588) );
  NOR2_X1 U530 ( .A1(n541), .A2(n622), .ZN(n542) );
  XNOR2_X1 U531 ( .A(n690), .B(n689), .ZN(n691) );
  XNOR2_X1 U532 ( .A(n684), .B(n683), .ZN(n685) );
  INV_X1 U533 ( .A(KEYINPUT32), .ZN(n553) );
  BUF_X1 U534 ( .A(n499), .Z(n514) );
  XNOR2_X1 U535 ( .A(n597), .B(KEYINPUT90), .ZN(n598) );
  XNOR2_X1 U536 ( .A(n686), .B(n685), .ZN(n687) );
  INV_X1 U537 ( .A(KEYINPUT2), .ZN(n668) );
  XNOR2_X1 U538 ( .A(G902), .B(KEYINPUT15), .ZN(n543) );
  XOR2_X1 U539 ( .A(KEYINPUT85), .B(n543), .Z(n421) );
  XOR2_X1 U540 ( .A(KEYINPUT14), .B(n422), .Z(n659) );
  INV_X1 U541 ( .A(n659), .ZN(n503) );
  XOR2_X1 U542 ( .A(G137), .B(G140), .Z(n454) );
  NAND2_X1 U543 ( .A1(n722), .A2(G234), .ZN(n425) );
  XNOR2_X1 U544 ( .A(KEYINPUT69), .B(KEYINPUT8), .ZN(n424) );
  XNOR2_X1 U545 ( .A(n425), .B(n424), .ZN(n480) );
  XNOR2_X1 U546 ( .A(n427), .B(n426), .ZN(n428) );
  XOR2_X1 U547 ( .A(n428), .B(KEYINPUT24), .Z(n430) );
  XNOR2_X1 U548 ( .A(G128), .B(G110), .ZN(n429) );
  XOR2_X1 U549 ( .A(n430), .B(n429), .Z(n431) );
  NAND2_X1 U550 ( .A1(G234), .A2(n543), .ZN(n432) );
  XNOR2_X1 U551 ( .A(KEYINPUT20), .B(n432), .ZN(n436) );
  NAND2_X1 U552 ( .A1(G217), .A2(n436), .ZN(n433) );
  NAND2_X1 U553 ( .A1(n436), .A2(G221), .ZN(n437) );
  NAND2_X1 U554 ( .A1(G952), .A2(n664), .ZN(n546) );
  NOR2_X1 U555 ( .A1(G900), .A2(n369), .ZN(n438) );
  NAND2_X1 U556 ( .A1(G902), .A2(n438), .ZN(n439) );
  NAND2_X1 U557 ( .A1(n546), .A2(n439), .ZN(n502) );
  NAND2_X1 U558 ( .A1(n359), .A2(n502), .ZN(n440) );
  INV_X1 U559 ( .A(n441), .ZN(n443) );
  XNOR2_X1 U560 ( .A(KEYINPUT3), .B(G119), .ZN(n442) );
  XNOR2_X1 U561 ( .A(n443), .B(n442), .ZN(n464) );
  XNOR2_X1 U562 ( .A(KEYINPUT28), .B(KEYINPUT113), .ZN(n449) );
  XNOR2_X1 U563 ( .A(G101), .B(G110), .ZN(n450) );
  XNOR2_X1 U564 ( .A(n451), .B(n450), .ZN(n453) );
  XOR2_X1 U565 ( .A(n454), .B(KEYINPUT91), .Z(n456) );
  NAND2_X1 U566 ( .A1(G227), .A2(n369), .ZN(n455) );
  XNOR2_X1 U567 ( .A(n456), .B(n455), .ZN(n457) );
  NOR2_X1 U568 ( .A1(G902), .A2(n684), .ZN(n460) );
  INV_X1 U569 ( .A(G469), .ZN(n458) );
  NAND2_X1 U570 ( .A1(n461), .A2(n517), .ZN(n526) );
  XNOR2_X1 U571 ( .A(G110), .B(n492), .ZN(n463) );
  XOR2_X2 U572 ( .A(G122), .B(G107), .Z(n475) );
  XOR2_X1 U573 ( .A(KEYINPUT79), .B(KEYINPUT89), .Z(n466) );
  XNOR2_X1 U574 ( .A(n466), .B(n465), .ZN(n467) );
  XOR2_X1 U575 ( .A(KEYINPUT17), .B(KEYINPUT18), .Z(n469) );
  NAND2_X1 U576 ( .A1(G224), .A2(n722), .ZN(n468) );
  OR2_X1 U577 ( .A1(G237), .A2(G902), .ZN(n470) );
  NAND2_X1 U578 ( .A1(G214), .A2(n470), .ZN(n643) );
  INV_X1 U579 ( .A(n550), .ZN(n471) );
  XNOR2_X1 U580 ( .A(G116), .B(KEYINPUT9), .ZN(n473) );
  XNOR2_X1 U581 ( .A(n474), .B(n473), .ZN(n476) );
  XOR2_X1 U582 ( .A(n476), .B(n475), .Z(n479) );
  XNOR2_X1 U583 ( .A(n477), .B(G134), .ZN(n478) );
  XNOR2_X1 U584 ( .A(n479), .B(n478), .ZN(n482) );
  NAND2_X1 U585 ( .A1(n480), .A2(G217), .ZN(n481) );
  XOR2_X1 U586 ( .A(n482), .B(n481), .Z(n696) );
  NOR2_X1 U587 ( .A1(G902), .A2(n696), .ZN(n483) );
  XNOR2_X1 U588 ( .A(G143), .B(G140), .ZN(n484) );
  XNOR2_X1 U589 ( .A(n485), .B(n484), .ZN(n495) );
  XOR2_X1 U590 ( .A(KEYINPUT100), .B(KEYINPUT102), .Z(n487) );
  XNOR2_X1 U591 ( .A(KEYINPUT101), .B(KEYINPUT98), .ZN(n486) );
  XNOR2_X1 U592 ( .A(n487), .B(n486), .ZN(n491) );
  XOR2_X1 U593 ( .A(KEYINPUT99), .B(KEYINPUT12), .Z(n490) );
  NAND2_X1 U594 ( .A1(G214), .A2(n488), .ZN(n489) );
  NOR2_X1 U595 ( .A1(n690), .A2(G902), .ZN(n498) );
  XOR2_X1 U596 ( .A(KEYINPUT13), .B(KEYINPUT104), .Z(n497) );
  XNOR2_X1 U597 ( .A(KEYINPUT103), .B(G475), .ZN(n496) );
  INV_X1 U598 ( .A(n615), .ZN(n530) );
  NAND2_X1 U599 ( .A1(n500), .A2(n523), .ZN(n603) );
  NAND2_X1 U600 ( .A1(n530), .A2(n603), .ZN(n647) );
  INV_X1 U601 ( .A(n500), .ZN(n524) );
  NOR2_X1 U602 ( .A1(n523), .A2(n524), .ZN(n501) );
  XNOR2_X1 U603 ( .A(KEYINPUT108), .B(n501), .ZN(n565) );
  NAND2_X1 U604 ( .A1(n634), .A2(n643), .ZN(n505) );
  XOR2_X1 U605 ( .A(KEYINPUT30), .B(KEYINPUT112), .Z(n504) );
  XNOR2_X1 U606 ( .A(n505), .B(n504), .ZN(n507) );
  INV_X1 U607 ( .A(n585), .ZN(n628) );
  NAND2_X1 U608 ( .A1(n628), .A2(n359), .ZN(n625) );
  NOR2_X1 U609 ( .A1(n506), .A2(n625), .ZN(n573) );
  AND2_X1 U610 ( .A1(n565), .A2(n528), .ZN(n508) );
  NAND2_X1 U611 ( .A1(n514), .A2(n508), .ZN(n612) );
  XNOR2_X1 U612 ( .A(n509), .B(KEYINPUT82), .ZN(n521) );
  XOR2_X1 U613 ( .A(KEYINPUT47), .B(KEYINPUT68), .Z(n510) );
  XOR2_X1 U614 ( .A(KEYINPUT83), .B(n647), .Z(n568) );
  NAND2_X1 U615 ( .A1(n510), .A2(n568), .ZN(n511) );
  XNOR2_X1 U616 ( .A(n511), .B(KEYINPUT77), .ZN(n513) );
  BUF_X1 U617 ( .A(n512), .Z(n613) );
  NAND2_X1 U618 ( .A1(n513), .A2(n613), .ZN(n519) );
  XNOR2_X1 U619 ( .A(n555), .B(KEYINPUT6), .ZN(n561) );
  NOR2_X1 U620 ( .A1(n539), .A2(n536), .ZN(n516) );
  XNOR2_X1 U621 ( .A(n516), .B(KEYINPUT36), .ZN(n518) );
  INV_X1 U622 ( .A(n570), .ZN(n626) );
  NAND2_X1 U623 ( .A1(n518), .A2(n570), .ZN(n621) );
  NAND2_X1 U624 ( .A1(n519), .A2(n621), .ZN(n520) );
  NOR2_X1 U625 ( .A1(n521), .A2(n520), .ZN(n522) );
  XNOR2_X1 U626 ( .A(n522), .B(KEYINPUT72), .ZN(n533) );
  NAND2_X1 U627 ( .A1(n524), .A2(n523), .ZN(n646) );
  NAND2_X1 U628 ( .A1(n644), .A2(n643), .ZN(n648) );
  NOR2_X1 U629 ( .A1(n646), .A2(n648), .ZN(n525) );
  XNOR2_X1 U630 ( .A(KEYINPUT41), .B(n525), .ZN(n640) );
  NOR2_X1 U631 ( .A1(n526), .A2(n640), .ZN(n527) );
  XNOR2_X1 U632 ( .A(n527), .B(KEYINPUT42), .ZN(n732) );
  XOR2_X1 U633 ( .A(KEYINPUT74), .B(KEYINPUT39), .Z(n529) );
  NOR2_X1 U634 ( .A1(n540), .A2(n530), .ZN(n531) );
  XNOR2_X1 U635 ( .A(n531), .B(KEYINPUT40), .ZN(n731) );
  NOR2_X1 U636 ( .A1(n732), .A2(n731), .ZN(n532) );
  XNOR2_X1 U637 ( .A(KEYINPUT110), .B(n536), .ZN(n537) );
  NOR2_X1 U638 ( .A1(n570), .A2(n537), .ZN(n538) );
  NOR2_X1 U639 ( .A1(n540), .A2(n603), .ZN(n622) );
  INV_X1 U640 ( .A(n543), .ZN(n544) );
  NAND2_X1 U641 ( .A1(n585), .A2(n570), .ZN(n545) );
  XNOR2_X1 U642 ( .A(n545), .B(KEYINPUT107), .ZN(n552) );
  NOR2_X1 U643 ( .A1(G898), .A2(n664), .ZN(n704) );
  NAND2_X1 U644 ( .A1(n704), .A2(G902), .ZN(n547) );
  AND2_X1 U645 ( .A1(n547), .A2(n546), .ZN(n548) );
  NOR2_X1 U646 ( .A1(n548), .A2(n659), .ZN(n549) );
  INV_X1 U647 ( .A(n646), .ZN(n551) );
  NAND2_X1 U648 ( .A1(n552), .A2(n582), .ZN(n554) );
  XNOR2_X1 U649 ( .A(n554), .B(n553), .ZN(n730) );
  NOR2_X1 U650 ( .A1(n556), .A2(n570), .ZN(n557) );
  NAND2_X1 U651 ( .A1(n574), .A2(n557), .ZN(n558) );
  NOR2_X1 U652 ( .A1(n628), .A2(n558), .ZN(n609) );
  NOR2_X1 U653 ( .A1(n730), .A2(n609), .ZN(n560) );
  XNOR2_X1 U654 ( .A(n560), .B(n559), .ZN(n566) );
  INV_X1 U655 ( .A(n625), .ZN(n569) );
  AND2_X1 U656 ( .A1(n561), .A2(n569), .ZN(n562) );
  NOR2_X1 U657 ( .A1(n576), .A2(n652), .ZN(n564) );
  XOR2_X1 U658 ( .A(KEYINPUT75), .B(KEYINPUT34), .Z(n563) );
  XNOR2_X1 U659 ( .A(n567), .B(KEYINPUT44), .ZN(n589) );
  INV_X1 U660 ( .A(n568), .ZN(n579) );
  NOR2_X1 U661 ( .A1(n576), .A2(n574), .ZN(n571) );
  NAND2_X1 U662 ( .A1(n574), .A2(n573), .ZN(n575) );
  NOR2_X1 U663 ( .A1(n576), .A2(n575), .ZN(n604) );
  XOR2_X1 U664 ( .A(KEYINPUT97), .B(n577), .Z(n578) );
  NOR2_X1 U665 ( .A1(n579), .A2(n578), .ZN(n581) );
  XNOR2_X1 U666 ( .A(n581), .B(n580), .ZN(n587) );
  NAND2_X1 U667 ( .A1(n582), .A2(n626), .ZN(n583) );
  XOR2_X1 U668 ( .A(KEYINPUT87), .B(n583), .Z(n584) );
  NOR2_X1 U669 ( .A1(n585), .A2(n584), .ZN(n600) );
  NAND2_X1 U670 ( .A1(n688), .A2(G472), .ZN(n595) );
  XNOR2_X1 U671 ( .A(n593), .B(KEYINPUT62), .ZN(n594) );
  XNOR2_X1 U672 ( .A(n595), .B(n594), .ZN(n596) );
  INV_X1 U673 ( .A(KEYINPUT63), .ZN(n597) );
  XNOR2_X1 U674 ( .A(n599), .B(n598), .ZN(G57) );
  XOR2_X1 U675 ( .A(G101), .B(n600), .Z(G3) );
  NAND2_X1 U676 ( .A1(n604), .A2(n615), .ZN(n601) );
  XNOR2_X1 U677 ( .A(n601), .B(KEYINPUT114), .ZN(n602) );
  XNOR2_X1 U678 ( .A(G104), .B(n602), .ZN(G6) );
  XOR2_X1 U679 ( .A(KEYINPUT26), .B(KEYINPUT115), .Z(n606) );
  INV_X1 U680 ( .A(n603), .ZN(n618) );
  NAND2_X1 U681 ( .A1(n604), .A2(n618), .ZN(n605) );
  XNOR2_X1 U682 ( .A(n606), .B(n605), .ZN(n608) );
  XOR2_X1 U683 ( .A(G107), .B(KEYINPUT27), .Z(n607) );
  XNOR2_X1 U684 ( .A(n608), .B(n607), .ZN(G9) );
  XOR2_X1 U685 ( .A(G110), .B(n609), .Z(G12) );
  XOR2_X1 U686 ( .A(G128), .B(KEYINPUT29), .Z(n611) );
  NAND2_X1 U687 ( .A1(n618), .A2(n613), .ZN(n610) );
  XNOR2_X1 U688 ( .A(n611), .B(n610), .ZN(G30) );
  XNOR2_X1 U689 ( .A(G143), .B(n612), .ZN(G45) );
  NAND2_X1 U690 ( .A1(n613), .A2(n615), .ZN(n614) );
  XNOR2_X1 U691 ( .A(n614), .B(G146), .ZN(G48) );
  XNOR2_X1 U692 ( .A(G113), .B(KEYINPUT116), .ZN(n617) );
  XNOR2_X1 U693 ( .A(n617), .B(n616), .ZN(G15) );
  XNOR2_X1 U694 ( .A(n619), .B(G116), .ZN(G18) );
  XOR2_X1 U695 ( .A(G125), .B(KEYINPUT37), .Z(n620) );
  XNOR2_X1 U696 ( .A(n621), .B(n620), .ZN(G27) );
  XNOR2_X1 U697 ( .A(G134), .B(n622), .ZN(n623) );
  XNOR2_X1 U698 ( .A(n623), .B(KEYINPUT117), .ZN(G36) );
  XNOR2_X1 U699 ( .A(G140), .B(n624), .ZN(G42) );
  NOR2_X1 U700 ( .A1(n652), .A2(n640), .ZN(n662) );
  NAND2_X1 U701 ( .A1(n626), .A2(n625), .ZN(n627) );
  XNOR2_X1 U702 ( .A(KEYINPUT50), .B(n627), .ZN(n632) );
  NOR2_X1 U703 ( .A1(n359), .A2(n628), .ZN(n629) );
  XOR2_X1 U704 ( .A(KEYINPUT49), .B(n629), .Z(n630) );
  NOR2_X1 U705 ( .A1(n634), .A2(n630), .ZN(n631) );
  NAND2_X1 U706 ( .A1(n632), .A2(n631), .ZN(n633) );
  XNOR2_X1 U707 ( .A(n633), .B(KEYINPUT118), .ZN(n637) );
  NAND2_X1 U708 ( .A1(n635), .A2(n634), .ZN(n636) );
  NAND2_X1 U709 ( .A1(n637), .A2(n636), .ZN(n639) );
  XOR2_X1 U710 ( .A(KEYINPUT119), .B(KEYINPUT51), .Z(n638) );
  XNOR2_X1 U711 ( .A(n639), .B(n638), .ZN(n641) );
  NOR2_X1 U712 ( .A1(n641), .A2(n640), .ZN(n642) );
  XOR2_X1 U713 ( .A(KEYINPUT120), .B(n642), .Z(n656) );
  NOR2_X1 U714 ( .A1(n644), .A2(n643), .ZN(n645) );
  NOR2_X1 U715 ( .A1(n646), .A2(n645), .ZN(n651) );
  INV_X1 U716 ( .A(n647), .ZN(n649) );
  NOR2_X1 U717 ( .A1(n649), .A2(n648), .ZN(n650) );
  NOR2_X1 U718 ( .A1(n651), .A2(n650), .ZN(n653) );
  NOR2_X1 U719 ( .A1(n653), .A2(n652), .ZN(n654) );
  XNOR2_X1 U720 ( .A(KEYINPUT121), .B(n654), .ZN(n655) );
  NAND2_X1 U721 ( .A1(n656), .A2(n655), .ZN(n657) );
  XNOR2_X1 U722 ( .A(KEYINPUT52), .B(n657), .ZN(n658) );
  NAND2_X1 U723 ( .A1(n658), .A2(G952), .ZN(n660) );
  NOR2_X1 U724 ( .A1(n660), .A2(n659), .ZN(n661) );
  NOR2_X1 U725 ( .A1(n662), .A2(n661), .ZN(n663) );
  XNOR2_X1 U726 ( .A(n663), .B(KEYINPUT122), .ZN(n665) );
  NAND2_X1 U727 ( .A1(n665), .A2(n664), .ZN(n674) );
  INV_X1 U728 ( .A(n720), .ZN(n666) );
  NAND2_X1 U729 ( .A1(n666), .A2(n668), .ZN(n667) );
  XNOR2_X1 U730 ( .A(n667), .B(KEYINPUT84), .ZN(n670) );
  NAND2_X1 U731 ( .A1(n705), .A2(n668), .ZN(n669) );
  NAND2_X1 U732 ( .A1(n670), .A2(n669), .ZN(n671) );
  NOR2_X1 U733 ( .A1(n672), .A2(n671), .ZN(n673) );
  NOR2_X1 U734 ( .A1(n674), .A2(n673), .ZN(n675) );
  XNOR2_X1 U735 ( .A(KEYINPUT53), .B(n675), .ZN(G75) );
  XOR2_X1 U736 ( .A(KEYINPUT54), .B(KEYINPUT55), .Z(n678) );
  XNOR2_X1 U737 ( .A(n676), .B(KEYINPUT81), .ZN(n677) );
  XNOR2_X1 U738 ( .A(n678), .B(n677), .ZN(n680) );
  NAND2_X1 U739 ( .A1(n688), .A2(G210), .ZN(n679) );
  XNOR2_X1 U740 ( .A(n680), .B(n679), .ZN(n681) );
  XNOR2_X1 U741 ( .A(KEYINPUT56), .B(n682), .ZN(G51) );
  NAND2_X1 U742 ( .A1(n698), .A2(G469), .ZN(n686) );
  XOR2_X1 U743 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n683) );
  NOR2_X1 U744 ( .A1(n702), .A2(n687), .ZN(G54) );
  NAND2_X1 U745 ( .A1(n688), .A2(G475), .ZN(n692) );
  XOR2_X1 U746 ( .A(KEYINPUT59), .B(KEYINPUT66), .Z(n689) );
  XNOR2_X1 U747 ( .A(n692), .B(n691), .ZN(n693) );
  XNOR2_X1 U748 ( .A(KEYINPUT60), .B(n694), .ZN(G60) );
  NAND2_X1 U749 ( .A1(G478), .A2(n698), .ZN(n695) );
  XNOR2_X1 U750 ( .A(n696), .B(n695), .ZN(n697) );
  NOR2_X1 U751 ( .A1(n702), .A2(n697), .ZN(G63) );
  NAND2_X1 U752 ( .A1(G217), .A2(n698), .ZN(n699) );
  XNOR2_X1 U753 ( .A(n700), .B(n699), .ZN(n701) );
  NOR2_X1 U754 ( .A1(n702), .A2(n701), .ZN(G66) );
  NOR2_X1 U755 ( .A1(n704), .A2(n703), .ZN(n713) );
  NOR2_X1 U756 ( .A1(G953), .A2(n705), .ZN(n706) );
  XNOR2_X1 U757 ( .A(KEYINPUT123), .B(n706), .ZN(n710) );
  NAND2_X1 U758 ( .A1(G953), .A2(G224), .ZN(n707) );
  XNOR2_X1 U759 ( .A(KEYINPUT61), .B(n707), .ZN(n708) );
  NAND2_X1 U760 ( .A1(n708), .A2(G898), .ZN(n709) );
  NAND2_X1 U761 ( .A1(n710), .A2(n709), .ZN(n711) );
  XNOR2_X1 U762 ( .A(n711), .B(KEYINPUT124), .ZN(n712) );
  XNOR2_X1 U763 ( .A(n713), .B(n712), .ZN(G69) );
  BUF_X1 U764 ( .A(n714), .Z(n716) );
  XOR2_X1 U765 ( .A(n716), .B(n715), .Z(n717) );
  XNOR2_X1 U766 ( .A(KEYINPUT125), .B(n717), .ZN(n723) );
  INV_X1 U767 ( .A(n723), .ZN(n718) );
  XNOR2_X1 U768 ( .A(n718), .B(KEYINPUT126), .ZN(n719) );
  XNOR2_X1 U769 ( .A(n720), .B(n719), .ZN(n721) );
  NAND2_X1 U770 ( .A1(n369), .A2(n721), .ZN(n727) );
  XNOR2_X1 U771 ( .A(G227), .B(n723), .ZN(n724) );
  NAND2_X1 U772 ( .A1(n724), .A2(G900), .ZN(n725) );
  NAND2_X1 U773 ( .A1(G953), .A2(n725), .ZN(n726) );
  NAND2_X1 U774 ( .A1(n727), .A2(n726), .ZN(n728) );
  XOR2_X1 U775 ( .A(KEYINPUT127), .B(n728), .Z(G72) );
  XOR2_X1 U776 ( .A(G122), .B(n729), .Z(G24) );
  XOR2_X1 U777 ( .A(n730), .B(G119), .Z(G21) );
  XOR2_X1 U778 ( .A(G131), .B(n731), .Z(G33) );
  XOR2_X1 U779 ( .A(G137), .B(n732), .Z(G39) );
endmodule

