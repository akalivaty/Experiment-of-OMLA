//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 0 0 1 0 0 1 1 0 0 1 1 0 0 1 1 1 1 0 0 0 1 0 0 1 0 0 0 0 0 0 0 0 0 0 1 0 1 1 1 1 0 1 1 1 0 1 0 1 1 1 0 1 1 0 0 0 1 0 1 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:18:41 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n697, new_n698, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n732, new_n733, new_n734, new_n735, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n756, new_n757, new_n758, new_n759, new_n761, new_n762, new_n763,
    new_n764, new_n766, new_n767, new_n768, new_n770, new_n772, new_n773,
    new_n774, new_n775, new_n776, new_n777, new_n778, new_n779, new_n780,
    new_n781, new_n782, new_n783, new_n784, new_n785, new_n786, new_n787,
    new_n788, new_n789, new_n790, new_n791, new_n792, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n817,
    new_n818, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n855,
    new_n856, new_n858, new_n860, new_n861, new_n862, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n906, new_n907, new_n908, new_n910,
    new_n911, new_n912, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n921, new_n922, new_n924, new_n925, new_n926, new_n927,
    new_n928, new_n929, new_n931, new_n932, new_n933, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n947, new_n948, new_n949, new_n950, new_n951, new_n952,
    new_n953, new_n954, new_n955, new_n956, new_n957, new_n958, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965;
  XNOR2_X1  g000(.A(G1gat), .B(G29gat), .ZN(new_n202));
  XNOR2_X1  g001(.A(new_n202), .B(KEYINPUT0), .ZN(new_n203));
  XNOR2_X1  g002(.A(G57gat), .B(G85gat), .ZN(new_n204));
  XOR2_X1   g003(.A(new_n203), .B(new_n204), .Z(new_n205));
  INV_X1    g004(.A(KEYINPUT66), .ZN(new_n206));
  INV_X1    g005(.A(G134gat), .ZN(new_n207));
  INV_X1    g006(.A(G127gat), .ZN(new_n208));
  NAND2_X1  g007(.A1(new_n208), .A2(KEYINPUT65), .ZN(new_n209));
  INV_X1    g008(.A(KEYINPUT65), .ZN(new_n210));
  NAND2_X1  g009(.A1(new_n210), .A2(G127gat), .ZN(new_n211));
  AOI21_X1  g010(.A(new_n207), .B1(new_n209), .B2(new_n211), .ZN(new_n212));
  NOR2_X1   g011(.A1(G127gat), .A2(G134gat), .ZN(new_n213));
  OAI21_X1  g012(.A(new_n206), .B1(new_n212), .B2(new_n213), .ZN(new_n214));
  INV_X1    g013(.A(G120gat), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n215), .A2(G113gat), .ZN(new_n216));
  INV_X1    g015(.A(G113gat), .ZN(new_n217));
  NAND2_X1  g016(.A1(new_n217), .A2(G120gat), .ZN(new_n218));
  AOI21_X1  g017(.A(KEYINPUT1), .B1(new_n216), .B2(new_n218), .ZN(new_n219));
  INV_X1    g018(.A(new_n219), .ZN(new_n220));
  INV_X1    g019(.A(new_n213), .ZN(new_n221));
  XNOR2_X1  g020(.A(KEYINPUT65), .B(G127gat), .ZN(new_n222));
  OAI211_X1 g021(.A(KEYINPUT66), .B(new_n221), .C1(new_n222), .C2(new_n207), .ZN(new_n223));
  NAND3_X1  g022(.A1(new_n214), .A2(new_n220), .A3(new_n223), .ZN(new_n224));
  XNOR2_X1  g023(.A(G127gat), .B(G134gat), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n219), .A2(new_n225), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n224), .A2(new_n226), .ZN(new_n227));
  NAND2_X1  g026(.A1(G155gat), .A2(G162gat), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n228), .A2(KEYINPUT2), .ZN(new_n229));
  OR2_X1    g028(.A1(G141gat), .A2(G148gat), .ZN(new_n230));
  NAND2_X1  g029(.A1(G141gat), .A2(G148gat), .ZN(new_n231));
  NAND3_X1  g030(.A1(new_n229), .A2(new_n230), .A3(new_n231), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n232), .A2(KEYINPUT75), .ZN(new_n233));
  XNOR2_X1  g032(.A(G155gat), .B(G162gat), .ZN(new_n234));
  INV_X1    g033(.A(new_n234), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n233), .A2(new_n235), .ZN(new_n236));
  NAND3_X1  g035(.A1(new_n232), .A2(KEYINPUT75), .A3(new_n234), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n236), .A2(new_n237), .ZN(new_n238));
  INV_X1    g037(.A(new_n238), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n227), .A2(new_n239), .ZN(new_n240));
  NAND3_X1  g039(.A1(new_n238), .A2(new_n224), .A3(new_n226), .ZN(new_n241));
  NAND3_X1  g040(.A1(new_n240), .A2(KEYINPUT76), .A3(new_n241), .ZN(new_n242));
  NAND2_X1  g041(.A1(G225gat), .A2(G233gat), .ZN(new_n243));
  INV_X1    g042(.A(new_n243), .ZN(new_n244));
  INV_X1    g043(.A(KEYINPUT76), .ZN(new_n245));
  NAND3_X1  g044(.A1(new_n227), .A2(new_n239), .A3(new_n245), .ZN(new_n246));
  NAND3_X1  g045(.A1(new_n242), .A2(new_n244), .A3(new_n246), .ZN(new_n247));
  INV_X1    g046(.A(KEYINPUT3), .ZN(new_n248));
  AND3_X1   g047(.A1(new_n232), .A2(KEYINPUT75), .A3(new_n234), .ZN(new_n249));
  AOI21_X1  g048(.A(new_n234), .B1(new_n232), .B2(KEYINPUT75), .ZN(new_n250));
  OAI21_X1  g049(.A(new_n248), .B1(new_n249), .B2(new_n250), .ZN(new_n251));
  NAND3_X1  g050(.A1(new_n236), .A2(KEYINPUT3), .A3(new_n237), .ZN(new_n252));
  NAND3_X1  g051(.A1(new_n227), .A2(new_n251), .A3(new_n252), .ZN(new_n253));
  INV_X1    g052(.A(KEYINPUT4), .ZN(new_n254));
  OAI21_X1  g053(.A(new_n221), .B1(new_n222), .B2(new_n207), .ZN(new_n255));
  AOI21_X1  g054(.A(new_n219), .B1(new_n255), .B2(new_n206), .ZN(new_n256));
  AOI22_X1  g055(.A1(new_n256), .A2(new_n223), .B1(new_n225), .B2(new_n219), .ZN(new_n257));
  AOI21_X1  g056(.A(new_n254), .B1(new_n257), .B2(new_n238), .ZN(new_n258));
  NAND4_X1  g057(.A1(new_n238), .A2(new_n224), .A3(new_n254), .A4(new_n226), .ZN(new_n259));
  INV_X1    g058(.A(new_n259), .ZN(new_n260));
  OAI211_X1 g059(.A(new_n253), .B(new_n243), .C1(new_n258), .C2(new_n260), .ZN(new_n261));
  NAND3_X1  g060(.A1(new_n247), .A2(new_n261), .A3(KEYINPUT5), .ZN(new_n262));
  AND2_X1   g061(.A1(new_n253), .A2(new_n243), .ZN(new_n263));
  NAND2_X1  g062(.A1(new_n241), .A2(KEYINPUT4), .ZN(new_n264));
  INV_X1    g063(.A(KEYINPUT77), .ZN(new_n265));
  NAND3_X1  g064(.A1(new_n264), .A2(new_n265), .A3(new_n259), .ZN(new_n266));
  INV_X1    g065(.A(KEYINPUT5), .ZN(new_n267));
  NAND3_X1  g066(.A1(new_n241), .A2(KEYINPUT77), .A3(KEYINPUT4), .ZN(new_n268));
  NAND4_X1  g067(.A1(new_n263), .A2(new_n266), .A3(new_n267), .A4(new_n268), .ZN(new_n269));
  AOI21_X1  g068(.A(new_n205), .B1(new_n262), .B2(new_n269), .ZN(new_n270));
  INV_X1    g069(.A(new_n270), .ZN(new_n271));
  NAND3_X1  g070(.A1(new_n266), .A2(new_n268), .A3(new_n253), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n272), .A2(new_n244), .ZN(new_n273));
  INV_X1    g072(.A(KEYINPUT39), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n242), .A2(new_n246), .ZN(new_n275));
  AOI21_X1  g074(.A(new_n274), .B1(new_n275), .B2(new_n243), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n273), .A2(new_n276), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n277), .A2(KEYINPUT40), .ZN(new_n278));
  NAND3_X1  g077(.A1(new_n272), .A2(new_n274), .A3(new_n244), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n279), .A2(new_n205), .ZN(new_n280));
  OAI21_X1  g079(.A(new_n271), .B1(new_n278), .B2(new_n280), .ZN(new_n281));
  XNOR2_X1  g080(.A(KEYINPUT80), .B(KEYINPUT40), .ZN(new_n282));
  AND2_X1   g081(.A1(new_n279), .A2(new_n205), .ZN(new_n283));
  AOI21_X1  g082(.A(new_n282), .B1(new_n283), .B2(new_n277), .ZN(new_n284));
  NOR2_X1   g083(.A1(new_n281), .A2(new_n284), .ZN(new_n285));
  AND2_X1   g084(.A1(G211gat), .A2(G218gat), .ZN(new_n286));
  NOR2_X1   g085(.A1(new_n286), .A2(KEYINPUT22), .ZN(new_n287));
  INV_X1    g086(.A(new_n287), .ZN(new_n288));
  INV_X1    g087(.A(G197gat), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n289), .A2(KEYINPUT71), .ZN(new_n290));
  INV_X1    g089(.A(KEYINPUT71), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n291), .A2(G197gat), .ZN(new_n292));
  AND3_X1   g091(.A1(new_n290), .A2(new_n292), .A3(G204gat), .ZN(new_n293));
  AOI21_X1  g092(.A(G204gat), .B1(new_n290), .B2(new_n292), .ZN(new_n294));
  OAI21_X1  g093(.A(new_n288), .B1(new_n293), .B2(new_n294), .ZN(new_n295));
  NOR2_X1   g094(.A1(G211gat), .A2(G218gat), .ZN(new_n296));
  NOR2_X1   g095(.A1(new_n286), .A2(new_n296), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n295), .A2(new_n297), .ZN(new_n298));
  INV_X1    g097(.A(new_n297), .ZN(new_n299));
  OAI211_X1 g098(.A(new_n299), .B(new_n288), .C1(new_n293), .C2(new_n294), .ZN(new_n300));
  NAND3_X1  g099(.A1(new_n298), .A2(KEYINPUT72), .A3(new_n300), .ZN(new_n301));
  INV_X1    g100(.A(G204gat), .ZN(new_n302));
  NOR2_X1   g101(.A1(new_n291), .A2(G197gat), .ZN(new_n303));
  NOR2_X1   g102(.A1(new_n289), .A2(KEYINPUT71), .ZN(new_n304));
  OAI21_X1  g103(.A(new_n302), .B1(new_n303), .B2(new_n304), .ZN(new_n305));
  NAND3_X1  g104(.A1(new_n290), .A2(new_n292), .A3(G204gat), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n305), .A2(new_n306), .ZN(new_n307));
  AOI21_X1  g106(.A(new_n299), .B1(new_n307), .B2(new_n288), .ZN(new_n308));
  INV_X1    g107(.A(KEYINPUT72), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n308), .A2(new_n309), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n301), .A2(new_n310), .ZN(new_n311));
  INV_X1    g110(.A(G226gat), .ZN(new_n312));
  INV_X1    g111(.A(G233gat), .ZN(new_n313));
  NOR2_X1   g112(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  INV_X1    g113(.A(new_n314), .ZN(new_n315));
  INV_X1    g114(.A(KEYINPUT25), .ZN(new_n316));
  OAI21_X1  g115(.A(KEYINPUT23), .B1(G169gat), .B2(G176gat), .ZN(new_n317));
  INV_X1    g116(.A(new_n317), .ZN(new_n318));
  NOR3_X1   g117(.A1(KEYINPUT23), .A2(G169gat), .A3(G176gat), .ZN(new_n319));
  NAND3_X1  g118(.A1(KEYINPUT64), .A2(G169gat), .A3(G176gat), .ZN(new_n320));
  INV_X1    g119(.A(new_n320), .ZN(new_n321));
  AOI21_X1  g120(.A(KEYINPUT64), .B1(G169gat), .B2(G176gat), .ZN(new_n322));
  OAI22_X1  g121(.A1(new_n318), .A2(new_n319), .B1(new_n321), .B2(new_n322), .ZN(new_n323));
  NAND2_X1  g122(.A1(KEYINPUT24), .A2(G183gat), .ZN(new_n324));
  INV_X1    g123(.A(G190gat), .ZN(new_n325));
  NOR2_X1   g124(.A1(new_n324), .A2(new_n325), .ZN(new_n326));
  OAI21_X1  g125(.A(G190gat), .B1(KEYINPUT24), .B2(G183gat), .ZN(new_n327));
  AOI21_X1  g126(.A(new_n326), .B1(new_n324), .B2(new_n327), .ZN(new_n328));
  OAI21_X1  g127(.A(new_n316), .B1(new_n323), .B2(new_n328), .ZN(new_n329));
  NOR2_X1   g128(.A1(G169gat), .A2(G176gat), .ZN(new_n330));
  INV_X1    g129(.A(KEYINPUT23), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n330), .A2(new_n331), .ZN(new_n332));
  NAND2_X1  g131(.A1(G169gat), .A2(G176gat), .ZN(new_n333));
  INV_X1    g132(.A(KEYINPUT64), .ZN(new_n334));
  NAND2_X1  g133(.A1(new_n333), .A2(new_n334), .ZN(new_n335));
  AOI22_X1  g134(.A1(new_n332), .A2(new_n317), .B1(new_n335), .B2(new_n320), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n327), .A2(new_n324), .ZN(new_n337));
  OAI21_X1  g136(.A(new_n337), .B1(new_n325), .B2(new_n324), .ZN(new_n338));
  NAND3_X1  g137(.A1(new_n336), .A2(new_n338), .A3(KEYINPUT25), .ZN(new_n339));
  INV_X1    g138(.A(G183gat), .ZN(new_n340));
  NOR2_X1   g139(.A1(new_n340), .A2(new_n325), .ZN(new_n341));
  INV_X1    g140(.A(KEYINPUT26), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n330), .A2(new_n342), .ZN(new_n343));
  OAI21_X1  g142(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n344));
  AND2_X1   g143(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n335), .A2(new_n320), .ZN(new_n346));
  AOI21_X1  g145(.A(new_n341), .B1(new_n345), .B2(new_n346), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n340), .A2(KEYINPUT27), .ZN(new_n348));
  INV_X1    g147(.A(KEYINPUT27), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n349), .A2(G183gat), .ZN(new_n350));
  NAND3_X1  g149(.A1(new_n348), .A2(new_n350), .A3(new_n325), .ZN(new_n351));
  INV_X1    g150(.A(KEYINPUT28), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n351), .A2(new_n352), .ZN(new_n353));
  XNOR2_X1  g152(.A(KEYINPUT27), .B(G183gat), .ZN(new_n354));
  NAND3_X1  g153(.A1(new_n354), .A2(KEYINPUT28), .A3(new_n325), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n353), .A2(new_n355), .ZN(new_n356));
  AOI22_X1  g155(.A1(new_n329), .A2(new_n339), .B1(new_n347), .B2(new_n356), .ZN(new_n357));
  OAI21_X1  g156(.A(new_n315), .B1(new_n357), .B2(KEYINPUT29), .ZN(new_n358));
  NAND3_X1  g157(.A1(new_n346), .A2(new_n344), .A3(new_n343), .ZN(new_n359));
  INV_X1    g158(.A(new_n341), .ZN(new_n360));
  AOI21_X1  g159(.A(KEYINPUT28), .B1(new_n354), .B2(new_n325), .ZN(new_n361));
  AND4_X1   g160(.A1(KEYINPUT28), .A2(new_n348), .A3(new_n350), .A4(new_n325), .ZN(new_n362));
  OAI211_X1 g161(.A(new_n359), .B(new_n360), .C1(new_n361), .C2(new_n362), .ZN(new_n363));
  NOR3_X1   g162(.A1(new_n323), .A2(new_n328), .A3(new_n316), .ZN(new_n364));
  AOI21_X1  g163(.A(KEYINPUT25), .B1(new_n336), .B2(new_n338), .ZN(new_n365));
  OAI21_X1  g164(.A(new_n363), .B1(new_n364), .B2(new_n365), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n366), .A2(new_n314), .ZN(new_n367));
  AOI21_X1  g166(.A(KEYINPUT73), .B1(new_n358), .B2(new_n367), .ZN(new_n368));
  INV_X1    g167(.A(KEYINPUT29), .ZN(new_n369));
  AOI21_X1  g168(.A(new_n314), .B1(new_n366), .B2(new_n369), .ZN(new_n370));
  INV_X1    g169(.A(KEYINPUT73), .ZN(new_n371));
  NOR2_X1   g170(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  OAI21_X1  g171(.A(new_n311), .B1(new_n368), .B2(new_n372), .ZN(new_n373));
  XNOR2_X1  g172(.A(G8gat), .B(G36gat), .ZN(new_n374));
  XNOR2_X1  g173(.A(G64gat), .B(G92gat), .ZN(new_n375));
  XOR2_X1   g174(.A(new_n374), .B(new_n375), .Z(new_n376));
  NOR2_X1   g175(.A1(new_n357), .A2(new_n315), .ZN(new_n377));
  NOR3_X1   g176(.A1(new_n370), .A2(new_n377), .A3(new_n311), .ZN(new_n378));
  INV_X1    g177(.A(new_n378), .ZN(new_n379));
  NAND3_X1  g178(.A1(new_n373), .A2(new_n376), .A3(new_n379), .ZN(new_n380));
  INV_X1    g179(.A(KEYINPUT74), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n380), .A2(new_n381), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n382), .A2(KEYINPUT30), .ZN(new_n383));
  INV_X1    g182(.A(KEYINPUT30), .ZN(new_n384));
  NAND3_X1  g183(.A1(new_n380), .A2(new_n381), .A3(new_n384), .ZN(new_n385));
  AOI21_X1  g184(.A(new_n376), .B1(new_n373), .B2(new_n379), .ZN(new_n386));
  INV_X1    g185(.A(new_n386), .ZN(new_n387));
  NAND3_X1  g186(.A1(new_n383), .A2(new_n385), .A3(new_n387), .ZN(new_n388));
  XNOR2_X1  g187(.A(KEYINPUT31), .B(G50gat), .ZN(new_n389));
  INV_X1    g188(.A(new_n389), .ZN(new_n390));
  NAND2_X1  g189(.A1(G228gat), .A2(G233gat), .ZN(new_n391));
  XNOR2_X1  g190(.A(new_n391), .B(KEYINPUT79), .ZN(new_n392));
  AOI211_X1 g191(.A(new_n297), .B(new_n287), .C1(new_n305), .C2(new_n306), .ZN(new_n393));
  OAI21_X1  g192(.A(new_n369), .B1(new_n308), .B2(new_n393), .ZN(new_n394));
  AOI21_X1  g193(.A(new_n238), .B1(new_n394), .B2(new_n248), .ZN(new_n395));
  AOI22_X1  g194(.A1(new_n301), .A2(new_n310), .B1(new_n369), .B2(new_n251), .ZN(new_n396));
  OAI21_X1  g195(.A(new_n392), .B1(new_n395), .B2(new_n396), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n251), .A2(new_n369), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n311), .A2(new_n398), .ZN(new_n399));
  INV_X1    g198(.A(new_n391), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n399), .A2(new_n400), .ZN(new_n401));
  NAND3_X1  g200(.A1(new_n301), .A2(new_n369), .A3(new_n310), .ZN(new_n402));
  AOI21_X1  g201(.A(new_n238), .B1(new_n402), .B2(new_n248), .ZN(new_n403));
  OAI21_X1  g202(.A(new_n397), .B1(new_n401), .B2(new_n403), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n404), .A2(G22gat), .ZN(new_n405));
  INV_X1    g204(.A(G22gat), .ZN(new_n406));
  OAI211_X1 g205(.A(new_n397), .B(new_n406), .C1(new_n401), .C2(new_n403), .ZN(new_n407));
  XNOR2_X1  g206(.A(G78gat), .B(G106gat), .ZN(new_n408));
  INV_X1    g207(.A(new_n408), .ZN(new_n409));
  AND3_X1   g208(.A1(new_n405), .A2(new_n407), .A3(new_n409), .ZN(new_n410));
  AOI21_X1  g209(.A(new_n409), .B1(new_n405), .B2(new_n407), .ZN(new_n411));
  OAI21_X1  g210(.A(new_n390), .B1(new_n410), .B2(new_n411), .ZN(new_n412));
  INV_X1    g211(.A(new_n407), .ZN(new_n413));
  NAND2_X1  g212(.A1(new_n402), .A2(new_n248), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n414), .A2(new_n239), .ZN(new_n415));
  NOR2_X1   g214(.A1(new_n396), .A2(new_n391), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n415), .A2(new_n416), .ZN(new_n417));
  AOI21_X1  g216(.A(new_n406), .B1(new_n417), .B2(new_n397), .ZN(new_n418));
  OAI21_X1  g217(.A(new_n408), .B1(new_n413), .B2(new_n418), .ZN(new_n419));
  NAND3_X1  g218(.A1(new_n405), .A2(new_n407), .A3(new_n409), .ZN(new_n420));
  NAND3_X1  g219(.A1(new_n419), .A2(new_n389), .A3(new_n420), .ZN(new_n421));
  AOI22_X1  g220(.A1(new_n285), .A2(new_n388), .B1(new_n412), .B2(new_n421), .ZN(new_n422));
  INV_X1    g221(.A(KEYINPUT78), .ZN(new_n423));
  NAND4_X1  g222(.A1(new_n262), .A2(new_n423), .A3(new_n269), .A4(new_n205), .ZN(new_n424));
  INV_X1    g223(.A(KEYINPUT6), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n426), .A2(new_n271), .ZN(new_n427));
  NAND3_X1  g226(.A1(new_n262), .A2(new_n269), .A3(new_n205), .ZN(new_n428));
  AOI21_X1  g227(.A(new_n270), .B1(KEYINPUT78), .B2(new_n428), .ZN(new_n429));
  OAI21_X1  g228(.A(new_n427), .B1(new_n429), .B2(KEYINPUT6), .ZN(new_n430));
  INV_X1    g229(.A(new_n311), .ZN(new_n431));
  OAI21_X1  g230(.A(new_n371), .B1(new_n370), .B2(new_n377), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n358), .A2(KEYINPUT73), .ZN(new_n433));
  AOI21_X1  g232(.A(new_n431), .B1(new_n432), .B2(new_n433), .ZN(new_n434));
  OAI21_X1  g233(.A(KEYINPUT37), .B1(new_n434), .B2(new_n378), .ZN(new_n435));
  INV_X1    g234(.A(KEYINPUT37), .ZN(new_n436));
  NOR2_X1   g235(.A1(new_n376), .A2(new_n436), .ZN(new_n437));
  OAI21_X1  g236(.A(new_n435), .B1(new_n386), .B2(new_n437), .ZN(new_n438));
  NOR2_X1   g237(.A1(new_n434), .A2(new_n378), .ZN(new_n439));
  AOI22_X1  g238(.A1(new_n438), .A2(KEYINPUT38), .B1(new_n376), .B2(new_n439), .ZN(new_n440));
  INV_X1    g239(.A(KEYINPUT82), .ZN(new_n441));
  INV_X1    g240(.A(KEYINPUT38), .ZN(new_n442));
  OAI21_X1  g241(.A(new_n442), .B1(new_n386), .B2(new_n437), .ZN(new_n443));
  INV_X1    g242(.A(KEYINPUT81), .ZN(new_n444));
  NAND4_X1  g243(.A1(new_n432), .A2(new_n444), .A3(new_n431), .A4(new_n433), .ZN(new_n445));
  NOR3_X1   g244(.A1(new_n368), .A2(new_n372), .A3(new_n311), .ZN(new_n446));
  OAI21_X1  g245(.A(new_n311), .B1(new_n370), .B2(new_n377), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n447), .A2(KEYINPUT81), .ZN(new_n448));
  OAI211_X1 g247(.A(KEYINPUT37), .B(new_n445), .C1(new_n446), .C2(new_n448), .ZN(new_n449));
  INV_X1    g248(.A(new_n449), .ZN(new_n450));
  OAI21_X1  g249(.A(new_n441), .B1(new_n443), .B2(new_n450), .ZN(new_n451));
  AOI21_X1  g250(.A(new_n376), .B1(new_n439), .B2(new_n436), .ZN(new_n452));
  NAND4_X1  g251(.A1(new_n452), .A2(new_n449), .A3(KEYINPUT82), .A4(new_n442), .ZN(new_n453));
  NAND4_X1  g252(.A1(new_n430), .A2(new_n440), .A3(new_n451), .A4(new_n453), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n422), .A2(new_n454), .ZN(new_n455));
  INV_X1    g254(.A(KEYINPUT83), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n455), .A2(new_n456), .ZN(new_n457));
  NAND3_X1  g256(.A1(new_n422), .A2(new_n454), .A3(KEYINPUT83), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n366), .A2(new_n257), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n357), .A2(new_n227), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  INV_X1    g261(.A(KEYINPUT34), .ZN(new_n463));
  NAND2_X1  g262(.A1(G227gat), .A2(G233gat), .ZN(new_n464));
  NAND3_X1  g263(.A1(new_n462), .A2(new_n463), .A3(new_n464), .ZN(new_n465));
  OR2_X1    g264(.A1(new_n465), .A2(KEYINPUT70), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n462), .A2(new_n464), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n467), .A2(KEYINPUT34), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n465), .A2(KEYINPUT70), .ZN(new_n469));
  NAND3_X1  g268(.A1(new_n466), .A2(new_n468), .A3(new_n469), .ZN(new_n470));
  INV_X1    g269(.A(new_n470), .ZN(new_n471));
  INV_X1    g270(.A(KEYINPUT32), .ZN(new_n472));
  INV_X1    g271(.A(new_n464), .ZN(new_n473));
  NAND3_X1  g272(.A1(new_n460), .A2(new_n461), .A3(new_n473), .ZN(new_n474));
  INV_X1    g273(.A(KEYINPUT67), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  NAND4_X1  g275(.A1(new_n460), .A2(new_n461), .A3(KEYINPUT67), .A4(new_n473), .ZN(new_n477));
  AOI21_X1  g276(.A(new_n472), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  XNOR2_X1  g277(.A(G15gat), .B(G43gat), .ZN(new_n479));
  XNOR2_X1  g278(.A(G71gat), .B(G99gat), .ZN(new_n480));
  XOR2_X1   g279(.A(new_n479), .B(new_n480), .Z(new_n481));
  OAI21_X1  g280(.A(KEYINPUT33), .B1(new_n481), .B2(KEYINPUT69), .ZN(new_n482));
  AOI21_X1  g281(.A(new_n482), .B1(KEYINPUT69), .B2(new_n481), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n478), .A2(new_n483), .ZN(new_n484));
  INV_X1    g283(.A(new_n481), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n476), .A2(new_n477), .ZN(new_n486));
  INV_X1    g285(.A(KEYINPUT33), .ZN(new_n487));
  AOI21_X1  g286(.A(new_n485), .B1(new_n486), .B2(new_n487), .ZN(new_n488));
  INV_X1    g287(.A(KEYINPUT68), .ZN(new_n489));
  AOI21_X1  g288(.A(new_n484), .B1(new_n488), .B2(new_n489), .ZN(new_n490));
  AOI21_X1  g289(.A(new_n478), .B1(new_n488), .B2(KEYINPUT68), .ZN(new_n491));
  OAI21_X1  g290(.A(new_n471), .B1(new_n490), .B2(new_n491), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n486), .A2(new_n487), .ZN(new_n493));
  NAND3_X1  g292(.A1(new_n493), .A2(KEYINPUT68), .A3(new_n481), .ZN(new_n494));
  INV_X1    g293(.A(new_n478), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  NAND3_X1  g295(.A1(new_n493), .A2(new_n489), .A3(new_n481), .ZN(new_n497));
  AND2_X1   g296(.A1(new_n478), .A2(new_n483), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  NAND3_X1  g298(.A1(new_n496), .A2(new_n499), .A3(new_n470), .ZN(new_n500));
  AND3_X1   g299(.A1(new_n492), .A2(new_n500), .A3(KEYINPUT36), .ZN(new_n501));
  AOI21_X1  g300(.A(KEYINPUT36), .B1(new_n492), .B2(new_n500), .ZN(new_n502));
  NOR2_X1   g301(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  NOR2_X1   g302(.A1(new_n430), .A2(new_n388), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n412), .A2(new_n421), .ZN(new_n505));
  NOR2_X1   g304(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  NOR2_X1   g305(.A1(new_n503), .A2(new_n506), .ZN(new_n507));
  NOR3_X1   g306(.A1(new_n410), .A2(new_n411), .A3(new_n390), .ZN(new_n508));
  AOI21_X1  g307(.A(new_n389), .B1(new_n419), .B2(new_n420), .ZN(new_n509));
  OAI211_X1 g308(.A(new_n500), .B(new_n492), .C1(new_n508), .C2(new_n509), .ZN(new_n510));
  AND2_X1   g309(.A1(new_n428), .A2(KEYINPUT78), .ZN(new_n511));
  OAI21_X1  g310(.A(new_n425), .B1(new_n511), .B2(new_n270), .ZN(new_n512));
  AOI21_X1  g311(.A(new_n386), .B1(new_n382), .B2(KEYINPUT30), .ZN(new_n513));
  NAND4_X1  g312(.A1(new_n512), .A2(new_n427), .A3(new_n513), .A4(new_n385), .ZN(new_n514));
  OAI21_X1  g313(.A(KEYINPUT35), .B1(new_n510), .B2(new_n514), .ZN(new_n515));
  NOR3_X1   g314(.A1(new_n490), .A2(new_n491), .A3(new_n471), .ZN(new_n516));
  AOI21_X1  g315(.A(new_n470), .B1(new_n496), .B2(new_n499), .ZN(new_n517));
  NOR2_X1   g316(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  INV_X1    g317(.A(KEYINPUT35), .ZN(new_n519));
  NAND4_X1  g318(.A1(new_n518), .A2(new_n504), .A3(new_n519), .A4(new_n505), .ZN(new_n520));
  AOI22_X1  g319(.A1(new_n459), .A2(new_n507), .B1(new_n515), .B2(new_n520), .ZN(new_n521));
  INV_X1    g320(.A(G8gat), .ZN(new_n522));
  XNOR2_X1  g321(.A(G15gat), .B(G22gat), .ZN(new_n523));
  INV_X1    g322(.A(G1gat), .ZN(new_n524));
  NOR2_X1   g323(.A1(new_n524), .A2(KEYINPUT88), .ZN(new_n525));
  INV_X1    g324(.A(KEYINPUT88), .ZN(new_n526));
  OAI21_X1  g325(.A(KEYINPUT16), .B1(new_n526), .B2(G1gat), .ZN(new_n527));
  OAI21_X1  g326(.A(new_n523), .B1(new_n525), .B2(new_n527), .ZN(new_n528));
  INV_X1    g327(.A(KEYINPUT89), .ZN(new_n529));
  AOI21_X1  g328(.A(new_n522), .B1(new_n528), .B2(new_n529), .ZN(new_n530));
  OAI21_X1  g329(.A(new_n528), .B1(G1gat), .B2(new_n523), .ZN(new_n531));
  XOR2_X1   g330(.A(new_n530), .B(new_n531), .Z(new_n532));
  XNOR2_X1  g331(.A(new_n532), .B(KEYINPUT90), .ZN(new_n533));
  XOR2_X1   g332(.A(G43gat), .B(G50gat), .Z(new_n534));
  INV_X1    g333(.A(KEYINPUT15), .ZN(new_n535));
  OR2_X1    g334(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  OAI21_X1  g335(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n537));
  OR3_X1    g336(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n538));
  AOI22_X1  g337(.A1(new_n534), .A2(new_n535), .B1(new_n537), .B2(new_n538), .ZN(new_n539));
  XNOR2_X1  g338(.A(KEYINPUT86), .B(G29gat), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n540), .A2(G36gat), .ZN(new_n541));
  NAND3_X1  g340(.A1(new_n536), .A2(new_n539), .A3(new_n541), .ZN(new_n542));
  OR2_X1    g341(.A1(new_n537), .A2(KEYINPUT85), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n537), .A2(KEYINPUT85), .ZN(new_n544));
  NAND3_X1  g343(.A1(new_n543), .A2(new_n538), .A3(new_n544), .ZN(new_n545));
  AND2_X1   g344(.A1(new_n545), .A2(new_n541), .ZN(new_n546));
  OAI21_X1  g345(.A(new_n542), .B1(new_n546), .B2(new_n536), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n533), .A2(new_n547), .ZN(new_n548));
  INV_X1    g347(.A(KEYINPUT91), .ZN(new_n549));
  XNOR2_X1  g348(.A(new_n548), .B(new_n549), .ZN(new_n550));
  OAI21_X1  g349(.A(new_n550), .B1(new_n547), .B2(new_n533), .ZN(new_n551));
  NAND2_X1  g350(.A1(G229gat), .A2(G233gat), .ZN(new_n552));
  XOR2_X1   g351(.A(new_n552), .B(KEYINPUT13), .Z(new_n553));
  NAND2_X1  g352(.A1(new_n551), .A2(new_n553), .ZN(new_n554));
  INV_X1    g353(.A(KEYINPUT87), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n547), .A2(new_n555), .ZN(new_n556));
  XOR2_X1   g355(.A(new_n556), .B(KEYINPUT17), .Z(new_n557));
  NAND2_X1  g356(.A1(new_n557), .A2(new_n532), .ZN(new_n558));
  NAND3_X1  g357(.A1(new_n550), .A2(new_n552), .A3(new_n558), .ZN(new_n559));
  INV_X1    g358(.A(KEYINPUT18), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  NAND4_X1  g360(.A1(new_n550), .A2(KEYINPUT18), .A3(new_n552), .A4(new_n558), .ZN(new_n562));
  NAND3_X1  g361(.A1(new_n554), .A2(new_n561), .A3(new_n562), .ZN(new_n563));
  XNOR2_X1  g362(.A(G113gat), .B(G141gat), .ZN(new_n564));
  XNOR2_X1  g363(.A(new_n564), .B(G197gat), .ZN(new_n565));
  XOR2_X1   g364(.A(KEYINPUT11), .B(G169gat), .Z(new_n566));
  XNOR2_X1  g365(.A(new_n565), .B(new_n566), .ZN(new_n567));
  XNOR2_X1  g366(.A(KEYINPUT84), .B(KEYINPUT12), .ZN(new_n568));
  XOR2_X1   g367(.A(new_n567), .B(new_n568), .Z(new_n569));
  INV_X1    g368(.A(new_n569), .ZN(new_n570));
  NAND2_X1  g369(.A1(new_n563), .A2(new_n570), .ZN(new_n571));
  NAND4_X1  g370(.A1(new_n554), .A2(new_n561), .A3(new_n569), .A4(new_n562), .ZN(new_n572));
  NAND2_X1  g371(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  NAND2_X1  g372(.A1(new_n573), .A2(KEYINPUT92), .ZN(new_n574));
  INV_X1    g373(.A(KEYINPUT92), .ZN(new_n575));
  NAND3_X1  g374(.A1(new_n571), .A2(new_n575), .A3(new_n572), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n574), .A2(new_n576), .ZN(new_n577));
  NOR2_X1   g376(.A1(new_n521), .A2(new_n577), .ZN(new_n578));
  XNOR2_X1  g377(.A(G190gat), .B(G218gat), .ZN(new_n579));
  INV_X1    g378(.A(KEYINPUT98), .ZN(new_n580));
  NAND3_X1  g379(.A1(new_n580), .A2(G85gat), .A3(G92gat), .ZN(new_n581));
  XNOR2_X1  g380(.A(new_n581), .B(KEYINPUT7), .ZN(new_n582));
  INV_X1    g381(.A(KEYINPUT8), .ZN(new_n583));
  NAND2_X1  g382(.A1(G99gat), .A2(G106gat), .ZN(new_n584));
  AOI21_X1  g383(.A(new_n583), .B1(new_n584), .B2(KEYINPUT99), .ZN(new_n585));
  OAI21_X1  g384(.A(new_n585), .B1(KEYINPUT99), .B2(new_n584), .ZN(new_n586));
  XNOR2_X1  g385(.A(KEYINPUT100), .B(G92gat), .ZN(new_n587));
  OAI211_X1 g386(.A(new_n582), .B(new_n586), .C1(G85gat), .C2(new_n587), .ZN(new_n588));
  XNOR2_X1  g387(.A(new_n588), .B(KEYINPUT101), .ZN(new_n589));
  XOR2_X1   g388(.A(G99gat), .B(G106gat), .Z(new_n590));
  XNOR2_X1  g389(.A(new_n589), .B(new_n590), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n591), .A2(KEYINPUT102), .ZN(new_n592));
  INV_X1    g391(.A(new_n590), .ZN(new_n593));
  XNOR2_X1  g392(.A(new_n589), .B(new_n593), .ZN(new_n594));
  INV_X1    g393(.A(KEYINPUT102), .ZN(new_n595));
  NAND2_X1  g394(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  NAND3_X1  g395(.A1(new_n592), .A2(new_n596), .A3(new_n557), .ZN(new_n597));
  INV_X1    g396(.A(KEYINPUT103), .ZN(new_n598));
  AND2_X1   g397(.A1(G232gat), .A2(G233gat), .ZN(new_n599));
  AOI22_X1  g398(.A1(new_n591), .A2(new_n547), .B1(KEYINPUT41), .B2(new_n599), .ZN(new_n600));
  NAND3_X1  g399(.A1(new_n597), .A2(new_n598), .A3(new_n600), .ZN(new_n601));
  INV_X1    g400(.A(new_n601), .ZN(new_n602));
  AOI21_X1  g401(.A(new_n598), .B1(new_n597), .B2(new_n600), .ZN(new_n603));
  OAI21_X1  g402(.A(new_n579), .B1(new_n602), .B2(new_n603), .ZN(new_n604));
  INV_X1    g403(.A(new_n603), .ZN(new_n605));
  INV_X1    g404(.A(new_n579), .ZN(new_n606));
  NAND3_X1  g405(.A1(new_n605), .A2(new_n601), .A3(new_n606), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n604), .A2(new_n607), .ZN(new_n608));
  NOR2_X1   g407(.A1(new_n599), .A2(KEYINPUT41), .ZN(new_n609));
  XNOR2_X1  g408(.A(new_n609), .B(KEYINPUT97), .ZN(new_n610));
  XOR2_X1   g409(.A(G134gat), .B(G162gat), .Z(new_n611));
  XNOR2_X1  g410(.A(new_n610), .B(new_n611), .ZN(new_n612));
  NAND2_X1  g411(.A1(new_n612), .A2(KEYINPUT104), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n608), .A2(new_n613), .ZN(new_n614));
  XNOR2_X1  g413(.A(new_n612), .B(KEYINPUT104), .ZN(new_n615));
  NAND3_X1  g414(.A1(new_n604), .A2(new_n607), .A3(new_n615), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n614), .A2(new_n616), .ZN(new_n617));
  INV_X1    g416(.A(new_n617), .ZN(new_n618));
  AND2_X1   g417(.A1(G71gat), .A2(G78gat), .ZN(new_n619));
  INV_X1    g418(.A(new_n619), .ZN(new_n620));
  NOR2_X1   g419(.A1(G71gat), .A2(G78gat), .ZN(new_n621));
  INV_X1    g420(.A(new_n621), .ZN(new_n622));
  INV_X1    g421(.A(G57gat), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n623), .A2(G64gat), .ZN(new_n624));
  INV_X1    g423(.A(G64gat), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n625), .A2(G57gat), .ZN(new_n626));
  AND2_X1   g425(.A1(new_n624), .A2(new_n626), .ZN(new_n627));
  INV_X1    g426(.A(KEYINPUT9), .ZN(new_n628));
  OAI211_X1 g427(.A(new_n620), .B(new_n622), .C1(new_n627), .C2(new_n628), .ZN(new_n629));
  OR2_X1    g428(.A1(new_n629), .A2(KEYINPUT93), .ZN(new_n630));
  OAI21_X1  g429(.A(new_n620), .B1(new_n622), .B2(new_n628), .ZN(new_n631));
  NAND2_X1  g430(.A1(new_n626), .A2(KEYINPUT94), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n632), .A2(new_n624), .ZN(new_n633));
  NOR2_X1   g432(.A1(new_n626), .A2(KEYINPUT94), .ZN(new_n634));
  OAI21_X1  g433(.A(new_n631), .B1(new_n633), .B2(new_n634), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n629), .A2(KEYINPUT93), .ZN(new_n636));
  NAND3_X1  g435(.A1(new_n630), .A2(new_n635), .A3(new_n636), .ZN(new_n637));
  XNOR2_X1  g436(.A(KEYINPUT95), .B(KEYINPUT21), .ZN(new_n638));
  NAND2_X1  g437(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  NAND2_X1  g438(.A1(G231gat), .A2(G233gat), .ZN(new_n640));
  XNOR2_X1  g439(.A(new_n639), .B(new_n640), .ZN(new_n641));
  XOR2_X1   g440(.A(G127gat), .B(G155gat), .Z(new_n642));
  XNOR2_X1  g441(.A(new_n642), .B(KEYINPUT20), .ZN(new_n643));
  XNOR2_X1  g442(.A(new_n641), .B(new_n643), .ZN(new_n644));
  XOR2_X1   g443(.A(G183gat), .B(G211gat), .Z(new_n645));
  XNOR2_X1  g444(.A(new_n644), .B(new_n645), .ZN(new_n646));
  INV_X1    g445(.A(new_n533), .ZN(new_n647));
  INV_X1    g446(.A(KEYINPUT21), .ZN(new_n648));
  OAI21_X1  g447(.A(new_n647), .B1(new_n648), .B2(new_n637), .ZN(new_n649));
  XNOR2_X1  g448(.A(KEYINPUT96), .B(KEYINPUT19), .ZN(new_n650));
  XNOR2_X1  g449(.A(new_n649), .B(new_n650), .ZN(new_n651));
  XNOR2_X1  g450(.A(new_n646), .B(new_n651), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n618), .A2(new_n652), .ZN(new_n653));
  INV_X1    g452(.A(G230gat), .ZN(new_n654));
  NOR2_X1   g453(.A1(new_n654), .A2(new_n313), .ZN(new_n655));
  OR2_X1    g454(.A1(new_n594), .A2(new_n637), .ZN(new_n656));
  INV_X1    g455(.A(KEYINPUT10), .ZN(new_n657));
  NAND2_X1  g456(.A1(new_n594), .A2(new_n637), .ZN(new_n658));
  NAND3_X1  g457(.A1(new_n656), .A2(new_n657), .A3(new_n658), .ZN(new_n659));
  OR3_X1    g458(.A1(new_n594), .A2(new_n657), .A3(new_n637), .ZN(new_n660));
  AOI21_X1  g459(.A(new_n655), .B1(new_n659), .B2(new_n660), .ZN(new_n661));
  INV_X1    g460(.A(new_n661), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n656), .A2(new_n658), .ZN(new_n663));
  NAND2_X1  g462(.A1(new_n663), .A2(new_n655), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n662), .A2(new_n664), .ZN(new_n665));
  XOR2_X1   g464(.A(G120gat), .B(G148gat), .Z(new_n666));
  XNOR2_X1  g465(.A(new_n666), .B(KEYINPUT105), .ZN(new_n667));
  XNOR2_X1  g466(.A(G176gat), .B(G204gat), .ZN(new_n668));
  XOR2_X1   g467(.A(new_n667), .B(new_n668), .Z(new_n669));
  NAND2_X1  g468(.A1(new_n665), .A2(new_n669), .ZN(new_n670));
  INV_X1    g469(.A(new_n669), .ZN(new_n671));
  NAND3_X1  g470(.A1(new_n662), .A2(new_n664), .A3(new_n671), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n670), .A2(new_n672), .ZN(new_n673));
  NOR2_X1   g472(.A1(new_n653), .A2(new_n673), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n578), .A2(new_n674), .ZN(new_n675));
  INV_X1    g474(.A(new_n430), .ZN(new_n676));
  NOR2_X1   g475(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  XNOR2_X1  g476(.A(new_n677), .B(new_n524), .ZN(G1324gat));
  INV_X1    g477(.A(new_n388), .ZN(new_n679));
  NOR2_X1   g478(.A1(new_n675), .A2(new_n679), .ZN(new_n680));
  XOR2_X1   g479(.A(KEYINPUT16), .B(G8gat), .Z(new_n681));
  NAND2_X1  g480(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  OAI21_X1  g481(.A(new_n682), .B1(new_n522), .B2(new_n680), .ZN(new_n683));
  MUX2_X1   g482(.A(new_n682), .B(new_n683), .S(KEYINPUT42), .Z(G1325gat));
  INV_X1    g483(.A(KEYINPUT106), .ZN(new_n685));
  NOR3_X1   g484(.A1(new_n501), .A2(new_n502), .A3(new_n685), .ZN(new_n686));
  INV_X1    g485(.A(KEYINPUT36), .ZN(new_n687));
  OAI21_X1  g486(.A(new_n687), .B1(new_n516), .B2(new_n517), .ZN(new_n688));
  NAND3_X1  g487(.A1(new_n492), .A2(new_n500), .A3(KEYINPUT36), .ZN(new_n689));
  AOI21_X1  g488(.A(KEYINPUT106), .B1(new_n688), .B2(new_n689), .ZN(new_n690));
  NOR2_X1   g489(.A1(new_n686), .A2(new_n690), .ZN(new_n691));
  XOR2_X1   g490(.A(new_n691), .B(KEYINPUT107), .Z(new_n692));
  OAI21_X1  g491(.A(G15gat), .B1(new_n675), .B2(new_n692), .ZN(new_n693));
  INV_X1    g492(.A(new_n518), .ZN(new_n694));
  OR2_X1    g493(.A1(new_n694), .A2(G15gat), .ZN(new_n695));
  OAI21_X1  g494(.A(new_n693), .B1(new_n675), .B2(new_n695), .ZN(G1326gat));
  NOR2_X1   g495(.A1(new_n675), .A2(new_n505), .ZN(new_n697));
  XOR2_X1   g496(.A(KEYINPUT43), .B(G22gat), .Z(new_n698));
  XNOR2_X1  g497(.A(new_n697), .B(new_n698), .ZN(G1327gat));
  INV_X1    g498(.A(new_n673), .ZN(new_n700));
  INV_X1    g499(.A(new_n652), .ZN(new_n701));
  NAND3_X1  g500(.A1(new_n617), .A2(new_n700), .A3(new_n701), .ZN(new_n702));
  XOR2_X1   g501(.A(new_n702), .B(KEYINPUT108), .Z(new_n703));
  NAND2_X1  g502(.A1(new_n703), .A2(new_n578), .ZN(new_n704));
  NOR3_X1   g503(.A1(new_n704), .A2(new_n676), .A3(new_n540), .ZN(new_n705));
  XOR2_X1   g504(.A(new_n705), .B(KEYINPUT45), .Z(new_n706));
  OAI21_X1  g505(.A(KEYINPUT44), .B1(new_n521), .B2(new_n618), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n515), .A2(new_n520), .ZN(new_n708));
  NAND2_X1  g507(.A1(new_n708), .A2(KEYINPUT110), .ZN(new_n709));
  INV_X1    g508(.A(KEYINPUT110), .ZN(new_n710));
  NAND3_X1  g509(.A1(new_n515), .A2(new_n520), .A3(new_n710), .ZN(new_n711));
  INV_X1    g510(.A(new_n506), .ZN(new_n712));
  OAI21_X1  g511(.A(new_n712), .B1(new_n686), .B2(new_n690), .ZN(new_n713));
  AND3_X1   g512(.A1(new_n422), .A2(new_n454), .A3(KEYINPUT83), .ZN(new_n714));
  AOI21_X1  g513(.A(KEYINPUT83), .B1(new_n422), .B2(new_n454), .ZN(new_n715));
  NOR2_X1   g514(.A1(new_n714), .A2(new_n715), .ZN(new_n716));
  OAI211_X1 g515(.A(new_n709), .B(new_n711), .C1(new_n713), .C2(new_n716), .ZN(new_n717));
  NAND2_X1  g516(.A1(new_n617), .A2(KEYINPUT111), .ZN(new_n718));
  INV_X1    g517(.A(KEYINPUT111), .ZN(new_n719));
  NAND3_X1  g518(.A1(new_n614), .A2(new_n719), .A3(new_n616), .ZN(new_n720));
  AOI21_X1  g519(.A(KEYINPUT44), .B1(new_n718), .B2(new_n720), .ZN(new_n721));
  AND3_X1   g520(.A1(new_n717), .A2(KEYINPUT112), .A3(new_n721), .ZN(new_n722));
  AOI21_X1  g521(.A(KEYINPUT112), .B1(new_n717), .B2(new_n721), .ZN(new_n723));
  OAI21_X1  g522(.A(new_n707), .B1(new_n722), .B2(new_n723), .ZN(new_n724));
  XNOR2_X1  g523(.A(new_n673), .B(KEYINPUT109), .ZN(new_n725));
  INV_X1    g524(.A(new_n573), .ZN(new_n726));
  NOR3_X1   g525(.A1(new_n725), .A2(new_n726), .A3(new_n652), .ZN(new_n727));
  AND2_X1   g526(.A1(new_n724), .A2(new_n727), .ZN(new_n728));
  INV_X1    g527(.A(new_n728), .ZN(new_n729));
  OAI21_X1  g528(.A(new_n540), .B1(new_n729), .B2(new_n676), .ZN(new_n730));
  NAND2_X1  g529(.A1(new_n706), .A2(new_n730), .ZN(G1328gat));
  OAI21_X1  g530(.A(G36gat), .B1(new_n729), .B2(new_n679), .ZN(new_n732));
  NOR3_X1   g531(.A1(new_n704), .A2(G36gat), .A3(new_n679), .ZN(new_n733));
  XNOR2_X1  g532(.A(new_n733), .B(KEYINPUT46), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n732), .A2(new_n734), .ZN(new_n735));
  XNOR2_X1  g534(.A(new_n735), .B(KEYINPUT113), .ZN(G1329gat));
  INV_X1    g535(.A(new_n691), .ZN(new_n737));
  OAI21_X1  g536(.A(G43gat), .B1(new_n729), .B2(new_n737), .ZN(new_n738));
  NOR3_X1   g537(.A1(new_n704), .A2(G43gat), .A3(new_n694), .ZN(new_n739));
  INV_X1    g538(.A(KEYINPUT47), .ZN(new_n740));
  NOR2_X1   g539(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  NAND2_X1  g540(.A1(new_n738), .A2(new_n741), .ZN(new_n742));
  INV_X1    g541(.A(new_n692), .ZN(new_n743));
  NAND2_X1  g542(.A1(new_n728), .A2(new_n743), .ZN(new_n744));
  AND3_X1   g543(.A1(new_n744), .A2(KEYINPUT114), .A3(G43gat), .ZN(new_n745));
  AOI21_X1  g544(.A(KEYINPUT114), .B1(new_n744), .B2(G43gat), .ZN(new_n746));
  NOR3_X1   g545(.A1(new_n745), .A2(new_n746), .A3(new_n739), .ZN(new_n747));
  OAI21_X1  g546(.A(new_n742), .B1(new_n747), .B2(KEYINPUT47), .ZN(G1330gat));
  NOR2_X1   g547(.A1(new_n505), .A2(G50gat), .ZN(new_n749));
  XOR2_X1   g548(.A(new_n749), .B(KEYINPUT115), .Z(new_n750));
  NOR2_X1   g549(.A1(new_n704), .A2(new_n750), .ZN(new_n751));
  INV_X1    g550(.A(new_n505), .ZN(new_n752));
  NAND2_X1  g551(.A1(new_n728), .A2(new_n752), .ZN(new_n753));
  AOI21_X1  g552(.A(new_n751), .B1(new_n753), .B2(G50gat), .ZN(new_n754));
  XNOR2_X1  g553(.A(new_n754), .B(KEYINPUT48), .ZN(G1331gat));
  INV_X1    g554(.A(new_n725), .ZN(new_n756));
  NOR3_X1   g555(.A1(new_n756), .A2(new_n653), .A3(new_n573), .ZN(new_n757));
  AND2_X1   g556(.A1(new_n757), .A2(new_n717), .ZN(new_n758));
  NAND2_X1  g557(.A1(new_n758), .A2(new_n430), .ZN(new_n759));
  XNOR2_X1  g558(.A(new_n759), .B(G57gat), .ZN(G1332gat));
  AOI21_X1  g559(.A(new_n679), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n761));
  NAND2_X1  g560(.A1(new_n758), .A2(new_n761), .ZN(new_n762));
  XNOR2_X1  g561(.A(new_n762), .B(KEYINPUT116), .ZN(new_n763));
  NOR2_X1   g562(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n764));
  XNOR2_X1  g563(.A(new_n763), .B(new_n764), .ZN(G1333gat));
  NAND2_X1  g564(.A1(new_n758), .A2(new_n743), .ZN(new_n766));
  NOR2_X1   g565(.A1(new_n694), .A2(G71gat), .ZN(new_n767));
  AOI22_X1  g566(.A1(new_n766), .A2(G71gat), .B1(new_n758), .B2(new_n767), .ZN(new_n768));
  XNOR2_X1  g567(.A(new_n768), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g568(.A1(new_n758), .A2(new_n752), .ZN(new_n770));
  XNOR2_X1  g569(.A(new_n770), .B(G78gat), .ZN(G1335gat));
  NOR3_X1   g570(.A1(new_n573), .A2(new_n700), .A3(new_n652), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n724), .A2(new_n772), .ZN(new_n773));
  OAI21_X1  g572(.A(G85gat), .B1(new_n773), .B2(new_n676), .ZN(new_n774));
  INV_X1    g573(.A(KEYINPUT117), .ZN(new_n775));
  NAND3_X1  g574(.A1(new_n726), .A2(new_n617), .A3(new_n701), .ZN(new_n776));
  AND3_X1   g575(.A1(new_n515), .A2(new_n520), .A3(new_n710), .ZN(new_n777));
  AOI21_X1  g576(.A(new_n710), .B1(new_n515), .B2(new_n520), .ZN(new_n778));
  NOR2_X1   g577(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  OAI21_X1  g578(.A(new_n685), .B1(new_n501), .B2(new_n502), .ZN(new_n780));
  NAND3_X1  g579(.A1(new_n688), .A2(KEYINPUT106), .A3(new_n689), .ZN(new_n781));
  AOI21_X1  g580(.A(new_n506), .B1(new_n780), .B2(new_n781), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n459), .A2(new_n782), .ZN(new_n783));
  AOI21_X1  g582(.A(new_n776), .B1(new_n779), .B2(new_n783), .ZN(new_n784));
  AOI21_X1  g583(.A(new_n775), .B1(new_n784), .B2(KEYINPUT51), .ZN(new_n785));
  INV_X1    g584(.A(new_n776), .ZN(new_n786));
  AND4_X1   g585(.A1(new_n775), .A2(new_n717), .A3(KEYINPUT51), .A4(new_n786), .ZN(new_n787));
  NOR2_X1   g586(.A1(new_n785), .A2(new_n787), .ZN(new_n788));
  INV_X1    g587(.A(KEYINPUT51), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n717), .A2(new_n786), .ZN(new_n790));
  AOI21_X1  g589(.A(new_n788), .B1(new_n789), .B2(new_n790), .ZN(new_n791));
  OR3_X1    g590(.A1(new_n700), .A2(G85gat), .A3(new_n676), .ZN(new_n792));
  OAI21_X1  g591(.A(new_n774), .B1(new_n791), .B2(new_n792), .ZN(G1336gat));
  NOR3_X1   g592(.A1(new_n756), .A2(G92gat), .A3(new_n679), .ZN(new_n794));
  OAI21_X1  g593(.A(KEYINPUT119), .B1(new_n784), .B2(KEYINPUT51), .ZN(new_n795));
  INV_X1    g594(.A(KEYINPUT119), .ZN(new_n796));
  NAND3_X1  g595(.A1(new_n790), .A2(new_n796), .A3(new_n789), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n795), .A2(new_n797), .ZN(new_n798));
  OAI21_X1  g597(.A(new_n794), .B1(new_n788), .B2(new_n798), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n799), .A2(KEYINPUT120), .ZN(new_n800));
  NAND3_X1  g599(.A1(new_n724), .A2(new_n388), .A3(new_n772), .ZN(new_n801));
  NAND3_X1  g600(.A1(new_n801), .A2(KEYINPUT118), .A3(new_n587), .ZN(new_n802));
  INV_X1    g601(.A(KEYINPUT120), .ZN(new_n803));
  OAI211_X1 g602(.A(new_n803), .B(new_n794), .C1(new_n788), .C2(new_n798), .ZN(new_n804));
  NAND3_X1  g603(.A1(new_n800), .A2(new_n802), .A3(new_n804), .ZN(new_n805));
  AOI21_X1  g604(.A(KEYINPUT118), .B1(new_n801), .B2(new_n587), .ZN(new_n806));
  OAI21_X1  g605(.A(KEYINPUT52), .B1(new_n805), .B2(new_n806), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n801), .A2(new_n587), .ZN(new_n808));
  INV_X1    g607(.A(KEYINPUT52), .ZN(new_n809));
  INV_X1    g608(.A(new_n794), .ZN(new_n810));
  OAI211_X1 g609(.A(new_n808), .B(new_n809), .C1(new_n791), .C2(new_n810), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n807), .A2(new_n811), .ZN(new_n812));
  INV_X1    g611(.A(KEYINPUT121), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n812), .A2(new_n813), .ZN(new_n814));
  NAND3_X1  g613(.A1(new_n807), .A2(KEYINPUT121), .A3(new_n811), .ZN(new_n815));
  NAND2_X1  g614(.A1(new_n814), .A2(new_n815), .ZN(G1337gat));
  OAI21_X1  g615(.A(G99gat), .B1(new_n773), .B2(new_n692), .ZN(new_n817));
  OR3_X1    g616(.A1(new_n700), .A2(G99gat), .A3(new_n694), .ZN(new_n818));
  OAI21_X1  g617(.A(new_n817), .B1(new_n791), .B2(new_n818), .ZN(G1338gat));
  NAND3_X1  g618(.A1(new_n724), .A2(new_n752), .A3(new_n772), .ZN(new_n820));
  AND2_X1   g619(.A1(new_n820), .A2(G106gat), .ZN(new_n821));
  OR2_X1    g620(.A1(new_n788), .A2(new_n798), .ZN(new_n822));
  NOR3_X1   g621(.A1(new_n756), .A2(G106gat), .A3(new_n505), .ZN(new_n823));
  AOI21_X1  g622(.A(new_n821), .B1(new_n822), .B2(new_n823), .ZN(new_n824));
  INV_X1    g623(.A(KEYINPUT53), .ZN(new_n825));
  INV_X1    g624(.A(new_n823), .ZN(new_n826));
  OAI21_X1  g625(.A(new_n825), .B1(new_n791), .B2(new_n826), .ZN(new_n827));
  OAI22_X1  g626(.A1(new_n824), .A2(new_n825), .B1(new_n821), .B2(new_n827), .ZN(G1339gat));
  NAND3_X1  g627(.A1(new_n659), .A2(new_n660), .A3(new_n655), .ZN(new_n829));
  NAND3_X1  g628(.A1(new_n662), .A2(KEYINPUT54), .A3(new_n829), .ZN(new_n830));
  INV_X1    g629(.A(KEYINPUT54), .ZN(new_n831));
  AOI21_X1  g630(.A(new_n671), .B1(new_n661), .B2(new_n831), .ZN(new_n832));
  NAND3_X1  g631(.A1(new_n830), .A2(KEYINPUT55), .A3(new_n832), .ZN(new_n833));
  NAND2_X1  g632(.A1(new_n833), .A2(new_n672), .ZN(new_n834));
  AOI21_X1  g633(.A(KEYINPUT55), .B1(new_n830), .B2(new_n832), .ZN(new_n835));
  NOR2_X1   g634(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  NOR2_X1   g635(.A1(new_n551), .A2(new_n553), .ZN(new_n837));
  AOI21_X1  g636(.A(new_n552), .B1(new_n550), .B2(new_n558), .ZN(new_n838));
  OAI21_X1  g637(.A(new_n567), .B1(new_n837), .B2(new_n838), .ZN(new_n839));
  NAND3_X1  g638(.A1(new_n836), .A2(new_n572), .A3(new_n839), .ZN(new_n840));
  AOI21_X1  g639(.A(new_n840), .B1(new_n718), .B2(new_n720), .ZN(new_n841));
  NAND2_X1  g640(.A1(new_n718), .A2(new_n720), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n836), .A2(new_n573), .ZN(new_n843));
  NAND3_X1  g642(.A1(new_n673), .A2(new_n572), .A3(new_n839), .ZN(new_n844));
  AOI21_X1  g643(.A(new_n842), .B1(new_n843), .B2(new_n844), .ZN(new_n845));
  OAI21_X1  g644(.A(new_n701), .B1(new_n841), .B2(new_n845), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n674), .A2(new_n726), .ZN(new_n847));
  AOI21_X1  g646(.A(new_n510), .B1(new_n846), .B2(new_n847), .ZN(new_n848));
  NOR2_X1   g647(.A1(new_n676), .A2(new_n388), .ZN(new_n849));
  NAND2_X1  g648(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  NOR3_X1   g649(.A1(new_n850), .A2(new_n217), .A3(new_n577), .ZN(new_n851));
  INV_X1    g650(.A(new_n850), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n852), .A2(new_n573), .ZN(new_n853));
  AOI21_X1  g652(.A(new_n851), .B1(new_n217), .B2(new_n853), .ZN(G1340gat));
  NOR3_X1   g653(.A1(new_n850), .A2(new_n215), .A3(new_n756), .ZN(new_n855));
  NAND2_X1  g654(.A1(new_n852), .A2(new_n673), .ZN(new_n856));
  AOI21_X1  g655(.A(new_n855), .B1(new_n215), .B2(new_n856), .ZN(G1341gat));
  NOR2_X1   g656(.A1(new_n850), .A2(new_n701), .ZN(new_n858));
  XNOR2_X1  g657(.A(new_n858), .B(new_n222), .ZN(G1342gat));
  NAND4_X1  g658(.A1(new_n848), .A2(new_n207), .A3(new_n617), .A4(new_n849), .ZN(new_n860));
  XOR2_X1   g659(.A(new_n860), .B(KEYINPUT56), .Z(new_n861));
  OAI21_X1  g660(.A(G134gat), .B1(new_n850), .B2(new_n618), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n861), .A2(new_n862), .ZN(G1343gat));
  NAND2_X1  g662(.A1(new_n737), .A2(new_n849), .ZN(new_n864));
  AOI21_X1  g663(.A(new_n505), .B1(new_n846), .B2(new_n847), .ZN(new_n865));
  NOR2_X1   g664(.A1(new_n865), .A2(KEYINPUT57), .ZN(new_n866));
  INV_X1    g665(.A(new_n866), .ZN(new_n867));
  INV_X1    g666(.A(KEYINPUT57), .ZN(new_n868));
  NOR2_X1   g667(.A1(new_n505), .A2(new_n868), .ZN(new_n869));
  INV_X1    g668(.A(new_n869), .ZN(new_n870));
  NAND3_X1  g669(.A1(new_n574), .A2(new_n836), .A3(new_n576), .ZN(new_n871));
  AOI21_X1  g670(.A(new_n617), .B1(new_n871), .B2(new_n844), .ZN(new_n872));
  OAI21_X1  g671(.A(new_n701), .B1(new_n841), .B2(new_n872), .ZN(new_n873));
  AOI21_X1  g672(.A(new_n870), .B1(new_n873), .B2(new_n847), .ZN(new_n874));
  INV_X1    g673(.A(new_n874), .ZN(new_n875));
  AOI21_X1  g674(.A(new_n864), .B1(new_n867), .B2(new_n875), .ZN(new_n876));
  INV_X1    g675(.A(new_n577), .ZN(new_n877));
  AND2_X1   g676(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  INV_X1    g677(.A(G141gat), .ZN(new_n879));
  NOR2_X1   g678(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n865), .A2(new_n692), .ZN(new_n881));
  INV_X1    g680(.A(new_n881), .ZN(new_n882));
  NAND4_X1  g681(.A1(new_n882), .A2(new_n879), .A3(new_n877), .A4(new_n849), .ZN(new_n883));
  INV_X1    g682(.A(KEYINPUT58), .ZN(new_n884));
  NAND2_X1  g683(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  INV_X1    g684(.A(new_n864), .ZN(new_n886));
  OAI211_X1 g685(.A(new_n573), .B(new_n886), .C1(new_n866), .C2(new_n874), .ZN(new_n887));
  NAND2_X1  g686(.A1(new_n887), .A2(G141gat), .ZN(new_n888));
  AND3_X1   g687(.A1(new_n888), .A2(KEYINPUT122), .A3(new_n883), .ZN(new_n889));
  OAI21_X1  g688(.A(KEYINPUT58), .B1(new_n888), .B2(KEYINPUT122), .ZN(new_n890));
  OAI22_X1  g689(.A1(new_n880), .A2(new_n885), .B1(new_n889), .B2(new_n890), .ZN(G1344gat));
  NOR2_X1   g690(.A1(new_n840), .A2(new_n618), .ZN(new_n892));
  OAI21_X1  g691(.A(new_n701), .B1(new_n872), .B2(new_n892), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n674), .A2(new_n577), .ZN(new_n894));
  NAND2_X1  g693(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  AOI21_X1  g694(.A(KEYINPUT57), .B1(new_n895), .B2(new_n752), .ZN(new_n896));
  AOI21_X1  g695(.A(new_n870), .B1(new_n846), .B2(new_n847), .ZN(new_n897));
  OR2_X1    g696(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  NAND3_X1  g697(.A1(new_n898), .A2(new_n673), .A3(new_n886), .ZN(new_n899));
  NAND3_X1  g698(.A1(new_n899), .A2(KEYINPUT59), .A3(G148gat), .ZN(new_n900));
  INV_X1    g699(.A(KEYINPUT59), .ZN(new_n901));
  NAND3_X1  g700(.A1(new_n876), .A2(new_n901), .A3(new_n673), .ZN(new_n902));
  NOR3_X1   g701(.A1(new_n881), .A2(new_n676), .A3(new_n388), .ZN(new_n903));
  AOI21_X1  g702(.A(new_n901), .B1(new_n903), .B2(new_n673), .ZN(new_n904));
  OAI211_X1 g703(.A(new_n900), .B(new_n902), .C1(G148gat), .C2(new_n904), .ZN(G1345gat));
  INV_X1    g704(.A(G155gat), .ZN(new_n906));
  NAND3_X1  g705(.A1(new_n903), .A2(new_n906), .A3(new_n652), .ZN(new_n907));
  AND2_X1   g706(.A1(new_n876), .A2(new_n652), .ZN(new_n908));
  OAI21_X1  g707(.A(new_n907), .B1(new_n908), .B2(new_n906), .ZN(G1346gat));
  INV_X1    g708(.A(G162gat), .ZN(new_n910));
  NAND4_X1  g709(.A1(new_n882), .A2(new_n910), .A3(new_n617), .A4(new_n849), .ZN(new_n911));
  AND2_X1   g710(.A1(new_n876), .A2(new_n842), .ZN(new_n912));
  OAI21_X1  g711(.A(new_n911), .B1(new_n912), .B2(new_n910), .ZN(G1347gat));
  NOR2_X1   g712(.A1(new_n679), .A2(new_n430), .ZN(new_n914));
  NAND2_X1  g713(.A1(new_n848), .A2(new_n914), .ZN(new_n915));
  INV_X1    g714(.A(G169gat), .ZN(new_n916));
  NOR3_X1   g715(.A1(new_n915), .A2(new_n916), .A3(new_n577), .ZN(new_n917));
  INV_X1    g716(.A(new_n915), .ZN(new_n918));
  NAND2_X1  g717(.A1(new_n918), .A2(new_n573), .ZN(new_n919));
  AOI21_X1  g718(.A(new_n917), .B1(new_n916), .B2(new_n919), .ZN(G1348gat));
  OAI21_X1  g719(.A(G176gat), .B1(new_n915), .B2(new_n756), .ZN(new_n921));
  OR2_X1    g720(.A1(new_n700), .A2(G176gat), .ZN(new_n922));
  OAI21_X1  g721(.A(new_n921), .B1(new_n915), .B2(new_n922), .ZN(G1349gat));
  OAI21_X1  g722(.A(new_n340), .B1(new_n915), .B2(new_n701), .ZN(new_n924));
  INV_X1    g723(.A(KEYINPUT60), .ZN(new_n925));
  NAND2_X1  g724(.A1(new_n925), .A2(KEYINPUT123), .ZN(new_n926));
  NAND2_X1  g725(.A1(new_n918), .A2(new_n652), .ZN(new_n927));
  OAI211_X1 g726(.A(new_n924), .B(new_n926), .C1(new_n927), .C2(new_n354), .ZN(new_n928));
  NOR2_X1   g727(.A1(new_n925), .A2(KEYINPUT123), .ZN(new_n929));
  XOR2_X1   g728(.A(new_n928), .B(new_n929), .Z(G1350gat));
  OAI21_X1  g729(.A(G190gat), .B1(new_n915), .B2(new_n618), .ZN(new_n931));
  XNOR2_X1  g730(.A(new_n931), .B(KEYINPUT61), .ZN(new_n932));
  NAND3_X1  g731(.A1(new_n918), .A2(new_n325), .A3(new_n842), .ZN(new_n933));
  NAND2_X1  g732(.A1(new_n932), .A2(new_n933), .ZN(G1351gat));
  AND2_X1   g733(.A1(new_n692), .A2(new_n914), .ZN(new_n935));
  NAND2_X1  g734(.A1(new_n898), .A2(new_n935), .ZN(new_n936));
  NOR3_X1   g735(.A1(new_n936), .A2(new_n289), .A3(new_n577), .ZN(new_n937));
  AND2_X1   g736(.A1(new_n865), .A2(new_n935), .ZN(new_n938));
  AOI21_X1  g737(.A(G197gat), .B1(new_n938), .B2(new_n573), .ZN(new_n939));
  NOR2_X1   g738(.A1(new_n937), .A2(new_n939), .ZN(G1352gat));
  NAND3_X1  g739(.A1(new_n938), .A2(new_n302), .A3(new_n673), .ZN(new_n941));
  AOI21_X1  g740(.A(new_n941), .B1(KEYINPUT124), .B2(KEYINPUT62), .ZN(new_n942));
  XNOR2_X1  g741(.A(KEYINPUT124), .B(KEYINPUT62), .ZN(new_n943));
  AOI21_X1  g742(.A(new_n942), .B1(new_n941), .B2(new_n943), .ZN(new_n944));
  OAI21_X1  g743(.A(G204gat), .B1(new_n936), .B2(new_n756), .ZN(new_n945));
  NAND2_X1  g744(.A1(new_n944), .A2(new_n945), .ZN(G1353gat));
  INV_X1    g745(.A(G211gat), .ZN(new_n947));
  NAND3_X1  g746(.A1(new_n938), .A2(new_n947), .A3(new_n652), .ZN(new_n948));
  OAI211_X1 g747(.A(new_n652), .B(new_n935), .C1(new_n896), .C2(new_n897), .ZN(new_n949));
  INV_X1    g748(.A(KEYINPUT63), .ZN(new_n950));
  NOR2_X1   g749(.A1(new_n950), .A2(KEYINPUT125), .ZN(new_n951));
  AOI21_X1  g750(.A(new_n947), .B1(KEYINPUT125), .B2(new_n950), .ZN(new_n952));
  AND3_X1   g751(.A1(new_n949), .A2(new_n951), .A3(new_n952), .ZN(new_n953));
  AOI21_X1  g752(.A(new_n951), .B1(new_n949), .B2(new_n952), .ZN(new_n954));
  OAI21_X1  g753(.A(new_n948), .B1(new_n953), .B2(new_n954), .ZN(new_n955));
  INV_X1    g754(.A(KEYINPUT126), .ZN(new_n956));
  NAND2_X1  g755(.A1(new_n955), .A2(new_n956), .ZN(new_n957));
  OAI211_X1 g756(.A(KEYINPUT126), .B(new_n948), .C1(new_n953), .C2(new_n954), .ZN(new_n958));
  NAND2_X1  g757(.A1(new_n957), .A2(new_n958), .ZN(G1354gat));
  INV_X1    g758(.A(G218gat), .ZN(new_n960));
  NAND3_X1  g759(.A1(new_n938), .A2(new_n960), .A3(new_n842), .ZN(new_n961));
  NAND2_X1  g760(.A1(new_n936), .A2(KEYINPUT127), .ZN(new_n962));
  INV_X1    g761(.A(KEYINPUT127), .ZN(new_n963));
  NAND3_X1  g762(.A1(new_n898), .A2(new_n963), .A3(new_n935), .ZN(new_n964));
  AND3_X1   g763(.A1(new_n962), .A2(new_n617), .A3(new_n964), .ZN(new_n965));
  OAI21_X1  g764(.A(new_n961), .B1(new_n965), .B2(new_n960), .ZN(G1355gat));
endmodule


