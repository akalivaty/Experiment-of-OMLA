//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 1 1 1 1 1 1 0 1 1 1 0 1 1 1 0 1 1 0 1 1 0 0 0 0 0 1 1 0 0 0 1 0 0 1 1 1 0 0 0 0 0 0 0 1 0 1 0 1 0 0 0 1 1 1 1 1 0 1 1 0 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:30:25 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n443, new_n448, new_n449, new_n453, new_n454, new_n455,
    new_n456, new_n457, new_n460, new_n461, new_n462, new_n463, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n529, new_n530, new_n531, new_n532,
    new_n533, new_n534, new_n535, new_n536, new_n537, new_n539, new_n540,
    new_n541, new_n542, new_n543, new_n544, new_n545, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n554, new_n556, new_n557,
    new_n558, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n570, new_n571, new_n572, new_n574, new_n575, new_n576,
    new_n578, new_n579, new_n580, new_n581, new_n582, new_n583, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n606, new_n607, new_n610, new_n611,
    new_n613, new_n614, new_n615, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1171, new_n1172,
    new_n1173, new_n1174, new_n1175, new_n1176, new_n1177, new_n1178,
    new_n1179, new_n1181;
  BUF_X1    g000(.A(G452), .Z(G350));
  XNOR2_X1  g001(.A(KEYINPUT64), .B(G452), .ZN(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(new_n436));
  XNOR2_X1  g011(.A(new_n436), .B(KEYINPUT65), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  XOR2_X1   g013(.A(KEYINPUT66), .B(G69), .Z(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  XOR2_X1   g016(.A(KEYINPUT67), .B(G108), .Z(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(new_n443));
  XNOR2_X1  g018(.A(new_n443), .B(KEYINPUT68), .ZN(G158));
  NAND3_X1  g019(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g020(.A(G452), .Z(G391));
  AND2_X1   g021(.A1(G94), .A2(G452), .ZN(G173));
  XNOR2_X1  g022(.A(KEYINPUT69), .B(KEYINPUT1), .ZN(new_n448));
  AND2_X1   g023(.A1(G7), .A2(G661), .ZN(new_n449));
  XNOR2_X1  g024(.A(new_n448), .B(new_n449), .ZN(G223));
  NAND2_X1  g025(.A1(new_n449), .A2(G567), .ZN(G234));
  NAND2_X1  g026(.A1(new_n449), .A2(G2106), .ZN(G217));
  OR4_X1    g027(.A1(G218), .A2(G220), .A3(G221), .A4(G219), .ZN(new_n453));
  XNOR2_X1  g028(.A(new_n453), .B(KEYINPUT2), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR4_X1   g030(.A1(G238), .A2(G235), .A3(G237), .A4(G236), .ZN(new_n456));
  NAND2_X1  g031(.A1(new_n455), .A2(new_n456), .ZN(new_n457));
  XNOR2_X1  g032(.A(new_n457), .B(KEYINPUT70), .ZN(G261));
  INV_X1    g033(.A(G261), .ZN(G325));
  NAND2_X1  g034(.A1(new_n454), .A2(G2106), .ZN(new_n460));
  INV_X1    g035(.A(G567), .ZN(new_n461));
  OR2_X1    g036(.A1(new_n456), .A2(new_n461), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n460), .A2(new_n462), .ZN(new_n463));
  INV_X1    g038(.A(new_n463), .ZN(G319));
  INV_X1    g039(.A(G2105), .ZN(new_n465));
  INV_X1    g040(.A(KEYINPUT3), .ZN(new_n466));
  INV_X1    g041(.A(G2104), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  NAND2_X1  g043(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n470), .A2(G125), .ZN(new_n471));
  NAND2_X1  g046(.A1(G113), .A2(G2104), .ZN(new_n472));
  AOI21_X1  g047(.A(new_n465), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  NAND3_X1  g048(.A1(new_n470), .A2(G137), .A3(new_n465), .ZN(new_n474));
  NOR2_X1   g049(.A1(new_n467), .A2(G2105), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n475), .A2(G101), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n474), .A2(new_n476), .ZN(new_n477));
  NOR2_X1   g052(.A1(new_n473), .A2(new_n477), .ZN(G160));
  NAND2_X1  g053(.A1(new_n470), .A2(new_n465), .ZN(new_n479));
  INV_X1    g054(.A(new_n479), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n480), .A2(G136), .ZN(new_n481));
  NOR2_X1   g056(.A1(G100), .A2(G2105), .ZN(new_n482));
  XOR2_X1   g057(.A(new_n482), .B(KEYINPUT72), .Z(new_n483));
  OAI21_X1  g058(.A(G2104), .B1(new_n465), .B2(G112), .ZN(new_n484));
  OAI21_X1  g059(.A(new_n481), .B1(new_n483), .B2(new_n484), .ZN(new_n485));
  NAND3_X1  g060(.A1(new_n470), .A2(KEYINPUT71), .A3(G2105), .ZN(new_n486));
  INV_X1    g061(.A(new_n486), .ZN(new_n487));
  AOI21_X1  g062(.A(KEYINPUT71), .B1(new_n470), .B2(G2105), .ZN(new_n488));
  NOR2_X1   g063(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  INV_X1    g064(.A(new_n489), .ZN(new_n490));
  AOI21_X1  g065(.A(new_n485), .B1(G124), .B2(new_n490), .ZN(new_n491));
  XNOR2_X1  g066(.A(new_n491), .B(KEYINPUT73), .ZN(G162));
  INV_X1    g067(.A(G126), .ZN(new_n493));
  AOI21_X1  g068(.A(new_n493), .B1(new_n468), .B2(new_n469), .ZN(new_n494));
  AND2_X1   g069(.A1(G114), .A2(G2104), .ZN(new_n495));
  OAI21_X1  g070(.A(G2105), .B1(new_n494), .B2(new_n495), .ZN(new_n496));
  NAND2_X1  g071(.A1(KEYINPUT4), .A2(G138), .ZN(new_n497));
  AOI21_X1  g072(.A(new_n497), .B1(new_n468), .B2(new_n469), .ZN(new_n498));
  NAND2_X1  g073(.A1(G102), .A2(G2104), .ZN(new_n499));
  INV_X1    g074(.A(new_n499), .ZN(new_n500));
  OAI21_X1  g075(.A(new_n465), .B1(new_n498), .B2(new_n500), .ZN(new_n501));
  AND2_X1   g076(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n502));
  NOR2_X1   g077(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n503));
  OAI211_X1 g078(.A(G138), .B(new_n465), .C1(new_n502), .C2(new_n503), .ZN(new_n504));
  INV_X1    g079(.A(KEYINPUT4), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  NAND3_X1  g081(.A1(new_n496), .A2(new_n501), .A3(new_n506), .ZN(new_n507));
  INV_X1    g082(.A(new_n507), .ZN(G164));
  INV_X1    g083(.A(G62), .ZN(new_n509));
  OR2_X1    g084(.A1(KEYINPUT5), .A2(G543), .ZN(new_n510));
  NAND2_X1  g085(.A1(KEYINPUT5), .A2(G543), .ZN(new_n511));
  AOI21_X1  g086(.A(new_n509), .B1(new_n510), .B2(new_n511), .ZN(new_n512));
  NAND2_X1  g087(.A1(G75), .A2(G543), .ZN(new_n513));
  INV_X1    g088(.A(new_n513), .ZN(new_n514));
  OAI21_X1  g089(.A(G651), .B1(new_n512), .B2(new_n514), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n510), .A2(new_n511), .ZN(new_n516));
  OR2_X1    g091(.A1(KEYINPUT6), .A2(G651), .ZN(new_n517));
  NAND2_X1  g092(.A1(KEYINPUT6), .A2(G651), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  NAND3_X1  g094(.A1(new_n516), .A2(new_n519), .A3(G88), .ZN(new_n520));
  INV_X1    g095(.A(G543), .ZN(new_n521));
  AOI21_X1  g096(.A(new_n521), .B1(new_n517), .B2(new_n518), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n522), .A2(G50), .ZN(new_n523));
  NAND3_X1  g098(.A1(new_n515), .A2(new_n520), .A3(new_n523), .ZN(new_n524));
  INV_X1    g099(.A(KEYINPUT74), .ZN(new_n525));
  NAND2_X1  g100(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  NAND4_X1  g101(.A1(new_n515), .A2(KEYINPUT74), .A3(new_n520), .A4(new_n523), .ZN(new_n527));
  NAND2_X1  g102(.A1(new_n526), .A2(new_n527), .ZN(G166));
  INV_X1    g103(.A(new_n516), .ZN(new_n529));
  NAND2_X1  g104(.A1(new_n519), .A2(G89), .ZN(new_n530));
  NAND2_X1  g105(.A1(G63), .A2(G651), .ZN(new_n531));
  AOI21_X1  g106(.A(new_n529), .B1(new_n530), .B2(new_n531), .ZN(new_n532));
  NAND3_X1  g107(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n533));
  XNOR2_X1  g108(.A(new_n533), .B(KEYINPUT7), .ZN(new_n534));
  NAND2_X1  g109(.A1(new_n519), .A2(G543), .ZN(new_n535));
  INV_X1    g110(.A(G51), .ZN(new_n536));
  OAI21_X1  g111(.A(new_n534), .B1(new_n535), .B2(new_n536), .ZN(new_n537));
  NOR2_X1   g112(.A1(new_n532), .A2(new_n537), .ZN(G168));
  NAND2_X1  g113(.A1(new_n522), .A2(G52), .ZN(new_n539));
  INV_X1    g114(.A(G90), .ZN(new_n540));
  NAND2_X1  g115(.A1(new_n516), .A2(new_n519), .ZN(new_n541));
  OAI21_X1  g116(.A(new_n539), .B1(new_n540), .B2(new_n541), .ZN(new_n542));
  AOI22_X1  g117(.A1(new_n516), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n543));
  INV_X1    g118(.A(G651), .ZN(new_n544));
  NOR2_X1   g119(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  NOR2_X1   g120(.A1(new_n542), .A2(new_n545), .ZN(G171));
  NAND2_X1  g121(.A1(new_n522), .A2(G43), .ZN(new_n547));
  INV_X1    g122(.A(G81), .ZN(new_n548));
  OAI21_X1  g123(.A(new_n547), .B1(new_n548), .B2(new_n541), .ZN(new_n549));
  AOI22_X1  g124(.A1(new_n516), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n550));
  NOR2_X1   g125(.A1(new_n550), .A2(new_n544), .ZN(new_n551));
  NOR2_X1   g126(.A1(new_n549), .A2(new_n551), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n552), .A2(G860), .ZN(G153));
  AND3_X1   g128(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n554), .A2(G36), .ZN(G176));
  NAND2_X1  g130(.A1(G1), .A2(G3), .ZN(new_n556));
  XNOR2_X1  g131(.A(new_n556), .B(KEYINPUT75), .ZN(new_n557));
  XNOR2_X1  g132(.A(new_n557), .B(KEYINPUT8), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n554), .A2(new_n558), .ZN(G188));
  NAND2_X1  g134(.A1(new_n522), .A2(G53), .ZN(new_n560));
  XNOR2_X1  g135(.A(new_n560), .B(KEYINPUT9), .ZN(new_n561));
  INV_X1    g136(.A(G91), .ZN(new_n562));
  OR3_X1    g137(.A1(new_n541), .A2(KEYINPUT76), .A3(new_n562), .ZN(new_n563));
  AOI22_X1  g138(.A1(new_n516), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n564));
  OR2_X1    g139(.A1(new_n564), .A2(new_n544), .ZN(new_n565));
  OAI21_X1  g140(.A(KEYINPUT76), .B1(new_n541), .B2(new_n562), .ZN(new_n566));
  NAND4_X1  g141(.A1(new_n561), .A2(new_n563), .A3(new_n565), .A4(new_n566), .ZN(G299));
  XOR2_X1   g142(.A(G171), .B(KEYINPUT77), .Z(G301));
  INV_X1    g143(.A(G168), .ZN(G286));
  INV_X1    g144(.A(KEYINPUT78), .ZN(new_n570));
  AND3_X1   g145(.A1(new_n526), .A2(new_n570), .A3(new_n527), .ZN(new_n571));
  AOI21_X1  g146(.A(new_n570), .B1(new_n526), .B2(new_n527), .ZN(new_n572));
  NOR2_X1   g147(.A1(new_n571), .A2(new_n572), .ZN(G303));
  OAI21_X1  g148(.A(G651), .B1(new_n516), .B2(G74), .ZN(new_n574));
  NAND2_X1  g149(.A1(new_n522), .A2(G49), .ZN(new_n575));
  NAND3_X1  g150(.A1(new_n516), .A2(new_n519), .A3(G87), .ZN(new_n576));
  NAND3_X1  g151(.A1(new_n574), .A2(new_n575), .A3(new_n576), .ZN(G288));
  NAND2_X1  g152(.A1(new_n522), .A2(G48), .ZN(new_n578));
  INV_X1    g153(.A(G86), .ZN(new_n579));
  OAI21_X1  g154(.A(new_n578), .B1(new_n579), .B2(new_n541), .ZN(new_n580));
  AOI22_X1  g155(.A1(new_n516), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n581));
  NOR2_X1   g156(.A1(new_n581), .A2(new_n544), .ZN(new_n582));
  NOR2_X1   g157(.A1(new_n580), .A2(new_n582), .ZN(new_n583));
  INV_X1    g158(.A(new_n583), .ZN(G305));
  NAND2_X1  g159(.A1(new_n522), .A2(G47), .ZN(new_n585));
  INV_X1    g160(.A(G85), .ZN(new_n586));
  OAI21_X1  g161(.A(new_n585), .B1(new_n586), .B2(new_n541), .ZN(new_n587));
  AOI22_X1  g162(.A1(new_n516), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n588));
  NOR2_X1   g163(.A1(new_n588), .A2(new_n544), .ZN(new_n589));
  OR3_X1    g164(.A1(new_n587), .A2(new_n589), .A3(KEYINPUT79), .ZN(new_n590));
  OAI21_X1  g165(.A(KEYINPUT79), .B1(new_n587), .B2(new_n589), .ZN(new_n591));
  NAND2_X1  g166(.A1(new_n590), .A2(new_n591), .ZN(G290));
  NAND3_X1  g167(.A1(new_n516), .A2(new_n519), .A3(G92), .ZN(new_n593));
  XOR2_X1   g168(.A(new_n593), .B(KEYINPUT10), .Z(new_n594));
  NAND2_X1  g169(.A1(G79), .A2(G543), .ZN(new_n595));
  INV_X1    g170(.A(G66), .ZN(new_n596));
  OAI21_X1  g171(.A(new_n595), .B1(new_n529), .B2(new_n596), .ZN(new_n597));
  AOI22_X1  g172(.A1(new_n597), .A2(G651), .B1(G54), .B2(new_n522), .ZN(new_n598));
  AND2_X1   g173(.A1(new_n594), .A2(new_n598), .ZN(new_n599));
  INV_X1    g174(.A(new_n599), .ZN(new_n600));
  INV_X1    g175(.A(G868), .ZN(new_n601));
  NAND2_X1  g176(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  XNOR2_X1  g177(.A(G171), .B(KEYINPUT77), .ZN(new_n603));
  OAI21_X1  g178(.A(new_n602), .B1(new_n603), .B2(new_n601), .ZN(G284));
  XOR2_X1   g179(.A(G284), .B(KEYINPUT80), .Z(G321));
  NOR2_X1   g180(.A1(G286), .A2(new_n601), .ZN(new_n606));
  INV_X1    g181(.A(G299), .ZN(new_n607));
  AOI21_X1  g182(.A(new_n606), .B1(new_n607), .B2(new_n601), .ZN(G297));
  AOI21_X1  g183(.A(new_n606), .B1(new_n607), .B2(new_n601), .ZN(G280));
  INV_X1    g184(.A(G559), .ZN(new_n610));
  OAI21_X1  g185(.A(new_n599), .B1(new_n610), .B2(G860), .ZN(new_n611));
  XNOR2_X1  g186(.A(new_n611), .B(KEYINPUT81), .ZN(G148));
  NAND3_X1  g187(.A1(new_n599), .A2(new_n610), .A3(G868), .ZN(new_n613));
  NAND2_X1  g188(.A1(new_n552), .A2(new_n601), .ZN(new_n614));
  NAND2_X1  g189(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  XOR2_X1   g190(.A(new_n615), .B(KEYINPUT11), .Z(G282));
  INV_X1    g191(.A(new_n615), .ZN(G323));
  NOR2_X1   g192(.A1(new_n479), .A2(new_n467), .ZN(new_n618));
  XOR2_X1   g193(.A(KEYINPUT82), .B(KEYINPUT12), .Z(new_n619));
  XNOR2_X1  g194(.A(new_n618), .B(new_n619), .ZN(new_n620));
  XNOR2_X1  g195(.A(KEYINPUT13), .B(G2100), .ZN(new_n621));
  XNOR2_X1  g196(.A(new_n620), .B(new_n621), .ZN(new_n622));
  NAND2_X1  g197(.A1(new_n490), .A2(G123), .ZN(new_n623));
  INV_X1    g198(.A(G2096), .ZN(new_n624));
  MUX2_X1   g199(.A(G99), .B(G111), .S(G2105), .Z(new_n625));
  AOI22_X1  g200(.A1(new_n480), .A2(G135), .B1(G2104), .B2(new_n625), .ZN(new_n626));
  NAND3_X1  g201(.A1(new_n623), .A2(new_n624), .A3(new_n626), .ZN(new_n627));
  NAND2_X1  g202(.A1(new_n623), .A2(new_n626), .ZN(new_n628));
  NAND2_X1  g203(.A1(new_n628), .A2(G2096), .ZN(new_n629));
  NAND3_X1  g204(.A1(new_n622), .A2(new_n627), .A3(new_n629), .ZN(G156));
  INV_X1    g205(.A(KEYINPUT14), .ZN(new_n631));
  XNOR2_X1  g206(.A(KEYINPUT15), .B(G2435), .ZN(new_n632));
  XNOR2_X1  g207(.A(new_n632), .B(G2438), .ZN(new_n633));
  XNOR2_X1  g208(.A(G2427), .B(G2430), .ZN(new_n634));
  AOI21_X1  g209(.A(new_n631), .B1(new_n633), .B2(new_n634), .ZN(new_n635));
  XNOR2_X1  g210(.A(new_n635), .B(KEYINPUT84), .ZN(new_n636));
  OAI21_X1  g211(.A(new_n636), .B1(new_n633), .B2(new_n634), .ZN(new_n637));
  XOR2_X1   g212(.A(KEYINPUT83), .B(KEYINPUT16), .Z(new_n638));
  XNOR2_X1  g213(.A(new_n637), .B(new_n638), .ZN(new_n639));
  XNOR2_X1  g214(.A(G1341), .B(G1348), .ZN(new_n640));
  XNOR2_X1  g215(.A(new_n639), .B(new_n640), .ZN(new_n641));
  XNOR2_X1  g216(.A(G2451), .B(G2454), .ZN(new_n642));
  XNOR2_X1  g217(.A(G2443), .B(G2446), .ZN(new_n643));
  XOR2_X1   g218(.A(new_n642), .B(new_n643), .Z(new_n644));
  INV_X1    g219(.A(new_n644), .ZN(new_n645));
  NAND2_X1  g220(.A1(new_n641), .A2(new_n645), .ZN(new_n646));
  NAND2_X1  g221(.A1(new_n646), .A2(G14), .ZN(new_n647));
  NOR2_X1   g222(.A1(new_n641), .A2(new_n645), .ZN(new_n648));
  NOR2_X1   g223(.A1(new_n647), .A2(new_n648), .ZN(G401));
  XNOR2_X1  g224(.A(G2072), .B(G2078), .ZN(new_n650));
  XOR2_X1   g225(.A(new_n650), .B(KEYINPUT17), .Z(new_n651));
  XNOR2_X1  g226(.A(G2067), .B(G2678), .ZN(new_n652));
  INV_X1    g227(.A(new_n652), .ZN(new_n653));
  XNOR2_X1  g228(.A(G2084), .B(G2090), .ZN(new_n654));
  INV_X1    g229(.A(new_n654), .ZN(new_n655));
  NAND3_X1  g230(.A1(new_n651), .A2(new_n653), .A3(new_n655), .ZN(new_n656));
  INV_X1    g231(.A(KEYINPUT86), .ZN(new_n657));
  XNOR2_X1  g232(.A(new_n656), .B(new_n657), .ZN(new_n658));
  XOR2_X1   g233(.A(new_n650), .B(KEYINPUT85), .Z(new_n659));
  NAND2_X1  g234(.A1(new_n659), .A2(new_n653), .ZN(new_n660));
  OAI211_X1 g235(.A(new_n660), .B(new_n654), .C1(new_n651), .C2(new_n653), .ZN(new_n661));
  NAND3_X1  g236(.A1(new_n655), .A2(new_n650), .A3(new_n652), .ZN(new_n662));
  XOR2_X1   g237(.A(new_n662), .B(KEYINPUT18), .Z(new_n663));
  NAND3_X1  g238(.A1(new_n658), .A2(new_n661), .A3(new_n663), .ZN(new_n664));
  XNOR2_X1  g239(.A(new_n664), .B(new_n624), .ZN(new_n665));
  XNOR2_X1  g240(.A(new_n665), .B(G2100), .ZN(G227));
  XNOR2_X1  g241(.A(G1956), .B(G2474), .ZN(new_n667));
  XNOR2_X1  g242(.A(new_n667), .B(KEYINPUT87), .ZN(new_n668));
  XOR2_X1   g243(.A(G1961), .B(G1966), .Z(new_n669));
  NAND2_X1  g244(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  XNOR2_X1  g245(.A(new_n670), .B(KEYINPUT88), .ZN(new_n671));
  XNOR2_X1  g246(.A(G1971), .B(G1976), .ZN(new_n672));
  XNOR2_X1  g247(.A(new_n672), .B(KEYINPUT19), .ZN(new_n673));
  INV_X1    g248(.A(new_n673), .ZN(new_n674));
  NAND2_X1  g249(.A1(new_n671), .A2(new_n674), .ZN(new_n675));
  XNOR2_X1  g250(.A(new_n675), .B(KEYINPUT20), .ZN(new_n676));
  NAND2_X1  g251(.A1(new_n670), .A2(new_n673), .ZN(new_n677));
  NOR2_X1   g252(.A1(new_n668), .A2(new_n669), .ZN(new_n678));
  MUX2_X1   g253(.A(new_n677), .B(new_n673), .S(new_n678), .Z(new_n679));
  NAND2_X1  g254(.A1(new_n676), .A2(new_n679), .ZN(new_n680));
  XNOR2_X1  g255(.A(G1981), .B(G1986), .ZN(new_n681));
  INV_X1    g256(.A(new_n681), .ZN(new_n682));
  NAND2_X1  g257(.A1(new_n680), .A2(new_n682), .ZN(new_n683));
  NAND3_X1  g258(.A1(new_n676), .A2(new_n679), .A3(new_n681), .ZN(new_n684));
  XNOR2_X1  g259(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n685));
  XNOR2_X1  g260(.A(new_n685), .B(KEYINPUT89), .ZN(new_n686));
  XNOR2_X1  g261(.A(new_n686), .B(KEYINPUT90), .ZN(new_n687));
  XOR2_X1   g262(.A(G1991), .B(G1996), .Z(new_n688));
  XNOR2_X1  g263(.A(new_n687), .B(new_n688), .ZN(new_n689));
  AND3_X1   g264(.A1(new_n683), .A2(new_n684), .A3(new_n689), .ZN(new_n690));
  AOI21_X1  g265(.A(new_n689), .B1(new_n683), .B2(new_n684), .ZN(new_n691));
  OR2_X1    g266(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  INV_X1    g267(.A(new_n692), .ZN(G229));
  INV_X1    g268(.A(G16), .ZN(new_n694));
  NAND2_X1  g269(.A1(new_n694), .A2(G20), .ZN(new_n695));
  XNOR2_X1  g270(.A(new_n695), .B(KEYINPUT23), .ZN(new_n696));
  OAI21_X1  g271(.A(new_n696), .B1(new_n607), .B2(new_n694), .ZN(new_n697));
  XNOR2_X1  g272(.A(new_n697), .B(G1956), .ZN(new_n698));
  INV_X1    g273(.A(G29), .ZN(new_n699));
  NAND2_X1  g274(.A1(new_n699), .A2(G26), .ZN(new_n700));
  XNOR2_X1  g275(.A(new_n700), .B(KEYINPUT28), .ZN(new_n701));
  MUX2_X1   g276(.A(G104), .B(G116), .S(G2105), .Z(new_n702));
  NAND2_X1  g277(.A1(new_n702), .A2(G2104), .ZN(new_n703));
  XOR2_X1   g278(.A(new_n703), .B(KEYINPUT94), .Z(new_n704));
  INV_X1    g279(.A(G140), .ZN(new_n705));
  OAI21_X1  g280(.A(new_n704), .B1(new_n705), .B2(new_n479), .ZN(new_n706));
  AND2_X1   g281(.A1(new_n490), .A2(G128), .ZN(new_n707));
  NOR2_X1   g282(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  OAI21_X1  g283(.A(new_n701), .B1(new_n708), .B2(new_n699), .ZN(new_n709));
  INV_X1    g284(.A(G2067), .ZN(new_n710));
  XNOR2_X1  g285(.A(new_n709), .B(new_n710), .ZN(new_n711));
  NOR2_X1   g286(.A1(G16), .A2(G19), .ZN(new_n712));
  AOI21_X1  g287(.A(new_n712), .B1(new_n552), .B2(G16), .ZN(new_n713));
  XNOR2_X1  g288(.A(new_n713), .B(G1341), .ZN(new_n714));
  XNOR2_X1  g289(.A(KEYINPUT93), .B(G1348), .ZN(new_n715));
  INV_X1    g290(.A(new_n715), .ZN(new_n716));
  NOR2_X1   g291(.A1(G4), .A2(G16), .ZN(new_n717));
  AOI21_X1  g292(.A(new_n717), .B1(new_n599), .B2(G16), .ZN(new_n718));
  AOI21_X1  g293(.A(new_n714), .B1(new_n716), .B2(new_n718), .ZN(new_n719));
  OR2_X1    g294(.A1(new_n718), .A2(new_n716), .ZN(new_n720));
  NAND3_X1  g295(.A1(new_n711), .A2(new_n719), .A3(new_n720), .ZN(new_n721));
  NOR2_X1   g296(.A1(G29), .A2(G35), .ZN(new_n722));
  AOI21_X1  g297(.A(new_n722), .B1(G162), .B2(G29), .ZN(new_n723));
  XOR2_X1   g298(.A(KEYINPUT99), .B(KEYINPUT29), .Z(new_n724));
  XNOR2_X1  g299(.A(new_n723), .B(new_n724), .ZN(new_n725));
  INV_X1    g300(.A(G2090), .ZN(new_n726));
  AOI211_X1 g301(.A(new_n698), .B(new_n721), .C1(new_n725), .C2(new_n726), .ZN(new_n727));
  NAND2_X1  g302(.A1(new_n699), .A2(G33), .ZN(new_n728));
  INV_X1    g303(.A(new_n475), .ZN(new_n729));
  INV_X1    g304(.A(G103), .ZN(new_n730));
  OR3_X1    g305(.A1(new_n729), .A2(KEYINPUT25), .A3(new_n730), .ZN(new_n731));
  OAI21_X1  g306(.A(KEYINPUT25), .B1(new_n729), .B2(new_n730), .ZN(new_n732));
  INV_X1    g307(.A(G139), .ZN(new_n733));
  OAI211_X1 g308(.A(new_n731), .B(new_n732), .C1(new_n479), .C2(new_n733), .ZN(new_n734));
  XOR2_X1   g309(.A(new_n734), .B(KEYINPUT95), .Z(new_n735));
  AOI22_X1  g310(.A1(new_n470), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n736));
  NOR2_X1   g311(.A1(new_n736), .A2(new_n465), .ZN(new_n737));
  NOR2_X1   g312(.A1(new_n735), .A2(new_n737), .ZN(new_n738));
  OAI21_X1  g313(.A(new_n728), .B1(new_n738), .B2(new_n699), .ZN(new_n739));
  XOR2_X1   g314(.A(new_n739), .B(G2072), .Z(new_n740));
  NOR2_X1   g315(.A1(G27), .A2(G29), .ZN(new_n741));
  AOI21_X1  g316(.A(new_n741), .B1(G164), .B2(G29), .ZN(new_n742));
  XNOR2_X1  g317(.A(KEYINPUT97), .B(G2078), .ZN(new_n743));
  XNOR2_X1  g318(.A(new_n742), .B(new_n743), .ZN(new_n744));
  NAND2_X1  g319(.A1(new_n699), .A2(G32), .ZN(new_n745));
  AOI22_X1  g320(.A1(new_n480), .A2(G141), .B1(G105), .B2(new_n475), .ZN(new_n746));
  NAND3_X1  g321(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n747));
  XOR2_X1   g322(.A(new_n747), .B(KEYINPUT26), .Z(new_n748));
  NAND2_X1  g323(.A1(new_n746), .A2(new_n748), .ZN(new_n749));
  AOI21_X1  g324(.A(new_n749), .B1(G129), .B2(new_n490), .ZN(new_n750));
  OAI21_X1  g325(.A(new_n745), .B1(new_n750), .B2(new_n699), .ZN(new_n751));
  XNOR2_X1  g326(.A(KEYINPUT27), .B(G1996), .ZN(new_n752));
  XNOR2_X1  g327(.A(new_n751), .B(new_n752), .ZN(new_n753));
  OR2_X1    g328(.A1(KEYINPUT24), .A2(G34), .ZN(new_n754));
  NAND2_X1  g329(.A1(KEYINPUT24), .A2(G34), .ZN(new_n755));
  AOI21_X1  g330(.A(G29), .B1(new_n754), .B2(new_n755), .ZN(new_n756));
  AOI21_X1  g331(.A(new_n756), .B1(G160), .B2(G29), .ZN(new_n757));
  XOR2_X1   g332(.A(new_n757), .B(G2084), .Z(new_n758));
  NAND2_X1  g333(.A1(new_n694), .A2(G5), .ZN(new_n759));
  OAI21_X1  g334(.A(new_n759), .B1(G171), .B2(new_n694), .ZN(new_n760));
  OAI21_X1  g335(.A(new_n758), .B1(G1961), .B2(new_n760), .ZN(new_n761));
  NAND2_X1  g336(.A1(new_n694), .A2(G21), .ZN(new_n762));
  OAI21_X1  g337(.A(new_n762), .B1(G168), .B2(new_n694), .ZN(new_n763));
  NOR2_X1   g338(.A1(new_n763), .A2(G1966), .ZN(new_n764));
  XOR2_X1   g339(.A(KEYINPUT96), .B(G28), .Z(new_n765));
  AOI21_X1  g340(.A(G29), .B1(new_n765), .B2(KEYINPUT30), .ZN(new_n766));
  OAI21_X1  g341(.A(new_n766), .B1(KEYINPUT30), .B2(new_n765), .ZN(new_n767));
  XNOR2_X1  g342(.A(KEYINPUT31), .B(G11), .ZN(new_n768));
  OAI211_X1 g343(.A(new_n767), .B(new_n768), .C1(new_n628), .C2(new_n699), .ZN(new_n769));
  NAND2_X1  g344(.A1(new_n760), .A2(G1961), .ZN(new_n770));
  INV_X1    g345(.A(G1966), .ZN(new_n771));
  INV_X1    g346(.A(new_n763), .ZN(new_n772));
  OAI21_X1  g347(.A(new_n770), .B1(new_n771), .B2(new_n772), .ZN(new_n773));
  NOR4_X1   g348(.A1(new_n761), .A2(new_n764), .A3(new_n769), .A4(new_n773), .ZN(new_n774));
  NAND4_X1  g349(.A1(new_n740), .A2(new_n744), .A3(new_n753), .A4(new_n774), .ZN(new_n775));
  XNOR2_X1  g350(.A(new_n775), .B(KEYINPUT98), .ZN(new_n776));
  OAI211_X1 g351(.A(new_n727), .B(new_n776), .C1(new_n726), .C2(new_n725), .ZN(new_n777));
  NAND2_X1  g352(.A1(new_n694), .A2(G22), .ZN(new_n778));
  OAI21_X1  g353(.A(new_n778), .B1(G166), .B2(new_n694), .ZN(new_n779));
  XNOR2_X1  g354(.A(KEYINPUT91), .B(G1971), .ZN(new_n780));
  OR2_X1    g355(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  NOR2_X1   g356(.A1(G6), .A2(G16), .ZN(new_n782));
  AOI21_X1  g357(.A(new_n782), .B1(new_n583), .B2(G16), .ZN(new_n783));
  XOR2_X1   g358(.A(KEYINPUT32), .B(G1981), .Z(new_n784));
  XNOR2_X1  g359(.A(new_n783), .B(new_n784), .ZN(new_n785));
  NAND2_X1  g360(.A1(new_n694), .A2(G23), .ZN(new_n786));
  INV_X1    g361(.A(G288), .ZN(new_n787));
  OAI21_X1  g362(.A(new_n786), .B1(new_n787), .B2(new_n694), .ZN(new_n788));
  XNOR2_X1  g363(.A(KEYINPUT33), .B(G1976), .ZN(new_n789));
  XNOR2_X1  g364(.A(new_n788), .B(new_n789), .ZN(new_n790));
  NAND3_X1  g365(.A1(new_n781), .A2(new_n785), .A3(new_n790), .ZN(new_n791));
  AOI21_X1  g366(.A(new_n791), .B1(new_n779), .B2(new_n780), .ZN(new_n792));
  INV_X1    g367(.A(KEYINPUT34), .ZN(new_n793));
  OR2_X1    g368(.A1(new_n792), .A2(new_n793), .ZN(new_n794));
  AND2_X1   g369(.A1(new_n590), .A2(new_n591), .ZN(new_n795));
  NAND2_X1  g370(.A1(new_n795), .A2(G16), .ZN(new_n796));
  OAI21_X1  g371(.A(new_n796), .B1(G16), .B2(G24), .ZN(new_n797));
  INV_X1    g372(.A(G1986), .ZN(new_n798));
  AND2_X1   g373(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  NOR2_X1   g374(.A1(new_n797), .A2(new_n798), .ZN(new_n800));
  INV_X1    g375(.A(KEYINPUT36), .ZN(new_n801));
  NOR2_X1   g376(.A1(new_n801), .A2(KEYINPUT92), .ZN(new_n802));
  MUX2_X1   g377(.A(G95), .B(G107), .S(G2105), .Z(new_n803));
  AOI22_X1  g378(.A1(new_n480), .A2(G131), .B1(G2104), .B2(new_n803), .ZN(new_n804));
  INV_X1    g379(.A(G119), .ZN(new_n805));
  OAI21_X1  g380(.A(new_n804), .B1(new_n489), .B2(new_n805), .ZN(new_n806));
  MUX2_X1   g381(.A(G25), .B(new_n806), .S(G29), .Z(new_n807));
  XNOR2_X1  g382(.A(KEYINPUT35), .B(G1991), .ZN(new_n808));
  XNOR2_X1  g383(.A(new_n807), .B(new_n808), .ZN(new_n809));
  NOR4_X1   g384(.A1(new_n799), .A2(new_n800), .A3(new_n802), .A4(new_n809), .ZN(new_n810));
  NAND2_X1  g385(.A1(new_n792), .A2(new_n793), .ZN(new_n811));
  NAND3_X1  g386(.A1(new_n794), .A2(new_n810), .A3(new_n811), .ZN(new_n812));
  NAND3_X1  g387(.A1(new_n812), .A2(KEYINPUT92), .A3(new_n801), .ZN(new_n813));
  INV_X1    g388(.A(new_n813), .ZN(new_n814));
  AOI21_X1  g389(.A(new_n812), .B1(KEYINPUT92), .B2(new_n801), .ZN(new_n815));
  NOR3_X1   g390(.A1(new_n777), .A2(new_n814), .A3(new_n815), .ZN(G311));
  INV_X1    g391(.A(G311), .ZN(G150));
  NAND2_X1  g392(.A1(new_n522), .A2(G55), .ZN(new_n818));
  INV_X1    g393(.A(G93), .ZN(new_n819));
  OAI21_X1  g394(.A(new_n818), .B1(new_n819), .B2(new_n541), .ZN(new_n820));
  AOI22_X1  g395(.A1(new_n516), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n821));
  NOR2_X1   g396(.A1(new_n821), .A2(new_n544), .ZN(new_n822));
  NOR2_X1   g397(.A1(new_n820), .A2(new_n822), .ZN(new_n823));
  INV_X1    g398(.A(new_n823), .ZN(new_n824));
  NAND2_X1  g399(.A1(new_n824), .A2(G860), .ZN(new_n825));
  XOR2_X1   g400(.A(new_n825), .B(KEYINPUT37), .Z(new_n826));
  NAND2_X1  g401(.A1(new_n599), .A2(G559), .ZN(new_n827));
  XNOR2_X1  g402(.A(new_n827), .B(KEYINPUT38), .ZN(new_n828));
  OR2_X1    g403(.A1(new_n552), .A2(KEYINPUT100), .ZN(new_n829));
  NAND2_X1  g404(.A1(new_n552), .A2(KEYINPUT100), .ZN(new_n830));
  NAND3_X1  g405(.A1(new_n829), .A2(new_n830), .A3(new_n824), .ZN(new_n831));
  NAND3_X1  g406(.A1(new_n552), .A2(new_n823), .A3(KEYINPUT100), .ZN(new_n832));
  NAND2_X1  g407(.A1(new_n831), .A2(new_n832), .ZN(new_n833));
  INV_X1    g408(.A(new_n833), .ZN(new_n834));
  XNOR2_X1  g409(.A(new_n828), .B(new_n834), .ZN(new_n835));
  NOR2_X1   g410(.A1(new_n835), .A2(KEYINPUT39), .ZN(new_n836));
  XOR2_X1   g411(.A(new_n836), .B(KEYINPUT101), .Z(new_n837));
  AOI21_X1  g412(.A(G860), .B1(new_n835), .B2(KEYINPUT39), .ZN(new_n838));
  NAND3_X1  g413(.A1(new_n837), .A2(KEYINPUT102), .A3(new_n838), .ZN(new_n839));
  INV_X1    g414(.A(new_n839), .ZN(new_n840));
  AOI21_X1  g415(.A(KEYINPUT102), .B1(new_n837), .B2(new_n838), .ZN(new_n841));
  OAI21_X1  g416(.A(new_n826), .B1(new_n840), .B2(new_n841), .ZN(G145));
  MUX2_X1   g417(.A(G106), .B(G118), .S(G2105), .Z(new_n843));
  AOI22_X1  g418(.A1(new_n480), .A2(G142), .B1(G2104), .B2(new_n843), .ZN(new_n844));
  INV_X1    g419(.A(G130), .ZN(new_n845));
  OAI21_X1  g420(.A(new_n844), .B1(new_n489), .B2(new_n845), .ZN(new_n846));
  XNOR2_X1  g421(.A(new_n806), .B(new_n846), .ZN(new_n847));
  XNOR2_X1  g422(.A(new_n847), .B(new_n620), .ZN(new_n848));
  XNOR2_X1  g423(.A(new_n708), .B(G164), .ZN(new_n849));
  XNOR2_X1  g424(.A(new_n848), .B(new_n849), .ZN(new_n850));
  XNOR2_X1  g425(.A(new_n738), .B(new_n750), .ZN(new_n851));
  OR2_X1    g426(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n850), .A2(new_n851), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  XNOR2_X1  g429(.A(G162), .B(G160), .ZN(new_n855));
  XNOR2_X1  g430(.A(new_n628), .B(KEYINPUT103), .ZN(new_n856));
  XNOR2_X1  g431(.A(new_n855), .B(new_n856), .ZN(new_n857));
  INV_X1    g432(.A(new_n857), .ZN(new_n858));
  NAND2_X1  g433(.A1(new_n854), .A2(new_n858), .ZN(new_n859));
  INV_X1    g434(.A(G37), .ZN(new_n860));
  NAND3_X1  g435(.A1(new_n852), .A2(new_n857), .A3(new_n853), .ZN(new_n861));
  NAND3_X1  g436(.A1(new_n859), .A2(new_n860), .A3(new_n861), .ZN(new_n862));
  XNOR2_X1  g437(.A(new_n862), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g438(.A1(new_n599), .A2(new_n610), .ZN(new_n864));
  XNOR2_X1  g439(.A(new_n833), .B(new_n864), .ZN(new_n865));
  XNOR2_X1  g440(.A(new_n599), .B(G299), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  XNOR2_X1  g442(.A(new_n866), .B(KEYINPUT41), .ZN(new_n868));
  OAI21_X1  g443(.A(new_n867), .B1(new_n868), .B2(new_n865), .ZN(new_n869));
  OR2_X1    g444(.A1(new_n869), .A2(KEYINPUT42), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n869), .A2(KEYINPUT42), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  XNOR2_X1  g447(.A(G290), .B(G288), .ZN(new_n873));
  XNOR2_X1  g448(.A(G166), .B(new_n583), .ZN(new_n874));
  XNOR2_X1  g449(.A(new_n873), .B(new_n874), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n872), .A2(new_n875), .ZN(new_n876));
  INV_X1    g451(.A(new_n875), .ZN(new_n877));
  NAND3_X1  g452(.A1(new_n870), .A2(new_n877), .A3(new_n871), .ZN(new_n878));
  NAND3_X1  g453(.A1(new_n876), .A2(G868), .A3(new_n878), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n879), .A2(KEYINPUT104), .ZN(new_n880));
  INV_X1    g455(.A(KEYINPUT104), .ZN(new_n881));
  NAND4_X1  g456(.A1(new_n876), .A2(new_n881), .A3(G868), .A4(new_n878), .ZN(new_n882));
  OAI211_X1 g457(.A(new_n880), .B(new_n882), .C1(G868), .C2(new_n823), .ZN(G295));
  OAI211_X1 g458(.A(new_n880), .B(new_n882), .C1(G868), .C2(new_n823), .ZN(G331));
  INV_X1    g459(.A(KEYINPUT43), .ZN(new_n885));
  INV_X1    g460(.A(G171), .ZN(new_n886));
  NOR2_X1   g461(.A1(new_n886), .A2(G168), .ZN(new_n887));
  INV_X1    g462(.A(new_n887), .ZN(new_n888));
  OAI21_X1  g463(.A(new_n888), .B1(new_n603), .B2(G286), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n834), .A2(new_n889), .ZN(new_n890));
  OAI211_X1 g465(.A(new_n833), .B(new_n888), .C1(G286), .C2(new_n603), .ZN(new_n891));
  NAND3_X1  g466(.A1(new_n890), .A2(new_n891), .A3(new_n866), .ZN(new_n892));
  AND2_X1   g467(.A1(new_n890), .A2(new_n891), .ZN(new_n893));
  OAI21_X1  g468(.A(new_n892), .B1(new_n893), .B2(new_n868), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n894), .A2(new_n877), .ZN(new_n895));
  INV_X1    g470(.A(KEYINPUT106), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  NAND3_X1  g472(.A1(new_n894), .A2(KEYINPUT106), .A3(new_n877), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  INV_X1    g474(.A(KEYINPUT105), .ZN(new_n900));
  OAI21_X1  g475(.A(new_n900), .B1(new_n894), .B2(new_n877), .ZN(new_n901));
  XOR2_X1   g476(.A(new_n866), .B(KEYINPUT41), .Z(new_n902));
  NAND2_X1  g477(.A1(new_n890), .A2(new_n891), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  NAND4_X1  g479(.A1(new_n904), .A2(KEYINPUT105), .A3(new_n875), .A4(new_n892), .ZN(new_n905));
  AOI21_X1  g480(.A(G37), .B1(new_n901), .B2(new_n905), .ZN(new_n906));
  AOI21_X1  g481(.A(new_n885), .B1(new_n899), .B2(new_n906), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n901), .A2(new_n905), .ZN(new_n908));
  AOI21_X1  g483(.A(G37), .B1(new_n894), .B2(new_n877), .ZN(new_n909));
  AND3_X1   g484(.A1(new_n908), .A2(new_n909), .A3(new_n885), .ZN(new_n910));
  OAI21_X1  g485(.A(KEYINPUT44), .B1(new_n907), .B2(new_n910), .ZN(new_n911));
  INV_X1    g486(.A(KEYINPUT44), .ZN(new_n912));
  AOI21_X1  g487(.A(KEYINPUT43), .B1(new_n899), .B2(new_n906), .ZN(new_n913));
  AND3_X1   g488(.A1(new_n908), .A2(new_n909), .A3(KEYINPUT43), .ZN(new_n914));
  OAI21_X1  g489(.A(new_n912), .B1(new_n913), .B2(new_n914), .ZN(new_n915));
  AND2_X1   g490(.A1(new_n911), .A2(new_n915), .ZN(G397));
  INV_X1    g491(.A(G1384), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n507), .A2(new_n917), .ZN(new_n918));
  INV_X1    g493(.A(G40), .ZN(new_n919));
  NOR3_X1   g494(.A1(new_n473), .A2(new_n477), .A3(new_n919), .ZN(new_n920));
  XNOR2_X1  g495(.A(KEYINPUT107), .B(KEYINPUT45), .ZN(new_n921));
  NAND3_X1  g496(.A1(new_n918), .A2(new_n920), .A3(new_n921), .ZN(new_n922));
  INV_X1    g497(.A(new_n922), .ZN(new_n923));
  NOR2_X1   g498(.A1(new_n708), .A2(new_n710), .ZN(new_n924));
  NOR3_X1   g499(.A1(new_n706), .A2(new_n707), .A3(G2067), .ZN(new_n925));
  NOR2_X1   g500(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  XNOR2_X1  g501(.A(new_n750), .B(G1996), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  AND2_X1   g503(.A1(new_n806), .A2(new_n808), .ZN(new_n929));
  NOR2_X1   g504(.A1(new_n806), .A2(new_n808), .ZN(new_n930));
  OR3_X1    g505(.A1(new_n928), .A2(new_n929), .A3(new_n930), .ZN(new_n931));
  XNOR2_X1  g506(.A(G290), .B(G1986), .ZN(new_n932));
  OAI21_X1  g507(.A(new_n923), .B1(new_n931), .B2(new_n932), .ZN(new_n933));
  INV_X1    g508(.A(KEYINPUT123), .ZN(new_n934));
  NOR2_X1   g509(.A1(new_n502), .A2(new_n503), .ZN(new_n935));
  INV_X1    g510(.A(G125), .ZN(new_n936));
  OAI21_X1  g511(.A(new_n472), .B1(new_n935), .B2(new_n936), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n937), .A2(G2105), .ZN(new_n938));
  NAND4_X1  g513(.A1(new_n938), .A2(G40), .A3(new_n476), .A4(new_n474), .ZN(new_n939));
  NOR2_X1   g514(.A1(new_n918), .A2(new_n939), .ZN(new_n940));
  INV_X1    g515(.A(G8), .ZN(new_n941));
  NOR2_X1   g516(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  NOR3_X1   g517(.A1(new_n580), .A2(new_n582), .A3(G1981), .ZN(new_n943));
  INV_X1    g518(.A(new_n943), .ZN(new_n944));
  OAI21_X1  g519(.A(G1981), .B1(new_n580), .B2(new_n582), .ZN(new_n945));
  NAND3_X1  g520(.A1(new_n944), .A2(KEYINPUT49), .A3(new_n945), .ZN(new_n946));
  INV_X1    g521(.A(KEYINPUT49), .ZN(new_n947));
  INV_X1    g522(.A(new_n945), .ZN(new_n948));
  OAI21_X1  g523(.A(new_n947), .B1(new_n948), .B2(new_n943), .ZN(new_n949));
  NAND3_X1  g524(.A1(new_n946), .A2(new_n949), .A3(new_n942), .ZN(new_n950));
  INV_X1    g525(.A(G1976), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n787), .A2(new_n951), .ZN(new_n952));
  XNOR2_X1  g527(.A(new_n952), .B(KEYINPUT110), .ZN(new_n953));
  AND2_X1   g528(.A1(new_n950), .A2(new_n953), .ZN(new_n954));
  OAI21_X1  g529(.A(new_n942), .B1(new_n954), .B2(new_n943), .ZN(new_n955));
  INV_X1    g530(.A(KEYINPUT109), .ZN(new_n956));
  INV_X1    g531(.A(KEYINPUT55), .ZN(new_n957));
  NOR2_X1   g532(.A1(new_n956), .A2(new_n957), .ZN(new_n958));
  INV_X1    g533(.A(new_n958), .ZN(new_n959));
  OAI21_X1  g534(.A(G8), .B1(KEYINPUT109), .B2(KEYINPUT55), .ZN(new_n960));
  INV_X1    g535(.A(new_n960), .ZN(new_n961));
  AOI21_X1  g536(.A(new_n959), .B1(G303), .B2(new_n961), .ZN(new_n962));
  NOR4_X1   g537(.A1(new_n571), .A2(new_n572), .A3(new_n960), .A4(new_n958), .ZN(new_n963));
  NOR2_X1   g538(.A1(new_n962), .A2(new_n963), .ZN(new_n964));
  AOI21_X1  g539(.A(new_n939), .B1(new_n918), .B2(new_n921), .ZN(new_n965));
  AND2_X1   g540(.A1(KEYINPUT4), .A2(G138), .ZN(new_n966));
  OAI21_X1  g541(.A(new_n966), .B1(new_n502), .B2(new_n503), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n967), .A2(new_n499), .ZN(new_n968));
  AOI22_X1  g543(.A1(new_n968), .A2(new_n465), .B1(new_n505), .B2(new_n504), .ZN(new_n969));
  AOI21_X1  g544(.A(G1384), .B1(new_n969), .B2(new_n496), .ZN(new_n970));
  AOI21_X1  g545(.A(KEYINPUT108), .B1(new_n970), .B2(KEYINPUT45), .ZN(new_n971));
  AND4_X1   g546(.A1(KEYINPUT108), .A2(new_n507), .A3(KEYINPUT45), .A4(new_n917), .ZN(new_n972));
  OAI21_X1  g547(.A(new_n965), .B1(new_n971), .B2(new_n972), .ZN(new_n973));
  INV_X1    g548(.A(G1971), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n973), .A2(new_n974), .ZN(new_n975));
  INV_X1    g550(.A(KEYINPUT50), .ZN(new_n976));
  OAI21_X1  g551(.A(new_n920), .B1(new_n970), .B2(new_n976), .ZN(new_n977));
  NAND3_X1  g552(.A1(new_n507), .A2(new_n976), .A3(new_n917), .ZN(new_n978));
  INV_X1    g553(.A(new_n978), .ZN(new_n979));
  NOR2_X1   g554(.A1(new_n977), .A2(new_n979), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n980), .A2(new_n726), .ZN(new_n981));
  AOI21_X1  g556(.A(new_n941), .B1(new_n975), .B2(new_n981), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n964), .A2(new_n982), .ZN(new_n983));
  NAND2_X1  g558(.A1(new_n787), .A2(G1976), .ZN(new_n984));
  AOI21_X1  g559(.A(KEYINPUT52), .B1(G288), .B2(new_n951), .ZN(new_n985));
  NAND3_X1  g560(.A1(new_n942), .A2(new_n984), .A3(new_n985), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n970), .A2(new_n920), .ZN(new_n987));
  NAND3_X1  g562(.A1(new_n987), .A2(G8), .A3(new_n984), .ZN(new_n988));
  NAND2_X1  g563(.A1(new_n988), .A2(KEYINPUT52), .ZN(new_n989));
  NAND3_X1  g564(.A1(new_n950), .A2(new_n986), .A3(new_n989), .ZN(new_n990));
  OAI21_X1  g565(.A(new_n955), .B1(new_n983), .B2(new_n990), .ZN(new_n991));
  AOI21_X1  g566(.A(new_n990), .B1(new_n964), .B2(new_n982), .ZN(new_n992));
  AOI21_X1  g567(.A(KEYINPUT45), .B1(new_n507), .B2(new_n917), .ZN(new_n993));
  OAI21_X1  g568(.A(KEYINPUT113), .B1(new_n993), .B2(new_n939), .ZN(new_n994));
  INV_X1    g569(.A(KEYINPUT113), .ZN(new_n995));
  OAI211_X1 g570(.A(new_n920), .B(new_n995), .C1(new_n970), .C2(KEYINPUT45), .ZN(new_n996));
  OR2_X1    g571(.A1(new_n918), .A2(new_n921), .ZN(new_n997));
  NAND3_X1  g572(.A1(new_n994), .A2(new_n996), .A3(new_n997), .ZN(new_n998));
  XOR2_X1   g573(.A(KEYINPUT114), .B(G2084), .Z(new_n999));
  INV_X1    g574(.A(new_n999), .ZN(new_n1000));
  AOI22_X1  g575(.A1(new_n998), .A2(new_n771), .B1(new_n980), .B2(new_n1000), .ZN(new_n1001));
  NOR3_X1   g576(.A1(new_n1001), .A2(new_n941), .A3(G286), .ZN(new_n1002));
  INV_X1    g577(.A(KEYINPUT112), .ZN(new_n1003));
  AOI21_X1  g578(.A(new_n939), .B1(new_n918), .B2(KEYINPUT50), .ZN(new_n1004));
  INV_X1    g579(.A(KEYINPUT111), .ZN(new_n1005));
  AOI21_X1  g580(.A(new_n1005), .B1(new_n970), .B2(new_n976), .ZN(new_n1006));
  NAND4_X1  g581(.A1(new_n507), .A2(new_n1005), .A3(new_n976), .A4(new_n917), .ZN(new_n1007));
  INV_X1    g582(.A(new_n1007), .ZN(new_n1008));
  OAI211_X1 g583(.A(new_n1003), .B(new_n1004), .C1(new_n1006), .C2(new_n1008), .ZN(new_n1009));
  INV_X1    g584(.A(new_n1009), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n978), .A2(KEYINPUT111), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n1011), .A2(new_n1007), .ZN(new_n1012));
  AOI21_X1  g587(.A(new_n1003), .B1(new_n1012), .B2(new_n1004), .ZN(new_n1013));
  OAI21_X1  g588(.A(new_n726), .B1(new_n1010), .B2(new_n1013), .ZN(new_n1014));
  AOI21_X1  g589(.A(new_n941), .B1(new_n1014), .B2(new_n975), .ZN(new_n1015));
  OAI211_X1 g590(.A(new_n992), .B(new_n1002), .C1(new_n1015), .C2(new_n964), .ZN(new_n1016));
  XNOR2_X1  g591(.A(KEYINPUT115), .B(KEYINPUT63), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n1016), .A2(new_n1017), .ZN(new_n1018));
  OR2_X1    g593(.A1(new_n964), .A2(new_n982), .ZN(new_n1019));
  NAND4_X1  g594(.A1(new_n1019), .A2(new_n992), .A3(KEYINPUT63), .A4(new_n1002), .ZN(new_n1020));
  AOI21_X1  g595(.A(new_n991), .B1(new_n1018), .B2(new_n1020), .ZN(new_n1021));
  AOI21_X1  g596(.A(new_n716), .B1(new_n1004), .B2(new_n978), .ZN(new_n1022));
  NOR2_X1   g597(.A1(new_n987), .A2(G2067), .ZN(new_n1023));
  OAI21_X1  g598(.A(KEYINPUT116), .B1(new_n1022), .B2(new_n1023), .ZN(new_n1024));
  OAI21_X1  g599(.A(new_n715), .B1(new_n977), .B2(new_n979), .ZN(new_n1025));
  INV_X1    g600(.A(KEYINPUT116), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n940), .A2(new_n710), .ZN(new_n1027));
  NAND3_X1  g602(.A1(new_n1025), .A2(new_n1026), .A3(new_n1027), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n1024), .A2(new_n1028), .ZN(new_n1029));
  INV_X1    g604(.A(new_n1029), .ZN(new_n1030));
  INV_X1    g605(.A(KEYINPUT57), .ZN(new_n1031));
  XNOR2_X1  g606(.A(G299), .B(new_n1031), .ZN(new_n1032));
  XNOR2_X1  g607(.A(KEYINPUT56), .B(G2072), .ZN(new_n1033));
  OAI211_X1 g608(.A(new_n965), .B(new_n1033), .C1(new_n971), .C2(new_n972), .ZN(new_n1034));
  AOI21_X1  g609(.A(new_n977), .B1(new_n1011), .B2(new_n1007), .ZN(new_n1035));
  OAI211_X1 g610(.A(new_n1032), .B(new_n1034), .C1(G1956), .C2(new_n1035), .ZN(new_n1036));
  NAND3_X1  g611(.A1(new_n1030), .A2(new_n599), .A3(new_n1036), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n1012), .A2(new_n1004), .ZN(new_n1038));
  INV_X1    g613(.A(G1956), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n1038), .A2(new_n1039), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n1040), .A2(new_n1034), .ZN(new_n1041));
  INV_X1    g616(.A(new_n1032), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n1041), .A2(new_n1042), .ZN(new_n1043));
  NAND2_X1  g618(.A1(new_n1037), .A2(new_n1043), .ZN(new_n1044));
  NOR3_X1   g619(.A1(new_n1022), .A2(KEYINPUT116), .A3(new_n1023), .ZN(new_n1045));
  AOI21_X1  g620(.A(new_n1026), .B1(new_n1025), .B2(new_n1027), .ZN(new_n1046));
  OAI21_X1  g621(.A(KEYINPUT60), .B1(new_n1045), .B2(new_n1046), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n1047), .A2(new_n599), .ZN(new_n1048));
  NAND3_X1  g623(.A1(new_n1029), .A2(KEYINPUT60), .A3(new_n600), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n1048), .A2(new_n1049), .ZN(new_n1050));
  INV_X1    g625(.A(KEYINPUT60), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n1030), .A2(new_n1051), .ZN(new_n1052));
  INV_X1    g627(.A(new_n1036), .ZN(new_n1053));
  AOI21_X1  g628(.A(new_n1032), .B1(new_n1040), .B2(new_n1034), .ZN(new_n1054));
  OAI21_X1  g629(.A(KEYINPUT61), .B1(new_n1053), .B2(new_n1054), .ZN(new_n1055));
  INV_X1    g630(.A(KEYINPUT61), .ZN(new_n1056));
  NAND3_X1  g631(.A1(new_n1043), .A2(new_n1056), .A3(new_n1036), .ZN(new_n1057));
  AOI22_X1  g632(.A1(new_n1050), .A2(new_n1052), .B1(new_n1055), .B2(new_n1057), .ZN(new_n1058));
  INV_X1    g633(.A(KEYINPUT118), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n1059), .A2(KEYINPUT59), .ZN(new_n1060));
  NOR2_X1   g635(.A1(new_n1059), .A2(KEYINPUT59), .ZN(new_n1061));
  INV_X1    g636(.A(new_n1061), .ZN(new_n1062));
  OAI21_X1  g637(.A(KEYINPUT117), .B1(new_n973), .B2(G1996), .ZN(new_n1063));
  NAND3_X1  g638(.A1(new_n507), .A2(KEYINPUT45), .A3(new_n917), .ZN(new_n1064));
  INV_X1    g639(.A(KEYINPUT108), .ZN(new_n1065));
  XNOR2_X1  g640(.A(new_n1064), .B(new_n1065), .ZN(new_n1066));
  INV_X1    g641(.A(KEYINPUT117), .ZN(new_n1067));
  INV_X1    g642(.A(G1996), .ZN(new_n1068));
  NAND4_X1  g643(.A1(new_n1066), .A2(new_n1067), .A3(new_n1068), .A4(new_n965), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n1063), .A2(new_n1069), .ZN(new_n1070));
  XOR2_X1   g645(.A(KEYINPUT58), .B(G1341), .Z(new_n1071));
  NAND2_X1  g646(.A1(new_n987), .A2(new_n1071), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n1070), .A2(new_n1072), .ZN(new_n1073));
  AOI21_X1  g648(.A(new_n1062), .B1(new_n1073), .B2(new_n552), .ZN(new_n1074));
  AOI22_X1  g649(.A1(new_n1063), .A2(new_n1069), .B1(new_n987), .B2(new_n1071), .ZN(new_n1075));
  INV_X1    g650(.A(new_n552), .ZN(new_n1076));
  NOR3_X1   g651(.A1(new_n1075), .A2(new_n1076), .A3(new_n1061), .ZN(new_n1077));
  OAI21_X1  g652(.A(new_n1060), .B1(new_n1074), .B2(new_n1077), .ZN(new_n1078));
  AOI21_X1  g653(.A(new_n1044), .B1(new_n1058), .B2(new_n1078), .ZN(new_n1079));
  OAI21_X1  g654(.A(new_n992), .B1(new_n1015), .B2(new_n964), .ZN(new_n1080));
  INV_X1    g655(.A(G2078), .ZN(new_n1081));
  OAI211_X1 g656(.A(new_n1081), .B(new_n965), .C1(new_n971), .C2(new_n972), .ZN(new_n1082));
  INV_X1    g657(.A(KEYINPUT53), .ZN(new_n1083));
  INV_X1    g658(.A(G1961), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n1004), .A2(new_n978), .ZN(new_n1085));
  AOI22_X1  g660(.A1(new_n1082), .A2(new_n1083), .B1(new_n1084), .B2(new_n1085), .ZN(new_n1086));
  NOR2_X1   g661(.A1(new_n918), .A2(new_n921), .ZN(new_n1087));
  OAI21_X1  g662(.A(new_n920), .B1(new_n970), .B2(KEYINPUT45), .ZN(new_n1088));
  AOI21_X1  g663(.A(new_n1087), .B1(new_n1088), .B2(KEYINPUT113), .ZN(new_n1089));
  NAND4_X1  g664(.A1(new_n1089), .A2(KEYINPUT53), .A3(new_n1081), .A4(new_n996), .ZN(new_n1090));
  AND3_X1   g665(.A1(new_n1086), .A2(G301), .A3(new_n1090), .ZN(new_n1091));
  NAND4_X1  g666(.A1(new_n1066), .A2(KEYINPUT53), .A3(new_n1081), .A4(new_n965), .ZN(new_n1092));
  AOI21_X1  g667(.A(new_n886), .B1(new_n1086), .B2(new_n1092), .ZN(new_n1093));
  INV_X1    g668(.A(KEYINPUT54), .ZN(new_n1094));
  NOR3_X1   g669(.A1(new_n1091), .A2(new_n1093), .A3(new_n1094), .ZN(new_n1095));
  NOR2_X1   g670(.A1(new_n1080), .A2(new_n1095), .ZN(new_n1096));
  OAI21_X1  g671(.A(KEYINPUT122), .B1(new_n1001), .B2(new_n941), .ZN(new_n1097));
  INV_X1    g672(.A(KEYINPUT122), .ZN(new_n1098));
  AOI21_X1  g673(.A(G1966), .B1(new_n1089), .B2(new_n996), .ZN(new_n1099));
  NOR2_X1   g674(.A1(new_n1085), .A2(new_n999), .ZN(new_n1100));
  OAI211_X1 g675(.A(new_n1098), .B(G8), .C1(new_n1099), .C2(new_n1100), .ZN(new_n1101));
  NAND3_X1  g676(.A1(G286), .A2(KEYINPUT119), .A3(G8), .ZN(new_n1102));
  INV_X1    g677(.A(KEYINPUT119), .ZN(new_n1103));
  OAI21_X1  g678(.A(new_n1103), .B1(G168), .B2(new_n941), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n1102), .A2(new_n1104), .ZN(new_n1105));
  NOR2_X1   g680(.A1(new_n1105), .A2(KEYINPUT51), .ZN(new_n1106));
  NAND3_X1  g681(.A1(new_n1097), .A2(new_n1101), .A3(new_n1106), .ZN(new_n1107));
  XNOR2_X1  g682(.A(KEYINPUT120), .B(KEYINPUT51), .ZN(new_n1108));
  NAND2_X1  g683(.A1(new_n998), .A2(new_n771), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n980), .A2(new_n1000), .ZN(new_n1110));
  AOI21_X1  g685(.A(new_n941), .B1(new_n1109), .B2(new_n1110), .ZN(new_n1111));
  XNOR2_X1  g686(.A(new_n1105), .B(KEYINPUT121), .ZN(new_n1112));
  OAI21_X1  g687(.A(new_n1108), .B1(new_n1111), .B2(new_n1112), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n1107), .A2(new_n1113), .ZN(new_n1114));
  AOI21_X1  g689(.A(new_n1001), .B1(new_n1102), .B2(new_n1104), .ZN(new_n1115));
  INV_X1    g690(.A(new_n1115), .ZN(new_n1116));
  NAND2_X1  g691(.A1(new_n1114), .A2(new_n1116), .ZN(new_n1117));
  AND3_X1   g692(.A1(new_n1086), .A2(G301), .A3(new_n1092), .ZN(new_n1118));
  AOI21_X1  g693(.A(G301), .B1(new_n1086), .B2(new_n1090), .ZN(new_n1119));
  OAI21_X1  g694(.A(new_n1094), .B1(new_n1118), .B2(new_n1119), .ZN(new_n1120));
  NAND3_X1  g695(.A1(new_n1096), .A2(new_n1117), .A3(new_n1120), .ZN(new_n1121));
  OAI211_X1 g696(.A(new_n934), .B(new_n1021), .C1(new_n1079), .C2(new_n1121), .ZN(new_n1122));
  OR2_X1    g697(.A1(new_n1117), .A2(KEYINPUT62), .ZN(new_n1123));
  INV_X1    g698(.A(new_n1080), .ZN(new_n1124));
  NAND2_X1  g699(.A1(new_n1117), .A2(KEYINPUT62), .ZN(new_n1125));
  NAND4_X1  g700(.A1(new_n1123), .A2(new_n1119), .A3(new_n1124), .A4(new_n1125), .ZN(new_n1126));
  NAND2_X1  g701(.A1(new_n1122), .A2(new_n1126), .ZN(new_n1127));
  INV_X1    g702(.A(new_n964), .ZN(new_n1128));
  AND2_X1   g703(.A1(new_n1014), .A2(new_n975), .ZN(new_n1129));
  OAI21_X1  g704(.A(new_n1128), .B1(new_n1129), .B2(new_n941), .ZN(new_n1130));
  NAND3_X1  g705(.A1(new_n1086), .A2(G301), .A3(new_n1090), .ZN(new_n1131));
  AND2_X1   g706(.A1(new_n1086), .A2(new_n1092), .ZN(new_n1132));
  OAI211_X1 g707(.A(KEYINPUT54), .B(new_n1131), .C1(new_n1132), .C2(new_n886), .ZN(new_n1133));
  NAND4_X1  g708(.A1(new_n1130), .A2(new_n1120), .A3(new_n1133), .A4(new_n992), .ZN(new_n1134));
  AOI21_X1  g709(.A(new_n1115), .B1(new_n1107), .B2(new_n1113), .ZN(new_n1135));
  NOR2_X1   g710(.A1(new_n1134), .A2(new_n1135), .ZN(new_n1136));
  INV_X1    g711(.A(new_n1044), .ZN(new_n1137));
  NAND2_X1  g712(.A1(new_n1055), .A2(new_n1057), .ZN(new_n1138));
  AOI21_X1  g713(.A(new_n600), .B1(new_n1029), .B2(KEYINPUT60), .ZN(new_n1139));
  AOI211_X1 g714(.A(new_n1051), .B(new_n599), .C1(new_n1024), .C2(new_n1028), .ZN(new_n1140));
  OAI21_X1  g715(.A(new_n1052), .B1(new_n1139), .B2(new_n1140), .ZN(new_n1141));
  NAND2_X1  g716(.A1(new_n1138), .A2(new_n1141), .ZN(new_n1142));
  NAND3_X1  g717(.A1(new_n1073), .A2(new_n552), .A3(new_n1062), .ZN(new_n1143));
  OAI21_X1  g718(.A(new_n1061), .B1(new_n1075), .B2(new_n1076), .ZN(new_n1144));
  AOI22_X1  g719(.A1(new_n1143), .A2(new_n1144), .B1(new_n1059), .B2(KEYINPUT59), .ZN(new_n1145));
  OAI21_X1  g720(.A(new_n1137), .B1(new_n1142), .B2(new_n1145), .ZN(new_n1146));
  NAND2_X1  g721(.A1(new_n1136), .A2(new_n1146), .ZN(new_n1147));
  AOI21_X1  g722(.A(new_n934), .B1(new_n1147), .B2(new_n1021), .ZN(new_n1148));
  OAI21_X1  g723(.A(new_n933), .B1(new_n1127), .B2(new_n1148), .ZN(new_n1149));
  AOI21_X1  g724(.A(new_n922), .B1(new_n926), .B2(new_n750), .ZN(new_n1150));
  XNOR2_X1  g725(.A(new_n1150), .B(KEYINPUT126), .ZN(new_n1151));
  INV_X1    g726(.A(KEYINPUT125), .ZN(new_n1152));
  INV_X1    g727(.A(KEYINPUT46), .ZN(new_n1153));
  OAI211_X1 g728(.A(new_n1152), .B(new_n1153), .C1(new_n922), .C2(G1996), .ZN(new_n1154));
  OAI22_X1  g729(.A1(new_n922), .A2(G1996), .B1(new_n1152), .B2(new_n1153), .ZN(new_n1155));
  OAI21_X1  g730(.A(new_n1155), .B1(KEYINPUT125), .B2(KEYINPUT46), .ZN(new_n1156));
  NAND3_X1  g731(.A1(new_n1151), .A2(new_n1154), .A3(new_n1156), .ZN(new_n1157));
  XNOR2_X1  g732(.A(new_n1157), .B(KEYINPUT47), .ZN(new_n1158));
  NAND2_X1  g733(.A1(new_n928), .A2(new_n923), .ZN(new_n1159));
  AOI21_X1  g734(.A(new_n925), .B1(new_n1159), .B2(new_n930), .ZN(new_n1160));
  OR2_X1    g735(.A1(new_n1160), .A2(KEYINPUT124), .ZN(new_n1161));
  AOI21_X1  g736(.A(new_n922), .B1(new_n1160), .B2(KEYINPUT124), .ZN(new_n1162));
  NOR2_X1   g737(.A1(G290), .A2(G1986), .ZN(new_n1163));
  AOI21_X1  g738(.A(KEYINPUT48), .B1(new_n1163), .B2(new_n923), .ZN(new_n1164));
  AOI21_X1  g739(.A(new_n1164), .B1(new_n931), .B2(new_n923), .ZN(new_n1165));
  NAND3_X1  g740(.A1(new_n1163), .A2(KEYINPUT48), .A3(new_n923), .ZN(new_n1166));
  AOI22_X1  g741(.A1(new_n1161), .A2(new_n1162), .B1(new_n1165), .B2(new_n1166), .ZN(new_n1167));
  AND2_X1   g742(.A1(new_n1158), .A2(new_n1167), .ZN(new_n1168));
  NAND2_X1  g743(.A1(new_n1149), .A2(new_n1168), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g744(.A1(G227), .A2(new_n463), .ZN(new_n1171));
  NAND2_X1  g745(.A1(new_n692), .A2(new_n1171), .ZN(new_n1172));
  OAI21_X1  g746(.A(KEYINPUT127), .B1(G401), .B2(new_n1172), .ZN(new_n1173));
  INV_X1    g747(.A(new_n641), .ZN(new_n1174));
  NAND2_X1  g748(.A1(new_n1174), .A2(new_n644), .ZN(new_n1175));
  NAND3_X1  g749(.A1(new_n1175), .A2(new_n646), .A3(G14), .ZN(new_n1176));
  INV_X1    g750(.A(KEYINPUT127), .ZN(new_n1177));
  NAND4_X1  g751(.A1(new_n1176), .A2(new_n1177), .A3(new_n692), .A4(new_n1171), .ZN(new_n1178));
  NAND3_X1  g752(.A1(new_n1173), .A2(new_n862), .A3(new_n1178), .ZN(new_n1179));
  NOR3_X1   g753(.A1(new_n1179), .A2(new_n913), .A3(new_n914), .ZN(G308));
  NOR2_X1   g754(.A1(new_n913), .A2(new_n914), .ZN(new_n1181));
  NAND4_X1  g755(.A1(new_n1181), .A2(new_n862), .A3(new_n1178), .A4(new_n1173), .ZN(G225));
endmodule


