//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 0 1 0 1 0 1 1 1 0 1 1 0 0 1 1 1 0 1 1 1 0 1 1 0 0 0 0 0 0 0 0 0 0 0 1 1 1 1 1 0 0 0 1 1 0 0 1 1 0 1 0 1 0 1 1 0 0 1 0 0 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:35:04 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n205, new_n206, new_n207, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n236, new_n237,
    new_n238, new_n240, new_n241, new_n242, new_n243, new_n244, new_n245,
    new_n246, new_n247, new_n249, new_n250, new_n251, new_n252, new_n253,
    new_n254, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1185, new_n1186, new_n1187,
    new_n1188, new_n1189, new_n1190, new_n1191, new_n1192, new_n1193,
    new_n1194, new_n1195, new_n1196, new_n1197, new_n1198, new_n1199,
    new_n1200, new_n1201, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1217, new_n1218,
    new_n1219, new_n1220, new_n1221, new_n1222, new_n1223, new_n1224,
    new_n1225, new_n1226, new_n1227, new_n1228, new_n1229, new_n1231,
    new_n1232, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1290, new_n1291, new_n1292, new_n1293,
    new_n1294, new_n1295, new_n1296, new_n1297;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  INV_X1    g0004(.A(G97), .ZN(new_n205));
  INV_X1    g0005(.A(G107), .ZN(new_n206));
  NAND2_X1  g0006(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  NAND2_X1  g0007(.A1(new_n207), .A2(G87), .ZN(G355));
  INV_X1    g0008(.A(G1), .ZN(new_n209));
  INV_X1    g0009(.A(G20), .ZN(new_n210));
  NOR2_X1   g0010(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  INV_X1    g0011(.A(new_n211), .ZN(new_n212));
  AOI22_X1  g0012(.A1(G77), .A2(G244), .B1(G97), .B2(G257), .ZN(new_n213));
  INV_X1    g0013(.A(G87), .ZN(new_n214));
  INV_X1    g0014(.A(G250), .ZN(new_n215));
  INV_X1    g0015(.A(G116), .ZN(new_n216));
  INV_X1    g0016(.A(G270), .ZN(new_n217));
  OAI221_X1 g0017(.A(new_n213), .B1(new_n214), .B2(new_n215), .C1(new_n216), .C2(new_n217), .ZN(new_n218));
  AOI21_X1  g0018(.A(new_n218), .B1(G50), .B2(G226), .ZN(new_n219));
  INV_X1    g0019(.A(G58), .ZN(new_n220));
  INV_X1    g0020(.A(G232), .ZN(new_n221));
  INV_X1    g0021(.A(G264), .ZN(new_n222));
  OAI221_X1 g0022(.A(new_n219), .B1(new_n220), .B2(new_n221), .C1(new_n206), .C2(new_n222), .ZN(new_n223));
  INV_X1    g0023(.A(G68), .ZN(new_n224));
  INV_X1    g0024(.A(G238), .ZN(new_n225));
  NOR2_X1   g0025(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  OAI21_X1  g0026(.A(new_n212), .B1(new_n223), .B2(new_n226), .ZN(new_n227));
  XNOR2_X1  g0027(.A(new_n227), .B(KEYINPUT64), .ZN(new_n228));
  XNOR2_X1  g0028(.A(new_n228), .B(KEYINPUT1), .ZN(new_n229));
  NOR2_X1   g0029(.A1(new_n212), .A2(G13), .ZN(new_n230));
  OAI211_X1 g0030(.A(new_n230), .B(G250), .C1(G257), .C2(G264), .ZN(new_n231));
  XOR2_X1   g0031(.A(new_n231), .B(KEYINPUT0), .Z(new_n232));
  NAND2_X1  g0032(.A1(G1), .A2(G13), .ZN(new_n233));
  NOR2_X1   g0033(.A1(new_n233), .A2(new_n210), .ZN(new_n234));
  OAI21_X1  g0034(.A(G50), .B1(G58), .B2(G68), .ZN(new_n235));
  INV_X1    g0035(.A(new_n235), .ZN(new_n236));
  AOI21_X1  g0036(.A(new_n232), .B1(new_n234), .B2(new_n236), .ZN(new_n237));
  NAND2_X1  g0037(.A1(new_n229), .A2(new_n237), .ZN(new_n238));
  XOR2_X1   g0038(.A(new_n238), .B(KEYINPUT65), .Z(G361));
  XNOR2_X1  g0039(.A(G238), .B(G244), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n240), .B(new_n221), .ZN(new_n241));
  XOR2_X1   g0041(.A(KEYINPUT2), .B(G226), .Z(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XNOR2_X1  g0043(.A(G250), .B(G257), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n244), .B(new_n217), .ZN(new_n245));
  XOR2_X1   g0045(.A(KEYINPUT66), .B(G264), .Z(new_n246));
  XNOR2_X1  g0046(.A(new_n245), .B(new_n246), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n243), .B(new_n247), .ZN(G358));
  XOR2_X1   g0048(.A(G87), .B(G97), .Z(new_n249));
  XNOR2_X1  g0049(.A(G107), .B(G116), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n249), .B(new_n250), .ZN(new_n251));
  XOR2_X1   g0051(.A(G68), .B(G77), .Z(new_n252));
  XNOR2_X1  g0052(.A(G50), .B(G58), .ZN(new_n253));
  XNOR2_X1  g0053(.A(new_n252), .B(new_n253), .ZN(new_n254));
  XNOR2_X1  g0054(.A(new_n251), .B(new_n254), .ZN(G351));
  NOR2_X1   g0055(.A1(KEYINPUT3), .A2(G33), .ZN(new_n256));
  XNOR2_X1  g0056(.A(KEYINPUT72), .B(KEYINPUT3), .ZN(new_n257));
  AOI21_X1  g0057(.A(new_n256), .B1(new_n257), .B2(G33), .ZN(new_n258));
  INV_X1    g0058(.A(KEYINPUT7), .ZN(new_n259));
  NAND3_X1  g0059(.A1(new_n258), .A2(new_n259), .A3(new_n210), .ZN(new_n260));
  INV_X1    g0060(.A(KEYINPUT3), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n261), .A2(KEYINPUT72), .ZN(new_n262));
  INV_X1    g0062(.A(KEYINPUT72), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n263), .A2(KEYINPUT3), .ZN(new_n264));
  NAND3_X1  g0064(.A1(new_n262), .A2(new_n264), .A3(G33), .ZN(new_n265));
  INV_X1    g0065(.A(G33), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n261), .A2(new_n266), .ZN(new_n267));
  NAND3_X1  g0067(.A1(new_n265), .A2(new_n210), .A3(new_n267), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n268), .A2(KEYINPUT7), .ZN(new_n269));
  NAND3_X1  g0069(.A1(new_n260), .A2(new_n269), .A3(G68), .ZN(new_n270));
  NOR2_X1   g0070(.A1(new_n220), .A2(new_n224), .ZN(new_n271));
  OR2_X1    g0071(.A1(new_n271), .A2(new_n201), .ZN(new_n272));
  NOR2_X1   g0072(.A1(G20), .A2(G33), .ZN(new_n273));
  AOI22_X1  g0073(.A1(new_n272), .A2(G20), .B1(G159), .B2(new_n273), .ZN(new_n274));
  NAND3_X1  g0074(.A1(new_n270), .A2(KEYINPUT16), .A3(new_n274), .ZN(new_n275));
  NOR2_X1   g0075(.A1(new_n263), .A2(KEYINPUT3), .ZN(new_n276));
  NOR2_X1   g0076(.A1(new_n261), .A2(KEYINPUT72), .ZN(new_n277));
  OAI21_X1  g0077(.A(new_n266), .B1(new_n276), .B2(new_n277), .ZN(new_n278));
  AND2_X1   g0078(.A1(KEYINPUT3), .A2(G33), .ZN(new_n279));
  NOR3_X1   g0079(.A1(new_n279), .A2(new_n259), .A3(G20), .ZN(new_n280));
  NAND2_X1  g0080(.A1(KEYINPUT3), .A2(G33), .ZN(new_n281));
  NAND3_X1  g0081(.A1(new_n267), .A2(new_n210), .A3(new_n281), .ZN(new_n282));
  AOI22_X1  g0082(.A1(new_n278), .A2(new_n280), .B1(new_n259), .B2(new_n282), .ZN(new_n283));
  OAI21_X1  g0083(.A(new_n274), .B1(new_n283), .B2(new_n224), .ZN(new_n284));
  INV_X1    g0084(.A(KEYINPUT16), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  AOI22_X1  g0086(.A1(new_n211), .A2(G33), .B1(G1), .B2(G13), .ZN(new_n287));
  INV_X1    g0087(.A(new_n287), .ZN(new_n288));
  NAND3_X1  g0088(.A1(new_n275), .A2(new_n286), .A3(new_n288), .ZN(new_n289));
  XNOR2_X1  g0089(.A(KEYINPUT8), .B(G58), .ZN(new_n290));
  INV_X1    g0090(.A(new_n290), .ZN(new_n291));
  NAND3_X1  g0091(.A1(new_n209), .A2(G13), .A3(G20), .ZN(new_n292));
  INV_X1    g0092(.A(new_n292), .ZN(new_n293));
  NOR2_X1   g0093(.A1(new_n291), .A2(new_n293), .ZN(new_n294));
  NOR2_X1   g0094(.A1(new_n210), .A2(G1), .ZN(new_n295));
  INV_X1    g0095(.A(new_n295), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n287), .A2(new_n296), .ZN(new_n297));
  AOI21_X1  g0097(.A(new_n294), .B1(new_n297), .B2(new_n291), .ZN(new_n298));
  INV_X1    g0098(.A(new_n298), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n289), .A2(new_n299), .ZN(new_n300));
  OAI21_X1  g0100(.A(new_n209), .B1(G41), .B2(G45), .ZN(new_n301));
  INV_X1    g0101(.A(G274), .ZN(new_n302));
  OR2_X1    g0102(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  INV_X1    g0103(.A(G41), .ZN(new_n304));
  OAI211_X1 g0104(.A(G1), .B(G13), .C1(new_n266), .C2(new_n304), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n305), .A2(new_n301), .ZN(new_n306));
  INV_X1    g0106(.A(new_n306), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n307), .A2(G232), .ZN(new_n308));
  NOR2_X1   g0108(.A1(new_n266), .A2(new_n214), .ZN(new_n309));
  NOR2_X1   g0109(.A1(G223), .A2(G1698), .ZN(new_n310));
  AOI21_X1  g0110(.A(new_n310), .B1(new_n265), .B2(new_n267), .ZN(new_n311));
  INV_X1    g0111(.A(G226), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n312), .A2(G1698), .ZN(new_n313));
  AOI21_X1  g0113(.A(new_n309), .B1(new_n311), .B2(new_n313), .ZN(new_n314));
  OAI211_X1 g0114(.A(new_n303), .B(new_n308), .C1(new_n314), .C2(new_n305), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n315), .A2(G169), .ZN(new_n316));
  INV_X1    g0116(.A(G179), .ZN(new_n317));
  OAI21_X1  g0117(.A(new_n316), .B1(new_n317), .B2(new_n315), .ZN(new_n318));
  NAND3_X1  g0118(.A1(new_n300), .A2(new_n318), .A3(KEYINPUT18), .ZN(new_n319));
  INV_X1    g0119(.A(KEYINPUT73), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  NAND4_X1  g0121(.A1(new_n300), .A2(new_n318), .A3(KEYINPUT73), .A4(KEYINPUT18), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n300), .A2(new_n318), .ZN(new_n323));
  INV_X1    g0123(.A(KEYINPUT18), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n323), .A2(new_n324), .ZN(new_n325));
  AND3_X1   g0125(.A1(new_n321), .A2(new_n322), .A3(new_n325), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n315), .A2(G200), .ZN(new_n327));
  AND3_X1   g0127(.A1(new_n289), .A2(new_n299), .A3(new_n327), .ZN(new_n328));
  XOR2_X1   g0128(.A(KEYINPUT74), .B(G190), .Z(new_n329));
  INV_X1    g0129(.A(new_n329), .ZN(new_n330));
  OR2_X1    g0130(.A1(new_n315), .A2(new_n330), .ZN(new_n331));
  NAND4_X1  g0131(.A1(new_n328), .A2(KEYINPUT75), .A3(KEYINPUT17), .A4(new_n331), .ZN(new_n332));
  INV_X1    g0132(.A(KEYINPUT17), .ZN(new_n333));
  NAND4_X1  g0133(.A1(new_n331), .A2(new_n289), .A3(new_n299), .A4(new_n327), .ZN(new_n334));
  INV_X1    g0134(.A(KEYINPUT75), .ZN(new_n335));
  OAI21_X1  g0135(.A(new_n333), .B1(new_n334), .B2(new_n335), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n332), .A2(new_n336), .ZN(new_n337));
  NOR2_X1   g0137(.A1(new_n326), .A2(new_n337), .ZN(new_n338));
  NOR2_X1   g0138(.A1(new_n279), .A2(new_n256), .ZN(new_n339));
  AOI21_X1  g0139(.A(new_n339), .B1(new_n221), .B2(G1698), .ZN(new_n340));
  INV_X1    g0140(.A(G1698), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n312), .A2(new_n341), .ZN(new_n342));
  AOI22_X1  g0142(.A1(new_n340), .A2(new_n342), .B1(G33), .B2(G97), .ZN(new_n343));
  OAI221_X1 g0143(.A(new_n303), .B1(new_n225), .B2(new_n306), .C1(new_n343), .C2(new_n305), .ZN(new_n344));
  INV_X1    g0144(.A(KEYINPUT13), .ZN(new_n345));
  XNOR2_X1  g0145(.A(new_n344), .B(new_n345), .ZN(new_n346));
  INV_X1    g0146(.A(G169), .ZN(new_n347));
  OAI21_X1  g0147(.A(KEYINPUT14), .B1(new_n346), .B2(new_n347), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n346), .A2(G179), .ZN(new_n349));
  XNOR2_X1  g0149(.A(new_n344), .B(KEYINPUT13), .ZN(new_n350));
  INV_X1    g0150(.A(KEYINPUT14), .ZN(new_n351));
  NAND3_X1  g0151(.A1(new_n350), .A2(new_n351), .A3(G169), .ZN(new_n352));
  NAND3_X1  g0152(.A1(new_n348), .A2(new_n349), .A3(new_n352), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n210), .A2(G33), .ZN(new_n354));
  INV_X1    g0154(.A(G77), .ZN(new_n355));
  OAI22_X1  g0155(.A1(new_n354), .A2(new_n355), .B1(new_n210), .B2(G68), .ZN(new_n356));
  XNOR2_X1  g0156(.A(new_n356), .B(KEYINPUT71), .ZN(new_n357));
  INV_X1    g0157(.A(new_n273), .ZN(new_n358));
  NOR2_X1   g0158(.A1(new_n358), .A2(new_n202), .ZN(new_n359));
  OAI21_X1  g0159(.A(new_n288), .B1(new_n357), .B2(new_n359), .ZN(new_n360));
  XOR2_X1   g0160(.A(new_n360), .B(KEYINPUT11), .Z(new_n361));
  INV_X1    g0161(.A(KEYINPUT12), .ZN(new_n362));
  AOI21_X1  g0162(.A(new_n362), .B1(new_n293), .B2(new_n224), .ZN(new_n363));
  NOR3_X1   g0163(.A1(new_n292), .A2(KEYINPUT12), .A3(G68), .ZN(new_n364));
  OAI22_X1  g0164(.A1(new_n297), .A2(new_n224), .B1(new_n363), .B2(new_n364), .ZN(new_n365));
  NOR2_X1   g0165(.A1(new_n361), .A2(new_n365), .ZN(new_n366));
  INV_X1    g0166(.A(new_n366), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n353), .A2(new_n367), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n350), .A2(G200), .ZN(new_n369));
  AND2_X1   g0169(.A1(new_n369), .A2(new_n366), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n346), .A2(G190), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  NOR2_X1   g0172(.A1(new_n297), .A2(new_n355), .ZN(new_n373));
  AOI22_X1  g0173(.A1(new_n291), .A2(new_n273), .B1(G20), .B2(G77), .ZN(new_n374));
  XOR2_X1   g0174(.A(KEYINPUT15), .B(G87), .Z(new_n375));
  INV_X1    g0175(.A(new_n375), .ZN(new_n376));
  OAI21_X1  g0176(.A(new_n374), .B1(new_n354), .B2(new_n376), .ZN(new_n377));
  AOI21_X1  g0177(.A(new_n373), .B1(new_n377), .B2(new_n288), .ZN(new_n378));
  OAI21_X1  g0178(.A(new_n378), .B1(G77), .B2(new_n292), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n267), .A2(new_n281), .ZN(new_n380));
  NAND3_X1  g0180(.A1(new_n380), .A2(G232), .A3(new_n341), .ZN(new_n381));
  NAND3_X1  g0181(.A1(new_n380), .A2(G238), .A3(G1698), .ZN(new_n382));
  OAI211_X1 g0182(.A(new_n381), .B(new_n382), .C1(new_n206), .C2(new_n380), .ZN(new_n383));
  INV_X1    g0183(.A(new_n305), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n307), .A2(G244), .ZN(new_n386));
  NAND3_X1  g0186(.A1(new_n385), .A2(new_n303), .A3(new_n386), .ZN(new_n387));
  AOI21_X1  g0187(.A(new_n379), .B1(G200), .B2(new_n387), .ZN(new_n388));
  INV_X1    g0188(.A(G190), .ZN(new_n389));
  OAI21_X1  g0189(.A(new_n388), .B1(new_n389), .B2(new_n387), .ZN(new_n390));
  NAND4_X1  g0190(.A1(new_n338), .A2(new_n368), .A3(new_n372), .A4(new_n390), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n293), .A2(new_n202), .ZN(new_n392));
  OR3_X1    g0192(.A1(new_n295), .A2(KEYINPUT67), .A3(new_n202), .ZN(new_n393));
  OAI21_X1  g0193(.A(KEYINPUT67), .B1(new_n295), .B2(new_n202), .ZN(new_n394));
  NAND4_X1  g0194(.A1(new_n393), .A2(new_n287), .A3(new_n292), .A4(new_n394), .ZN(new_n395));
  INV_X1    g0195(.A(G150), .ZN(new_n396));
  OAI22_X1  g0196(.A1(new_n290), .A2(new_n354), .B1(new_n396), .B2(new_n358), .ZN(new_n397));
  AOI21_X1  g0197(.A(new_n397), .B1(G20), .B2(new_n203), .ZN(new_n398));
  OAI211_X1 g0198(.A(new_n392), .B(new_n395), .C1(new_n398), .C2(new_n287), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n339), .A2(new_n355), .ZN(new_n400));
  MUX2_X1   g0200(.A(G222), .B(G223), .S(G1698), .Z(new_n401));
  OAI211_X1 g0201(.A(new_n400), .B(new_n384), .C1(new_n339), .C2(new_n401), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n307), .A2(G226), .ZN(new_n403));
  NAND3_X1  g0203(.A1(new_n402), .A2(new_n403), .A3(new_n303), .ZN(new_n404));
  INV_X1    g0204(.A(new_n404), .ZN(new_n405));
  OAI21_X1  g0205(.A(new_n399), .B1(new_n405), .B2(G169), .ZN(new_n406));
  XNOR2_X1  g0206(.A(new_n406), .B(KEYINPUT68), .ZN(new_n407));
  OAI21_X1  g0207(.A(new_n407), .B1(G179), .B2(new_n404), .ZN(new_n408));
  XNOR2_X1  g0208(.A(new_n399), .B(KEYINPUT69), .ZN(new_n409));
  XNOR2_X1  g0209(.A(new_n409), .B(KEYINPUT9), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n405), .A2(G190), .ZN(new_n411));
  XNOR2_X1  g0211(.A(new_n411), .B(KEYINPUT70), .ZN(new_n412));
  AOI21_X1  g0212(.A(new_n412), .B1(G200), .B2(new_n404), .ZN(new_n413));
  INV_X1    g0213(.A(KEYINPUT10), .ZN(new_n414));
  NAND3_X1  g0214(.A1(new_n410), .A2(new_n413), .A3(new_n414), .ZN(new_n415));
  INV_X1    g0215(.A(new_n415), .ZN(new_n416));
  AOI21_X1  g0216(.A(new_n414), .B1(new_n410), .B2(new_n413), .ZN(new_n417));
  OAI21_X1  g0217(.A(new_n408), .B1(new_n416), .B2(new_n417), .ZN(new_n418));
  INV_X1    g0218(.A(new_n387), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n419), .A2(new_n317), .ZN(new_n420));
  OAI211_X1 g0220(.A(new_n420), .B(new_n379), .C1(G169), .C2(new_n419), .ZN(new_n421));
  INV_X1    g0221(.A(new_n421), .ZN(new_n422));
  NOR3_X1   g0222(.A1(new_n391), .A2(new_n418), .A3(new_n422), .ZN(new_n423));
  INV_X1    g0223(.A(KEYINPUT83), .ZN(new_n424));
  INV_X1    g0224(.A(KEYINPUT22), .ZN(new_n425));
  NAND3_X1  g0225(.A1(new_n425), .A2(new_n210), .A3(G87), .ZN(new_n426));
  OAI21_X1  g0226(.A(new_n424), .B1(new_n339), .B2(new_n426), .ZN(new_n427));
  INV_X1    g0227(.A(new_n426), .ZN(new_n428));
  NAND3_X1  g0228(.A1(new_n428), .A2(new_n380), .A3(KEYINPUT83), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n427), .A2(new_n429), .ZN(new_n430));
  INV_X1    g0230(.A(new_n430), .ZN(new_n431));
  NOR3_X1   g0231(.A1(new_n258), .A2(G20), .A3(new_n214), .ZN(new_n432));
  OAI21_X1  g0232(.A(new_n431), .B1(new_n432), .B2(new_n425), .ZN(new_n433));
  INV_X1    g0233(.A(KEYINPUT24), .ZN(new_n434));
  NOR2_X1   g0234(.A1(new_n210), .A2(G107), .ZN(new_n435));
  XNOR2_X1  g0235(.A(new_n435), .B(KEYINPUT23), .ZN(new_n436));
  NOR2_X1   g0236(.A1(new_n266), .A2(new_n216), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n437), .A2(new_n210), .ZN(new_n438));
  NAND4_X1  g0238(.A1(new_n433), .A2(new_n434), .A3(new_n436), .A4(new_n438), .ZN(new_n439));
  AOI21_X1  g0239(.A(G20), .B1(new_n265), .B2(new_n267), .ZN(new_n440));
  AOI21_X1  g0240(.A(new_n425), .B1(new_n440), .B2(G87), .ZN(new_n441));
  OAI211_X1 g0241(.A(new_n436), .B(new_n438), .C1(new_n441), .C2(new_n430), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n442), .A2(KEYINPUT24), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n439), .A2(new_n443), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n444), .A2(new_n288), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n211), .A2(G33), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n209), .A2(G33), .ZN(new_n447));
  NAND4_X1  g0247(.A1(new_n446), .A2(new_n233), .A3(new_n292), .A4(new_n447), .ZN(new_n448));
  INV_X1    g0248(.A(new_n448), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n449), .A2(G107), .ZN(new_n450));
  NOR2_X1   g0250(.A1(new_n292), .A2(G107), .ZN(new_n451));
  XNOR2_X1  g0251(.A(new_n451), .B(KEYINPUT25), .ZN(new_n452));
  NAND3_X1  g0252(.A1(new_n445), .A2(new_n450), .A3(new_n452), .ZN(new_n453));
  OAI211_X1 g0253(.A(new_n209), .B(G45), .C1(new_n304), .C2(KEYINPUT5), .ZN(new_n454));
  INV_X1    g0254(.A(KEYINPUT5), .ZN(new_n455));
  NOR2_X1   g0255(.A1(new_n455), .A2(G41), .ZN(new_n456));
  OAI21_X1  g0256(.A(new_n305), .B1(new_n454), .B2(new_n456), .ZN(new_n457));
  INV_X1    g0257(.A(new_n457), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n458), .A2(G264), .ZN(new_n459));
  INV_X1    g0259(.A(new_n456), .ZN(new_n460));
  INV_X1    g0260(.A(KEYINPUT78), .ZN(new_n461));
  OAI211_X1 g0261(.A(new_n305), .B(new_n460), .C1(new_n454), .C2(new_n461), .ZN(new_n462));
  INV_X1    g0262(.A(new_n462), .ZN(new_n463));
  AOI21_X1  g0263(.A(new_n302), .B1(new_n454), .B2(new_n461), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  AOI22_X1  g0265(.A1(new_n265), .A2(new_n267), .B1(new_n215), .B2(new_n341), .ZN(new_n466));
  INV_X1    g0266(.A(G257), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n467), .A2(G1698), .ZN(new_n468));
  AOI22_X1  g0268(.A1(new_n466), .A2(new_n468), .B1(G33), .B2(G294), .ZN(new_n469));
  OAI211_X1 g0269(.A(new_n459), .B(new_n465), .C1(new_n469), .C2(new_n305), .ZN(new_n470));
  INV_X1    g0270(.A(new_n470), .ZN(new_n471));
  NOR2_X1   g0271(.A1(new_n471), .A2(G169), .ZN(new_n472));
  INV_X1    g0272(.A(new_n472), .ZN(new_n473));
  NOR2_X1   g0273(.A1(new_n470), .A2(G179), .ZN(new_n474));
  INV_X1    g0274(.A(new_n474), .ZN(new_n475));
  NAND3_X1  g0275(.A1(new_n453), .A2(new_n473), .A3(new_n475), .ZN(new_n476));
  NOR2_X1   g0276(.A1(new_n375), .A2(new_n292), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n440), .A2(G68), .ZN(new_n478));
  NAND3_X1  g0278(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n479), .A2(new_n210), .ZN(new_n480));
  NAND3_X1  g0280(.A1(new_n214), .A2(new_n205), .A3(new_n206), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  INV_X1    g0282(.A(KEYINPUT19), .ZN(new_n483));
  OAI21_X1  g0283(.A(new_n483), .B1(new_n354), .B2(new_n205), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n482), .A2(new_n484), .ZN(new_n485));
  INV_X1    g0285(.A(new_n485), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n478), .A2(new_n486), .ZN(new_n487));
  AOI21_X1  g0287(.A(new_n477), .B1(new_n487), .B2(new_n288), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n449), .A2(new_n375), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n209), .A2(G45), .ZN(new_n490));
  NOR2_X1   g0290(.A1(new_n490), .A2(new_n302), .ZN(new_n491));
  INV_X1    g0291(.A(new_n491), .ZN(new_n492));
  NAND3_X1  g0292(.A1(new_n305), .A2(G250), .A3(new_n490), .ZN(new_n493));
  NOR2_X1   g0293(.A1(new_n341), .A2(G244), .ZN(new_n494));
  AOI21_X1  g0294(.A(new_n494), .B1(new_n265), .B2(new_n267), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n225), .A2(new_n341), .ZN(new_n496));
  AOI21_X1  g0296(.A(new_n437), .B1(new_n495), .B2(new_n496), .ZN(new_n497));
  OAI211_X1 g0297(.A(new_n492), .B(new_n493), .C1(new_n497), .C2(new_n305), .ZN(new_n498));
  AOI22_X1  g0298(.A1(new_n488), .A2(new_n489), .B1(new_n498), .B2(new_n347), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n265), .A2(new_n267), .ZN(new_n500));
  INV_X1    g0300(.A(new_n494), .ZN(new_n501));
  NAND3_X1  g0301(.A1(new_n500), .A2(new_n496), .A3(new_n501), .ZN(new_n502));
  INV_X1    g0302(.A(new_n437), .ZN(new_n503));
  AOI21_X1  g0303(.A(new_n305), .B1(new_n502), .B2(new_n503), .ZN(new_n504));
  INV_X1    g0304(.A(new_n504), .ZN(new_n505));
  NAND4_X1  g0305(.A1(new_n505), .A2(new_n317), .A3(new_n492), .A4(new_n493), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n449), .A2(G87), .ZN(new_n507));
  INV_X1    g0307(.A(new_n477), .ZN(new_n508));
  AOI21_X1  g0308(.A(new_n485), .B1(new_n440), .B2(G68), .ZN(new_n509));
  OAI211_X1 g0309(.A(new_n507), .B(new_n508), .C1(new_n509), .C2(new_n287), .ZN(new_n510));
  AOI21_X1  g0310(.A(new_n510), .B1(G200), .B2(new_n498), .ZN(new_n511));
  INV_X1    g0311(.A(new_n498), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n512), .A2(G190), .ZN(new_n513));
  AOI22_X1  g0313(.A1(new_n499), .A2(new_n506), .B1(new_n511), .B2(new_n513), .ZN(new_n514));
  AND2_X1   g0314(.A1(new_n476), .A2(new_n514), .ZN(new_n515));
  INV_X1    g0315(.A(G200), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n470), .A2(new_n516), .ZN(new_n517));
  OAI21_X1  g0317(.A(new_n517), .B1(G190), .B2(new_n470), .ZN(new_n518));
  NAND4_X1  g0318(.A1(new_n445), .A2(new_n450), .A3(new_n452), .A4(new_n518), .ZN(new_n519));
  NOR2_X1   g0319(.A1(new_n292), .A2(G97), .ZN(new_n520));
  INV_X1    g0320(.A(new_n520), .ZN(new_n521));
  OAI21_X1  g0321(.A(new_n521), .B1(new_n448), .B2(new_n205), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n273), .A2(G77), .ZN(new_n523));
  INV_X1    g0323(.A(KEYINPUT76), .ZN(new_n524));
  NAND2_X1  g0324(.A1(KEYINPUT6), .A2(G97), .ZN(new_n525));
  OAI21_X1  g0325(.A(new_n524), .B1(new_n525), .B2(G107), .ZN(new_n526));
  NAND4_X1  g0326(.A1(new_n206), .A2(KEYINPUT76), .A3(KEYINPUT6), .A4(G97), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  NAND2_X1  g0328(.A1(G97), .A2(G107), .ZN(new_n529));
  AOI21_X1  g0329(.A(KEYINPUT6), .B1(new_n207), .B2(new_n529), .ZN(new_n530));
  OAI21_X1  g0330(.A(G20), .B1(new_n528), .B2(new_n530), .ZN(new_n531));
  OAI211_X1 g0331(.A(new_n523), .B(new_n531), .C1(new_n283), .C2(new_n206), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n532), .A2(new_n288), .ZN(new_n533));
  INV_X1    g0333(.A(KEYINPUT77), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  NAND3_X1  g0335(.A1(new_n532), .A2(KEYINPUT77), .A3(new_n288), .ZN(new_n536));
  AOI21_X1  g0336(.A(new_n522), .B1(new_n535), .B2(new_n536), .ZN(new_n537));
  INV_X1    g0337(.A(new_n464), .ZN(new_n538));
  OAI22_X1  g0338(.A1(new_n538), .A2(new_n462), .B1(new_n467), .B2(new_n457), .ZN(new_n539));
  OAI211_X1 g0339(.A(G250), .B(G1698), .C1(new_n279), .C2(new_n256), .ZN(new_n540));
  AND2_X1   g0340(.A1(KEYINPUT4), .A2(G244), .ZN(new_n541));
  OAI211_X1 g0341(.A(new_n341), .B(new_n541), .C1(new_n279), .C2(new_n256), .ZN(new_n542));
  NAND2_X1  g0342(.A1(G33), .A2(G283), .ZN(new_n543));
  NAND3_X1  g0343(.A1(new_n540), .A2(new_n542), .A3(new_n543), .ZN(new_n544));
  INV_X1    g0344(.A(new_n544), .ZN(new_n545));
  INV_X1    g0345(.A(G244), .ZN(new_n546));
  AOI211_X1 g0346(.A(new_n546), .B(G1698), .C1(new_n265), .C2(new_n267), .ZN(new_n547));
  OAI21_X1  g0347(.A(new_n545), .B1(new_n547), .B2(KEYINPUT4), .ZN(new_n548));
  AOI21_X1  g0348(.A(new_n539), .B1(new_n548), .B2(new_n384), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n549), .A2(G190), .ZN(new_n550));
  OAI211_X1 g0350(.A(new_n537), .B(new_n550), .C1(new_n516), .C2(new_n549), .ZN(new_n551));
  AOI21_X1  g0351(.A(G1698), .B1(new_n265), .B2(new_n267), .ZN(new_n552));
  AOI21_X1  g0352(.A(KEYINPUT4), .B1(new_n552), .B2(G244), .ZN(new_n553));
  OAI21_X1  g0353(.A(new_n384), .B1(new_n553), .B2(new_n544), .ZN(new_n554));
  INV_X1    g0354(.A(new_n539), .ZN(new_n555));
  NAND3_X1  g0355(.A1(new_n554), .A2(new_n317), .A3(new_n555), .ZN(new_n556));
  OAI21_X1  g0356(.A(new_n556), .B1(new_n549), .B2(G169), .ZN(new_n557));
  NOR3_X1   g0357(.A1(new_n537), .A2(new_n557), .A3(KEYINPUT79), .ZN(new_n558));
  INV_X1    g0358(.A(KEYINPUT79), .ZN(new_n559));
  AOI211_X1 g0359(.A(G179), .B(new_n539), .C1(new_n548), .C2(new_n384), .ZN(new_n560));
  AOI21_X1  g0360(.A(G169), .B1(new_n554), .B2(new_n555), .ZN(new_n561));
  NOR2_X1   g0361(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  INV_X1    g0362(.A(new_n522), .ZN(new_n563));
  AND3_X1   g0363(.A1(new_n532), .A2(KEYINPUT77), .A3(new_n288), .ZN(new_n564));
  AOI21_X1  g0364(.A(KEYINPUT77), .B1(new_n532), .B2(new_n288), .ZN(new_n565));
  OAI21_X1  g0365(.A(new_n563), .B1(new_n564), .B2(new_n565), .ZN(new_n566));
  AOI21_X1  g0366(.A(new_n559), .B1(new_n562), .B2(new_n566), .ZN(new_n567));
  OAI211_X1 g0367(.A(new_n519), .B(new_n551), .C1(new_n558), .C2(new_n567), .ZN(new_n568));
  INV_X1    g0368(.A(new_n568), .ZN(new_n569));
  INV_X1    g0369(.A(KEYINPUT80), .ZN(new_n570));
  NAND2_X1  g0370(.A1(G264), .A2(G1698), .ZN(new_n571));
  OAI21_X1  g0371(.A(new_n570), .B1(new_n258), .B2(new_n571), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n339), .A2(G303), .ZN(new_n573));
  NAND3_X1  g0373(.A1(new_n500), .A2(G257), .A3(new_n341), .ZN(new_n574));
  INV_X1    g0374(.A(new_n571), .ZN(new_n575));
  NAND3_X1  g0375(.A1(new_n500), .A2(KEYINPUT80), .A3(new_n575), .ZN(new_n576));
  NAND4_X1  g0376(.A1(new_n572), .A2(new_n573), .A3(new_n574), .A4(new_n576), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n577), .A2(new_n384), .ZN(new_n578));
  OAI22_X1  g0378(.A1(new_n538), .A2(new_n462), .B1(new_n217), .B2(new_n457), .ZN(new_n579));
  INV_X1    g0379(.A(new_n579), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n578), .A2(new_n580), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n293), .A2(new_n216), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n449), .A2(G116), .ZN(new_n583));
  AOI22_X1  g0383(.A1(new_n446), .A2(new_n233), .B1(G20), .B2(new_n216), .ZN(new_n584));
  OAI211_X1 g0384(.A(new_n543), .B(new_n210), .C1(G33), .C2(new_n205), .ZN(new_n585));
  AND3_X1   g0385(.A1(new_n584), .A2(KEYINPUT20), .A3(new_n585), .ZN(new_n586));
  AOI21_X1  g0386(.A(KEYINPUT20), .B1(new_n584), .B2(new_n585), .ZN(new_n587));
  OAI211_X1 g0387(.A(new_n582), .B(new_n583), .C1(new_n586), .C2(new_n587), .ZN(new_n588));
  NAND3_X1  g0388(.A1(new_n581), .A2(G169), .A3(new_n588), .ZN(new_n589));
  INV_X1    g0389(.A(KEYINPUT21), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  INV_X1    g0391(.A(new_n588), .ZN(new_n592));
  AOI21_X1  g0392(.A(new_n579), .B1(new_n577), .B2(new_n384), .ZN(new_n593));
  OAI21_X1  g0393(.A(new_n592), .B1(new_n593), .B2(new_n516), .ZN(new_n594));
  INV_X1    g0394(.A(KEYINPUT82), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n593), .A2(new_n329), .ZN(new_n597));
  OAI211_X1 g0397(.A(new_n592), .B(KEYINPUT82), .C1(new_n593), .C2(new_n516), .ZN(new_n598));
  NAND3_X1  g0398(.A1(new_n596), .A2(new_n597), .A3(new_n598), .ZN(new_n599));
  INV_X1    g0399(.A(KEYINPUT81), .ZN(new_n600));
  AOI21_X1  g0400(.A(KEYINPUT80), .B1(new_n500), .B2(new_n575), .ZN(new_n601));
  AOI211_X1 g0401(.A(new_n570), .B(new_n571), .C1(new_n265), .C2(new_n267), .ZN(new_n602));
  NOR2_X1   g0402(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  AOI22_X1  g0403(.A1(new_n552), .A2(G257), .B1(G303), .B2(new_n339), .ZN(new_n604));
  AOI21_X1  g0404(.A(new_n305), .B1(new_n603), .B2(new_n604), .ZN(new_n605));
  OAI211_X1 g0405(.A(KEYINPUT21), .B(G169), .C1(new_n605), .C2(new_n579), .ZN(new_n606));
  NAND3_X1  g0406(.A1(new_n578), .A2(G179), .A3(new_n580), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  AOI21_X1  g0408(.A(new_n600), .B1(new_n608), .B2(new_n588), .ZN(new_n609));
  AOI211_X1 g0409(.A(KEYINPUT81), .B(new_n592), .C1(new_n606), .C2(new_n607), .ZN(new_n610));
  OAI211_X1 g0410(.A(new_n591), .B(new_n599), .C1(new_n609), .C2(new_n610), .ZN(new_n611));
  INV_X1    g0411(.A(new_n611), .ZN(new_n612));
  AND4_X1   g0412(.A1(new_n423), .A2(new_n515), .A3(new_n569), .A4(new_n612), .ZN(G372));
  INV_X1    g0413(.A(new_n408), .ZN(new_n614));
  AND2_X1   g0414(.A1(new_n325), .A2(new_n319), .ZN(new_n615));
  INV_X1    g0415(.A(new_n615), .ZN(new_n616));
  AOI22_X1  g0416(.A1(new_n353), .A2(new_n367), .B1(new_n372), .B2(new_n422), .ZN(new_n617));
  OAI211_X1 g0417(.A(KEYINPUT85), .B(new_n616), .C1(new_n617), .C2(new_n337), .ZN(new_n618));
  OR2_X1    g0418(.A1(new_n416), .A2(new_n417), .ZN(new_n619));
  AND2_X1   g0419(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  OAI21_X1  g0420(.A(new_n616), .B1(new_n617), .B2(new_n337), .ZN(new_n621));
  INV_X1    g0421(.A(KEYINPUT85), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  AOI21_X1  g0423(.A(new_n614), .B1(new_n620), .B2(new_n623), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n488), .A2(new_n489), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n498), .A2(new_n347), .ZN(new_n626));
  AND3_X1   g0426(.A1(new_n506), .A2(new_n625), .A3(new_n626), .ZN(new_n627));
  NOR2_X1   g0427(.A1(new_n498), .A2(new_n389), .ZN(new_n628));
  INV_X1    g0428(.A(KEYINPUT84), .ZN(new_n629));
  AOI21_X1  g0429(.A(new_n628), .B1(new_n511), .B2(new_n629), .ZN(new_n630));
  INV_X1    g0430(.A(new_n510), .ZN(new_n631));
  OAI21_X1  g0431(.A(new_n631), .B1(new_n512), .B2(new_n516), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n632), .A2(KEYINPUT84), .ZN(new_n633));
  AOI21_X1  g0433(.A(new_n627), .B1(new_n630), .B2(new_n633), .ZN(new_n634));
  INV_X1    g0434(.A(KEYINPUT26), .ZN(new_n635));
  NOR2_X1   g0435(.A1(new_n537), .A2(new_n557), .ZN(new_n636));
  NAND3_X1  g0436(.A1(new_n634), .A2(new_n635), .A3(new_n636), .ZN(new_n637));
  OAI21_X1  g0437(.A(KEYINPUT79), .B1(new_n537), .B2(new_n557), .ZN(new_n638));
  NAND3_X1  g0438(.A1(new_n562), .A2(new_n566), .A3(new_n559), .ZN(new_n639));
  NAND3_X1  g0439(.A1(new_n638), .A2(new_n514), .A3(new_n639), .ZN(new_n640));
  AOI21_X1  g0440(.A(new_n627), .B1(new_n640), .B2(KEYINPUT26), .ZN(new_n641));
  AOI211_X1 g0441(.A(new_n317), .B(new_n579), .C1(new_n577), .C2(new_n384), .ZN(new_n642));
  NOR2_X1   g0442(.A1(new_n593), .A2(new_n347), .ZN(new_n643));
  AOI21_X1  g0443(.A(new_n642), .B1(new_n643), .B2(KEYINPUT21), .ZN(new_n644));
  OAI21_X1  g0444(.A(new_n591), .B1(new_n644), .B2(new_n592), .ZN(new_n645));
  AOI22_X1  g0445(.A1(new_n444), .A2(new_n288), .B1(G107), .B2(new_n449), .ZN(new_n646));
  AOI21_X1  g0446(.A(new_n472), .B1(new_n646), .B2(new_n452), .ZN(new_n647));
  AOI21_X1  g0447(.A(new_n645), .B1(new_n647), .B2(new_n475), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n638), .A2(new_n639), .ZN(new_n649));
  NAND4_X1  g0449(.A1(new_n649), .A2(new_n634), .A3(new_n551), .A4(new_n519), .ZN(new_n650));
  OAI211_X1 g0450(.A(new_n637), .B(new_n641), .C1(new_n648), .C2(new_n650), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n423), .A2(new_n651), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n624), .A2(new_n652), .ZN(G369));
  INV_X1    g0453(.A(G13), .ZN(new_n654));
  NOR2_X1   g0454(.A1(new_n654), .A2(G20), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n655), .A2(new_n209), .ZN(new_n656));
  OR2_X1    g0456(.A1(new_n656), .A2(KEYINPUT27), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n656), .A2(KEYINPUT27), .ZN(new_n658));
  NAND3_X1  g0458(.A1(new_n657), .A2(G213), .A3(new_n658), .ZN(new_n659));
  INV_X1    g0459(.A(G343), .ZN(new_n660));
  NOR2_X1   g0460(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  INV_X1    g0461(.A(new_n661), .ZN(new_n662));
  OAI21_X1  g0462(.A(new_n612), .B1(new_n592), .B2(new_n662), .ZN(new_n663));
  NAND3_X1  g0463(.A1(new_n645), .A2(new_n588), .A3(new_n661), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n664), .A2(KEYINPUT86), .ZN(new_n665));
  OR2_X1    g0465(.A1(new_n664), .A2(KEYINPUT86), .ZN(new_n666));
  NAND3_X1  g0466(.A1(new_n663), .A2(new_n665), .A3(new_n666), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n667), .A2(G330), .ZN(new_n668));
  NOR2_X1   g0468(.A1(new_n476), .A2(new_n661), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n453), .A2(new_n661), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n670), .A2(new_n519), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n671), .A2(new_n476), .ZN(new_n672));
  INV_X1    g0472(.A(new_n672), .ZN(new_n673));
  NOR3_X1   g0473(.A1(new_n668), .A2(new_n669), .A3(new_n673), .ZN(new_n674));
  INV_X1    g0474(.A(new_n674), .ZN(new_n675));
  OAI21_X1  g0475(.A(new_n591), .B1(new_n609), .B2(new_n610), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n676), .A2(new_n662), .ZN(new_n677));
  INV_X1    g0477(.A(new_n677), .ZN(new_n678));
  AOI21_X1  g0478(.A(new_n669), .B1(new_n678), .B2(new_n672), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n675), .A2(new_n679), .ZN(G399));
  NAND2_X1  g0480(.A1(new_n230), .A2(new_n304), .ZN(new_n681));
  NOR2_X1   g0481(.A1(new_n481), .A2(G116), .ZN(new_n682));
  NAND3_X1  g0482(.A1(new_n681), .A2(G1), .A3(new_n682), .ZN(new_n683));
  OAI21_X1  g0483(.A(new_n683), .B1(new_n235), .B2(new_n681), .ZN(new_n684));
  XNOR2_X1  g0484(.A(new_n684), .B(KEYINPUT28), .ZN(new_n685));
  INV_X1    g0485(.A(KEYINPUT29), .ZN(new_n686));
  INV_X1    g0486(.A(KEYINPUT88), .ZN(new_n687));
  AND3_X1   g0487(.A1(new_n651), .A2(new_n687), .A3(new_n662), .ZN(new_n688));
  AOI21_X1  g0488(.A(new_n687), .B1(new_n651), .B2(new_n662), .ZN(new_n689));
  OAI21_X1  g0489(.A(new_n686), .B1(new_n688), .B2(new_n689), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n690), .A2(KEYINPUT89), .ZN(new_n691));
  AOI211_X1 g0491(.A(new_n472), .B(new_n474), .C1(new_n646), .C2(new_n452), .ZN(new_n692));
  NOR2_X1   g0492(.A1(new_n676), .A2(new_n692), .ZN(new_n693));
  OAI21_X1  g0493(.A(KEYINPUT90), .B1(new_n693), .B2(new_n650), .ZN(new_n694));
  OR2_X1    g0494(.A1(new_n640), .A2(KEYINPUT26), .ZN(new_n695));
  OAI211_X1 g0495(.A(new_n476), .B(new_n591), .C1(new_n609), .C2(new_n610), .ZN(new_n696));
  INV_X1    g0496(.A(KEYINPUT90), .ZN(new_n697));
  NAND4_X1  g0497(.A1(new_n696), .A2(new_n569), .A3(new_n697), .A4(new_n634), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n634), .A2(new_n636), .ZN(new_n699));
  AOI21_X1  g0499(.A(new_n627), .B1(new_n699), .B2(KEYINPUT26), .ZN(new_n700));
  NAND4_X1  g0500(.A1(new_n694), .A2(new_n695), .A3(new_n698), .A4(new_n700), .ZN(new_n701));
  NAND3_X1  g0501(.A1(new_n701), .A2(KEYINPUT29), .A3(new_n662), .ZN(new_n702));
  INV_X1    g0502(.A(KEYINPUT89), .ZN(new_n703));
  OAI211_X1 g0503(.A(new_n703), .B(new_n686), .C1(new_n688), .C2(new_n689), .ZN(new_n704));
  NAND3_X1  g0504(.A1(new_n691), .A2(new_n702), .A3(new_n704), .ZN(new_n705));
  NAND4_X1  g0505(.A1(new_n612), .A2(new_n515), .A3(new_n569), .A4(new_n662), .ZN(new_n706));
  OAI21_X1  g0506(.A(new_n459), .B1(new_n469), .B2(new_n305), .ZN(new_n707));
  NOR2_X1   g0507(.A1(new_n707), .A2(new_n498), .ZN(new_n708));
  NAND3_X1  g0508(.A1(new_n642), .A2(new_n549), .A3(new_n708), .ZN(new_n709));
  INV_X1    g0509(.A(KEYINPUT30), .ZN(new_n710));
  AND2_X1   g0510(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  NOR2_X1   g0511(.A1(new_n549), .A2(G179), .ZN(new_n712));
  NAND4_X1  g0512(.A1(new_n712), .A2(new_n498), .A3(new_n470), .A4(new_n581), .ZN(new_n713));
  NAND4_X1  g0513(.A1(new_n642), .A2(new_n708), .A3(KEYINPUT30), .A4(new_n549), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  OAI211_X1 g0515(.A(KEYINPUT31), .B(new_n661), .C1(new_n711), .C2(new_n715), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n466), .A2(new_n468), .ZN(new_n717));
  NAND2_X1  g0517(.A1(G33), .A2(G294), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  AOI22_X1  g0519(.A1(new_n719), .A2(new_n384), .B1(G264), .B2(new_n458), .ZN(new_n720));
  NAND3_X1  g0520(.A1(new_n512), .A2(new_n549), .A3(new_n720), .ZN(new_n721));
  OAI211_X1 g0521(.A(KEYINPUT87), .B(new_n710), .C1(new_n721), .C2(new_n607), .ZN(new_n722));
  NAND3_X1  g0522(.A1(new_n722), .A2(new_n714), .A3(new_n713), .ZN(new_n723));
  AOI21_X1  g0523(.A(KEYINPUT87), .B1(new_n709), .B2(new_n710), .ZN(new_n724));
  OAI21_X1  g0524(.A(new_n661), .B1(new_n723), .B2(new_n724), .ZN(new_n725));
  INV_X1    g0525(.A(KEYINPUT31), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  NAND3_X1  g0527(.A1(new_n706), .A2(new_n716), .A3(new_n727), .ZN(new_n728));
  NAND2_X1  g0528(.A1(new_n728), .A2(G330), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n705), .A2(new_n729), .ZN(new_n730));
  NAND2_X1  g0530(.A1(new_n730), .A2(KEYINPUT91), .ZN(new_n731));
  INV_X1    g0531(.A(KEYINPUT91), .ZN(new_n732));
  NAND3_X1  g0532(.A1(new_n705), .A2(new_n732), .A3(new_n729), .ZN(new_n733));
  NAND2_X1  g0533(.A1(new_n731), .A2(new_n733), .ZN(new_n734));
  OAI21_X1  g0534(.A(new_n685), .B1(new_n734), .B2(G1), .ZN(G364));
  INV_X1    g0535(.A(new_n667), .ZN(new_n736));
  NOR2_X1   g0536(.A1(G13), .A2(G33), .ZN(new_n737));
  INV_X1    g0537(.A(new_n737), .ZN(new_n738));
  NOR2_X1   g0538(.A1(new_n738), .A2(G20), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n736), .A2(new_n739), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n655), .A2(G45), .ZN(new_n741));
  NAND3_X1  g0541(.A1(new_n681), .A2(G1), .A3(new_n741), .ZN(new_n742));
  INV_X1    g0542(.A(new_n742), .ZN(new_n743));
  NAND2_X1  g0543(.A1(new_n258), .A2(new_n230), .ZN(new_n744));
  INV_X1    g0544(.A(new_n744), .ZN(new_n745));
  INV_X1    g0545(.A(G45), .ZN(new_n746));
  NAND2_X1  g0546(.A1(new_n236), .A2(new_n746), .ZN(new_n747));
  OAI211_X1 g0547(.A(new_n745), .B(new_n747), .C1(new_n254), .C2(new_n746), .ZN(new_n748));
  NAND3_X1  g0548(.A1(new_n230), .A2(G355), .A3(new_n380), .ZN(new_n749));
  OAI211_X1 g0549(.A(new_n748), .B(new_n749), .C1(G116), .C2(new_n230), .ZN(new_n750));
  AOI21_X1  g0550(.A(new_n233), .B1(G20), .B2(new_n347), .ZN(new_n751));
  NOR2_X1   g0551(.A1(new_n739), .A2(new_n751), .ZN(new_n752));
  NAND2_X1  g0552(.A1(new_n750), .A2(new_n752), .ZN(new_n753));
  NAND2_X1  g0553(.A1(G20), .A2(G179), .ZN(new_n754));
  XNOR2_X1  g0554(.A(new_n754), .B(KEYINPUT92), .ZN(new_n755));
  NAND3_X1  g0555(.A1(new_n755), .A2(new_n329), .A3(new_n516), .ZN(new_n756));
  INV_X1    g0556(.A(new_n756), .ZN(new_n757));
  AOI21_X1  g0557(.A(new_n380), .B1(new_n757), .B2(G322), .ZN(new_n758));
  NOR2_X1   g0558(.A1(new_n210), .A2(G179), .ZN(new_n759));
  NAND3_X1  g0559(.A1(new_n759), .A2(new_n389), .A3(G200), .ZN(new_n760));
  INV_X1    g0560(.A(G283), .ZN(new_n761));
  NAND3_X1  g0561(.A1(new_n759), .A2(G190), .A3(G200), .ZN(new_n762));
  INV_X1    g0562(.A(G303), .ZN(new_n763));
  OAI22_X1  g0563(.A1(new_n760), .A2(new_n761), .B1(new_n762), .B2(new_n763), .ZN(new_n764));
  NOR2_X1   g0564(.A1(G190), .A2(G200), .ZN(new_n765));
  NAND2_X1  g0565(.A1(new_n755), .A2(new_n765), .ZN(new_n766));
  INV_X1    g0566(.A(new_n766), .ZN(new_n767));
  AOI21_X1  g0567(.A(new_n764), .B1(new_n767), .B2(G311), .ZN(new_n768));
  NAND3_X1  g0568(.A1(new_n755), .A2(new_n389), .A3(G200), .ZN(new_n769));
  XOR2_X1   g0569(.A(KEYINPUT33), .B(G317), .Z(new_n770));
  OAI211_X1 g0570(.A(new_n758), .B(new_n768), .C1(new_n769), .C2(new_n770), .ZN(new_n771));
  NAND2_X1  g0571(.A1(new_n759), .A2(new_n765), .ZN(new_n772));
  INV_X1    g0572(.A(new_n772), .ZN(new_n773));
  NAND2_X1  g0573(.A1(new_n773), .A2(G329), .ZN(new_n774));
  NAND3_X1  g0574(.A1(new_n755), .A2(new_n329), .A3(G200), .ZN(new_n775));
  XNOR2_X1  g0575(.A(new_n775), .B(KEYINPUT94), .ZN(new_n776));
  INV_X1    g0576(.A(new_n776), .ZN(new_n777));
  INV_X1    g0577(.A(G326), .ZN(new_n778));
  OAI21_X1  g0578(.A(new_n774), .B1(new_n777), .B2(new_n778), .ZN(new_n779));
  NOR3_X1   g0579(.A1(new_n389), .A2(G179), .A3(G200), .ZN(new_n780));
  NOR2_X1   g0580(.A1(new_n780), .A2(new_n210), .ZN(new_n781));
  INV_X1    g0581(.A(new_n781), .ZN(new_n782));
  AOI211_X1 g0582(.A(new_n771), .B(new_n779), .C1(G294), .C2(new_n782), .ZN(new_n783));
  XNOR2_X1  g0583(.A(new_n766), .B(KEYINPUT93), .ZN(new_n784));
  INV_X1    g0584(.A(new_n784), .ZN(new_n785));
  OAI221_X1 g0585(.A(new_n380), .B1(new_n220), .B2(new_n756), .C1(new_n785), .C2(new_n355), .ZN(new_n786));
  INV_X1    g0586(.A(new_n775), .ZN(new_n787));
  INV_X1    g0587(.A(new_n760), .ZN(new_n788));
  AOI22_X1  g0588(.A1(new_n787), .A2(G50), .B1(G107), .B2(new_n788), .ZN(new_n789));
  OAI221_X1 g0589(.A(new_n789), .B1(new_n224), .B2(new_n769), .C1(new_n214), .C2(new_n762), .ZN(new_n790));
  INV_X1    g0590(.A(G159), .ZN(new_n791));
  NOR3_X1   g0591(.A1(new_n772), .A2(KEYINPUT32), .A3(new_n791), .ZN(new_n792));
  OAI21_X1  g0592(.A(KEYINPUT32), .B1(new_n772), .B2(new_n791), .ZN(new_n793));
  OAI21_X1  g0593(.A(new_n793), .B1(new_n205), .B2(new_n781), .ZN(new_n794));
  NOR4_X1   g0594(.A1(new_n786), .A2(new_n790), .A3(new_n792), .A4(new_n794), .ZN(new_n795));
  OAI21_X1  g0595(.A(new_n751), .B1(new_n783), .B2(new_n795), .ZN(new_n796));
  NAND4_X1  g0596(.A1(new_n740), .A2(new_n743), .A3(new_n753), .A4(new_n796), .ZN(new_n797));
  INV_X1    g0597(.A(G330), .ZN(new_n798));
  NAND2_X1  g0598(.A1(new_n736), .A2(new_n798), .ZN(new_n799));
  NAND3_X1  g0599(.A1(new_n799), .A2(new_n668), .A3(new_n742), .ZN(new_n800));
  NAND2_X1  g0600(.A1(new_n797), .A2(new_n800), .ZN(G396));
  NAND2_X1  g0601(.A1(new_n379), .A2(new_n661), .ZN(new_n802));
  AOI21_X1  g0602(.A(new_n422), .B1(new_n390), .B2(new_n802), .ZN(new_n803));
  NOR2_X1   g0603(.A1(new_n421), .A2(new_n661), .ZN(new_n804));
  NOR2_X1   g0604(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  NAND3_X1  g0605(.A1(new_n651), .A2(new_n662), .A3(new_n805), .ZN(new_n806));
  INV_X1    g0606(.A(new_n806), .ZN(new_n807));
  OR2_X1    g0607(.A1(new_n688), .A2(new_n689), .ZN(new_n808));
  INV_X1    g0608(.A(new_n805), .ZN(new_n809));
  AOI21_X1  g0609(.A(new_n807), .B1(new_n808), .B2(new_n809), .ZN(new_n810));
  XNOR2_X1  g0610(.A(new_n810), .B(new_n729), .ZN(new_n811));
  NAND2_X1  g0611(.A1(new_n811), .A2(new_n742), .ZN(new_n812));
  NOR2_X1   g0612(.A1(new_n751), .A2(new_n737), .ZN(new_n813));
  XOR2_X1   g0613(.A(new_n813), .B(KEYINPUT95), .Z(new_n814));
  AOI22_X1  g0614(.A1(new_n809), .A2(new_n737), .B1(new_n355), .B2(new_n814), .ZN(new_n815));
  OAI21_X1  g0615(.A(new_n339), .B1(new_n785), .B2(new_n216), .ZN(new_n816));
  NOR2_X1   g0616(.A1(new_n775), .A2(new_n763), .ZN(new_n817));
  INV_X1    g0617(.A(G294), .ZN(new_n818));
  OAI22_X1  g0618(.A1(new_n761), .A2(new_n769), .B1(new_n756), .B2(new_n818), .ZN(new_n819));
  OAI22_X1  g0619(.A1(new_n760), .A2(new_n214), .B1(new_n762), .B2(new_n206), .ZN(new_n820));
  AOI21_X1  g0620(.A(new_n820), .B1(G311), .B2(new_n773), .ZN(new_n821));
  OAI21_X1  g0621(.A(new_n821), .B1(new_n205), .B2(new_n781), .ZN(new_n822));
  NOR4_X1   g0622(.A1(new_n816), .A2(new_n817), .A3(new_n819), .A4(new_n822), .ZN(new_n823));
  INV_X1    g0623(.A(new_n769), .ZN(new_n824));
  AOI22_X1  g0624(.A1(new_n824), .A2(G150), .B1(new_n757), .B2(G143), .ZN(new_n825));
  INV_X1    g0625(.A(G137), .ZN(new_n826));
  OAI21_X1  g0626(.A(new_n825), .B1(new_n826), .B2(new_n775), .ZN(new_n827));
  AOI21_X1  g0627(.A(new_n827), .B1(G159), .B2(new_n784), .ZN(new_n828));
  XNOR2_X1  g0628(.A(new_n828), .B(KEYINPUT97), .ZN(new_n829));
  XOR2_X1   g0629(.A(KEYINPUT96), .B(KEYINPUT34), .Z(new_n830));
  INV_X1    g0630(.A(new_n830), .ZN(new_n831));
  NAND2_X1  g0631(.A1(new_n829), .A2(new_n831), .ZN(new_n832));
  INV_X1    g0632(.A(G132), .ZN(new_n833));
  OAI21_X1  g0633(.A(new_n832), .B1(new_n833), .B2(new_n772), .ZN(new_n834));
  OAI22_X1  g0634(.A1(new_n829), .A2(new_n831), .B1(new_n220), .B2(new_n781), .ZN(new_n835));
  NOR2_X1   g0635(.A1(new_n760), .A2(new_n224), .ZN(new_n836));
  NOR4_X1   g0636(.A1(new_n834), .A2(new_n835), .A3(new_n258), .A4(new_n836), .ZN(new_n837));
  INV_X1    g0637(.A(new_n762), .ZN(new_n838));
  NAND2_X1  g0638(.A1(new_n838), .A2(G50), .ZN(new_n839));
  AOI21_X1  g0639(.A(new_n823), .B1(new_n837), .B2(new_n839), .ZN(new_n840));
  INV_X1    g0640(.A(new_n751), .ZN(new_n841));
  OAI211_X1 g0641(.A(new_n743), .B(new_n815), .C1(new_n840), .C2(new_n841), .ZN(new_n842));
  NAND2_X1  g0642(.A1(new_n812), .A2(new_n842), .ZN(G384));
  NAND4_X1  g0643(.A1(new_n691), .A2(new_n423), .A3(new_n702), .A4(new_n704), .ZN(new_n844));
  AND2_X1   g0644(.A1(new_n844), .A2(new_n624), .ZN(new_n845));
  NOR2_X1   g0645(.A1(new_n368), .A2(new_n661), .ZN(new_n846));
  INV_X1    g0646(.A(KEYINPUT39), .ZN(new_n847));
  INV_X1    g0647(.A(new_n659), .ZN(new_n848));
  NAND2_X1  g0648(.A1(new_n275), .A2(new_n288), .ZN(new_n849));
  AOI21_X1  g0649(.A(KEYINPUT16), .B1(new_n270), .B2(new_n274), .ZN(new_n850));
  OAI21_X1  g0650(.A(new_n299), .B1(new_n849), .B2(new_n850), .ZN(new_n851));
  OAI211_X1 g0651(.A(new_n848), .B(new_n851), .C1(new_n326), .C2(new_n337), .ZN(new_n852));
  OAI21_X1  g0652(.A(new_n300), .B1(new_n318), .B2(new_n848), .ZN(new_n853));
  INV_X1    g0653(.A(KEYINPUT37), .ZN(new_n854));
  NAND3_X1  g0654(.A1(new_n853), .A2(new_n854), .A3(new_n334), .ZN(new_n855));
  OAI21_X1  g0655(.A(new_n851), .B1(new_n318), .B2(new_n848), .ZN(new_n856));
  AND2_X1   g0656(.A1(new_n856), .A2(new_n334), .ZN(new_n857));
  OAI21_X1  g0657(.A(new_n855), .B1(new_n857), .B2(new_n854), .ZN(new_n858));
  AOI21_X1  g0658(.A(KEYINPUT38), .B1(new_n852), .B2(new_n858), .ZN(new_n859));
  INV_X1    g0659(.A(new_n859), .ZN(new_n860));
  NAND3_X1  g0660(.A1(new_n852), .A2(KEYINPUT38), .A3(new_n858), .ZN(new_n861));
  AOI21_X1  g0661(.A(new_n847), .B1(new_n860), .B2(new_n861), .ZN(new_n862));
  OAI211_X1 g0662(.A(new_n300), .B(new_n848), .C1(new_n615), .C2(new_n337), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n853), .A2(new_n334), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n864), .A2(KEYINPUT37), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n865), .A2(new_n855), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n863), .A2(new_n866), .ZN(new_n867));
  INV_X1    g0667(.A(KEYINPUT38), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  NAND3_X1  g0669(.A1(new_n869), .A2(new_n847), .A3(new_n861), .ZN(new_n870));
  INV_X1    g0670(.A(new_n870), .ZN(new_n871));
  OAI21_X1  g0671(.A(new_n846), .B1(new_n862), .B2(new_n871), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n367), .A2(new_n661), .ZN(new_n873));
  NAND3_X1  g0673(.A1(new_n368), .A2(new_n372), .A3(new_n873), .ZN(new_n874));
  NAND3_X1  g0674(.A1(new_n353), .A2(new_n367), .A3(new_n661), .ZN(new_n875));
  AND2_X1   g0675(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  XNOR2_X1  g0676(.A(new_n804), .B(KEYINPUT98), .ZN(new_n877));
  AOI21_X1  g0677(.A(new_n876), .B1(new_n806), .B2(new_n877), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n860), .A2(new_n861), .ZN(new_n879));
  AOI22_X1  g0679(.A1(new_n878), .A2(new_n879), .B1(new_n615), .B2(new_n659), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n872), .A2(new_n880), .ZN(new_n881));
  XNOR2_X1  g0681(.A(new_n845), .B(new_n881), .ZN(new_n882));
  OAI211_X1 g0682(.A(KEYINPUT31), .B(new_n661), .C1(new_n723), .C2(new_n724), .ZN(new_n883));
  INV_X1    g0683(.A(KEYINPUT99), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n885), .A2(new_n727), .ZN(new_n886));
  NAND3_X1  g0686(.A1(new_n725), .A2(new_n884), .A3(new_n726), .ZN(new_n887));
  NAND3_X1  g0687(.A1(new_n706), .A2(new_n886), .A3(new_n887), .ZN(new_n888));
  AOI21_X1  g0688(.A(new_n809), .B1(new_n874), .B2(new_n875), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n890), .A2(KEYINPUT100), .ZN(new_n891));
  INV_X1    g0691(.A(KEYINPUT100), .ZN(new_n892));
  NAND3_X1  g0692(.A1(new_n888), .A2(new_n892), .A3(new_n889), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n869), .A2(new_n861), .ZN(new_n894));
  NAND4_X1  g0694(.A1(new_n891), .A2(KEYINPUT40), .A3(new_n893), .A4(new_n894), .ZN(new_n895));
  AND3_X1   g0695(.A1(new_n852), .A2(KEYINPUT38), .A3(new_n858), .ZN(new_n896));
  OAI211_X1 g0696(.A(new_n888), .B(new_n889), .C1(new_n896), .C2(new_n859), .ZN(new_n897));
  INV_X1    g0697(.A(KEYINPUT40), .ZN(new_n898));
  AOI21_X1  g0698(.A(new_n798), .B1(new_n897), .B2(new_n898), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n895), .A2(new_n899), .ZN(new_n900));
  AND2_X1   g0700(.A1(new_n423), .A2(new_n888), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n901), .A2(G330), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n900), .A2(new_n902), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n897), .A2(new_n898), .ZN(new_n904));
  NAND3_X1  g0704(.A1(new_n895), .A2(new_n904), .A3(new_n901), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n903), .A2(new_n905), .ZN(new_n906));
  XNOR2_X1  g0706(.A(new_n882), .B(new_n906), .ZN(new_n907));
  OAI21_X1  g0707(.A(new_n907), .B1(new_n209), .B2(new_n655), .ZN(new_n908));
  OR2_X1    g0708(.A1(new_n528), .A2(new_n530), .ZN(new_n909));
  AOI21_X1  g0709(.A(new_n216), .B1(new_n909), .B2(KEYINPUT35), .ZN(new_n910));
  OAI211_X1 g0710(.A(new_n910), .B(new_n234), .C1(KEYINPUT35), .C2(new_n909), .ZN(new_n911));
  XNOR2_X1  g0711(.A(new_n911), .B(KEYINPUT36), .ZN(new_n912));
  OAI21_X1  g0712(.A(G77), .B1(new_n220), .B2(new_n224), .ZN(new_n913));
  OAI22_X1  g0713(.A1(new_n913), .A2(new_n235), .B1(G50), .B2(new_n224), .ZN(new_n914));
  NAND3_X1  g0714(.A1(new_n914), .A2(G1), .A3(new_n654), .ZN(new_n915));
  NAND3_X1  g0715(.A1(new_n908), .A2(new_n912), .A3(new_n915), .ZN(G367));
  NAND2_X1  g0716(.A1(new_n784), .A2(G283), .ZN(new_n917));
  NAND3_X1  g0717(.A1(new_n838), .A2(KEYINPUT46), .A3(G116), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n773), .A2(G317), .ZN(new_n919));
  NAND3_X1  g0719(.A1(new_n917), .A2(new_n918), .A3(new_n919), .ZN(new_n920));
  NOR2_X1   g0720(.A1(new_n769), .A2(new_n818), .ZN(new_n921));
  NOR2_X1   g0721(.A1(new_n756), .A2(new_n763), .ZN(new_n922));
  AOI21_X1  g0722(.A(KEYINPUT46), .B1(new_n838), .B2(G116), .ZN(new_n923));
  NOR4_X1   g0723(.A1(new_n920), .A2(new_n921), .A3(new_n922), .A4(new_n923), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n776), .A2(G311), .ZN(new_n925));
  AOI21_X1  g0725(.A(new_n500), .B1(G97), .B2(new_n788), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n782), .A2(G107), .ZN(new_n927));
  NAND4_X1  g0727(.A1(new_n924), .A2(new_n925), .A3(new_n926), .A4(new_n927), .ZN(new_n928));
  XOR2_X1   g0728(.A(new_n928), .B(KEYINPUT105), .Z(new_n929));
  NAND2_X1  g0729(.A1(new_n776), .A2(G143), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n784), .A2(G50), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n782), .A2(G68), .ZN(new_n932));
  NAND3_X1  g0732(.A1(new_n930), .A2(new_n931), .A3(new_n932), .ZN(new_n933));
  NOR2_X1   g0733(.A1(new_n760), .A2(new_n355), .ZN(new_n934));
  OAI22_X1  g0734(.A1(new_n762), .A2(new_n220), .B1(new_n772), .B2(new_n826), .ZN(new_n935));
  NOR3_X1   g0735(.A1(new_n933), .A2(new_n934), .A3(new_n935), .ZN(new_n936));
  AOI21_X1  g0736(.A(new_n339), .B1(new_n757), .B2(G150), .ZN(new_n937));
  OAI211_X1 g0737(.A(new_n936), .B(new_n937), .C1(new_n791), .C2(new_n769), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n929), .A2(new_n938), .ZN(new_n939));
  XOR2_X1   g0739(.A(new_n939), .B(KEYINPUT106), .Z(new_n940));
  XNOR2_X1  g0740(.A(new_n940), .B(KEYINPUT47), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n941), .A2(new_n751), .ZN(new_n942));
  NOR2_X1   g0742(.A1(new_n631), .A2(new_n662), .ZN(new_n943));
  MUX2_X1   g0743(.A(new_n634), .B(new_n627), .S(new_n943), .Z(new_n944));
  XNOR2_X1  g0744(.A(new_n944), .B(KEYINPUT101), .ZN(new_n945));
  INV_X1    g0745(.A(new_n739), .ZN(new_n946));
  OR2_X1    g0746(.A1(new_n945), .A2(new_n946), .ZN(new_n947));
  OAI221_X1 g0747(.A(new_n752), .B1(new_n230), .B2(new_n376), .C1(new_n247), .C2(new_n744), .ZN(new_n948));
  NAND4_X1  g0748(.A1(new_n942), .A2(new_n743), .A3(new_n947), .A4(new_n948), .ZN(new_n949));
  INV_X1    g0749(.A(KEYINPUT107), .ZN(new_n950));
  XNOR2_X1  g0750(.A(new_n949), .B(new_n950), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n741), .A2(G1), .ZN(new_n952));
  INV_X1    g0752(.A(KEYINPUT44), .ZN(new_n953));
  OAI211_X1 g0753(.A(new_n649), .B(new_n551), .C1(new_n537), .C2(new_n662), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n636), .A2(new_n661), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n954), .A2(new_n955), .ZN(new_n956));
  OAI21_X1  g0756(.A(new_n953), .B1(new_n679), .B2(new_n956), .ZN(new_n957));
  INV_X1    g0757(.A(new_n669), .ZN(new_n958));
  OAI21_X1  g0758(.A(new_n958), .B1(new_n673), .B2(new_n677), .ZN(new_n959));
  INV_X1    g0759(.A(new_n956), .ZN(new_n960));
  NAND3_X1  g0760(.A1(new_n959), .A2(KEYINPUT44), .A3(new_n960), .ZN(new_n961));
  NAND3_X1  g0761(.A1(new_n957), .A2(KEYINPUT104), .A3(new_n961), .ZN(new_n962));
  INV_X1    g0762(.A(KEYINPUT104), .ZN(new_n963));
  OAI211_X1 g0763(.A(new_n963), .B(new_n953), .C1(new_n679), .C2(new_n956), .ZN(new_n964));
  AOI21_X1  g0764(.A(KEYINPUT45), .B1(new_n679), .B2(new_n956), .ZN(new_n965));
  AND3_X1   g0765(.A1(new_n679), .A2(KEYINPUT45), .A3(new_n956), .ZN(new_n966));
  OAI211_X1 g0766(.A(new_n962), .B(new_n964), .C1(new_n965), .C2(new_n966), .ZN(new_n967));
  XNOR2_X1  g0767(.A(new_n967), .B(new_n674), .ZN(new_n968));
  NOR2_X1   g0768(.A1(new_n673), .A2(new_n669), .ZN(new_n969));
  XNOR2_X1  g0769(.A(new_n969), .B(new_n678), .ZN(new_n970));
  XNOR2_X1  g0770(.A(new_n970), .B(new_n668), .ZN(new_n971));
  OAI21_X1  g0771(.A(new_n734), .B1(new_n968), .B2(new_n971), .ZN(new_n972));
  XOR2_X1   g0772(.A(new_n681), .B(KEYINPUT41), .Z(new_n973));
  AOI21_X1  g0773(.A(new_n952), .B1(new_n972), .B2(new_n973), .ZN(new_n974));
  NAND3_X1  g0774(.A1(new_n678), .A2(new_n672), .A3(new_n958), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n649), .A2(new_n551), .ZN(new_n976));
  OR3_X1    g0776(.A1(new_n975), .A2(KEYINPUT42), .A3(new_n976), .ZN(new_n977));
  OAI21_X1  g0777(.A(new_n649), .B1(new_n960), .B2(new_n476), .ZN(new_n978));
  NAND2_X1  g0778(.A1(new_n978), .A2(new_n662), .ZN(new_n979));
  OAI21_X1  g0779(.A(KEYINPUT42), .B1(new_n975), .B2(new_n976), .ZN(new_n980));
  NAND3_X1  g0780(.A1(new_n977), .A2(new_n979), .A3(new_n980), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n981), .A2(KEYINPUT102), .ZN(new_n982));
  NOR2_X1   g0782(.A1(new_n945), .A2(KEYINPUT43), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n982), .A2(new_n983), .ZN(new_n984));
  INV_X1    g0784(.A(KEYINPUT103), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n984), .A2(new_n985), .ZN(new_n986));
  INV_X1    g0786(.A(KEYINPUT102), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n945), .A2(KEYINPUT43), .ZN(new_n988));
  AOI21_X1  g0788(.A(new_n983), .B1(new_n987), .B2(new_n988), .ZN(new_n989));
  OAI211_X1 g0789(.A(new_n989), .B(new_n981), .C1(new_n987), .C2(new_n988), .ZN(new_n990));
  NAND3_X1  g0790(.A1(new_n982), .A2(KEYINPUT103), .A3(new_n983), .ZN(new_n991));
  NAND3_X1  g0791(.A1(new_n986), .A2(new_n990), .A3(new_n991), .ZN(new_n992));
  NOR2_X1   g0792(.A1(new_n675), .A2(new_n960), .ZN(new_n993));
  INV_X1    g0793(.A(new_n993), .ZN(new_n994));
  XNOR2_X1  g0794(.A(new_n992), .B(new_n994), .ZN(new_n995));
  OAI21_X1  g0795(.A(new_n951), .B1(new_n974), .B2(new_n995), .ZN(G387));
  INV_X1    g0796(.A(new_n971), .ZN(new_n997));
  NAND2_X1  g0797(.A1(new_n734), .A2(new_n997), .ZN(new_n998));
  INV_X1    g0798(.A(KEYINPUT112), .ZN(new_n999));
  XOR2_X1   g0799(.A(new_n681), .B(KEYINPUT111), .Z(new_n1000));
  INV_X1    g0800(.A(new_n1000), .ZN(new_n1001));
  NAND3_X1  g0801(.A1(new_n998), .A2(new_n999), .A3(new_n1001), .ZN(new_n1002));
  AOI21_X1  g0802(.A(new_n971), .B1(new_n731), .B2(new_n733), .ZN(new_n1003));
  OAI21_X1  g0803(.A(KEYINPUT112), .B1(new_n1003), .B2(new_n1000), .ZN(new_n1004));
  OAI211_X1 g0804(.A(new_n1002), .B(new_n1004), .C1(new_n734), .C2(new_n997), .ZN(new_n1005));
  OAI21_X1  g0805(.A(new_n743), .B1(new_n969), .B2(new_n946), .ZN(new_n1006));
  AOI22_X1  g0806(.A1(new_n776), .A2(G322), .B1(new_n784), .B2(G303), .ZN(new_n1007));
  INV_X1    g0807(.A(G311), .ZN(new_n1008));
  INV_X1    g0808(.A(G317), .ZN(new_n1009));
  OAI221_X1 g0809(.A(new_n1007), .B1(new_n1008), .B2(new_n769), .C1(new_n1009), .C2(new_n756), .ZN(new_n1010));
  XNOR2_X1  g0810(.A(new_n1010), .B(KEYINPUT48), .ZN(new_n1011));
  OAI221_X1 g0811(.A(new_n1011), .B1(new_n761), .B2(new_n781), .C1(new_n818), .C2(new_n762), .ZN(new_n1012));
  XNOR2_X1  g0812(.A(new_n1012), .B(KEYINPUT49), .ZN(new_n1013));
  OAI221_X1 g0813(.A(new_n258), .B1(new_n216), .B2(new_n760), .C1(new_n778), .C2(new_n772), .ZN(new_n1014));
  XNOR2_X1  g0814(.A(new_n1014), .B(KEYINPUT110), .ZN(new_n1015));
  NAND2_X1  g0815(.A1(new_n1013), .A2(new_n1015), .ZN(new_n1016));
  NAND2_X1  g0816(.A1(new_n787), .A2(G159), .ZN(new_n1017));
  XOR2_X1   g0817(.A(new_n1017), .B(KEYINPUT109), .Z(new_n1018));
  NAND2_X1  g0818(.A1(new_n782), .A2(new_n375), .ZN(new_n1019));
  OAI221_X1 g0819(.A(new_n1019), .B1(new_n355), .B2(new_n762), .C1(new_n205), .C2(new_n760), .ZN(new_n1020));
  OAI22_X1  g0820(.A1(new_n756), .A2(new_n202), .B1(new_n766), .B2(new_n224), .ZN(new_n1021));
  NOR4_X1   g0821(.A1(new_n1018), .A2(new_n258), .A3(new_n1020), .A4(new_n1021), .ZN(new_n1022));
  OAI221_X1 g0822(.A(new_n1022), .B1(new_n396), .B2(new_n772), .C1(new_n290), .C2(new_n769), .ZN(new_n1023));
  AOI21_X1  g0823(.A(new_n841), .B1(new_n1016), .B2(new_n1023), .ZN(new_n1024));
  NOR3_X1   g0824(.A1(new_n290), .A2(KEYINPUT50), .A3(G50), .ZN(new_n1025));
  INV_X1    g0825(.A(new_n682), .ZN(new_n1026));
  NOR2_X1   g0826(.A1(new_n1025), .A2(new_n1026), .ZN(new_n1027));
  NAND2_X1  g0827(.A1(G68), .A2(G77), .ZN(new_n1028));
  OAI21_X1  g0828(.A(KEYINPUT50), .B1(new_n290), .B2(G50), .ZN(new_n1029));
  NAND4_X1  g0829(.A1(new_n1027), .A2(new_n746), .A3(new_n1028), .A4(new_n1029), .ZN(new_n1030));
  OAI211_X1 g0830(.A(new_n745), .B(new_n1030), .C1(new_n243), .C2(new_n746), .ZN(new_n1031));
  NAND3_X1  g0831(.A1(new_n1026), .A2(new_n230), .A3(new_n380), .ZN(new_n1032));
  OAI211_X1 g0832(.A(new_n1031), .B(new_n1032), .C1(G107), .C2(new_n230), .ZN(new_n1033));
  XNOR2_X1  g0833(.A(new_n1033), .B(KEYINPUT108), .ZN(new_n1034));
  AOI211_X1 g0834(.A(new_n1006), .B(new_n1024), .C1(new_n752), .C2(new_n1034), .ZN(new_n1035));
  AOI21_X1  g0835(.A(new_n1035), .B1(new_n997), .B2(new_n952), .ZN(new_n1036));
  NAND2_X1  g0836(.A1(new_n1005), .A2(new_n1036), .ZN(G393));
  XNOR2_X1  g0837(.A(new_n967), .B(new_n675), .ZN(new_n1038));
  AOI21_X1  g0838(.A(new_n1000), .B1(new_n1003), .B2(new_n1038), .ZN(new_n1039));
  OAI21_X1  g0839(.A(new_n1039), .B1(new_n1038), .B2(new_n1003), .ZN(new_n1040));
  AOI21_X1  g0840(.A(new_n742), .B1(new_n960), .B2(new_n739), .ZN(new_n1041));
  OAI21_X1  g0841(.A(new_n339), .B1(new_n781), .B2(new_n216), .ZN(new_n1042));
  OAI22_X1  g0842(.A1(new_n1008), .A2(new_n756), .B1(new_n775), .B2(new_n1009), .ZN(new_n1043));
  XNOR2_X1  g0843(.A(new_n1043), .B(KEYINPUT52), .ZN(new_n1044));
  INV_X1    g0844(.A(G322), .ZN(new_n1045));
  OAI22_X1  g0845(.A1(new_n762), .A2(new_n761), .B1(new_n772), .B2(new_n1045), .ZN(new_n1046));
  AOI21_X1  g0846(.A(new_n1046), .B1(new_n824), .B2(G303), .ZN(new_n1047));
  OAI211_X1 g0847(.A(new_n1044), .B(new_n1047), .C1(new_n818), .C2(new_n766), .ZN(new_n1048));
  AOI211_X1 g0848(.A(new_n1042), .B(new_n1048), .C1(G107), .C2(new_n788), .ZN(new_n1049));
  OAI22_X1  g0849(.A1(new_n396), .A2(new_n775), .B1(new_n756), .B2(new_n791), .ZN(new_n1050));
  XOR2_X1   g0850(.A(new_n1050), .B(KEYINPUT51), .Z(new_n1051));
  AOI22_X1  g0851(.A1(new_n838), .A2(G68), .B1(new_n773), .B2(G143), .ZN(new_n1052));
  OAI211_X1 g0852(.A(new_n1052), .B(new_n500), .C1(new_n214), .C2(new_n760), .ZN(new_n1053));
  XNOR2_X1  g0853(.A(new_n1053), .B(KEYINPUT113), .ZN(new_n1054));
  OAI22_X1  g0854(.A1(new_n785), .A2(new_n290), .B1(new_n202), .B2(new_n769), .ZN(new_n1055));
  NOR2_X1   g0855(.A1(new_n781), .A2(new_n355), .ZN(new_n1056));
  NOR4_X1   g0856(.A1(new_n1051), .A2(new_n1054), .A3(new_n1055), .A4(new_n1056), .ZN(new_n1057));
  OAI21_X1  g0857(.A(new_n751), .B1(new_n1049), .B2(new_n1057), .ZN(new_n1058));
  OAI221_X1 g0858(.A(new_n752), .B1(new_n205), .B2(new_n230), .C1(new_n251), .C2(new_n744), .ZN(new_n1059));
  AND3_X1   g0859(.A1(new_n1041), .A2(new_n1058), .A3(new_n1059), .ZN(new_n1060));
  AOI21_X1  g0860(.A(new_n1060), .B1(new_n1038), .B2(new_n952), .ZN(new_n1061));
  NAND2_X1  g0861(.A1(new_n1040), .A2(new_n1061), .ZN(G390));
  NAND2_X1  g0862(.A1(new_n806), .A2(new_n877), .ZN(new_n1063));
  NAND2_X1  g0863(.A1(new_n874), .A2(new_n875), .ZN(new_n1064));
  NOR2_X1   g0864(.A1(new_n809), .A2(new_n798), .ZN(new_n1065));
  NAND3_X1  g0865(.A1(new_n888), .A2(new_n1064), .A3(new_n1065), .ZN(new_n1066));
  INV_X1    g0866(.A(new_n1066), .ZN(new_n1067));
  AOI21_X1  g0867(.A(new_n1064), .B1(new_n728), .B2(new_n1065), .ZN(new_n1068));
  OAI21_X1  g0868(.A(new_n1063), .B1(new_n1067), .B2(new_n1068), .ZN(new_n1069));
  NAND2_X1  g0869(.A1(new_n888), .A2(new_n1065), .ZN(new_n1070));
  NAND2_X1  g0870(.A1(new_n1070), .A2(new_n876), .ZN(new_n1071));
  NAND3_X1  g0871(.A1(new_n701), .A2(new_n662), .A3(new_n805), .ZN(new_n1072));
  NAND3_X1  g0872(.A1(new_n728), .A2(new_n1064), .A3(new_n1065), .ZN(new_n1073));
  NAND4_X1  g0873(.A1(new_n1071), .A2(new_n877), .A3(new_n1072), .A4(new_n1073), .ZN(new_n1074));
  NAND2_X1  g0874(.A1(new_n1069), .A2(new_n1074), .ZN(new_n1075));
  NAND4_X1  g0875(.A1(new_n1075), .A2(new_n844), .A3(new_n624), .A4(new_n902), .ZN(new_n1076));
  INV_X1    g0876(.A(new_n1076), .ZN(new_n1077));
  OAI21_X1  g0877(.A(KEYINPUT39), .B1(new_n896), .B2(new_n859), .ZN(new_n1078));
  OAI211_X1 g0878(.A(new_n1078), .B(new_n870), .C1(new_n878), .C2(new_n846), .ZN(new_n1079));
  AOI21_X1  g0879(.A(new_n876), .B1(new_n1072), .B2(new_n877), .ZN(new_n1080));
  OAI21_X1  g0880(.A(new_n894), .B1(new_n368), .B2(new_n661), .ZN(new_n1081));
  OAI21_X1  g0881(.A(new_n1079), .B1(new_n1080), .B2(new_n1081), .ZN(new_n1082));
  NAND2_X1  g0882(.A1(new_n1082), .A2(new_n1066), .ZN(new_n1083));
  INV_X1    g0883(.A(new_n1073), .ZN(new_n1084));
  OAI211_X1 g0884(.A(new_n1084), .B(new_n1079), .C1(new_n1080), .C2(new_n1081), .ZN(new_n1085));
  NAND2_X1  g0885(.A1(new_n1083), .A2(new_n1085), .ZN(new_n1086));
  NAND2_X1  g0886(.A1(new_n1077), .A2(new_n1086), .ZN(new_n1087));
  NAND3_X1  g0887(.A1(new_n1076), .A2(new_n1083), .A3(new_n1085), .ZN(new_n1088));
  AND3_X1   g0888(.A1(new_n1087), .A2(new_n1001), .A3(new_n1088), .ZN(new_n1089));
  INV_X1    g0889(.A(new_n1089), .ZN(new_n1090));
  NAND2_X1  g0890(.A1(new_n1086), .A2(new_n952), .ZN(new_n1091));
  NAND3_X1  g0891(.A1(new_n1078), .A2(new_n737), .A3(new_n870), .ZN(new_n1092));
  AOI21_X1  g0892(.A(new_n380), .B1(new_n784), .B2(G97), .ZN(new_n1093));
  OAI22_X1  g0893(.A1(new_n206), .A2(new_n769), .B1(new_n756), .B2(new_n216), .ZN(new_n1094));
  AOI21_X1  g0894(.A(new_n1094), .B1(G283), .B2(new_n787), .ZN(new_n1095));
  AOI211_X1 g0895(.A(new_n836), .B(new_n1056), .C1(G87), .C2(new_n838), .ZN(new_n1096));
  NAND3_X1  g0896(.A1(new_n1093), .A2(new_n1095), .A3(new_n1096), .ZN(new_n1097));
  AOI21_X1  g0897(.A(new_n1097), .B1(G294), .B2(new_n773), .ZN(new_n1098));
  XNOR2_X1  g0898(.A(new_n1098), .B(KEYINPUT115), .ZN(new_n1099));
  OAI22_X1  g0899(.A1(new_n833), .A2(new_n756), .B1(new_n769), .B2(new_n826), .ZN(new_n1100));
  NOR2_X1   g0900(.A1(new_n762), .A2(new_n396), .ZN(new_n1101));
  XNOR2_X1  g0901(.A(new_n1101), .B(KEYINPUT114), .ZN(new_n1102));
  NOR2_X1   g0902(.A1(new_n1102), .A2(KEYINPUT53), .ZN(new_n1103));
  AOI211_X1 g0903(.A(new_n1100), .B(new_n1103), .C1(G128), .C2(new_n787), .ZN(new_n1104));
  XOR2_X1   g0904(.A(KEYINPUT54), .B(G143), .Z(new_n1105));
  AOI22_X1  g0905(.A1(new_n784), .A2(new_n1105), .B1(new_n1102), .B2(KEYINPUT53), .ZN(new_n1106));
  OAI21_X1  g0906(.A(new_n380), .B1(new_n781), .B2(new_n791), .ZN(new_n1107));
  AOI21_X1  g0907(.A(new_n1107), .B1(G50), .B2(new_n788), .ZN(new_n1108));
  NAND3_X1  g0908(.A1(new_n1104), .A2(new_n1106), .A3(new_n1108), .ZN(new_n1109));
  AOI21_X1  g0909(.A(new_n1109), .B1(G125), .B2(new_n773), .ZN(new_n1110));
  OAI21_X1  g0910(.A(new_n751), .B1(new_n1099), .B2(new_n1110), .ZN(new_n1111));
  NAND2_X1  g0911(.A1(new_n814), .A2(new_n290), .ZN(new_n1112));
  NAND4_X1  g0912(.A1(new_n1092), .A2(new_n743), .A3(new_n1111), .A4(new_n1112), .ZN(new_n1113));
  NAND3_X1  g0913(.A1(new_n1091), .A2(KEYINPUT116), .A3(new_n1113), .ZN(new_n1114));
  INV_X1    g0914(.A(KEYINPUT116), .ZN(new_n1115));
  INV_X1    g0915(.A(new_n952), .ZN(new_n1116));
  AOI21_X1  g0916(.A(new_n1116), .B1(new_n1083), .B2(new_n1085), .ZN(new_n1117));
  INV_X1    g0917(.A(new_n1113), .ZN(new_n1118));
  OAI21_X1  g0918(.A(new_n1115), .B1(new_n1117), .B2(new_n1118), .ZN(new_n1119));
  NAND3_X1  g0919(.A1(new_n1114), .A2(KEYINPUT117), .A3(new_n1119), .ZN(new_n1120));
  INV_X1    g0920(.A(new_n1120), .ZN(new_n1121));
  AOI21_X1  g0921(.A(KEYINPUT117), .B1(new_n1114), .B2(new_n1119), .ZN(new_n1122));
  OAI21_X1  g0922(.A(new_n1090), .B1(new_n1121), .B2(new_n1122), .ZN(G378));
  INV_X1    g0923(.A(new_n881), .ZN(new_n1124));
  NAND2_X1  g0924(.A1(new_n409), .A2(new_n848), .ZN(new_n1125));
  NAND3_X1  g0925(.A1(new_n619), .A2(new_n408), .A3(new_n1125), .ZN(new_n1126));
  INV_X1    g0926(.A(new_n1125), .ZN(new_n1127));
  NAND2_X1  g0927(.A1(new_n418), .A2(new_n1127), .ZN(new_n1128));
  XNOR2_X1  g0928(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1129));
  AND3_X1   g0929(.A1(new_n1126), .A2(new_n1128), .A3(new_n1129), .ZN(new_n1130));
  AOI21_X1  g0930(.A(new_n1129), .B1(new_n1126), .B2(new_n1128), .ZN(new_n1131));
  NOR2_X1   g0931(.A1(new_n1130), .A2(new_n1131), .ZN(new_n1132));
  AND3_X1   g0932(.A1(new_n895), .A2(new_n899), .A3(new_n1132), .ZN(new_n1133));
  AOI21_X1  g0933(.A(new_n1132), .B1(new_n895), .B2(new_n899), .ZN(new_n1134));
  OAI21_X1  g0934(.A(new_n1124), .B1(new_n1133), .B2(new_n1134), .ZN(new_n1135));
  INV_X1    g0935(.A(new_n1132), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n900), .A2(new_n1136), .ZN(new_n1137));
  NAND3_X1  g0937(.A1(new_n895), .A2(new_n899), .A3(new_n1132), .ZN(new_n1138));
  NAND3_X1  g0938(.A1(new_n1137), .A2(new_n881), .A3(new_n1138), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n1135), .A2(new_n1139), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n1140), .A2(new_n952), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n1132), .A2(new_n737), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n787), .A2(G116), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n757), .A2(G107), .ZN(new_n1144));
  NAND4_X1  g0944(.A1(new_n1143), .A2(new_n1144), .A3(new_n267), .A4(new_n932), .ZN(new_n1145));
  NAND2_X1  g0945(.A1(new_n265), .A2(new_n304), .ZN(new_n1146));
  NOR2_X1   g0946(.A1(new_n772), .A2(new_n761), .ZN(new_n1147));
  AOI211_X1 g0947(.A(new_n1146), .B(new_n1147), .C1(G77), .C2(new_n838), .ZN(new_n1148));
  NOR2_X1   g0948(.A1(new_n760), .A2(new_n220), .ZN(new_n1149));
  XNOR2_X1  g0949(.A(new_n1149), .B(KEYINPUT118), .ZN(new_n1150));
  OAI211_X1 g0950(.A(new_n1148), .B(new_n1150), .C1(new_n205), .C2(new_n769), .ZN(new_n1151));
  AOI211_X1 g0951(.A(new_n1145), .B(new_n1151), .C1(new_n375), .C2(new_n767), .ZN(new_n1152));
  XNOR2_X1  g0952(.A(new_n1152), .B(KEYINPUT119), .ZN(new_n1153));
  OR2_X1    g0953(.A1(new_n1153), .A2(KEYINPUT58), .ZN(new_n1154));
  NAND2_X1  g0954(.A1(new_n1153), .A2(KEYINPUT58), .ZN(new_n1155));
  INV_X1    g0955(.A(G124), .ZN(new_n1156));
  OAI21_X1  g0956(.A(new_n266), .B1(new_n772), .B2(new_n1156), .ZN(new_n1157));
  OAI22_X1  g0957(.A1(new_n769), .A2(new_n833), .B1(new_n766), .B2(new_n826), .ZN(new_n1158));
  AOI21_X1  g0958(.A(new_n1158), .B1(G128), .B2(new_n757), .ZN(new_n1159));
  AOI22_X1  g0959(.A1(new_n787), .A2(G125), .B1(new_n838), .B2(new_n1105), .ZN(new_n1160));
  OAI211_X1 g0960(.A(new_n1159), .B(new_n1160), .C1(new_n396), .C2(new_n781), .ZN(new_n1161));
  AOI211_X1 g0961(.A(G41), .B(new_n1157), .C1(new_n1161), .C2(KEYINPUT59), .ZN(new_n1162));
  OAI221_X1 g0962(.A(new_n1162), .B1(KEYINPUT59), .B2(new_n1161), .C1(new_n791), .C2(new_n760), .ZN(new_n1163));
  NAND2_X1  g0963(.A1(new_n1146), .A2(new_n202), .ZN(new_n1164));
  NAND4_X1  g0964(.A1(new_n1154), .A2(new_n1155), .A3(new_n1163), .A4(new_n1164), .ZN(new_n1165));
  NAND2_X1  g0965(.A1(new_n1165), .A2(new_n751), .ZN(new_n1166));
  NAND2_X1  g0966(.A1(new_n813), .A2(new_n202), .ZN(new_n1167));
  NAND4_X1  g0967(.A1(new_n1142), .A2(new_n743), .A3(new_n1166), .A4(new_n1167), .ZN(new_n1168));
  NAND2_X1  g0968(.A1(new_n1141), .A2(new_n1168), .ZN(new_n1169));
  INV_X1    g0969(.A(new_n1169), .ZN(new_n1170));
  INV_X1    g0970(.A(KEYINPUT57), .ZN(new_n1171));
  AND2_X1   g0971(.A1(new_n1135), .A2(new_n1139), .ZN(new_n1172));
  NAND3_X1  g0972(.A1(new_n844), .A2(new_n624), .A3(new_n902), .ZN(new_n1173));
  AOI21_X1  g0973(.A(new_n1173), .B1(new_n1086), .B2(new_n1075), .ZN(new_n1174));
  OAI21_X1  g0974(.A(new_n1171), .B1(new_n1172), .B2(new_n1174), .ZN(new_n1175));
  NAND2_X1  g0975(.A1(new_n1175), .A2(new_n1001), .ZN(new_n1176));
  AOI21_X1  g0976(.A(new_n1076), .B1(new_n1083), .B2(new_n1085), .ZN(new_n1177));
  OAI21_X1  g0977(.A(KEYINPUT57), .B1(new_n1177), .B2(new_n1173), .ZN(new_n1178));
  NAND3_X1  g0978(.A1(new_n1135), .A2(new_n1139), .A3(KEYINPUT120), .ZN(new_n1179));
  INV_X1    g0979(.A(KEYINPUT120), .ZN(new_n1180));
  OAI211_X1 g0980(.A(new_n1180), .B(new_n1124), .C1(new_n1133), .C2(new_n1134), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n1179), .A2(new_n1181), .ZN(new_n1182));
  NOR2_X1   g0982(.A1(new_n1178), .A2(new_n1182), .ZN(new_n1183));
  OAI21_X1  g0983(.A(new_n1170), .B1(new_n1176), .B2(new_n1183), .ZN(G375));
  INV_X1    g0984(.A(KEYINPUT122), .ZN(new_n1185));
  XOR2_X1   g0985(.A(new_n952), .B(KEYINPUT121), .Z(new_n1186));
  AND3_X1   g0986(.A1(new_n1075), .A2(new_n1185), .A3(new_n1186), .ZN(new_n1187));
  AOI21_X1  g0987(.A(new_n1185), .B1(new_n1075), .B2(new_n1186), .ZN(new_n1188));
  NAND2_X1  g0988(.A1(new_n814), .A2(new_n224), .ZN(new_n1189));
  OAI21_X1  g0989(.A(new_n1189), .B1(new_n1064), .B2(new_n738), .ZN(new_n1190));
  INV_X1    g0990(.A(G128), .ZN(new_n1191));
  OAI21_X1  g0991(.A(new_n500), .B1(new_n1191), .B2(new_n772), .ZN(new_n1192));
  OAI221_X1 g0992(.A(new_n1150), .B1(new_n396), .B2(new_n766), .C1(new_n791), .C2(new_n762), .ZN(new_n1193));
  AOI211_X1 g0993(.A(new_n1192), .B(new_n1193), .C1(G50), .C2(new_n782), .ZN(new_n1194));
  INV_X1    g0994(.A(new_n1194), .ZN(new_n1195));
  AOI22_X1  g0995(.A1(new_n1195), .A2(KEYINPUT123), .B1(G137), .B2(new_n757), .ZN(new_n1196));
  INV_X1    g0996(.A(KEYINPUT123), .ZN(new_n1197));
  AOI22_X1  g0997(.A1(new_n1194), .A2(new_n1197), .B1(new_n824), .B2(new_n1105), .ZN(new_n1198));
  OAI211_X1 g0998(.A(new_n1196), .B(new_n1198), .C1(new_n833), .C2(new_n775), .ZN(new_n1199));
  NOR2_X1   g0999(.A1(new_n775), .A2(new_n818), .ZN(new_n1200));
  OAI21_X1  g1000(.A(new_n1019), .B1(new_n205), .B2(new_n762), .ZN(new_n1201));
  AOI211_X1 g1001(.A(new_n934), .B(new_n1201), .C1(G303), .C2(new_n773), .ZN(new_n1202));
  AOI21_X1  g1002(.A(new_n380), .B1(new_n784), .B2(G107), .ZN(new_n1203));
  AOI22_X1  g1003(.A1(new_n824), .A2(G116), .B1(new_n757), .B2(G283), .ZN(new_n1204));
  NAND3_X1  g1004(.A1(new_n1202), .A2(new_n1203), .A3(new_n1204), .ZN(new_n1205));
  OAI21_X1  g1005(.A(new_n1199), .B1(new_n1200), .B2(new_n1205), .ZN(new_n1206));
  AOI211_X1 g1006(.A(new_n742), .B(new_n1190), .C1(new_n751), .C2(new_n1206), .ZN(new_n1207));
  NOR3_X1   g1007(.A1(new_n1187), .A2(new_n1188), .A3(new_n1207), .ZN(new_n1208));
  INV_X1    g1008(.A(new_n1075), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(new_n1173), .A2(new_n1209), .ZN(new_n1210));
  NAND3_X1  g1010(.A1(new_n1210), .A2(new_n973), .A3(new_n1076), .ZN(new_n1211));
  NAND2_X1  g1011(.A1(new_n1208), .A2(new_n1211), .ZN(G381));
  OR2_X1    g1012(.A1(new_n1178), .A2(new_n1182), .ZN(new_n1213));
  OAI21_X1  g1013(.A(new_n1140), .B1(new_n1177), .B2(new_n1173), .ZN(new_n1214));
  AOI21_X1  g1014(.A(new_n1000), .B1(new_n1214), .B2(new_n1171), .ZN(new_n1215));
  AOI21_X1  g1015(.A(new_n1169), .B1(new_n1213), .B2(new_n1215), .ZN(new_n1216));
  AOI21_X1  g1016(.A(KEYINPUT116), .B1(new_n1091), .B2(new_n1113), .ZN(new_n1217));
  NOR3_X1   g1017(.A1(new_n1117), .A2(new_n1115), .A3(new_n1118), .ZN(new_n1218));
  NOR3_X1   g1018(.A1(new_n1089), .A2(new_n1217), .A3(new_n1218), .ZN(new_n1219));
  AND2_X1   g1019(.A1(new_n1216), .A2(new_n1219), .ZN(new_n1220));
  NOR2_X1   g1020(.A1(G381), .A2(G384), .ZN(new_n1221));
  AOI22_X1  g1021(.A1(new_n1038), .A2(new_n997), .B1(new_n731), .B2(new_n733), .ZN(new_n1222));
  INV_X1    g1022(.A(new_n973), .ZN(new_n1223));
  OAI21_X1  g1023(.A(new_n1116), .B1(new_n1222), .B2(new_n1223), .ZN(new_n1224));
  XNOR2_X1  g1024(.A(new_n992), .B(new_n993), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(new_n1224), .A2(new_n1225), .ZN(new_n1226));
  NAND4_X1  g1026(.A1(new_n1226), .A2(new_n1040), .A3(new_n951), .A4(new_n1061), .ZN(new_n1227));
  INV_X1    g1027(.A(new_n1227), .ZN(new_n1228));
  NOR2_X1   g1028(.A1(G393), .A2(G396), .ZN(new_n1229));
  NAND4_X1  g1029(.A1(new_n1220), .A2(new_n1221), .A3(new_n1228), .A4(new_n1229), .ZN(G407));
  INV_X1    g1030(.A(G213), .ZN(new_n1231));
  AOI21_X1  g1031(.A(new_n1231), .B1(new_n1220), .B2(new_n660), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(new_n1232), .A2(G407), .ZN(G409));
  NAND2_X1  g1033(.A1(G387), .A2(G390), .ZN(new_n1234));
  INV_X1    g1034(.A(KEYINPUT125), .ZN(new_n1235));
  AND3_X1   g1035(.A1(new_n1234), .A2(new_n1235), .A3(new_n1227), .ZN(new_n1236));
  AOI21_X1  g1036(.A(new_n1235), .B1(new_n1234), .B2(new_n1227), .ZN(new_n1237));
  AOI22_X1  g1037(.A1(new_n1005), .A2(new_n1036), .B1(new_n797), .B2(new_n800), .ZN(new_n1238));
  OAI22_X1  g1038(.A1(new_n1236), .A2(new_n1237), .B1(new_n1229), .B2(new_n1238), .ZN(new_n1239));
  NAND2_X1  g1039(.A1(new_n1234), .A2(new_n1227), .ZN(new_n1240));
  NAND2_X1  g1040(.A1(new_n1240), .A2(KEYINPUT125), .ZN(new_n1241));
  NOR2_X1   g1041(.A1(new_n1229), .A2(new_n1238), .ZN(new_n1242));
  NAND3_X1  g1042(.A1(new_n1234), .A2(new_n1235), .A3(new_n1227), .ZN(new_n1243));
  NAND3_X1  g1043(.A1(new_n1241), .A2(new_n1242), .A3(new_n1243), .ZN(new_n1244));
  NAND3_X1  g1044(.A1(new_n1179), .A2(new_n1181), .A3(new_n1186), .ZN(new_n1245));
  OAI211_X1 g1045(.A(new_n1245), .B(new_n1168), .C1(new_n1214), .C2(new_n1223), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(new_n1219), .A2(new_n1246), .ZN(new_n1247));
  INV_X1    g1047(.A(KEYINPUT117), .ZN(new_n1248));
  OAI21_X1  g1048(.A(new_n1248), .B1(new_n1217), .B2(new_n1218), .ZN(new_n1249));
  AOI21_X1  g1049(.A(new_n1089), .B1(new_n1249), .B2(new_n1120), .ZN(new_n1250));
  OAI21_X1  g1050(.A(new_n1247), .B1(G375), .B2(new_n1250), .ZN(new_n1251));
  INV_X1    g1051(.A(KEYINPUT60), .ZN(new_n1252));
  OAI211_X1 g1052(.A(new_n1001), .B(new_n1076), .C1(new_n1210), .C2(new_n1252), .ZN(new_n1253));
  AOI21_X1  g1053(.A(KEYINPUT60), .B1(new_n1173), .B2(new_n1209), .ZN(new_n1254));
  OAI21_X1  g1054(.A(new_n1208), .B1(new_n1253), .B2(new_n1254), .ZN(new_n1255));
  INV_X1    g1055(.A(G384), .ZN(new_n1256));
  OR2_X1    g1056(.A1(new_n1255), .A2(new_n1256), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(new_n1255), .A2(new_n1256), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(new_n1257), .A2(new_n1258), .ZN(new_n1259));
  INV_X1    g1059(.A(new_n1259), .ZN(new_n1260));
  NOR2_X1   g1060(.A1(new_n1231), .A2(G343), .ZN(new_n1261));
  INV_X1    g1061(.A(new_n1261), .ZN(new_n1262));
  NAND4_X1  g1062(.A1(new_n1251), .A2(new_n1260), .A3(KEYINPUT63), .A4(new_n1262), .ZN(new_n1263));
  AND3_X1   g1063(.A1(new_n1239), .A2(new_n1244), .A3(new_n1263), .ZN(new_n1264));
  INV_X1    g1064(.A(KEYINPUT61), .ZN(new_n1265));
  INV_X1    g1065(.A(KEYINPUT63), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(new_n1251), .A2(KEYINPUT124), .ZN(new_n1267));
  INV_X1    g1067(.A(KEYINPUT124), .ZN(new_n1268));
  OAI211_X1 g1068(.A(new_n1268), .B(new_n1247), .C1(G375), .C2(new_n1250), .ZN(new_n1269));
  NAND3_X1  g1069(.A1(new_n1267), .A2(new_n1262), .A3(new_n1269), .ZN(new_n1270));
  INV_X1    g1070(.A(G2897), .ZN(new_n1271));
  NOR3_X1   g1071(.A1(new_n1259), .A2(new_n1271), .A3(new_n1262), .ZN(new_n1272));
  AOI22_X1  g1072(.A1(new_n1257), .A2(new_n1258), .B1(G2897), .B2(new_n1261), .ZN(new_n1273));
  OR2_X1    g1073(.A1(new_n1272), .A2(new_n1273), .ZN(new_n1274));
  AOI21_X1  g1074(.A(new_n1266), .B1(new_n1270), .B2(new_n1274), .ZN(new_n1275));
  NAND4_X1  g1075(.A1(new_n1267), .A2(new_n1262), .A3(new_n1260), .A4(new_n1269), .ZN(new_n1276));
  INV_X1    g1076(.A(new_n1276), .ZN(new_n1277));
  OAI211_X1 g1077(.A(new_n1264), .B(new_n1265), .C1(new_n1275), .C2(new_n1277), .ZN(new_n1278));
  NAND2_X1  g1078(.A1(new_n1239), .A2(new_n1244), .ZN(new_n1279));
  AOI22_X1  g1079(.A1(new_n1216), .A2(G378), .B1(new_n1219), .B2(new_n1246), .ZN(new_n1280));
  NAND3_X1  g1080(.A1(new_n1257), .A2(KEYINPUT62), .A3(new_n1258), .ZN(new_n1281));
  NOR3_X1   g1081(.A1(new_n1280), .A2(new_n1261), .A3(new_n1281), .ZN(new_n1282));
  XNOR2_X1  g1082(.A(KEYINPUT126), .B(KEYINPUT62), .ZN(new_n1283));
  AOI21_X1  g1083(.A(new_n1282), .B1(new_n1276), .B2(new_n1283), .ZN(new_n1284));
  NOR2_X1   g1084(.A1(new_n1272), .A2(new_n1273), .ZN(new_n1285));
  NOR2_X1   g1085(.A1(new_n1280), .A2(new_n1261), .ZN(new_n1286));
  OAI21_X1  g1086(.A(new_n1265), .B1(new_n1285), .B2(new_n1286), .ZN(new_n1287));
  OAI21_X1  g1087(.A(new_n1279), .B1(new_n1284), .B2(new_n1287), .ZN(new_n1288));
  NAND2_X1  g1088(.A1(new_n1278), .A2(new_n1288), .ZN(G405));
  NAND2_X1  g1089(.A1(new_n1279), .A2(KEYINPUT127), .ZN(new_n1290));
  NAND2_X1  g1090(.A1(G375), .A2(new_n1219), .ZN(new_n1291));
  OAI21_X1  g1091(.A(new_n1291), .B1(new_n1250), .B2(G375), .ZN(new_n1292));
  XNOR2_X1  g1092(.A(new_n1292), .B(new_n1260), .ZN(new_n1293));
  INV_X1    g1093(.A(KEYINPUT127), .ZN(new_n1294));
  NAND3_X1  g1094(.A1(new_n1239), .A2(new_n1244), .A3(new_n1294), .ZN(new_n1295));
  NAND3_X1  g1095(.A1(new_n1290), .A2(new_n1293), .A3(new_n1295), .ZN(new_n1296));
  OR2_X1    g1096(.A1(new_n1293), .A2(new_n1295), .ZN(new_n1297));
  NAND2_X1  g1097(.A1(new_n1296), .A2(new_n1297), .ZN(G402));
endmodule


