

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360,
         n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371,
         n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382,
         n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393,
         n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404,
         n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415,
         n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426,
         n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437,
         n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448,
         n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459,
         n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470,
         n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481,
         n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492,
         n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503,
         n504, n505, n506, n507, n508, n509, n510, n511, n512, n513, n514,
         n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525,
         n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536,
         n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547,
         n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558,
         n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569,
         n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580,
         n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591,
         n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602,
         n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613,
         n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624,
         n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635,
         n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646,
         n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657,
         n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668,
         n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679,
         n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690,
         n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701,
         n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712,
         n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723,
         n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734,
         n735, n736, n737, n738, n739, n740, n741, n742, n743;

  XNOR2_X1 U371 ( .A(n375), .B(G107), .ZN(n450) );
  INV_X1 U372 ( .A(G116), .ZN(n375) );
  INV_X1 U373 ( .A(G953), .ZN(n737) );
  OR2_X2 U374 ( .A1(n509), .A2(n578), .ZN(n510) );
  XNOR2_X2 U375 ( .A(n422), .B(n421), .ZN(n553) );
  XOR2_X2 U376 ( .A(KEYINPUT77), .B(G110), .Z(n494) );
  AND2_X1 U377 ( .A1(n619), .A2(n634), .ZN(n540) );
  NAND2_X1 U378 ( .A1(n523), .A2(n564), .ZN(n503) );
  INV_X1 U379 ( .A(G119), .ZN(n365) );
  NOR2_X1 U380 ( .A1(n614), .A2(n718), .ZN(n615) );
  NOR2_X1 U381 ( .A1(n706), .A2(n718), .ZN(n708) );
  NOR2_X1 U382 ( .A1(n626), .A2(n718), .ZN(n628) );
  BUF_X1 U383 ( .A(n702), .Z(n712) );
  XNOR2_X1 U384 ( .A(n369), .B(n368), .ZN(n535) );
  XNOR2_X1 U385 ( .A(n376), .B(KEYINPUT32), .ZN(n619) );
  XNOR2_X1 U386 ( .A(n463), .B(n462), .ZN(n534) );
  XNOR2_X1 U387 ( .A(n396), .B(KEYINPUT39), .ZN(n595) );
  XNOR2_X1 U388 ( .A(n374), .B(KEYINPUT0), .ZN(n504) );
  AND2_X1 U389 ( .A1(n406), .A2(n405), .ZN(n404) );
  XNOR2_X1 U390 ( .A(n472), .B(n394), .ZN(n665) );
  XNOR2_X1 U391 ( .A(n364), .B(n363), .ZN(n476) );
  XNOR2_X1 U392 ( .A(n365), .B(KEYINPUT3), .ZN(n364) );
  XNOR2_X1 U393 ( .A(n400), .B(G146), .ZN(n434) );
  XNOR2_X1 U394 ( .A(G143), .B(G128), .ZN(n451) );
  XNOR2_X1 U395 ( .A(G101), .B(G113), .ZN(n363) );
  NAND2_X2 U396 ( .A1(n404), .A2(n401), .ZN(n639) );
  XNOR2_X1 U397 ( .A(n391), .B(KEYINPUT108), .ZN(n547) );
  NAND2_X1 U398 ( .A1(n549), .A2(n358), .ZN(n391) );
  XOR2_X1 U399 ( .A(KEYINPUT10), .B(n434), .Z(n468) );
  NOR2_X1 U400 ( .A1(G237), .A2(G953), .ZN(n439) );
  XNOR2_X1 U401 ( .A(n587), .B(n586), .ZN(n390) );
  XNOR2_X1 U402 ( .A(KEYINPUT85), .B(KEYINPUT48), .ZN(n586) );
  INV_X1 U403 ( .A(G237), .ZN(n419) );
  XNOR2_X1 U404 ( .A(n379), .B(KEYINPUT71), .ZN(n566) );
  NAND2_X1 U405 ( .A1(n392), .A2(n574), .ZN(n379) );
  AND2_X1 U406 ( .A1(n665), .A2(n393), .ZN(n392) );
  NOR2_X1 U407 ( .A1(G902), .A2(n697), .ZN(n526) );
  NAND2_X1 U408 ( .A1(n639), .A2(n431), .ZN(n374) );
  AND2_X1 U409 ( .A1(n513), .A2(n512), .ZN(n518) );
  AND2_X1 U410 ( .A1(n540), .A2(KEYINPUT64), .ZN(n511) );
  XOR2_X1 U411 ( .A(G137), .B(KEYINPUT99), .Z(n478) );
  XNOR2_X1 U412 ( .A(n475), .B(n474), .ZN(n729) );
  XOR2_X1 U413 ( .A(n467), .B(KEYINPUT70), .Z(n490) );
  XNOR2_X1 U414 ( .A(G137), .B(G140), .ZN(n467) );
  XNOR2_X1 U415 ( .A(n729), .B(G146), .ZN(n496) );
  INV_X1 U416 ( .A(G125), .ZN(n400) );
  XNOR2_X1 U417 ( .A(n395), .B(KEYINPUT79), .ZN(n574) );
  NOR2_X1 U418 ( .A1(n551), .A2(n550), .ZN(n395) );
  XNOR2_X1 U419 ( .A(n381), .B(KEYINPUT97), .ZN(n380) );
  XNOR2_X1 U420 ( .A(G119), .B(G110), .ZN(n381) );
  XNOR2_X1 U421 ( .A(n384), .B(n383), .ZN(n382) );
  XNOR2_X1 U422 ( .A(KEYINPUT24), .B(G128), .ZN(n384) );
  XNOR2_X1 U423 ( .A(KEYINPUT23), .B(KEYINPUT96), .ZN(n383) );
  XNOR2_X1 U424 ( .A(n443), .B(n442), .ZN(n703) );
  XNOR2_X1 U425 ( .A(n441), .B(n440), .ZN(n442) );
  AND2_X2 U426 ( .A1(n357), .A2(n366), .ZN(n702) );
  AND2_X1 U427 ( .A1(n390), .A2(n596), .ZN(n735) );
  INV_X1 U428 ( .A(KEYINPUT19), .ZN(n402) );
  NAND2_X1 U429 ( .A1(n424), .A2(KEYINPUT19), .ZN(n405) );
  INV_X1 U430 ( .A(n553), .ZN(n403) );
  XNOR2_X1 U431 ( .A(n526), .B(n353), .ZN(n589) );
  XNOR2_X1 U432 ( .A(n471), .B(n473), .ZN(n394) );
  NAND2_X1 U433 ( .A1(n371), .A2(n370), .ZN(n369) );
  INV_X1 U434 ( .A(n629), .ZN(n370) );
  INV_X1 U435 ( .A(n682), .ZN(n372) );
  INV_X1 U436 ( .A(KEYINPUT104), .ZN(n368) );
  XNOR2_X1 U437 ( .A(G143), .B(G113), .ZN(n432) );
  XNOR2_X1 U438 ( .A(n492), .B(n491), .ZN(n493) );
  INV_X1 U439 ( .A(G104), .ZN(n491) );
  XNOR2_X1 U440 ( .A(n386), .B(KEYINPUT75), .ZN(n523) );
  XNOR2_X1 U441 ( .A(n399), .B(n398), .ZN(n623) );
  INV_X1 U442 ( .A(n496), .ZN(n398) );
  XNOR2_X1 U443 ( .A(n479), .B(n485), .ZN(n399) );
  XOR2_X1 U444 ( .A(G122), .B(G104), .Z(n438) );
  XNOR2_X1 U445 ( .A(n496), .B(n387), .ZN(n697) );
  XNOR2_X1 U446 ( .A(n389), .B(n388), .ZN(n387) );
  XNOR2_X1 U447 ( .A(n493), .B(G101), .ZN(n388) );
  XNOR2_X1 U448 ( .A(n495), .B(n490), .ZN(n389) );
  XNOR2_X1 U449 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n413) );
  XNOR2_X1 U450 ( .A(n377), .B(KEYINPUT83), .ZN(n385) );
  NAND2_X1 U451 ( .A1(n390), .A2(n607), .ZN(n377) );
  XNOR2_X1 U452 ( .A(n428), .B(n429), .ZN(n549) );
  NAND2_X1 U453 ( .A1(n351), .A2(n397), .ZN(n396) );
  AND2_X1 U454 ( .A1(n552), .A2(n679), .ZN(n397) );
  XNOR2_X1 U455 ( .A(n378), .B(KEYINPUT28), .ZN(n557) );
  BUF_X1 U456 ( .A(n504), .Z(n530) );
  XNOR2_X1 U457 ( .A(n382), .B(n380), .ZN(n466) );
  XNOR2_X1 U458 ( .A(n703), .B(n407), .ZN(n704) );
  AND2_X1 U459 ( .A1(n613), .A2(G953), .ZN(n718) );
  NAND2_X1 U460 ( .A1(n534), .A2(n356), .ZN(n376) );
  NAND2_X1 U461 ( .A1(n403), .A2(n359), .ZN(n401) );
  AND2_X1 U462 ( .A1(n534), .A2(n665), .ZN(n501) );
  NOR2_X1 U463 ( .A1(n521), .A2(n520), .ZN(n350) );
  XOR2_X1 U464 ( .A(n546), .B(KEYINPUT30), .Z(n351) );
  NOR2_X1 U465 ( .A1(n530), .A2(n529), .ZN(n352) );
  XOR2_X1 U466 ( .A(n525), .B(KEYINPUT1), .Z(n353) );
  OR2_X1 U467 ( .A1(n521), .A2(n507), .ZN(n354) );
  NOR2_X1 U468 ( .A1(n589), .A2(n556), .ZN(n355) );
  AND2_X1 U469 ( .A1(n499), .A2(n665), .ZN(n356) );
  NAND2_X1 U470 ( .A1(n655), .A2(n385), .ZN(n357) );
  AND2_X1 U471 ( .A1(G953), .A2(G902), .ZN(n358) );
  AND2_X1 U472 ( .A1(n678), .A2(n402), .ZN(n359) );
  XOR2_X1 U473 ( .A(KEYINPUT84), .B(KEYINPUT35), .Z(n360) );
  XOR2_X1 U474 ( .A(n699), .B(n698), .Z(n361) );
  AND2_X1 U475 ( .A1(n604), .A2(n603), .ZN(n362) );
  NAND2_X1 U476 ( .A1(n367), .A2(n362), .ZN(n366) );
  NAND2_X1 U477 ( .A1(n655), .A2(n598), .ZN(n367) );
  XNOR2_X2 U478 ( .A(n545), .B(n544), .ZN(n655) );
  NAND2_X1 U479 ( .A1(n373), .A2(n372), .ZN(n371) );
  OR2_X1 U480 ( .A1(n646), .A2(n352), .ZN(n373) );
  NAND2_X1 U481 ( .A1(n566), .A2(n556), .ZN(n378) );
  INV_X1 U482 ( .A(n589), .ZN(n661) );
  NAND2_X1 U483 ( .A1(n527), .A2(n589), .ZN(n386) );
  INV_X1 U484 ( .A(n666), .ZN(n393) );
  NAND2_X1 U485 ( .A1(n595), .A2(n644), .ZN(n555) );
  NAND2_X1 U486 ( .A1(n403), .A2(n678), .ZN(n567) );
  NAND2_X1 U487 ( .A1(n553), .A2(KEYINPUT19), .ZN(n406) );
  XNOR2_X1 U488 ( .A(n700), .B(n361), .ZN(n701) );
  NAND2_X1 U489 ( .A1(n712), .A2(G469), .ZN(n700) );
  XNOR2_X1 U490 ( .A(n714), .B(n713), .ZN(n715) );
  BUF_X1 U491 ( .A(n553), .Z(n593) );
  XNOR2_X1 U492 ( .A(KEYINPUT59), .B(KEYINPUT65), .ZN(n407) );
  XNOR2_X1 U493 ( .A(n561), .B(KEYINPUT86), .ZN(n562) );
  XNOR2_X1 U494 ( .A(G131), .B(KEYINPUT12), .ZN(n435) );
  XNOR2_X1 U495 ( .A(n468), .B(n435), .ZN(n436) );
  XNOR2_X1 U496 ( .A(n484), .B(n483), .ZN(n485) );
  XNOR2_X1 U497 ( .A(n445), .B(n444), .ZN(n521) );
  XNOR2_X1 U498 ( .A(n555), .B(n554), .ZN(n741) );
  XNOR2_X1 U499 ( .A(n716), .B(n715), .ZN(n717) );
  XNOR2_X1 U500 ( .A(n494), .B(n450), .ZN(n408) );
  XNOR2_X1 U501 ( .A(n408), .B(n476), .ZN(n410) );
  XOR2_X1 U502 ( .A(KEYINPUT16), .B(n438), .Z(n409) );
  XNOR2_X1 U503 ( .A(n410), .B(n409), .ZN(n719) );
  INV_X1 U504 ( .A(KEYINPUT4), .ZN(n411) );
  XNOR2_X1 U505 ( .A(n451), .B(n411), .ZN(n475) );
  NAND2_X1 U506 ( .A1(n737), .A2(G224), .ZN(n412) );
  XNOR2_X1 U507 ( .A(n412), .B(KEYINPUT93), .ZN(n415) );
  XNOR2_X1 U508 ( .A(n434), .B(n413), .ZN(n414) );
  XNOR2_X1 U509 ( .A(n415), .B(n414), .ZN(n416) );
  XNOR2_X1 U510 ( .A(n475), .B(n416), .ZN(n417) );
  XNOR2_X1 U511 ( .A(n719), .B(n417), .ZN(n610) );
  XNOR2_X1 U512 ( .A(G902), .B(KEYINPUT92), .ZN(n418) );
  XNOR2_X1 U513 ( .A(n418), .B(KEYINPUT15), .ZN(n601) );
  NAND2_X1 U514 ( .A1(n610), .A2(n601), .ZN(n422) );
  INV_X1 U515 ( .A(G902), .ZN(n486) );
  NAND2_X1 U516 ( .A1(n486), .A2(n419), .ZN(n423) );
  NAND2_X1 U517 ( .A1(n423), .A2(G210), .ZN(n420) );
  XNOR2_X1 U518 ( .A(n420), .B(KEYINPUT94), .ZN(n421) );
  NAND2_X1 U519 ( .A1(n423), .A2(G214), .ZN(n678) );
  INV_X1 U520 ( .A(n678), .ZN(n424) );
  NOR2_X1 U521 ( .A1(G898), .A2(n737), .ZN(n720) );
  NAND2_X1 U522 ( .A1(n720), .A2(G902), .ZN(n426) );
  NAND2_X1 U523 ( .A1(n737), .A2(G952), .ZN(n425) );
  NAND2_X1 U524 ( .A1(n426), .A2(n425), .ZN(n430) );
  XOR2_X1 U525 ( .A(KEYINPUT95), .B(KEYINPUT14), .Z(n429) );
  NAND2_X1 U526 ( .A1(G234), .A2(G237), .ZN(n427) );
  XNOR2_X1 U527 ( .A(n427), .B(KEYINPUT74), .ZN(n428) );
  AND2_X1 U528 ( .A1(n430), .A2(n549), .ZN(n431) );
  INV_X1 U529 ( .A(n504), .ZN(n461) );
  XOR2_X1 U530 ( .A(KEYINPUT11), .B(KEYINPUT102), .Z(n433) );
  XNOR2_X1 U531 ( .A(n433), .B(n432), .ZN(n437) );
  XOR2_X1 U532 ( .A(n437), .B(n436), .Z(n443) );
  XNOR2_X1 U533 ( .A(n438), .B(G140), .ZN(n441) );
  XNOR2_X1 U534 ( .A(n439), .B(KEYINPUT78), .ZN(n482) );
  NAND2_X1 U535 ( .A1(G214), .A2(n482), .ZN(n440) );
  NOR2_X1 U536 ( .A1(G902), .A2(n703), .ZN(n445) );
  XNOR2_X1 U537 ( .A(KEYINPUT13), .B(G475), .ZN(n444) );
  XOR2_X1 U538 ( .A(G122), .B(KEYINPUT9), .Z(n449) );
  NAND2_X1 U539 ( .A1(n737), .A2(G234), .ZN(n447) );
  XNOR2_X1 U540 ( .A(KEYINPUT69), .B(KEYINPUT8), .ZN(n446) );
  XNOR2_X1 U541 ( .A(n447), .B(n446), .ZN(n464) );
  NAND2_X1 U542 ( .A1(G217), .A2(n464), .ZN(n448) );
  XNOR2_X1 U543 ( .A(n449), .B(n448), .ZN(n455) );
  XOR2_X1 U544 ( .A(KEYINPUT7), .B(n450), .Z(n453) );
  XOR2_X1 U545 ( .A(n451), .B(G134), .Z(n452) );
  XNOR2_X1 U546 ( .A(n453), .B(n452), .ZN(n454) );
  XNOR2_X1 U547 ( .A(n455), .B(n454), .ZN(n709) );
  NOR2_X1 U548 ( .A1(G902), .A2(n709), .ZN(n456) );
  XNOR2_X1 U549 ( .A(G478), .B(n456), .ZN(n520) );
  INV_X1 U550 ( .A(n520), .ZN(n507) );
  NAND2_X1 U551 ( .A1(G234), .A2(n601), .ZN(n457) );
  XNOR2_X1 U552 ( .A(n457), .B(KEYINPUT20), .ZN(n470) );
  AND2_X1 U553 ( .A1(n470), .A2(G221), .ZN(n459) );
  INV_X1 U554 ( .A(KEYINPUT21), .ZN(n458) );
  XNOR2_X1 U555 ( .A(n459), .B(n458), .ZN(n666) );
  NOR2_X1 U556 ( .A1(n354), .A2(n666), .ZN(n460) );
  NAND2_X1 U557 ( .A1(n461), .A2(n460), .ZN(n463) );
  INV_X1 U558 ( .A(KEYINPUT22), .ZN(n462) );
  NAND2_X1 U559 ( .A1(G221), .A2(n464), .ZN(n465) );
  XNOR2_X1 U560 ( .A(n466), .B(n465), .ZN(n469) );
  XNOR2_X1 U561 ( .A(n468), .B(n490), .ZN(n728) );
  XNOR2_X1 U562 ( .A(n469), .B(n728), .ZN(n714) );
  NOR2_X1 U563 ( .A1(G902), .A2(n714), .ZN(n472) );
  NAND2_X1 U564 ( .A1(n470), .A2(G217), .ZN(n471) );
  INV_X1 U565 ( .A(KEYINPUT25), .ZN(n473) );
  XNOR2_X1 U566 ( .A(G131), .B(G134), .ZN(n474) );
  XNOR2_X1 U567 ( .A(G116), .B(n476), .ZN(n477) );
  XNOR2_X1 U568 ( .A(n478), .B(n477), .ZN(n479) );
  XOR2_X1 U569 ( .A(KEYINPUT100), .B(KEYINPUT98), .Z(n481) );
  XNOR2_X1 U570 ( .A(KEYINPUT76), .B(KEYINPUT5), .ZN(n480) );
  XOR2_X1 U571 ( .A(n481), .B(n480), .Z(n484) );
  NAND2_X1 U572 ( .A1(G210), .A2(n482), .ZN(n483) );
  NAND2_X1 U573 ( .A1(n623), .A2(n486), .ZN(n488) );
  XOR2_X1 U574 ( .A(G472), .B(KEYINPUT101), .Z(n487) );
  XNOR2_X2 U575 ( .A(n488), .B(n487), .ZN(n522) );
  INV_X1 U576 ( .A(KEYINPUT6), .ZN(n489) );
  XNOR2_X1 U577 ( .A(n522), .B(n489), .ZN(n564) );
  INV_X1 U578 ( .A(n564), .ZN(n498) );
  NAND2_X1 U579 ( .A1(G227), .A2(n737), .ZN(n492) );
  XNOR2_X1 U580 ( .A(n494), .B(G107), .ZN(n495) );
  XNOR2_X1 U581 ( .A(KEYINPUT72), .B(G469), .ZN(n525) );
  INV_X1 U582 ( .A(KEYINPUT90), .ZN(n497) );
  XNOR2_X1 U583 ( .A(n661), .B(n497), .ZN(n569) );
  AND2_X1 U584 ( .A1(n498), .A2(n569), .ZN(n499) );
  INV_X1 U585 ( .A(KEYINPUT105), .ZN(n500) );
  XNOR2_X1 U586 ( .A(n522), .B(n500), .ZN(n556) );
  NAND2_X1 U587 ( .A1(n501), .A2(n355), .ZN(n634) );
  NOR2_X1 U588 ( .A1(n666), .A2(n665), .ZN(n527) );
  XOR2_X1 U589 ( .A(KEYINPUT106), .B(KEYINPUT33), .Z(n502) );
  XNOR2_X2 U590 ( .A(n503), .B(n502), .ZN(n687) );
  NOR2_X1 U591 ( .A1(n687), .A2(n530), .ZN(n506) );
  XNOR2_X1 U592 ( .A(KEYINPUT73), .B(KEYINPUT34), .ZN(n505) );
  XNOR2_X1 U593 ( .A(n506), .B(n505), .ZN(n509) );
  NAND2_X1 U594 ( .A1(n507), .A2(n521), .ZN(n508) );
  XOR2_X1 U595 ( .A(KEYINPUT107), .B(n508), .Z(n578) );
  XNOR2_X2 U596 ( .A(n510), .B(n360), .ZN(n538) );
  NAND2_X1 U597 ( .A1(n511), .A2(n538), .ZN(n513) );
  OR2_X1 U598 ( .A1(n514), .A2(KEYINPUT44), .ZN(n512) );
  INV_X1 U599 ( .A(KEYINPUT64), .ZN(n514) );
  NAND2_X1 U600 ( .A1(n514), .A2(KEYINPUT44), .ZN(n515) );
  NOR2_X1 U601 ( .A1(n515), .A2(n540), .ZN(n516) );
  NAND2_X1 U602 ( .A1(n538), .A2(n516), .ZN(n517) );
  NAND2_X1 U603 ( .A1(n518), .A2(n517), .ZN(n536) );
  NAND2_X1 U604 ( .A1(n520), .A2(n521), .ZN(n519) );
  XNOR2_X1 U605 ( .A(n519), .B(KEYINPUT103), .ZN(n644) );
  NOR2_X1 U606 ( .A1(n644), .A2(n350), .ZN(n682) );
  NAND2_X1 U607 ( .A1(n523), .A2(n522), .ZN(n672) );
  NOR2_X1 U608 ( .A1(n672), .A2(n530), .ZN(n524) );
  XOR2_X1 U609 ( .A(KEYINPUT31), .B(n524), .Z(n646) );
  XNOR2_X1 U610 ( .A(n526), .B(n525), .ZN(n558) );
  INV_X1 U611 ( .A(n527), .ZN(n662) );
  NOR2_X1 U612 ( .A1(n558), .A2(n662), .ZN(n576) );
  INV_X1 U613 ( .A(n522), .ZN(n528) );
  NAND2_X1 U614 ( .A1(n576), .A2(n528), .ZN(n529) );
  INV_X1 U615 ( .A(n665), .ZN(n531) );
  NAND2_X1 U616 ( .A1(n661), .A2(n531), .ZN(n532) );
  NOR2_X1 U617 ( .A1(n564), .A2(n532), .ZN(n533) );
  AND2_X1 U618 ( .A1(n534), .A2(n533), .ZN(n629) );
  NAND2_X1 U619 ( .A1(n536), .A2(n535), .ZN(n537) );
  XNOR2_X1 U620 ( .A(n537), .B(KEYINPUT87), .ZN(n543) );
  INV_X1 U621 ( .A(n538), .ZN(n743) );
  NOR2_X1 U622 ( .A1(n743), .A2(KEYINPUT44), .ZN(n539) );
  XNOR2_X1 U623 ( .A(n539), .B(KEYINPUT68), .ZN(n541) );
  NAND2_X1 U624 ( .A1(n541), .A2(n540), .ZN(n542) );
  NAND2_X1 U625 ( .A1(n543), .A2(n542), .ZN(n545) );
  XNOR2_X1 U626 ( .A(KEYINPUT82), .B(KEYINPUT45), .ZN(n544) );
  NAND2_X1 U627 ( .A1(n556), .A2(n678), .ZN(n546) );
  NOR2_X1 U628 ( .A1(G900), .A2(n547), .ZN(n548) );
  XOR2_X1 U629 ( .A(KEYINPUT109), .B(n548), .Z(n551) );
  NAND2_X1 U630 ( .A1(G952), .A2(n549), .ZN(n693) );
  NOR2_X1 U631 ( .A1(G953), .A2(n693), .ZN(n550) );
  AND2_X1 U632 ( .A1(n574), .A2(n576), .ZN(n552) );
  XNOR2_X1 U633 ( .A(n593), .B(KEYINPUT38), .ZN(n679) );
  XOR2_X1 U634 ( .A(KEYINPUT111), .B(KEYINPUT40), .Z(n554) );
  NOR2_X1 U635 ( .A1(n558), .A2(n557), .ZN(n635) );
  NAND2_X1 U636 ( .A1(n679), .A2(n678), .ZN(n683) );
  NOR2_X1 U637 ( .A1(n354), .A2(n683), .ZN(n559) );
  XOR2_X1 U638 ( .A(KEYINPUT41), .B(n559), .Z(n653) );
  NAND2_X1 U639 ( .A1(n635), .A2(n653), .ZN(n560) );
  XNOR2_X1 U640 ( .A(n560), .B(KEYINPUT42), .ZN(n742) );
  NAND2_X1 U641 ( .A1(n741), .A2(n742), .ZN(n563) );
  INV_X1 U642 ( .A(KEYINPUT46), .ZN(n561) );
  XNOR2_X1 U643 ( .A(n563), .B(n562), .ZN(n585) );
  AND2_X1 U644 ( .A1(n564), .A2(n644), .ZN(n565) );
  NAND2_X1 U645 ( .A1(n566), .A2(n565), .ZN(n588) );
  NOR2_X1 U646 ( .A1(n588), .A2(n567), .ZN(n568) );
  XNOR2_X1 U647 ( .A(n568), .B(KEYINPUT36), .ZN(n570) );
  NAND2_X1 U648 ( .A1(n570), .A2(n569), .ZN(n649) );
  INV_X1 U649 ( .A(n649), .ZN(n583) );
  INV_X1 U650 ( .A(n639), .ZN(n571) );
  NOR2_X1 U651 ( .A1(n571), .A2(n682), .ZN(n572) );
  NAND2_X1 U652 ( .A1(n635), .A2(n572), .ZN(n573) );
  XOR2_X1 U653 ( .A(KEYINPUT47), .B(n573), .Z(n581) );
  AND2_X1 U654 ( .A1(n351), .A2(n574), .ZN(n575) );
  NAND2_X1 U655 ( .A1(n576), .A2(n575), .ZN(n577) );
  NOR2_X1 U656 ( .A1(n578), .A2(n577), .ZN(n580) );
  INV_X1 U657 ( .A(n593), .ZN(n579) );
  NAND2_X1 U658 ( .A1(n580), .A2(n579), .ZN(n616) );
  NAND2_X1 U659 ( .A1(n581), .A2(n616), .ZN(n582) );
  NOR2_X1 U660 ( .A1(n583), .A2(n582), .ZN(n584) );
  NAND2_X1 U661 ( .A1(n585), .A2(n584), .ZN(n587) );
  NOR2_X1 U662 ( .A1(n589), .A2(n588), .ZN(n590) );
  NAND2_X1 U663 ( .A1(n678), .A2(n590), .ZN(n591) );
  XNOR2_X1 U664 ( .A(n591), .B(KEYINPUT43), .ZN(n592) );
  XNOR2_X1 U665 ( .A(KEYINPUT110), .B(n592), .ZN(n594) );
  NAND2_X1 U666 ( .A1(n594), .A2(n593), .ZN(n618) );
  NAND2_X1 U667 ( .A1(n595), .A2(n350), .ZN(n652) );
  AND2_X1 U668 ( .A1(n618), .A2(n652), .ZN(n596) );
  INV_X1 U669 ( .A(n601), .ZN(n597) );
  AND2_X1 U670 ( .A1(n735), .A2(n597), .ZN(n598) );
  NAND2_X1 U671 ( .A1(KEYINPUT66), .A2(KEYINPUT2), .ZN(n599) );
  OR2_X1 U672 ( .A1(n601), .A2(n599), .ZN(n604) );
  INV_X1 U673 ( .A(KEYINPUT2), .ZN(n600) );
  NOR2_X1 U674 ( .A1(n601), .A2(n600), .ZN(n602) );
  OR2_X1 U675 ( .A1(n602), .A2(KEYINPUT66), .ZN(n603) );
  NAND2_X1 U676 ( .A1(KEYINPUT2), .A2(n652), .ZN(n605) );
  XOR2_X1 U677 ( .A(KEYINPUT80), .B(n605), .Z(n606) );
  AND2_X1 U678 ( .A1(n618), .A2(n606), .ZN(n607) );
  NAND2_X1 U679 ( .A1(n702), .A2(G210), .ZN(n612) );
  XNOR2_X1 U680 ( .A(KEYINPUT55), .B(KEYINPUT88), .ZN(n608) );
  XNOR2_X1 U681 ( .A(n608), .B(KEYINPUT54), .ZN(n609) );
  XNOR2_X1 U682 ( .A(n610), .B(n609), .ZN(n611) );
  XNOR2_X1 U683 ( .A(n612), .B(n611), .ZN(n614) );
  INV_X1 U684 ( .A(G952), .ZN(n613) );
  XNOR2_X1 U685 ( .A(n615), .B(KEYINPUT56), .ZN(G51) );
  XNOR2_X1 U686 ( .A(n616), .B(G143), .ZN(G45) );
  XNOR2_X1 U687 ( .A(G140), .B(KEYINPUT116), .ZN(n617) );
  XNOR2_X1 U688 ( .A(n618), .B(n617), .ZN(G42) );
  BUF_X1 U689 ( .A(n619), .Z(n620) );
  XNOR2_X1 U690 ( .A(n620), .B(G119), .ZN(G21) );
  NAND2_X1 U691 ( .A1(n702), .A2(G472), .ZN(n625) );
  XNOR2_X1 U692 ( .A(KEYINPUT89), .B(KEYINPUT112), .ZN(n621) );
  XNOR2_X1 U693 ( .A(n621), .B(KEYINPUT62), .ZN(n622) );
  XNOR2_X1 U694 ( .A(n623), .B(n622), .ZN(n624) );
  XNOR2_X1 U695 ( .A(n625), .B(n624), .ZN(n626) );
  XNOR2_X1 U696 ( .A(KEYINPUT91), .B(KEYINPUT63), .ZN(n627) );
  XNOR2_X1 U697 ( .A(n628), .B(n627), .ZN(G57) );
  XOR2_X1 U698 ( .A(G101), .B(n629), .Z(G3) );
  NAND2_X1 U699 ( .A1(n352), .A2(n644), .ZN(n630) );
  XNOR2_X1 U700 ( .A(n630), .B(G104), .ZN(G6) );
  XOR2_X1 U701 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n632) );
  NAND2_X1 U702 ( .A1(n352), .A2(n350), .ZN(n631) );
  XNOR2_X1 U703 ( .A(n632), .B(n631), .ZN(n633) );
  XNOR2_X1 U704 ( .A(G107), .B(n633), .ZN(G9) );
  XNOR2_X1 U705 ( .A(G110), .B(n634), .ZN(G12) );
  INV_X1 U706 ( .A(n635), .ZN(n641) );
  NAND2_X1 U707 ( .A1(n350), .A2(n639), .ZN(n636) );
  NOR2_X1 U708 ( .A1(n641), .A2(n636), .ZN(n638) );
  XNOR2_X1 U709 ( .A(G128), .B(KEYINPUT29), .ZN(n637) );
  XNOR2_X1 U710 ( .A(n638), .B(n637), .ZN(G30) );
  NAND2_X1 U711 ( .A1(n644), .A2(n639), .ZN(n640) );
  NOR2_X1 U712 ( .A1(n641), .A2(n640), .ZN(n643) );
  XNOR2_X1 U713 ( .A(G146), .B(KEYINPUT113), .ZN(n642) );
  XNOR2_X1 U714 ( .A(n643), .B(n642), .ZN(G48) );
  NAND2_X1 U715 ( .A1(n646), .A2(n644), .ZN(n645) );
  XNOR2_X1 U716 ( .A(n645), .B(G113), .ZN(G15) );
  NAND2_X1 U717 ( .A1(n646), .A2(n350), .ZN(n647) );
  XNOR2_X1 U718 ( .A(n647), .B(KEYINPUT114), .ZN(n648) );
  XNOR2_X1 U719 ( .A(G116), .B(n648), .ZN(G18) );
  XNOR2_X1 U720 ( .A(KEYINPUT37), .B(KEYINPUT115), .ZN(n650) );
  XNOR2_X1 U721 ( .A(n650), .B(n649), .ZN(n651) );
  XNOR2_X1 U722 ( .A(G125), .B(n651), .ZN(G27) );
  XNOR2_X1 U723 ( .A(G134), .B(n652), .ZN(G36) );
  INV_X1 U724 ( .A(n653), .ZN(n676) );
  NOR2_X1 U725 ( .A1(n687), .A2(n676), .ZN(n654) );
  NOR2_X1 U726 ( .A1(G953), .A2(n654), .ZN(n660) );
  NAND2_X1 U727 ( .A1(n735), .A2(n655), .ZN(n657) );
  XNOR2_X1 U728 ( .A(KEYINPUT81), .B(KEYINPUT2), .ZN(n656) );
  NAND2_X1 U729 ( .A1(n657), .A2(n656), .ZN(n658) );
  NAND2_X1 U730 ( .A1(n357), .A2(n658), .ZN(n659) );
  NAND2_X1 U731 ( .A1(n660), .A2(n659), .ZN(n695) );
  NAND2_X1 U732 ( .A1(n662), .A2(n661), .ZN(n663) );
  XNOR2_X1 U733 ( .A(n663), .B(KEYINPUT50), .ZN(n664) );
  XNOR2_X1 U734 ( .A(n664), .B(KEYINPUT118), .ZN(n671) );
  NAND2_X1 U735 ( .A1(n666), .A2(n665), .ZN(n667) );
  XNOR2_X1 U736 ( .A(KEYINPUT49), .B(n667), .ZN(n668) );
  NOR2_X1 U737 ( .A1(n522), .A2(n668), .ZN(n669) );
  XOR2_X1 U738 ( .A(KEYINPUT117), .B(n669), .Z(n670) );
  NAND2_X1 U739 ( .A1(n671), .A2(n670), .ZN(n673) );
  NAND2_X1 U740 ( .A1(n673), .A2(n672), .ZN(n675) );
  XOR2_X1 U741 ( .A(KEYINPUT51), .B(KEYINPUT119), .Z(n674) );
  XNOR2_X1 U742 ( .A(n675), .B(n674), .ZN(n677) );
  NOR2_X1 U743 ( .A1(n677), .A2(n676), .ZN(n689) );
  NOR2_X1 U744 ( .A1(n679), .A2(n678), .ZN(n680) );
  NOR2_X1 U745 ( .A1(n354), .A2(n680), .ZN(n681) );
  XNOR2_X1 U746 ( .A(n681), .B(KEYINPUT120), .ZN(n685) );
  NOR2_X1 U747 ( .A1(n683), .A2(n682), .ZN(n684) );
  NOR2_X1 U748 ( .A1(n685), .A2(n684), .ZN(n686) );
  NOR2_X1 U749 ( .A1(n687), .A2(n686), .ZN(n688) );
  NOR2_X1 U750 ( .A1(n689), .A2(n688), .ZN(n690) );
  XOR2_X1 U751 ( .A(n690), .B(KEYINPUT121), .Z(n691) );
  XNOR2_X1 U752 ( .A(KEYINPUT52), .B(n691), .ZN(n692) );
  NOR2_X1 U753 ( .A1(n693), .A2(n692), .ZN(n694) );
  NOR2_X1 U754 ( .A1(n695), .A2(n694), .ZN(n696) );
  XNOR2_X1 U755 ( .A(n696), .B(KEYINPUT53), .ZN(G75) );
  XNOR2_X1 U756 ( .A(KEYINPUT58), .B(KEYINPUT122), .ZN(n699) );
  XNOR2_X1 U757 ( .A(n697), .B(KEYINPUT57), .ZN(n698) );
  NOR2_X1 U758 ( .A1(n718), .A2(n701), .ZN(G54) );
  NAND2_X1 U759 ( .A1(n702), .A2(G475), .ZN(n705) );
  XNOR2_X1 U760 ( .A(n705), .B(n704), .ZN(n706) );
  XOR2_X1 U761 ( .A(KEYINPUT67), .B(KEYINPUT60), .Z(n707) );
  XNOR2_X1 U762 ( .A(n708), .B(n707), .ZN(G60) );
  NAND2_X1 U763 ( .A1(n712), .A2(G478), .ZN(n710) );
  XNOR2_X1 U764 ( .A(n710), .B(n709), .ZN(n711) );
  NOR2_X1 U765 ( .A1(n718), .A2(n711), .ZN(G63) );
  NAND2_X1 U766 ( .A1(n712), .A2(G217), .ZN(n716) );
  INV_X1 U767 ( .A(KEYINPUT123), .ZN(n713) );
  NOR2_X1 U768 ( .A1(n718), .A2(n717), .ZN(G66) );
  NOR2_X1 U769 ( .A1(n719), .A2(n720), .ZN(n727) );
  NAND2_X1 U770 ( .A1(n655), .A2(n737), .ZN(n725) );
  NAND2_X1 U771 ( .A1(G953), .A2(G224), .ZN(n721) );
  XNOR2_X1 U772 ( .A(KEYINPUT61), .B(n721), .ZN(n722) );
  NAND2_X1 U773 ( .A1(n722), .A2(G898), .ZN(n723) );
  XNOR2_X1 U774 ( .A(n723), .B(KEYINPUT124), .ZN(n724) );
  NAND2_X1 U775 ( .A1(n725), .A2(n724), .ZN(n726) );
  XNOR2_X1 U776 ( .A(n727), .B(n726), .ZN(G69) );
  XNOR2_X1 U777 ( .A(n729), .B(n728), .ZN(n736) );
  XNOR2_X1 U778 ( .A(n736), .B(G227), .ZN(n730) );
  XNOR2_X1 U779 ( .A(n730), .B(KEYINPUT125), .ZN(n731) );
  NAND2_X1 U780 ( .A1(n731), .A2(G900), .ZN(n732) );
  XOR2_X1 U781 ( .A(KEYINPUT126), .B(n732), .Z(n733) );
  NOR2_X1 U782 ( .A1(n737), .A2(n733), .ZN(n734) );
  XNOR2_X1 U783 ( .A(n734), .B(KEYINPUT127), .ZN(n740) );
  XNOR2_X1 U784 ( .A(n736), .B(n735), .ZN(n738) );
  NAND2_X1 U785 ( .A1(n738), .A2(n737), .ZN(n739) );
  NAND2_X1 U786 ( .A1(n740), .A2(n739), .ZN(G72) );
  XNOR2_X1 U787 ( .A(G131), .B(n741), .ZN(G33) );
  XNOR2_X1 U788 ( .A(G137), .B(n742), .ZN(G39) );
  XOR2_X1 U789 ( .A(G122), .B(n743), .Z(G24) );
endmodule

