

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352,
         n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
         n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
         n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
         n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396,
         n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407,
         n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418,
         n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429,
         n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440,
         n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451,
         n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462,
         n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473,
         n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484,
         n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495,
         n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506,
         n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517,
         n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583,
         n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594,
         n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605,
         n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616,
         n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627,
         n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638,
         n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649,
         n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660,
         n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671,
         n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682,
         n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693,
         n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704,
         n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715,
         n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726,
         n727, n728, n729, n730, n731, n732, n733, n734, n735, n736;

  NOR2_X1 U364 ( .A1(n541), .A2(n545), .ZN(n668) );
  INV_X1 U365 ( .A(n544), .ZN(n541) );
  XNOR2_X1 U366 ( .A(n457), .B(n456), .ZN(n552) );
  NOR2_X1 U367 ( .A1(n571), .A2(n639), .ZN(n349) );
  XNOR2_X1 U368 ( .A(n535), .B(KEYINPUT42), .ZN(n736) );
  NOR2_X2 U369 ( .A1(n706), .A2(n707), .ZN(n374) );
  XNOR2_X2 U370 ( .A(n413), .B(KEYINPUT33), .ZN(n665) );
  XNOR2_X2 U371 ( .A(G110), .B(G119), .ZN(n471) );
  XNOR2_X2 U372 ( .A(n366), .B(n589), .ZN(n732) );
  NAND2_X2 U373 ( .A1(n599), .A2(n588), .ZN(n366) );
  INV_X1 U374 ( .A(n734), .ZN(n352) );
  NOR2_X1 U375 ( .A1(n391), .A2(n736), .ZN(n420) );
  NOR2_X1 U376 ( .A1(n697), .A2(G902), .ZN(n511) );
  INV_X2 U377 ( .A(G953), .ZN(n727) );
  INV_X4 U378 ( .A(G125), .ZN(n354) );
  INV_X4 U379 ( .A(G128), .ZN(n357) );
  NOR2_X1 U380 ( .A1(n421), .A2(n418), .ZN(n563) );
  OR2_X1 U381 ( .A1(n650), .A2(n552), .ZN(n605) );
  NAND2_X1 U382 ( .A1(n388), .A2(n387), .ZN(n650) );
  OR2_X1 U383 ( .A1(n666), .A2(n667), .ZN(n534) );
  XNOR2_X1 U384 ( .A(n407), .B(G478), .ZN(n545) );
  XNOR2_X1 U385 ( .A(n483), .B(n482), .ZN(n590) );
  OR2_X1 U386 ( .A1(n702), .A2(G902), .ZN(n407) );
  XOR2_X1 U387 ( .A(n476), .B(n475), .Z(n705) );
  XNOR2_X1 U388 ( .A(n519), .B(n446), .ZN(n721) );
  XNOR2_X1 U389 ( .A(n520), .B(n469), .ZN(n503) );
  XNOR2_X1 U390 ( .A(n362), .B(n491), .ZN(n524) );
  XNOR2_X1 U391 ( .A(n363), .B(G113), .ZN(n362) );
  INV_X1 U392 ( .A(G101), .ZN(n363) );
  XNOR2_X1 U393 ( .A(G119), .B(KEYINPUT3), .ZN(n491) );
  NOR2_X1 U394 ( .A1(G953), .A2(G237), .ZN(n497) );
  XNOR2_X1 U395 ( .A(G137), .B(KEYINPUT66), .ZN(n470) );
  AND2_X1 U396 ( .A1(G227), .A2(n727), .ZN(n451) );
  NOR2_X1 U397 ( .A1(KEYINPUT44), .A2(KEYINPUT79), .ZN(n594) );
  XNOR2_X1 U398 ( .A(n468), .B(G140), .ZN(n469) );
  INV_X1 U399 ( .A(KEYINPUT10), .ZN(n468) );
  XNOR2_X1 U400 ( .A(n721), .B(G146), .ZN(n490) );
  NAND2_X1 U401 ( .A1(G237), .A2(G234), .ZN(n464) );
  AND2_X1 U402 ( .A1(n568), .A2(n378), .ZN(n557) );
  NOR2_X1 U403 ( .A1(n639), .A2(n556), .ZN(n564) );
  NOR2_X1 U404 ( .A1(n554), .A2(n553), .ZN(n555) );
  NOR2_X1 U405 ( .A1(n342), .A2(n644), .ZN(n424) );
  XOR2_X1 U406 ( .A(KEYINPUT11), .B(KEYINPUT95), .Z(n499) );
  XOR2_X1 U407 ( .A(KEYINPUT93), .B(KEYINPUT94), .Z(n496) );
  XNOR2_X1 U408 ( .A(KEYINPUT51), .B(KEYINPUT117), .ZN(n361) );
  INV_X1 U409 ( .A(KEYINPUT44), .ZN(n351) );
  XNOR2_X1 U410 ( .A(n568), .B(KEYINPUT38), .ZN(n666) );
  XNOR2_X1 U411 ( .A(n606), .B(KEYINPUT6), .ZN(n553) );
  XNOR2_X1 U412 ( .A(n573), .B(n385), .ZN(n602) );
  INV_X1 U413 ( .A(KEYINPUT70), .ZN(n385) );
  NOR2_X1 U414 ( .A1(n650), .A2(n572), .ZN(n573) );
  XNOR2_X1 U415 ( .A(n481), .B(n480), .ZN(n482) );
  XNOR2_X1 U416 ( .A(KEYINPUT21), .B(n461), .ZN(n655) );
  INV_X1 U417 ( .A(n553), .ZN(n587) );
  XNOR2_X1 U418 ( .A(n552), .B(KEYINPUT1), .ZN(n572) );
  XNOR2_X1 U419 ( .A(n489), .B(n395), .ZN(n394) );
  INV_X1 U420 ( .A(n524), .ZN(n395) );
  XNOR2_X1 U421 ( .A(G122), .B(G104), .ZN(n526) );
  INV_X1 U422 ( .A(KEYINPUT16), .ZN(n444) );
  INV_X1 U423 ( .A(KEYINPUT23), .ZN(n384) );
  XNOR2_X1 U424 ( .A(n503), .B(n367), .ZN(n719) );
  INV_X1 U425 ( .A(n470), .ZN(n367) );
  XNOR2_X1 U426 ( .A(n406), .B(G107), .ZN(n525) );
  INV_X1 U427 ( .A(G116), .ZN(n406) );
  XNOR2_X1 U428 ( .A(G122), .B(KEYINPUT98), .ZN(n405) );
  INV_X1 U429 ( .A(G134), .ZN(n447) );
  XNOR2_X1 U430 ( .A(KEYINPUT9), .B(KEYINPUT7), .ZN(n512) );
  XOR2_X1 U431 ( .A(KEYINPUT96), .B(KEYINPUT97), .Z(n513) );
  XNOR2_X1 U432 ( .A(n506), .B(n505), .ZN(n507) );
  INV_X1 U433 ( .A(G143), .ZN(n505) );
  XNOR2_X1 U434 ( .A(n714), .B(n437), .ZN(n689) );
  XNOR2_X1 U435 ( .A(n523), .B(n438), .ZN(n437) );
  XNOR2_X1 U436 ( .A(n521), .B(n439), .ZN(n438) );
  XNOR2_X1 U437 ( .A(n430), .B(n429), .ZN(n685) );
  INV_X1 U438 ( .A(KEYINPUT41), .ZN(n429) );
  INV_X1 U439 ( .A(n537), .ZN(n375) );
  XNOR2_X1 U440 ( .A(n557), .B(n343), .ZN(n576) );
  AND2_X1 U441 ( .A1(n426), .A2(n425), .ZN(n548) );
  XNOR2_X1 U442 ( .A(n493), .B(n372), .ZN(n426) );
  XNOR2_X1 U443 ( .A(n494), .B(n427), .ZN(n372) );
  INV_X1 U444 ( .A(n606), .ZN(n652) );
  OR2_X1 U445 ( .A1(n682), .A2(n404), .ZN(n403) );
  OR2_X1 U446 ( .A1(n620), .A2(n434), .ZN(n404) );
  AND2_X1 U447 ( .A1(n402), .A2(n401), .ZN(n400) );
  NAND2_X1 U448 ( .A1(n620), .A2(n434), .ZN(n402) );
  NAND2_X1 U449 ( .A1(n435), .A2(G475), .ZN(n432) );
  XNOR2_X1 U450 ( .A(n490), .B(n416), .ZN(n695) );
  XNOR2_X1 U451 ( .A(n417), .B(n450), .ZN(n416) );
  XNOR2_X1 U452 ( .A(n452), .B(n453), .ZN(n417) );
  NAND2_X1 U453 ( .A1(n435), .A2(G210), .ZN(n431) );
  INV_X1 U454 ( .A(KEYINPUT99), .ZN(n396) );
  XNOR2_X1 U455 ( .A(n670), .B(KEYINPUT74), .ZN(n609) );
  INV_X1 U456 ( .A(KEYINPUT46), .ZN(n419) );
  NAND2_X1 U457 ( .A1(n560), .A2(n559), .ZN(n423) );
  XNOR2_X1 U458 ( .A(n546), .B(n365), .ZN(n670) );
  INV_X1 U459 ( .A(KEYINPUT100), .ZN(n365) );
  AND2_X1 U460 ( .A1(n641), .A2(n639), .ZN(n546) );
  XNOR2_X1 U461 ( .A(n459), .B(n458), .ZN(n477) );
  XNOR2_X1 U462 ( .A(G137), .B(G116), .ZN(n485) );
  XOR2_X1 U463 ( .A(KEYINPUT71), .B(KEYINPUT5), .Z(n486) );
  XNOR2_X1 U464 ( .A(G131), .B(KEYINPUT12), .ZN(n495) );
  XOR2_X1 U465 ( .A(KEYINPUT4), .B(G131), .Z(n446) );
  XNOR2_X1 U466 ( .A(n441), .B(n440), .ZN(n439) );
  INV_X1 U467 ( .A(KEYINPUT17), .ZN(n440) );
  XNOR2_X1 U468 ( .A(KEYINPUT82), .B(KEYINPUT18), .ZN(n441) );
  INV_X1 U469 ( .A(KEYINPUT118), .ZN(n359) );
  XNOR2_X1 U470 ( .A(n662), .B(n361), .ZN(n663) );
  OR2_X1 U471 ( .A1(G902), .A2(G237), .ZN(n532) );
  INV_X1 U472 ( .A(n655), .ZN(n387) );
  INV_X1 U473 ( .A(n590), .ZN(n388) );
  NAND2_X1 U474 ( .A1(n435), .A2(G472), .ZN(n434) );
  NAND2_X1 U475 ( .A1(n373), .A2(n392), .ZN(n722) );
  XNOR2_X1 U476 ( .A(n393), .B(KEYINPUT77), .ZN(n373) );
  INV_X1 U477 ( .A(G104), .ZN(n448) );
  XNOR2_X1 U478 ( .A(n451), .B(G140), .ZN(n452) );
  XOR2_X1 U479 ( .A(G107), .B(G101), .Z(n453) );
  BUF_X1 U480 ( .A(n665), .Z(n683) );
  NOR2_X1 U481 ( .A1(n666), .A2(n542), .ZN(n540) );
  XNOR2_X1 U482 ( .A(n511), .B(n510), .ZN(n544) );
  INV_X1 U483 ( .A(KEYINPUT13), .ZN(n509) );
  BUF_X1 U484 ( .A(n590), .Z(n353) );
  OR2_X1 U485 ( .A1(n619), .A2(G902), .ZN(n492) );
  INV_X1 U486 ( .A(KEYINPUT0), .ZN(n355) );
  AND2_X1 U487 ( .A1(n577), .A2(n578), .ZN(n382) );
  XNOR2_X1 U488 ( .A(n442), .B(n527), .ZN(n714) );
  XNOR2_X1 U489 ( .A(n524), .B(n443), .ZN(n442) );
  XNOR2_X1 U490 ( .A(n526), .B(n444), .ZN(n443) );
  NAND2_X1 U491 ( .A1(n435), .A2(G217), .ZN(n433) );
  XNOR2_X1 U492 ( .A(n525), .B(n405), .ZN(n515) );
  BUF_X1 U493 ( .A(n685), .Z(n364) );
  AND2_X1 U494 ( .A1(n428), .A2(n548), .ZN(n535) );
  AND2_X1 U495 ( .A1(n350), .A2(n601), .ZN(n644) );
  XNOR2_X1 U496 ( .A(n558), .B(n344), .ZN(n350) );
  INV_X1 U497 ( .A(n580), .ZN(n410) );
  NOR2_X1 U498 ( .A1(n543), .A2(n580), .ZN(n635) );
  NOR2_X1 U499 ( .A1(n399), .A2(n398), .ZN(n621) );
  INV_X1 U500 ( .A(KEYINPUT60), .ZN(n370) );
  XNOR2_X1 U501 ( .A(n693), .B(n386), .ZN(n696) );
  XNOR2_X1 U502 ( .A(n695), .B(n694), .ZN(n386) );
  INV_X1 U503 ( .A(KEYINPUT56), .ZN(n368) );
  INV_X1 U504 ( .A(n639), .ZN(n636) );
  XNOR2_X1 U505 ( .A(KEYINPUT15), .B(G902), .ZN(n618) );
  INV_X1 U506 ( .A(n667), .ZN(n378) );
  NAND2_X1 U507 ( .A1(n551), .A2(n550), .ZN(n342) );
  INV_X1 U508 ( .A(n601), .ZN(n649) );
  XOR2_X1 U509 ( .A(KEYINPUT72), .B(KEYINPUT19), .Z(n343) );
  XOR2_X1 U510 ( .A(KEYINPUT80), .B(KEYINPUT36), .Z(n344) );
  XOR2_X1 U511 ( .A(KEYINPUT35), .B(KEYINPUT76), .Z(n345) );
  XOR2_X1 U512 ( .A(n699), .B(n698), .Z(n346) );
  XNOR2_X1 U513 ( .A(n691), .B(n690), .ZN(n347) );
  INV_X1 U514 ( .A(n618), .ZN(n435) );
  NOR2_X1 U515 ( .A1(G952), .A2(n727), .ZN(n707) );
  INV_X1 U516 ( .A(n707), .ZN(n401) );
  XNOR2_X1 U517 ( .A(n490), .B(n394), .ZN(n619) );
  NAND2_X1 U518 ( .A1(n348), .A2(n376), .ZN(n542) );
  AND2_X1 U519 ( .A1(n389), .A2(n375), .ZN(n348) );
  XNOR2_X1 U520 ( .A(n635), .B(KEYINPUT75), .ZN(n551) );
  NAND2_X1 U521 ( .A1(n477), .A2(G221), .ZN(n460) );
  XNOR2_X2 U522 ( .A(n349), .B(KEYINPUT40), .ZN(n391) );
  NAND2_X1 U523 ( .A1(n352), .A2(n351), .ZN(n597) );
  XNOR2_X2 U524 ( .A(n354), .B(G146), .ZN(n520) );
  XNOR2_X2 U525 ( .A(n356), .B(n355), .ZN(n584) );
  NAND2_X1 U526 ( .A1(n576), .A2(n382), .ZN(n356) );
  XNOR2_X2 U527 ( .A(n522), .B(n447), .ZN(n519) );
  XNOR2_X2 U528 ( .A(n357), .B(G143), .ZN(n522) );
  NAND2_X1 U529 ( .A1(n358), .A2(n675), .ZN(n676) );
  XNOR2_X1 U530 ( .A(n664), .B(n359), .ZN(n358) );
  XNOR2_X1 U531 ( .A(n360), .B(KEYINPUT53), .ZN(G75) );
  AND2_X1 U532 ( .A1(n688), .A2(n727), .ZN(n360) );
  OR2_X2 U533 ( .A1(n682), .A2(n433), .ZN(n704) );
  XNOR2_X1 U534 ( .A(n420), .B(n419), .ZN(n418) );
  INV_X1 U535 ( .A(n605), .ZN(n376) );
  XNOR2_X2 U536 ( .A(n531), .B(n530), .ZN(n568) );
  XNOR2_X1 U537 ( .A(n508), .B(n507), .ZN(n697) );
  XNOR2_X1 U538 ( .A(n390), .B(n538), .ZN(n389) );
  NAND2_X1 U539 ( .A1(n536), .A2(n541), .ZN(n397) );
  XNOR2_X1 U540 ( .A(n602), .B(n415), .ZN(n414) );
  XNOR2_X1 U541 ( .A(n369), .B(n368), .ZN(G51) );
  NAND2_X1 U542 ( .A1(n379), .A2(n401), .ZN(n369) );
  XNOR2_X1 U543 ( .A(n371), .B(n370), .ZN(G60) );
  NAND2_X1 U544 ( .A1(n380), .A2(n401), .ZN(n371) );
  XNOR2_X1 U545 ( .A(n374), .B(KEYINPUT122), .ZN(G66) );
  XNOR2_X1 U546 ( .A(n471), .B(n384), .ZN(n383) );
  XNOR2_X1 U547 ( .A(n383), .B(n472), .ZN(n473) );
  NAND2_X1 U548 ( .A1(n377), .A2(n597), .ZN(n614) );
  NAND2_X1 U549 ( .A1(n596), .A2(n734), .ZN(n377) );
  INV_X1 U550 ( .A(n568), .ZN(n547) );
  XNOR2_X1 U551 ( .A(n692), .B(n347), .ZN(n379) );
  XNOR2_X1 U552 ( .A(n616), .B(n615), .ZN(n708) );
  XNOR2_X1 U553 ( .A(n700), .B(n346), .ZN(n380) );
  XNOR2_X2 U554 ( .A(n381), .B(KEYINPUT2), .ZN(n682) );
  NOR2_X2 U555 ( .A1(n722), .A2(n617), .ZN(n381) );
  NAND2_X1 U556 ( .A1(n614), .A2(n613), .ZN(n616) );
  NOR2_X2 U557 ( .A1(n592), .A2(n587), .ZN(n599) );
  NAND2_X1 U558 ( .A1(n606), .A2(n378), .ZN(n390) );
  XNOR2_X1 U559 ( .A(n391), .B(n735), .ZN(G33) );
  INV_X1 U560 ( .A(n647), .ZN(n392) );
  NAND2_X1 U561 ( .A1(n570), .A2(n569), .ZN(n393) );
  XNOR2_X2 U562 ( .A(n397), .B(n396), .ZN(n639) );
  AND2_X1 U563 ( .A1(n682), .A2(n620), .ZN(n398) );
  NAND2_X1 U564 ( .A1(n403), .A2(n400), .ZN(n399) );
  XNOR2_X1 U565 ( .A(n518), .B(n408), .ZN(n702) );
  XNOR2_X1 U566 ( .A(n519), .B(n517), .ZN(n408) );
  XNOR2_X2 U567 ( .A(n409), .B(n345), .ZN(n734) );
  NAND2_X1 U568 ( .A1(n411), .A2(n410), .ZN(n409) );
  XNOR2_X1 U569 ( .A(n579), .B(n412), .ZN(n411) );
  INV_X1 U570 ( .A(KEYINPUT34), .ZN(n412) );
  NAND2_X1 U571 ( .A1(n414), .A2(n587), .ZN(n413) );
  INV_X1 U572 ( .A(KEYINPUT106), .ZN(n415) );
  NAND2_X1 U573 ( .A1(n424), .A2(n422), .ZN(n421) );
  NAND2_X1 U574 ( .A1(n423), .A2(n562), .ZN(n422) );
  INV_X1 U575 ( .A(n552), .ZN(n425) );
  INV_X1 U576 ( .A(KEYINPUT28), .ZN(n427) );
  INV_X1 U577 ( .A(n685), .ZN(n428) );
  NAND2_X1 U578 ( .A1(n671), .A2(n668), .ZN(n430) );
  XNOR2_X2 U579 ( .A(n534), .B(KEYINPUT111), .ZN(n671) );
  NOR2_X1 U580 ( .A1(n682), .A2(n618), .ZN(n436) );
  OR2_X1 U581 ( .A1(n682), .A2(n431), .ZN(n692) );
  OR2_X1 U582 ( .A1(n682), .A2(n432), .ZN(n700) );
  NAND2_X1 U583 ( .A1(n436), .A2(G469), .ZN(n693) );
  NAND2_X1 U584 ( .A1(n436), .A2(G478), .ZN(n701) );
  XNOR2_X1 U585 ( .A(n619), .B(KEYINPUT62), .ZN(n620) );
  AND2_X1 U586 ( .A1(G224), .A2(n727), .ZN(n445) );
  INV_X1 U587 ( .A(n648), .ZN(n569) );
  XNOR2_X1 U588 ( .A(n488), .B(n487), .ZN(n489) );
  XNOR2_X1 U589 ( .A(n449), .B(n448), .ZN(n450) );
  XNOR2_X1 U590 ( .A(n509), .B(G475), .ZN(n510) );
  XOR2_X1 U591 ( .A(n470), .B(G110), .Z(n449) );
  NOR2_X1 U592 ( .A1(n695), .A2(G902), .ZN(n457) );
  XOR2_X1 U593 ( .A(KEYINPUT67), .B(KEYINPUT69), .Z(n455) );
  XNOR2_X1 U594 ( .A(KEYINPUT68), .B(G469), .ZN(n454) );
  XOR2_X1 U595 ( .A(n455), .B(n454), .Z(n456) );
  XOR2_X1 U596 ( .A(KEYINPUT110), .B(KEYINPUT109), .Z(n494) );
  NAND2_X1 U597 ( .A1(n618), .A2(G234), .ZN(n459) );
  XNOR2_X1 U598 ( .A(KEYINPUT88), .B(KEYINPUT20), .ZN(n458) );
  XOR2_X1 U599 ( .A(KEYINPUT91), .B(n460), .Z(n461) );
  NOR2_X1 U600 ( .A1(G900), .A2(n727), .ZN(n462) );
  NAND2_X1 U601 ( .A1(n462), .A2(G902), .ZN(n463) );
  NAND2_X1 U602 ( .A1(G952), .A2(n727), .ZN(n574) );
  NAND2_X1 U603 ( .A1(n463), .A2(n574), .ZN(n466) );
  XOR2_X1 U604 ( .A(KEYINPUT14), .B(KEYINPUT85), .Z(n465) );
  XNOR2_X1 U605 ( .A(n465), .B(n464), .ZN(n578) );
  NAND2_X1 U606 ( .A1(n466), .A2(n578), .ZN(n537) );
  NOR2_X1 U607 ( .A1(n655), .A2(n537), .ZN(n484) );
  NAND2_X1 U608 ( .A1(G234), .A2(n727), .ZN(n467) );
  XOR2_X1 U609 ( .A(KEYINPUT8), .B(n467), .Z(n516) );
  NAND2_X1 U610 ( .A1(n516), .A2(G221), .ZN(n476) );
  XOR2_X1 U611 ( .A(KEYINPUT86), .B(G128), .Z(n472) );
  XNOR2_X1 U612 ( .A(n473), .B(KEYINPUT24), .ZN(n474) );
  XNOR2_X1 U613 ( .A(n474), .B(n719), .ZN(n475) );
  NOR2_X1 U614 ( .A1(n705), .A2(G902), .ZN(n483) );
  NAND2_X1 U615 ( .A1(G217), .A2(n477), .ZN(n481) );
  XOR2_X1 U616 ( .A(KEYINPUT87), .B(KEYINPUT89), .Z(n479) );
  XNOR2_X1 U617 ( .A(KEYINPUT25), .B(KEYINPUT90), .ZN(n478) );
  XNOR2_X1 U618 ( .A(n479), .B(n478), .ZN(n480) );
  NAND2_X1 U619 ( .A1(n484), .A2(n590), .ZN(n554) );
  XOR2_X1 U620 ( .A(n486), .B(n485), .Z(n488) );
  NAND2_X1 U621 ( .A1(n497), .A2(G210), .ZN(n487) );
  XNOR2_X2 U622 ( .A(n492), .B(G472), .ZN(n606) );
  OR2_X1 U623 ( .A1(n554), .A2(n652), .ZN(n493) );
  XNOR2_X1 U624 ( .A(n496), .B(n495), .ZN(n501) );
  NAND2_X1 U625 ( .A1(n497), .A2(G214), .ZN(n498) );
  XNOR2_X1 U626 ( .A(n499), .B(n498), .ZN(n500) );
  XOR2_X1 U627 ( .A(n501), .B(n500), .Z(n502) );
  XNOR2_X1 U628 ( .A(n503), .B(n502), .ZN(n508) );
  INV_X1 U629 ( .A(n526), .ZN(n504) );
  XNOR2_X1 U630 ( .A(n504), .B(G113), .ZN(n506) );
  XNOR2_X1 U631 ( .A(n513), .B(n512), .ZN(n514) );
  XOR2_X1 U632 ( .A(n515), .B(n514), .Z(n518) );
  NAND2_X1 U633 ( .A1(G217), .A2(n516), .ZN(n517) );
  XNOR2_X1 U634 ( .A(n520), .B(KEYINPUT4), .ZN(n521) );
  XNOR2_X1 U635 ( .A(n522), .B(n445), .ZN(n523) );
  XNOR2_X1 U636 ( .A(G110), .B(n525), .ZN(n527) );
  NAND2_X1 U637 ( .A1(n689), .A2(n618), .ZN(n531) );
  XOR2_X1 U638 ( .A(KEYINPUT83), .B(KEYINPUT73), .Z(n529) );
  NAND2_X1 U639 ( .A1(G210), .A2(n532), .ZN(n528) );
  XNOR2_X1 U640 ( .A(n529), .B(n528), .ZN(n530) );
  NAND2_X1 U641 ( .A1(n532), .A2(G214), .ZN(n533) );
  XOR2_X1 U642 ( .A(n533), .B(KEYINPUT84), .Z(n667) );
  INV_X1 U643 ( .A(n545), .ZN(n536) );
  XOR2_X1 U644 ( .A(KEYINPUT30), .B(KEYINPUT108), .Z(n538) );
  XNOR2_X1 U645 ( .A(KEYINPUT39), .B(KEYINPUT78), .ZN(n539) );
  XNOR2_X1 U646 ( .A(n540), .B(n539), .ZN(n571) );
  NAND2_X1 U647 ( .A1(n541), .A2(n545), .ZN(n580) );
  OR2_X1 U648 ( .A1(n547), .A2(n542), .ZN(n543) );
  NAND2_X1 U649 ( .A1(n545), .A2(n544), .ZN(n641) );
  INV_X1 U650 ( .A(n641), .ZN(n632) );
  NOR2_X1 U651 ( .A1(KEYINPUT74), .A2(n670), .ZN(n549) );
  AND2_X1 U652 ( .A1(n576), .A2(n548), .ZN(n637) );
  NAND2_X1 U653 ( .A1(n549), .A2(n637), .ZN(n550) );
  INV_X1 U654 ( .A(n572), .ZN(n601) );
  XNOR2_X1 U655 ( .A(n555), .B(KEYINPUT107), .ZN(n556) );
  NAND2_X1 U656 ( .A1(n564), .A2(n557), .ZN(n558) );
  AND2_X1 U657 ( .A1(n637), .A2(n670), .ZN(n561) );
  NAND2_X1 U658 ( .A1(n561), .A2(KEYINPUT74), .ZN(n560) );
  INV_X1 U659 ( .A(KEYINPUT47), .ZN(n559) );
  NAND2_X1 U660 ( .A1(n561), .A2(KEYINPUT47), .ZN(n562) );
  XNOR2_X1 U661 ( .A(n563), .B(KEYINPUT48), .ZN(n570) );
  NAND2_X1 U662 ( .A1(n564), .A2(n649), .ZN(n565) );
  NOR2_X1 U663 ( .A1(n667), .A2(n565), .ZN(n566) );
  XNOR2_X1 U664 ( .A(n566), .B(KEYINPUT43), .ZN(n567) );
  NOR2_X1 U665 ( .A1(n568), .A2(n567), .ZN(n648) );
  NOR2_X1 U666 ( .A1(n571), .A2(n641), .ZN(n647) );
  NOR2_X1 U667 ( .A1(G898), .A2(n727), .ZN(n716) );
  NAND2_X1 U668 ( .A1(G902), .A2(n716), .ZN(n575) );
  NAND2_X1 U669 ( .A1(n575), .A2(n574), .ZN(n577) );
  INV_X1 U670 ( .A(n578), .ZN(n679) );
  NAND2_X1 U671 ( .A1(n665), .A2(n584), .ZN(n579) );
  XNOR2_X1 U672 ( .A(n353), .B(KEYINPUT103), .ZN(n598) );
  INV_X1 U673 ( .A(n598), .ZN(n654) );
  NAND2_X1 U674 ( .A1(n601), .A2(n654), .ZN(n581) );
  XNOR2_X1 U675 ( .A(KEYINPUT105), .B(n581), .ZN(n588) );
  INV_X1 U676 ( .A(n668), .ZN(n582) );
  NOR2_X1 U677 ( .A1(n655), .A2(n582), .ZN(n583) );
  XNOR2_X1 U678 ( .A(KEYINPUT102), .B(n583), .ZN(n585) );
  NAND2_X1 U679 ( .A1(n585), .A2(n584), .ZN(n586) );
  XNOR2_X1 U680 ( .A(n586), .B(KEYINPUT22), .ZN(n592) );
  XOR2_X1 U681 ( .A(KEYINPUT65), .B(KEYINPUT32), .Z(n589) );
  NAND2_X1 U682 ( .A1(n353), .A2(n649), .ZN(n591) );
  NOR2_X1 U683 ( .A1(n592), .A2(n591), .ZN(n593) );
  NAND2_X1 U684 ( .A1(n593), .A2(n652), .ZN(n631) );
  NAND2_X1 U685 ( .A1(n732), .A2(n631), .ZN(n595) );
  XNOR2_X1 U686 ( .A(n595), .B(n594), .ZN(n596) );
  NAND2_X1 U687 ( .A1(n599), .A2(n598), .ZN(n600) );
  NOR2_X1 U688 ( .A1(n601), .A2(n600), .ZN(n622) );
  XOR2_X1 U689 ( .A(KEYINPUT92), .B(KEYINPUT31), .Z(n604) );
  NOR2_X1 U690 ( .A1(n602), .A2(n652), .ZN(n661) );
  NAND2_X1 U691 ( .A1(n661), .A2(n584), .ZN(n603) );
  XNOR2_X1 U692 ( .A(n604), .B(n603), .ZN(n642) );
  NOR2_X1 U693 ( .A1(n606), .A2(n605), .ZN(n607) );
  NAND2_X1 U694 ( .A1(n607), .A2(n584), .ZN(n626) );
  NAND2_X1 U695 ( .A1(n642), .A2(n626), .ZN(n608) );
  NAND2_X1 U696 ( .A1(n609), .A2(n608), .ZN(n610) );
  XNOR2_X1 U697 ( .A(KEYINPUT101), .B(n610), .ZN(n611) );
  NOR2_X1 U698 ( .A1(n622), .A2(n611), .ZN(n612) );
  XNOR2_X1 U699 ( .A(n612), .B(KEYINPUT104), .ZN(n613) );
  XNOR2_X1 U700 ( .A(KEYINPUT45), .B(KEYINPUT64), .ZN(n615) );
  INV_X1 U701 ( .A(n708), .ZN(n617) );
  XOR2_X1 U702 ( .A(KEYINPUT63), .B(n621), .Z(G57) );
  XOR2_X1 U703 ( .A(G101), .B(n622), .Z(G3) );
  NOR2_X1 U704 ( .A1(n639), .A2(n626), .ZN(n623) );
  XOR2_X1 U705 ( .A(G104), .B(n623), .Z(G6) );
  XOR2_X1 U706 ( .A(KEYINPUT114), .B(KEYINPUT113), .Z(n625) );
  XNOR2_X1 U707 ( .A(KEYINPUT112), .B(KEYINPUT27), .ZN(n624) );
  XNOR2_X1 U708 ( .A(n625), .B(n624), .ZN(n630) );
  NOR2_X1 U709 ( .A1(n641), .A2(n626), .ZN(n628) );
  XNOR2_X1 U710 ( .A(G107), .B(KEYINPUT26), .ZN(n627) );
  XNOR2_X1 U711 ( .A(n628), .B(n627), .ZN(n629) );
  XNOR2_X1 U712 ( .A(n630), .B(n629), .ZN(G9) );
  XNOR2_X1 U713 ( .A(G110), .B(n631), .ZN(G12) );
  XOR2_X1 U714 ( .A(G128), .B(KEYINPUT29), .Z(n634) );
  NAND2_X1 U715 ( .A1(n637), .A2(n632), .ZN(n633) );
  XNOR2_X1 U716 ( .A(n634), .B(n633), .ZN(G30) );
  XOR2_X1 U717 ( .A(G143), .B(n635), .Z(G45) );
  NAND2_X1 U718 ( .A1(n637), .A2(n636), .ZN(n638) );
  XNOR2_X1 U719 ( .A(n638), .B(G146), .ZN(G48) );
  NOR2_X1 U720 ( .A1(n642), .A2(n639), .ZN(n640) );
  XOR2_X1 U721 ( .A(G113), .B(n640), .Z(G15) );
  NOR2_X1 U722 ( .A1(n642), .A2(n641), .ZN(n643) );
  XOR2_X1 U723 ( .A(G116), .B(n643), .Z(G18) );
  XOR2_X1 U724 ( .A(KEYINPUT115), .B(KEYINPUT37), .Z(n646) );
  XNOR2_X1 U725 ( .A(n644), .B(G125), .ZN(n645) );
  XNOR2_X1 U726 ( .A(n646), .B(n645), .ZN(G27) );
  XOR2_X1 U727 ( .A(G134), .B(n647), .Z(G36) );
  XOR2_X1 U728 ( .A(G140), .B(n648), .Z(G42) );
  NAND2_X1 U729 ( .A1(n650), .A2(n649), .ZN(n651) );
  XNOR2_X1 U730 ( .A(n651), .B(KEYINPUT50), .ZN(n653) );
  NAND2_X1 U731 ( .A1(n653), .A2(n652), .ZN(n658) );
  NAND2_X1 U732 ( .A1(n655), .A2(n654), .ZN(n656) );
  XNOR2_X1 U733 ( .A(KEYINPUT49), .B(n656), .ZN(n657) );
  NOR2_X1 U734 ( .A1(n658), .A2(n657), .ZN(n659) );
  XNOR2_X1 U735 ( .A(n659), .B(KEYINPUT116), .ZN(n660) );
  NOR2_X1 U736 ( .A1(n661), .A2(n660), .ZN(n662) );
  NOR2_X1 U737 ( .A1(n364), .A2(n663), .ZN(n664) );
  NAND2_X1 U738 ( .A1(n667), .A2(n666), .ZN(n669) );
  NAND2_X1 U739 ( .A1(n669), .A2(n668), .ZN(n673) );
  NAND2_X1 U740 ( .A1(n671), .A2(n670), .ZN(n672) );
  NAND2_X1 U741 ( .A1(n673), .A2(n672), .ZN(n674) );
  NAND2_X1 U742 ( .A1(n683), .A2(n674), .ZN(n675) );
  XNOR2_X1 U743 ( .A(KEYINPUT52), .B(n676), .ZN(n677) );
  NAND2_X1 U744 ( .A1(n677), .A2(G952), .ZN(n678) );
  NOR2_X1 U745 ( .A1(n679), .A2(n678), .ZN(n680) );
  XNOR2_X1 U746 ( .A(n680), .B(KEYINPUT119), .ZN(n681) );
  NAND2_X1 U747 ( .A1(n682), .A2(n681), .ZN(n687) );
  INV_X1 U748 ( .A(n683), .ZN(n684) );
  NOR2_X1 U749 ( .A1(n364), .A2(n684), .ZN(n686) );
  NOR2_X1 U750 ( .A1(n687), .A2(n686), .ZN(n688) );
  XOR2_X1 U751 ( .A(KEYINPUT120), .B(KEYINPUT54), .Z(n691) );
  XNOR2_X1 U752 ( .A(n689), .B(KEYINPUT55), .ZN(n690) );
  XOR2_X1 U753 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n694) );
  NOR2_X1 U754 ( .A1(n707), .A2(n696), .ZN(G54) );
  XOR2_X1 U755 ( .A(KEYINPUT59), .B(KEYINPUT121), .Z(n699) );
  XNOR2_X1 U756 ( .A(n697), .B(KEYINPUT81), .ZN(n698) );
  XNOR2_X1 U757 ( .A(n702), .B(n701), .ZN(n703) );
  NOR2_X1 U758 ( .A1(n707), .A2(n703), .ZN(G63) );
  XNOR2_X1 U759 ( .A(n704), .B(n705), .ZN(n706) );
  BUF_X1 U760 ( .A(n708), .Z(n709) );
  NAND2_X1 U761 ( .A1(n727), .A2(n709), .ZN(n713) );
  NAND2_X1 U762 ( .A1(G953), .A2(G224), .ZN(n710) );
  XNOR2_X1 U763 ( .A(KEYINPUT61), .B(n710), .ZN(n711) );
  NAND2_X1 U764 ( .A1(n711), .A2(G898), .ZN(n712) );
  NAND2_X1 U765 ( .A1(n713), .A2(n712), .ZN(n718) );
  XNOR2_X1 U766 ( .A(KEYINPUT123), .B(n714), .ZN(n715) );
  NOR2_X1 U767 ( .A1(n716), .A2(n715), .ZN(n717) );
  XNOR2_X1 U768 ( .A(n718), .B(n717), .ZN(G69) );
  XOR2_X1 U769 ( .A(n719), .B(KEYINPUT124), .Z(n720) );
  XNOR2_X1 U770 ( .A(n721), .B(n720), .ZN(n725) );
  INV_X1 U771 ( .A(n722), .ZN(n723) );
  XNOR2_X1 U772 ( .A(n725), .B(n723), .ZN(n724) );
  NAND2_X1 U773 ( .A1(n724), .A2(n727), .ZN(n730) );
  XOR2_X1 U774 ( .A(G227), .B(n725), .Z(n726) );
  NOR2_X1 U775 ( .A1(n727), .A2(n726), .ZN(n728) );
  NAND2_X1 U776 ( .A1(G900), .A2(n728), .ZN(n729) );
  NAND2_X1 U777 ( .A1(n730), .A2(n729), .ZN(n731) );
  XNOR2_X1 U778 ( .A(KEYINPUT125), .B(n731), .ZN(G72) );
  XNOR2_X1 U779 ( .A(n732), .B(G119), .ZN(n733) );
  XNOR2_X1 U780 ( .A(n733), .B(KEYINPUT126), .ZN(G21) );
  XNOR2_X1 U781 ( .A(n734), .B(G122), .ZN(G24) );
  XNOR2_X1 U782 ( .A(G131), .B(KEYINPUT127), .ZN(n735) );
  XOR2_X1 U783 ( .A(n736), .B(G137), .Z(G39) );
endmodule

