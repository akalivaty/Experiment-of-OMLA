//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 0 0 0 0 0 1 1 0 0 1 1 0 1 0 0 0 1 0 1 0 1 1 0 1 1 1 1 1 0 0 0 0 1 1 0 0 0 1 1 0 0 1 1 0 1 0 0 0 1 0 0 1 1 0 0 1 0 1 0 0 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:35:25 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n206, new_n207, new_n208,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n605,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n681, new_n682, new_n683, new_n684, new_n685,
    new_n686, new_n687, new_n688, new_n689, new_n690, new_n691, new_n692,
    new_n693, new_n694, new_n695, new_n696, new_n697, new_n698, new_n699,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n753, new_n754, new_n755, new_n756,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n799,
    new_n800, new_n801, new_n802, new_n803, new_n804, new_n805, new_n806,
    new_n807, new_n808, new_n809, new_n810, new_n811, new_n812, new_n813,
    new_n814, new_n815, new_n816, new_n817, new_n818, new_n819, new_n820,
    new_n821, new_n822, new_n823, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n898,
    new_n899, new_n900, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n965, new_n966, new_n967, new_n968, new_n969,
    new_n970, new_n971, new_n972, new_n973, new_n974, new_n975, new_n976,
    new_n977, new_n978, new_n979, new_n980, new_n981, new_n982, new_n983,
    new_n984, new_n985, new_n986, new_n987, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1010,
    new_n1011, new_n1012, new_n1013, new_n1014, new_n1015, new_n1016,
    new_n1017, new_n1018, new_n1019, new_n1020, new_n1021, new_n1022,
    new_n1023, new_n1024, new_n1025, new_n1026, new_n1027, new_n1028,
    new_n1029, new_n1030, new_n1032, new_n1033, new_n1034, new_n1035,
    new_n1036, new_n1037, new_n1038, new_n1039, new_n1040, new_n1041,
    new_n1042, new_n1043, new_n1044, new_n1045, new_n1046, new_n1047,
    new_n1048, new_n1049, new_n1050, new_n1051, new_n1052, new_n1053,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1102,
    new_n1103, new_n1104, new_n1105, new_n1106, new_n1107, new_n1108,
    new_n1109, new_n1110, new_n1111, new_n1112, new_n1113, new_n1114,
    new_n1115, new_n1116, new_n1117, new_n1118, new_n1119, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1164, new_n1165, new_n1166, new_n1167, new_n1168, new_n1169,
    new_n1170, new_n1171, new_n1172, new_n1173, new_n1174, new_n1175,
    new_n1176, new_n1177, new_n1178, new_n1179, new_n1180, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1187, new_n1188, new_n1189,
    new_n1190, new_n1192, new_n1193, new_n1194, new_n1195, new_n1196,
    new_n1197, new_n1198, new_n1199, new_n1200, new_n1201, new_n1202,
    new_n1203, new_n1204, new_n1205, new_n1206, new_n1207, new_n1208,
    new_n1209, new_n1210, new_n1211, new_n1212, new_n1213, new_n1214,
    new_n1215, new_n1216, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1263,
    new_n1264, new_n1265, new_n1266, new_n1267, new_n1268, new_n1269,
    new_n1270;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  XOR2_X1   g0003(.A(new_n203), .B(KEYINPUT64), .Z(new_n204));
  NOR2_X1   g0004(.A1(new_n204), .A2(G77), .ZN(G353));
  NOR2_X1   g0005(.A1(G97), .A2(G107), .ZN(new_n206));
  INV_X1    g0006(.A(new_n206), .ZN(new_n207));
  NAND2_X1  g0007(.A1(new_n207), .A2(G87), .ZN(new_n208));
  XOR2_X1   g0008(.A(new_n208), .B(KEYINPUT65), .Z(G355));
  INV_X1    g0009(.A(G1), .ZN(new_n210));
  INV_X1    g0010(.A(G20), .ZN(new_n211));
  NOR2_X1   g0011(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  INV_X1    g0012(.A(new_n212), .ZN(new_n213));
  NOR2_X1   g0013(.A1(new_n213), .A2(G13), .ZN(new_n214));
  OAI211_X1 g0014(.A(new_n214), .B(G250), .C1(G257), .C2(G264), .ZN(new_n215));
  XNOR2_X1  g0015(.A(new_n215), .B(KEYINPUT0), .ZN(new_n216));
  NAND2_X1  g0016(.A1(G1), .A2(G13), .ZN(new_n217));
  NOR2_X1   g0017(.A1(new_n217), .A2(new_n211), .ZN(new_n218));
  INV_X1    g0018(.A(new_n218), .ZN(new_n219));
  INV_X1    g0019(.A(new_n201), .ZN(new_n220));
  NAND2_X1  g0020(.A1(new_n220), .A2(G50), .ZN(new_n221));
  AOI22_X1  g0021(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n222));
  INV_X1    g0022(.A(G68), .ZN(new_n223));
  INV_X1    g0023(.A(G238), .ZN(new_n224));
  INV_X1    g0024(.A(G87), .ZN(new_n225));
  INV_X1    g0025(.A(G250), .ZN(new_n226));
  OAI221_X1 g0026(.A(new_n222), .B1(new_n223), .B2(new_n224), .C1(new_n225), .C2(new_n226), .ZN(new_n227));
  AOI22_X1  g0027(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n228));
  AOI22_X1  g0028(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n229));
  NAND2_X1  g0029(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  OAI21_X1  g0030(.A(new_n213), .B1(new_n227), .B2(new_n230), .ZN(new_n231));
  OAI221_X1 g0031(.A(new_n216), .B1(new_n219), .B2(new_n221), .C1(KEYINPUT1), .C2(new_n231), .ZN(new_n232));
  AOI21_X1  g0032(.A(new_n232), .B1(KEYINPUT1), .B2(new_n231), .ZN(G361));
  XOR2_X1   g0033(.A(G238), .B(G244), .Z(new_n234));
  XNOR2_X1  g0034(.A(new_n234), .B(G232), .ZN(new_n235));
  XOR2_X1   g0035(.A(KEYINPUT2), .B(G226), .Z(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XNOR2_X1  g0037(.A(G250), .B(G257), .ZN(new_n238));
  XNOR2_X1  g0038(.A(G264), .B(G270), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XOR2_X1   g0040(.A(new_n237), .B(new_n240), .Z(G358));
  XOR2_X1   g0041(.A(G87), .B(G97), .Z(new_n242));
  XNOR2_X1  g0042(.A(G107), .B(G116), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  NAND2_X1  g0044(.A1(new_n202), .A2(G68), .ZN(new_n245));
  NAND2_X1  g0045(.A1(new_n223), .A2(G50), .ZN(new_n246));
  NAND2_X1  g0046(.A1(new_n245), .A2(new_n246), .ZN(new_n247));
  XNOR2_X1  g0047(.A(G58), .B(G77), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n247), .B(new_n248), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n244), .B(new_n249), .ZN(G351));
  INV_X1    g0050(.A(KEYINPUT73), .ZN(new_n251));
  AOI21_X1  g0051(.A(new_n217), .B1(G33), .B2(G41), .ZN(new_n252));
  INV_X1    g0052(.A(G274), .ZN(new_n253));
  OAI21_X1  g0053(.A(new_n210), .B1(G41), .B2(G45), .ZN(new_n254));
  NOR3_X1   g0054(.A1(new_n252), .A2(new_n253), .A3(new_n254), .ZN(new_n255));
  INV_X1    g0055(.A(new_n255), .ZN(new_n256));
  INV_X1    g0056(.A(new_n254), .ZN(new_n257));
  NOR2_X1   g0057(.A1(new_n252), .A2(new_n257), .ZN(new_n258));
  INV_X1    g0058(.A(new_n258), .ZN(new_n259));
  INV_X1    g0059(.A(G226), .ZN(new_n260));
  OAI21_X1  g0060(.A(new_n256), .B1(new_n259), .B2(new_n260), .ZN(new_n261));
  AND2_X1   g0061(.A1(KEYINPUT3), .A2(G33), .ZN(new_n262));
  NOR2_X1   g0062(.A1(KEYINPUT3), .A2(G33), .ZN(new_n263));
  NOR2_X1   g0063(.A1(new_n262), .A2(new_n263), .ZN(new_n264));
  INV_X1    g0064(.A(G1698), .ZN(new_n265));
  NOR2_X1   g0065(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  AOI22_X1  g0066(.A1(new_n266), .A2(G223), .B1(G77), .B2(new_n264), .ZN(new_n267));
  INV_X1    g0067(.A(G222), .ZN(new_n268));
  INV_X1    g0068(.A(KEYINPUT3), .ZN(new_n269));
  INV_X1    g0069(.A(G33), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  NAND2_X1  g0071(.A1(KEYINPUT3), .A2(G33), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n273), .A2(new_n265), .ZN(new_n274));
  OAI21_X1  g0074(.A(new_n267), .B1(new_n268), .B2(new_n274), .ZN(new_n275));
  AOI21_X1  g0075(.A(new_n261), .B1(new_n275), .B2(new_n252), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n276), .A2(G190), .ZN(new_n277));
  INV_X1    g0077(.A(G200), .ZN(new_n278));
  OAI21_X1  g0078(.A(new_n277), .B1(new_n278), .B2(new_n276), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n212), .A2(G33), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n280), .A2(new_n217), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n204), .A2(G20), .ZN(new_n282));
  INV_X1    g0082(.A(G58), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n283), .A2(KEYINPUT8), .ZN(new_n284));
  INV_X1    g0084(.A(KEYINPUT8), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n285), .A2(G58), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n284), .A2(new_n286), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n287), .A2(KEYINPUT66), .ZN(new_n288));
  XNOR2_X1  g0088(.A(KEYINPUT8), .B(G58), .ZN(new_n289));
  INV_X1    g0089(.A(KEYINPUT66), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  NOR2_X1   g0091(.A1(new_n270), .A2(G20), .ZN(new_n292));
  NAND3_X1  g0092(.A1(new_n288), .A2(new_n291), .A3(new_n292), .ZN(new_n293));
  NOR2_X1   g0093(.A1(G20), .A2(G33), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n294), .A2(G150), .ZN(new_n295));
  NAND3_X1  g0095(.A1(new_n293), .A2(KEYINPUT67), .A3(new_n295), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n282), .A2(new_n296), .ZN(new_n297));
  AOI21_X1  g0097(.A(KEYINPUT67), .B1(new_n293), .B2(new_n295), .ZN(new_n298));
  OAI21_X1  g0098(.A(new_n281), .B1(new_n297), .B2(new_n298), .ZN(new_n299));
  INV_X1    g0099(.A(G13), .ZN(new_n300));
  NOR2_X1   g0100(.A1(new_n300), .A2(G1), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n301), .A2(G20), .ZN(new_n302));
  NOR2_X1   g0102(.A1(new_n302), .A2(G50), .ZN(new_n303));
  NOR2_X1   g0103(.A1(new_n211), .A2(G1), .ZN(new_n304));
  NOR2_X1   g0104(.A1(new_n281), .A2(new_n304), .ZN(new_n305));
  AOI21_X1  g0105(.A(new_n303), .B1(new_n305), .B2(G50), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n299), .A2(new_n306), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n307), .A2(KEYINPUT9), .ZN(new_n308));
  INV_X1    g0108(.A(KEYINPUT9), .ZN(new_n309));
  NAND3_X1  g0109(.A1(new_n299), .A2(new_n309), .A3(new_n306), .ZN(new_n310));
  AOI21_X1  g0110(.A(new_n279), .B1(new_n308), .B2(new_n310), .ZN(new_n311));
  INV_X1    g0111(.A(KEYINPUT10), .ZN(new_n312));
  OAI21_X1  g0112(.A(new_n251), .B1(new_n311), .B2(new_n312), .ZN(new_n313));
  INV_X1    g0113(.A(new_n310), .ZN(new_n314));
  AOI21_X1  g0114(.A(new_n309), .B1(new_n299), .B2(new_n306), .ZN(new_n315));
  NOR2_X1   g0115(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  OAI211_X1 g0116(.A(KEYINPUT73), .B(KEYINPUT10), .C1(new_n316), .C2(new_n279), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n313), .A2(new_n317), .ZN(new_n318));
  OAI21_X1  g0118(.A(KEYINPUT72), .B1(new_n314), .B2(new_n315), .ZN(new_n319));
  INV_X1    g0119(.A(KEYINPUT72), .ZN(new_n320));
  NAND3_X1  g0120(.A1(new_n308), .A2(new_n320), .A3(new_n310), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n319), .A2(new_n321), .ZN(new_n322));
  NOR2_X1   g0122(.A1(new_n279), .A2(KEYINPUT10), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n318), .A2(new_n324), .ZN(new_n325));
  NAND3_X1  g0125(.A1(new_n273), .A2(G232), .A3(new_n265), .ZN(new_n326));
  INV_X1    g0126(.A(G107), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n273), .A2(G1698), .ZN(new_n328));
  OAI221_X1 g0128(.A(new_n326), .B1(new_n327), .B2(new_n273), .C1(new_n328), .C2(new_n224), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n329), .A2(new_n252), .ZN(new_n330));
  AOI21_X1  g0130(.A(new_n255), .B1(G244), .B2(new_n258), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n330), .A2(new_n331), .ZN(new_n332));
  INV_X1    g0132(.A(new_n332), .ZN(new_n333));
  INV_X1    g0133(.A(G179), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n333), .A2(new_n334), .ZN(new_n335));
  AOI22_X1  g0135(.A1(new_n287), .A2(new_n294), .B1(G20), .B2(G77), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n336), .A2(KEYINPUT68), .ZN(new_n337));
  INV_X1    g0137(.A(new_n292), .ZN(new_n338));
  XNOR2_X1  g0138(.A(KEYINPUT15), .B(G87), .ZN(new_n339));
  OAI21_X1  g0139(.A(new_n337), .B1(new_n338), .B2(new_n339), .ZN(new_n340));
  NOR2_X1   g0140(.A1(new_n336), .A2(KEYINPUT68), .ZN(new_n341));
  OAI21_X1  g0141(.A(new_n281), .B1(new_n340), .B2(new_n341), .ZN(new_n342));
  INV_X1    g0142(.A(KEYINPUT69), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n302), .A2(new_n343), .ZN(new_n344));
  NOR3_X1   g0144(.A1(new_n300), .A2(new_n211), .A3(G1), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n345), .A2(KEYINPUT69), .ZN(new_n346));
  AOI21_X1  g0146(.A(new_n281), .B1(new_n344), .B2(new_n346), .ZN(new_n347));
  INV_X1    g0147(.A(G77), .ZN(new_n348));
  AND2_X1   g0148(.A1(new_n344), .A2(new_n346), .ZN(new_n349));
  NOR2_X1   g0149(.A1(new_n304), .A2(new_n348), .ZN(new_n350));
  OAI22_X1  g0150(.A1(new_n347), .A2(new_n348), .B1(new_n349), .B2(new_n350), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n342), .A2(new_n351), .ZN(new_n352));
  INV_X1    g0152(.A(G169), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n332), .A2(new_n353), .ZN(new_n354));
  NAND3_X1  g0154(.A1(new_n335), .A2(new_n352), .A3(new_n354), .ZN(new_n355));
  OAI211_X1 g0155(.A(new_n342), .B(new_n351), .C1(new_n333), .C2(new_n278), .ZN(new_n356));
  INV_X1    g0156(.A(KEYINPUT70), .ZN(new_n357));
  INV_X1    g0157(.A(G190), .ZN(new_n358));
  OAI22_X1  g0158(.A1(new_n356), .A2(new_n357), .B1(new_n358), .B2(new_n332), .ZN(new_n359));
  AND2_X1   g0159(.A1(new_n356), .A2(new_n357), .ZN(new_n360));
  OAI21_X1  g0160(.A(new_n355), .B1(new_n359), .B2(new_n360), .ZN(new_n361));
  INV_X1    g0161(.A(KEYINPUT71), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n361), .A2(new_n362), .ZN(new_n363));
  OAI211_X1 g0163(.A(KEYINPUT71), .B(new_n355), .C1(new_n359), .C2(new_n360), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n363), .A2(new_n364), .ZN(new_n365));
  NOR2_X1   g0165(.A1(new_n276), .A2(G169), .ZN(new_n366));
  AOI21_X1  g0166(.A(new_n366), .B1(new_n334), .B2(new_n276), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n367), .A2(new_n307), .ZN(new_n368));
  NAND3_X1  g0168(.A1(new_n325), .A2(new_n365), .A3(new_n368), .ZN(new_n369));
  INV_X1    g0169(.A(KEYINPUT74), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n369), .A2(new_n370), .ZN(new_n371));
  NAND4_X1  g0171(.A1(new_n325), .A2(new_n365), .A3(KEYINPUT74), .A4(new_n368), .ZN(new_n372));
  AND2_X1   g0172(.A1(KEYINPUT78), .A2(G169), .ZN(new_n373));
  NAND3_X1  g0173(.A1(new_n273), .A2(G232), .A3(G1698), .ZN(new_n374));
  NAND3_X1  g0174(.A1(new_n273), .A2(G226), .A3(new_n265), .ZN(new_n375));
  NAND2_X1  g0175(.A1(G33), .A2(G97), .ZN(new_n376));
  NAND3_X1  g0176(.A1(new_n374), .A2(new_n375), .A3(new_n376), .ZN(new_n377));
  INV_X1    g0177(.A(KEYINPUT75), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n377), .A2(new_n378), .ZN(new_n379));
  NAND4_X1  g0179(.A1(new_n374), .A2(new_n375), .A3(KEYINPUT75), .A4(new_n376), .ZN(new_n380));
  NAND3_X1  g0180(.A1(new_n379), .A2(new_n252), .A3(new_n380), .ZN(new_n381));
  INV_X1    g0181(.A(KEYINPUT13), .ZN(new_n382));
  AOI21_X1  g0182(.A(new_n255), .B1(G238), .B2(new_n258), .ZN(new_n383));
  AND3_X1   g0183(.A1(new_n381), .A2(new_n382), .A3(new_n383), .ZN(new_n384));
  AOI21_X1  g0184(.A(new_n382), .B1(new_n381), .B2(new_n383), .ZN(new_n385));
  OAI21_X1  g0185(.A(new_n373), .B1(new_n384), .B2(new_n385), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n386), .A2(KEYINPUT14), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n381), .A2(new_n383), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n388), .A2(KEYINPUT13), .ZN(new_n389));
  NAND3_X1  g0189(.A1(new_n381), .A2(new_n382), .A3(new_n383), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n389), .A2(new_n390), .ZN(new_n391));
  INV_X1    g0191(.A(KEYINPUT14), .ZN(new_n392));
  NAND3_X1  g0192(.A1(new_n391), .A2(new_n392), .A3(new_n373), .ZN(new_n393));
  INV_X1    g0193(.A(KEYINPUT76), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n390), .A2(new_n394), .ZN(new_n395));
  NAND4_X1  g0195(.A1(new_n381), .A2(KEYINPUT76), .A3(new_n382), .A4(new_n383), .ZN(new_n396));
  NAND4_X1  g0196(.A1(new_n395), .A2(new_n389), .A3(G179), .A4(new_n396), .ZN(new_n397));
  NAND3_X1  g0197(.A1(new_n387), .A2(new_n393), .A3(new_n397), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n294), .A2(G50), .ZN(new_n399));
  OAI221_X1 g0199(.A(new_n399), .B1(new_n211), .B2(G68), .C1(new_n348), .C2(new_n338), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n400), .A2(new_n281), .ZN(new_n401));
  INV_X1    g0201(.A(KEYINPUT11), .ZN(new_n402));
  XNOR2_X1  g0202(.A(new_n401), .B(new_n402), .ZN(new_n403));
  NOR2_X1   g0203(.A1(new_n304), .A2(new_n223), .ZN(new_n404));
  AOI21_X1  g0204(.A(new_n403), .B1(new_n347), .B2(new_n404), .ZN(new_n405));
  INV_X1    g0205(.A(KEYINPUT12), .ZN(new_n406));
  AOI21_X1  g0206(.A(new_n406), .B1(new_n349), .B2(new_n223), .ZN(new_n407));
  XNOR2_X1  g0207(.A(new_n407), .B(KEYINPUT77), .ZN(new_n408));
  NAND4_X1  g0208(.A1(new_n301), .A2(new_n406), .A3(G20), .A4(new_n223), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n408), .A2(new_n409), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n405), .A2(new_n410), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n398), .A2(new_n411), .ZN(new_n412));
  AND2_X1   g0212(.A1(new_n405), .A2(new_n410), .ZN(new_n413));
  NAND4_X1  g0213(.A1(new_n395), .A2(new_n389), .A3(G190), .A4(new_n396), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n391), .A2(G200), .ZN(new_n415));
  NAND3_X1  g0215(.A1(new_n413), .A2(new_n414), .A3(new_n415), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n412), .A2(new_n416), .ZN(new_n417));
  NAND3_X1  g0217(.A1(new_n273), .A2(G223), .A3(new_n265), .ZN(new_n418));
  NAND2_X1  g0218(.A1(G33), .A2(G87), .ZN(new_n419));
  OAI211_X1 g0219(.A(new_n418), .B(new_n419), .C1(new_n328), .C2(new_n260), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n420), .A2(new_n252), .ZN(new_n421));
  AOI21_X1  g0221(.A(new_n255), .B1(G232), .B2(new_n258), .ZN(new_n422));
  AND3_X1   g0222(.A1(new_n421), .A2(G179), .A3(new_n422), .ZN(new_n423));
  AOI21_X1  g0223(.A(new_n353), .B1(new_n421), .B2(new_n422), .ZN(new_n424));
  NOR2_X1   g0224(.A1(new_n423), .A2(new_n424), .ZN(new_n425));
  NOR2_X1   g0225(.A1(new_n283), .A2(new_n223), .ZN(new_n426));
  OR2_X1    g0226(.A1(new_n426), .A2(new_n201), .ZN(new_n427));
  AOI22_X1  g0227(.A1(new_n427), .A2(G20), .B1(G159), .B2(new_n294), .ZN(new_n428));
  NAND3_X1  g0228(.A1(new_n271), .A2(new_n211), .A3(new_n272), .ZN(new_n429));
  INV_X1    g0229(.A(KEYINPUT7), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n429), .A2(new_n430), .ZN(new_n431));
  NAND4_X1  g0231(.A1(new_n271), .A2(KEYINPUT7), .A3(new_n211), .A4(new_n272), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n431), .A2(new_n432), .ZN(new_n433));
  AOI21_X1  g0233(.A(KEYINPUT79), .B1(new_n433), .B2(G68), .ZN(new_n434));
  INV_X1    g0234(.A(KEYINPUT79), .ZN(new_n435));
  AOI211_X1 g0235(.A(new_n435), .B(new_n223), .C1(new_n431), .C2(new_n432), .ZN(new_n436));
  OAI211_X1 g0236(.A(KEYINPUT16), .B(new_n428), .C1(new_n434), .C2(new_n436), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n433), .A2(G68), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n438), .A2(new_n428), .ZN(new_n439));
  INV_X1    g0239(.A(KEYINPUT16), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n439), .A2(new_n440), .ZN(new_n441));
  NAND3_X1  g0241(.A1(new_n437), .A2(new_n281), .A3(new_n441), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n288), .A2(new_n291), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n443), .A2(new_n302), .ZN(new_n444));
  OAI21_X1  g0244(.A(new_n444), .B1(new_n443), .B2(new_n305), .ZN(new_n445));
  AOI21_X1  g0245(.A(new_n425), .B1(new_n442), .B2(new_n445), .ZN(new_n446));
  XNOR2_X1  g0246(.A(new_n446), .B(KEYINPUT18), .ZN(new_n447));
  NAND3_X1  g0247(.A1(new_n421), .A2(new_n358), .A3(new_n422), .ZN(new_n448));
  AND2_X1   g0248(.A1(new_n421), .A2(new_n422), .ZN(new_n449));
  OAI21_X1  g0249(.A(new_n448), .B1(new_n449), .B2(G200), .ZN(new_n450));
  NAND3_X1  g0250(.A1(new_n450), .A2(new_n442), .A3(new_n445), .ZN(new_n451));
  XNOR2_X1  g0251(.A(new_n451), .B(KEYINPUT17), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n447), .A2(new_n452), .ZN(new_n453));
  NOR2_X1   g0253(.A1(new_n417), .A2(new_n453), .ZN(new_n454));
  NAND3_X1  g0254(.A1(new_n371), .A2(new_n372), .A3(new_n454), .ZN(new_n455));
  INV_X1    g0255(.A(new_n455), .ZN(new_n456));
  INV_X1    g0256(.A(KEYINPUT80), .ZN(new_n457));
  INV_X1    g0257(.A(G41), .ZN(new_n458));
  OAI21_X1  g0258(.A(new_n457), .B1(new_n458), .B2(KEYINPUT5), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n458), .A2(KEYINPUT5), .ZN(new_n460));
  AND2_X1   g0260(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  INV_X1    g0261(.A(G45), .ZN(new_n462));
  NOR2_X1   g0262(.A1(new_n462), .A2(G1), .ZN(new_n463));
  OAI21_X1  g0263(.A(new_n463), .B1(new_n460), .B2(KEYINPUT80), .ZN(new_n464));
  NOR2_X1   g0264(.A1(new_n461), .A2(new_n464), .ZN(new_n465));
  NOR2_X1   g0265(.A1(new_n252), .A2(new_n253), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  INV_X1    g0267(.A(new_n252), .ZN(new_n468));
  OAI211_X1 g0268(.A(G257), .B(new_n468), .C1(new_n461), .C2(new_n464), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n467), .A2(new_n469), .ZN(new_n470));
  INV_X1    g0270(.A(KEYINPUT4), .ZN(new_n471));
  INV_X1    g0271(.A(G244), .ZN(new_n472));
  OAI21_X1  g0272(.A(new_n471), .B1(new_n274), .B2(new_n472), .ZN(new_n473));
  NOR2_X1   g0273(.A1(new_n264), .A2(G1698), .ZN(new_n474));
  NAND3_X1  g0274(.A1(new_n474), .A2(KEYINPUT4), .A3(G244), .ZN(new_n475));
  NAND2_X1  g0275(.A1(G33), .A2(G283), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n266), .A2(G250), .ZN(new_n477));
  NAND4_X1  g0277(.A1(new_n473), .A2(new_n475), .A3(new_n476), .A4(new_n477), .ZN(new_n478));
  AOI21_X1  g0278(.A(new_n470), .B1(new_n478), .B2(new_n252), .ZN(new_n479));
  OR2_X1    g0279(.A1(new_n479), .A2(G169), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n479), .A2(new_n334), .ZN(new_n481));
  INV_X1    g0281(.A(G97), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n345), .A2(new_n482), .ZN(new_n483));
  AOI21_X1  g0283(.A(new_n345), .B1(new_n210), .B2(G33), .ZN(new_n484));
  NAND3_X1  g0284(.A1(new_n484), .A2(new_n217), .A3(new_n280), .ZN(new_n485));
  OAI21_X1  g0285(.A(new_n483), .B1(new_n485), .B2(new_n482), .ZN(new_n486));
  NAND3_X1  g0286(.A1(new_n327), .A2(KEYINPUT6), .A3(G97), .ZN(new_n487));
  NOR2_X1   g0287(.A1(new_n482), .A2(new_n327), .ZN(new_n488));
  NOR2_X1   g0288(.A1(new_n488), .A2(new_n206), .ZN(new_n489));
  OAI21_X1  g0289(.A(new_n487), .B1(new_n489), .B2(KEYINPUT6), .ZN(new_n490));
  AOI22_X1  g0290(.A1(new_n490), .A2(G20), .B1(G77), .B2(new_n294), .ZN(new_n491));
  INV_X1    g0291(.A(new_n433), .ZN(new_n492));
  OAI21_X1  g0292(.A(new_n491), .B1(new_n492), .B2(new_n327), .ZN(new_n493));
  AOI21_X1  g0293(.A(new_n486), .B1(new_n493), .B2(new_n281), .ZN(new_n494));
  INV_X1    g0294(.A(new_n494), .ZN(new_n495));
  NAND3_X1  g0295(.A1(new_n480), .A2(new_n481), .A3(new_n495), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n479), .A2(G190), .ZN(new_n497));
  OAI211_X1 g0297(.A(new_n497), .B(new_n494), .C1(new_n278), .C2(new_n479), .ZN(new_n498));
  OR3_X1    g0298(.A1(new_n302), .A2(KEYINPUT25), .A3(G107), .ZN(new_n499));
  OAI21_X1  g0299(.A(KEYINPUT25), .B1(new_n302), .B2(G107), .ZN(new_n500));
  OAI211_X1 g0300(.A(new_n499), .B(new_n500), .C1(new_n485), .C2(new_n327), .ZN(new_n501));
  INV_X1    g0301(.A(KEYINPUT84), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  AND2_X1   g0303(.A1(new_n499), .A2(new_n500), .ZN(new_n504));
  OAI211_X1 g0304(.A(new_n504), .B(KEYINPUT84), .C1(new_n327), .C2(new_n485), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n503), .A2(new_n505), .ZN(new_n506));
  INV_X1    g0306(.A(KEYINPUT23), .ZN(new_n507));
  OAI21_X1  g0307(.A(new_n507), .B1(new_n211), .B2(G107), .ZN(new_n508));
  NAND3_X1  g0308(.A1(new_n327), .A2(KEYINPUT23), .A3(G20), .ZN(new_n509));
  NAND2_X1  g0309(.A1(G33), .A2(G116), .ZN(new_n510));
  INV_X1    g0310(.A(new_n510), .ZN(new_n511));
  AOI22_X1  g0311(.A1(new_n508), .A2(new_n509), .B1(new_n511), .B2(new_n211), .ZN(new_n512));
  INV_X1    g0312(.A(new_n512), .ZN(new_n513));
  NAND3_X1  g0313(.A1(new_n273), .A2(new_n211), .A3(G87), .ZN(new_n514));
  NOR2_X1   g0314(.A1(new_n514), .A2(KEYINPUT22), .ZN(new_n515));
  INV_X1    g0315(.A(new_n515), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n514), .A2(KEYINPUT22), .ZN(new_n517));
  AOI21_X1  g0317(.A(new_n513), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  OAI21_X1  g0318(.A(new_n281), .B1(new_n518), .B2(KEYINPUT24), .ZN(new_n519));
  INV_X1    g0319(.A(KEYINPUT24), .ZN(new_n520));
  AOI211_X1 g0320(.A(new_n520), .B(new_n513), .C1(new_n516), .C2(new_n517), .ZN(new_n521));
  NAND3_X1  g0321(.A1(new_n273), .A2(G257), .A3(G1698), .ZN(new_n522));
  INV_X1    g0322(.A(G294), .ZN(new_n523));
  OAI221_X1 g0323(.A(new_n522), .B1(new_n270), .B2(new_n523), .C1(new_n274), .C2(new_n226), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n524), .A2(new_n252), .ZN(new_n525));
  INV_X1    g0325(.A(new_n465), .ZN(new_n526));
  NAND3_X1  g0326(.A1(new_n526), .A2(G264), .A3(new_n468), .ZN(new_n527));
  NAND3_X1  g0327(.A1(new_n525), .A2(new_n467), .A3(new_n527), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n528), .A2(new_n278), .ZN(new_n529));
  OAI221_X1 g0329(.A(new_n506), .B1(new_n519), .B2(new_n521), .C1(new_n529), .C2(KEYINPUT86), .ZN(new_n530));
  NOR2_X1   g0330(.A1(new_n465), .A2(new_n252), .ZN(new_n531));
  AOI22_X1  g0331(.A1(new_n252), .A2(new_n524), .B1(new_n531), .B2(G264), .ZN(new_n532));
  NAND3_X1  g0332(.A1(new_n532), .A2(new_n358), .A3(new_n467), .ZN(new_n533));
  AND3_X1   g0333(.A1(new_n529), .A2(new_n533), .A3(KEYINPUT86), .ZN(new_n534));
  OAI211_X1 g0334(.A(new_n496), .B(new_n498), .C1(new_n530), .C2(new_n534), .ZN(new_n535));
  AOI21_X1  g0335(.A(new_n511), .B1(new_n266), .B2(G244), .ZN(new_n536));
  AOI21_X1  g0336(.A(KEYINPUT81), .B1(new_n474), .B2(G238), .ZN(new_n537));
  INV_X1    g0337(.A(KEYINPUT81), .ZN(new_n538));
  NOR3_X1   g0338(.A1(new_n274), .A2(new_n538), .A3(new_n224), .ZN(new_n539));
  OAI21_X1  g0339(.A(new_n536), .B1(new_n537), .B2(new_n539), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n540), .A2(new_n252), .ZN(new_n541));
  OAI211_X1 g0341(.A(new_n468), .B(G250), .C1(G1), .C2(new_n462), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n466), .A2(new_n463), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  INV_X1    g0344(.A(new_n544), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n541), .A2(new_n545), .ZN(new_n546));
  OAI21_X1  g0346(.A(KEYINPUT83), .B1(new_n546), .B2(new_n358), .ZN(new_n547));
  INV_X1    g0347(.A(KEYINPUT19), .ZN(new_n548));
  OAI21_X1  g0348(.A(new_n548), .B1(new_n338), .B2(new_n482), .ZN(new_n549));
  NAND3_X1  g0349(.A1(new_n273), .A2(new_n211), .A3(G68), .ZN(new_n550));
  OAI21_X1  g0350(.A(new_n211), .B1(new_n376), .B2(new_n548), .ZN(new_n551));
  OAI21_X1  g0351(.A(new_n551), .B1(G87), .B2(new_n207), .ZN(new_n552));
  NAND3_X1  g0352(.A1(new_n549), .A2(new_n550), .A3(new_n552), .ZN(new_n553));
  AOI22_X1  g0353(.A1(new_n281), .A2(new_n553), .B1(new_n349), .B2(new_n339), .ZN(new_n554));
  OAI21_X1  g0354(.A(new_n554), .B1(new_n225), .B2(new_n485), .ZN(new_n555));
  AOI21_X1  g0355(.A(new_n555), .B1(new_n546), .B2(G200), .ZN(new_n556));
  AOI21_X1  g0356(.A(new_n544), .B1(new_n540), .B2(new_n252), .ZN(new_n557));
  INV_X1    g0357(.A(KEYINPUT83), .ZN(new_n558));
  NAND3_X1  g0358(.A1(new_n557), .A2(new_n558), .A3(G190), .ZN(new_n559));
  NAND3_X1  g0359(.A1(new_n547), .A2(new_n556), .A3(new_n559), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n546), .A2(new_n353), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n557), .A2(new_n334), .ZN(new_n562));
  XNOR2_X1  g0362(.A(new_n339), .B(KEYINPUT82), .ZN(new_n563));
  OAI21_X1  g0363(.A(new_n554), .B1(new_n485), .B2(new_n563), .ZN(new_n564));
  NAND3_X1  g0364(.A1(new_n561), .A2(new_n562), .A3(new_n564), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n560), .A2(new_n565), .ZN(new_n566));
  NOR2_X1   g0366(.A1(new_n535), .A2(new_n566), .ZN(new_n567));
  OAI21_X1  g0367(.A(new_n506), .B1(new_n519), .B2(new_n521), .ZN(new_n568));
  INV_X1    g0368(.A(KEYINPUT85), .ZN(new_n569));
  NAND3_X1  g0369(.A1(new_n528), .A2(new_n569), .A3(G169), .ZN(new_n570));
  OAI21_X1  g0370(.A(new_n570), .B1(new_n334), .B2(new_n528), .ZN(new_n571));
  AOI21_X1  g0371(.A(new_n569), .B1(new_n528), .B2(G169), .ZN(new_n572));
  OAI21_X1  g0372(.A(new_n568), .B1(new_n571), .B2(new_n572), .ZN(new_n573));
  INV_X1    g0373(.A(G116), .ZN(new_n574));
  AOI21_X1  g0374(.A(new_n574), .B1(new_n210), .B2(G33), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n347), .A2(new_n575), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n349), .A2(new_n574), .ZN(new_n577));
  AOI22_X1  g0377(.A1(new_n280), .A2(new_n217), .B1(G20), .B2(new_n574), .ZN(new_n578));
  OAI211_X1 g0378(.A(new_n476), .B(new_n211), .C1(G33), .C2(new_n482), .ZN(new_n579));
  NAND3_X1  g0379(.A1(new_n578), .A2(KEYINPUT20), .A3(new_n579), .ZN(new_n580));
  INV_X1    g0380(.A(new_n580), .ZN(new_n581));
  AOI21_X1  g0381(.A(KEYINPUT20), .B1(new_n578), .B2(new_n579), .ZN(new_n582));
  OAI211_X1 g0382(.A(new_n576), .B(new_n577), .C1(new_n581), .C2(new_n582), .ZN(new_n583));
  NAND3_X1  g0383(.A1(new_n273), .A2(G257), .A3(new_n265), .ZN(new_n584));
  INV_X1    g0384(.A(G303), .ZN(new_n585));
  INV_X1    g0385(.A(G264), .ZN(new_n586));
  OAI221_X1 g0386(.A(new_n584), .B1(new_n585), .B2(new_n273), .C1(new_n328), .C2(new_n586), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n587), .A2(new_n252), .ZN(new_n588));
  NAND3_X1  g0388(.A1(new_n526), .A2(G270), .A3(new_n468), .ZN(new_n589));
  NAND3_X1  g0389(.A1(new_n588), .A2(new_n467), .A3(new_n589), .ZN(new_n590));
  NAND4_X1  g0390(.A1(new_n583), .A2(new_n590), .A3(KEYINPUT21), .A4(G169), .ZN(new_n591));
  AOI22_X1  g0391(.A1(new_n531), .A2(G270), .B1(new_n466), .B2(new_n465), .ZN(new_n592));
  NAND4_X1  g0392(.A1(new_n583), .A2(new_n592), .A3(G179), .A4(new_n588), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n591), .A2(new_n593), .ZN(new_n594));
  INV_X1    g0394(.A(new_n582), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n595), .A2(new_n580), .ZN(new_n596));
  AOI22_X1  g0396(.A1(new_n347), .A2(new_n575), .B1(new_n349), .B2(new_n574), .ZN(new_n597));
  AOI21_X1  g0397(.A(new_n353), .B1(new_n596), .B2(new_n597), .ZN(new_n598));
  AOI21_X1  g0398(.A(KEYINPUT21), .B1(new_n598), .B2(new_n590), .ZN(new_n599));
  NOR2_X1   g0399(.A1(new_n594), .A2(new_n599), .ZN(new_n600));
  AOI21_X1  g0400(.A(new_n583), .B1(G200), .B2(new_n590), .ZN(new_n601));
  OAI21_X1  g0401(.A(new_n601), .B1(new_n358), .B2(new_n590), .ZN(new_n602));
  AND3_X1   g0402(.A1(new_n573), .A2(new_n600), .A3(new_n602), .ZN(new_n603));
  AND3_X1   g0403(.A1(new_n456), .A2(new_n567), .A3(new_n603), .ZN(G372));
  INV_X1    g0404(.A(new_n565), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n573), .A2(new_n600), .ZN(new_n606));
  AOI21_X1  g0406(.A(new_n605), .B1(new_n567), .B2(new_n606), .ZN(new_n607));
  INV_X1    g0407(.A(new_n566), .ZN(new_n608));
  AND3_X1   g0408(.A1(new_n480), .A2(new_n481), .A3(new_n495), .ZN(new_n609));
  NAND4_X1  g0409(.A1(new_n608), .A2(KEYINPUT87), .A3(KEYINPUT26), .A4(new_n609), .ZN(new_n610));
  INV_X1    g0410(.A(KEYINPUT87), .ZN(new_n611));
  NAND3_X1  g0411(.A1(new_n609), .A2(new_n560), .A3(new_n565), .ZN(new_n612));
  INV_X1    g0412(.A(KEYINPUT26), .ZN(new_n613));
  OAI21_X1  g0413(.A(new_n611), .B1(new_n612), .B2(new_n613), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n612), .A2(new_n613), .ZN(new_n615));
  NAND3_X1  g0415(.A1(new_n610), .A2(new_n614), .A3(new_n615), .ZN(new_n616));
  AOI21_X1  g0416(.A(new_n455), .B1(new_n607), .B2(new_n616), .ZN(new_n617));
  INV_X1    g0417(.A(new_n447), .ZN(new_n618));
  AND3_X1   g0418(.A1(new_n413), .A2(new_n414), .A3(new_n415), .ZN(new_n619));
  OAI21_X1  g0419(.A(new_n412), .B1(new_n355), .B2(new_n619), .ZN(new_n620));
  AOI21_X1  g0420(.A(new_n618), .B1(new_n620), .B2(new_n452), .ZN(new_n621));
  AOI22_X1  g0421(.A1(new_n313), .A2(new_n317), .B1(new_n322), .B2(new_n323), .ZN(new_n622));
  OAI21_X1  g0422(.A(new_n368), .B1(new_n621), .B2(new_n622), .ZN(new_n623));
  OR2_X1    g0423(.A1(new_n617), .A2(new_n623), .ZN(G369));
  NAND2_X1  g0424(.A1(new_n301), .A2(new_n211), .ZN(new_n625));
  OR2_X1    g0425(.A1(new_n625), .A2(KEYINPUT27), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n625), .A2(KEYINPUT27), .ZN(new_n627));
  NAND3_X1  g0427(.A1(new_n626), .A2(G213), .A3(new_n627), .ZN(new_n628));
  INV_X1    g0428(.A(G343), .ZN(new_n629));
  NOR2_X1   g0429(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n583), .A2(new_n630), .ZN(new_n631));
  XNOR2_X1  g0431(.A(new_n600), .B(new_n631), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n632), .A2(new_n602), .ZN(new_n633));
  INV_X1    g0433(.A(new_n633), .ZN(new_n634));
  OR2_X1    g0434(.A1(new_n573), .A2(new_n630), .ZN(new_n635));
  INV_X1    g0435(.A(new_n635), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n568), .A2(new_n630), .ZN(new_n637));
  OAI21_X1  g0437(.A(new_n637), .B1(new_n530), .B2(new_n534), .ZN(new_n638));
  AND2_X1   g0438(.A1(new_n638), .A2(new_n573), .ZN(new_n639));
  NOR2_X1   g0439(.A1(new_n636), .A2(new_n639), .ZN(new_n640));
  NAND3_X1  g0440(.A1(new_n634), .A2(G330), .A3(new_n640), .ZN(new_n641));
  NOR2_X1   g0441(.A1(new_n600), .A2(new_n630), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n640), .A2(new_n642), .ZN(new_n643));
  NAND3_X1  g0443(.A1(new_n641), .A2(new_n635), .A3(new_n643), .ZN(G399));
  INV_X1    g0444(.A(new_n214), .ZN(new_n645));
  NOR2_X1   g0445(.A1(new_n645), .A2(G41), .ZN(new_n646));
  INV_X1    g0446(.A(new_n646), .ZN(new_n647));
  NOR3_X1   g0447(.A1(new_n207), .A2(G87), .A3(G116), .ZN(new_n648));
  NAND3_X1  g0448(.A1(new_n647), .A2(G1), .A3(new_n648), .ZN(new_n649));
  OAI21_X1  g0449(.A(new_n649), .B1(new_n221), .B2(new_n647), .ZN(new_n650));
  XNOR2_X1  g0450(.A(new_n650), .B(KEYINPUT28), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n616), .A2(new_n607), .ZN(new_n652));
  INV_X1    g0452(.A(new_n630), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  XNOR2_X1  g0454(.A(KEYINPUT88), .B(KEYINPUT29), .ZN(new_n655));
  XNOR2_X1  g0455(.A(new_n612), .B(new_n613), .ZN(new_n656));
  AOI21_X1  g0456(.A(new_n630), .B1(new_n607), .B2(new_n656), .ZN(new_n657));
  AOI22_X1  g0457(.A1(new_n654), .A2(new_n655), .B1(KEYINPUT29), .B2(new_n657), .ZN(new_n658));
  INV_X1    g0458(.A(G330), .ZN(new_n659));
  NOR2_X1   g0459(.A1(new_n530), .A2(new_n534), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n496), .A2(new_n498), .ZN(new_n661));
  NOR2_X1   g0461(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  NAND4_X1  g0462(.A1(new_n603), .A2(new_n662), .A3(new_n608), .A4(new_n653), .ZN(new_n663));
  NOR2_X1   g0463(.A1(new_n479), .A2(new_n557), .ZN(new_n664));
  NAND4_X1  g0464(.A1(new_n664), .A2(new_n334), .A3(new_n528), .A4(new_n590), .ZN(new_n665));
  INV_X1    g0465(.A(KEYINPUT30), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n479), .A2(new_n557), .ZN(new_n667));
  NAND4_X1  g0467(.A1(new_n532), .A2(new_n592), .A3(G179), .A4(new_n588), .ZN(new_n668));
  OAI21_X1  g0468(.A(new_n666), .B1(new_n667), .B2(new_n668), .ZN(new_n669));
  NAND4_X1  g0469(.A1(new_n588), .A2(new_n589), .A3(G179), .A4(new_n467), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n525), .A2(new_n527), .ZN(new_n671));
  NOR2_X1   g0471(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  NAND4_X1  g0472(.A1(new_n672), .A2(KEYINPUT30), .A3(new_n557), .A4(new_n479), .ZN(new_n673));
  NAND3_X1  g0473(.A1(new_n665), .A2(new_n669), .A3(new_n673), .ZN(new_n674));
  AND3_X1   g0474(.A1(new_n674), .A2(KEYINPUT31), .A3(new_n630), .ZN(new_n675));
  AOI21_X1  g0475(.A(KEYINPUT31), .B1(new_n674), .B2(new_n630), .ZN(new_n676));
  NOR2_X1   g0476(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  AOI21_X1  g0477(.A(new_n659), .B1(new_n663), .B2(new_n677), .ZN(new_n678));
  NOR2_X1   g0478(.A1(new_n658), .A2(new_n678), .ZN(new_n679));
  OAI21_X1  g0479(.A(new_n651), .B1(new_n679), .B2(G1), .ZN(G364));
  NOR2_X1   g0480(.A1(new_n300), .A2(G20), .ZN(new_n681));
  AOI21_X1  g0481(.A(new_n210), .B1(new_n681), .B2(G45), .ZN(new_n682));
  INV_X1    g0482(.A(new_n682), .ZN(new_n683));
  NOR2_X1   g0483(.A1(new_n646), .A2(new_n683), .ZN(new_n684));
  INV_X1    g0484(.A(new_n684), .ZN(new_n685));
  NOR2_X1   g0485(.A1(new_n645), .A2(new_n264), .ZN(new_n686));
  AOI22_X1  g0486(.A1(G355), .A2(new_n686), .B1(new_n574), .B2(new_n645), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n214), .A2(new_n264), .ZN(new_n688));
  XOR2_X1   g0488(.A(new_n688), .B(KEYINPUT90), .Z(new_n689));
  OAI21_X1  g0489(.A(new_n689), .B1(G45), .B2(new_n221), .ZN(new_n690));
  NOR2_X1   g0490(.A1(new_n249), .A2(new_n462), .ZN(new_n691));
  OAI21_X1  g0491(.A(new_n687), .B1(new_n690), .B2(new_n691), .ZN(new_n692));
  NOR2_X1   g0492(.A1(G13), .A2(G33), .ZN(new_n693));
  INV_X1    g0493(.A(new_n693), .ZN(new_n694));
  NOR2_X1   g0494(.A1(new_n694), .A2(G20), .ZN(new_n695));
  AOI21_X1  g0495(.A(new_n217), .B1(G20), .B2(new_n353), .ZN(new_n696));
  NOR2_X1   g0496(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  AOI21_X1  g0497(.A(new_n685), .B1(new_n692), .B2(new_n697), .ZN(new_n698));
  INV_X1    g0498(.A(new_n696), .ZN(new_n699));
  NOR2_X1   g0499(.A1(new_n211), .A2(new_n334), .ZN(new_n700));
  NOR2_X1   g0500(.A1(G190), .A2(G200), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  NOR2_X1   g0502(.A1(new_n211), .A2(G179), .ZN(new_n703));
  NAND3_X1  g0503(.A1(new_n703), .A2(G190), .A3(G200), .ZN(new_n704));
  OAI221_X1 g0504(.A(new_n273), .B1(new_n702), .B2(new_n348), .C1(new_n225), .C2(new_n704), .ZN(new_n705));
  NAND3_X1  g0505(.A1(new_n703), .A2(new_n358), .A3(G200), .ZN(new_n706));
  NOR2_X1   g0506(.A1(new_n706), .A2(new_n327), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n700), .A2(G200), .ZN(new_n708));
  NOR2_X1   g0508(.A1(new_n708), .A2(G190), .ZN(new_n709));
  AOI21_X1  g0509(.A(new_n707), .B1(G68), .B2(new_n709), .ZN(new_n710));
  NOR2_X1   g0510(.A1(new_n708), .A2(new_n358), .ZN(new_n711));
  INV_X1    g0511(.A(new_n711), .ZN(new_n712));
  NOR2_X1   g0512(.A1(new_n358), .A2(G200), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n713), .A2(new_n334), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n714), .A2(G20), .ZN(new_n715));
  INV_X1    g0515(.A(new_n715), .ZN(new_n716));
  OAI221_X1 g0516(.A(new_n710), .B1(new_n202), .B2(new_n712), .C1(new_n482), .C2(new_n716), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n700), .A2(new_n713), .ZN(new_n718));
  INV_X1    g0518(.A(KEYINPUT91), .ZN(new_n719));
  NAND2_X1  g0519(.A1(new_n718), .A2(new_n719), .ZN(new_n720));
  INV_X1    g0520(.A(new_n720), .ZN(new_n721));
  NOR2_X1   g0521(.A1(new_n718), .A2(new_n719), .ZN(new_n722));
  NOR2_X1   g0522(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  INV_X1    g0523(.A(new_n723), .ZN(new_n724));
  AOI211_X1 g0524(.A(new_n705), .B(new_n717), .C1(G58), .C2(new_n724), .ZN(new_n725));
  NAND2_X1  g0525(.A1(new_n703), .A2(new_n701), .ZN(new_n726));
  OR2_X1    g0526(.A1(new_n726), .A2(KEYINPUT92), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n726), .A2(KEYINPUT92), .ZN(new_n728));
  NAND2_X1  g0528(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  XOR2_X1   g0529(.A(KEYINPUT93), .B(G159), .Z(new_n730));
  NOR2_X1   g0530(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  XNOR2_X1  g0531(.A(new_n731), .B(KEYINPUT32), .ZN(new_n732));
  INV_X1    g0532(.A(G283), .ZN(new_n733));
  NOR2_X1   g0533(.A1(new_n706), .A2(new_n733), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n711), .A2(G326), .ZN(new_n735));
  OAI21_X1  g0535(.A(new_n735), .B1(new_n523), .B2(new_n716), .ZN(new_n736));
  XNOR2_X1  g0536(.A(KEYINPUT33), .B(G317), .ZN(new_n737));
  AOI211_X1 g0537(.A(new_n734), .B(new_n736), .C1(new_n709), .C2(new_n737), .ZN(new_n738));
  INV_X1    g0538(.A(G311), .ZN(new_n739));
  OAI221_X1 g0539(.A(new_n264), .B1(new_n702), .B2(new_n739), .C1(new_n585), .C2(new_n704), .ZN(new_n740));
  INV_X1    g0540(.A(G322), .ZN(new_n741));
  NOR2_X1   g0541(.A1(new_n723), .A2(new_n741), .ZN(new_n742));
  INV_X1    g0542(.A(new_n729), .ZN(new_n743));
  AOI211_X1 g0543(.A(new_n740), .B(new_n742), .C1(G329), .C2(new_n743), .ZN(new_n744));
  AOI22_X1  g0544(.A1(new_n725), .A2(new_n732), .B1(new_n738), .B2(new_n744), .ZN(new_n745));
  INV_X1    g0545(.A(new_n695), .ZN(new_n746));
  OAI221_X1 g0546(.A(new_n698), .B1(new_n699), .B2(new_n745), .C1(new_n634), .C2(new_n746), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n633), .A2(new_n659), .ZN(new_n748));
  XOR2_X1   g0548(.A(new_n748), .B(KEYINPUT89), .Z(new_n749));
  NAND2_X1  g0549(.A1(new_n634), .A2(G330), .ZN(new_n750));
  NAND2_X1  g0550(.A1(new_n750), .A2(new_n685), .ZN(new_n751));
  OAI21_X1  g0551(.A(new_n747), .B1(new_n749), .B2(new_n751), .ZN(G396));
  INV_X1    g0552(.A(new_n355), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n753), .A2(new_n653), .ZN(new_n754));
  INV_X1    g0554(.A(new_n754), .ZN(new_n755));
  NAND2_X1  g0555(.A1(new_n352), .A2(new_n630), .ZN(new_n756));
  OAI21_X1  g0556(.A(new_n756), .B1(new_n359), .B2(new_n360), .ZN(new_n757));
  AOI21_X1  g0557(.A(new_n755), .B1(new_n757), .B2(new_n355), .ZN(new_n758));
  INV_X1    g0558(.A(new_n758), .ZN(new_n759));
  NAND2_X1  g0559(.A1(new_n654), .A2(new_n759), .ZN(new_n760));
  AOI21_X1  g0560(.A(new_n630), .B1(new_n616), .B2(new_n607), .ZN(new_n761));
  NAND2_X1  g0561(.A1(new_n761), .A2(new_n758), .ZN(new_n762));
  NAND2_X1  g0562(.A1(new_n760), .A2(new_n762), .ZN(new_n763));
  INV_X1    g0563(.A(new_n678), .ZN(new_n764));
  AOI21_X1  g0564(.A(new_n684), .B1(new_n763), .B2(new_n764), .ZN(new_n765));
  NAND3_X1  g0565(.A1(new_n760), .A2(new_n678), .A3(new_n762), .ZN(new_n766));
  AND2_X1   g0566(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  NOR2_X1   g0567(.A1(new_n696), .A2(new_n693), .ZN(new_n768));
  INV_X1    g0568(.A(new_n768), .ZN(new_n769));
  OAI21_X1  g0569(.A(new_n684), .B1(G77), .B2(new_n769), .ZN(new_n770));
  INV_X1    g0570(.A(new_n709), .ZN(new_n771));
  OAI22_X1  g0571(.A1(new_n733), .A2(new_n771), .B1(new_n712), .B2(new_n585), .ZN(new_n772));
  INV_X1    g0572(.A(new_n706), .ZN(new_n773));
  AOI21_X1  g0573(.A(new_n772), .B1(G87), .B2(new_n773), .ZN(new_n774));
  OAI21_X1  g0574(.A(new_n264), .B1(new_n704), .B2(new_n327), .ZN(new_n775));
  XNOR2_X1  g0575(.A(new_n775), .B(KEYINPUT94), .ZN(new_n776));
  NAND2_X1  g0576(.A1(new_n724), .A2(G294), .ZN(new_n777));
  OAI22_X1  g0577(.A1(new_n716), .A2(new_n482), .B1(new_n702), .B2(new_n574), .ZN(new_n778));
  AOI21_X1  g0578(.A(new_n778), .B1(new_n743), .B2(G311), .ZN(new_n779));
  NAND4_X1  g0579(.A1(new_n774), .A2(new_n776), .A3(new_n777), .A4(new_n779), .ZN(new_n780));
  OAI21_X1  g0580(.A(new_n273), .B1(new_n704), .B2(new_n202), .ZN(new_n781));
  OAI22_X1  g0581(.A1(new_n716), .A2(new_n283), .B1(new_n706), .B2(new_n223), .ZN(new_n782));
  AOI211_X1 g0582(.A(new_n781), .B(new_n782), .C1(G132), .C2(new_n743), .ZN(new_n783));
  INV_X1    g0583(.A(new_n730), .ZN(new_n784));
  INV_X1    g0584(.A(new_n702), .ZN(new_n785));
  AOI22_X1  g0585(.A1(new_n711), .A2(G137), .B1(new_n784), .B2(new_n785), .ZN(new_n786));
  INV_X1    g0586(.A(G150), .ZN(new_n787));
  INV_X1    g0587(.A(G143), .ZN(new_n788));
  OAI221_X1 g0588(.A(new_n786), .B1(new_n787), .B2(new_n771), .C1(new_n723), .C2(new_n788), .ZN(new_n789));
  INV_X1    g0589(.A(new_n789), .ZN(new_n790));
  OAI21_X1  g0590(.A(new_n783), .B1(new_n790), .B2(KEYINPUT34), .ZN(new_n791));
  INV_X1    g0591(.A(KEYINPUT34), .ZN(new_n792));
  NOR2_X1   g0592(.A1(new_n789), .A2(new_n792), .ZN(new_n793));
  OAI21_X1  g0593(.A(new_n780), .B1(new_n791), .B2(new_n793), .ZN(new_n794));
  AOI21_X1  g0594(.A(new_n770), .B1(new_n794), .B2(new_n696), .ZN(new_n795));
  OAI21_X1  g0595(.A(new_n795), .B1(new_n758), .B2(new_n694), .ZN(new_n796));
  XNOR2_X1  g0596(.A(new_n796), .B(KEYINPUT95), .ZN(new_n797));
  OR2_X1    g0597(.A1(new_n767), .A2(new_n797), .ZN(G384));
  AOI211_X1 g0598(.A(new_n574), .B(new_n219), .C1(new_n490), .C2(KEYINPUT35), .ZN(new_n799));
  OAI21_X1  g0599(.A(new_n799), .B1(KEYINPUT35), .B2(new_n490), .ZN(new_n800));
  XOR2_X1   g0600(.A(new_n800), .B(KEYINPUT36), .Z(new_n801));
  OR3_X1    g0601(.A1(new_n221), .A2(new_n348), .A3(new_n426), .ZN(new_n802));
  XOR2_X1   g0602(.A(new_n245), .B(KEYINPUT96), .Z(new_n803));
  AOI211_X1 g0603(.A(new_n210), .B(G13), .C1(new_n802), .C2(new_n803), .ZN(new_n804));
  NOR2_X1   g0604(.A1(new_n801), .A2(new_n804), .ZN(new_n805));
  AOI21_X1  g0605(.A(new_n755), .B1(new_n761), .B2(new_n758), .ZN(new_n806));
  INV_X1    g0606(.A(new_n806), .ZN(new_n807));
  INV_X1    g0607(.A(KEYINPUT38), .ZN(new_n808));
  INV_X1    g0608(.A(KEYINPUT99), .ZN(new_n809));
  INV_X1    g0609(.A(new_n445), .ZN(new_n810));
  OAI21_X1  g0610(.A(new_n428), .B1(new_n434), .B2(new_n436), .ZN(new_n811));
  INV_X1    g0611(.A(KEYINPUT98), .ZN(new_n812));
  NAND2_X1  g0612(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  OAI211_X1 g0613(.A(KEYINPUT98), .B(new_n428), .C1(new_n434), .C2(new_n436), .ZN(new_n814));
  NAND3_X1  g0614(.A1(new_n813), .A2(new_n440), .A3(new_n814), .ZN(new_n815));
  NAND2_X1  g0615(.A1(new_n437), .A2(new_n281), .ZN(new_n816));
  INV_X1    g0616(.A(new_n816), .ZN(new_n817));
  AOI21_X1  g0617(.A(new_n810), .B1(new_n815), .B2(new_n817), .ZN(new_n818));
  OAI21_X1  g0618(.A(new_n809), .B1(new_n818), .B2(new_n628), .ZN(new_n819));
  INV_X1    g0619(.A(new_n628), .ZN(new_n820));
  AOI21_X1  g0620(.A(KEYINPUT16), .B1(new_n811), .B2(new_n812), .ZN(new_n821));
  AOI21_X1  g0621(.A(new_n816), .B1(new_n821), .B2(new_n814), .ZN(new_n822));
  OAI211_X1 g0622(.A(KEYINPUT99), .B(new_n820), .C1(new_n822), .C2(new_n810), .ZN(new_n823));
  NAND2_X1  g0623(.A1(new_n819), .A2(new_n823), .ZN(new_n824));
  NAND2_X1  g0624(.A1(new_n453), .A2(new_n824), .ZN(new_n825));
  INV_X1    g0625(.A(new_n825), .ZN(new_n826));
  INV_X1    g0626(.A(new_n425), .ZN(new_n827));
  OAI21_X1  g0627(.A(new_n827), .B1(new_n822), .B2(new_n810), .ZN(new_n828));
  NAND4_X1  g0628(.A1(new_n819), .A2(new_n451), .A3(new_n823), .A4(new_n828), .ZN(new_n829));
  INV_X1    g0629(.A(new_n451), .ZN(new_n830));
  NOR2_X1   g0630(.A1(new_n830), .A2(new_n446), .ZN(new_n831));
  INV_X1    g0631(.A(KEYINPUT37), .ZN(new_n832));
  NAND2_X1  g0632(.A1(new_n442), .A2(new_n445), .ZN(new_n833));
  NAND2_X1  g0633(.A1(new_n833), .A2(new_n820), .ZN(new_n834));
  NAND4_X1  g0634(.A1(new_n831), .A2(KEYINPUT100), .A3(new_n832), .A4(new_n834), .ZN(new_n835));
  NAND2_X1  g0635(.A1(new_n833), .A2(new_n827), .ZN(new_n836));
  NAND4_X1  g0636(.A1(new_n836), .A2(new_n834), .A3(new_n832), .A4(new_n451), .ZN(new_n837));
  INV_X1    g0637(.A(KEYINPUT100), .ZN(new_n838));
  NAND2_X1  g0638(.A1(new_n837), .A2(new_n838), .ZN(new_n839));
  AOI22_X1  g0639(.A1(new_n829), .A2(KEYINPUT37), .B1(new_n835), .B2(new_n839), .ZN(new_n840));
  OAI21_X1  g0640(.A(new_n808), .B1(new_n826), .B2(new_n840), .ZN(new_n841));
  NAND2_X1  g0641(.A1(new_n829), .A2(KEYINPUT37), .ZN(new_n842));
  NAND2_X1  g0642(.A1(new_n835), .A2(new_n839), .ZN(new_n843));
  NAND2_X1  g0643(.A1(new_n842), .A2(new_n843), .ZN(new_n844));
  NAND3_X1  g0644(.A1(new_n844), .A2(KEYINPUT38), .A3(new_n825), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n841), .A2(new_n845), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n411), .A2(new_n630), .ZN(new_n847));
  OAI21_X1  g0647(.A(new_n847), .B1(new_n417), .B2(KEYINPUT97), .ZN(new_n848));
  NOR3_X1   g0648(.A1(new_n619), .A2(new_n398), .A3(new_n847), .ZN(new_n849));
  NAND3_X1  g0649(.A1(new_n412), .A2(KEYINPUT97), .A3(new_n416), .ZN(new_n850));
  NAND2_X1  g0650(.A1(new_n849), .A2(new_n850), .ZN(new_n851));
  AND2_X1   g0651(.A1(new_n848), .A2(new_n851), .ZN(new_n852));
  NAND3_X1  g0652(.A1(new_n807), .A2(new_n846), .A3(new_n852), .ZN(new_n853));
  NAND2_X1  g0653(.A1(new_n618), .A2(new_n628), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  INV_X1    g0655(.A(KEYINPUT39), .ZN(new_n856));
  AOI21_X1  g0656(.A(new_n832), .B1(new_n831), .B2(new_n834), .ZN(new_n857));
  AOI21_X1  g0657(.A(new_n857), .B1(new_n839), .B2(new_n835), .ZN(new_n858));
  AOI21_X1  g0658(.A(new_n834), .B1(new_n447), .B2(new_n452), .ZN(new_n859));
  OAI21_X1  g0659(.A(new_n808), .B1(new_n858), .B2(new_n859), .ZN(new_n860));
  NAND3_X1  g0660(.A1(new_n845), .A2(new_n856), .A3(new_n860), .ZN(new_n861));
  INV_X1    g0661(.A(KEYINPUT102), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  NAND4_X1  g0663(.A1(new_n845), .A2(KEYINPUT102), .A3(new_n860), .A4(new_n856), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  AOI21_X1  g0665(.A(KEYINPUT101), .B1(new_n846), .B2(KEYINPUT39), .ZN(new_n866));
  INV_X1    g0666(.A(KEYINPUT101), .ZN(new_n867));
  AOI211_X1 g0667(.A(new_n867), .B(new_n856), .C1(new_n841), .C2(new_n845), .ZN(new_n868));
  OAI21_X1  g0668(.A(new_n865), .B1(new_n866), .B2(new_n868), .ZN(new_n869));
  NOR2_X1   g0669(.A1(new_n412), .A2(new_n630), .ZN(new_n870));
  AOI21_X1  g0670(.A(new_n855), .B1(new_n869), .B2(new_n870), .ZN(new_n871));
  INV_X1    g0671(.A(KEYINPUT103), .ZN(new_n872));
  NAND3_X1  g0672(.A1(new_n456), .A2(new_n658), .A3(new_n872), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n607), .A2(new_n656), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n874), .A2(new_n653), .ZN(new_n875));
  INV_X1    g0675(.A(KEYINPUT29), .ZN(new_n876));
  INV_X1    g0676(.A(new_n655), .ZN(new_n877));
  OAI22_X1  g0677(.A1(new_n875), .A2(new_n876), .B1(new_n761), .B2(new_n877), .ZN(new_n878));
  OAI21_X1  g0678(.A(KEYINPUT103), .B1(new_n878), .B2(new_n455), .ZN(new_n879));
  AOI21_X1  g0679(.A(new_n623), .B1(new_n873), .B2(new_n879), .ZN(new_n880));
  XNOR2_X1  g0680(.A(new_n871), .B(new_n880), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n663), .A2(new_n677), .ZN(new_n882));
  NAND4_X1  g0682(.A1(new_n882), .A2(new_n848), .A3(new_n851), .A4(new_n758), .ZN(new_n883));
  INV_X1    g0683(.A(new_n883), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n846), .A2(new_n884), .ZN(new_n885));
  INV_X1    g0685(.A(KEYINPUT40), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n845), .A2(new_n860), .ZN(new_n888));
  NAND3_X1  g0688(.A1(new_n884), .A2(new_n888), .A3(KEYINPUT40), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n887), .A2(new_n889), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n456), .A2(new_n882), .ZN(new_n891));
  AOI21_X1  g0691(.A(new_n659), .B1(new_n890), .B2(new_n891), .ZN(new_n892));
  OAI21_X1  g0692(.A(new_n892), .B1(new_n891), .B2(new_n890), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n881), .A2(new_n893), .ZN(new_n894));
  OAI21_X1  g0694(.A(new_n894), .B1(new_n210), .B2(new_n681), .ZN(new_n895));
  NOR2_X1   g0695(.A1(new_n881), .A2(new_n893), .ZN(new_n896));
  OAI21_X1  g0696(.A(new_n805), .B1(new_n895), .B2(new_n896), .ZN(G367));
  NAND2_X1  g0697(.A1(new_n689), .A2(new_n240), .ZN(new_n898));
  NOR2_X1   g0698(.A1(new_n214), .A2(new_n339), .ZN(new_n899));
  NOR3_X1   g0699(.A1(new_n899), .A2(new_n695), .A3(new_n696), .ZN(new_n900));
  AOI21_X1  g0700(.A(new_n685), .B1(new_n898), .B2(new_n900), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n555), .A2(new_n630), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n608), .A2(new_n902), .ZN(new_n903));
  OAI21_X1  g0703(.A(new_n903), .B1(new_n565), .B2(new_n902), .ZN(new_n904));
  AOI22_X1  g0704(.A1(new_n724), .A2(G303), .B1(new_n743), .B2(G317), .ZN(new_n905));
  OAI22_X1  g0705(.A1(new_n712), .A2(new_n739), .B1(new_n706), .B2(new_n482), .ZN(new_n906));
  AOI21_X1  g0706(.A(new_n906), .B1(G294), .B2(new_n709), .ZN(new_n907));
  INV_X1    g0707(.A(KEYINPUT46), .ZN(new_n908));
  OAI21_X1  g0708(.A(new_n908), .B1(new_n704), .B2(new_n574), .ZN(new_n909));
  XOR2_X1   g0709(.A(new_n909), .B(KEYINPUT105), .Z(new_n910));
  OAI21_X1  g0710(.A(new_n264), .B1(new_n702), .B2(new_n733), .ZN(new_n911));
  NOR3_X1   g0711(.A1(new_n704), .A2(new_n908), .A3(new_n574), .ZN(new_n912));
  AOI211_X1 g0712(.A(new_n911), .B(new_n912), .C1(G107), .C2(new_n715), .ZN(new_n913));
  NAND4_X1  g0713(.A1(new_n905), .A2(new_n907), .A3(new_n910), .A4(new_n913), .ZN(new_n914));
  XOR2_X1   g0714(.A(new_n914), .B(KEYINPUT106), .Z(new_n915));
  XNOR2_X1  g0715(.A(KEYINPUT107), .B(G137), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n743), .A2(new_n916), .ZN(new_n917));
  OAI21_X1  g0717(.A(new_n917), .B1(new_n283), .B2(new_n704), .ZN(new_n918));
  NOR2_X1   g0718(.A1(new_n918), .A2(KEYINPUT108), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n918), .A2(KEYINPUT108), .ZN(new_n920));
  OAI22_X1  g0720(.A1(new_n771), .A2(new_n730), .B1(new_n712), .B2(new_n788), .ZN(new_n921));
  NOR2_X1   g0721(.A1(new_n706), .A2(new_n348), .ZN(new_n922));
  NOR2_X1   g0722(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n724), .A2(G150), .ZN(new_n924));
  NOR2_X1   g0724(.A1(new_n716), .A2(new_n223), .ZN(new_n925));
  AOI211_X1 g0725(.A(new_n264), .B(new_n925), .C1(G50), .C2(new_n785), .ZN(new_n926));
  NAND4_X1  g0726(.A1(new_n920), .A2(new_n923), .A3(new_n924), .A4(new_n926), .ZN(new_n927));
  OAI21_X1  g0727(.A(new_n915), .B1(new_n919), .B2(new_n927), .ZN(new_n928));
  XOR2_X1   g0728(.A(new_n928), .B(KEYINPUT47), .Z(new_n929));
  OAI221_X1 g0729(.A(new_n901), .B1(new_n746), .B2(new_n904), .C1(new_n929), .C2(new_n699), .ZN(new_n930));
  OAI211_X1 g0730(.A(new_n496), .B(new_n498), .C1(new_n494), .C2(new_n653), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n609), .A2(new_n630), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n931), .A2(new_n932), .ZN(new_n933));
  NAND3_X1  g0733(.A1(new_n643), .A2(new_n635), .A3(new_n933), .ZN(new_n934));
  XOR2_X1   g0734(.A(new_n934), .B(KEYINPUT45), .Z(new_n935));
  AOI21_X1  g0735(.A(new_n933), .B1(new_n643), .B2(new_n635), .ZN(new_n936));
  NOR2_X1   g0736(.A1(new_n936), .A2(KEYINPUT44), .ZN(new_n937));
  AND2_X1   g0737(.A1(new_n936), .A2(KEYINPUT44), .ZN(new_n938));
  OAI211_X1 g0738(.A(new_n935), .B(new_n641), .C1(new_n937), .C2(new_n938), .ZN(new_n939));
  INV_X1    g0739(.A(new_n641), .ZN(new_n940));
  NOR2_X1   g0740(.A1(new_n938), .A2(new_n937), .ZN(new_n941));
  XNOR2_X1  g0741(.A(new_n934), .B(KEYINPUT45), .ZN(new_n942));
  OAI21_X1  g0742(.A(new_n940), .B1(new_n941), .B2(new_n942), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n939), .A2(new_n943), .ZN(new_n944));
  XNOR2_X1  g0744(.A(new_n640), .B(new_n642), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n750), .A2(KEYINPUT104), .ZN(new_n946));
  XNOR2_X1  g0746(.A(new_n945), .B(new_n946), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n947), .A2(new_n679), .ZN(new_n948));
  OAI21_X1  g0748(.A(new_n679), .B1(new_n944), .B2(new_n948), .ZN(new_n949));
  XOR2_X1   g0749(.A(new_n646), .B(KEYINPUT41), .Z(new_n950));
  INV_X1    g0750(.A(new_n950), .ZN(new_n951));
  AOI21_X1  g0751(.A(new_n683), .B1(new_n949), .B2(new_n951), .ZN(new_n952));
  NAND3_X1  g0752(.A1(new_n640), .A2(new_n642), .A3(new_n933), .ZN(new_n953));
  OAI21_X1  g0753(.A(new_n496), .B1(new_n931), .B2(new_n573), .ZN(new_n954));
  AOI22_X1  g0754(.A1(new_n953), .A2(KEYINPUT42), .B1(new_n653), .B2(new_n954), .ZN(new_n955));
  OAI21_X1  g0755(.A(new_n955), .B1(KEYINPUT42), .B2(new_n953), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n904), .A2(KEYINPUT43), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n956), .A2(new_n957), .ZN(new_n958));
  NOR2_X1   g0758(.A1(new_n904), .A2(KEYINPUT43), .ZN(new_n959));
  XNOR2_X1  g0759(.A(new_n958), .B(new_n959), .ZN(new_n960));
  INV_X1    g0760(.A(new_n933), .ZN(new_n961));
  NOR2_X1   g0761(.A1(new_n641), .A2(new_n961), .ZN(new_n962));
  XOR2_X1   g0762(.A(new_n960), .B(new_n962), .Z(new_n963));
  OAI21_X1  g0763(.A(new_n930), .B1(new_n952), .B2(new_n963), .ZN(G387));
  NAND2_X1  g0764(.A1(new_n947), .A2(new_n683), .ZN(new_n965));
  INV_X1    g0765(.A(new_n689), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n287), .A2(new_n202), .ZN(new_n967));
  XNOR2_X1  g0767(.A(new_n967), .B(KEYINPUT50), .ZN(new_n968));
  INV_X1    g0768(.A(new_n968), .ZN(new_n969));
  INV_X1    g0769(.A(new_n648), .ZN(new_n970));
  AOI211_X1 g0770(.A(G45), .B(new_n970), .C1(G68), .C2(G77), .ZN(new_n971));
  AOI21_X1  g0771(.A(new_n966), .B1(new_n969), .B2(new_n971), .ZN(new_n972));
  OAI21_X1  g0772(.A(new_n972), .B1(new_n462), .B2(new_n237), .ZN(new_n973));
  AOI22_X1  g0773(.A1(new_n686), .A2(new_n970), .B1(new_n327), .B2(new_n645), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n973), .A2(new_n974), .ZN(new_n975));
  AOI21_X1  g0775(.A(new_n685), .B1(new_n975), .B2(new_n697), .ZN(new_n976));
  NOR2_X1   g0776(.A1(new_n771), .A2(new_n443), .ZN(new_n977));
  AOI21_X1  g0777(.A(new_n977), .B1(new_n724), .B2(G50), .ZN(new_n978));
  INV_X1    g0778(.A(new_n563), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n979), .A2(new_n715), .ZN(new_n980));
  OAI211_X1 g0780(.A(new_n978), .B(new_n980), .C1(new_n787), .C2(new_n729), .ZN(new_n981));
  OAI221_X1 g0781(.A(new_n273), .B1(new_n702), .B2(new_n223), .C1(new_n482), .C2(new_n706), .ZN(new_n982));
  INV_X1    g0782(.A(G159), .ZN(new_n983));
  NOR2_X1   g0783(.A1(new_n712), .A2(new_n983), .ZN(new_n984));
  NOR2_X1   g0784(.A1(new_n704), .A2(new_n348), .ZN(new_n985));
  NOR4_X1   g0785(.A1(new_n981), .A2(new_n982), .A3(new_n984), .A4(new_n985), .ZN(new_n986));
  OAI21_X1  g0786(.A(new_n264), .B1(new_n706), .B2(new_n574), .ZN(new_n987));
  AOI22_X1  g0787(.A1(new_n709), .A2(G311), .B1(new_n785), .B2(G303), .ZN(new_n988));
  INV_X1    g0788(.A(G317), .ZN(new_n989));
  OAI221_X1 g0789(.A(new_n988), .B1(new_n741), .B2(new_n712), .C1(new_n723), .C2(new_n989), .ZN(new_n990));
  INV_X1    g0790(.A(KEYINPUT48), .ZN(new_n991));
  OR2_X1    g0791(.A1(new_n990), .A2(new_n991), .ZN(new_n992));
  NAND2_X1  g0792(.A1(new_n990), .A2(new_n991), .ZN(new_n993));
  INV_X1    g0793(.A(new_n704), .ZN(new_n994));
  AOI22_X1  g0794(.A1(new_n994), .A2(G294), .B1(new_n715), .B2(G283), .ZN(new_n995));
  NAND3_X1  g0795(.A1(new_n992), .A2(new_n993), .A3(new_n995), .ZN(new_n996));
  INV_X1    g0796(.A(KEYINPUT49), .ZN(new_n997));
  NOR2_X1   g0797(.A1(new_n996), .A2(new_n997), .ZN(new_n998));
  AOI211_X1 g0798(.A(new_n987), .B(new_n998), .C1(G326), .C2(new_n743), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n996), .A2(new_n997), .ZN(new_n1000));
  AOI21_X1  g0800(.A(new_n986), .B1(new_n999), .B2(new_n1000), .ZN(new_n1001));
  OAI21_X1  g0801(.A(new_n976), .B1(new_n1001), .B2(new_n699), .ZN(new_n1002));
  INV_X1    g0802(.A(KEYINPUT109), .ZN(new_n1003));
  NOR2_X1   g0803(.A1(new_n1002), .A2(new_n1003), .ZN(new_n1004));
  NAND2_X1  g0804(.A1(new_n1002), .A2(new_n1003), .ZN(new_n1005));
  OAI21_X1  g0805(.A(new_n1005), .B1(new_n640), .B2(new_n746), .ZN(new_n1006));
  NAND2_X1  g0806(.A1(new_n948), .A2(new_n646), .ZN(new_n1007));
  NOR2_X1   g0807(.A1(new_n947), .A2(new_n679), .ZN(new_n1008));
  OAI221_X1 g0808(.A(new_n965), .B1(new_n1004), .B2(new_n1006), .C1(new_n1007), .C2(new_n1008), .ZN(G393));
  NAND3_X1  g0809(.A1(new_n939), .A2(new_n683), .A3(new_n943), .ZN(new_n1010));
  OAI221_X1 g0810(.A(new_n697), .B1(new_n482), .B2(new_n214), .C1(new_n966), .C2(new_n244), .ZN(new_n1011));
  AND2_X1   g0811(.A1(new_n1011), .A2(new_n684), .ZN(new_n1012));
  OAI22_X1  g0812(.A1(new_n771), .A2(new_n585), .B1(new_n704), .B2(new_n733), .ZN(new_n1013));
  AOI211_X1 g0813(.A(new_n273), .B(new_n707), .C1(G294), .C2(new_n785), .ZN(new_n1014));
  OAI21_X1  g0814(.A(new_n1014), .B1(new_n741), .B2(new_n729), .ZN(new_n1015));
  AOI211_X1 g0815(.A(new_n1013), .B(new_n1015), .C1(G116), .C2(new_n715), .ZN(new_n1016));
  OAI22_X1  g0816(.A1(new_n723), .A2(new_n739), .B1(new_n989), .B2(new_n712), .ZN(new_n1017));
  XNOR2_X1  g0817(.A(new_n1017), .B(KEYINPUT52), .ZN(new_n1018));
  OAI22_X1  g0818(.A1(new_n723), .A2(new_n983), .B1(new_n787), .B2(new_n712), .ZN(new_n1019));
  XNOR2_X1  g0819(.A(new_n1019), .B(KEYINPUT51), .ZN(new_n1020));
  AOI21_X1  g0820(.A(new_n264), .B1(new_n785), .B2(new_n287), .ZN(new_n1021));
  OAI221_X1 g0821(.A(new_n1021), .B1(new_n225), .B2(new_n706), .C1(new_n729), .C2(new_n788), .ZN(new_n1022));
  NOR2_X1   g0822(.A1(new_n716), .A2(new_n348), .ZN(new_n1023));
  OAI22_X1  g0823(.A1(new_n771), .A2(new_n202), .B1(new_n704), .B2(new_n223), .ZN(new_n1024));
  NOR3_X1   g0824(.A1(new_n1022), .A2(new_n1023), .A3(new_n1024), .ZN(new_n1025));
  AOI22_X1  g0825(.A1(new_n1016), .A2(new_n1018), .B1(new_n1020), .B2(new_n1025), .ZN(new_n1026));
  XNOR2_X1  g0826(.A(new_n1026), .B(KEYINPUT110), .ZN(new_n1027));
  OAI221_X1 g0827(.A(new_n1012), .B1(new_n746), .B2(new_n933), .C1(new_n1027), .C2(new_n699), .ZN(new_n1028));
  AND2_X1   g0828(.A1(new_n944), .A2(new_n948), .ZN(new_n1029));
  OAI21_X1  g0829(.A(new_n646), .B1(new_n944), .B2(new_n948), .ZN(new_n1030));
  OAI211_X1 g0830(.A(new_n1010), .B(new_n1028), .C1(new_n1029), .C2(new_n1030), .ZN(G390));
  INV_X1    g0831(.A(new_n870), .ZN(new_n1032));
  NAND2_X1  g0832(.A1(new_n848), .A2(new_n851), .ZN(new_n1033));
  OAI21_X1  g0833(.A(new_n1032), .B1(new_n806), .B2(new_n1033), .ZN(new_n1034));
  OAI211_X1 g0834(.A(new_n865), .B(new_n1034), .C1(new_n866), .C2(new_n868), .ZN(new_n1035));
  NAND2_X1  g0835(.A1(new_n757), .A2(new_n355), .ZN(new_n1036));
  AOI21_X1  g0836(.A(new_n755), .B1(new_n657), .B2(new_n1036), .ZN(new_n1037));
  OAI211_X1 g0837(.A(new_n1032), .B(new_n888), .C1(new_n1037), .C2(new_n1033), .ZN(new_n1038));
  NAND2_X1  g0838(.A1(new_n1035), .A2(new_n1038), .ZN(new_n1039));
  NAND4_X1  g0839(.A1(new_n678), .A2(new_n758), .A3(new_n848), .A4(new_n851), .ZN(new_n1040));
  INV_X1    g0840(.A(KEYINPUT111), .ZN(new_n1041));
  NAND2_X1  g0841(.A1(new_n1040), .A2(new_n1041), .ZN(new_n1042));
  NAND4_X1  g0842(.A1(new_n852), .A2(KEYINPUT111), .A3(new_n678), .A4(new_n758), .ZN(new_n1043));
  NAND2_X1  g0843(.A1(new_n1042), .A2(new_n1043), .ZN(new_n1044));
  INV_X1    g0844(.A(new_n1044), .ZN(new_n1045));
  NAND2_X1  g0845(.A1(new_n1039), .A2(new_n1045), .ZN(new_n1046));
  AND2_X1   g0846(.A1(new_n1038), .A2(new_n1040), .ZN(new_n1047));
  AND3_X1   g0847(.A1(new_n1035), .A2(KEYINPUT112), .A3(new_n1047), .ZN(new_n1048));
  AOI21_X1  g0848(.A(KEYINPUT112), .B1(new_n1035), .B2(new_n1047), .ZN(new_n1049));
  OAI21_X1  g0849(.A(new_n1046), .B1(new_n1048), .B2(new_n1049), .ZN(new_n1050));
  OAI21_X1  g0850(.A(KEYINPUT114), .B1(new_n1050), .B2(new_n682), .ZN(new_n1051));
  AOI21_X1  g0851(.A(new_n1044), .B1(new_n1035), .B2(new_n1038), .ZN(new_n1052));
  NAND2_X1  g0852(.A1(new_n1035), .A2(new_n1047), .ZN(new_n1053));
  INV_X1    g0853(.A(KEYINPUT112), .ZN(new_n1054));
  NAND2_X1  g0854(.A1(new_n1053), .A2(new_n1054), .ZN(new_n1055));
  NAND3_X1  g0855(.A1(new_n1035), .A2(KEYINPUT112), .A3(new_n1047), .ZN(new_n1056));
  AOI21_X1  g0856(.A(new_n1052), .B1(new_n1055), .B2(new_n1056), .ZN(new_n1057));
  INV_X1    g0857(.A(KEYINPUT114), .ZN(new_n1058));
  NAND3_X1  g0858(.A1(new_n1057), .A2(new_n1058), .A3(new_n683), .ZN(new_n1059));
  NAND2_X1  g0859(.A1(new_n1051), .A2(new_n1059), .ZN(new_n1060));
  AOI22_X1  g0860(.A1(new_n678), .A2(new_n758), .B1(new_n848), .B2(new_n851), .ZN(new_n1061));
  INV_X1    g0861(.A(new_n1061), .ZN(new_n1062));
  NAND3_X1  g0862(.A1(new_n1062), .A2(new_n1040), .A3(new_n1037), .ZN(new_n1063));
  AOI21_X1  g0863(.A(new_n1061), .B1(new_n1042), .B2(new_n1043), .ZN(new_n1064));
  OAI21_X1  g0864(.A(new_n1063), .B1(new_n1064), .B2(new_n806), .ZN(new_n1065));
  NAND4_X1  g0865(.A1(new_n371), .A2(new_n372), .A3(new_n454), .A4(new_n678), .ZN(new_n1066));
  INV_X1    g0866(.A(KEYINPUT113), .ZN(new_n1067));
  XNOR2_X1  g0867(.A(new_n1066), .B(new_n1067), .ZN(new_n1068));
  NAND3_X1  g0868(.A1(new_n880), .A2(new_n1065), .A3(new_n1068), .ZN(new_n1069));
  NAND2_X1  g0869(.A1(new_n1050), .A2(new_n1069), .ZN(new_n1070));
  AND3_X1   g0870(.A1(new_n880), .A2(new_n1065), .A3(new_n1068), .ZN(new_n1071));
  OAI211_X1 g0871(.A(new_n1071), .B(new_n1046), .C1(new_n1048), .C2(new_n1049), .ZN(new_n1072));
  NAND3_X1  g0872(.A1(new_n1070), .A2(new_n646), .A3(new_n1072), .ZN(new_n1073));
  AOI21_X1  g0873(.A(new_n685), .B1(new_n443), .B2(new_n768), .ZN(new_n1074));
  OAI22_X1  g0874(.A1(new_n327), .A2(new_n771), .B1(new_n712), .B2(new_n733), .ZN(new_n1075));
  AOI211_X1 g0875(.A(new_n1023), .B(new_n1075), .C1(G68), .C2(new_n773), .ZN(new_n1076));
  OAI221_X1 g0876(.A(new_n264), .B1(new_n702), .B2(new_n482), .C1(new_n225), .C2(new_n704), .ZN(new_n1077));
  NOR2_X1   g0877(.A1(new_n729), .A2(new_n523), .ZN(new_n1078));
  AOI211_X1 g0878(.A(new_n1077), .B(new_n1078), .C1(G116), .C2(new_n724), .ZN(new_n1079));
  INV_X1    g0879(.A(G132), .ZN(new_n1080));
  INV_X1    g0880(.A(G125), .ZN(new_n1081));
  OAI22_X1  g0881(.A1(new_n723), .A2(new_n1080), .B1(new_n729), .B2(new_n1081), .ZN(new_n1082));
  NAND2_X1  g0882(.A1(new_n994), .A2(G150), .ZN(new_n1083));
  XNOR2_X1  g0883(.A(new_n1083), .B(KEYINPUT53), .ZN(new_n1084));
  INV_X1    g0884(.A(G128), .ZN(new_n1085));
  OAI221_X1 g0885(.A(new_n273), .B1(new_n202), .B2(new_n706), .C1(new_n712), .C2(new_n1085), .ZN(new_n1086));
  NOR3_X1   g0886(.A1(new_n1082), .A2(new_n1084), .A3(new_n1086), .ZN(new_n1087));
  XOR2_X1   g0887(.A(KEYINPUT54), .B(G143), .Z(new_n1088));
  AOI22_X1  g0888(.A1(G159), .A2(new_n715), .B1(new_n785), .B2(new_n1088), .ZN(new_n1089));
  NAND2_X1  g0889(.A1(new_n709), .A2(new_n916), .ZN(new_n1090));
  NAND2_X1  g0890(.A1(new_n1089), .A2(new_n1090), .ZN(new_n1091));
  XNOR2_X1  g0891(.A(new_n1091), .B(KEYINPUT115), .ZN(new_n1092));
  AOI22_X1  g0892(.A1(new_n1076), .A2(new_n1079), .B1(new_n1087), .B2(new_n1092), .ZN(new_n1093));
  OAI21_X1  g0893(.A(new_n1074), .B1(new_n1093), .B2(new_n699), .ZN(new_n1094));
  NAND2_X1  g0894(.A1(new_n846), .A2(KEYINPUT39), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n1095), .A2(new_n867), .ZN(new_n1096));
  NAND3_X1  g0896(.A1(new_n846), .A2(KEYINPUT101), .A3(KEYINPUT39), .ZN(new_n1097));
  AOI22_X1  g0897(.A1(new_n1096), .A2(new_n1097), .B1(new_n863), .B2(new_n864), .ZN(new_n1098));
  AOI21_X1  g0898(.A(new_n1094), .B1(new_n1098), .B2(new_n693), .ZN(new_n1099));
  INV_X1    g0899(.A(new_n1099), .ZN(new_n1100));
  NAND3_X1  g0900(.A1(new_n1060), .A2(new_n1073), .A3(new_n1100), .ZN(G378));
  AOI21_X1  g0901(.A(new_n883), .B1(new_n841), .B2(new_n845), .ZN(new_n1102));
  OAI211_X1 g0902(.A(new_n889), .B(G330), .C1(new_n1102), .C2(KEYINPUT40), .ZN(new_n1103));
  XOR2_X1   g0903(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1104));
  NAND2_X1  g0904(.A1(new_n307), .A2(new_n820), .ZN(new_n1105));
  XOR2_X1   g0905(.A(new_n1105), .B(KEYINPUT116), .Z(new_n1106));
  INV_X1    g0906(.A(new_n1106), .ZN(new_n1107));
  NAND3_X1  g0907(.A1(new_n325), .A2(new_n368), .A3(new_n1107), .ZN(new_n1108));
  INV_X1    g0908(.A(new_n368), .ZN(new_n1109));
  OAI21_X1  g0909(.A(new_n1106), .B1(new_n622), .B2(new_n1109), .ZN(new_n1110));
  AOI21_X1  g0910(.A(new_n1104), .B1(new_n1108), .B2(new_n1110), .ZN(new_n1111));
  INV_X1    g0911(.A(new_n1111), .ZN(new_n1112));
  NAND3_X1  g0912(.A1(new_n1108), .A2(new_n1110), .A3(new_n1104), .ZN(new_n1113));
  NAND2_X1  g0913(.A1(new_n1112), .A2(new_n1113), .ZN(new_n1114));
  NAND2_X1  g0914(.A1(new_n1103), .A2(new_n1114), .ZN(new_n1115));
  NAND3_X1  g0915(.A1(new_n1112), .A2(KEYINPUT117), .A3(new_n1113), .ZN(new_n1116));
  INV_X1    g0916(.A(KEYINPUT117), .ZN(new_n1117));
  INV_X1    g0917(.A(new_n1113), .ZN(new_n1118));
  OAI21_X1  g0918(.A(new_n1117), .B1(new_n1118), .B2(new_n1111), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n1116), .A2(new_n1119), .ZN(new_n1120));
  NAND4_X1  g0920(.A1(new_n1120), .A2(G330), .A3(new_n887), .A4(new_n889), .ZN(new_n1121));
  NOR2_X1   g0921(.A1(new_n1098), .A2(new_n1032), .ZN(new_n1122));
  OAI211_X1 g0922(.A(new_n1115), .B(new_n1121), .C1(new_n1122), .C2(new_n855), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n1121), .A2(new_n1115), .ZN(new_n1124));
  NAND2_X1  g0924(.A1(new_n1124), .A2(new_n871), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n1123), .A2(new_n1125), .ZN(new_n1126));
  NAND2_X1  g0926(.A1(new_n1126), .A2(new_n683), .ZN(new_n1127));
  NAND2_X1  g0927(.A1(new_n1120), .A2(new_n693), .ZN(new_n1128));
  AOI21_X1  g0928(.A(new_n685), .B1(new_n202), .B2(new_n768), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n785), .A2(G137), .ZN(new_n1130));
  OAI21_X1  g0930(.A(new_n1130), .B1(new_n771), .B2(new_n1080), .ZN(new_n1131));
  AOI22_X1  g0931(.A1(new_n994), .A2(new_n1088), .B1(new_n715), .B2(G150), .ZN(new_n1132));
  OAI21_X1  g0932(.A(new_n1132), .B1(new_n1081), .B2(new_n712), .ZN(new_n1133));
  AOI211_X1 g0933(.A(new_n1131), .B(new_n1133), .C1(G128), .C2(new_n724), .ZN(new_n1134));
  INV_X1    g0934(.A(KEYINPUT59), .ZN(new_n1135));
  OR2_X1    g0935(.A1(new_n1134), .A2(new_n1135), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n1134), .A2(new_n1135), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n743), .A2(G124), .ZN(new_n1138));
  AOI211_X1 g0938(.A(G33), .B(G41), .C1(new_n784), .C2(new_n773), .ZN(new_n1139));
  NAND4_X1  g0939(.A1(new_n1136), .A2(new_n1137), .A3(new_n1138), .A4(new_n1139), .ZN(new_n1140));
  AOI22_X1  g0940(.A1(new_n724), .A2(G107), .B1(new_n743), .B2(G283), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n264), .A2(new_n458), .ZN(new_n1142));
  NOR2_X1   g0942(.A1(new_n925), .A2(new_n1142), .ZN(new_n1143));
  OAI211_X1 g0943(.A(new_n1141), .B(new_n1143), .C1(new_n563), .C2(new_n702), .ZN(new_n1144));
  NOR2_X1   g0944(.A1(new_n706), .A2(new_n283), .ZN(new_n1145));
  OAI22_X1  g0945(.A1(new_n482), .A2(new_n771), .B1(new_n712), .B2(new_n574), .ZN(new_n1146));
  NOR4_X1   g0946(.A1(new_n1144), .A2(new_n985), .A3(new_n1145), .A4(new_n1146), .ZN(new_n1147));
  OR2_X1    g0947(.A1(new_n1147), .A2(KEYINPUT58), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n1147), .A2(KEYINPUT58), .ZN(new_n1149));
  OAI211_X1 g0949(.A(new_n1142), .B(new_n202), .C1(G33), .C2(G41), .ZN(new_n1150));
  AND4_X1   g0950(.A1(new_n1140), .A2(new_n1148), .A3(new_n1149), .A4(new_n1150), .ZN(new_n1151));
  OAI211_X1 g0951(.A(new_n1128), .B(new_n1129), .C1(new_n699), .C2(new_n1151), .ZN(new_n1152));
  AND2_X1   g0952(.A1(new_n1127), .A2(new_n1152), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n880), .A2(new_n1068), .ZN(new_n1154));
  AOI21_X1  g0954(.A(new_n1154), .B1(new_n1057), .B2(new_n1071), .ZN(new_n1155));
  AND2_X1   g0955(.A1(new_n1124), .A2(new_n871), .ZN(new_n1156));
  NOR2_X1   g0956(.A1(new_n1124), .A2(new_n871), .ZN(new_n1157));
  OAI21_X1  g0957(.A(KEYINPUT57), .B1(new_n1156), .B2(new_n1157), .ZN(new_n1158));
  OAI21_X1  g0958(.A(new_n646), .B1(new_n1155), .B2(new_n1158), .ZN(new_n1159));
  INV_X1    g0959(.A(new_n1154), .ZN(new_n1160));
  NAND2_X1  g0960(.A1(new_n1072), .A2(new_n1160), .ZN(new_n1161));
  AOI21_X1  g0961(.A(KEYINPUT57), .B1(new_n1161), .B2(new_n1126), .ZN(new_n1162));
  OAI21_X1  g0962(.A(new_n1153), .B1(new_n1159), .B2(new_n1162), .ZN(G375));
  OAI221_X1 g0963(.A(new_n273), .B1(new_n702), .B2(new_n787), .C1(new_n283), .C2(new_n706), .ZN(new_n1164));
  AOI22_X1  g0964(.A1(G132), .A2(new_n711), .B1(new_n709), .B2(new_n1088), .ZN(new_n1165));
  OAI21_X1  g0965(.A(new_n1165), .B1(new_n202), .B2(new_n716), .ZN(new_n1166));
  AOI211_X1 g0966(.A(new_n1164), .B(new_n1166), .C1(new_n724), .C2(new_n916), .ZN(new_n1167));
  OAI22_X1  g0967(.A1(new_n729), .A2(new_n1085), .B1(new_n983), .B2(new_n704), .ZN(new_n1168));
  XOR2_X1   g0968(.A(new_n1168), .B(KEYINPUT118), .Z(new_n1169));
  AOI22_X1  g0969(.A1(new_n724), .A2(G283), .B1(new_n743), .B2(G303), .ZN(new_n1170));
  AOI211_X1 g0970(.A(new_n273), .B(new_n922), .C1(G107), .C2(new_n785), .ZN(new_n1171));
  AND3_X1   g0971(.A1(new_n1170), .A2(new_n1171), .A3(new_n980), .ZN(new_n1172));
  OAI22_X1  g0972(.A1(new_n771), .A2(new_n574), .B1(new_n704), .B2(new_n482), .ZN(new_n1173));
  AOI21_X1  g0973(.A(new_n1173), .B1(G294), .B2(new_n711), .ZN(new_n1174));
  AOI22_X1  g0974(.A1(new_n1167), .A2(new_n1169), .B1(new_n1172), .B2(new_n1174), .ZN(new_n1175));
  OAI221_X1 g0975(.A(new_n684), .B1(G68), .B2(new_n769), .C1(new_n1175), .C2(new_n699), .ZN(new_n1176));
  AOI21_X1  g0976(.A(new_n1176), .B1(new_n1033), .B2(new_n693), .ZN(new_n1177));
  AOI21_X1  g0977(.A(new_n1177), .B1(new_n1065), .B2(new_n683), .ZN(new_n1178));
  NAND2_X1  g0978(.A1(new_n1069), .A2(new_n951), .ZN(new_n1179));
  AOI21_X1  g0979(.A(new_n1065), .B1(new_n880), .B2(new_n1068), .ZN(new_n1180));
  OAI21_X1  g0980(.A(new_n1178), .B1(new_n1179), .B2(new_n1180), .ZN(G381));
  INV_X1    g0981(.A(G390), .ZN(new_n1182));
  INV_X1    g0982(.A(G384), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n1182), .A2(new_n1183), .ZN(new_n1184));
  OR4_X1    g0984(.A1(G396), .A2(new_n1184), .A3(G387), .A4(G393), .ZN(new_n1185));
  OR4_X1    g0985(.A1(G378), .A2(new_n1185), .A3(G375), .A4(G381), .ZN(G407));
  AND3_X1   g0986(.A1(new_n1060), .A2(new_n1073), .A3(new_n1100), .ZN(new_n1187));
  NAND2_X1  g0987(.A1(new_n629), .A2(G213), .ZN(new_n1188));
  INV_X1    g0988(.A(new_n1188), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n1187), .A2(new_n1189), .ZN(new_n1190));
  OAI211_X1 g0990(.A(G407), .B(G213), .C1(G375), .C2(new_n1190), .ZN(G409));
  NAND2_X1  g0991(.A1(G387), .A2(new_n1182), .ZN(new_n1192));
  OAI211_X1 g0992(.A(G390), .B(new_n930), .C1(new_n952), .C2(new_n963), .ZN(new_n1193));
  NAND2_X1  g0993(.A1(new_n1192), .A2(new_n1193), .ZN(new_n1194));
  XOR2_X1   g0994(.A(G393), .B(G396), .Z(new_n1195));
  INV_X1    g0995(.A(new_n1195), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(new_n1194), .A2(new_n1196), .ZN(new_n1197));
  NAND3_X1  g0997(.A1(new_n1192), .A2(new_n1195), .A3(new_n1193), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(new_n1197), .A2(new_n1198), .ZN(new_n1199));
  INV_X1    g0999(.A(KEYINPUT124), .ZN(new_n1200));
  XNOR2_X1  g1000(.A(new_n1199), .B(new_n1200), .ZN(new_n1201));
  AOI21_X1  g1001(.A(new_n647), .B1(new_n1050), .B2(new_n1069), .ZN(new_n1202));
  AOI21_X1  g1002(.A(new_n1099), .B1(new_n1202), .B2(new_n1072), .ZN(new_n1203));
  AOI221_X4 g1003(.A(new_n950), .B1(new_n1123), .B2(new_n1125), .C1(new_n1072), .C2(new_n1160), .ZN(new_n1204));
  NAND2_X1  g1004(.A1(new_n1127), .A2(new_n1152), .ZN(new_n1205));
  OAI211_X1 g1005(.A(new_n1203), .B(new_n1060), .C1(new_n1204), .C2(new_n1205), .ZN(new_n1206));
  OAI21_X1  g1006(.A(new_n1206), .B1(G375), .B2(new_n1187), .ZN(new_n1207));
  INV_X1    g1007(.A(KEYINPUT62), .ZN(new_n1208));
  INV_X1    g1008(.A(new_n1065), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(new_n1154), .A2(new_n1209), .ZN(new_n1210));
  INV_X1    g1010(.A(KEYINPUT60), .ZN(new_n1211));
  OAI21_X1  g1011(.A(new_n1210), .B1(new_n1071), .B2(new_n1211), .ZN(new_n1212));
  NAND3_X1  g1012(.A1(new_n1154), .A2(new_n1209), .A3(KEYINPUT60), .ZN(new_n1213));
  NAND3_X1  g1013(.A1(new_n1212), .A2(new_n646), .A3(new_n1213), .ZN(new_n1214));
  AOI21_X1  g1014(.A(G384), .B1(new_n1214), .B2(new_n1178), .ZN(new_n1215));
  AOI21_X1  g1015(.A(new_n1180), .B1(KEYINPUT60), .B2(new_n1069), .ZN(new_n1216));
  NAND2_X1  g1016(.A1(new_n1213), .A2(new_n646), .ZN(new_n1217));
  OAI211_X1 g1017(.A(G384), .B(new_n1178), .C1(new_n1216), .C2(new_n1217), .ZN(new_n1218));
  INV_X1    g1018(.A(new_n1218), .ZN(new_n1219));
  NOR2_X1   g1019(.A1(new_n1215), .A2(new_n1219), .ZN(new_n1220));
  NAND4_X1  g1020(.A1(new_n1207), .A2(new_n1208), .A3(new_n1188), .A4(new_n1220), .ZN(new_n1221));
  INV_X1    g1021(.A(KEYINPUT61), .ZN(new_n1222));
  INV_X1    g1022(.A(KEYINPUT57), .ZN(new_n1223));
  AOI21_X1  g1023(.A(new_n1223), .B1(new_n1123), .B2(new_n1125), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(new_n1161), .A2(new_n1224), .ZN(new_n1225));
  AOI22_X1  g1025(.A1(new_n1072), .A2(new_n1160), .B1(new_n1125), .B2(new_n1123), .ZN(new_n1226));
  OAI211_X1 g1026(.A(new_n1225), .B(new_n646), .C1(KEYINPUT57), .C2(new_n1226), .ZN(new_n1227));
  NAND3_X1  g1027(.A1(new_n1227), .A2(G378), .A3(new_n1153), .ZN(new_n1228));
  AOI21_X1  g1028(.A(new_n1189), .B1(new_n1228), .B2(new_n1206), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n1214), .A2(new_n1178), .ZN(new_n1230));
  NAND2_X1  g1030(.A1(new_n1230), .A2(new_n1183), .ZN(new_n1231));
  NAND2_X1  g1031(.A1(new_n1189), .A2(G2897), .ZN(new_n1232));
  XOR2_X1   g1032(.A(new_n1232), .B(KEYINPUT121), .Z(new_n1233));
  INV_X1    g1033(.A(new_n1233), .ZN(new_n1234));
  NAND3_X1  g1034(.A1(new_n1231), .A2(new_n1218), .A3(new_n1234), .ZN(new_n1235));
  OAI21_X1  g1035(.A(new_n1233), .B1(new_n1215), .B2(new_n1219), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n1235), .A2(new_n1236), .ZN(new_n1237));
  OAI211_X1 g1037(.A(new_n1221), .B(new_n1222), .C1(new_n1229), .C2(new_n1237), .ZN(new_n1238));
  AOI21_X1  g1038(.A(new_n1208), .B1(new_n1229), .B2(new_n1220), .ZN(new_n1239));
  OAI21_X1  g1039(.A(new_n1201), .B1(new_n1238), .B2(new_n1239), .ZN(new_n1240));
  NAND3_X1  g1040(.A1(new_n1197), .A2(new_n1222), .A3(new_n1198), .ZN(new_n1241));
  AOI21_X1  g1041(.A(new_n1237), .B1(new_n1207), .B2(new_n1188), .ZN(new_n1242));
  INV_X1    g1042(.A(KEYINPUT122), .ZN(new_n1243));
  AOI21_X1  g1043(.A(new_n1241), .B1(new_n1242), .B2(new_n1243), .ZN(new_n1244));
  OAI21_X1  g1044(.A(KEYINPUT122), .B1(new_n1229), .B2(new_n1237), .ZN(new_n1245));
  NAND4_X1  g1045(.A1(new_n1207), .A2(KEYINPUT63), .A3(new_n1188), .A4(new_n1220), .ZN(new_n1246));
  INV_X1    g1046(.A(KEYINPUT123), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n1246), .A2(new_n1247), .ZN(new_n1248));
  NAND4_X1  g1048(.A1(new_n1229), .A2(KEYINPUT123), .A3(KEYINPUT63), .A4(new_n1220), .ZN(new_n1249));
  NAND4_X1  g1049(.A1(new_n1244), .A2(new_n1245), .A3(new_n1248), .A4(new_n1249), .ZN(new_n1250));
  INV_X1    g1050(.A(KEYINPUT120), .ZN(new_n1251));
  XOR2_X1   g1051(.A(KEYINPUT119), .B(KEYINPUT63), .Z(new_n1252));
  AOI211_X1 g1052(.A(new_n1251), .B(new_n1252), .C1(new_n1229), .C2(new_n1220), .ZN(new_n1253));
  NAND3_X1  g1053(.A1(new_n1207), .A2(new_n1188), .A3(new_n1220), .ZN(new_n1254));
  INV_X1    g1054(.A(new_n1252), .ZN(new_n1255));
  AOI21_X1  g1055(.A(KEYINPUT120), .B1(new_n1254), .B2(new_n1255), .ZN(new_n1256));
  NOR2_X1   g1056(.A1(new_n1253), .A2(new_n1256), .ZN(new_n1257));
  OAI21_X1  g1057(.A(new_n1240), .B1(new_n1250), .B2(new_n1257), .ZN(new_n1258));
  INV_X1    g1058(.A(KEYINPUT125), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(new_n1258), .A2(new_n1259), .ZN(new_n1260));
  OAI211_X1 g1060(.A(new_n1240), .B(KEYINPUT125), .C1(new_n1250), .C2(new_n1257), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(new_n1260), .A2(new_n1261), .ZN(G405));
  NAND2_X1  g1062(.A1(G375), .A2(new_n1187), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n1263), .A2(new_n1228), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(new_n1220), .A2(KEYINPUT126), .ZN(new_n1265));
  XNOR2_X1  g1065(.A(new_n1264), .B(new_n1265), .ZN(new_n1266));
  INV_X1    g1066(.A(KEYINPUT127), .ZN(new_n1267));
  AOI21_X1  g1067(.A(new_n1266), .B1(new_n1267), .B2(new_n1199), .ZN(new_n1268));
  INV_X1    g1068(.A(new_n1199), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n1269), .A2(KEYINPUT127), .ZN(new_n1270));
  XNOR2_X1  g1070(.A(new_n1268), .B(new_n1270), .ZN(G402));
endmodule


