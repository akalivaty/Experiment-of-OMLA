//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 1 0 0 0 1 0 1 1 0 0 0 1 0 0 1 1 1 1 0 0 0 0 0 0 0 0 1 0 1 0 0 1 0 0 0 0 1 0 1 0 0 1 1 0 1 0 1 0 1 1 0 1 1 0 1 1 0 0 0 1 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:40:28 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1113, new_n1114, new_n1115, new_n1116, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1190, new_n1191,
    new_n1192, new_n1193, new_n1194, new_n1195, new_n1196, new_n1197,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1255, new_n1256, new_n1257, new_n1258,
    new_n1259, new_n1260, new_n1261, new_n1262, new_n1263, new_n1264,
    new_n1265, new_n1266, new_n1267, new_n1268, new_n1270, new_n1271,
    new_n1272, new_n1273, new_n1274, new_n1275, new_n1276, new_n1277,
    new_n1278, new_n1279, new_n1280, new_n1281, new_n1282, new_n1283,
    new_n1284, new_n1285, new_n1286, new_n1287, new_n1288, new_n1289,
    new_n1291, new_n1292, new_n1294, new_n1295, new_n1296, new_n1297,
    new_n1298, new_n1299, new_n1300, new_n1301, new_n1302, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1350, new_n1351, new_n1352,
    new_n1353, new_n1354, new_n1355, new_n1357, new_n1358, new_n1359,
    new_n1360, new_n1361, new_n1362, new_n1363;
  XNOR2_X1  g0000(.A(KEYINPUT64), .B(G50), .ZN(new_n201));
  INV_X1    g0001(.A(new_n201), .ZN(new_n202));
  NOR2_X1   g0002(.A1(G58), .A2(G68), .ZN(new_n203));
  INV_X1    g0003(.A(new_n203), .ZN(new_n204));
  NOR3_X1   g0004(.A1(new_n202), .A2(G77), .A3(new_n204), .ZN(G353));
  OAI21_X1  g0005(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0006(.A(G1), .ZN(new_n207));
  INV_X1    g0007(.A(G20), .ZN(new_n208));
  NOR2_X1   g0008(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  INV_X1    g0009(.A(new_n209), .ZN(new_n210));
  NOR2_X1   g0010(.A1(new_n210), .A2(G13), .ZN(new_n211));
  OAI211_X1 g0011(.A(new_n211), .B(G250), .C1(G257), .C2(G264), .ZN(new_n212));
  XNOR2_X1  g0012(.A(new_n212), .B(KEYINPUT0), .ZN(new_n213));
  NAND2_X1  g0013(.A1(G1), .A2(G13), .ZN(new_n214));
  NOR2_X1   g0014(.A1(new_n214), .A2(new_n208), .ZN(new_n215));
  INV_X1    g0015(.A(new_n215), .ZN(new_n216));
  NAND2_X1  g0016(.A1(new_n204), .A2(G50), .ZN(new_n217));
  AOI22_X1  g0017(.A1(G107), .A2(G264), .B1(G116), .B2(G270), .ZN(new_n218));
  INV_X1    g0018(.A(G77), .ZN(new_n219));
  INV_X1    g0019(.A(G244), .ZN(new_n220));
  INV_X1    g0020(.A(G87), .ZN(new_n221));
  INV_X1    g0021(.A(G250), .ZN(new_n222));
  OAI221_X1 g0022(.A(new_n218), .B1(new_n219), .B2(new_n220), .C1(new_n221), .C2(new_n222), .ZN(new_n223));
  AOI22_X1  g0023(.A1(G50), .A2(G226), .B1(G97), .B2(G257), .ZN(new_n224));
  INV_X1    g0024(.A(G58), .ZN(new_n225));
  INV_X1    g0025(.A(G232), .ZN(new_n226));
  INV_X1    g0026(.A(G68), .ZN(new_n227));
  INV_X1    g0027(.A(G238), .ZN(new_n228));
  OAI221_X1 g0028(.A(new_n224), .B1(new_n225), .B2(new_n226), .C1(new_n227), .C2(new_n228), .ZN(new_n229));
  OAI21_X1  g0029(.A(new_n210), .B1(new_n223), .B2(new_n229), .ZN(new_n230));
  OAI221_X1 g0030(.A(new_n213), .B1(new_n216), .B2(new_n217), .C1(KEYINPUT1), .C2(new_n230), .ZN(new_n231));
  NAND2_X1  g0031(.A1(new_n230), .A2(KEYINPUT1), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n232), .B(KEYINPUT65), .ZN(new_n233));
  NOR2_X1   g0033(.A1(new_n231), .A2(new_n233), .ZN(G361));
  XNOR2_X1  g0034(.A(G238), .B(G244), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n235), .B(KEYINPUT2), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n236), .B(G226), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n237), .B(new_n226), .ZN(new_n238));
  XNOR2_X1  g0038(.A(G250), .B(G257), .ZN(new_n239));
  XNOR2_X1  g0039(.A(G264), .B(G270), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n238), .B(new_n241), .ZN(G358));
  XOR2_X1   g0042(.A(G50), .B(G58), .Z(new_n243));
  XNOR2_X1  g0043(.A(new_n243), .B(KEYINPUT66), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n244), .B(KEYINPUT67), .ZN(new_n245));
  XOR2_X1   g0045(.A(G68), .B(G77), .Z(new_n246));
  XNOR2_X1  g0046(.A(new_n245), .B(new_n246), .ZN(new_n247));
  XNOR2_X1  g0047(.A(G87), .B(G97), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n248), .B(KEYINPUT68), .ZN(new_n249));
  XNOR2_X1  g0049(.A(G107), .B(G116), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n249), .B(new_n250), .ZN(new_n251));
  XNOR2_X1  g0051(.A(new_n247), .B(new_n251), .ZN(G351));
  AND2_X1   g0052(.A1(KEYINPUT3), .A2(G33), .ZN(new_n253));
  NOR2_X1   g0053(.A1(KEYINPUT3), .A2(G33), .ZN(new_n254));
  OAI211_X1 g0054(.A(G232), .B(G1698), .C1(new_n253), .C2(new_n254), .ZN(new_n255));
  INV_X1    g0055(.A(G1698), .ZN(new_n256));
  OAI211_X1 g0056(.A(G226), .B(new_n256), .C1(new_n253), .C2(new_n254), .ZN(new_n257));
  INV_X1    g0057(.A(G33), .ZN(new_n258));
  INV_X1    g0058(.A(G97), .ZN(new_n259));
  OAI211_X1 g0059(.A(new_n255), .B(new_n257), .C1(new_n258), .C2(new_n259), .ZN(new_n260));
  AOI21_X1  g0060(.A(new_n214), .B1(G33), .B2(G41), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  INV_X1    g0062(.A(new_n214), .ZN(new_n263));
  NAND2_X1  g0063(.A1(G33), .A2(G41), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  OAI21_X1  g0065(.A(new_n207), .B1(G41), .B2(G45), .ZN(new_n266));
  AND2_X1   g0066(.A1(new_n265), .A2(new_n266), .ZN(new_n267));
  INV_X1    g0067(.A(G45), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n268), .A2(KEYINPUT69), .ZN(new_n269));
  INV_X1    g0069(.A(KEYINPUT69), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n270), .A2(G45), .ZN(new_n271));
  INV_X1    g0071(.A(G41), .ZN(new_n272));
  NAND3_X1  g0072(.A1(new_n269), .A2(new_n271), .A3(new_n272), .ZN(new_n273));
  INV_X1    g0073(.A(G274), .ZN(new_n274));
  NOR2_X1   g0074(.A1(new_n274), .A2(G1), .ZN(new_n275));
  AOI22_X1  g0075(.A1(new_n267), .A2(G238), .B1(new_n273), .B2(new_n275), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n262), .A2(new_n276), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n277), .A2(KEYINPUT13), .ZN(new_n278));
  INV_X1    g0078(.A(KEYINPUT13), .ZN(new_n279));
  NAND3_X1  g0079(.A1(new_n262), .A2(new_n276), .A3(new_n279), .ZN(new_n280));
  NAND3_X1  g0080(.A1(new_n278), .A2(KEYINPUT72), .A3(new_n280), .ZN(new_n281));
  OR3_X1    g0081(.A1(new_n277), .A2(KEYINPUT72), .A3(KEYINPUT13), .ZN(new_n282));
  NAND3_X1  g0082(.A1(new_n281), .A2(new_n282), .A3(G169), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n283), .A2(KEYINPUT14), .ZN(new_n284));
  INV_X1    g0084(.A(KEYINPUT14), .ZN(new_n285));
  NAND4_X1  g0085(.A1(new_n281), .A2(new_n282), .A3(new_n285), .A4(G169), .ZN(new_n286));
  NAND3_X1  g0086(.A1(new_n278), .A2(G179), .A3(new_n280), .ZN(new_n287));
  NAND3_X1  g0087(.A1(new_n284), .A2(new_n286), .A3(new_n287), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n227), .A2(G20), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n208), .A2(G33), .ZN(new_n290));
  NOR2_X1   g0090(.A1(G20), .A2(G33), .ZN(new_n291));
  INV_X1    g0091(.A(new_n291), .ZN(new_n292));
  INV_X1    g0092(.A(G50), .ZN(new_n293));
  OAI221_X1 g0093(.A(new_n289), .B1(new_n290), .B2(new_n219), .C1(new_n292), .C2(new_n293), .ZN(new_n294));
  NAND3_X1  g0094(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n295), .A2(new_n214), .ZN(new_n296));
  AND2_X1   g0096(.A1(new_n294), .A2(new_n296), .ZN(new_n297));
  OR2_X1    g0097(.A1(new_n297), .A2(KEYINPUT11), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n297), .A2(KEYINPUT11), .ZN(new_n299));
  INV_X1    g0099(.A(KEYINPUT12), .ZN(new_n300));
  INV_X1    g0100(.A(G13), .ZN(new_n301));
  NOR3_X1   g0101(.A1(new_n300), .A2(new_n301), .A3(G1), .ZN(new_n302));
  INV_X1    g0102(.A(new_n289), .ZN(new_n303));
  NAND3_X1  g0103(.A1(new_n207), .A2(G13), .A3(G20), .ZN(new_n304));
  AOI22_X1  g0104(.A1(new_n302), .A2(new_n303), .B1(new_n300), .B2(new_n304), .ZN(new_n305));
  OAI211_X1 g0105(.A(new_n295), .B(new_n214), .C1(G1), .C2(new_n208), .ZN(new_n306));
  INV_X1    g0106(.A(new_n306), .ZN(new_n307));
  OAI21_X1  g0107(.A(G68), .B1(new_n307), .B2(new_n300), .ZN(new_n308));
  NAND4_X1  g0108(.A1(new_n298), .A2(new_n299), .A3(new_n305), .A4(new_n308), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n288), .A2(new_n309), .ZN(new_n310));
  AND2_X1   g0110(.A1(new_n280), .A2(G190), .ZN(new_n311));
  AOI21_X1  g0111(.A(new_n309), .B1(new_n311), .B2(new_n278), .ZN(new_n312));
  NAND3_X1  g0112(.A1(new_n281), .A2(new_n282), .A3(G200), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n310), .A2(new_n314), .ZN(new_n315));
  XNOR2_X1  g0115(.A(KEYINPUT8), .B(G58), .ZN(new_n316));
  INV_X1    g0116(.A(G150), .ZN(new_n317));
  OAI22_X1  g0117(.A1(new_n316), .A2(new_n290), .B1(new_n317), .B2(new_n292), .ZN(new_n318));
  AOI21_X1  g0118(.A(new_n208), .B1(new_n201), .B2(new_n203), .ZN(new_n319));
  OAI21_X1  g0119(.A(new_n296), .B1(new_n318), .B2(new_n319), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n307), .A2(G50), .ZN(new_n321));
  OAI211_X1 g0121(.A(new_n320), .B(new_n321), .C1(G50), .C2(new_n304), .ZN(new_n322));
  XNOR2_X1  g0122(.A(new_n322), .B(KEYINPUT9), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n267), .A2(G226), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n273), .A2(new_n275), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n324), .A2(new_n325), .ZN(new_n326));
  INV_X1    g0126(.A(new_n326), .ZN(new_n327));
  INV_X1    g0127(.A(KEYINPUT3), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n328), .A2(new_n258), .ZN(new_n329));
  NAND2_X1  g0129(.A1(KEYINPUT3), .A2(G33), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  NAND3_X1  g0131(.A1(new_n331), .A2(G222), .A3(new_n256), .ZN(new_n332));
  XNOR2_X1  g0132(.A(new_n332), .B(KEYINPUT70), .ZN(new_n333));
  NOR2_X1   g0133(.A1(new_n253), .A2(new_n254), .ZN(new_n334));
  NOR2_X1   g0134(.A1(new_n334), .A2(new_n256), .ZN(new_n335));
  AOI22_X1  g0135(.A1(new_n335), .A2(G223), .B1(G77), .B2(new_n334), .ZN(new_n336));
  AND2_X1   g0136(.A1(new_n333), .A2(new_n336), .ZN(new_n337));
  OAI211_X1 g0137(.A(G190), .B(new_n327), .C1(new_n337), .C2(new_n265), .ZN(new_n338));
  AOI21_X1  g0138(.A(new_n265), .B1(new_n333), .B2(new_n336), .ZN(new_n339));
  OAI21_X1  g0139(.A(G200), .B1(new_n339), .B2(new_n326), .ZN(new_n340));
  NAND3_X1  g0140(.A1(new_n323), .A2(new_n338), .A3(new_n340), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n341), .A2(KEYINPUT10), .ZN(new_n342));
  INV_X1    g0142(.A(KEYINPUT10), .ZN(new_n343));
  NAND4_X1  g0143(.A1(new_n323), .A2(new_n338), .A3(new_n343), .A4(new_n340), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n342), .A2(new_n344), .ZN(new_n345));
  OAI21_X1  g0145(.A(new_n327), .B1(new_n337), .B2(new_n265), .ZN(new_n346));
  OR2_X1    g0146(.A1(new_n346), .A2(G179), .ZN(new_n347));
  INV_X1    g0147(.A(G169), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n346), .A2(new_n348), .ZN(new_n349));
  NAND3_X1  g0149(.A1(new_n347), .A2(new_n349), .A3(new_n322), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n345), .A2(new_n350), .ZN(new_n351));
  INV_X1    g0151(.A(G223), .ZN(new_n352));
  NOR2_X1   g0152(.A1(new_n352), .A2(G1698), .ZN(new_n353));
  OAI21_X1  g0153(.A(new_n353), .B1(new_n253), .B2(new_n254), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n354), .A2(KEYINPUT74), .ZN(new_n355));
  NAND2_X1  g0155(.A1(G33), .A2(G87), .ZN(new_n356));
  OAI211_X1 g0156(.A(G226), .B(G1698), .C1(new_n253), .C2(new_n254), .ZN(new_n357));
  INV_X1    g0157(.A(KEYINPUT74), .ZN(new_n358));
  OAI211_X1 g0158(.A(new_n353), .B(new_n358), .C1(new_n254), .C2(new_n253), .ZN(new_n359));
  NAND4_X1  g0159(.A1(new_n355), .A2(new_n356), .A3(new_n357), .A4(new_n359), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n360), .A2(new_n261), .ZN(new_n361));
  NAND3_X1  g0161(.A1(new_n265), .A2(G232), .A3(new_n266), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n325), .A2(new_n362), .ZN(new_n363));
  INV_X1    g0163(.A(new_n363), .ZN(new_n364));
  AOI21_X1  g0164(.A(G169), .B1(new_n361), .B2(new_n364), .ZN(new_n365));
  AOI211_X1 g0165(.A(G179), .B(new_n363), .C1(new_n360), .C2(new_n261), .ZN(new_n366));
  NOR2_X1   g0166(.A1(new_n365), .A2(new_n366), .ZN(new_n367));
  INV_X1    g0167(.A(KEYINPUT16), .ZN(new_n368));
  NAND3_X1  g0168(.A1(new_n329), .A2(new_n208), .A3(new_n330), .ZN(new_n369));
  INV_X1    g0169(.A(KEYINPUT7), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n369), .A2(new_n370), .ZN(new_n371));
  NAND4_X1  g0171(.A1(new_n329), .A2(KEYINPUT7), .A3(new_n208), .A4(new_n330), .ZN(new_n372));
  AOI21_X1  g0172(.A(new_n227), .B1(new_n371), .B2(new_n372), .ZN(new_n373));
  NOR2_X1   g0173(.A1(new_n225), .A2(new_n227), .ZN(new_n374));
  OAI21_X1  g0174(.A(G20), .B1(new_n374), .B2(new_n203), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n291), .A2(G159), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n375), .A2(new_n376), .ZN(new_n377));
  OAI21_X1  g0177(.A(new_n368), .B1(new_n373), .B2(new_n377), .ZN(new_n378));
  AOI21_X1  g0178(.A(KEYINPUT7), .B1(new_n334), .B2(new_n208), .ZN(new_n379));
  INV_X1    g0179(.A(new_n372), .ZN(new_n380));
  OAI21_X1  g0180(.A(G68), .B1(new_n379), .B2(new_n380), .ZN(new_n381));
  INV_X1    g0181(.A(new_n377), .ZN(new_n382));
  NAND3_X1  g0182(.A1(new_n381), .A2(KEYINPUT16), .A3(new_n382), .ZN(new_n383));
  NAND3_X1  g0183(.A1(new_n378), .A2(new_n383), .A3(new_n296), .ZN(new_n384));
  XOR2_X1   g0184(.A(KEYINPUT8), .B(G58), .Z(new_n385));
  NAND2_X1  g0185(.A1(new_n385), .A2(new_n306), .ZN(new_n386));
  INV_X1    g0186(.A(KEYINPUT73), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n316), .A2(new_n304), .ZN(new_n388));
  AND3_X1   g0188(.A1(new_n386), .A2(new_n387), .A3(new_n388), .ZN(new_n389));
  AOI21_X1  g0189(.A(new_n387), .B1(new_n386), .B2(new_n388), .ZN(new_n390));
  NOR2_X1   g0190(.A1(new_n389), .A2(new_n390), .ZN(new_n391));
  INV_X1    g0191(.A(new_n391), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n384), .A2(new_n392), .ZN(new_n393));
  INV_X1    g0193(.A(KEYINPUT18), .ZN(new_n394));
  AND3_X1   g0194(.A1(new_n367), .A2(new_n393), .A3(new_n394), .ZN(new_n395));
  AOI21_X1  g0195(.A(new_n394), .B1(new_n367), .B2(new_n393), .ZN(new_n396));
  NOR2_X1   g0196(.A1(new_n395), .A2(new_n396), .ZN(new_n397));
  AOI21_X1  g0197(.A(new_n363), .B1(new_n360), .B2(new_n261), .ZN(new_n398));
  INV_X1    g0198(.A(G200), .ZN(new_n399));
  OR2_X1    g0199(.A1(new_n398), .A2(new_n399), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n398), .A2(G190), .ZN(new_n401));
  NAND4_X1  g0201(.A1(new_n400), .A2(new_n384), .A3(new_n392), .A4(new_n401), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n402), .A2(KEYINPUT17), .ZN(new_n403));
  INV_X1    g0203(.A(new_n296), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n381), .A2(new_n382), .ZN(new_n405));
  AOI21_X1  g0205(.A(new_n404), .B1(new_n405), .B2(new_n368), .ZN(new_n406));
  AOI21_X1  g0206(.A(new_n391), .B1(new_n406), .B2(new_n383), .ZN(new_n407));
  INV_X1    g0207(.A(KEYINPUT17), .ZN(new_n408));
  NAND4_X1  g0208(.A1(new_n407), .A2(new_n408), .A3(new_n400), .A4(new_n401), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n403), .A2(new_n409), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n397), .A2(new_n410), .ZN(new_n411));
  OAI211_X1 g0211(.A(G232), .B(new_n256), .C1(new_n253), .C2(new_n254), .ZN(new_n412));
  OAI211_X1 g0212(.A(G238), .B(G1698), .C1(new_n253), .C2(new_n254), .ZN(new_n413));
  INV_X1    g0213(.A(G107), .ZN(new_n414));
  OAI211_X1 g0214(.A(new_n412), .B(new_n413), .C1(new_n414), .C2(new_n331), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n415), .A2(new_n261), .ZN(new_n416));
  AOI22_X1  g0216(.A1(new_n267), .A2(G244), .B1(new_n273), .B2(new_n275), .ZN(new_n417));
  INV_X1    g0217(.A(KEYINPUT71), .ZN(new_n418));
  NAND3_X1  g0218(.A1(new_n416), .A2(new_n417), .A3(new_n418), .ZN(new_n419));
  INV_X1    g0219(.A(new_n419), .ZN(new_n420));
  AOI21_X1  g0220(.A(new_n418), .B1(new_n416), .B2(new_n417), .ZN(new_n421));
  NOR2_X1   g0221(.A1(new_n420), .A2(new_n421), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n422), .A2(G200), .ZN(new_n423));
  XOR2_X1   g0223(.A(KEYINPUT15), .B(G87), .Z(new_n424));
  INV_X1    g0224(.A(new_n290), .ZN(new_n425));
  AOI22_X1  g0225(.A1(new_n424), .A2(new_n425), .B1(G20), .B2(G77), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n385), .A2(new_n291), .ZN(new_n427));
  AOI21_X1  g0227(.A(new_n404), .B1(new_n426), .B2(new_n427), .ZN(new_n428));
  INV_X1    g0228(.A(new_n304), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n429), .A2(new_n219), .ZN(new_n430));
  OAI21_X1  g0230(.A(new_n430), .B1(new_n219), .B2(new_n306), .ZN(new_n431));
  NOR2_X1   g0231(.A1(new_n428), .A2(new_n431), .ZN(new_n432));
  INV_X1    g0232(.A(G190), .ZN(new_n433));
  OAI211_X1 g0233(.A(new_n423), .B(new_n432), .C1(new_n433), .C2(new_n422), .ZN(new_n434));
  INV_X1    g0234(.A(new_n421), .ZN(new_n435));
  NAND3_X1  g0235(.A1(new_n435), .A2(new_n348), .A3(new_n419), .ZN(new_n436));
  INV_X1    g0236(.A(G179), .ZN(new_n437));
  OAI21_X1  g0237(.A(new_n437), .B1(new_n420), .B2(new_n421), .ZN(new_n438));
  INV_X1    g0238(.A(new_n432), .ZN(new_n439));
  NAND3_X1  g0239(.A1(new_n436), .A2(new_n438), .A3(new_n439), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n434), .A2(new_n440), .ZN(new_n441));
  NOR4_X1   g0241(.A1(new_n315), .A2(new_n351), .A3(new_n411), .A4(new_n441), .ZN(new_n442));
  INV_X1    g0242(.A(KEYINPUT4), .ZN(new_n443));
  NOR2_X1   g0243(.A1(new_n443), .A2(G1698), .ZN(new_n444));
  OAI211_X1 g0244(.A(new_n444), .B(G244), .C1(new_n254), .C2(new_n253), .ZN(new_n445));
  NAND2_X1  g0245(.A1(G33), .A2(G283), .ZN(new_n446));
  AOI21_X1  g0246(.A(new_n220), .B1(new_n329), .B2(new_n330), .ZN(new_n447));
  OAI211_X1 g0247(.A(new_n445), .B(new_n446), .C1(new_n447), .C2(KEYINPUT4), .ZN(new_n448));
  OAI21_X1  g0248(.A(G250), .B1(new_n253), .B2(new_n254), .ZN(new_n449));
  AOI21_X1  g0249(.A(new_n256), .B1(new_n449), .B2(KEYINPUT4), .ZN(new_n450));
  OAI21_X1  g0250(.A(new_n261), .B1(new_n448), .B2(new_n450), .ZN(new_n451));
  XNOR2_X1  g0251(.A(KEYINPUT5), .B(G41), .ZN(new_n452));
  NOR3_X1   g0252(.A1(new_n268), .A2(new_n274), .A3(G1), .ZN(new_n453));
  NAND3_X1  g0253(.A1(new_n265), .A2(new_n452), .A3(new_n453), .ZN(new_n454));
  INV_X1    g0254(.A(new_n454), .ZN(new_n455));
  NOR2_X1   g0255(.A1(new_n268), .A2(G1), .ZN(new_n456));
  INV_X1    g0256(.A(KEYINPUT5), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n457), .A2(G41), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n272), .A2(KEYINPUT5), .ZN(new_n459));
  NAND3_X1  g0259(.A1(new_n456), .A2(new_n458), .A3(new_n459), .ZN(new_n460));
  NAND3_X1  g0260(.A1(new_n460), .A2(G257), .A3(new_n265), .ZN(new_n461));
  INV_X1    g0261(.A(KEYINPUT75), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  NAND4_X1  g0263(.A1(new_n460), .A2(KEYINPUT75), .A3(G257), .A4(new_n265), .ZN(new_n464));
  AOI21_X1  g0264(.A(new_n455), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  OAI21_X1  g0265(.A(new_n451), .B1(new_n465), .B2(KEYINPUT76), .ZN(new_n466));
  INV_X1    g0266(.A(KEYINPUT76), .ZN(new_n467));
  AOI211_X1 g0267(.A(new_n467), .B(new_n455), .C1(new_n463), .C2(new_n464), .ZN(new_n468));
  NOR3_X1   g0268(.A1(new_n466), .A2(new_n468), .A3(G179), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n465), .A2(new_n451), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n470), .A2(new_n348), .ZN(new_n471));
  OAI21_X1  g0271(.A(G107), .B1(new_n379), .B2(new_n380), .ZN(new_n472));
  INV_X1    g0272(.A(KEYINPUT6), .ZN(new_n473));
  AND2_X1   g0273(.A1(G97), .A2(G107), .ZN(new_n474));
  NOR2_X1   g0274(.A1(G97), .A2(G107), .ZN(new_n475));
  OAI21_X1  g0275(.A(new_n473), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  NAND3_X1  g0276(.A1(new_n414), .A2(KEYINPUT6), .A3(G97), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  AOI22_X1  g0278(.A1(new_n478), .A2(G20), .B1(G77), .B2(new_n291), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n472), .A2(new_n479), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n480), .A2(new_n296), .ZN(new_n481));
  NOR2_X1   g0281(.A1(new_n304), .A2(G97), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n207), .A2(G33), .ZN(new_n483));
  NAND4_X1  g0283(.A1(new_n304), .A2(new_n483), .A3(new_n214), .A4(new_n295), .ZN(new_n484));
  INV_X1    g0284(.A(new_n484), .ZN(new_n485));
  AOI21_X1  g0285(.A(new_n482), .B1(new_n485), .B2(G97), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n481), .A2(new_n486), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n471), .A2(new_n487), .ZN(new_n488));
  NOR2_X1   g0288(.A1(new_n469), .A2(new_n488), .ZN(new_n489));
  OAI21_X1  g0289(.A(G200), .B1(new_n466), .B2(new_n468), .ZN(new_n490));
  INV_X1    g0290(.A(new_n486), .ZN(new_n491));
  AOI21_X1  g0291(.A(new_n491), .B1(new_n480), .B2(new_n296), .ZN(new_n492));
  NAND3_X1  g0292(.A1(new_n465), .A2(new_n451), .A3(G190), .ZN(new_n493));
  AND2_X1   g0293(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n490), .A2(new_n494), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n495), .A2(KEYINPUT77), .ZN(new_n496));
  INV_X1    g0296(.A(KEYINPUT77), .ZN(new_n497));
  NAND3_X1  g0297(.A1(new_n490), .A2(new_n494), .A3(new_n497), .ZN(new_n498));
  AOI21_X1  g0298(.A(new_n489), .B1(new_n496), .B2(new_n498), .ZN(new_n499));
  INV_X1    g0299(.A(KEYINPUT83), .ZN(new_n500));
  NAND3_X1  g0300(.A1(new_n429), .A2(KEYINPUT25), .A3(new_n414), .ZN(new_n501));
  INV_X1    g0301(.A(KEYINPUT25), .ZN(new_n502));
  OAI21_X1  g0302(.A(new_n502), .B1(new_n304), .B2(G107), .ZN(new_n503));
  AOI22_X1  g0303(.A1(G107), .A2(new_n485), .B1(new_n501), .B2(new_n503), .ZN(new_n504));
  INV_X1    g0304(.A(new_n504), .ZN(new_n505));
  AOI21_X1  g0305(.A(KEYINPUT23), .B1(new_n414), .B2(G20), .ZN(new_n506));
  INV_X1    g0306(.A(new_n506), .ZN(new_n507));
  NAND3_X1  g0307(.A1(new_n414), .A2(KEYINPUT23), .A3(G20), .ZN(new_n508));
  AOI22_X1  g0308(.A1(new_n507), .A2(new_n508), .B1(new_n425), .B2(G116), .ZN(new_n509));
  NAND3_X1  g0309(.A1(new_n208), .A2(KEYINPUT82), .A3(G87), .ZN(new_n510));
  NOR3_X1   g0310(.A1(new_n334), .A2(KEYINPUT22), .A3(new_n510), .ZN(new_n511));
  INV_X1    g0311(.A(KEYINPUT22), .ZN(new_n512));
  AND3_X1   g0312(.A1(new_n208), .A2(KEYINPUT82), .A3(G87), .ZN(new_n513));
  AOI21_X1  g0313(.A(new_n512), .B1(new_n331), .B2(new_n513), .ZN(new_n514));
  OAI21_X1  g0314(.A(new_n509), .B1(new_n511), .B2(new_n514), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n515), .A2(KEYINPUT24), .ZN(new_n516));
  OAI21_X1  g0316(.A(KEYINPUT22), .B1(new_n334), .B2(new_n510), .ZN(new_n517));
  NAND3_X1  g0317(.A1(new_n331), .A2(new_n512), .A3(new_n513), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  INV_X1    g0319(.A(KEYINPUT24), .ZN(new_n520));
  NAND3_X1  g0320(.A1(new_n519), .A2(new_n520), .A3(new_n509), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n516), .A2(new_n521), .ZN(new_n522));
  AOI21_X1  g0322(.A(new_n505), .B1(new_n522), .B2(new_n296), .ZN(new_n523));
  OAI211_X1 g0323(.A(G250), .B(new_n256), .C1(new_n253), .C2(new_n254), .ZN(new_n524));
  OAI211_X1 g0324(.A(G257), .B(G1698), .C1(new_n253), .C2(new_n254), .ZN(new_n525));
  NAND2_X1  g0325(.A1(G33), .A2(G294), .ZN(new_n526));
  NAND3_X1  g0326(.A1(new_n524), .A2(new_n525), .A3(new_n526), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n527), .A2(new_n261), .ZN(new_n528));
  AOI22_X1  g0328(.A1(new_n452), .A2(new_n456), .B1(new_n263), .B2(new_n264), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n529), .A2(G264), .ZN(new_n530));
  NAND3_X1  g0330(.A1(new_n528), .A2(new_n454), .A3(new_n530), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n531), .A2(new_n348), .ZN(new_n532));
  AOI22_X1  g0332(.A1(new_n527), .A2(new_n261), .B1(new_n529), .B2(G264), .ZN(new_n533));
  NAND3_X1  g0333(.A1(new_n533), .A2(new_n437), .A3(new_n454), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n532), .A2(new_n534), .ZN(new_n535));
  OAI21_X1  g0335(.A(new_n500), .B1(new_n523), .B2(new_n535), .ZN(new_n536));
  NAND3_X1  g0336(.A1(new_n208), .A2(G33), .A3(G116), .ZN(new_n537));
  AND3_X1   g0337(.A1(new_n414), .A2(KEYINPUT23), .A3(G20), .ZN(new_n538));
  OAI21_X1  g0338(.A(new_n537), .B1(new_n538), .B2(new_n506), .ZN(new_n539));
  AOI211_X1 g0339(.A(KEYINPUT24), .B(new_n539), .C1(new_n517), .C2(new_n518), .ZN(new_n540));
  AOI21_X1  g0340(.A(new_n520), .B1(new_n519), .B2(new_n509), .ZN(new_n541));
  OAI21_X1  g0341(.A(new_n296), .B1(new_n540), .B2(new_n541), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n542), .A2(new_n504), .ZN(new_n543));
  AND4_X1   g0343(.A1(new_n437), .A2(new_n528), .A3(new_n454), .A4(new_n530), .ZN(new_n544));
  AOI21_X1  g0344(.A(G169), .B1(new_n533), .B2(new_n454), .ZN(new_n545));
  NOR2_X1   g0345(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  NAND3_X1  g0346(.A1(new_n543), .A2(new_n546), .A3(KEYINPUT83), .ZN(new_n547));
  NAND3_X1  g0347(.A1(new_n533), .A2(G190), .A3(new_n454), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n531), .A2(G200), .ZN(new_n549));
  NAND4_X1  g0349(.A1(new_n542), .A2(new_n504), .A3(new_n548), .A4(new_n549), .ZN(new_n550));
  NAND3_X1  g0350(.A1(new_n536), .A2(new_n547), .A3(new_n550), .ZN(new_n551));
  INV_X1    g0351(.A(new_n551), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n256), .A2(G257), .ZN(new_n553));
  NAND2_X1  g0353(.A1(G264), .A2(G1698), .ZN(new_n554));
  OAI211_X1 g0354(.A(new_n553), .B(new_n554), .C1(new_n253), .C2(new_n254), .ZN(new_n555));
  OAI211_X1 g0355(.A(new_n555), .B(new_n261), .C1(G303), .C2(new_n331), .ZN(new_n556));
  NAND3_X1  g0356(.A1(new_n460), .A2(G270), .A3(new_n265), .ZN(new_n557));
  NAND3_X1  g0357(.A1(new_n556), .A2(new_n454), .A3(new_n557), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n558), .A2(G169), .ZN(new_n559));
  INV_X1    g0359(.A(G116), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n429), .A2(new_n560), .ZN(new_n561));
  OAI21_X1  g0361(.A(new_n561), .B1(new_n484), .B2(new_n560), .ZN(new_n562));
  OAI211_X1 g0362(.A(new_n446), .B(new_n208), .C1(G33), .C2(new_n259), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n560), .A2(G20), .ZN(new_n564));
  NAND3_X1  g0364(.A1(new_n563), .A2(new_n296), .A3(new_n564), .ZN(new_n565));
  INV_X1    g0365(.A(KEYINPUT20), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  NAND4_X1  g0367(.A1(new_n563), .A2(KEYINPUT20), .A3(new_n296), .A4(new_n564), .ZN(new_n568));
  AOI21_X1  g0368(.A(new_n562), .B1(new_n567), .B2(new_n568), .ZN(new_n569));
  OAI21_X1  g0369(.A(KEYINPUT81), .B1(new_n559), .B2(new_n569), .ZN(new_n570));
  INV_X1    g0370(.A(KEYINPUT21), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  OAI211_X1 g0372(.A(KEYINPUT81), .B(KEYINPUT21), .C1(new_n559), .C2(new_n569), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  INV_X1    g0374(.A(new_n558), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n575), .A2(G179), .ZN(new_n576));
  OAI21_X1  g0376(.A(KEYINPUT80), .B1(new_n576), .B2(new_n569), .ZN(new_n577));
  INV_X1    g0377(.A(new_n569), .ZN(new_n578));
  NOR2_X1   g0378(.A1(new_n558), .A2(new_n437), .ZN(new_n579));
  INV_X1    g0379(.A(KEYINPUT80), .ZN(new_n580));
  NAND3_X1  g0380(.A1(new_n578), .A2(new_n579), .A3(new_n580), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n577), .A2(new_n581), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n558), .A2(G200), .ZN(new_n583));
  OAI211_X1 g0383(.A(new_n583), .B(new_n569), .C1(new_n433), .C2(new_n558), .ZN(new_n584));
  NAND3_X1  g0384(.A1(new_n574), .A2(new_n582), .A3(new_n584), .ZN(new_n585));
  NOR2_X1   g0385(.A1(new_n424), .A2(new_n304), .ZN(new_n586));
  NAND3_X1  g0386(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n587), .A2(new_n208), .ZN(new_n588));
  NAND3_X1  g0388(.A1(new_n221), .A2(new_n259), .A3(new_n414), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  NOR2_X1   g0390(.A1(new_n227), .A2(G20), .ZN(new_n591));
  OAI21_X1  g0391(.A(new_n591), .B1(new_n253), .B2(new_n254), .ZN(new_n592));
  INV_X1    g0392(.A(KEYINPUT19), .ZN(new_n593));
  OAI21_X1  g0393(.A(new_n593), .B1(new_n290), .B2(new_n259), .ZN(new_n594));
  NAND3_X1  g0394(.A1(new_n590), .A2(new_n592), .A3(new_n594), .ZN(new_n595));
  AOI21_X1  g0395(.A(new_n586), .B1(new_n595), .B2(new_n296), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n485), .A2(G87), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  NOR2_X1   g0398(.A1(new_n228), .A2(G1698), .ZN(new_n599));
  OAI21_X1  g0399(.A(new_n599), .B1(new_n253), .B2(new_n254), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n600), .A2(KEYINPUT78), .ZN(new_n601));
  NAND3_X1  g0401(.A1(new_n331), .A2(G244), .A3(G1698), .ZN(new_n602));
  NAND2_X1  g0402(.A1(G33), .A2(G116), .ZN(new_n603));
  INV_X1    g0403(.A(KEYINPUT78), .ZN(new_n604));
  OAI211_X1 g0404(.A(new_n599), .B(new_n604), .C1(new_n254), .C2(new_n253), .ZN(new_n605));
  NAND4_X1  g0405(.A1(new_n601), .A2(new_n602), .A3(new_n603), .A4(new_n605), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n606), .A2(new_n261), .ZN(new_n607));
  NOR2_X1   g0407(.A1(new_n456), .A2(new_n222), .ZN(new_n608));
  OAI21_X1  g0408(.A(new_n265), .B1(new_n608), .B2(new_n453), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n607), .A2(new_n609), .ZN(new_n610));
  AOI21_X1  g0410(.A(new_n598), .B1(new_n610), .B2(G200), .ZN(new_n611));
  INV_X1    g0411(.A(new_n609), .ZN(new_n612));
  AOI21_X1  g0412(.A(new_n612), .B1(new_n606), .B2(new_n261), .ZN(new_n613));
  AND3_X1   g0413(.A1(new_n613), .A2(KEYINPUT79), .A3(G190), .ZN(new_n614));
  AOI21_X1  g0414(.A(KEYINPUT79), .B1(new_n613), .B2(G190), .ZN(new_n615));
  OAI21_X1  g0415(.A(new_n611), .B1(new_n614), .B2(new_n615), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n485), .A2(new_n424), .ZN(new_n617));
  AOI22_X1  g0417(.A1(new_n610), .A2(new_n348), .B1(new_n596), .B2(new_n617), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n613), .A2(new_n437), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n616), .A2(new_n620), .ZN(new_n621));
  NOR2_X1   g0421(.A1(new_n585), .A2(new_n621), .ZN(new_n622));
  AND4_X1   g0422(.A1(new_n442), .A2(new_n499), .A3(new_n552), .A4(new_n622), .ZN(G372));
  NAND2_X1  g0423(.A1(new_n595), .A2(new_n296), .ZN(new_n624));
  INV_X1    g0424(.A(new_n586), .ZN(new_n625));
  AND4_X1   g0425(.A1(KEYINPUT84), .A2(new_n624), .A3(new_n625), .A4(new_n597), .ZN(new_n626));
  AOI21_X1  g0426(.A(KEYINPUT84), .B1(new_n596), .B2(new_n597), .ZN(new_n627));
  NOR2_X1   g0427(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n610), .A2(G200), .ZN(new_n629));
  OAI211_X1 g0429(.A(new_n628), .B(new_n629), .C1(new_n614), .C2(new_n615), .ZN(new_n630));
  AND3_X1   g0430(.A1(new_n630), .A2(new_n550), .A3(new_n620), .ZN(new_n631));
  AOI22_X1  g0431(.A1(new_n572), .A2(new_n573), .B1(new_n577), .B2(new_n581), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n543), .A2(new_n546), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n631), .A2(new_n634), .ZN(new_n635));
  INV_X1    g0435(.A(new_n466), .ZN(new_n636));
  INV_X1    g0436(.A(new_n468), .ZN(new_n637));
  NAND3_X1  g0437(.A1(new_n636), .A2(new_n437), .A3(new_n637), .ZN(new_n638));
  AOI21_X1  g0438(.A(new_n492), .B1(new_n348), .B2(new_n470), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  INV_X1    g0440(.A(new_n498), .ZN(new_n641));
  AOI21_X1  g0441(.A(new_n497), .B1(new_n490), .B2(new_n494), .ZN(new_n642));
  OAI21_X1  g0442(.A(new_n640), .B1(new_n641), .B2(new_n642), .ZN(new_n643));
  OAI21_X1  g0443(.A(KEYINPUT85), .B1(new_n635), .B2(new_n643), .ZN(new_n644));
  OAI21_X1  g0444(.A(KEYINPUT26), .B1(new_n621), .B2(new_n640), .ZN(new_n645));
  INV_X1    g0445(.A(KEYINPUT26), .ZN(new_n646));
  NAND4_X1  g0446(.A1(new_n489), .A2(new_n646), .A3(new_n620), .A4(new_n630), .ZN(new_n647));
  NAND3_X1  g0447(.A1(new_n645), .A2(new_n647), .A3(new_n620), .ZN(new_n648));
  INV_X1    g0448(.A(new_n648), .ZN(new_n649));
  INV_X1    g0449(.A(KEYINPUT85), .ZN(new_n650));
  NAND4_X1  g0450(.A1(new_n499), .A2(new_n650), .A3(new_n634), .A4(new_n631), .ZN(new_n651));
  NAND3_X1  g0451(.A1(new_n644), .A2(new_n649), .A3(new_n651), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n442), .A2(new_n652), .ZN(new_n653));
  INV_X1    g0453(.A(new_n350), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n398), .A2(new_n437), .ZN(new_n655));
  OAI21_X1  g0455(.A(new_n655), .B1(G169), .B2(new_n398), .ZN(new_n656));
  OAI21_X1  g0456(.A(KEYINPUT18), .B1(new_n407), .B2(new_n656), .ZN(new_n657));
  NAND3_X1  g0457(.A1(new_n367), .A2(new_n393), .A3(new_n394), .ZN(new_n658));
  NAND3_X1  g0458(.A1(new_n657), .A2(KEYINPUT86), .A3(new_n658), .ZN(new_n659));
  INV_X1    g0459(.A(KEYINPUT86), .ZN(new_n660));
  OAI21_X1  g0460(.A(new_n660), .B1(new_n395), .B2(new_n396), .ZN(new_n661));
  INV_X1    g0461(.A(new_n440), .ZN(new_n662));
  AOI22_X1  g0462(.A1(new_n288), .A2(new_n309), .B1(new_n314), .B2(new_n662), .ZN(new_n663));
  INV_X1    g0463(.A(new_n410), .ZN(new_n664));
  OAI211_X1 g0464(.A(new_n659), .B(new_n661), .C1(new_n663), .C2(new_n664), .ZN(new_n665));
  INV_X1    g0465(.A(KEYINPUT87), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n345), .A2(new_n666), .ZN(new_n667));
  NAND3_X1  g0467(.A1(new_n342), .A2(KEYINPUT87), .A3(new_n344), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  AOI21_X1  g0469(.A(new_n654), .B1(new_n665), .B2(new_n669), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n653), .A2(new_n670), .ZN(G369));
  INV_X1    g0471(.A(G330), .ZN(new_n672));
  INV_X1    g0472(.A(KEYINPUT89), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n585), .A2(new_n673), .ZN(new_n674));
  NAND3_X1  g0474(.A1(new_n632), .A2(KEYINPUT89), .A3(new_n584), .ZN(new_n675));
  NAND3_X1  g0475(.A1(new_n207), .A2(new_n208), .A3(G13), .ZN(new_n676));
  OR2_X1    g0476(.A1(new_n676), .A2(KEYINPUT27), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n676), .A2(KEYINPUT27), .ZN(new_n678));
  NAND3_X1  g0478(.A1(new_n677), .A2(new_n678), .A3(G213), .ZN(new_n679));
  INV_X1    g0479(.A(G343), .ZN(new_n680));
  NOR2_X1   g0480(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  INV_X1    g0481(.A(new_n681), .ZN(new_n682));
  NOR2_X1   g0482(.A1(new_n682), .A2(new_n569), .ZN(new_n683));
  INV_X1    g0483(.A(new_n683), .ZN(new_n684));
  NAND3_X1  g0484(.A1(new_n674), .A2(new_n675), .A3(new_n684), .ZN(new_n685));
  INV_X1    g0485(.A(KEYINPUT88), .ZN(new_n686));
  OAI21_X1  g0486(.A(new_n686), .B1(new_n632), .B2(new_n684), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n574), .A2(new_n582), .ZN(new_n688));
  NAND3_X1  g0488(.A1(new_n688), .A2(KEYINPUT88), .A3(new_n683), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n687), .A2(new_n689), .ZN(new_n690));
  AOI21_X1  g0490(.A(new_n672), .B1(new_n685), .B2(new_n690), .ZN(new_n691));
  OAI21_X1  g0491(.A(new_n552), .B1(new_n523), .B2(new_n682), .ZN(new_n692));
  OAI21_X1  g0492(.A(new_n692), .B1(new_n633), .B2(new_n682), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n691), .A2(new_n693), .ZN(new_n694));
  INV_X1    g0494(.A(KEYINPUT90), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  NAND3_X1  g0496(.A1(new_n691), .A2(new_n693), .A3(KEYINPUT90), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n688), .A2(new_n682), .ZN(new_n699));
  NOR2_X1   g0499(.A1(new_n699), .A2(new_n551), .ZN(new_n700));
  INV_X1    g0500(.A(new_n633), .ZN(new_n701));
  AOI21_X1  g0501(.A(new_n700), .B1(new_n701), .B2(new_n682), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n698), .A2(new_n702), .ZN(G399));
  INV_X1    g0503(.A(new_n211), .ZN(new_n704));
  NOR2_X1   g0504(.A1(new_n704), .A2(G41), .ZN(new_n705));
  INV_X1    g0505(.A(new_n705), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n706), .A2(G1), .ZN(new_n707));
  OR2_X1    g0507(.A1(new_n589), .A2(G116), .ZN(new_n708));
  OAI22_X1  g0508(.A1(new_n707), .A2(new_n708), .B1(new_n217), .B2(new_n706), .ZN(new_n709));
  XOR2_X1   g0509(.A(KEYINPUT91), .B(KEYINPUT28), .Z(new_n710));
  XNOR2_X1  g0510(.A(new_n709), .B(new_n710), .ZN(new_n711));
  NAND3_X1  g0511(.A1(new_n579), .A2(new_n533), .A3(new_n613), .ZN(new_n712));
  INV_X1    g0512(.A(KEYINPUT30), .ZN(new_n713));
  OR3_X1    g0513(.A1(new_n712), .A2(new_n713), .A3(new_n470), .ZN(new_n714));
  NOR3_X1   g0514(.A1(new_n613), .A2(new_n575), .A3(G179), .ZN(new_n715));
  OAI211_X1 g0515(.A(new_n715), .B(new_n531), .C1(new_n468), .C2(new_n466), .ZN(new_n716));
  OAI21_X1  g0516(.A(new_n713), .B1(new_n712), .B2(new_n470), .ZN(new_n717));
  NAND3_X1  g0517(.A1(new_n714), .A2(new_n716), .A3(new_n717), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n718), .A2(new_n681), .ZN(new_n719));
  XOR2_X1   g0519(.A(KEYINPUT92), .B(KEYINPUT31), .Z(new_n720));
  NOR2_X1   g0520(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  AOI21_X1  g0521(.A(KEYINPUT31), .B1(new_n718), .B2(new_n681), .ZN(new_n722));
  NOR2_X1   g0522(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  NAND4_X1  g0523(.A1(new_n499), .A2(new_n622), .A3(new_n552), .A4(new_n682), .ZN(new_n724));
  AOI21_X1  g0524(.A(new_n672), .B1(new_n723), .B2(new_n724), .ZN(new_n725));
  INV_X1    g0525(.A(new_n620), .ZN(new_n726));
  NAND3_X1  g0526(.A1(new_n630), .A2(new_n550), .A3(new_n620), .ZN(new_n727));
  NOR3_X1   g0527(.A1(new_n523), .A2(new_n535), .A3(new_n500), .ZN(new_n728));
  AOI21_X1  g0528(.A(KEYINPUT83), .B1(new_n543), .B2(new_n546), .ZN(new_n729));
  NOR2_X1   g0529(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  AOI21_X1  g0530(.A(new_n727), .B1(new_n730), .B2(new_n632), .ZN(new_n731));
  AOI21_X1  g0531(.A(new_n726), .B1(new_n731), .B2(new_n499), .ZN(new_n732));
  NAND4_X1  g0532(.A1(new_n630), .A2(new_n638), .A3(new_n639), .A4(new_n620), .ZN(new_n733));
  OAI21_X1  g0533(.A(KEYINPUT93), .B1(new_n733), .B2(new_n646), .ZN(new_n734));
  INV_X1    g0534(.A(new_n615), .ZN(new_n735));
  NAND3_X1  g0535(.A1(new_n613), .A2(KEYINPUT79), .A3(G190), .ZN(new_n736));
  NAND2_X1  g0536(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  NOR2_X1   g0537(.A1(new_n613), .A2(new_n399), .ZN(new_n738));
  NOR3_X1   g0538(.A1(new_n738), .A2(new_n627), .A3(new_n626), .ZN(new_n739));
  AOI22_X1  g0539(.A1(new_n737), .A2(new_n739), .B1(new_n619), .B2(new_n618), .ZN(new_n740));
  INV_X1    g0540(.A(KEYINPUT93), .ZN(new_n741));
  NAND4_X1  g0541(.A1(new_n740), .A2(new_n741), .A3(KEYINPUT26), .A4(new_n489), .ZN(new_n742));
  OAI21_X1  g0542(.A(new_n646), .B1(new_n621), .B2(new_n640), .ZN(new_n743));
  NAND3_X1  g0543(.A1(new_n734), .A2(new_n742), .A3(new_n743), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n732), .A2(new_n744), .ZN(new_n745));
  AOI21_X1  g0545(.A(KEYINPUT94), .B1(new_n745), .B2(new_n682), .ZN(new_n746));
  INV_X1    g0546(.A(KEYINPUT94), .ZN(new_n747));
  AOI211_X1 g0547(.A(new_n747), .B(new_n681), .C1(new_n732), .C2(new_n744), .ZN(new_n748));
  OAI21_X1  g0548(.A(KEYINPUT29), .B1(new_n746), .B2(new_n748), .ZN(new_n749));
  NAND2_X1  g0549(.A1(new_n652), .A2(new_n682), .ZN(new_n750));
  INV_X1    g0550(.A(KEYINPUT29), .ZN(new_n751));
  NAND2_X1  g0551(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  AOI21_X1  g0552(.A(new_n725), .B1(new_n749), .B2(new_n752), .ZN(new_n753));
  OAI21_X1  g0553(.A(new_n711), .B1(new_n753), .B2(G1), .ZN(G364));
  NOR2_X1   g0554(.A1(new_n301), .A2(G20), .ZN(new_n755));
  NAND2_X1  g0555(.A1(new_n755), .A2(G45), .ZN(new_n756));
  NAND3_X1  g0556(.A1(new_n706), .A2(G1), .A3(new_n756), .ZN(new_n757));
  XNOR2_X1  g0557(.A(new_n757), .B(KEYINPUT95), .ZN(new_n758));
  NOR2_X1   g0558(.A1(G179), .A2(G200), .ZN(new_n759));
  AOI21_X1  g0559(.A(new_n208), .B1(new_n759), .B2(G190), .ZN(new_n760));
  INV_X1    g0560(.A(G294), .ZN(new_n761));
  INV_X1    g0561(.A(G283), .ZN(new_n762));
  NOR2_X1   g0562(.A1(new_n208), .A2(G190), .ZN(new_n763));
  NOR2_X1   g0563(.A1(new_n399), .A2(G179), .ZN(new_n764));
  NAND2_X1  g0564(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  OAI221_X1 g0565(.A(new_n334), .B1(new_n760), .B2(new_n761), .C1(new_n762), .C2(new_n765), .ZN(new_n766));
  NOR2_X1   g0566(.A1(new_n208), .A2(new_n433), .ZN(new_n767));
  NOR2_X1   g0567(.A1(new_n437), .A2(G200), .ZN(new_n768));
  NAND2_X1  g0568(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  INV_X1    g0569(.A(new_n769), .ZN(new_n770));
  NAND2_X1  g0570(.A1(new_n763), .A2(new_n759), .ZN(new_n771));
  INV_X1    g0571(.A(new_n771), .ZN(new_n772));
  AOI22_X1  g0572(.A1(G322), .A2(new_n770), .B1(new_n772), .B2(G329), .ZN(new_n773));
  INV_X1    g0573(.A(G303), .ZN(new_n774));
  NAND2_X1  g0574(.A1(new_n767), .A2(new_n764), .ZN(new_n775));
  INV_X1    g0575(.A(G311), .ZN(new_n776));
  NAND2_X1  g0576(.A1(new_n763), .A2(new_n768), .ZN(new_n777));
  OAI221_X1 g0577(.A(new_n773), .B1(new_n774), .B2(new_n775), .C1(new_n776), .C2(new_n777), .ZN(new_n778));
  NOR2_X1   g0578(.A1(new_n208), .A2(new_n437), .ZN(new_n779));
  NAND3_X1  g0579(.A1(new_n779), .A2(new_n433), .A3(G200), .ZN(new_n780));
  INV_X1    g0580(.A(new_n780), .ZN(new_n781));
  XNOR2_X1  g0581(.A(KEYINPUT33), .B(G317), .ZN(new_n782));
  AOI211_X1 g0582(.A(new_n766), .B(new_n778), .C1(new_n781), .C2(new_n782), .ZN(new_n783));
  NAND3_X1  g0583(.A1(new_n779), .A2(G190), .A3(G200), .ZN(new_n784));
  XOR2_X1   g0584(.A(new_n784), .B(KEYINPUT98), .Z(new_n785));
  INV_X1    g0585(.A(new_n785), .ZN(new_n786));
  NAND2_X1  g0586(.A1(new_n786), .A2(G326), .ZN(new_n787));
  XOR2_X1   g0587(.A(new_n760), .B(KEYINPUT97), .Z(new_n788));
  NAND2_X1  g0588(.A1(new_n788), .A2(G97), .ZN(new_n789));
  NAND2_X1  g0589(.A1(new_n772), .A2(G159), .ZN(new_n790));
  NAND2_X1  g0590(.A1(new_n790), .A2(KEYINPUT32), .ZN(new_n791));
  OAI221_X1 g0591(.A(new_n791), .B1(new_n293), .B2(new_n784), .C1(new_n227), .C2(new_n780), .ZN(new_n792));
  INV_X1    g0592(.A(new_n775), .ZN(new_n793));
  INV_X1    g0593(.A(new_n765), .ZN(new_n794));
  AOI22_X1  g0594(.A1(G87), .A2(new_n793), .B1(new_n794), .B2(G107), .ZN(new_n795));
  OAI21_X1  g0595(.A(new_n795), .B1(new_n225), .B2(new_n769), .ZN(new_n796));
  OAI221_X1 g0596(.A(new_n331), .B1(new_n219), .B2(new_n777), .C1(new_n790), .C2(KEYINPUT32), .ZN(new_n797));
  NOR3_X1   g0597(.A1(new_n792), .A2(new_n796), .A3(new_n797), .ZN(new_n798));
  AOI22_X1  g0598(.A1(new_n783), .A2(new_n787), .B1(new_n789), .B2(new_n798), .ZN(new_n799));
  AOI21_X1  g0599(.A(new_n214), .B1(G20), .B2(new_n348), .ZN(new_n800));
  INV_X1    g0600(.A(new_n800), .ZN(new_n801));
  OAI21_X1  g0601(.A(new_n758), .B1(new_n799), .B2(new_n801), .ZN(new_n802));
  NOR2_X1   g0602(.A1(new_n704), .A2(new_n331), .ZN(new_n803));
  AND2_X1   g0603(.A1(new_n269), .A2(new_n271), .ZN(new_n804));
  INV_X1    g0604(.A(new_n804), .ZN(new_n805));
  OAI221_X1 g0605(.A(new_n803), .B1(new_n217), .B2(new_n805), .C1(new_n247), .C2(new_n268), .ZN(new_n806));
  NOR2_X1   g0606(.A1(new_n704), .A2(new_n334), .ZN(new_n807));
  AOI22_X1  g0607(.A1(new_n807), .A2(G355), .B1(new_n560), .B2(new_n704), .ZN(new_n808));
  NAND2_X1  g0608(.A1(new_n806), .A2(new_n808), .ZN(new_n809));
  OR2_X1    g0609(.A1(new_n809), .A2(KEYINPUT96), .ZN(new_n810));
  NOR2_X1   g0610(.A1(G13), .A2(G33), .ZN(new_n811));
  INV_X1    g0611(.A(new_n811), .ZN(new_n812));
  NOR2_X1   g0612(.A1(new_n812), .A2(G20), .ZN(new_n813));
  NOR2_X1   g0613(.A1(new_n813), .A2(new_n800), .ZN(new_n814));
  INV_X1    g0614(.A(new_n814), .ZN(new_n815));
  AOI21_X1  g0615(.A(new_n815), .B1(new_n809), .B2(KEYINPUT96), .ZN(new_n816));
  AOI21_X1  g0616(.A(new_n802), .B1(new_n810), .B2(new_n816), .ZN(new_n817));
  NAND3_X1  g0617(.A1(new_n685), .A2(new_n690), .A3(new_n813), .ZN(new_n818));
  NAND2_X1  g0618(.A1(new_n817), .A2(new_n818), .ZN(new_n819));
  NOR2_X1   g0619(.A1(new_n691), .A2(new_n758), .ZN(new_n820));
  NAND3_X1  g0620(.A1(new_n685), .A2(new_n690), .A3(new_n672), .ZN(new_n821));
  NAND2_X1  g0621(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  AND2_X1   g0622(.A1(new_n819), .A2(new_n822), .ZN(new_n823));
  INV_X1    g0623(.A(new_n823), .ZN(G396));
  NAND2_X1  g0624(.A1(new_n496), .A2(new_n498), .ZN(new_n825));
  NAND4_X1  g0625(.A1(new_n825), .A2(new_n640), .A3(new_n634), .A4(new_n631), .ZN(new_n826));
  AOI21_X1  g0626(.A(new_n648), .B1(new_n826), .B2(KEYINPUT85), .ZN(new_n827));
  AOI21_X1  g0627(.A(new_n681), .B1(new_n827), .B2(new_n651), .ZN(new_n828));
  NAND2_X1  g0628(.A1(new_n440), .A2(KEYINPUT101), .ZN(new_n829));
  NAND2_X1  g0629(.A1(new_n439), .A2(new_n681), .ZN(new_n830));
  XNOR2_X1  g0630(.A(new_n830), .B(KEYINPUT102), .ZN(new_n831));
  INV_X1    g0631(.A(KEYINPUT101), .ZN(new_n832));
  NAND4_X1  g0632(.A1(new_n436), .A2(new_n438), .A3(new_n832), .A4(new_n439), .ZN(new_n833));
  NAND4_X1  g0633(.A1(new_n829), .A2(new_n434), .A3(new_n831), .A4(new_n833), .ZN(new_n834));
  NAND2_X1  g0634(.A1(new_n662), .A2(new_n681), .ZN(new_n835));
  NAND2_X1  g0635(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  OAI21_X1  g0636(.A(KEYINPUT103), .B1(new_n828), .B2(new_n836), .ZN(new_n837));
  INV_X1    g0637(.A(KEYINPUT103), .ZN(new_n838));
  INV_X1    g0638(.A(new_n836), .ZN(new_n839));
  NAND3_X1  g0639(.A1(new_n750), .A2(new_n838), .A3(new_n839), .ZN(new_n840));
  INV_X1    g0640(.A(new_n834), .ZN(new_n841));
  NAND3_X1  g0641(.A1(new_n652), .A2(new_n682), .A3(new_n841), .ZN(new_n842));
  NAND3_X1  g0642(.A1(new_n837), .A2(new_n840), .A3(new_n842), .ZN(new_n843));
  INV_X1    g0643(.A(new_n725), .ZN(new_n844));
  AOI21_X1  g0644(.A(new_n758), .B1(new_n843), .B2(new_n844), .ZN(new_n845));
  OAI21_X1  g0645(.A(new_n845), .B1(new_n844), .B2(new_n843), .ZN(new_n846));
  NOR2_X1   g0646(.A1(new_n800), .A2(new_n811), .ZN(new_n847));
  XNOR2_X1  g0647(.A(new_n847), .B(KEYINPUT99), .ZN(new_n848));
  OAI21_X1  g0648(.A(new_n758), .B1(G77), .B2(new_n848), .ZN(new_n849));
  XNOR2_X1  g0649(.A(new_n849), .B(KEYINPUT100), .ZN(new_n850));
  INV_X1    g0650(.A(new_n777), .ZN(new_n851));
  AOI22_X1  g0651(.A1(G143), .A2(new_n770), .B1(new_n851), .B2(G159), .ZN(new_n852));
  OAI21_X1  g0652(.A(new_n852), .B1(new_n317), .B2(new_n780), .ZN(new_n853));
  INV_X1    g0653(.A(new_n784), .ZN(new_n854));
  AOI21_X1  g0654(.A(new_n853), .B1(G137), .B2(new_n854), .ZN(new_n855));
  XOR2_X1   g0655(.A(new_n855), .B(KEYINPUT34), .Z(new_n856));
  INV_X1    g0656(.A(G132), .ZN(new_n857));
  OAI22_X1  g0657(.A1(new_n775), .A2(new_n293), .B1(new_n771), .B2(new_n857), .ZN(new_n858));
  NOR2_X1   g0658(.A1(new_n765), .A2(new_n227), .ZN(new_n859));
  NOR3_X1   g0659(.A1(new_n858), .A2(new_n334), .A3(new_n859), .ZN(new_n860));
  OAI211_X1 g0660(.A(new_n856), .B(new_n860), .C1(new_n225), .C2(new_n760), .ZN(new_n861));
  OAI221_X1 g0661(.A(new_n334), .B1(new_n769), .B2(new_n761), .C1(new_n774), .C2(new_n784), .ZN(new_n862));
  AOI21_X1  g0662(.A(new_n862), .B1(G283), .B2(new_n781), .ZN(new_n863));
  AOI22_X1  g0663(.A1(G107), .A2(new_n793), .B1(new_n851), .B2(G116), .ZN(new_n864));
  AOI22_X1  g0664(.A1(new_n794), .A2(G87), .B1(new_n772), .B2(G311), .ZN(new_n865));
  NAND4_X1  g0665(.A1(new_n863), .A2(new_n789), .A3(new_n864), .A4(new_n865), .ZN(new_n866));
  AND2_X1   g0666(.A1(new_n861), .A2(new_n866), .ZN(new_n867));
  OAI221_X1 g0667(.A(new_n850), .B1(new_n836), .B2(new_n812), .C1(new_n801), .C2(new_n867), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n846), .A2(new_n868), .ZN(G384));
  AOI211_X1 g0669(.A(new_n560), .B(new_n216), .C1(new_n478), .C2(KEYINPUT35), .ZN(new_n870));
  OAI21_X1  g0670(.A(new_n870), .B1(KEYINPUT35), .B2(new_n478), .ZN(new_n871));
  XOR2_X1   g0671(.A(new_n871), .B(KEYINPUT36), .Z(new_n872));
  OR3_X1    g0672(.A1(new_n217), .A2(new_n219), .A3(new_n374), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n201), .A2(G68), .ZN(new_n874));
  AOI211_X1 g0674(.A(new_n207), .B(G13), .C1(new_n873), .C2(new_n874), .ZN(new_n875));
  NOR2_X1   g0675(.A1(new_n872), .A2(new_n875), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n309), .A2(new_n681), .ZN(new_n877));
  NAND3_X1  g0677(.A1(new_n310), .A2(new_n314), .A3(new_n877), .ZN(new_n878));
  INV_X1    g0678(.A(new_n314), .ZN(new_n879));
  OAI211_X1 g0679(.A(new_n309), .B(new_n681), .C1(new_n288), .C2(new_n879), .ZN(new_n880));
  AOI21_X1  g0680(.A(new_n839), .B1(new_n878), .B2(new_n880), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n719), .A2(new_n720), .ZN(new_n882));
  INV_X1    g0682(.A(KEYINPUT31), .ZN(new_n883));
  OAI211_X1 g0683(.A(new_n724), .B(new_n882), .C1(new_n883), .C2(new_n719), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n881), .A2(new_n884), .ZN(new_n885));
  INV_X1    g0685(.A(KEYINPUT38), .ZN(new_n886));
  INV_X1    g0686(.A(KEYINPUT104), .ZN(new_n887));
  OAI21_X1  g0687(.A(new_n887), .B1(new_n407), .B2(new_n679), .ZN(new_n888));
  INV_X1    g0688(.A(new_n679), .ZN(new_n889));
  NAND3_X1  g0689(.A1(new_n393), .A2(KEYINPUT104), .A3(new_n889), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n888), .A2(new_n890), .ZN(new_n891));
  AOI21_X1  g0691(.A(new_n886), .B1(new_n411), .B2(new_n891), .ZN(new_n892));
  INV_X1    g0692(.A(KEYINPUT37), .ZN(new_n893));
  AOI21_X1  g0693(.A(KEYINPUT104), .B1(new_n393), .B2(new_n889), .ZN(new_n894));
  AOI211_X1 g0694(.A(new_n887), .B(new_n679), .C1(new_n384), .C2(new_n392), .ZN(new_n895));
  NOR2_X1   g0695(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n367), .A2(new_n393), .ZN(new_n897));
  AND2_X1   g0697(.A1(new_n897), .A2(new_n402), .ZN(new_n898));
  AOI21_X1  g0698(.A(new_n893), .B1(new_n896), .B2(new_n898), .ZN(new_n899));
  INV_X1    g0699(.A(KEYINPUT105), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n897), .A2(new_n402), .ZN(new_n901));
  NOR2_X1   g0701(.A1(new_n407), .A2(new_n679), .ZN(new_n902));
  NOR3_X1   g0702(.A1(new_n901), .A2(KEYINPUT37), .A3(new_n902), .ZN(new_n903));
  NOR3_X1   g0703(.A1(new_n899), .A2(new_n900), .A3(new_n903), .ZN(new_n904));
  OAI21_X1  g0704(.A(KEYINPUT37), .B1(new_n891), .B2(new_n901), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n393), .A2(new_n889), .ZN(new_n906));
  NAND3_X1  g0706(.A1(new_n898), .A2(new_n893), .A3(new_n906), .ZN(new_n907));
  AOI21_X1  g0707(.A(KEYINPUT105), .B1(new_n905), .B2(new_n907), .ZN(new_n908));
  OAI21_X1  g0708(.A(new_n892), .B1(new_n904), .B2(new_n908), .ZN(new_n909));
  OAI21_X1  g0709(.A(new_n900), .B1(new_n899), .B2(new_n903), .ZN(new_n910));
  NAND3_X1  g0710(.A1(new_n905), .A2(KEYINPUT105), .A3(new_n907), .ZN(new_n911));
  AOI22_X1  g0711(.A1(new_n910), .A2(new_n911), .B1(new_n411), .B2(new_n891), .ZN(new_n912));
  OAI21_X1  g0712(.A(new_n909), .B1(new_n912), .B2(KEYINPUT38), .ZN(new_n913));
  INV_X1    g0713(.A(KEYINPUT106), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  OAI211_X1 g0715(.A(new_n909), .B(KEYINPUT106), .C1(new_n912), .C2(KEYINPUT38), .ZN(new_n916));
  AOI21_X1  g0716(.A(new_n885), .B1(new_n915), .B2(new_n916), .ZN(new_n917));
  INV_X1    g0717(.A(KEYINPUT40), .ZN(new_n918));
  NAND3_X1  g0718(.A1(new_n661), .A2(new_n410), .A3(new_n659), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n919), .A2(new_n902), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n402), .A2(new_n906), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n897), .A2(new_n660), .ZN(new_n922));
  NAND3_X1  g0722(.A1(new_n367), .A2(new_n393), .A3(KEYINPUT86), .ZN(new_n923));
  AOI21_X1  g0723(.A(new_n921), .B1(new_n922), .B2(new_n923), .ZN(new_n924));
  OAI21_X1  g0724(.A(new_n907), .B1(new_n924), .B2(new_n893), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n920), .A2(new_n925), .ZN(new_n926));
  XOR2_X1   g0726(.A(KEYINPUT107), .B(KEYINPUT38), .Z(new_n927));
  NAND2_X1  g0727(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  AOI21_X1  g0728(.A(new_n918), .B1(new_n928), .B2(new_n909), .ZN(new_n929));
  INV_X1    g0729(.A(new_n929), .ZN(new_n930));
  OAI22_X1  g0730(.A1(new_n917), .A2(KEYINPUT40), .B1(new_n885), .B2(new_n930), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n442), .A2(new_n884), .ZN(new_n932));
  OR2_X1    g0732(.A1(new_n931), .A2(new_n932), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n933), .A2(G330), .ZN(new_n934));
  AOI21_X1  g0734(.A(new_n934), .B1(new_n931), .B2(new_n932), .ZN(new_n935));
  AOI21_X1  g0735(.A(new_n889), .B1(new_n661), .B2(new_n659), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n915), .A2(new_n916), .ZN(new_n937));
  INV_X1    g0737(.A(new_n829), .ZN(new_n938));
  INV_X1    g0738(.A(new_n833), .ZN(new_n939));
  OAI21_X1  g0739(.A(new_n682), .B1(new_n938), .B2(new_n939), .ZN(new_n940));
  INV_X1    g0740(.A(new_n940), .ZN(new_n941));
  AOI21_X1  g0741(.A(new_n941), .B1(new_n828), .B2(new_n841), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n878), .A2(new_n880), .ZN(new_n943));
  INV_X1    g0743(.A(new_n943), .ZN(new_n944));
  NOR2_X1   g0744(.A1(new_n942), .A2(new_n944), .ZN(new_n945));
  AOI21_X1  g0745(.A(new_n936), .B1(new_n937), .B2(new_n945), .ZN(new_n946));
  INV_X1    g0746(.A(KEYINPUT39), .ZN(new_n947));
  NAND3_X1  g0747(.A1(new_n928), .A2(new_n909), .A3(new_n947), .ZN(new_n948));
  INV_X1    g0748(.A(KEYINPUT108), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n948), .A2(new_n949), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n910), .A2(new_n911), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n411), .A2(new_n891), .ZN(new_n952));
  AOI21_X1  g0752(.A(KEYINPUT38), .B1(new_n951), .B2(new_n952), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n952), .A2(KEYINPUT38), .ZN(new_n954));
  AOI21_X1  g0754(.A(new_n954), .B1(new_n910), .B2(new_n911), .ZN(new_n955));
  OAI21_X1  g0755(.A(KEYINPUT39), .B1(new_n953), .B2(new_n955), .ZN(new_n956));
  NAND4_X1  g0756(.A1(new_n928), .A2(new_n909), .A3(KEYINPUT108), .A4(new_n947), .ZN(new_n957));
  NAND3_X1  g0757(.A1(new_n950), .A2(new_n956), .A3(new_n957), .ZN(new_n958));
  NOR2_X1   g0758(.A1(new_n310), .A2(new_n681), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n958), .A2(new_n959), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n946), .A2(new_n960), .ZN(new_n961));
  NAND3_X1  g0761(.A1(new_n749), .A2(new_n442), .A3(new_n752), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n962), .A2(new_n670), .ZN(new_n963));
  XNOR2_X1  g0763(.A(new_n961), .B(new_n963), .ZN(new_n964));
  INV_X1    g0764(.A(new_n964), .ZN(new_n965));
  OAI22_X1  g0765(.A1(new_n935), .A2(new_n965), .B1(new_n207), .B2(new_n755), .ZN(new_n966));
  AND2_X1   g0766(.A1(new_n935), .A2(new_n965), .ZN(new_n967));
  OAI21_X1  g0767(.A(new_n876), .B1(new_n966), .B2(new_n967), .ZN(G367));
  INV_X1    g0768(.A(new_n758), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n803), .A2(new_n241), .ZN(new_n970));
  AOI21_X1  g0770(.A(new_n815), .B1(new_n704), .B2(new_n424), .ZN(new_n971));
  AOI21_X1  g0771(.A(new_n969), .B1(new_n970), .B2(new_n971), .ZN(new_n972));
  NOR2_X1   g0772(.A1(new_n628), .A2(new_n682), .ZN(new_n973));
  MUX2_X1   g0773(.A(new_n740), .B(new_n726), .S(new_n973), .Z(new_n974));
  INV_X1    g0774(.A(new_n813), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n786), .A2(G143), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n788), .A2(G68), .ZN(new_n977));
  OAI22_X1  g0777(.A1(new_n775), .A2(new_n225), .B1(new_n777), .B2(new_n201), .ZN(new_n978));
  XOR2_X1   g0778(.A(KEYINPUT114), .B(G137), .Z(new_n979));
  OAI22_X1  g0779(.A1(new_n979), .A2(new_n771), .B1(new_n765), .B2(new_n219), .ZN(new_n980));
  NOR2_X1   g0780(.A1(new_n978), .A2(new_n980), .ZN(new_n981));
  OAI21_X1  g0781(.A(new_n331), .B1(new_n769), .B2(new_n317), .ZN(new_n982));
  AOI21_X1  g0782(.A(new_n982), .B1(G159), .B2(new_n781), .ZN(new_n983));
  NAND4_X1  g0783(.A1(new_n976), .A2(new_n977), .A3(new_n981), .A4(new_n983), .ZN(new_n984));
  AOI21_X1  g0784(.A(KEYINPUT46), .B1(new_n793), .B2(G116), .ZN(new_n985));
  AND3_X1   g0785(.A1(new_n793), .A2(KEYINPUT46), .A3(G116), .ZN(new_n986));
  AOI211_X1 g0786(.A(new_n985), .B(new_n986), .C1(G294), .C2(new_n781), .ZN(new_n987));
  OAI22_X1  g0787(.A1(new_n769), .A2(new_n774), .B1(new_n777), .B2(new_n762), .ZN(new_n988));
  INV_X1    g0788(.A(new_n760), .ZN(new_n989));
  AOI21_X1  g0789(.A(new_n988), .B1(G107), .B2(new_n989), .ZN(new_n990));
  OAI211_X1 g0790(.A(new_n987), .B(new_n990), .C1(new_n776), .C2(new_n785), .ZN(new_n991));
  NOR2_X1   g0791(.A1(new_n765), .A2(new_n259), .ZN(new_n992));
  XNOR2_X1  g0792(.A(KEYINPUT112), .B(G317), .ZN(new_n993));
  AOI211_X1 g0793(.A(new_n331), .B(new_n992), .C1(new_n772), .C2(new_n993), .ZN(new_n994));
  XNOR2_X1  g0794(.A(new_n994), .B(KEYINPUT113), .ZN(new_n995));
  OAI21_X1  g0795(.A(new_n984), .B1(new_n991), .B2(new_n995), .ZN(new_n996));
  XOR2_X1   g0796(.A(new_n996), .B(KEYINPUT47), .Z(new_n997));
  OAI221_X1 g0797(.A(new_n972), .B1(new_n974), .B2(new_n975), .C1(new_n997), .C2(new_n801), .ZN(new_n998));
  NAND2_X1  g0798(.A1(new_n756), .A2(G1), .ZN(new_n999));
  INV_X1    g0799(.A(KEYINPUT111), .ZN(new_n1000));
  NAND3_X1  g0800(.A1(new_n696), .A2(KEYINPUT110), .A3(new_n697), .ZN(new_n1001));
  INV_X1    g0801(.A(new_n1001), .ZN(new_n1002));
  OAI221_X1 g0802(.A(new_n640), .B1(new_n492), .B2(new_n682), .C1(new_n641), .C2(new_n642), .ZN(new_n1003));
  NAND2_X1  g0803(.A1(new_n489), .A2(new_n681), .ZN(new_n1004));
  NAND2_X1  g0804(.A1(new_n1003), .A2(new_n1004), .ZN(new_n1005));
  INV_X1    g0805(.A(new_n1005), .ZN(new_n1006));
  INV_X1    g0806(.A(new_n699), .ZN(new_n1007));
  NAND2_X1  g0807(.A1(new_n1007), .A2(new_n552), .ZN(new_n1008));
  OAI21_X1  g0808(.A(new_n1008), .B1(new_n633), .B2(new_n681), .ZN(new_n1009));
  INV_X1    g0809(.A(KEYINPUT109), .ZN(new_n1010));
  NAND3_X1  g0810(.A1(new_n1006), .A2(new_n1009), .A3(new_n1010), .ZN(new_n1011));
  OAI21_X1  g0811(.A(KEYINPUT109), .B1(new_n702), .B2(new_n1005), .ZN(new_n1012));
  NAND3_X1  g0812(.A1(new_n1011), .A2(new_n1012), .A3(KEYINPUT44), .ZN(new_n1013));
  INV_X1    g0813(.A(KEYINPUT45), .ZN(new_n1014));
  OAI21_X1  g0814(.A(new_n1014), .B1(new_n1006), .B2(new_n1009), .ZN(new_n1015));
  NAND3_X1  g0815(.A1(new_n702), .A2(new_n1005), .A3(KEYINPUT45), .ZN(new_n1016));
  NAND2_X1  g0816(.A1(new_n1015), .A2(new_n1016), .ZN(new_n1017));
  NAND2_X1  g0817(.A1(new_n1013), .A2(new_n1017), .ZN(new_n1018));
  AOI21_X1  g0818(.A(KEYINPUT44), .B1(new_n1011), .B2(new_n1012), .ZN(new_n1019));
  OAI21_X1  g0819(.A(new_n1002), .B1(new_n1018), .B2(new_n1019), .ZN(new_n1020));
  NAND2_X1  g0820(.A1(new_n1011), .A2(new_n1012), .ZN(new_n1021));
  INV_X1    g0821(.A(KEYINPUT44), .ZN(new_n1022));
  NAND2_X1  g0822(.A1(new_n1021), .A2(new_n1022), .ZN(new_n1023));
  NAND4_X1  g0823(.A1(new_n1023), .A2(new_n1001), .A3(new_n1013), .A4(new_n1017), .ZN(new_n1024));
  NAND2_X1  g0824(.A1(new_n1020), .A2(new_n1024), .ZN(new_n1025));
  OAI21_X1  g0825(.A(new_n1008), .B1(new_n693), .B2(new_n1007), .ZN(new_n1026));
  XNOR2_X1  g0826(.A(new_n1026), .B(new_n691), .ZN(new_n1027));
  NAND2_X1  g0827(.A1(new_n753), .A2(new_n1027), .ZN(new_n1028));
  OAI21_X1  g0828(.A(new_n1000), .B1(new_n1025), .B2(new_n1028), .ZN(new_n1029));
  INV_X1    g0829(.A(new_n1029), .ZN(new_n1030));
  NOR3_X1   g0830(.A1(new_n1025), .A2(new_n1028), .A3(new_n1000), .ZN(new_n1031));
  OAI21_X1  g0831(.A(new_n753), .B1(new_n1030), .B2(new_n1031), .ZN(new_n1032));
  XOR2_X1   g0832(.A(new_n705), .B(KEYINPUT41), .Z(new_n1033));
  INV_X1    g0833(.A(new_n1033), .ZN(new_n1034));
  AOI21_X1  g0834(.A(new_n999), .B1(new_n1032), .B2(new_n1034), .ZN(new_n1035));
  NAND2_X1  g0835(.A1(new_n1005), .A2(new_n700), .ZN(new_n1036));
  OR2_X1    g0836(.A1(new_n1036), .A2(KEYINPUT42), .ZN(new_n1037));
  OAI21_X1  g0837(.A(new_n640), .B1(new_n1003), .B2(new_n730), .ZN(new_n1038));
  AOI22_X1  g0838(.A1(new_n1036), .A2(KEYINPUT42), .B1(new_n1038), .B2(new_n682), .ZN(new_n1039));
  AOI22_X1  g0839(.A1(new_n1037), .A2(new_n1039), .B1(KEYINPUT43), .B2(new_n974), .ZN(new_n1040));
  NOR2_X1   g0840(.A1(new_n974), .A2(KEYINPUT43), .ZN(new_n1041));
  XOR2_X1   g0841(.A(new_n1040), .B(new_n1041), .Z(new_n1042));
  NOR2_X1   g0842(.A1(new_n698), .A2(new_n1006), .ZN(new_n1043));
  XNOR2_X1  g0843(.A(new_n1042), .B(new_n1043), .ZN(new_n1044));
  INV_X1    g0844(.A(new_n1044), .ZN(new_n1045));
  OAI21_X1  g0845(.A(new_n998), .B1(new_n1035), .B2(new_n1045), .ZN(G387));
  NOR2_X1   g0846(.A1(new_n693), .A2(new_n975), .ZN(new_n1047));
  AOI211_X1 g0847(.A(new_n334), .B(new_n992), .C1(G159), .C2(new_n854), .ZN(new_n1048));
  NAND2_X1  g0848(.A1(new_n788), .A2(new_n424), .ZN(new_n1049));
  OAI22_X1  g0849(.A1(new_n769), .A2(new_n293), .B1(new_n777), .B2(new_n227), .ZN(new_n1050));
  OAI22_X1  g0850(.A1(new_n775), .A2(new_n219), .B1(new_n771), .B2(new_n317), .ZN(new_n1051));
  NOR2_X1   g0851(.A1(new_n1050), .A2(new_n1051), .ZN(new_n1052));
  NAND2_X1  g0852(.A1(new_n781), .A2(new_n385), .ZN(new_n1053));
  NAND4_X1  g0853(.A1(new_n1048), .A2(new_n1049), .A3(new_n1052), .A4(new_n1053), .ZN(new_n1054));
  AOI22_X1  g0854(.A1(new_n770), .A2(new_n993), .B1(new_n851), .B2(G303), .ZN(new_n1055));
  XNOR2_X1  g0855(.A(KEYINPUT116), .B(G322), .ZN(new_n1056));
  OAI221_X1 g0856(.A(new_n1055), .B1(new_n776), .B2(new_n780), .C1(new_n785), .C2(new_n1056), .ZN(new_n1057));
  INV_X1    g0857(.A(KEYINPUT48), .ZN(new_n1058));
  OR2_X1    g0858(.A1(new_n1057), .A2(new_n1058), .ZN(new_n1059));
  OAI22_X1  g0859(.A1(new_n775), .A2(new_n761), .B1(new_n760), .B2(new_n762), .ZN(new_n1060));
  AOI21_X1  g0860(.A(new_n1060), .B1(new_n1057), .B2(new_n1058), .ZN(new_n1061));
  NAND3_X1  g0861(.A1(new_n1059), .A2(KEYINPUT49), .A3(new_n1061), .ZN(new_n1062));
  AOI21_X1  g0862(.A(new_n331), .B1(new_n772), .B2(G326), .ZN(new_n1063));
  OAI211_X1 g0863(.A(new_n1062), .B(new_n1063), .C1(new_n560), .C2(new_n765), .ZN(new_n1064));
  AOI21_X1  g0864(.A(KEYINPUT49), .B1(new_n1059), .B2(new_n1061), .ZN(new_n1065));
  OAI21_X1  g0865(.A(new_n1054), .B1(new_n1064), .B2(new_n1065), .ZN(new_n1066));
  NAND2_X1  g0866(.A1(new_n1066), .A2(new_n800), .ZN(new_n1067));
  INV_X1    g0867(.A(new_n803), .ZN(new_n1068));
  AOI21_X1  g0868(.A(new_n1068), .B1(new_n238), .B2(new_n805), .ZN(new_n1069));
  AOI21_X1  g0869(.A(new_n1069), .B1(new_n708), .B2(new_n807), .ZN(new_n1070));
  NAND2_X1  g0870(.A1(new_n385), .A2(new_n293), .ZN(new_n1071));
  XNOR2_X1  g0871(.A(new_n1071), .B(KEYINPUT50), .ZN(new_n1072));
  OAI21_X1  g0872(.A(new_n268), .B1(new_n227), .B2(new_n219), .ZN(new_n1073));
  NOR3_X1   g0873(.A1(new_n1072), .A2(new_n708), .A3(new_n1073), .ZN(new_n1074));
  OAI22_X1  g0874(.A1(new_n1070), .A2(new_n1074), .B1(G107), .B2(new_n211), .ZN(new_n1075));
  AOI21_X1  g0875(.A(new_n969), .B1(new_n1075), .B2(new_n814), .ZN(new_n1076));
  INV_X1    g0876(.A(KEYINPUT115), .ZN(new_n1077));
  OAI21_X1  g0877(.A(new_n1067), .B1(new_n1076), .B2(new_n1077), .ZN(new_n1078));
  AOI211_X1 g0878(.A(new_n1047), .B(new_n1078), .C1(new_n1077), .C2(new_n1076), .ZN(new_n1079));
  AOI21_X1  g0879(.A(new_n1079), .B1(new_n999), .B2(new_n1027), .ZN(new_n1080));
  NAND2_X1  g0880(.A1(new_n1028), .A2(new_n705), .ZN(new_n1081));
  NOR2_X1   g0881(.A1(new_n753), .A2(new_n1027), .ZN(new_n1082));
  OAI21_X1  g0882(.A(new_n1080), .B1(new_n1081), .B2(new_n1082), .ZN(G393));
  AOI22_X1  g0883(.A1(G68), .A2(new_n793), .B1(new_n772), .B2(G143), .ZN(new_n1084));
  XOR2_X1   g0884(.A(new_n1084), .B(KEYINPUT118), .Z(new_n1085));
  INV_X1    g0885(.A(G159), .ZN(new_n1086));
  OAI22_X1  g0886(.A1(new_n784), .A2(new_n317), .B1(new_n769), .B2(new_n1086), .ZN(new_n1087));
  XNOR2_X1  g0887(.A(KEYINPUT117), .B(KEYINPUT51), .ZN(new_n1088));
  INV_X1    g0888(.A(new_n1088), .ZN(new_n1089));
  AOI21_X1  g0889(.A(new_n1085), .B1(new_n1087), .B2(new_n1089), .ZN(new_n1090));
  NAND2_X1  g0890(.A1(new_n788), .A2(G77), .ZN(new_n1091));
  OAI221_X1 g0891(.A(new_n331), .B1(new_n777), .B2(new_n316), .C1(new_n221), .C2(new_n765), .ZN(new_n1092));
  AOI21_X1  g0892(.A(new_n1092), .B1(new_n202), .B2(new_n781), .ZN(new_n1093));
  OR2_X1    g0893(.A1(new_n1087), .A2(new_n1089), .ZN(new_n1094));
  NAND4_X1  g0894(.A1(new_n1090), .A2(new_n1091), .A3(new_n1093), .A4(new_n1094), .ZN(new_n1095));
  AOI21_X1  g0895(.A(new_n331), .B1(new_n794), .B2(G107), .ZN(new_n1096));
  OAI221_X1 g0896(.A(new_n1096), .B1(new_n762), .B2(new_n775), .C1(new_n771), .C2(new_n1056), .ZN(new_n1097));
  XNOR2_X1  g0897(.A(new_n1097), .B(KEYINPUT119), .ZN(new_n1098));
  AOI22_X1  g0898(.A1(new_n854), .A2(G317), .B1(new_n770), .B2(G311), .ZN(new_n1099));
  XOR2_X1   g0899(.A(new_n1099), .B(KEYINPUT52), .Z(new_n1100));
  OAI22_X1  g0900(.A1(new_n780), .A2(new_n774), .B1(new_n777), .B2(new_n761), .ZN(new_n1101));
  AOI21_X1  g0901(.A(new_n1101), .B1(G116), .B2(new_n989), .ZN(new_n1102));
  NAND3_X1  g0902(.A1(new_n1098), .A2(new_n1100), .A3(new_n1102), .ZN(new_n1103));
  AOI21_X1  g0903(.A(new_n801), .B1(new_n1095), .B2(new_n1103), .ZN(new_n1104));
  OR2_X1    g0904(.A1(new_n251), .A2(new_n1068), .ZN(new_n1105));
  AOI21_X1  g0905(.A(new_n815), .B1(G97), .B2(new_n704), .ZN(new_n1106));
  AOI211_X1 g0906(.A(new_n969), .B(new_n1104), .C1(new_n1105), .C2(new_n1106), .ZN(new_n1107));
  OAI21_X1  g0907(.A(new_n1107), .B1(new_n1005), .B2(new_n975), .ZN(new_n1108));
  NOR2_X1   g0908(.A1(new_n1018), .A2(new_n1019), .ZN(new_n1109));
  XNOR2_X1  g0909(.A(new_n1109), .B(new_n698), .ZN(new_n1110));
  INV_X1    g0910(.A(new_n999), .ZN(new_n1111));
  OAI21_X1  g0911(.A(new_n1108), .B1(new_n1110), .B2(new_n1111), .ZN(new_n1112));
  INV_X1    g0912(.A(new_n1031), .ZN(new_n1113));
  NAND2_X1  g0913(.A1(new_n1113), .A2(new_n1029), .ZN(new_n1114));
  AOI21_X1  g0914(.A(new_n706), .B1(new_n1110), .B2(new_n1028), .ZN(new_n1115));
  AOI21_X1  g0915(.A(new_n1112), .B1(new_n1114), .B2(new_n1115), .ZN(new_n1116));
  INV_X1    g0916(.A(new_n1116), .ZN(G390));
  OAI21_X1  g0917(.A(new_n836), .B1(new_n746), .B2(new_n748), .ZN(new_n1118));
  AOI21_X1  g0918(.A(new_n944), .B1(new_n1118), .B2(new_n940), .ZN(new_n1119));
  AOI21_X1  g0919(.A(new_n959), .B1(new_n928), .B2(new_n909), .ZN(new_n1120));
  INV_X1    g0920(.A(new_n1120), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n842), .A2(new_n940), .ZN(new_n1122));
  AOI21_X1  g0922(.A(new_n959), .B1(new_n1122), .B2(new_n943), .ZN(new_n1123));
  OAI22_X1  g0923(.A1(new_n1119), .A2(new_n1121), .B1(new_n958), .B2(new_n1123), .ZN(new_n1124));
  NAND2_X1  g0924(.A1(new_n884), .A2(G330), .ZN(new_n1125));
  NOR3_X1   g0925(.A1(new_n1125), .A2(new_n839), .A3(new_n944), .ZN(new_n1126));
  NAND2_X1  g0926(.A1(new_n1124), .A2(new_n1126), .ZN(new_n1127));
  AND3_X1   g0927(.A1(new_n734), .A2(new_n742), .A3(new_n743), .ZN(new_n1128));
  NAND3_X1  g0928(.A1(new_n632), .A2(new_n536), .A3(new_n547), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n1129), .A2(new_n631), .ZN(new_n1130));
  OAI21_X1  g0930(.A(new_n620), .B1(new_n1130), .B2(new_n643), .ZN(new_n1131));
  OAI21_X1  g0931(.A(new_n682), .B1(new_n1128), .B2(new_n1131), .ZN(new_n1132));
  NAND2_X1  g0932(.A1(new_n1132), .A2(new_n747), .ZN(new_n1133));
  NAND3_X1  g0933(.A1(new_n745), .A2(KEYINPUT94), .A3(new_n682), .ZN(new_n1134));
  NAND2_X1  g0934(.A1(new_n1133), .A2(new_n1134), .ZN(new_n1135));
  AOI21_X1  g0935(.A(new_n941), .B1(new_n1135), .B2(new_n836), .ZN(new_n1136));
  OAI21_X1  g0936(.A(new_n1120), .B1(new_n1136), .B2(new_n944), .ZN(new_n1137));
  INV_X1    g0937(.A(new_n959), .ZN(new_n1138));
  OAI21_X1  g0938(.A(new_n1138), .B1(new_n942), .B2(new_n944), .ZN(new_n1139));
  AOI22_X1  g0939(.A1(KEYINPUT39), .A2(new_n913), .B1(new_n948), .B2(new_n949), .ZN(new_n1140));
  NAND3_X1  g0940(.A1(new_n1139), .A2(new_n1140), .A3(new_n957), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n881), .A2(new_n725), .ZN(new_n1142));
  NAND3_X1  g0942(.A1(new_n1137), .A2(new_n1141), .A3(new_n1142), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n1127), .A2(new_n1143), .ZN(new_n1144));
  AOI21_X1  g0944(.A(new_n943), .B1(new_n725), .B2(new_n836), .ZN(new_n1145));
  OAI21_X1  g0945(.A(new_n1122), .B1(new_n1126), .B2(new_n1145), .ZN(new_n1146));
  INV_X1    g0946(.A(KEYINPUT120), .ZN(new_n1147));
  INV_X1    g0947(.A(new_n724), .ZN(new_n1148));
  OAI21_X1  g0948(.A(new_n882), .B1(new_n883), .B2(new_n719), .ZN(new_n1149));
  OAI211_X1 g0949(.A(G330), .B(new_n836), .C1(new_n1148), .C2(new_n1149), .ZN(new_n1150));
  AOI22_X1  g0950(.A1(new_n944), .A2(new_n1150), .B1(new_n881), .B2(new_n725), .ZN(new_n1151));
  AOI21_X1  g0951(.A(new_n1147), .B1(new_n1136), .B2(new_n1151), .ZN(new_n1152));
  AND4_X1   g0952(.A1(new_n1147), .A2(new_n1118), .A3(new_n1151), .A4(new_n940), .ZN(new_n1153));
  OAI21_X1  g0953(.A(new_n1146), .B1(new_n1152), .B2(new_n1153), .ZN(new_n1154));
  INV_X1    g0954(.A(new_n1125), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n1155), .A2(new_n442), .ZN(new_n1156));
  NAND3_X1  g0956(.A1(new_n962), .A2(new_n670), .A3(new_n1156), .ZN(new_n1157));
  INV_X1    g0957(.A(new_n1157), .ZN(new_n1158));
  NAND2_X1  g0958(.A1(new_n1154), .A2(new_n1158), .ZN(new_n1159));
  AOI21_X1  g0959(.A(new_n706), .B1(new_n1144), .B2(new_n1159), .ZN(new_n1160));
  INV_X1    g0960(.A(new_n1142), .ZN(new_n1161));
  NOR2_X1   g0961(.A1(new_n1124), .A2(new_n1161), .ZN(new_n1162));
  INV_X1    g0962(.A(new_n1126), .ZN(new_n1163));
  AOI21_X1  g0963(.A(new_n1163), .B1(new_n1137), .B2(new_n1141), .ZN(new_n1164));
  NOR2_X1   g0964(.A1(new_n1162), .A2(new_n1164), .ZN(new_n1165));
  NAND3_X1  g0965(.A1(new_n1136), .A2(new_n1147), .A3(new_n1151), .ZN(new_n1166));
  NAND3_X1  g0966(.A1(new_n1118), .A2(new_n1151), .A3(new_n940), .ZN(new_n1167));
  NAND2_X1  g0967(.A1(new_n1167), .A2(KEYINPUT120), .ZN(new_n1168));
  NAND2_X1  g0968(.A1(new_n1166), .A2(new_n1168), .ZN(new_n1169));
  AOI21_X1  g0969(.A(new_n1157), .B1(new_n1169), .B2(new_n1146), .ZN(new_n1170));
  NAND2_X1  g0970(.A1(new_n1165), .A2(new_n1170), .ZN(new_n1171));
  NAND2_X1  g0971(.A1(new_n1160), .A2(new_n1171), .ZN(new_n1172));
  NAND3_X1  g0972(.A1(new_n1140), .A2(new_n811), .A3(new_n957), .ZN(new_n1173));
  OAI21_X1  g0973(.A(new_n758), .B1(new_n385), .B2(new_n848), .ZN(new_n1174));
  XNOR2_X1  g0974(.A(new_n1174), .B(KEYINPUT121), .ZN(new_n1175));
  OAI22_X1  g0975(.A1(new_n777), .A2(new_n259), .B1(new_n771), .B2(new_n761), .ZN(new_n1176));
  AOI211_X1 g0976(.A(new_n859), .B(new_n1176), .C1(G116), .C2(new_n770), .ZN(new_n1177));
  OAI221_X1 g0977(.A(new_n334), .B1(new_n775), .B2(new_n221), .C1(new_n762), .C2(new_n784), .ZN(new_n1178));
  AOI21_X1  g0978(.A(new_n1178), .B1(G107), .B2(new_n781), .ZN(new_n1179));
  NAND3_X1  g0979(.A1(new_n1177), .A2(new_n1179), .A3(new_n1091), .ZN(new_n1180));
  INV_X1    g0980(.A(G128), .ZN(new_n1181));
  OAI22_X1  g0981(.A1(new_n780), .A2(new_n979), .B1(new_n784), .B2(new_n1181), .ZN(new_n1182));
  INV_X1    g0982(.A(G125), .ZN(new_n1183));
  OAI22_X1  g0983(.A1(new_n769), .A2(new_n857), .B1(new_n771), .B2(new_n1183), .ZN(new_n1184));
  XNOR2_X1  g0984(.A(KEYINPUT54), .B(G143), .ZN(new_n1185));
  NOR2_X1   g0985(.A1(new_n777), .A2(new_n1185), .ZN(new_n1186));
  NOR3_X1   g0986(.A1(new_n1182), .A2(new_n1184), .A3(new_n1186), .ZN(new_n1187));
  INV_X1    g0987(.A(new_n788), .ZN(new_n1188));
  OAI21_X1  g0988(.A(new_n1187), .B1(new_n1188), .B2(new_n1086), .ZN(new_n1189));
  OAI21_X1  g0989(.A(new_n331), .B1(new_n765), .B2(new_n201), .ZN(new_n1190));
  XNOR2_X1  g0990(.A(new_n1190), .B(KEYINPUT122), .ZN(new_n1191));
  NOR2_X1   g0991(.A1(new_n775), .A2(new_n317), .ZN(new_n1192));
  XNOR2_X1  g0992(.A(new_n1192), .B(KEYINPUT53), .ZN(new_n1193));
  NAND2_X1  g0993(.A1(new_n1191), .A2(new_n1193), .ZN(new_n1194));
  OAI21_X1  g0994(.A(new_n1180), .B1(new_n1189), .B2(new_n1194), .ZN(new_n1195));
  AOI21_X1  g0995(.A(new_n1175), .B1(new_n800), .B2(new_n1195), .ZN(new_n1196));
  AOI22_X1  g0996(.A1(new_n1165), .A2(new_n999), .B1(new_n1173), .B2(new_n1196), .ZN(new_n1197));
  NAND2_X1  g0997(.A1(new_n1172), .A2(new_n1197), .ZN(G378));
  INV_X1    g0998(.A(KEYINPUT57), .ZN(new_n1199));
  AOI21_X1  g0999(.A(new_n1157), .B1(new_n1165), .B2(new_n1170), .ZN(new_n1200));
  INV_X1    g1000(.A(KEYINPUT123), .ZN(new_n1201));
  AND3_X1   g1001(.A1(new_n342), .A2(KEYINPUT87), .A3(new_n344), .ZN(new_n1202));
  AOI21_X1  g1002(.A(KEYINPUT87), .B1(new_n342), .B2(new_n344), .ZN(new_n1203));
  OAI21_X1  g1003(.A(new_n350), .B1(new_n1202), .B2(new_n1203), .ZN(new_n1204));
  XNOR2_X1  g1004(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1205));
  NAND2_X1  g1005(.A1(new_n1204), .A2(new_n1205), .ZN(new_n1206));
  INV_X1    g1006(.A(new_n1205), .ZN(new_n1207));
  NAND3_X1  g1007(.A1(new_n669), .A2(new_n350), .A3(new_n1207), .ZN(new_n1208));
  NAND2_X1  g1008(.A1(new_n322), .A2(new_n889), .ZN(new_n1209));
  INV_X1    g1009(.A(new_n1209), .ZN(new_n1210));
  AND3_X1   g1010(.A1(new_n1206), .A2(new_n1208), .A3(new_n1210), .ZN(new_n1211));
  AOI21_X1  g1011(.A(new_n1210), .B1(new_n1206), .B2(new_n1208), .ZN(new_n1212));
  OAI21_X1  g1012(.A(new_n1201), .B1(new_n1211), .B2(new_n1212), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(new_n1206), .A2(new_n1208), .ZN(new_n1214));
  NAND2_X1  g1014(.A1(new_n1214), .A2(new_n1209), .ZN(new_n1215));
  NAND3_X1  g1015(.A1(new_n1206), .A2(new_n1208), .A3(new_n1210), .ZN(new_n1216));
  NAND3_X1  g1016(.A1(new_n1215), .A2(KEYINPUT123), .A3(new_n1216), .ZN(new_n1217));
  NAND2_X1  g1017(.A1(new_n1213), .A2(new_n1217), .ZN(new_n1218));
  INV_X1    g1018(.A(new_n885), .ZN(new_n1219));
  AOI21_X1  g1019(.A(new_n672), .B1(new_n1219), .B2(new_n929), .ZN(new_n1220));
  OAI211_X1 g1020(.A(new_n1218), .B(new_n1220), .C1(new_n917), .C2(KEYINPUT40), .ZN(new_n1221));
  OAI21_X1  g1021(.A(G330), .B1(new_n930), .B2(new_n885), .ZN(new_n1222));
  NAND2_X1  g1022(.A1(new_n951), .A2(new_n952), .ZN(new_n1223));
  NAND2_X1  g1023(.A1(new_n1223), .A2(new_n886), .ZN(new_n1224));
  AOI21_X1  g1024(.A(KEYINPUT106), .B1(new_n1224), .B2(new_n909), .ZN(new_n1225));
  INV_X1    g1025(.A(new_n916), .ZN(new_n1226));
  OAI21_X1  g1026(.A(new_n1219), .B1(new_n1225), .B2(new_n1226), .ZN(new_n1227));
  AOI21_X1  g1027(.A(new_n1222), .B1(new_n1227), .B2(new_n918), .ZN(new_n1228));
  NOR2_X1   g1028(.A1(new_n1211), .A2(new_n1212), .ZN(new_n1229));
  INV_X1    g1029(.A(new_n1229), .ZN(new_n1230));
  OAI21_X1  g1030(.A(new_n1221), .B1(new_n1228), .B2(new_n1230), .ZN(new_n1231));
  INV_X1    g1031(.A(new_n961), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(new_n1231), .A2(new_n1232), .ZN(new_n1233));
  OAI21_X1  g1033(.A(new_n1220), .B1(new_n917), .B2(KEYINPUT40), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n1234), .A2(new_n1229), .ZN(new_n1235));
  NAND3_X1  g1035(.A1(new_n1235), .A2(new_n961), .A3(new_n1221), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n1233), .A2(new_n1236), .ZN(new_n1237));
  OAI21_X1  g1037(.A(new_n1199), .B1(new_n1200), .B2(new_n1237), .ZN(new_n1238));
  AND3_X1   g1038(.A1(new_n1235), .A2(new_n961), .A3(new_n1221), .ZN(new_n1239));
  AOI21_X1  g1039(.A(new_n961), .B1(new_n1235), .B2(new_n1221), .ZN(new_n1240));
  NOR2_X1   g1040(.A1(new_n1239), .A2(new_n1240), .ZN(new_n1241));
  OAI21_X1  g1041(.A(new_n1158), .B1(new_n1144), .B2(new_n1159), .ZN(new_n1242));
  NAND3_X1  g1042(.A1(new_n1241), .A2(new_n1242), .A3(KEYINPUT57), .ZN(new_n1243));
  NAND3_X1  g1043(.A1(new_n1238), .A2(new_n705), .A3(new_n1243), .ZN(new_n1244));
  NAND3_X1  g1044(.A1(new_n1213), .A2(new_n1217), .A3(new_n811), .ZN(new_n1245));
  OAI21_X1  g1045(.A(new_n758), .B1(new_n202), .B2(new_n848), .ZN(new_n1246));
  NOR2_X1   g1046(.A1(new_n331), .A2(G41), .ZN(new_n1247));
  AOI211_X1 g1047(.A(G50), .B(new_n1247), .C1(new_n258), .C2(new_n272), .ZN(new_n1248));
  OAI221_X1 g1048(.A(new_n1247), .B1(new_n219), .B2(new_n775), .C1(new_n259), .C2(new_n780), .ZN(new_n1249));
  AOI21_X1  g1049(.A(new_n1249), .B1(G116), .B2(new_n854), .ZN(new_n1250));
  NOR2_X1   g1050(.A1(new_n765), .A2(new_n225), .ZN(new_n1251));
  OAI22_X1  g1051(.A1(new_n769), .A2(new_n414), .B1(new_n771), .B2(new_n762), .ZN(new_n1252));
  AOI211_X1 g1052(.A(new_n1251), .B(new_n1252), .C1(new_n424), .C2(new_n851), .ZN(new_n1253));
  NAND3_X1  g1053(.A1(new_n1250), .A2(new_n977), .A3(new_n1253), .ZN(new_n1254));
  INV_X1    g1054(.A(KEYINPUT58), .ZN(new_n1255));
  AOI21_X1  g1055(.A(new_n1248), .B1(new_n1254), .B2(new_n1255), .ZN(new_n1256));
  OAI22_X1  g1056(.A1(new_n1181), .A2(new_n769), .B1(new_n775), .B2(new_n1185), .ZN(new_n1257));
  AOI21_X1  g1057(.A(new_n1257), .B1(G137), .B2(new_n851), .ZN(new_n1258));
  AOI22_X1  g1058(.A1(new_n781), .A2(G132), .B1(new_n854), .B2(G125), .ZN(new_n1259));
  OAI211_X1 g1059(.A(new_n1258), .B(new_n1259), .C1(new_n1188), .C2(new_n317), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(new_n1260), .A2(KEYINPUT59), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(new_n794), .A2(G159), .ZN(new_n1262));
  AOI211_X1 g1062(.A(G33), .B(G41), .C1(new_n772), .C2(G124), .ZN(new_n1263));
  NAND3_X1  g1063(.A1(new_n1261), .A2(new_n1262), .A3(new_n1263), .ZN(new_n1264));
  NOR2_X1   g1064(.A1(new_n1260), .A2(KEYINPUT59), .ZN(new_n1265));
  OAI221_X1 g1065(.A(new_n1256), .B1(new_n1255), .B2(new_n1254), .C1(new_n1264), .C2(new_n1265), .ZN(new_n1266));
  AOI21_X1  g1066(.A(new_n1246), .B1(new_n1266), .B2(new_n800), .ZN(new_n1267));
  AOI22_X1  g1067(.A1(new_n1241), .A2(new_n999), .B1(new_n1245), .B2(new_n1267), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1244), .A2(new_n1268), .ZN(G375));
  OAI211_X1 g1069(.A(new_n1157), .B(new_n1146), .C1(new_n1152), .C2(new_n1153), .ZN(new_n1270));
  NAND3_X1  g1070(.A1(new_n1159), .A2(new_n1034), .A3(new_n1270), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(new_n944), .A2(new_n811), .ZN(new_n1272));
  OAI21_X1  g1072(.A(new_n758), .B1(G68), .B2(new_n848), .ZN(new_n1273));
  OAI221_X1 g1073(.A(new_n334), .B1(new_n765), .B2(new_n219), .C1(new_n784), .C2(new_n761), .ZN(new_n1274));
  AOI21_X1  g1074(.A(new_n1274), .B1(G116), .B2(new_n781), .ZN(new_n1275));
  AOI22_X1  g1075(.A1(G283), .A2(new_n770), .B1(new_n851), .B2(G107), .ZN(new_n1276));
  AOI22_X1  g1076(.A1(G97), .A2(new_n793), .B1(new_n772), .B2(G303), .ZN(new_n1277));
  NAND4_X1  g1077(.A1(new_n1275), .A2(new_n1049), .A3(new_n1276), .A4(new_n1277), .ZN(new_n1278));
  NAND2_X1  g1078(.A1(new_n854), .A2(G132), .ZN(new_n1279));
  XNOR2_X1  g1079(.A(new_n1279), .B(KEYINPUT124), .ZN(new_n1280));
  OAI22_X1  g1080(.A1(new_n979), .A2(new_n769), .B1(new_n771), .B2(new_n1181), .ZN(new_n1281));
  OAI22_X1  g1081(.A1(new_n775), .A2(new_n1086), .B1(new_n777), .B2(new_n317), .ZN(new_n1282));
  NOR2_X1   g1082(.A1(new_n1281), .A2(new_n1282), .ZN(new_n1283));
  NOR2_X1   g1083(.A1(new_n780), .A2(new_n1185), .ZN(new_n1284));
  NOR3_X1   g1084(.A1(new_n1284), .A2(new_n1251), .A3(new_n334), .ZN(new_n1285));
  OAI211_X1 g1085(.A(new_n1283), .B(new_n1285), .C1(new_n1188), .C2(new_n293), .ZN(new_n1286));
  OAI21_X1  g1086(.A(new_n1278), .B1(new_n1280), .B2(new_n1286), .ZN(new_n1287));
  AOI21_X1  g1087(.A(new_n1273), .B1(new_n1287), .B2(new_n800), .ZN(new_n1288));
  AOI22_X1  g1088(.A1(new_n1154), .A2(new_n999), .B1(new_n1272), .B2(new_n1288), .ZN(new_n1289));
  NAND2_X1  g1089(.A1(new_n1271), .A2(new_n1289), .ZN(G381));
  OR4_X1    g1090(.A1(G396), .A2(G381), .A3(G384), .A4(G393), .ZN(new_n1291));
  OAI211_X1 g1091(.A(new_n998), .B(new_n1116), .C1(new_n1035), .C2(new_n1045), .ZN(new_n1292));
  OR4_X1    g1092(.A1(G378), .A2(G375), .A3(new_n1291), .A4(new_n1292), .ZN(G407));
  NAND2_X1  g1093(.A1(new_n1245), .A2(new_n1267), .ZN(new_n1294));
  OAI21_X1  g1094(.A(new_n1294), .B1(new_n1237), .B2(new_n1111), .ZN(new_n1295));
  NAND2_X1  g1095(.A1(new_n1241), .A2(new_n1242), .ZN(new_n1296));
  AOI21_X1  g1096(.A(new_n706), .B1(new_n1296), .B2(new_n1199), .ZN(new_n1297));
  AOI21_X1  g1097(.A(new_n1295), .B1(new_n1297), .B2(new_n1243), .ZN(new_n1298));
  INV_X1    g1098(.A(G378), .ZN(new_n1299));
  NAND2_X1  g1099(.A1(new_n680), .A2(G213), .ZN(new_n1300));
  INV_X1    g1100(.A(new_n1300), .ZN(new_n1301));
  NAND3_X1  g1101(.A1(new_n1298), .A2(new_n1299), .A3(new_n1301), .ZN(new_n1302));
  NAND3_X1  g1102(.A1(G407), .A2(G213), .A3(new_n1302), .ZN(G409));
  NAND3_X1  g1103(.A1(new_n1244), .A2(G378), .A3(new_n1268), .ZN(new_n1304));
  NAND3_X1  g1104(.A1(new_n1241), .A2(new_n1242), .A3(new_n1034), .ZN(new_n1305));
  NAND2_X1  g1105(.A1(new_n1268), .A2(new_n1305), .ZN(new_n1306));
  NAND2_X1  g1106(.A1(new_n1306), .A2(new_n1299), .ZN(new_n1307));
  NAND2_X1  g1107(.A1(new_n1304), .A2(new_n1307), .ZN(new_n1308));
  INV_X1    g1108(.A(KEYINPUT125), .ZN(new_n1309));
  INV_X1    g1109(.A(KEYINPUT60), .ZN(new_n1310));
  NAND2_X1  g1110(.A1(new_n1270), .A2(new_n1310), .ZN(new_n1311));
  NAND4_X1  g1111(.A1(new_n1169), .A2(KEYINPUT60), .A3(new_n1157), .A4(new_n1146), .ZN(new_n1312));
  NAND4_X1  g1112(.A1(new_n1311), .A2(new_n1159), .A3(new_n1312), .A4(new_n705), .ZN(new_n1313));
  AND3_X1   g1113(.A1(new_n1313), .A2(G384), .A3(new_n1289), .ZN(new_n1314));
  AOI21_X1  g1114(.A(G384), .B1(new_n1313), .B2(new_n1289), .ZN(new_n1315));
  OAI21_X1  g1115(.A(new_n1309), .B1(new_n1314), .B2(new_n1315), .ZN(new_n1316));
  NAND2_X1  g1116(.A1(new_n1313), .A2(new_n1289), .ZN(new_n1317));
  INV_X1    g1117(.A(G384), .ZN(new_n1318));
  NAND2_X1  g1118(.A1(new_n1317), .A2(new_n1318), .ZN(new_n1319));
  NAND3_X1  g1119(.A1(new_n1313), .A2(G384), .A3(new_n1289), .ZN(new_n1320));
  NAND3_X1  g1120(.A1(new_n1319), .A2(KEYINPUT125), .A3(new_n1320), .ZN(new_n1321));
  NAND2_X1  g1121(.A1(new_n1316), .A2(new_n1321), .ZN(new_n1322));
  NAND3_X1  g1122(.A1(new_n1308), .A2(new_n1300), .A3(new_n1322), .ZN(new_n1323));
  NAND2_X1  g1123(.A1(new_n1323), .A2(KEYINPUT62), .ZN(new_n1324));
  INV_X1    g1124(.A(KEYINPUT61), .ZN(new_n1325));
  NAND2_X1  g1125(.A1(new_n1301), .A2(G2897), .ZN(new_n1326));
  AOI21_X1  g1126(.A(new_n1326), .B1(new_n1319), .B2(new_n1320), .ZN(new_n1327));
  AOI21_X1  g1127(.A(new_n1327), .B1(new_n1322), .B2(new_n1326), .ZN(new_n1328));
  AOI21_X1  g1128(.A(G378), .B1(new_n1268), .B2(new_n1305), .ZN(new_n1329));
  AOI21_X1  g1129(.A(new_n1329), .B1(new_n1298), .B2(G378), .ZN(new_n1330));
  OAI21_X1  g1130(.A(new_n1328), .B1(new_n1330), .B2(new_n1301), .ZN(new_n1331));
  AOI21_X1  g1131(.A(new_n1301), .B1(new_n1304), .B2(new_n1307), .ZN(new_n1332));
  INV_X1    g1132(.A(KEYINPUT62), .ZN(new_n1333));
  NAND3_X1  g1133(.A1(new_n1332), .A2(new_n1333), .A3(new_n1322), .ZN(new_n1334));
  NAND4_X1  g1134(.A1(new_n1324), .A2(new_n1325), .A3(new_n1331), .A4(new_n1334), .ZN(new_n1335));
  XNOR2_X1  g1135(.A(G393), .B(new_n823), .ZN(new_n1336));
  AOI21_X1  g1136(.A(new_n1033), .B1(new_n1114), .B2(new_n753), .ZN(new_n1337));
  OAI21_X1  g1137(.A(new_n1044), .B1(new_n1337), .B2(new_n999), .ZN(new_n1338));
  AOI21_X1  g1138(.A(new_n1116), .B1(new_n1338), .B2(new_n998), .ZN(new_n1339));
  NAND2_X1  g1139(.A1(new_n1292), .A2(KEYINPUT126), .ZN(new_n1340));
  OAI21_X1  g1140(.A(new_n1336), .B1(new_n1339), .B2(new_n1340), .ZN(new_n1341));
  NAND2_X1  g1141(.A1(G387), .A2(G390), .ZN(new_n1342));
  INV_X1    g1142(.A(new_n1336), .ZN(new_n1343));
  NAND4_X1  g1143(.A1(new_n1342), .A2(new_n1343), .A3(KEYINPUT126), .A4(new_n1292), .ZN(new_n1344));
  AND3_X1   g1144(.A1(new_n1341), .A2(KEYINPUT127), .A3(new_n1344), .ZN(new_n1345));
  AOI21_X1  g1145(.A(KEYINPUT127), .B1(new_n1341), .B2(new_n1344), .ZN(new_n1346));
  NOR2_X1   g1146(.A1(new_n1345), .A2(new_n1346), .ZN(new_n1347));
  NAND2_X1  g1147(.A1(new_n1335), .A2(new_n1347), .ZN(new_n1348));
  INV_X1    g1148(.A(new_n1332), .ZN(new_n1349));
  AOI21_X1  g1149(.A(KEYINPUT61), .B1(new_n1349), .B2(new_n1328), .ZN(new_n1350));
  AND2_X1   g1150(.A1(new_n1341), .A2(new_n1344), .ZN(new_n1351));
  NOR2_X1   g1151(.A1(new_n1323), .A2(KEYINPUT63), .ZN(new_n1352));
  INV_X1    g1152(.A(KEYINPUT63), .ZN(new_n1353));
  AOI21_X1  g1153(.A(new_n1353), .B1(new_n1332), .B2(new_n1322), .ZN(new_n1354));
  OAI211_X1 g1154(.A(new_n1350), .B(new_n1351), .C1(new_n1352), .C2(new_n1354), .ZN(new_n1355));
  NAND2_X1  g1155(.A1(new_n1348), .A2(new_n1355), .ZN(G405));
  XNOR2_X1  g1156(.A(G375), .B(G378), .ZN(new_n1357));
  NAND2_X1  g1157(.A1(new_n1319), .A2(new_n1320), .ZN(new_n1358));
  NAND2_X1  g1158(.A1(new_n1357), .A2(new_n1358), .ZN(new_n1359));
  INV_X1    g1159(.A(new_n1322), .ZN(new_n1360));
  OAI21_X1  g1160(.A(new_n1359), .B1(new_n1360), .B2(new_n1357), .ZN(new_n1361));
  NAND2_X1  g1161(.A1(new_n1361), .A2(new_n1347), .ZN(new_n1362));
  OAI221_X1 g1162(.A(new_n1359), .B1(new_n1360), .B2(new_n1357), .C1(new_n1345), .C2(new_n1346), .ZN(new_n1363));
  NAND2_X1  g1163(.A1(new_n1362), .A2(new_n1363), .ZN(G402));
endmodule


