//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 0 0 1 1 0 1 0 0 0 0 0 0 0 1 0 0 0 1 1 1 1 0 0 0 0 1 1 0 0 0 1 1 0 1 1 1 1 0 1 0 1 0 1 1 0 0 0 0 1 0 0 1 1 1 1 1 0 1 1 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:19:47 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n683, new_n684, new_n685,
    new_n686, new_n687, new_n688, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n698, new_n699, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n728, new_n729, new_n730, new_n731,
    new_n732, new_n733, new_n734, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n780, new_n781, new_n782, new_n783, new_n785,
    new_n786, new_n787, new_n789, new_n791, new_n792, new_n793, new_n794,
    new_n795, new_n796, new_n797, new_n798, new_n799, new_n800, new_n801,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n814, new_n815, new_n816, new_n817,
    new_n818, new_n819, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n870, new_n871, new_n873, new_n874, new_n875, new_n877, new_n878,
    new_n879, new_n880, new_n881, new_n882, new_n883, new_n884, new_n885,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n936, new_n937,
    new_n939, new_n940, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n948, new_n949, new_n950, new_n952, new_n953, new_n954, new_n955,
    new_n956, new_n957, new_n959, new_n960, new_n961, new_n963, new_n964,
    new_n965, new_n966, new_n967, new_n968, new_n969, new_n970, new_n971,
    new_n972, new_n974, new_n975, new_n976, new_n977, new_n978, new_n980,
    new_n981, new_n982, new_n983, new_n984, new_n986, new_n987, new_n988;
  INV_X1    g000(.A(KEYINPUT35), .ZN(new_n202));
  INV_X1    g001(.A(KEYINPUT86), .ZN(new_n203));
  NAND2_X1  g002(.A1(G155gat), .A2(G162gat), .ZN(new_n204));
  INV_X1    g003(.A(G155gat), .ZN(new_n205));
  INV_X1    g004(.A(G162gat), .ZN(new_n206));
  NAND2_X1  g005(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  XNOR2_X1  g006(.A(G141gat), .B(G148gat), .ZN(new_n208));
  OAI211_X1 g007(.A(new_n204), .B(new_n207), .C1(new_n208), .C2(KEYINPUT2), .ZN(new_n209));
  AND2_X1   g008(.A1(G155gat), .A2(G162gat), .ZN(new_n210));
  NOR2_X1   g009(.A1(G155gat), .A2(G162gat), .ZN(new_n211));
  OAI21_X1  g010(.A(KEYINPUT80), .B1(new_n210), .B2(new_n211), .ZN(new_n212));
  INV_X1    g011(.A(KEYINPUT80), .ZN(new_n213));
  NAND3_X1  g012(.A1(new_n207), .A2(new_n213), .A3(new_n204), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n204), .A2(KEYINPUT2), .ZN(new_n215));
  NAND3_X1  g014(.A1(new_n212), .A2(new_n214), .A3(new_n215), .ZN(new_n216));
  INV_X1    g015(.A(G141gat), .ZN(new_n217));
  NAND2_X1  g016(.A1(new_n217), .A2(G148gat), .ZN(new_n218));
  INV_X1    g017(.A(new_n218), .ZN(new_n219));
  AND2_X1   g018(.A1(KEYINPUT79), .A2(G148gat), .ZN(new_n220));
  NOR2_X1   g019(.A1(KEYINPUT79), .A2(G148gat), .ZN(new_n221));
  NOR2_X1   g020(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  AOI21_X1  g021(.A(new_n219), .B1(new_n222), .B2(G141gat), .ZN(new_n223));
  OAI21_X1  g022(.A(new_n209), .B1(new_n216), .B2(new_n223), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n224), .A2(KEYINPUT81), .ZN(new_n225));
  INV_X1    g024(.A(KEYINPUT81), .ZN(new_n226));
  OAI211_X1 g025(.A(new_n226), .B(new_n209), .C1(new_n216), .C2(new_n223), .ZN(new_n227));
  AND2_X1   g026(.A1(new_n225), .A2(new_n227), .ZN(new_n228));
  INV_X1    g027(.A(KEYINPUT3), .ZN(new_n229));
  NAND2_X1  g028(.A1(G211gat), .A2(G218gat), .ZN(new_n230));
  INV_X1    g029(.A(KEYINPUT22), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n230), .A2(new_n231), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n232), .A2(KEYINPUT76), .ZN(new_n233));
  INV_X1    g032(.A(KEYINPUT76), .ZN(new_n234));
  NAND3_X1  g033(.A1(new_n230), .A2(new_n234), .A3(new_n231), .ZN(new_n235));
  XNOR2_X1  g034(.A(G197gat), .B(G204gat), .ZN(new_n236));
  NAND3_X1  g035(.A1(new_n233), .A2(new_n235), .A3(new_n236), .ZN(new_n237));
  XNOR2_X1  g036(.A(G211gat), .B(G218gat), .ZN(new_n238));
  INV_X1    g037(.A(new_n238), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n237), .A2(new_n239), .ZN(new_n240));
  NAND4_X1  g039(.A1(new_n233), .A2(new_n238), .A3(new_n236), .A4(new_n235), .ZN(new_n241));
  AOI21_X1  g040(.A(KEYINPUT29), .B1(new_n240), .B2(new_n241), .ZN(new_n242));
  OAI21_X1  g041(.A(new_n229), .B1(new_n242), .B2(KEYINPUT84), .ZN(new_n243));
  INV_X1    g042(.A(KEYINPUT84), .ZN(new_n244));
  AOI211_X1 g043(.A(new_n244), .B(KEYINPUT29), .C1(new_n240), .C2(new_n241), .ZN(new_n245));
  OAI21_X1  g044(.A(new_n228), .B1(new_n243), .B2(new_n245), .ZN(new_n246));
  NAND2_X1  g045(.A1(G228gat), .A2(G233gat), .ZN(new_n247));
  AND3_X1   g046(.A1(new_n240), .A2(KEYINPUT77), .A3(new_n241), .ZN(new_n248));
  AOI21_X1  g047(.A(KEYINPUT77), .B1(new_n240), .B2(new_n241), .ZN(new_n249));
  NOR2_X1   g048(.A1(new_n248), .A2(new_n249), .ZN(new_n250));
  OAI211_X1 g049(.A(new_n229), .B(new_n209), .C1(new_n216), .C2(new_n223), .ZN(new_n251));
  INV_X1    g050(.A(KEYINPUT29), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n251), .A2(new_n252), .ZN(new_n253));
  AOI21_X1  g052(.A(new_n247), .B1(new_n250), .B2(new_n253), .ZN(new_n254));
  NAND2_X1  g053(.A1(new_n246), .A2(new_n254), .ZN(new_n255));
  INV_X1    g054(.A(new_n249), .ZN(new_n256));
  NAND3_X1  g055(.A1(new_n240), .A2(KEYINPUT77), .A3(new_n241), .ZN(new_n257));
  NAND3_X1  g056(.A1(new_n256), .A2(new_n253), .A3(new_n257), .ZN(new_n258));
  OAI21_X1  g057(.A(new_n224), .B1(new_n242), .B2(KEYINPUT3), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n260), .A2(new_n247), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n255), .A2(new_n261), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n262), .A2(G22gat), .ZN(new_n263));
  XNOR2_X1  g062(.A(G78gat), .B(G106gat), .ZN(new_n264));
  XNOR2_X1  g063(.A(KEYINPUT31), .B(G50gat), .ZN(new_n265));
  XOR2_X1   g064(.A(new_n264), .B(new_n265), .Z(new_n266));
  INV_X1    g065(.A(new_n266), .ZN(new_n267));
  INV_X1    g066(.A(G22gat), .ZN(new_n268));
  NAND3_X1  g067(.A1(new_n255), .A2(new_n261), .A3(new_n268), .ZN(new_n269));
  NAND3_X1  g068(.A1(new_n263), .A2(new_n267), .A3(new_n269), .ZN(new_n270));
  NAND3_X1  g069(.A1(new_n263), .A2(KEYINPUT85), .A3(new_n269), .ZN(new_n271));
  AOI21_X1  g070(.A(new_n268), .B1(new_n255), .B2(new_n261), .ZN(new_n272));
  INV_X1    g071(.A(KEYINPUT85), .ZN(new_n273));
  AOI21_X1  g072(.A(new_n267), .B1(new_n272), .B2(new_n273), .ZN(new_n274));
  AOI22_X1  g073(.A1(new_n203), .A2(new_n270), .B1(new_n271), .B2(new_n274), .ZN(new_n275));
  OR2_X1    g074(.A1(new_n270), .A2(new_n203), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  INV_X1    g076(.A(G227gat), .ZN(new_n278));
  INV_X1    g077(.A(G233gat), .ZN(new_n279));
  NOR2_X1   g078(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  XNOR2_X1  g079(.A(new_n280), .B(KEYINPUT64), .ZN(new_n281));
  NAND2_X1  g080(.A1(G169gat), .A2(G176gat), .ZN(new_n282));
  INV_X1    g081(.A(G169gat), .ZN(new_n283));
  INV_X1    g082(.A(G176gat), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n285), .A2(KEYINPUT26), .ZN(new_n286));
  NAND3_X1  g085(.A1(new_n283), .A2(new_n284), .A3(KEYINPUT66), .ZN(new_n287));
  INV_X1    g086(.A(KEYINPUT66), .ZN(new_n288));
  OAI21_X1  g087(.A(new_n288), .B1(G169gat), .B2(G176gat), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n287), .A2(new_n289), .ZN(new_n290));
  OAI211_X1 g089(.A(new_n282), .B(new_n286), .C1(new_n290), .C2(KEYINPUT26), .ZN(new_n291));
  NAND2_X1  g090(.A1(G183gat), .A2(G190gat), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  INV_X1    g092(.A(KEYINPUT28), .ZN(new_n294));
  INV_X1    g093(.A(G183gat), .ZN(new_n295));
  OR3_X1    g094(.A1(new_n295), .A2(KEYINPUT70), .A3(KEYINPUT27), .ZN(new_n296));
  INV_X1    g095(.A(G190gat), .ZN(new_n297));
  OAI21_X1  g096(.A(KEYINPUT70), .B1(new_n295), .B2(KEYINPUT27), .ZN(new_n298));
  NAND3_X1  g097(.A1(new_n296), .A2(new_n297), .A3(new_n298), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n295), .A2(KEYINPUT67), .ZN(new_n300));
  INV_X1    g099(.A(KEYINPUT67), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n301), .A2(G183gat), .ZN(new_n302));
  AND3_X1   g101(.A1(new_n300), .A2(new_n302), .A3(KEYINPUT27), .ZN(new_n303));
  OAI21_X1  g102(.A(new_n294), .B1(new_n299), .B2(new_n303), .ZN(new_n304));
  XNOR2_X1  g103(.A(KEYINPUT27), .B(G183gat), .ZN(new_n305));
  NOR2_X1   g104(.A1(new_n294), .A2(G190gat), .ZN(new_n306));
  AND3_X1   g105(.A1(new_n305), .A2(KEYINPUT71), .A3(new_n306), .ZN(new_n307));
  AOI21_X1  g106(.A(KEYINPUT71), .B1(new_n305), .B2(new_n306), .ZN(new_n308));
  NOR2_X1   g107(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  AOI21_X1  g108(.A(new_n293), .B1(new_n304), .B2(new_n309), .ZN(new_n310));
  NAND3_X1  g109(.A1(new_n300), .A2(new_n302), .A3(new_n297), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n292), .A2(KEYINPUT24), .ZN(new_n312));
  INV_X1    g111(.A(KEYINPUT24), .ZN(new_n313));
  NAND3_X1  g112(.A1(new_n313), .A2(G183gat), .A3(G190gat), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n312), .A2(new_n314), .ZN(new_n315));
  AND3_X1   g114(.A1(new_n311), .A2(new_n315), .A3(KEYINPUT68), .ZN(new_n316));
  AOI21_X1  g115(.A(KEYINPUT68), .B1(new_n311), .B2(new_n315), .ZN(new_n317));
  INV_X1    g116(.A(KEYINPUT25), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n282), .A2(KEYINPUT23), .ZN(new_n319));
  AOI21_X1  g118(.A(new_n318), .B1(new_n319), .B2(new_n285), .ZN(new_n320));
  NAND3_X1  g119(.A1(new_n287), .A2(new_n289), .A3(KEYINPUT23), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n320), .A2(new_n321), .ZN(new_n322));
  NOR3_X1   g121(.A1(new_n316), .A2(new_n317), .A3(new_n322), .ZN(new_n323));
  NOR2_X1   g122(.A1(G169gat), .A2(G176gat), .ZN(new_n324));
  AOI21_X1  g123(.A(new_n324), .B1(KEYINPUT23), .B2(new_n282), .ZN(new_n325));
  OR2_X1    g124(.A1(KEYINPUT65), .A2(G176gat), .ZN(new_n326));
  NAND2_X1  g125(.A1(KEYINPUT65), .A2(G176gat), .ZN(new_n327));
  AND2_X1   g126(.A1(new_n326), .A2(new_n327), .ZN(new_n328));
  AND2_X1   g127(.A1(new_n283), .A2(KEYINPUT23), .ZN(new_n329));
  AOI21_X1  g128(.A(new_n325), .B1(new_n328), .B2(new_n329), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n295), .A2(new_n297), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n315), .A2(new_n331), .ZN(new_n332));
  AOI21_X1  g131(.A(KEYINPUT25), .B1(new_n330), .B2(new_n332), .ZN(new_n333));
  OAI21_X1  g132(.A(KEYINPUT69), .B1(new_n323), .B2(new_n333), .ZN(new_n334));
  NAND2_X1  g133(.A1(new_n311), .A2(new_n315), .ZN(new_n335));
  INV_X1    g134(.A(KEYINPUT68), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n335), .A2(new_n336), .ZN(new_n337));
  AND2_X1   g136(.A1(new_n320), .A2(new_n321), .ZN(new_n338));
  NAND3_X1  g137(.A1(new_n311), .A2(new_n315), .A3(KEYINPUT68), .ZN(new_n339));
  NAND3_X1  g138(.A1(new_n337), .A2(new_n338), .A3(new_n339), .ZN(new_n340));
  INV_X1    g139(.A(new_n332), .ZN(new_n341));
  NAND3_X1  g140(.A1(new_n329), .A2(new_n326), .A3(new_n327), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n319), .A2(new_n285), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n342), .A2(new_n343), .ZN(new_n344));
  OAI21_X1  g143(.A(new_n318), .B1(new_n341), .B2(new_n344), .ZN(new_n345));
  INV_X1    g144(.A(KEYINPUT69), .ZN(new_n346));
  NAND3_X1  g145(.A1(new_n340), .A2(new_n345), .A3(new_n346), .ZN(new_n347));
  AOI21_X1  g146(.A(new_n310), .B1(new_n334), .B2(new_n347), .ZN(new_n348));
  INV_X1    g147(.A(G120gat), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n349), .A2(G113gat), .ZN(new_n350));
  INV_X1    g149(.A(G113gat), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n351), .A2(G120gat), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n350), .A2(new_n352), .ZN(new_n353));
  INV_X1    g152(.A(KEYINPUT1), .ZN(new_n354));
  XNOR2_X1  g153(.A(G127gat), .B(G134gat), .ZN(new_n355));
  OAI211_X1 g154(.A(new_n353), .B(new_n354), .C1(new_n355), .C2(KEYINPUT72), .ZN(new_n356));
  INV_X1    g155(.A(G127gat), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n357), .A2(G134gat), .ZN(new_n358));
  INV_X1    g157(.A(G134gat), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n359), .A2(G127gat), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n358), .A2(new_n360), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n354), .A2(KEYINPUT72), .ZN(new_n362));
  XNOR2_X1  g161(.A(G113gat), .B(G120gat), .ZN(new_n363));
  OAI211_X1 g162(.A(new_n361), .B(new_n362), .C1(new_n363), .C2(KEYINPUT1), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n356), .A2(new_n364), .ZN(new_n365));
  INV_X1    g164(.A(KEYINPUT73), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n365), .A2(new_n366), .ZN(new_n367));
  NAND3_X1  g166(.A1(new_n356), .A2(new_n364), .A3(KEYINPUT73), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  INV_X1    g168(.A(new_n369), .ZN(new_n370));
  NOR2_X1   g169(.A1(new_n348), .A2(new_n370), .ZN(new_n371));
  AOI211_X1 g170(.A(new_n369), .B(new_n310), .C1(new_n334), .C2(new_n347), .ZN(new_n372));
  OAI21_X1  g171(.A(new_n281), .B1(new_n371), .B2(new_n372), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n373), .A2(KEYINPUT32), .ZN(new_n374));
  INV_X1    g173(.A(KEYINPUT33), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n373), .A2(new_n375), .ZN(new_n376));
  XNOR2_X1  g175(.A(KEYINPUT74), .B(G71gat), .ZN(new_n377));
  XNOR2_X1  g176(.A(new_n377), .B(G99gat), .ZN(new_n378));
  XOR2_X1   g177(.A(G15gat), .B(G43gat), .Z(new_n379));
  XOR2_X1   g178(.A(new_n378), .B(new_n379), .Z(new_n380));
  NAND3_X1  g179(.A1(new_n374), .A2(new_n376), .A3(new_n380), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n309), .A2(new_n304), .ZN(new_n382));
  NAND3_X1  g181(.A1(new_n382), .A2(new_n292), .A3(new_n291), .ZN(new_n383));
  AND3_X1   g182(.A1(new_n340), .A2(new_n346), .A3(new_n345), .ZN(new_n384));
  AOI21_X1  g183(.A(new_n346), .B1(new_n340), .B2(new_n345), .ZN(new_n385));
  OAI21_X1  g184(.A(new_n383), .B1(new_n384), .B2(new_n385), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n386), .A2(new_n369), .ZN(new_n387));
  OAI211_X1 g186(.A(new_n370), .B(new_n383), .C1(new_n384), .C2(new_n385), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n387), .A2(new_n388), .ZN(new_n389));
  INV_X1    g188(.A(new_n389), .ZN(new_n390));
  NOR2_X1   g189(.A1(new_n281), .A2(KEYINPUT34), .ZN(new_n391));
  OAI211_X1 g190(.A(new_n387), .B(new_n388), .C1(new_n278), .C2(new_n279), .ZN(new_n392));
  AOI22_X1  g191(.A1(new_n390), .A2(new_n391), .B1(new_n392), .B2(KEYINPUT34), .ZN(new_n393));
  INV_X1    g192(.A(new_n380), .ZN(new_n394));
  OAI211_X1 g193(.A(new_n373), .B(KEYINPUT32), .C1(new_n375), .C2(new_n394), .ZN(new_n395));
  NAND3_X1  g194(.A1(new_n381), .A2(new_n393), .A3(new_n395), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n390), .A2(new_n391), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n392), .A2(KEYINPUT34), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n397), .A2(new_n398), .ZN(new_n399));
  INV_X1    g198(.A(new_n281), .ZN(new_n400));
  AOI21_X1  g199(.A(new_n400), .B1(new_n387), .B2(new_n388), .ZN(new_n401));
  OAI21_X1  g200(.A(new_n380), .B1(new_n401), .B2(KEYINPUT33), .ZN(new_n402));
  INV_X1    g201(.A(KEYINPUT32), .ZN(new_n403));
  NOR2_X1   g202(.A1(new_n401), .A2(new_n403), .ZN(new_n404));
  NOR2_X1   g203(.A1(new_n402), .A2(new_n404), .ZN(new_n405));
  AOI221_X4 g204(.A(new_n403), .B1(KEYINPUT33), .B2(new_n380), .C1(new_n389), .C2(new_n281), .ZN(new_n406));
  OAI21_X1  g205(.A(new_n399), .B1(new_n405), .B2(new_n406), .ZN(new_n407));
  NAND3_X1  g206(.A1(new_n277), .A2(new_n396), .A3(new_n407), .ZN(new_n408));
  XNOR2_X1  g207(.A(G1gat), .B(G29gat), .ZN(new_n409));
  XNOR2_X1  g208(.A(new_n409), .B(KEYINPUT0), .ZN(new_n410));
  XNOR2_X1  g209(.A(G57gat), .B(G85gat), .ZN(new_n411));
  XNOR2_X1  g210(.A(new_n410), .B(new_n411), .ZN(new_n412));
  XOR2_X1   g211(.A(KEYINPUT83), .B(KEYINPUT6), .Z(new_n413));
  NOR2_X1   g212(.A1(new_n412), .A2(new_n413), .ZN(new_n414));
  AND2_X1   g213(.A1(new_n412), .A2(new_n413), .ZN(new_n415));
  XNOR2_X1  g214(.A(KEYINPUT82), .B(KEYINPUT5), .ZN(new_n416));
  NAND3_X1  g215(.A1(new_n225), .A2(new_n227), .A3(new_n365), .ZN(new_n417));
  INV_X1    g216(.A(new_n365), .ZN(new_n418));
  XNOR2_X1  g217(.A(KEYINPUT79), .B(G148gat), .ZN(new_n419));
  OAI21_X1  g218(.A(new_n218), .B1(new_n419), .B2(new_n217), .ZN(new_n420));
  NAND4_X1  g219(.A1(new_n420), .A2(new_n214), .A3(new_n215), .A4(new_n212), .ZN(new_n421));
  NAND3_X1  g220(.A1(new_n418), .A2(new_n209), .A3(new_n421), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n417), .A2(new_n422), .ZN(new_n423));
  NAND2_X1  g222(.A1(G225gat), .A2(G233gat), .ZN(new_n424));
  INV_X1    g223(.A(new_n424), .ZN(new_n425));
  AOI21_X1  g224(.A(new_n416), .B1(new_n423), .B2(new_n425), .ZN(new_n426));
  NAND3_X1  g225(.A1(new_n225), .A2(KEYINPUT3), .A3(new_n227), .ZN(new_n427));
  AND2_X1   g226(.A1(new_n251), .A2(new_n365), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n427), .A2(new_n428), .ZN(new_n429));
  INV_X1    g228(.A(KEYINPUT4), .ZN(new_n430));
  AOI21_X1  g229(.A(new_n425), .B1(new_n422), .B2(new_n430), .ZN(new_n431));
  INV_X1    g230(.A(new_n224), .ZN(new_n432));
  NAND4_X1  g231(.A1(new_n432), .A2(new_n367), .A3(KEYINPUT4), .A4(new_n368), .ZN(new_n433));
  NAND3_X1  g232(.A1(new_n429), .A2(new_n431), .A3(new_n433), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n426), .A2(new_n434), .ZN(new_n435));
  NOR3_X1   g234(.A1(new_n224), .A2(new_n365), .A3(new_n430), .ZN(new_n436));
  NAND3_X1  g235(.A1(new_n432), .A2(new_n367), .A3(new_n368), .ZN(new_n437));
  AOI21_X1  g236(.A(new_n436), .B1(new_n437), .B2(new_n430), .ZN(new_n438));
  NAND4_X1  g237(.A1(new_n438), .A2(new_n429), .A3(new_n424), .A4(new_n416), .ZN(new_n439));
  AOI211_X1 g238(.A(new_n414), .B(new_n415), .C1(new_n435), .C2(new_n439), .ZN(new_n440));
  AND4_X1   g239(.A1(new_n435), .A2(new_n439), .A3(new_n412), .A4(new_n413), .ZN(new_n441));
  NOR2_X1   g240(.A1(new_n440), .A2(new_n441), .ZN(new_n442));
  INV_X1    g241(.A(new_n442), .ZN(new_n443));
  XNOR2_X1  g242(.A(G8gat), .B(G36gat), .ZN(new_n444));
  XNOR2_X1  g243(.A(new_n444), .B(KEYINPUT78), .ZN(new_n445));
  XNOR2_X1  g244(.A(G64gat), .B(G92gat), .ZN(new_n446));
  XOR2_X1   g245(.A(new_n445), .B(new_n446), .Z(new_n447));
  AND2_X1   g246(.A1(G226gat), .A2(G233gat), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n340), .A2(new_n345), .ZN(new_n449));
  NAND3_X1  g248(.A1(new_n383), .A2(new_n448), .A3(new_n449), .ZN(new_n450));
  NOR2_X1   g249(.A1(new_n448), .A2(KEYINPUT29), .ZN(new_n451));
  INV_X1    g250(.A(new_n451), .ZN(new_n452));
  OAI211_X1 g251(.A(new_n250), .B(new_n450), .C1(new_n348), .C2(new_n452), .ZN(new_n453));
  INV_X1    g252(.A(new_n453), .ZN(new_n454));
  OAI211_X1 g253(.A(new_n448), .B(new_n383), .C1(new_n384), .C2(new_n385), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n383), .A2(new_n449), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n456), .A2(new_n451), .ZN(new_n457));
  AOI21_X1  g256(.A(new_n250), .B1(new_n455), .B2(new_n457), .ZN(new_n458));
  OAI21_X1  g257(.A(new_n447), .B1(new_n454), .B2(new_n458), .ZN(new_n459));
  INV_X1    g258(.A(new_n447), .ZN(new_n460));
  AOI22_X1  g259(.A1(new_n348), .A2(new_n448), .B1(new_n451), .B2(new_n456), .ZN(new_n461));
  OAI211_X1 g260(.A(new_n453), .B(new_n460), .C1(new_n461), .C2(new_n250), .ZN(new_n462));
  NAND3_X1  g261(.A1(new_n459), .A2(KEYINPUT30), .A3(new_n462), .ZN(new_n463));
  INV_X1    g262(.A(new_n458), .ZN(new_n464));
  INV_X1    g263(.A(KEYINPUT30), .ZN(new_n465));
  NAND4_X1  g264(.A1(new_n464), .A2(new_n465), .A3(new_n460), .A4(new_n453), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n463), .A2(new_n466), .ZN(new_n467));
  INV_X1    g266(.A(KEYINPUT90), .ZN(new_n468));
  NAND3_X1  g267(.A1(new_n443), .A2(new_n467), .A3(new_n468), .ZN(new_n469));
  OAI21_X1  g268(.A(new_n202), .B1(new_n408), .B2(new_n469), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n407), .A2(new_n396), .ZN(new_n471));
  INV_X1    g270(.A(new_n471), .ZN(new_n472));
  INV_X1    g271(.A(new_n469), .ZN(new_n473));
  NAND4_X1  g272(.A1(new_n472), .A2(new_n473), .A3(KEYINPUT35), .A4(new_n277), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n470), .A2(new_n474), .ZN(new_n475));
  INV_X1    g274(.A(KEYINPUT89), .ZN(new_n476));
  INV_X1    g275(.A(KEYINPUT88), .ZN(new_n477));
  INV_X1    g276(.A(KEYINPUT38), .ZN(new_n478));
  INV_X1    g277(.A(new_n250), .ZN(new_n479));
  OAI211_X1 g278(.A(new_n479), .B(new_n450), .C1(new_n348), .C2(new_n452), .ZN(new_n480));
  OAI211_X1 g279(.A(new_n480), .B(KEYINPUT37), .C1(new_n461), .C2(new_n479), .ZN(new_n481));
  INV_X1    g280(.A(KEYINPUT37), .ZN(new_n482));
  OAI211_X1 g281(.A(new_n453), .B(new_n482), .C1(new_n461), .C2(new_n250), .ZN(new_n483));
  AND4_X1   g282(.A1(new_n478), .A2(new_n481), .A3(new_n483), .A4(new_n447), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n435), .A2(new_n439), .ZN(new_n485));
  INV_X1    g284(.A(new_n414), .ZN(new_n486));
  INV_X1    g285(.A(new_n415), .ZN(new_n487));
  NAND3_X1  g286(.A1(new_n485), .A2(new_n486), .A3(new_n487), .ZN(new_n488));
  NAND4_X1  g287(.A1(new_n435), .A2(new_n439), .A3(new_n412), .A4(new_n413), .ZN(new_n489));
  NAND3_X1  g288(.A1(new_n488), .A2(new_n489), .A3(new_n462), .ZN(new_n490));
  OAI21_X1  g289(.A(new_n477), .B1(new_n484), .B2(new_n490), .ZN(new_n491));
  NAND4_X1  g290(.A1(new_n481), .A2(new_n483), .A3(new_n478), .A4(new_n447), .ZN(new_n492));
  NAND4_X1  g291(.A1(new_n442), .A2(KEYINPUT88), .A3(new_n492), .A4(new_n462), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n483), .A2(new_n447), .ZN(new_n494));
  AOI21_X1  g293(.A(new_n482), .B1(new_n464), .B2(new_n453), .ZN(new_n495));
  OAI21_X1  g294(.A(KEYINPUT38), .B1(new_n494), .B2(new_n495), .ZN(new_n496));
  AND3_X1   g295(.A1(new_n491), .A2(new_n493), .A3(new_n496), .ZN(new_n497));
  INV_X1    g296(.A(KEYINPUT87), .ZN(new_n498));
  AOI21_X1  g297(.A(new_n424), .B1(new_n438), .B2(new_n429), .ZN(new_n499));
  INV_X1    g298(.A(KEYINPUT39), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  INV_X1    g300(.A(new_n412), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  NAND3_X1  g302(.A1(new_n417), .A2(new_n424), .A3(new_n422), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n504), .A2(KEYINPUT39), .ZN(new_n505));
  NOR2_X1   g304(.A1(new_n499), .A2(new_n505), .ZN(new_n506));
  OAI21_X1  g305(.A(new_n498), .B1(new_n503), .B2(new_n506), .ZN(new_n507));
  INV_X1    g306(.A(KEYINPUT40), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  OR2_X1    g308(.A1(new_n499), .A2(new_n505), .ZN(new_n510));
  AOI21_X1  g309(.A(new_n412), .B1(new_n499), .B2(new_n500), .ZN(new_n511));
  AOI21_X1  g310(.A(KEYINPUT87), .B1(new_n510), .B2(new_n511), .ZN(new_n512));
  NAND2_X1  g311(.A1(new_n512), .A2(KEYINPUT40), .ZN(new_n513));
  AND2_X1   g312(.A1(new_n509), .A2(new_n513), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n485), .A2(new_n412), .ZN(new_n515));
  NAND3_X1  g314(.A1(new_n463), .A2(new_n466), .A3(new_n515), .ZN(new_n516));
  OAI21_X1  g315(.A(new_n277), .B1(new_n514), .B2(new_n516), .ZN(new_n517));
  OAI21_X1  g316(.A(new_n476), .B1(new_n497), .B2(new_n517), .ZN(new_n518));
  AND3_X1   g317(.A1(new_n463), .A2(new_n466), .A3(new_n515), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n509), .A2(new_n513), .ZN(new_n520));
  AOI22_X1  g319(.A1(new_n519), .A2(new_n520), .B1(new_n275), .B2(new_n276), .ZN(new_n521));
  NAND3_X1  g320(.A1(new_n491), .A2(new_n493), .A3(new_n496), .ZN(new_n522));
  NAND3_X1  g321(.A1(new_n521), .A2(new_n522), .A3(KEYINPUT89), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n518), .A2(new_n523), .ZN(new_n524));
  INV_X1    g323(.A(KEYINPUT75), .ZN(new_n525));
  AND3_X1   g324(.A1(new_n381), .A2(new_n393), .A3(new_n395), .ZN(new_n526));
  AOI21_X1  g325(.A(new_n393), .B1(new_n381), .B2(new_n395), .ZN(new_n527));
  OAI21_X1  g326(.A(new_n525), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  INV_X1    g327(.A(KEYINPUT36), .ZN(new_n529));
  NAND2_X1  g328(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  INV_X1    g329(.A(new_n467), .ZN(new_n531));
  OAI211_X1 g330(.A(new_n276), .B(new_n275), .C1(new_n531), .C2(new_n442), .ZN(new_n532));
  NAND3_X1  g331(.A1(new_n471), .A2(new_n525), .A3(KEYINPUT36), .ZN(new_n533));
  AND3_X1   g332(.A1(new_n530), .A2(new_n532), .A3(new_n533), .ZN(new_n534));
  AOI21_X1  g333(.A(new_n475), .B1(new_n524), .B2(new_n534), .ZN(new_n535));
  XNOR2_X1  g334(.A(G113gat), .B(G141gat), .ZN(new_n536));
  XNOR2_X1  g335(.A(new_n536), .B(G197gat), .ZN(new_n537));
  XOR2_X1   g336(.A(KEYINPUT11), .B(G169gat), .Z(new_n538));
  XNOR2_X1  g337(.A(new_n537), .B(new_n538), .ZN(new_n539));
  XNOR2_X1  g338(.A(new_n539), .B(KEYINPUT12), .ZN(new_n540));
  XNOR2_X1  g339(.A(G15gat), .B(G22gat), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n541), .A2(KEYINPUT92), .ZN(new_n542));
  INV_X1    g341(.A(G8gat), .ZN(new_n543));
  XNOR2_X1  g342(.A(new_n542), .B(new_n543), .ZN(new_n544));
  INV_X1    g343(.A(KEYINPUT16), .ZN(new_n545));
  AOI21_X1  g344(.A(G1gat), .B1(new_n541), .B2(new_n545), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n544), .A2(new_n546), .ZN(new_n547));
  XNOR2_X1  g346(.A(new_n542), .B(G8gat), .ZN(new_n548));
  INV_X1    g347(.A(new_n546), .ZN(new_n549));
  NAND2_X1  g348(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n547), .A2(new_n550), .ZN(new_n551));
  INV_X1    g350(.A(G29gat), .ZN(new_n552));
  NAND3_X1  g351(.A1(new_n552), .A2(KEYINPUT14), .A3(G36gat), .ZN(new_n553));
  XOR2_X1   g352(.A(KEYINPUT14), .B(G29gat), .Z(new_n554));
  OAI21_X1  g353(.A(new_n553), .B1(new_n554), .B2(G36gat), .ZN(new_n555));
  INV_X1    g354(.A(KEYINPUT15), .ZN(new_n556));
  OR2_X1    g355(.A1(G43gat), .A2(G50gat), .ZN(new_n557));
  NAND2_X1  g356(.A1(G43gat), .A2(G50gat), .ZN(new_n558));
  AOI21_X1  g357(.A(new_n556), .B1(new_n557), .B2(new_n558), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n555), .A2(new_n559), .ZN(new_n560));
  INV_X1    g359(.A(new_n560), .ZN(new_n561));
  XNOR2_X1  g360(.A(KEYINPUT91), .B(G43gat), .ZN(new_n562));
  OAI211_X1 g361(.A(new_n556), .B(new_n558), .C1(new_n562), .C2(G50gat), .ZN(new_n563));
  AOI21_X1  g362(.A(new_n559), .B1(new_n555), .B2(new_n563), .ZN(new_n564));
  OAI21_X1  g363(.A(KEYINPUT17), .B1(new_n561), .B2(new_n564), .ZN(new_n565));
  INV_X1    g364(.A(KEYINPUT17), .ZN(new_n566));
  AND2_X1   g365(.A1(new_n555), .A2(new_n563), .ZN(new_n567));
  OAI211_X1 g366(.A(new_n566), .B(new_n560), .C1(new_n567), .C2(new_n559), .ZN(new_n568));
  NAND3_X1  g367(.A1(new_n551), .A2(new_n565), .A3(new_n568), .ZN(new_n569));
  NAND2_X1  g368(.A1(G229gat), .A2(G233gat), .ZN(new_n570));
  NOR2_X1   g369(.A1(new_n561), .A2(new_n564), .ZN(new_n571));
  NAND3_X1  g370(.A1(new_n571), .A2(new_n547), .A3(new_n550), .ZN(new_n572));
  NAND3_X1  g371(.A1(new_n569), .A2(new_n570), .A3(new_n572), .ZN(new_n573));
  INV_X1    g372(.A(KEYINPUT18), .ZN(new_n574));
  OAI21_X1  g373(.A(new_n551), .B1(new_n564), .B2(new_n561), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n575), .A2(new_n572), .ZN(new_n576));
  XOR2_X1   g375(.A(new_n570), .B(KEYINPUT13), .Z(new_n577));
  AOI22_X1  g376(.A1(new_n573), .A2(new_n574), .B1(new_n576), .B2(new_n577), .ZN(new_n578));
  NAND4_X1  g377(.A1(new_n569), .A2(KEYINPUT18), .A3(new_n570), .A4(new_n572), .ZN(new_n579));
  AOI21_X1  g378(.A(new_n540), .B1(new_n578), .B2(new_n579), .ZN(new_n580));
  NAND2_X1  g379(.A1(new_n573), .A2(new_n574), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n576), .A2(new_n577), .ZN(new_n582));
  AND4_X1   g381(.A1(new_n540), .A2(new_n581), .A3(new_n579), .A4(new_n582), .ZN(new_n583));
  NOR2_X1   g382(.A1(new_n580), .A2(new_n583), .ZN(new_n584));
  NOR2_X1   g383(.A1(new_n535), .A2(new_n584), .ZN(new_n585));
  XOR2_X1   g384(.A(G71gat), .B(G78gat), .Z(new_n586));
  INV_X1    g385(.A(new_n586), .ZN(new_n587));
  INV_X1    g386(.A(KEYINPUT9), .ZN(new_n588));
  INV_X1    g387(.A(G71gat), .ZN(new_n589));
  INV_X1    g388(.A(G78gat), .ZN(new_n590));
  OAI21_X1  g389(.A(new_n588), .B1(new_n589), .B2(new_n590), .ZN(new_n591));
  XOR2_X1   g390(.A(G57gat), .B(G64gat), .Z(new_n592));
  NAND3_X1  g391(.A1(new_n587), .A2(new_n591), .A3(new_n592), .ZN(new_n593));
  NAND2_X1  g392(.A1(new_n592), .A2(new_n591), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n594), .A2(new_n586), .ZN(new_n595));
  NAND2_X1  g394(.A1(new_n593), .A2(new_n595), .ZN(new_n596));
  INV_X1    g395(.A(KEYINPUT93), .ZN(new_n597));
  XNOR2_X1  g396(.A(new_n596), .B(new_n597), .ZN(new_n598));
  INV_X1    g397(.A(KEYINPUT21), .ZN(new_n599));
  OAI21_X1  g398(.A(new_n551), .B1(new_n598), .B2(new_n599), .ZN(new_n600));
  XNOR2_X1  g399(.A(new_n600), .B(KEYINPUT94), .ZN(new_n601));
  XNOR2_X1  g400(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n602));
  XNOR2_X1  g401(.A(new_n602), .B(new_n205), .ZN(new_n603));
  XOR2_X1   g402(.A(new_n601), .B(new_n603), .Z(new_n604));
  NAND2_X1  g403(.A1(new_n596), .A2(new_n599), .ZN(new_n605));
  NAND2_X1  g404(.A1(G231gat), .A2(G233gat), .ZN(new_n606));
  XNOR2_X1  g405(.A(new_n605), .B(new_n606), .ZN(new_n607));
  XNOR2_X1  g406(.A(new_n607), .B(G127gat), .ZN(new_n608));
  XOR2_X1   g407(.A(G183gat), .B(G211gat), .Z(new_n609));
  OR2_X1    g408(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  NAND2_X1  g409(.A1(new_n608), .A2(new_n609), .ZN(new_n611));
  AND2_X1   g410(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  OR2_X1    g411(.A1(new_n604), .A2(new_n612), .ZN(new_n613));
  NAND3_X1  g412(.A1(new_n604), .A2(new_n610), .A3(new_n611), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  INV_X1    g414(.A(new_n615), .ZN(new_n616));
  XNOR2_X1  g415(.A(G190gat), .B(G218gat), .ZN(new_n617));
  AND3_X1   g416(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n618));
  INV_X1    g417(.A(KEYINPUT95), .ZN(new_n619));
  INV_X1    g418(.A(G85gat), .ZN(new_n620));
  INV_X1    g419(.A(G92gat), .ZN(new_n621));
  OAI21_X1  g420(.A(new_n619), .B1(new_n620), .B2(new_n621), .ZN(new_n622));
  NAND3_X1  g421(.A1(KEYINPUT95), .A2(G85gat), .A3(G92gat), .ZN(new_n623));
  NAND3_X1  g422(.A1(new_n622), .A2(KEYINPUT7), .A3(new_n623), .ZN(new_n624));
  INV_X1    g423(.A(KEYINPUT7), .ZN(new_n625));
  OAI211_X1 g424(.A(new_n619), .B(new_n625), .C1(new_n620), .C2(new_n621), .ZN(new_n626));
  NAND2_X1  g425(.A1(G99gat), .A2(G106gat), .ZN(new_n627));
  AOI22_X1  g426(.A1(KEYINPUT8), .A2(new_n627), .B1(new_n620), .B2(new_n621), .ZN(new_n628));
  NAND3_X1  g427(.A1(new_n624), .A2(new_n626), .A3(new_n628), .ZN(new_n629));
  OR2_X1    g428(.A1(G99gat), .A2(G106gat), .ZN(new_n630));
  NAND3_X1  g429(.A1(new_n629), .A2(new_n627), .A3(new_n630), .ZN(new_n631));
  NAND2_X1  g430(.A1(new_n630), .A2(new_n627), .ZN(new_n632));
  NAND4_X1  g431(.A1(new_n624), .A2(new_n632), .A3(new_n626), .A4(new_n628), .ZN(new_n633));
  AND2_X1   g432(.A1(new_n631), .A2(new_n633), .ZN(new_n634));
  AOI21_X1  g433(.A(new_n618), .B1(new_n634), .B2(new_n571), .ZN(new_n635));
  XNOR2_X1  g434(.A(new_n634), .B(KEYINPUT96), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n568), .A2(new_n565), .ZN(new_n637));
  OAI21_X1  g436(.A(new_n635), .B1(new_n636), .B2(new_n637), .ZN(new_n638));
  OAI21_X1  g437(.A(new_n617), .B1(new_n638), .B2(KEYINPUT97), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n638), .A2(KEYINPUT97), .ZN(new_n640));
  XNOR2_X1  g439(.A(new_n639), .B(new_n640), .ZN(new_n641));
  XNOR2_X1  g440(.A(G134gat), .B(G162gat), .ZN(new_n642));
  AOI21_X1  g441(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n643));
  XOR2_X1   g442(.A(new_n642), .B(new_n643), .Z(new_n644));
  INV_X1    g443(.A(new_n644), .ZN(new_n645));
  NOR2_X1   g444(.A1(new_n645), .A2(KEYINPUT98), .ZN(new_n646));
  OR2_X1    g445(.A1(new_n641), .A2(new_n646), .ZN(new_n647));
  AND2_X1   g446(.A1(new_n645), .A2(KEYINPUT98), .ZN(new_n648));
  OAI21_X1  g447(.A(new_n641), .B1(new_n648), .B2(new_n646), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n647), .A2(new_n649), .ZN(new_n650));
  NOR2_X1   g449(.A1(new_n616), .A2(new_n650), .ZN(new_n651));
  XNOR2_X1  g450(.A(G120gat), .B(G148gat), .ZN(new_n652));
  XNOR2_X1  g451(.A(G176gat), .B(G204gat), .ZN(new_n653));
  XOR2_X1   g452(.A(new_n652), .B(new_n653), .Z(new_n654));
  INV_X1    g453(.A(KEYINPUT10), .ZN(new_n655));
  NAND2_X1  g454(.A1(new_n631), .A2(new_n633), .ZN(new_n656));
  NOR3_X1   g455(.A1(new_n598), .A2(new_n655), .A3(new_n656), .ZN(new_n657));
  INV_X1    g456(.A(new_n657), .ZN(new_n658));
  INV_X1    g457(.A(new_n596), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n656), .A2(new_n659), .ZN(new_n660));
  NAND3_X1  g459(.A1(new_n596), .A2(new_n631), .A3(new_n633), .ZN(new_n661));
  NAND2_X1  g460(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  INV_X1    g461(.A(KEYINPUT99), .ZN(new_n663));
  NAND3_X1  g462(.A1(new_n662), .A2(new_n663), .A3(new_n655), .ZN(new_n664));
  INV_X1    g463(.A(new_n664), .ZN(new_n665));
  AOI21_X1  g464(.A(new_n663), .B1(new_n662), .B2(new_n655), .ZN(new_n666));
  OAI21_X1  g465(.A(new_n658), .B1(new_n665), .B2(new_n666), .ZN(new_n667));
  NAND2_X1  g466(.A1(G230gat), .A2(G233gat), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  NOR2_X1   g468(.A1(new_n662), .A2(new_n668), .ZN(new_n670));
  XOR2_X1   g469(.A(new_n670), .B(KEYINPUT100), .Z(new_n671));
  AOI21_X1  g470(.A(new_n654), .B1(new_n669), .B2(new_n671), .ZN(new_n672));
  INV_X1    g471(.A(new_n672), .ZN(new_n673));
  NAND3_X1  g472(.A1(new_n669), .A2(new_n671), .A3(new_n654), .ZN(new_n674));
  NAND3_X1  g473(.A1(new_n673), .A2(KEYINPUT101), .A3(new_n674), .ZN(new_n675));
  INV_X1    g474(.A(KEYINPUT101), .ZN(new_n676));
  INV_X1    g475(.A(new_n674), .ZN(new_n677));
  OAI21_X1  g476(.A(new_n676), .B1(new_n677), .B2(new_n672), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n675), .A2(new_n678), .ZN(new_n679));
  NAND3_X1  g478(.A1(new_n585), .A2(new_n651), .A3(new_n679), .ZN(new_n680));
  NOR2_X1   g479(.A1(new_n680), .A2(new_n443), .ZN(new_n681));
  XOR2_X1   g480(.A(new_n681), .B(G1gat), .Z(G1324gat));
  OR2_X1    g481(.A1(new_n680), .A2(new_n467), .ZN(new_n683));
  NOR2_X1   g482(.A1(new_n545), .A2(new_n543), .ZN(new_n684));
  NOR2_X1   g483(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n685));
  OR3_X1    g484(.A1(new_n683), .A2(new_n684), .A3(new_n685), .ZN(new_n686));
  NAND2_X1  g485(.A1(new_n683), .A2(G8gat), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  MUX2_X1   g487(.A(new_n686), .B(new_n688), .S(KEYINPUT42), .Z(G1325gat));
  AOI21_X1  g488(.A(KEYINPUT36), .B1(new_n471), .B2(new_n525), .ZN(new_n690));
  AOI211_X1 g489(.A(KEYINPUT75), .B(new_n529), .C1(new_n407), .C2(new_n396), .ZN(new_n691));
  NOR2_X1   g490(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  XOR2_X1   g491(.A(new_n692), .B(KEYINPUT102), .Z(new_n693));
  INV_X1    g492(.A(new_n693), .ZN(new_n694));
  OAI21_X1  g493(.A(G15gat), .B1(new_n680), .B2(new_n694), .ZN(new_n695));
  OR2_X1    g494(.A1(new_n471), .A2(G15gat), .ZN(new_n696));
  OAI21_X1  g495(.A(new_n695), .B1(new_n680), .B2(new_n696), .ZN(G1326gat));
  NOR2_X1   g496(.A1(new_n680), .A2(new_n277), .ZN(new_n698));
  XOR2_X1   g497(.A(KEYINPUT43), .B(G22gat), .Z(new_n699));
  XNOR2_X1  g498(.A(new_n698), .B(new_n699), .ZN(G1327gat));
  INV_X1    g499(.A(new_n650), .ZN(new_n701));
  NOR2_X1   g500(.A1(new_n535), .A2(new_n701), .ZN(new_n702));
  NAND2_X1  g501(.A1(new_n616), .A2(new_n679), .ZN(new_n703));
  NOR2_X1   g502(.A1(new_n703), .A2(new_n584), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n702), .A2(new_n704), .ZN(new_n705));
  NOR3_X1   g504(.A1(new_n705), .A2(G29gat), .A3(new_n443), .ZN(new_n706));
  XNOR2_X1  g505(.A(KEYINPUT103), .B(KEYINPUT45), .ZN(new_n707));
  XNOR2_X1  g506(.A(new_n706), .B(new_n707), .ZN(new_n708));
  INV_X1    g507(.A(KEYINPUT104), .ZN(new_n709));
  NOR2_X1   g508(.A1(new_n709), .A2(KEYINPUT44), .ZN(new_n710));
  INV_X1    g509(.A(new_n710), .ZN(new_n711));
  AND3_X1   g510(.A1(new_n521), .A2(new_n522), .A3(KEYINPUT89), .ZN(new_n712));
  AOI21_X1  g511(.A(KEYINPUT89), .B1(new_n521), .B2(new_n522), .ZN(new_n713));
  OAI211_X1 g512(.A(new_n692), .B(new_n532), .C1(new_n712), .C2(new_n713), .ZN(new_n714));
  INV_X1    g513(.A(new_n475), .ZN(new_n715));
  NAND2_X1  g514(.A1(new_n714), .A2(new_n715), .ZN(new_n716));
  AOI21_X1  g515(.A(new_n711), .B1(new_n716), .B2(new_n650), .ZN(new_n717));
  XNOR2_X1  g516(.A(KEYINPUT104), .B(KEYINPUT44), .ZN(new_n718));
  INV_X1    g517(.A(new_n718), .ZN(new_n719));
  AOI211_X1 g518(.A(new_n701), .B(new_n719), .C1(new_n714), .C2(new_n715), .ZN(new_n720));
  NOR2_X1   g519(.A1(new_n717), .A2(new_n720), .ZN(new_n721));
  AND2_X1   g520(.A1(new_n721), .A2(new_n704), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n722), .A2(new_n442), .ZN(new_n723));
  NAND2_X1  g522(.A1(new_n723), .A2(KEYINPUT105), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n724), .A2(G29gat), .ZN(new_n725));
  NOR2_X1   g524(.A1(new_n723), .A2(KEYINPUT105), .ZN(new_n726));
  OAI21_X1  g525(.A(new_n708), .B1(new_n725), .B2(new_n726), .ZN(G1328gat));
  AND2_X1   g526(.A1(KEYINPUT106), .A2(KEYINPUT46), .ZN(new_n728));
  NOR2_X1   g527(.A1(KEYINPUT106), .A2(KEYINPUT46), .ZN(new_n729));
  NOR2_X1   g528(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  NOR3_X1   g529(.A1(new_n705), .A2(G36gat), .A3(new_n467), .ZN(new_n731));
  MUX2_X1   g530(.A(new_n730), .B(new_n728), .S(new_n731), .Z(new_n732));
  INV_X1    g531(.A(new_n722), .ZN(new_n733));
  OAI21_X1  g532(.A(G36gat), .B1(new_n733), .B2(new_n467), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n732), .A2(new_n734), .ZN(G1329gat));
  NOR3_X1   g534(.A1(new_n705), .A2(new_n562), .A3(new_n471), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n722), .A2(new_n693), .ZN(new_n737));
  AOI21_X1  g536(.A(new_n736), .B1(new_n737), .B2(new_n562), .ZN(new_n738));
  INV_X1    g537(.A(new_n562), .ZN(new_n739));
  INV_X1    g538(.A(new_n692), .ZN(new_n740));
  AOI21_X1  g539(.A(new_n739), .B1(new_n722), .B2(new_n740), .ZN(new_n741));
  INV_X1    g540(.A(KEYINPUT47), .ZN(new_n742));
  OR2_X1    g541(.A1(new_n736), .A2(new_n742), .ZN(new_n743));
  OAI22_X1  g542(.A1(new_n738), .A2(KEYINPUT47), .B1(new_n741), .B2(new_n743), .ZN(G1330gat));
  INV_X1    g543(.A(KEYINPUT48), .ZN(new_n745));
  INV_X1    g544(.A(new_n277), .ZN(new_n746));
  NAND4_X1  g545(.A1(new_n721), .A2(KEYINPUT108), .A3(new_n746), .A4(new_n704), .ZN(new_n747));
  OAI21_X1  g546(.A(new_n710), .B1(new_n535), .B2(new_n701), .ZN(new_n748));
  NAND3_X1  g547(.A1(new_n530), .A2(new_n532), .A3(new_n533), .ZN(new_n749));
  AOI21_X1  g548(.A(new_n749), .B1(new_n518), .B2(new_n523), .ZN(new_n750));
  OAI211_X1 g549(.A(new_n650), .B(new_n718), .C1(new_n750), .C2(new_n475), .ZN(new_n751));
  NAND4_X1  g550(.A1(new_n748), .A2(new_n746), .A3(new_n704), .A4(new_n751), .ZN(new_n752));
  INV_X1    g551(.A(KEYINPUT108), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  NAND3_X1  g553(.A1(new_n747), .A2(G50gat), .A3(new_n754), .ZN(new_n755));
  NOR4_X1   g554(.A1(new_n703), .A2(new_n701), .A3(G50gat), .A4(new_n277), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n585), .A2(new_n756), .ZN(new_n757));
  AOI21_X1  g556(.A(new_n745), .B1(new_n755), .B2(new_n757), .ZN(new_n758));
  INV_X1    g557(.A(KEYINPUT107), .ZN(new_n759));
  NAND3_X1  g558(.A1(new_n752), .A2(new_n759), .A3(G50gat), .ZN(new_n760));
  AOI21_X1  g559(.A(KEYINPUT48), .B1(new_n585), .B2(new_n756), .ZN(new_n761));
  NAND2_X1  g560(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  AOI21_X1  g561(.A(new_n759), .B1(new_n752), .B2(G50gat), .ZN(new_n763));
  NOR2_X1   g562(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  NOR3_X1   g563(.A1(new_n758), .A2(KEYINPUT109), .A3(new_n764), .ZN(new_n765));
  INV_X1    g564(.A(KEYINPUT109), .ZN(new_n766));
  AND2_X1   g565(.A1(new_n752), .A2(new_n753), .ZN(new_n767));
  OAI21_X1  g566(.A(G50gat), .B1(new_n752), .B2(new_n753), .ZN(new_n768));
  OAI21_X1  g567(.A(new_n757), .B1(new_n767), .B2(new_n768), .ZN(new_n769));
  NAND2_X1  g568(.A1(new_n769), .A2(KEYINPUT48), .ZN(new_n770));
  OR2_X1    g569(.A1(new_n762), .A2(new_n763), .ZN(new_n771));
  AOI21_X1  g570(.A(new_n766), .B1(new_n770), .B2(new_n771), .ZN(new_n772));
  NOR2_X1   g571(.A1(new_n765), .A2(new_n772), .ZN(G1331gat));
  INV_X1    g572(.A(new_n584), .ZN(new_n774));
  NOR4_X1   g573(.A1(new_n616), .A2(new_n650), .A3(new_n679), .A4(new_n774), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n716), .A2(new_n775), .ZN(new_n776));
  INV_X1    g575(.A(new_n776), .ZN(new_n777));
  NAND2_X1  g576(.A1(new_n777), .A2(new_n442), .ZN(new_n778));
  XNOR2_X1  g577(.A(new_n778), .B(G57gat), .ZN(G1332gat));
  NOR2_X1   g578(.A1(new_n776), .A2(new_n467), .ZN(new_n780));
  NOR2_X1   g579(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n781));
  AND2_X1   g580(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n782));
  OAI21_X1  g581(.A(new_n780), .B1(new_n781), .B2(new_n782), .ZN(new_n783));
  OAI21_X1  g582(.A(new_n783), .B1(new_n780), .B2(new_n781), .ZN(G1333gat));
  NOR3_X1   g583(.A1(new_n776), .A2(G71gat), .A3(new_n471), .ZN(new_n785));
  NAND2_X1  g584(.A1(new_n777), .A2(new_n693), .ZN(new_n786));
  AOI21_X1  g585(.A(new_n785), .B1(G71gat), .B2(new_n786), .ZN(new_n787));
  XNOR2_X1  g586(.A(new_n787), .B(KEYINPUT50), .ZN(G1334gat));
  NOR2_X1   g587(.A1(new_n776), .A2(new_n277), .ZN(new_n789));
  XNOR2_X1  g588(.A(new_n789), .B(new_n590), .ZN(G1335gat));
  NOR2_X1   g589(.A1(new_n615), .A2(new_n774), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n702), .A2(new_n791), .ZN(new_n792));
  INV_X1    g591(.A(KEYINPUT51), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n792), .A2(new_n793), .ZN(new_n794));
  NAND3_X1  g593(.A1(new_n702), .A2(KEYINPUT51), .A3(new_n791), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  INV_X1    g595(.A(new_n679), .ZN(new_n797));
  NAND4_X1  g596(.A1(new_n796), .A2(new_n620), .A3(new_n442), .A4(new_n797), .ZN(new_n798));
  NOR3_X1   g597(.A1(new_n679), .A2(new_n615), .A3(new_n774), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n721), .A2(new_n799), .ZN(new_n800));
  OAI21_X1  g599(.A(G85gat), .B1(new_n800), .B2(new_n443), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n798), .A2(new_n801), .ZN(G1336gat));
  NOR2_X1   g601(.A1(new_n467), .A2(G92gat), .ZN(new_n803));
  AND3_X1   g602(.A1(new_n796), .A2(new_n797), .A3(new_n803), .ZN(new_n804));
  NOR2_X1   g603(.A1(new_n804), .A2(KEYINPUT52), .ZN(new_n805));
  NAND3_X1  g604(.A1(new_n721), .A2(new_n531), .A3(new_n799), .ZN(new_n806));
  NOR2_X1   g605(.A1(new_n806), .A2(KEYINPUT110), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n806), .A2(KEYINPUT110), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n808), .A2(G92gat), .ZN(new_n809));
  OAI21_X1  g608(.A(new_n805), .B1(new_n807), .B2(new_n809), .ZN(new_n810));
  AND2_X1   g609(.A1(new_n806), .A2(G92gat), .ZN(new_n811));
  OAI21_X1  g610(.A(KEYINPUT52), .B1(new_n804), .B2(new_n811), .ZN(new_n812));
  NAND2_X1  g611(.A1(new_n810), .A2(new_n812), .ZN(G1337gat));
  OAI21_X1  g612(.A(G99gat), .B1(new_n800), .B2(new_n694), .ZN(new_n814));
  INV_X1    g613(.A(new_n796), .ZN(new_n815));
  NOR2_X1   g614(.A1(new_n679), .A2(new_n471), .ZN(new_n816));
  INV_X1    g615(.A(new_n816), .ZN(new_n817));
  NOR2_X1   g616(.A1(new_n817), .A2(G99gat), .ZN(new_n818));
  XNOR2_X1  g617(.A(new_n818), .B(KEYINPUT111), .ZN(new_n819));
  OAI21_X1  g618(.A(new_n814), .B1(new_n815), .B2(new_n819), .ZN(G1338gat));
  INV_X1    g619(.A(KEYINPUT53), .ZN(new_n821));
  NOR2_X1   g620(.A1(new_n277), .A2(G106gat), .ZN(new_n822));
  NAND3_X1  g621(.A1(new_n796), .A2(new_n797), .A3(new_n822), .ZN(new_n823));
  AOI21_X1  g622(.A(new_n821), .B1(new_n823), .B2(KEYINPUT112), .ZN(new_n824));
  OAI21_X1  g623(.A(G106gat), .B1(new_n800), .B2(new_n277), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n823), .A2(new_n825), .ZN(new_n826));
  XNOR2_X1  g625(.A(new_n824), .B(new_n826), .ZN(G1339gat));
  INV_X1    g626(.A(new_n583), .ZN(new_n828));
  NOR2_X1   g627(.A1(new_n576), .A2(new_n577), .ZN(new_n829));
  AOI21_X1  g628(.A(new_n570), .B1(new_n569), .B2(new_n572), .ZN(new_n830));
  OAI21_X1  g629(.A(new_n539), .B1(new_n829), .B2(new_n830), .ZN(new_n831));
  NAND2_X1  g630(.A1(new_n828), .A2(new_n831), .ZN(new_n832));
  AOI21_X1  g631(.A(new_n832), .B1(new_n647), .B2(new_n649), .ZN(new_n833));
  INV_X1    g632(.A(KEYINPUT114), .ZN(new_n834));
  INV_X1    g633(.A(new_n654), .ZN(new_n835));
  XNOR2_X1  g634(.A(KEYINPUT113), .B(KEYINPUT54), .ZN(new_n836));
  NAND3_X1  g635(.A1(new_n667), .A2(new_n668), .A3(new_n836), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n662), .A2(new_n655), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n838), .A2(KEYINPUT99), .ZN(new_n839));
  AOI21_X1  g638(.A(new_n657), .B1(new_n839), .B2(new_n664), .ZN(new_n840));
  INV_X1    g639(.A(new_n668), .ZN(new_n841));
  OAI21_X1  g640(.A(KEYINPUT54), .B1(new_n840), .B2(new_n841), .ZN(new_n842));
  NOR2_X1   g641(.A1(new_n667), .A2(new_n668), .ZN(new_n843));
  OAI211_X1 g642(.A(new_n835), .B(new_n837), .C1(new_n842), .C2(new_n843), .ZN(new_n844));
  INV_X1    g643(.A(KEYINPUT55), .ZN(new_n845));
  OAI21_X1  g644(.A(new_n834), .B1(new_n844), .B2(new_n845), .ZN(new_n846));
  AND2_X1   g645(.A1(new_n837), .A2(new_n835), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n840), .A2(new_n841), .ZN(new_n848));
  NAND3_X1  g647(.A1(new_n669), .A2(new_n848), .A3(KEYINPUT54), .ZN(new_n849));
  NAND4_X1  g648(.A1(new_n847), .A2(new_n849), .A3(KEYINPUT114), .A4(KEYINPUT55), .ZN(new_n850));
  AND2_X1   g649(.A1(new_n850), .A2(new_n674), .ZN(new_n851));
  NAND2_X1  g650(.A1(new_n844), .A2(new_n845), .ZN(new_n852));
  NAND4_X1  g651(.A1(new_n833), .A2(new_n846), .A3(new_n851), .A4(new_n852), .ZN(new_n853));
  INV_X1    g652(.A(new_n853), .ZN(new_n854));
  AOI21_X1  g653(.A(new_n584), .B1(new_n844), .B2(new_n845), .ZN(new_n855));
  NAND4_X1  g654(.A1(new_n846), .A2(new_n855), .A3(new_n674), .A4(new_n850), .ZN(new_n856));
  NAND4_X1  g655(.A1(new_n675), .A2(new_n678), .A3(new_n828), .A4(new_n831), .ZN(new_n857));
  AOI21_X1  g656(.A(new_n650), .B1(new_n856), .B2(new_n857), .ZN(new_n858));
  OAI21_X1  g657(.A(new_n616), .B1(new_n854), .B2(new_n858), .ZN(new_n859));
  NAND3_X1  g658(.A1(new_n651), .A2(new_n584), .A3(new_n679), .ZN(new_n860));
  AOI21_X1  g659(.A(new_n746), .B1(new_n859), .B2(new_n860), .ZN(new_n861));
  NOR2_X1   g660(.A1(new_n531), .A2(new_n443), .ZN(new_n862));
  AND2_X1   g661(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n863), .A2(new_n472), .ZN(new_n864));
  NOR3_X1   g663(.A1(new_n864), .A2(new_n351), .A3(new_n584), .ZN(new_n865));
  AOI211_X1 g664(.A(new_n443), .B(new_n408), .C1(new_n859), .C2(new_n860), .ZN(new_n866));
  AND2_X1   g665(.A1(new_n866), .A2(new_n467), .ZN(new_n867));
  AOI21_X1  g666(.A(G113gat), .B1(new_n867), .B2(new_n774), .ZN(new_n868));
  NOR2_X1   g667(.A1(new_n865), .A2(new_n868), .ZN(G1340gat));
  AOI21_X1  g668(.A(G120gat), .B1(new_n867), .B2(new_n797), .ZN(new_n870));
  NOR2_X1   g669(.A1(new_n817), .A2(new_n349), .ZN(new_n871));
  AOI21_X1  g670(.A(new_n870), .B1(new_n863), .B2(new_n871), .ZN(G1341gat));
  OAI21_X1  g671(.A(G127gat), .B1(new_n864), .B2(new_n616), .ZN(new_n873));
  NAND3_X1  g672(.A1(new_n867), .A2(new_n357), .A3(new_n615), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  XOR2_X1   g674(.A(new_n875), .B(KEYINPUT115), .Z(G1342gat));
  NAND2_X1  g675(.A1(new_n650), .A2(new_n467), .ZN(new_n877));
  XOR2_X1   g676(.A(new_n877), .B(KEYINPUT116), .Z(new_n878));
  INV_X1    g677(.A(new_n878), .ZN(new_n879));
  NAND3_X1  g678(.A1(new_n866), .A2(new_n359), .A3(new_n879), .ZN(new_n880));
  XOR2_X1   g679(.A(KEYINPUT117), .B(KEYINPUT56), .Z(new_n881));
  XNOR2_X1  g680(.A(new_n880), .B(new_n881), .ZN(new_n882));
  OAI21_X1  g681(.A(G134gat), .B1(new_n864), .B2(new_n701), .ZN(new_n883));
  AND2_X1   g682(.A1(new_n883), .A2(KEYINPUT118), .ZN(new_n884));
  NOR2_X1   g683(.A1(new_n883), .A2(KEYINPUT118), .ZN(new_n885));
  OAI21_X1  g684(.A(new_n882), .B1(new_n884), .B2(new_n885), .ZN(G1343gat));
  NAND2_X1  g685(.A1(new_n692), .A2(new_n862), .ZN(new_n887));
  INV_X1    g686(.A(new_n887), .ZN(new_n888));
  INV_X1    g687(.A(KEYINPUT57), .ZN(new_n889));
  NOR2_X1   g688(.A1(new_n277), .A2(new_n889), .ZN(new_n890));
  INV_X1    g689(.A(new_n890), .ZN(new_n891));
  OAI21_X1  g690(.A(new_n853), .B1(new_n858), .B2(KEYINPUT119), .ZN(new_n892));
  INV_X1    g691(.A(KEYINPUT119), .ZN(new_n893));
  AOI211_X1 g692(.A(new_n893), .B(new_n650), .C1(new_n856), .C2(new_n857), .ZN(new_n894));
  OAI211_X1 g693(.A(KEYINPUT120), .B(new_n616), .C1(new_n892), .C2(new_n894), .ZN(new_n895));
  AND2_X1   g694(.A1(new_n895), .A2(new_n860), .ZN(new_n896));
  OAI21_X1  g695(.A(new_n616), .B1(new_n892), .B2(new_n894), .ZN(new_n897));
  INV_X1    g696(.A(KEYINPUT120), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  AOI21_X1  g698(.A(new_n891), .B1(new_n896), .B2(new_n899), .ZN(new_n900));
  NAND2_X1  g699(.A1(new_n859), .A2(new_n860), .ZN(new_n901));
  AOI21_X1  g700(.A(KEYINPUT57), .B1(new_n901), .B2(new_n746), .ZN(new_n902));
  OAI211_X1 g701(.A(new_n774), .B(new_n888), .C1(new_n900), .C2(new_n902), .ZN(new_n903));
  NAND2_X1  g702(.A1(new_n903), .A2(KEYINPUT122), .ZN(new_n904));
  AND2_X1   g703(.A1(new_n897), .A2(new_n898), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n895), .A2(new_n860), .ZN(new_n906));
  OAI21_X1  g705(.A(new_n890), .B1(new_n905), .B2(new_n906), .ZN(new_n907));
  INV_X1    g706(.A(new_n902), .ZN(new_n908));
  AOI21_X1  g707(.A(new_n887), .B1(new_n907), .B2(new_n908), .ZN(new_n909));
  INV_X1    g708(.A(KEYINPUT122), .ZN(new_n910));
  NAND3_X1  g709(.A1(new_n909), .A2(new_n910), .A3(new_n774), .ZN(new_n911));
  NAND3_X1  g710(.A1(new_n904), .A2(G141gat), .A3(new_n911), .ZN(new_n912));
  NAND4_X1  g711(.A1(new_n901), .A2(new_n442), .A3(new_n746), .A4(new_n694), .ZN(new_n913));
  NOR2_X1   g712(.A1(new_n913), .A2(new_n531), .ZN(new_n914));
  NOR2_X1   g713(.A1(new_n584), .A2(G141gat), .ZN(new_n915));
  XNOR2_X1  g714(.A(new_n915), .B(KEYINPUT121), .ZN(new_n916));
  AND2_X1   g715(.A1(new_n914), .A2(new_n916), .ZN(new_n917));
  NOR2_X1   g716(.A1(new_n917), .A2(KEYINPUT58), .ZN(new_n918));
  NAND2_X1  g717(.A1(new_n912), .A2(new_n918), .ZN(new_n919));
  AOI21_X1  g718(.A(new_n217), .B1(new_n909), .B2(new_n774), .ZN(new_n920));
  OAI21_X1  g719(.A(KEYINPUT58), .B1(new_n920), .B2(new_n917), .ZN(new_n921));
  NAND2_X1  g720(.A1(new_n919), .A2(new_n921), .ZN(G1344gat));
  NAND3_X1  g721(.A1(new_n914), .A2(new_n222), .A3(new_n797), .ZN(new_n923));
  INV_X1    g722(.A(KEYINPUT59), .ZN(new_n924));
  AOI21_X1  g723(.A(new_n891), .B1(new_n859), .B2(new_n860), .ZN(new_n925));
  OR2_X1    g724(.A1(new_n902), .A2(new_n925), .ZN(new_n926));
  NOR2_X1   g725(.A1(new_n887), .A2(new_n679), .ZN(new_n927));
  NAND2_X1  g726(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  INV_X1    g727(.A(KEYINPUT123), .ZN(new_n929));
  NAND2_X1  g728(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  OAI211_X1 g729(.A(KEYINPUT123), .B(new_n927), .C1(new_n902), .C2(new_n925), .ZN(new_n931));
  AND2_X1   g730(.A1(new_n931), .A2(G148gat), .ZN(new_n932));
  AOI21_X1  g731(.A(new_n924), .B1(new_n930), .B2(new_n932), .ZN(new_n933));
  AOI211_X1 g732(.A(KEYINPUT59), .B(new_n222), .C1(new_n909), .C2(new_n797), .ZN(new_n934));
  OAI21_X1  g733(.A(new_n923), .B1(new_n933), .B2(new_n934), .ZN(G1345gat));
  NAND3_X1  g734(.A1(new_n914), .A2(new_n205), .A3(new_n615), .ZN(new_n936));
  AND2_X1   g735(.A1(new_n909), .A2(new_n615), .ZN(new_n937));
  OAI21_X1  g736(.A(new_n936), .B1(new_n937), .B2(new_n205), .ZN(G1346gat));
  AND2_X1   g737(.A1(new_n909), .A2(new_n650), .ZN(new_n939));
  NAND2_X1  g738(.A1(new_n879), .A2(new_n206), .ZN(new_n940));
  OAI22_X1  g739(.A1(new_n939), .A2(new_n206), .B1(new_n913), .B2(new_n940), .ZN(G1347gat));
  NAND4_X1  g740(.A1(new_n861), .A2(new_n443), .A3(new_n531), .A4(new_n472), .ZN(new_n942));
  NOR3_X1   g741(.A1(new_n942), .A2(new_n283), .A3(new_n584), .ZN(new_n943));
  AOI21_X1  g742(.A(new_n442), .B1(new_n859), .B2(new_n860), .ZN(new_n944));
  AND4_X1   g743(.A1(new_n277), .A2(new_n944), .A3(new_n531), .A4(new_n472), .ZN(new_n945));
  NAND2_X1  g744(.A1(new_n945), .A2(new_n774), .ZN(new_n946));
  AOI21_X1  g745(.A(new_n943), .B1(new_n283), .B2(new_n946), .ZN(G1348gat));
  AOI21_X1  g746(.A(G176gat), .B1(new_n945), .B2(new_n797), .ZN(new_n948));
  XNOR2_X1  g747(.A(new_n948), .B(KEYINPUT124), .ZN(new_n949));
  NOR3_X1   g748(.A1(new_n942), .A2(new_n328), .A3(new_n679), .ZN(new_n950));
  NOR2_X1   g749(.A1(new_n949), .A2(new_n950), .ZN(G1349gat));
  NAND3_X1  g750(.A1(new_n945), .A2(new_n305), .A3(new_n615), .ZN(new_n952));
  NAND2_X1  g751(.A1(new_n300), .A2(new_n302), .ZN(new_n953));
  OAI21_X1  g752(.A(new_n953), .B1(new_n942), .B2(new_n616), .ZN(new_n954));
  INV_X1    g753(.A(KEYINPUT60), .ZN(new_n955));
  AOI22_X1  g754(.A1(new_n952), .A2(new_n954), .B1(KEYINPUT125), .B2(new_n955), .ZN(new_n956));
  NOR2_X1   g755(.A1(new_n955), .A2(KEYINPUT125), .ZN(new_n957));
  XNOR2_X1  g756(.A(new_n956), .B(new_n957), .ZN(G1350gat));
  OAI21_X1  g757(.A(G190gat), .B1(new_n942), .B2(new_n701), .ZN(new_n959));
  XNOR2_X1  g758(.A(new_n959), .B(KEYINPUT61), .ZN(new_n960));
  NAND3_X1  g759(.A1(new_n945), .A2(new_n297), .A3(new_n650), .ZN(new_n961));
  NAND2_X1  g760(.A1(new_n960), .A2(new_n961), .ZN(G1351gat));
  NAND3_X1  g761(.A1(new_n694), .A2(new_n443), .A3(new_n531), .ZN(new_n963));
  XNOR2_X1  g762(.A(new_n963), .B(KEYINPUT127), .ZN(new_n964));
  NAND2_X1  g763(.A1(new_n964), .A2(new_n926), .ZN(new_n965));
  INV_X1    g764(.A(G197gat), .ZN(new_n966));
  NOR3_X1   g765(.A1(new_n965), .A2(new_n966), .A3(new_n584), .ZN(new_n967));
  NOR3_X1   g766(.A1(new_n693), .A2(new_n277), .A3(new_n467), .ZN(new_n968));
  OR2_X1    g767(.A1(new_n968), .A2(KEYINPUT126), .ZN(new_n969));
  NAND2_X1  g768(.A1(new_n968), .A2(KEYINPUT126), .ZN(new_n970));
  AND3_X1   g769(.A1(new_n969), .A2(new_n944), .A3(new_n970), .ZN(new_n971));
  AOI21_X1  g770(.A(G197gat), .B1(new_n971), .B2(new_n774), .ZN(new_n972));
  NOR2_X1   g771(.A1(new_n967), .A2(new_n972), .ZN(G1352gat));
  NOR2_X1   g772(.A1(new_n679), .A2(G204gat), .ZN(new_n974));
  NAND2_X1  g773(.A1(new_n971), .A2(new_n974), .ZN(new_n975));
  OR2_X1    g774(.A1(new_n975), .A2(KEYINPUT62), .ZN(new_n976));
  OAI21_X1  g775(.A(G204gat), .B1(new_n965), .B2(new_n679), .ZN(new_n977));
  NAND2_X1  g776(.A1(new_n975), .A2(KEYINPUT62), .ZN(new_n978));
  NAND3_X1  g777(.A1(new_n976), .A2(new_n977), .A3(new_n978), .ZN(G1353gat));
  INV_X1    g778(.A(G211gat), .ZN(new_n980));
  NAND3_X1  g779(.A1(new_n971), .A2(new_n980), .A3(new_n615), .ZN(new_n981));
  NAND3_X1  g780(.A1(new_n964), .A2(new_n615), .A3(new_n926), .ZN(new_n982));
  AND3_X1   g781(.A1(new_n982), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n983));
  AOI21_X1  g782(.A(KEYINPUT63), .B1(new_n982), .B2(G211gat), .ZN(new_n984));
  OAI21_X1  g783(.A(new_n981), .B1(new_n983), .B2(new_n984), .ZN(G1354gat));
  OAI21_X1  g784(.A(G218gat), .B1(new_n965), .B2(new_n701), .ZN(new_n986));
  INV_X1    g785(.A(G218gat), .ZN(new_n987));
  NAND3_X1  g786(.A1(new_n971), .A2(new_n987), .A3(new_n650), .ZN(new_n988));
  NAND2_X1  g787(.A1(new_n986), .A2(new_n988), .ZN(G1355gat));
endmodule


