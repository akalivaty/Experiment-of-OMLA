

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n524, n525, n526, n527,
         n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538,
         n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549,
         n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560,
         n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571,
         n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582,
         n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593,
         n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604,
         n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615,
         n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626,
         n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637,
         n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648,
         n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659,
         n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670,
         n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681,
         n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692,
         n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703,
         n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714,
         n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725,
         n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736,
         n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747,
         n748, n749, n750, n751, n752, n753, n754, n755, n756, n757, n758,
         n759, n760, n761, n762, n763, n764, n765, n766, n767, n768, n769,
         n770, n771, n772, n773, n774, n775, n776, n777, n778, n779, n780,
         n781, n782, n783, n784, n785, n786, n787, n788, n789, n790, n791,
         n792, n793, n794, n795, n796, n797, n798, n799, n800, n801, n802,
         n803, n804, n805, n806, n807, n808, n809, n810, n811, n812, n813,
         n814, n815, n816, n817, n818, n819, n820, n821, n822, n823, n824,
         n825, n826, n827, n828, n829, n830, n831, n832, n833, n834, n835,
         n836, n837, n838, n839, n840, n841, n842, n843, n844, n845, n846,
         n847, n848, n849, n850, n851, n852, n853, n854, n855, n856, n857,
         n858, n859, n860, n861, n862, n863, n864, n865, n866, n867, n868,
         n869, n870, n871, n872, n873, n874, n875, n876, n877, n878, n879,
         n880, n881, n882, n883, n884, n885, n886, n887, n888, n889, n890,
         n891, n892, n893, n894, n895, n896, n897, n898, n899, n900, n901,
         n902, n903, n904, n905, n906, n907, n908, n909, n910, n911, n912,
         n913, n914, n915, n916, n917, n918, n919, n920, n921, n922, n923,
         n924, n925, n926, n927, n928, n929, n930, n931, n932, n933, n934,
         n935, n936, n937, n938, n939, n940, n941, n942, n943, n944, n945,
         n946, n947, n948, n949, n950, n951, n952, n953, n954, n955, n956,
         n957, n958, n959, n960, n961, n962, n963, n964, n965, n966, n967,
         n968, n969, n970, n971, n972, n973, n974, n975, n976, n977, n978,
         n979, n980, n981, n982, n983, n984, n985, n986, n987, n988, n989,
         n990, n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000,
         n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010,
         n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020,
         n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030,
         n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040,
         n1041;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  BUF_X1 U556 ( .A(n885), .Z(n524) );
  NAND2_X1 U557 ( .A1(n706), .A2(n802), .ZN(n735) );
  NOR2_X2 U558 ( .A1(n539), .A2(n538), .ZN(G160) );
  NOR2_X1 U559 ( .A1(n743), .A2(n742), .ZN(n745) );
  NOR2_X1 U560 ( .A1(G164), .A2(G1384), .ZN(n802) );
  XNOR2_X1 U561 ( .A(n530), .B(KEYINPUT23), .ZN(n531) );
  AND2_X2 U562 ( .A1(n535), .A2(G2104), .ZN(n882) );
  XNOR2_X2 U563 ( .A(n736), .B(KEYINPUT91), .ZN(n787) );
  XOR2_X2 U564 ( .A(KEYINPUT17), .B(n532), .Z(n881) );
  XNOR2_X1 U565 ( .A(n745), .B(n744), .ZN(n757) );
  XNOR2_X1 U566 ( .A(n729), .B(n728), .ZN(n734) );
  AND2_X1 U567 ( .A1(n792), .A2(n766), .ZN(n765) );
  AND2_X1 U568 ( .A1(n757), .A2(n751), .ZN(n750) );
  XOR2_X1 U569 ( .A(G543), .B(KEYINPUT0), .Z(n525) );
  AND2_X1 U570 ( .A1(n784), .A2(n783), .ZN(n526) );
  OR2_X1 U571 ( .A1(n773), .A2(KEYINPUT98), .ZN(n527) );
  NOR2_X1 U572 ( .A1(n529), .A2(n832), .ZN(n528) );
  AND2_X1 U573 ( .A1(n945), .A2(n844), .ZN(n529) );
  NOR2_X1 U574 ( .A1(n953), .A2(n717), .ZN(n718) );
  INV_X1 U575 ( .A(KEYINPUT29), .ZN(n728) );
  INV_X1 U576 ( .A(KEYINPUT31), .ZN(n744) );
  NOR2_X1 U577 ( .A1(n760), .A2(n759), .ZN(n763) );
  AND2_X1 U578 ( .A1(n754), .A2(n753), .ZN(n755) );
  INV_X1 U579 ( .A(n950), .ZN(n783) );
  XOR2_X1 U580 ( .A(KEYINPUT15), .B(n609), .Z(n953) );
  INV_X1 U581 ( .A(G2105), .ZN(n535) );
  NOR2_X1 U582 ( .A1(n549), .A2(n669), .ZN(n659) );
  NOR2_X1 U583 ( .A1(G2104), .A2(n535), .ZN(n885) );
  NOR2_X1 U584 ( .A1(G543), .A2(G651), .ZN(n660) );
  NOR2_X1 U585 ( .A1(G651), .A2(n669), .ZN(n667) );
  NAND2_X1 U586 ( .A1(G101), .A2(n882), .ZN(n530) );
  XNOR2_X1 U587 ( .A(n531), .B(KEYINPUT65), .ZN(n534) );
  NOR2_X1 U588 ( .A1(G2104), .A2(G2105), .ZN(n532) );
  NAND2_X1 U589 ( .A1(G137), .A2(n881), .ZN(n533) );
  NAND2_X1 U590 ( .A1(n534), .A2(n533), .ZN(n539) );
  NAND2_X1 U591 ( .A1(G125), .A2(n524), .ZN(n537) );
  AND2_X1 U592 ( .A1(G2104), .A2(G2105), .ZN(n886) );
  NAND2_X1 U593 ( .A1(G113), .A2(n886), .ZN(n536) );
  NAND2_X1 U594 ( .A1(n537), .A2(n536), .ZN(n538) );
  AND2_X1 U595 ( .A1(G102), .A2(n882), .ZN(n543) );
  NAND2_X1 U596 ( .A1(G126), .A2(n524), .ZN(n541) );
  NAND2_X1 U597 ( .A1(G114), .A2(n886), .ZN(n540) );
  NAND2_X1 U598 ( .A1(n541), .A2(n540), .ZN(n542) );
  NOR2_X1 U599 ( .A1(n543), .A2(n542), .ZN(n545) );
  NAND2_X1 U600 ( .A1(G138), .A2(n881), .ZN(n544) );
  AND2_X1 U601 ( .A1(n545), .A2(n544), .ZN(G164) );
  INV_X1 U602 ( .A(G651), .ZN(n549) );
  NOR2_X1 U603 ( .A1(G543), .A2(n549), .ZN(n546) );
  XOR2_X1 U604 ( .A(KEYINPUT1), .B(n546), .Z(n673) );
  NAND2_X1 U605 ( .A1(G64), .A2(n673), .ZN(n548) );
  XNOR2_X1 U606 ( .A(KEYINPUT66), .B(n525), .ZN(n669) );
  NAND2_X1 U607 ( .A1(G52), .A2(n667), .ZN(n547) );
  NAND2_X1 U608 ( .A1(n548), .A2(n547), .ZN(n554) );
  NAND2_X1 U609 ( .A1(G77), .A2(n659), .ZN(n551) );
  NAND2_X1 U610 ( .A1(G90), .A2(n660), .ZN(n550) );
  NAND2_X1 U611 ( .A1(n551), .A2(n550), .ZN(n552) );
  XOR2_X1 U612 ( .A(KEYINPUT9), .B(n552), .Z(n553) );
  NOR2_X1 U613 ( .A1(n554), .A2(n553), .ZN(G171) );
  XOR2_X1 U614 ( .A(KEYINPUT101), .B(KEYINPUT103), .Z(n556) );
  XNOR2_X1 U615 ( .A(G2446), .B(G2451), .ZN(n555) );
  XNOR2_X1 U616 ( .A(n556), .B(n555), .ZN(n557) );
  XOR2_X1 U617 ( .A(n557), .B(KEYINPUT102), .Z(n559) );
  XNOR2_X1 U618 ( .A(G1348), .B(G1341), .ZN(n558) );
  XNOR2_X1 U619 ( .A(n559), .B(n558), .ZN(n563) );
  XOR2_X1 U620 ( .A(G2435), .B(G2438), .Z(n561) );
  XNOR2_X1 U621 ( .A(G2454), .B(G2430), .ZN(n560) );
  XNOR2_X1 U622 ( .A(n561), .B(n560), .ZN(n562) );
  XOR2_X1 U623 ( .A(n563), .B(n562), .Z(n565) );
  XNOR2_X1 U624 ( .A(G2443), .B(G2427), .ZN(n564) );
  XNOR2_X1 U625 ( .A(n565), .B(n564), .ZN(n566) );
  AND2_X1 U626 ( .A1(n566), .A2(G14), .ZN(G401) );
  NAND2_X1 U627 ( .A1(G123), .A2(n524), .ZN(n567) );
  XNOR2_X1 U628 ( .A(n567), .B(KEYINPUT18), .ZN(n569) );
  NAND2_X1 U629 ( .A1(n882), .A2(G99), .ZN(n568) );
  NAND2_X1 U630 ( .A1(n569), .A2(n568), .ZN(n573) );
  NAND2_X1 U631 ( .A1(G135), .A2(n881), .ZN(n571) );
  NAND2_X1 U632 ( .A1(G111), .A2(n886), .ZN(n570) );
  NAND2_X1 U633 ( .A1(n571), .A2(n570), .ZN(n572) );
  NOR2_X1 U634 ( .A1(n573), .A2(n572), .ZN(n987) );
  XNOR2_X1 U635 ( .A(n987), .B(G2096), .ZN(n574) );
  XNOR2_X1 U636 ( .A(n574), .B(KEYINPUT81), .ZN(n575) );
  OR2_X1 U637 ( .A1(G2100), .A2(n575), .ZN(G156) );
  INV_X1 U638 ( .A(G132), .ZN(G219) );
  INV_X1 U639 ( .A(G82), .ZN(G220) );
  INV_X1 U640 ( .A(G57), .ZN(G237) );
  NAND2_X1 U641 ( .A1(G63), .A2(n673), .ZN(n577) );
  NAND2_X1 U642 ( .A1(G51), .A2(n667), .ZN(n576) );
  NAND2_X1 U643 ( .A1(n577), .A2(n576), .ZN(n578) );
  XNOR2_X1 U644 ( .A(KEYINPUT6), .B(n578), .ZN(n585) );
  NAND2_X1 U645 ( .A1(n660), .A2(G89), .ZN(n579) );
  XNOR2_X1 U646 ( .A(n579), .B(KEYINPUT4), .ZN(n581) );
  NAND2_X1 U647 ( .A1(G76), .A2(n659), .ZN(n580) );
  NAND2_X1 U648 ( .A1(n581), .A2(n580), .ZN(n582) );
  XOR2_X1 U649 ( .A(KEYINPUT5), .B(n582), .Z(n583) );
  XNOR2_X1 U650 ( .A(KEYINPUT76), .B(n583), .ZN(n584) );
  NOR2_X1 U651 ( .A1(n585), .A2(n584), .ZN(n587) );
  XNOR2_X1 U652 ( .A(KEYINPUT77), .B(KEYINPUT7), .ZN(n586) );
  XNOR2_X1 U653 ( .A(n587), .B(n586), .ZN(G168) );
  XOR2_X1 U654 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U655 ( .A1(G94), .A2(G452), .ZN(n588) );
  XNOR2_X1 U656 ( .A(n588), .B(KEYINPUT69), .ZN(G173) );
  NAND2_X1 U657 ( .A1(G7), .A2(G661), .ZN(n589) );
  XNOR2_X1 U658 ( .A(n589), .B(KEYINPUT10), .ZN(G223) );
  XNOR2_X1 U659 ( .A(G223), .B(KEYINPUT71), .ZN(n849) );
  NAND2_X1 U660 ( .A1(n849), .A2(G567), .ZN(n590) );
  XOR2_X1 U661 ( .A(KEYINPUT11), .B(n590), .Z(G234) );
  NAND2_X1 U662 ( .A1(G56), .A2(n673), .ZN(n591) );
  XOR2_X1 U663 ( .A(KEYINPUT14), .B(n591), .Z(n597) );
  NAND2_X1 U664 ( .A1(n660), .A2(G81), .ZN(n592) );
  XNOR2_X1 U665 ( .A(n592), .B(KEYINPUT12), .ZN(n594) );
  NAND2_X1 U666 ( .A1(G68), .A2(n659), .ZN(n593) );
  NAND2_X1 U667 ( .A1(n594), .A2(n593), .ZN(n595) );
  XOR2_X1 U668 ( .A(KEYINPUT13), .B(n595), .Z(n596) );
  NOR2_X1 U669 ( .A1(n597), .A2(n596), .ZN(n599) );
  NAND2_X1 U670 ( .A1(n667), .A2(G43), .ZN(n598) );
  NAND2_X1 U671 ( .A1(n599), .A2(n598), .ZN(n932) );
  INV_X1 U672 ( .A(G860), .ZN(n625) );
  NOR2_X1 U673 ( .A1(n932), .A2(n625), .ZN(n600) );
  XOR2_X1 U674 ( .A(KEYINPUT72), .B(n600), .Z(G153) );
  NAND2_X1 U675 ( .A1(G868), .A2(G171), .ZN(n611) );
  NAND2_X1 U676 ( .A1(G54), .A2(n667), .ZN(n601) );
  XNOR2_X1 U677 ( .A(n601), .B(KEYINPUT74), .ZN(n608) );
  NAND2_X1 U678 ( .A1(G66), .A2(n673), .ZN(n603) );
  NAND2_X1 U679 ( .A1(G92), .A2(n660), .ZN(n602) );
  NAND2_X1 U680 ( .A1(n603), .A2(n602), .ZN(n606) );
  NAND2_X1 U681 ( .A1(G79), .A2(n659), .ZN(n604) );
  XNOR2_X1 U682 ( .A(KEYINPUT73), .B(n604), .ZN(n605) );
  NOR2_X1 U683 ( .A1(n606), .A2(n605), .ZN(n607) );
  NAND2_X1 U684 ( .A1(n608), .A2(n607), .ZN(n609) );
  INV_X1 U685 ( .A(n953), .ZN(n632) );
  INV_X1 U686 ( .A(G868), .ZN(n621) );
  NAND2_X1 U687 ( .A1(n632), .A2(n621), .ZN(n610) );
  NAND2_X1 U688 ( .A1(n611), .A2(n610), .ZN(n612) );
  XNOR2_X1 U689 ( .A(n612), .B(KEYINPUT75), .ZN(G284) );
  NAND2_X1 U690 ( .A1(G65), .A2(n673), .ZN(n614) );
  NAND2_X1 U691 ( .A1(G91), .A2(n660), .ZN(n613) );
  NAND2_X1 U692 ( .A1(n614), .A2(n613), .ZN(n617) );
  NAND2_X1 U693 ( .A1(n659), .A2(G78), .ZN(n615) );
  XOR2_X1 U694 ( .A(KEYINPUT70), .B(n615), .Z(n616) );
  NOR2_X1 U695 ( .A1(n617), .A2(n616), .ZN(n619) );
  NAND2_X1 U696 ( .A1(n667), .A2(G53), .ZN(n618) );
  NAND2_X1 U697 ( .A1(n619), .A2(n618), .ZN(G299) );
  NOR2_X1 U698 ( .A1(G868), .A2(G299), .ZN(n620) );
  XNOR2_X1 U699 ( .A(n620), .B(KEYINPUT78), .ZN(n623) );
  NOR2_X1 U700 ( .A1(n621), .A2(G286), .ZN(n622) );
  NOR2_X1 U701 ( .A1(n623), .A2(n622), .ZN(n624) );
  XOR2_X1 U702 ( .A(KEYINPUT79), .B(n624), .Z(G297) );
  NAND2_X1 U703 ( .A1(n625), .A2(G559), .ZN(n626) );
  NAND2_X1 U704 ( .A1(n626), .A2(n632), .ZN(n627) );
  XNOR2_X1 U705 ( .A(n627), .B(KEYINPUT16), .ZN(n628) );
  XNOR2_X1 U706 ( .A(KEYINPUT80), .B(n628), .ZN(G148) );
  NOR2_X1 U707 ( .A1(G868), .A2(n932), .ZN(n631) );
  NAND2_X1 U708 ( .A1(G868), .A2(n632), .ZN(n629) );
  NOR2_X1 U709 ( .A1(G559), .A2(n629), .ZN(n630) );
  NOR2_X1 U710 ( .A1(n631), .A2(n630), .ZN(G282) );
  NAND2_X1 U711 ( .A1(n632), .A2(G559), .ZN(n682) );
  XNOR2_X1 U712 ( .A(n932), .B(n682), .ZN(n633) );
  NOR2_X1 U713 ( .A1(n633), .A2(G860), .ZN(n640) );
  NAND2_X1 U714 ( .A1(G67), .A2(n673), .ZN(n635) );
  NAND2_X1 U715 ( .A1(G93), .A2(n660), .ZN(n634) );
  NAND2_X1 U716 ( .A1(n635), .A2(n634), .ZN(n639) );
  NAND2_X1 U717 ( .A1(G55), .A2(n667), .ZN(n637) );
  NAND2_X1 U718 ( .A1(G80), .A2(n659), .ZN(n636) );
  NAND2_X1 U719 ( .A1(n637), .A2(n636), .ZN(n638) );
  NOR2_X1 U720 ( .A1(n639), .A2(n638), .ZN(n684) );
  XNOR2_X1 U721 ( .A(n640), .B(n684), .ZN(G145) );
  NAND2_X1 U722 ( .A1(G61), .A2(n673), .ZN(n642) );
  NAND2_X1 U723 ( .A1(G86), .A2(n660), .ZN(n641) );
  NAND2_X1 U724 ( .A1(n642), .A2(n641), .ZN(n643) );
  XNOR2_X1 U725 ( .A(n643), .B(KEYINPUT83), .ZN(n645) );
  NAND2_X1 U726 ( .A1(G48), .A2(n667), .ZN(n644) );
  NAND2_X1 U727 ( .A1(n645), .A2(n644), .ZN(n649) );
  XOR2_X1 U728 ( .A(KEYINPUT84), .B(KEYINPUT2), .Z(n647) );
  NAND2_X1 U729 ( .A1(G73), .A2(n659), .ZN(n646) );
  XNOR2_X1 U730 ( .A(n647), .B(n646), .ZN(n648) );
  NOR2_X1 U731 ( .A1(n649), .A2(n648), .ZN(n650) );
  XNOR2_X1 U732 ( .A(n650), .B(KEYINPUT85), .ZN(G305) );
  NAND2_X1 U733 ( .A1(n667), .A2(G47), .ZN(n652) );
  NAND2_X1 U734 ( .A1(n673), .A2(G60), .ZN(n651) );
  NAND2_X1 U735 ( .A1(n652), .A2(n651), .ZN(n653) );
  XNOR2_X1 U736 ( .A(KEYINPUT68), .B(n653), .ZN(n656) );
  NAND2_X1 U737 ( .A1(G72), .A2(n659), .ZN(n654) );
  XNOR2_X1 U738 ( .A(KEYINPUT67), .B(n654), .ZN(n655) );
  NOR2_X1 U739 ( .A1(n656), .A2(n655), .ZN(n658) );
  NAND2_X1 U740 ( .A1(n660), .A2(G85), .ZN(n657) );
  NAND2_X1 U741 ( .A1(n658), .A2(n657), .ZN(G290) );
  NAND2_X1 U742 ( .A1(G75), .A2(n659), .ZN(n662) );
  NAND2_X1 U743 ( .A1(G88), .A2(n660), .ZN(n661) );
  NAND2_X1 U744 ( .A1(n662), .A2(n661), .ZN(n666) );
  NAND2_X1 U745 ( .A1(G62), .A2(n673), .ZN(n664) );
  NAND2_X1 U746 ( .A1(G50), .A2(n667), .ZN(n663) );
  NAND2_X1 U747 ( .A1(n664), .A2(n663), .ZN(n665) );
  NOR2_X1 U748 ( .A1(n666), .A2(n665), .ZN(G166) );
  NAND2_X1 U749 ( .A1(G49), .A2(n667), .ZN(n668) );
  XNOR2_X1 U750 ( .A(n668), .B(KEYINPUT82), .ZN(n675) );
  NAND2_X1 U751 ( .A1(G651), .A2(G74), .ZN(n671) );
  NAND2_X1 U752 ( .A1(G87), .A2(n669), .ZN(n670) );
  NAND2_X1 U753 ( .A1(n671), .A2(n670), .ZN(n672) );
  NOR2_X1 U754 ( .A1(n673), .A2(n672), .ZN(n674) );
  NAND2_X1 U755 ( .A1(n675), .A2(n674), .ZN(G288) );
  INV_X1 U756 ( .A(G299), .ZN(n935) );
  XNOR2_X1 U757 ( .A(n935), .B(n684), .ZN(n680) );
  XNOR2_X1 U758 ( .A(G290), .B(n932), .ZN(n678) );
  XNOR2_X1 U759 ( .A(G166), .B(KEYINPUT19), .ZN(n676) );
  XNOR2_X1 U760 ( .A(n676), .B(G288), .ZN(n677) );
  XNOR2_X1 U761 ( .A(n678), .B(n677), .ZN(n679) );
  XNOR2_X1 U762 ( .A(n680), .B(n679), .ZN(n681) );
  XNOR2_X1 U763 ( .A(G305), .B(n681), .ZN(n854) );
  XNOR2_X1 U764 ( .A(n682), .B(n854), .ZN(n683) );
  NAND2_X1 U765 ( .A1(n683), .A2(G868), .ZN(n686) );
  OR2_X1 U766 ( .A1(n684), .A2(G868), .ZN(n685) );
  NAND2_X1 U767 ( .A1(n686), .A2(n685), .ZN(G295) );
  NAND2_X1 U768 ( .A1(G2078), .A2(G2084), .ZN(n687) );
  XOR2_X1 U769 ( .A(KEYINPUT20), .B(n687), .Z(n688) );
  NAND2_X1 U770 ( .A1(G2090), .A2(n688), .ZN(n689) );
  XNOR2_X1 U771 ( .A(KEYINPUT21), .B(n689), .ZN(n690) );
  NAND2_X1 U772 ( .A1(n690), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U773 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NAND2_X1 U774 ( .A1(G120), .A2(G69), .ZN(n691) );
  NOR2_X1 U775 ( .A1(G237), .A2(n691), .ZN(n692) );
  XNOR2_X1 U776 ( .A(KEYINPUT86), .B(n692), .ZN(n693) );
  NAND2_X1 U777 ( .A1(n693), .A2(G108), .ZN(n903) );
  NAND2_X1 U778 ( .A1(n903), .A2(G567), .ZN(n698) );
  NOR2_X1 U779 ( .A1(G220), .A2(G219), .ZN(n694) );
  XOR2_X1 U780 ( .A(KEYINPUT22), .B(n694), .Z(n695) );
  NOR2_X1 U781 ( .A1(G218), .A2(n695), .ZN(n696) );
  NAND2_X1 U782 ( .A1(G96), .A2(n696), .ZN(n904) );
  NAND2_X1 U783 ( .A1(n904), .A2(G2106), .ZN(n697) );
  NAND2_X1 U784 ( .A1(n698), .A2(n697), .ZN(n905) );
  NAND2_X1 U785 ( .A1(G483), .A2(G661), .ZN(n699) );
  NOR2_X1 U786 ( .A1(n905), .A2(n699), .ZN(n853) );
  NAND2_X1 U787 ( .A1(n853), .A2(G36), .ZN(G176) );
  XNOR2_X1 U788 ( .A(KEYINPUT87), .B(G166), .ZN(G303) );
  NAND2_X1 U789 ( .A1(G160), .A2(G40), .ZN(n801) );
  NAND2_X1 U790 ( .A1(n735), .A2(G1956), .ZN(n703) );
  AND2_X1 U791 ( .A1(n706), .A2(n802), .ZN(n700) );
  AND2_X1 U792 ( .A1(n700), .A2(G2072), .ZN(n701) );
  XNOR2_X1 U793 ( .A(KEYINPUT27), .B(n701), .ZN(n702) );
  NAND2_X1 U794 ( .A1(n703), .A2(n702), .ZN(n704) );
  XNOR2_X1 U795 ( .A(n704), .B(KEYINPUT93), .ZN(n713) );
  NAND2_X1 U796 ( .A1(n935), .A2(n713), .ZN(n723) );
  INV_X1 U797 ( .A(n723), .ZN(n712) );
  AND2_X1 U798 ( .A1(G160), .A2(G40), .ZN(n706) );
  AND2_X1 U799 ( .A1(G1996), .A2(n802), .ZN(n705) );
  NAND2_X1 U800 ( .A1(n706), .A2(n705), .ZN(n707) );
  XOR2_X1 U801 ( .A(n707), .B(KEYINPUT26), .Z(n708) );
  NOR2_X1 U802 ( .A1(n932), .A2(n708), .ZN(n710) );
  NAND2_X1 U803 ( .A1(G1341), .A2(n735), .ZN(n709) );
  NAND2_X1 U804 ( .A1(n710), .A2(n709), .ZN(n717) );
  NAND2_X1 U805 ( .A1(n953), .A2(n717), .ZN(n711) );
  OR2_X1 U806 ( .A1(n712), .A2(n711), .ZN(n716) );
  NOR2_X1 U807 ( .A1(n713), .A2(n935), .ZN(n714) );
  XOR2_X1 U808 ( .A(n714), .B(KEYINPUT28), .Z(n715) );
  AND2_X1 U809 ( .A1(n716), .A2(n715), .ZN(n727) );
  XOR2_X1 U810 ( .A(KEYINPUT94), .B(n718), .Z(n725) );
  NAND2_X1 U811 ( .A1(G1348), .A2(n735), .ZN(n720) );
  NAND2_X1 U812 ( .A1(G2067), .A2(n700), .ZN(n719) );
  NAND2_X1 U813 ( .A1(n720), .A2(n719), .ZN(n721) );
  XOR2_X1 U814 ( .A(KEYINPUT95), .B(n721), .Z(n722) );
  AND2_X1 U815 ( .A1(n723), .A2(n722), .ZN(n724) );
  NAND2_X1 U816 ( .A1(n725), .A2(n724), .ZN(n726) );
  NAND2_X1 U817 ( .A1(n727), .A2(n726), .ZN(n729) );
  XNOR2_X1 U818 ( .A(G2078), .B(KEYINPUT25), .ZN(n969) );
  NAND2_X1 U819 ( .A1(n700), .A2(n969), .ZN(n730) );
  XNOR2_X1 U820 ( .A(n730), .B(KEYINPUT92), .ZN(n732) );
  OR2_X1 U821 ( .A1(G1961), .A2(n700), .ZN(n731) );
  NAND2_X1 U822 ( .A1(n732), .A2(n731), .ZN(n741) );
  NAND2_X1 U823 ( .A1(n741), .A2(G171), .ZN(n733) );
  NAND2_X1 U824 ( .A1(n734), .A2(n733), .ZN(n758) );
  INV_X1 U825 ( .A(G1966), .ZN(n737) );
  NAND2_X1 U826 ( .A1(n735), .A2(G8), .ZN(n736) );
  AND2_X1 U827 ( .A1(n737), .A2(n787), .ZN(n760) );
  NOR2_X1 U828 ( .A1(G2084), .A2(n735), .ZN(n761) );
  NOR2_X1 U829 ( .A1(n760), .A2(n761), .ZN(n738) );
  NAND2_X1 U830 ( .A1(G8), .A2(n738), .ZN(n739) );
  XNOR2_X1 U831 ( .A(KEYINPUT30), .B(n739), .ZN(n740) );
  NOR2_X1 U832 ( .A1(G168), .A2(n740), .ZN(n743) );
  NOR2_X1 U833 ( .A1(G171), .A2(n741), .ZN(n742) );
  INV_X1 U834 ( .A(n787), .ZN(n773) );
  NOR2_X1 U835 ( .A1(G1971), .A2(n773), .ZN(n747) );
  NOR2_X1 U836 ( .A1(G2090), .A2(n735), .ZN(n746) );
  NOR2_X1 U837 ( .A1(n747), .A2(n746), .ZN(n748) );
  XOR2_X1 U838 ( .A(KEYINPUT97), .B(n748), .Z(n749) );
  NAND2_X1 U839 ( .A1(n749), .A2(G303), .ZN(n751) );
  NAND2_X1 U840 ( .A1(n758), .A2(n750), .ZN(n754) );
  INV_X1 U841 ( .A(n751), .ZN(n752) );
  OR2_X1 U842 ( .A1(n752), .A2(G286), .ZN(n753) );
  NAND2_X1 U843 ( .A1(G8), .A2(n755), .ZN(n756) );
  XNOR2_X1 U844 ( .A(n756), .B(KEYINPUT32), .ZN(n792) );
  NAND2_X1 U845 ( .A1(G1976), .A2(G288), .ZN(n936) );
  AND2_X1 U846 ( .A1(n787), .A2(n936), .ZN(n766) );
  AND2_X1 U847 ( .A1(n758), .A2(n757), .ZN(n759) );
  NAND2_X1 U848 ( .A1(G8), .A2(n761), .ZN(n762) );
  NAND2_X1 U849 ( .A1(n763), .A2(n762), .ZN(n764) );
  XNOR2_X1 U850 ( .A(KEYINPUT96), .B(n764), .ZN(n791) );
  NAND2_X1 U851 ( .A1(n765), .A2(n791), .ZN(n771) );
  INV_X1 U852 ( .A(n766), .ZN(n769) );
  NOR2_X1 U853 ( .A1(G1971), .A2(G303), .ZN(n767) );
  NOR2_X1 U854 ( .A1(G1976), .A2(G288), .ZN(n778) );
  NOR2_X1 U855 ( .A1(n767), .A2(n778), .ZN(n768) );
  OR2_X1 U856 ( .A1(n769), .A2(n768), .ZN(n770) );
  NAND2_X1 U857 ( .A1(n771), .A2(n770), .ZN(n772) );
  XNOR2_X1 U858 ( .A(n772), .B(KEYINPUT64), .ZN(n774) );
  AND2_X1 U859 ( .A1(n774), .A2(n527), .ZN(n775) );
  NOR2_X1 U860 ( .A1(KEYINPUT33), .A2(n775), .ZN(n776) );
  INV_X1 U861 ( .A(n776), .ZN(n785) );
  NAND2_X1 U862 ( .A1(n778), .A2(KEYINPUT33), .ZN(n777) );
  AND2_X1 U863 ( .A1(n777), .A2(KEYINPUT98), .ZN(n780) );
  INV_X1 U864 ( .A(n778), .ZN(n937) );
  NOR2_X1 U865 ( .A1(KEYINPUT98), .A2(n937), .ZN(n779) );
  NOR2_X1 U866 ( .A1(n780), .A2(n779), .ZN(n781) );
  NAND2_X1 U867 ( .A1(n781), .A2(n787), .ZN(n784) );
  OR2_X1 U868 ( .A1(G1981), .A2(G305), .ZN(n786) );
  NAND2_X1 U869 ( .A1(G1981), .A2(G305), .ZN(n782) );
  NAND2_X1 U870 ( .A1(n786), .A2(n782), .ZN(n950) );
  NAND2_X1 U871 ( .A1(n785), .A2(n526), .ZN(n790) );
  XOR2_X1 U872 ( .A(n786), .B(KEYINPUT24), .Z(n788) );
  NAND2_X1 U873 ( .A1(n788), .A2(n787), .ZN(n789) );
  NAND2_X1 U874 ( .A1(n790), .A2(n789), .ZN(n799) );
  AND2_X1 U875 ( .A1(n792), .A2(n791), .ZN(n796) );
  NOR2_X1 U876 ( .A1(G2090), .A2(G303), .ZN(n793) );
  NAND2_X1 U877 ( .A1(G8), .A2(n793), .ZN(n794) );
  XNOR2_X1 U878 ( .A(KEYINPUT99), .B(n794), .ZN(n795) );
  NOR2_X1 U879 ( .A1(n796), .A2(n795), .ZN(n797) );
  NOR2_X1 U880 ( .A1(n787), .A2(n797), .ZN(n798) );
  NOR2_X1 U881 ( .A1(n799), .A2(n798), .ZN(n800) );
  INV_X1 U882 ( .A(n800), .ZN(n833) );
  XNOR2_X1 U883 ( .A(G1986), .B(G290), .ZN(n945) );
  NOR2_X1 U884 ( .A1(n802), .A2(n801), .ZN(n844) );
  NAND2_X1 U885 ( .A1(G140), .A2(n881), .ZN(n804) );
  NAND2_X1 U886 ( .A1(G104), .A2(n882), .ZN(n803) );
  NAND2_X1 U887 ( .A1(n804), .A2(n803), .ZN(n805) );
  XNOR2_X1 U888 ( .A(KEYINPUT34), .B(n805), .ZN(n810) );
  NAND2_X1 U889 ( .A1(G128), .A2(n524), .ZN(n807) );
  NAND2_X1 U890 ( .A1(G116), .A2(n886), .ZN(n806) );
  NAND2_X1 U891 ( .A1(n807), .A2(n806), .ZN(n808) );
  XOR2_X1 U892 ( .A(KEYINPUT35), .B(n808), .Z(n809) );
  NOR2_X1 U893 ( .A1(n810), .A2(n809), .ZN(n811) );
  XNOR2_X1 U894 ( .A(KEYINPUT36), .B(n811), .ZN(n900) );
  XNOR2_X1 U895 ( .A(KEYINPUT37), .B(G2067), .ZN(n834) );
  NOR2_X1 U896 ( .A1(n900), .A2(n834), .ZN(n988) );
  NAND2_X1 U897 ( .A1(n844), .A2(n988), .ZN(n842) );
  NAND2_X1 U898 ( .A1(G131), .A2(n881), .ZN(n813) );
  NAND2_X1 U899 ( .A1(G95), .A2(n882), .ZN(n812) );
  NAND2_X1 U900 ( .A1(n813), .A2(n812), .ZN(n814) );
  XNOR2_X1 U901 ( .A(KEYINPUT88), .B(n814), .ZN(n818) );
  NAND2_X1 U902 ( .A1(G119), .A2(n524), .ZN(n816) );
  NAND2_X1 U903 ( .A1(G107), .A2(n886), .ZN(n815) );
  NAND2_X1 U904 ( .A1(n816), .A2(n815), .ZN(n817) );
  NOR2_X1 U905 ( .A1(n818), .A2(n817), .ZN(n893) );
  INV_X1 U906 ( .A(G1991), .ZN(n963) );
  NOR2_X1 U907 ( .A1(n893), .A2(n963), .ZN(n829) );
  NAND2_X1 U908 ( .A1(G129), .A2(n524), .ZN(n820) );
  NAND2_X1 U909 ( .A1(G117), .A2(n886), .ZN(n819) );
  NAND2_X1 U910 ( .A1(n820), .A2(n819), .ZN(n824) );
  NAND2_X1 U911 ( .A1(G105), .A2(n882), .ZN(n821) );
  XNOR2_X1 U912 ( .A(n821), .B(KEYINPUT89), .ZN(n822) );
  XNOR2_X1 U913 ( .A(n822), .B(KEYINPUT38), .ZN(n823) );
  NOR2_X1 U914 ( .A1(n824), .A2(n823), .ZN(n825) );
  XNOR2_X1 U915 ( .A(n825), .B(KEYINPUT90), .ZN(n827) );
  NAND2_X1 U916 ( .A1(G141), .A2(n881), .ZN(n826) );
  NAND2_X1 U917 ( .A1(n827), .A2(n826), .ZN(n897) );
  AND2_X1 U918 ( .A1(n897), .A2(G1996), .ZN(n828) );
  NOR2_X1 U919 ( .A1(n829), .A2(n828), .ZN(n993) );
  INV_X1 U920 ( .A(n844), .ZN(n830) );
  NOR2_X1 U921 ( .A1(n993), .A2(n830), .ZN(n837) );
  INV_X1 U922 ( .A(n837), .ZN(n831) );
  NAND2_X1 U923 ( .A1(n842), .A2(n831), .ZN(n832) );
  NAND2_X1 U924 ( .A1(n833), .A2(n528), .ZN(n847) );
  NAND2_X1 U925 ( .A1(n900), .A2(n834), .ZN(n992) );
  XOR2_X1 U926 ( .A(KEYINPUT39), .B(KEYINPUT100), .Z(n840) );
  NOR2_X1 U927 ( .A1(G1996), .A2(n897), .ZN(n1004) );
  NOR2_X1 U928 ( .A1(G1986), .A2(G290), .ZN(n835) );
  AND2_X1 U929 ( .A1(n963), .A2(n893), .ZN(n986) );
  NOR2_X1 U930 ( .A1(n835), .A2(n986), .ZN(n836) );
  NOR2_X1 U931 ( .A1(n837), .A2(n836), .ZN(n838) );
  NOR2_X1 U932 ( .A1(n1004), .A2(n838), .ZN(n839) );
  XOR2_X1 U933 ( .A(n840), .B(n839), .Z(n841) );
  NAND2_X1 U934 ( .A1(n842), .A2(n841), .ZN(n843) );
  NAND2_X1 U935 ( .A1(n992), .A2(n843), .ZN(n845) );
  NAND2_X1 U936 ( .A1(n845), .A2(n844), .ZN(n846) );
  NAND2_X1 U937 ( .A1(n847), .A2(n846), .ZN(n848) );
  XNOR2_X1 U938 ( .A(KEYINPUT40), .B(n848), .ZN(G329) );
  NAND2_X1 U939 ( .A1(n849), .A2(G2106), .ZN(n850) );
  XNOR2_X1 U940 ( .A(n850), .B(KEYINPUT104), .ZN(G217) );
  AND2_X1 U941 ( .A1(G15), .A2(G2), .ZN(n851) );
  NAND2_X1 U942 ( .A1(G661), .A2(n851), .ZN(G259) );
  NAND2_X1 U943 ( .A1(G3), .A2(G1), .ZN(n852) );
  NAND2_X1 U944 ( .A1(n853), .A2(n852), .ZN(G188) );
  XNOR2_X1 U945 ( .A(G286), .B(n953), .ZN(n855) );
  XNOR2_X1 U946 ( .A(n855), .B(n854), .ZN(n856) );
  XNOR2_X1 U947 ( .A(n856), .B(G171), .ZN(n857) );
  NOR2_X1 U948 ( .A1(G37), .A2(n857), .ZN(G397) );
  XOR2_X1 U949 ( .A(KEYINPUT44), .B(KEYINPUT108), .Z(n859) );
  NAND2_X1 U950 ( .A1(G124), .A2(n524), .ZN(n858) );
  XNOR2_X1 U951 ( .A(n859), .B(n858), .ZN(n860) );
  XNOR2_X1 U952 ( .A(n860), .B(KEYINPUT107), .ZN(n862) );
  NAND2_X1 U953 ( .A1(n882), .A2(G100), .ZN(n861) );
  NAND2_X1 U954 ( .A1(n862), .A2(n861), .ZN(n866) );
  NAND2_X1 U955 ( .A1(G136), .A2(n881), .ZN(n864) );
  NAND2_X1 U956 ( .A1(G112), .A2(n886), .ZN(n863) );
  NAND2_X1 U957 ( .A1(n864), .A2(n863), .ZN(n865) );
  NOR2_X1 U958 ( .A1(n866), .A2(n865), .ZN(G162) );
  XOR2_X1 U959 ( .A(KEYINPUT46), .B(KEYINPUT48), .Z(n877) );
  NAND2_X1 U960 ( .A1(G130), .A2(n524), .ZN(n868) );
  NAND2_X1 U961 ( .A1(G118), .A2(n886), .ZN(n867) );
  NAND2_X1 U962 ( .A1(n868), .A2(n867), .ZN(n874) );
  NAND2_X1 U963 ( .A1(G142), .A2(n881), .ZN(n870) );
  NAND2_X1 U964 ( .A1(G106), .A2(n882), .ZN(n869) );
  NAND2_X1 U965 ( .A1(n870), .A2(n869), .ZN(n871) );
  XNOR2_X1 U966 ( .A(KEYINPUT109), .B(n871), .ZN(n872) );
  XNOR2_X1 U967 ( .A(KEYINPUT45), .B(n872), .ZN(n873) );
  NOR2_X1 U968 ( .A1(n874), .A2(n873), .ZN(n875) );
  XNOR2_X1 U969 ( .A(n875), .B(KEYINPUT111), .ZN(n876) );
  XNOR2_X1 U970 ( .A(n877), .B(n876), .ZN(n878) );
  XOR2_X1 U971 ( .A(n878), .B(KEYINPUT112), .Z(n880) );
  XNOR2_X1 U972 ( .A(G164), .B(KEYINPUT110), .ZN(n879) );
  XNOR2_X1 U973 ( .A(n880), .B(n879), .ZN(n892) );
  NAND2_X1 U974 ( .A1(G139), .A2(n881), .ZN(n884) );
  NAND2_X1 U975 ( .A1(G103), .A2(n882), .ZN(n883) );
  NAND2_X1 U976 ( .A1(n884), .A2(n883), .ZN(n891) );
  NAND2_X1 U977 ( .A1(G127), .A2(n524), .ZN(n888) );
  NAND2_X1 U978 ( .A1(G115), .A2(n886), .ZN(n887) );
  NAND2_X1 U979 ( .A1(n888), .A2(n887), .ZN(n889) );
  XOR2_X1 U980 ( .A(KEYINPUT47), .B(n889), .Z(n890) );
  NOR2_X1 U981 ( .A1(n891), .A2(n890), .ZN(n994) );
  XOR2_X1 U982 ( .A(n892), .B(n994), .Z(n895) );
  XNOR2_X1 U983 ( .A(n893), .B(G162), .ZN(n894) );
  XNOR2_X1 U984 ( .A(n895), .B(n894), .ZN(n896) );
  XOR2_X1 U985 ( .A(n896), .B(n987), .Z(n899) );
  XOR2_X1 U986 ( .A(G160), .B(n897), .Z(n898) );
  XNOR2_X1 U987 ( .A(n899), .B(n898), .ZN(n901) );
  XOR2_X1 U988 ( .A(n901), .B(n900), .Z(n902) );
  NOR2_X1 U989 ( .A1(G37), .A2(n902), .ZN(G395) );
  INV_X1 U991 ( .A(G120), .ZN(G236) );
  INV_X1 U992 ( .A(G108), .ZN(G238) );
  INV_X1 U993 ( .A(G96), .ZN(G221) );
  INV_X1 U994 ( .A(G69), .ZN(G235) );
  NOR2_X1 U995 ( .A1(n904), .A2(n903), .ZN(G325) );
  INV_X1 U996 ( .A(G325), .ZN(G261) );
  INV_X1 U997 ( .A(n905), .ZN(G319) );
  XOR2_X1 U998 ( .A(KEYINPUT106), .B(KEYINPUT105), .Z(n907) );
  XNOR2_X1 U999 ( .A(G2678), .B(KEYINPUT43), .ZN(n906) );
  XNOR2_X1 U1000 ( .A(n907), .B(n906), .ZN(n911) );
  XOR2_X1 U1001 ( .A(KEYINPUT42), .B(G2090), .Z(n909) );
  XNOR2_X1 U1002 ( .A(G2067), .B(G2072), .ZN(n908) );
  XNOR2_X1 U1003 ( .A(n909), .B(n908), .ZN(n910) );
  XOR2_X1 U1004 ( .A(n911), .B(n910), .Z(n913) );
  XNOR2_X1 U1005 ( .A(G2096), .B(G2100), .ZN(n912) );
  XNOR2_X1 U1006 ( .A(n913), .B(n912), .ZN(n915) );
  XOR2_X1 U1007 ( .A(G2078), .B(G2084), .Z(n914) );
  XNOR2_X1 U1008 ( .A(n915), .B(n914), .ZN(G227) );
  XOR2_X1 U1009 ( .A(G1971), .B(G1961), .Z(n917) );
  XNOR2_X1 U1010 ( .A(G1986), .B(G1966), .ZN(n916) );
  XNOR2_X1 U1011 ( .A(n917), .B(n916), .ZN(n918) );
  XOR2_X1 U1012 ( .A(n918), .B(KEYINPUT41), .Z(n920) );
  XNOR2_X1 U1013 ( .A(G1956), .B(G1981), .ZN(n919) );
  XNOR2_X1 U1014 ( .A(n920), .B(n919), .ZN(n924) );
  XOR2_X1 U1015 ( .A(G2474), .B(G1976), .Z(n922) );
  XNOR2_X1 U1016 ( .A(G1996), .B(G1991), .ZN(n921) );
  XNOR2_X1 U1017 ( .A(n922), .B(n921), .ZN(n923) );
  XNOR2_X1 U1018 ( .A(n924), .B(n923), .ZN(G229) );
  NOR2_X1 U1019 ( .A1(G227), .A2(G229), .ZN(n926) );
  XNOR2_X1 U1020 ( .A(KEYINPUT113), .B(KEYINPUT49), .ZN(n925) );
  XNOR2_X1 U1021 ( .A(n926), .B(n925), .ZN(n929) );
  NOR2_X1 U1022 ( .A1(G397), .A2(G395), .ZN(n927) );
  XNOR2_X1 U1023 ( .A(n927), .B(KEYINPUT114), .ZN(n928) );
  NAND2_X1 U1024 ( .A1(n929), .A2(n928), .ZN(n930) );
  NOR2_X1 U1025 ( .A1(G401), .A2(n930), .ZN(n931) );
  NAND2_X1 U1026 ( .A1(G319), .A2(n931), .ZN(G225) );
  INV_X1 U1027 ( .A(G225), .ZN(G308) );
  INV_X1 U1028 ( .A(G171), .ZN(G301) );
  XOR2_X1 U1029 ( .A(G16), .B(KEYINPUT56), .Z(n959) );
  XNOR2_X1 U1030 ( .A(G301), .B(G1961), .ZN(n934) );
  XNOR2_X1 U1031 ( .A(n932), .B(G1341), .ZN(n933) );
  NOR2_X1 U1032 ( .A1(n934), .A2(n933), .ZN(n948) );
  XNOR2_X1 U1033 ( .A(n935), .B(G1956), .ZN(n943) );
  NAND2_X1 U1034 ( .A1(n937), .A2(n936), .ZN(n938) );
  XOR2_X1 U1035 ( .A(KEYINPUT121), .B(n938), .Z(n941) );
  XNOR2_X1 U1036 ( .A(G1971), .B(G303), .ZN(n939) );
  XNOR2_X1 U1037 ( .A(KEYINPUT122), .B(n939), .ZN(n940) );
  NOR2_X1 U1038 ( .A1(n941), .A2(n940), .ZN(n942) );
  NAND2_X1 U1039 ( .A1(n943), .A2(n942), .ZN(n944) );
  NOR2_X1 U1040 ( .A1(n945), .A2(n944), .ZN(n946) );
  XOR2_X1 U1041 ( .A(KEYINPUT123), .B(n946), .Z(n947) );
  NAND2_X1 U1042 ( .A1(n948), .A2(n947), .ZN(n957) );
  XOR2_X1 U1043 ( .A(G168), .B(G1966), .Z(n949) );
  NOR2_X1 U1044 ( .A1(n950), .A2(n949), .ZN(n951) );
  XOR2_X1 U1045 ( .A(KEYINPUT57), .B(n951), .Z(n955) );
  XOR2_X1 U1046 ( .A(G1348), .B(KEYINPUT120), .Z(n952) );
  XNOR2_X1 U1047 ( .A(n953), .B(n952), .ZN(n954) );
  NAND2_X1 U1048 ( .A1(n955), .A2(n954), .ZN(n956) );
  NOR2_X1 U1049 ( .A1(n957), .A2(n956), .ZN(n958) );
  NOR2_X1 U1050 ( .A1(n959), .A2(n958), .ZN(n984) );
  XNOR2_X1 U1051 ( .A(KEYINPUT55), .B(KEYINPUT117), .ZN(n1009) );
  XNOR2_X1 U1052 ( .A(G1996), .B(G32), .ZN(n961) );
  XNOR2_X1 U1053 ( .A(G33), .B(G2072), .ZN(n960) );
  NOR2_X1 U1054 ( .A1(n961), .A2(n960), .ZN(n968) );
  XOR2_X1 U1055 ( .A(G2067), .B(G26), .Z(n962) );
  NAND2_X1 U1056 ( .A1(n962), .A2(G28), .ZN(n966) );
  XOR2_X1 U1057 ( .A(G25), .B(n963), .Z(n964) );
  XNOR2_X1 U1058 ( .A(KEYINPUT118), .B(n964), .ZN(n965) );
  NOR2_X1 U1059 ( .A1(n966), .A2(n965), .ZN(n967) );
  NAND2_X1 U1060 ( .A1(n968), .A2(n967), .ZN(n971) );
  XOR2_X1 U1061 ( .A(G27), .B(n969), .Z(n970) );
  NOR2_X1 U1062 ( .A1(n971), .A2(n970), .ZN(n972) );
  XOR2_X1 U1063 ( .A(KEYINPUT53), .B(n972), .Z(n975) );
  XOR2_X1 U1064 ( .A(G34), .B(KEYINPUT54), .Z(n973) );
  XNOR2_X1 U1065 ( .A(G2084), .B(n973), .ZN(n974) );
  NAND2_X1 U1066 ( .A1(n975), .A2(n974), .ZN(n977) );
  XNOR2_X1 U1067 ( .A(G35), .B(G2090), .ZN(n976) );
  NOR2_X1 U1068 ( .A1(n977), .A2(n976), .ZN(n978) );
  XOR2_X1 U1069 ( .A(n1009), .B(n978), .Z(n980) );
  INV_X1 U1070 ( .A(G29), .ZN(n979) );
  NAND2_X1 U1071 ( .A1(n980), .A2(n979), .ZN(n981) );
  NAND2_X1 U1072 ( .A1(n981), .A2(G11), .ZN(n982) );
  XOR2_X1 U1073 ( .A(KEYINPUT119), .B(n982), .Z(n983) );
  NOR2_X1 U1074 ( .A1(n984), .A2(n983), .ZN(n1013) );
  XOR2_X1 U1075 ( .A(G160), .B(G2084), .Z(n985) );
  NOR2_X1 U1076 ( .A1(n986), .A2(n985), .ZN(n990) );
  NOR2_X1 U1077 ( .A1(n988), .A2(n987), .ZN(n989) );
  NAND2_X1 U1078 ( .A1(n990), .A2(n989), .ZN(n991) );
  XNOR2_X1 U1079 ( .A(KEYINPUT115), .B(n991), .ZN(n1002) );
  NAND2_X1 U1080 ( .A1(n993), .A2(n992), .ZN(n1000) );
  XOR2_X1 U1081 ( .A(G2072), .B(n994), .Z(n996) );
  XOR2_X1 U1082 ( .A(G164), .B(G2078), .Z(n995) );
  NOR2_X1 U1083 ( .A1(n996), .A2(n995), .ZN(n997) );
  XOR2_X1 U1084 ( .A(KEYINPUT50), .B(n997), .Z(n998) );
  XNOR2_X1 U1085 ( .A(KEYINPUT116), .B(n998), .ZN(n999) );
  NOR2_X1 U1086 ( .A1(n1000), .A2(n999), .ZN(n1001) );
  NAND2_X1 U1087 ( .A1(n1002), .A2(n1001), .ZN(n1007) );
  XOR2_X1 U1088 ( .A(G2090), .B(G162), .Z(n1003) );
  NOR2_X1 U1089 ( .A1(n1004), .A2(n1003), .ZN(n1005) );
  XNOR2_X1 U1090 ( .A(n1005), .B(KEYINPUT51), .ZN(n1006) );
  NOR2_X1 U1091 ( .A1(n1007), .A2(n1006), .ZN(n1008) );
  XNOR2_X1 U1092 ( .A(KEYINPUT52), .B(n1008), .ZN(n1010) );
  NAND2_X1 U1093 ( .A1(n1010), .A2(n1009), .ZN(n1011) );
  NAND2_X1 U1094 ( .A1(n1011), .A2(G29), .ZN(n1012) );
  NAND2_X1 U1095 ( .A1(n1013), .A2(n1012), .ZN(n1040) );
  XNOR2_X1 U1096 ( .A(G1348), .B(KEYINPUT59), .ZN(n1014) );
  XNOR2_X1 U1097 ( .A(n1014), .B(G4), .ZN(n1018) );
  XNOR2_X1 U1098 ( .A(G1341), .B(G19), .ZN(n1016) );
  XNOR2_X1 U1099 ( .A(G6), .B(G1981), .ZN(n1015) );
  NOR2_X1 U1100 ( .A1(n1016), .A2(n1015), .ZN(n1017) );
  NAND2_X1 U1101 ( .A1(n1018), .A2(n1017), .ZN(n1020) );
  XNOR2_X1 U1102 ( .A(G20), .B(G1956), .ZN(n1019) );
  NOR2_X1 U1103 ( .A1(n1020), .A2(n1019), .ZN(n1021) );
  XOR2_X1 U1104 ( .A(KEYINPUT60), .B(n1021), .Z(n1023) );
  XNOR2_X1 U1105 ( .A(G1966), .B(G21), .ZN(n1022) );
  NOR2_X1 U1106 ( .A1(n1023), .A2(n1022), .ZN(n1024) );
  XOR2_X1 U1107 ( .A(KEYINPUT125), .B(n1024), .Z(n1033) );
  XOR2_X1 U1108 ( .A(G1976), .B(KEYINPUT126), .Z(n1025) );
  XNOR2_X1 U1109 ( .A(G23), .B(n1025), .ZN(n1029) );
  XNOR2_X1 U1110 ( .A(G1986), .B(G24), .ZN(n1027) );
  XNOR2_X1 U1111 ( .A(G1971), .B(G22), .ZN(n1026) );
  NOR2_X1 U1112 ( .A1(n1027), .A2(n1026), .ZN(n1028) );
  NAND2_X1 U1113 ( .A1(n1029), .A2(n1028), .ZN(n1030) );
  XNOR2_X1 U1114 ( .A(n1030), .B(KEYINPUT127), .ZN(n1031) );
  XNOR2_X1 U1115 ( .A(KEYINPUT58), .B(n1031), .ZN(n1032) );
  NAND2_X1 U1116 ( .A1(n1033), .A2(n1032), .ZN(n1035) );
  XNOR2_X1 U1117 ( .A(G5), .B(G1961), .ZN(n1034) );
  NOR2_X1 U1118 ( .A1(n1035), .A2(n1034), .ZN(n1036) );
  XOR2_X1 U1119 ( .A(KEYINPUT61), .B(n1036), .Z(n1038) );
  XNOR2_X1 U1120 ( .A(KEYINPUT124), .B(G16), .ZN(n1037) );
  NOR2_X1 U1121 ( .A1(n1038), .A2(n1037), .ZN(n1039) );
  NOR2_X1 U1122 ( .A1(n1040), .A2(n1039), .ZN(n1041) );
  XNOR2_X1 U1123 ( .A(n1041), .B(KEYINPUT62), .ZN(G311) );
  INV_X1 U1124 ( .A(G311), .ZN(G150) );
endmodule

