

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n513, n514, n515, n516,
         n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527,
         n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538,
         n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549,
         n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560,
         n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571,
         n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582,
         n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593,
         n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604,
         n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615,
         n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626,
         n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637,
         n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648,
         n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659,
         n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670,
         n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681,
         n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692,
         n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703,
         n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714,
         n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725,
         n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736,
         n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747,
         n748, n749, n750, n751, n752, n753, n754, n755, n756, n757, n758,
         n759, n760, n761, n762, n763, n764, n765, n766, n767, n768, n769,
         n770, n771, n772, n773, n774, n775, n776, n777, n778, n779, n780,
         n781, n782, n783, n784, n785, n786, n787, n788, n789, n790, n791,
         n792, n793, n794, n795, n796, n797, n798, n799, n800, n801, n802,
         n803, n804, n805, n806, n807, n808, n809, n810, n811, n812, n813,
         n814, n815, n816, n817, n818, n819, n820, n821, n822, n823, n824,
         n825, n826, n827, n828, n829, n830, n831, n832, n833, n834, n835,
         n836, n837, n838, n839, n840, n841, n842, n843, n844, n845, n846,
         n847, n848, n849, n850, n851, n852, n853, n854, n855, n856, n857,
         n858, n859, n860, n861, n862, n863, n864, n865, n866, n867, n868,
         n869, n870, n871, n872, n873, n874, n875, n876, n877, n878, n879,
         n880, n881, n882, n883, n884, n885, n886, n887, n888, n889, n890,
         n891, n892, n893, n894, n895, n896, n897, n898, n899, n900, n901,
         n902, n903, n904, n905, n906, n907, n908, n909, n910, n911, n912,
         n913, n914, n915, n916, n917, n918, n919, n920, n921, n922, n923,
         n924, n925, n926, n927, n928, n929, n930, n931, n932, n933, n934,
         n935, n936, n937, n938, n939, n940, n941, n942, n943, n944, n945,
         n946, n947, n948, n949, n950, n951, n952, n953, n954, n955, n956,
         n957, n958, n959, n960, n961, n962, n963, n964, n965, n966, n967,
         n968, n969, n970, n971, n972, n973, n974, n975, n976, n977, n978,
         n979, n980, n981, n982, n983, n984, n985, n986, n987, n988, n989,
         n990, n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000,
         n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  INV_X1 U545 ( .A(n738), .ZN(n708) );
  XOR2_X2 U546 ( .A(KEYINPUT17), .B(n515), .Z(n965) );
  NOR2_X1 U547 ( .A1(n700), .A2(n699), .ZN(n717) );
  AND2_X1 U548 ( .A1(n745), .A2(n744), .ZN(n746) );
  NOR2_X1 U549 ( .A1(KEYINPUT33), .A2(n760), .ZN(n761) );
  NOR2_X1 U550 ( .A1(G2105), .A2(G2104), .ZN(n515) );
  XOR2_X1 U551 ( .A(n719), .B(KEYINPUT28), .Z(n513) );
  NOR2_X1 U552 ( .A1(n772), .A2(n758), .ZN(n514) );
  NOR2_X1 U553 ( .A1(n738), .A2(n989), .ZN(n702) );
  NOR2_X1 U554 ( .A1(n983), .A2(n705), .ZN(n706) );
  XNOR2_X1 U555 ( .A(KEYINPUT106), .B(KEYINPUT30), .ZN(n726) );
  XNOR2_X1 U556 ( .A(n727), .B(n726), .ZN(n728) );
  INV_X1 U557 ( .A(KEYINPUT29), .ZN(n721) );
  XNOR2_X1 U558 ( .A(n722), .B(n721), .ZN(n723) );
  AND2_X1 U559 ( .A1(n759), .A2(n514), .ZN(n760) );
  OR2_X2 U560 ( .A1(n690), .A2(n777), .ZN(n738) );
  NOR2_X1 U561 ( .A1(G2105), .A2(n521), .ZN(n966) );
  NOR2_X1 U562 ( .A1(n627), .A2(G651), .ZN(n649) );
  AND2_X1 U563 ( .A1(G2105), .A2(G2104), .ZN(n961) );
  NAND2_X1 U564 ( .A1(G113), .A2(n961), .ZN(n517) );
  NAND2_X1 U565 ( .A1(G137), .A2(n965), .ZN(n516) );
  NAND2_X1 U566 ( .A1(n517), .A2(n516), .ZN(n526) );
  XNOR2_X1 U567 ( .A(KEYINPUT65), .B(G2104), .ZN(n521) );
  NAND2_X1 U568 ( .A1(n966), .A2(G101), .ZN(n520) );
  XNOR2_X1 U569 ( .A(KEYINPUT23), .B(KEYINPUT68), .ZN(n518) );
  XNOR2_X1 U570 ( .A(n518), .B(KEYINPUT67), .ZN(n519) );
  XNOR2_X1 U571 ( .A(n520), .B(n519), .ZN(n524) );
  NAND2_X1 U572 ( .A1(n521), .A2(G2105), .ZN(n522) );
  XOR2_X2 U573 ( .A(KEYINPUT66), .B(n522), .Z(n962) );
  NAND2_X1 U574 ( .A1(G125), .A2(n962), .ZN(n523) );
  NAND2_X1 U575 ( .A1(n524), .A2(n523), .ZN(n525) );
  NOR2_X2 U576 ( .A1(n526), .A2(n525), .ZN(G160) );
  NAND2_X1 U577 ( .A1(n965), .A2(G138), .ZN(n528) );
  NAND2_X1 U578 ( .A1(n966), .A2(G102), .ZN(n527) );
  NAND2_X1 U579 ( .A1(n528), .A2(n527), .ZN(n529) );
  XNOR2_X1 U580 ( .A(n529), .B(KEYINPUT95), .ZN(n531) );
  NAND2_X1 U581 ( .A1(G114), .A2(n961), .ZN(n530) );
  NAND2_X1 U582 ( .A1(n531), .A2(n530), .ZN(n534) );
  NAND2_X1 U583 ( .A1(n962), .A2(G126), .ZN(n532) );
  XOR2_X1 U584 ( .A(n532), .B(KEYINPUT94), .Z(n533) );
  NOR2_X2 U585 ( .A1(n534), .A2(n533), .ZN(G164) );
  XOR2_X1 U586 ( .A(G2443), .B(G2451), .Z(n536) );
  XNOR2_X1 U587 ( .A(G2454), .B(G2435), .ZN(n535) );
  XNOR2_X1 U588 ( .A(n536), .B(n535), .ZN(n543) );
  XOR2_X1 U589 ( .A(G2427), .B(G2446), .Z(n538) );
  XNOR2_X1 U590 ( .A(G1341), .B(KEYINPUT111), .ZN(n537) );
  XNOR2_X1 U591 ( .A(n538), .B(n537), .ZN(n539) );
  XOR2_X1 U592 ( .A(n539), .B(G2438), .Z(n541) );
  INV_X1 U593 ( .A(G1348), .ZN(n843) );
  XOR2_X1 U594 ( .A(n843), .B(G2430), .Z(n540) );
  XNOR2_X1 U595 ( .A(n541), .B(n540), .ZN(n542) );
  XNOR2_X1 U596 ( .A(n543), .B(n542), .ZN(n544) );
  AND2_X1 U597 ( .A1(n544), .A2(G14), .ZN(G401) );
  XOR2_X1 U598 ( .A(KEYINPUT0), .B(G543), .Z(n627) );
  NAND2_X1 U599 ( .A1(n649), .A2(G52), .ZN(n548) );
  INV_X1 U600 ( .A(G651), .ZN(n550) );
  NOR2_X1 U601 ( .A1(G543), .A2(n550), .ZN(n545) );
  XOR2_X1 U602 ( .A(KEYINPUT1), .B(n545), .Z(n546) );
  XNOR2_X1 U603 ( .A(KEYINPUT70), .B(n546), .ZN(n653) );
  NAND2_X1 U604 ( .A1(G64), .A2(n653), .ZN(n547) );
  NAND2_X1 U605 ( .A1(n548), .A2(n547), .ZN(n556) );
  NOR2_X1 U606 ( .A1(G543), .A2(G651), .ZN(n648) );
  NAND2_X1 U607 ( .A1(n648), .A2(G90), .ZN(n549) );
  XNOR2_X1 U608 ( .A(n549), .B(KEYINPUT72), .ZN(n553) );
  OR2_X1 U609 ( .A1(n550), .A2(n627), .ZN(n551) );
  XNOR2_X1 U610 ( .A(KEYINPUT69), .B(n551), .ZN(n652) );
  NAND2_X1 U611 ( .A1(G77), .A2(n652), .ZN(n552) );
  NAND2_X1 U612 ( .A1(n553), .A2(n552), .ZN(n554) );
  XOR2_X1 U613 ( .A(KEYINPUT9), .B(n554), .Z(n555) );
  NOR2_X1 U614 ( .A1(n556), .A2(n555), .ZN(G171) );
  INV_X1 U615 ( .A(G171), .ZN(G301) );
  AND2_X1 U616 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U617 ( .A(G57), .ZN(G237) );
  INV_X1 U618 ( .A(G69), .ZN(G235) );
  INV_X1 U619 ( .A(G108), .ZN(G238) );
  INV_X1 U620 ( .A(G120), .ZN(G236) );
  INV_X1 U621 ( .A(G82), .ZN(G220) );
  NAND2_X1 U622 ( .A1(G89), .A2(n648), .ZN(n557) );
  XOR2_X1 U623 ( .A(KEYINPUT77), .B(n557), .Z(n558) );
  XNOR2_X1 U624 ( .A(n558), .B(KEYINPUT4), .ZN(n560) );
  NAND2_X1 U625 ( .A1(G76), .A2(n652), .ZN(n559) );
  NAND2_X1 U626 ( .A1(n560), .A2(n559), .ZN(n561) );
  XNOR2_X1 U627 ( .A(n561), .B(KEYINPUT5), .ZN(n566) );
  NAND2_X1 U628 ( .A1(n649), .A2(G51), .ZN(n563) );
  NAND2_X1 U629 ( .A1(G63), .A2(n653), .ZN(n562) );
  NAND2_X1 U630 ( .A1(n563), .A2(n562), .ZN(n564) );
  XOR2_X1 U631 ( .A(KEYINPUT6), .B(n564), .Z(n565) );
  NAND2_X1 U632 ( .A1(n566), .A2(n565), .ZN(n567) );
  XNOR2_X1 U633 ( .A(n567), .B(KEYINPUT7), .ZN(G168) );
  XOR2_X1 U634 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  XOR2_X1 U635 ( .A(KEYINPUT75), .B(KEYINPUT10), .Z(n569) );
  NAND2_X1 U636 ( .A1(G7), .A2(G661), .ZN(n568) );
  XNOR2_X1 U637 ( .A(n569), .B(n568), .ZN(G223) );
  XOR2_X1 U638 ( .A(G223), .B(KEYINPUT76), .Z(n826) );
  AND2_X1 U639 ( .A1(n826), .A2(G567), .ZN(n570) );
  XNOR2_X1 U640 ( .A(n570), .B(KEYINPUT11), .ZN(G234) );
  NAND2_X1 U641 ( .A1(n653), .A2(G56), .ZN(n571) );
  XOR2_X1 U642 ( .A(KEYINPUT14), .B(n571), .Z(n577) );
  NAND2_X1 U643 ( .A1(n648), .A2(G81), .ZN(n572) );
  XNOR2_X1 U644 ( .A(n572), .B(KEYINPUT12), .ZN(n574) );
  NAND2_X1 U645 ( .A1(G68), .A2(n652), .ZN(n573) );
  NAND2_X1 U646 ( .A1(n574), .A2(n573), .ZN(n575) );
  XOR2_X1 U647 ( .A(KEYINPUT13), .B(n575), .Z(n576) );
  NOR2_X1 U648 ( .A1(n577), .A2(n576), .ZN(n579) );
  NAND2_X1 U649 ( .A1(n649), .A2(G43), .ZN(n578) );
  NAND2_X1 U650 ( .A1(n579), .A2(n578), .ZN(n983) );
  INV_X1 U651 ( .A(G860), .ZN(n599) );
  OR2_X1 U652 ( .A1(n983), .A2(n599), .ZN(G153) );
  NAND2_X1 U653 ( .A1(G868), .A2(G301), .ZN(n588) );
  NAND2_X1 U654 ( .A1(n648), .A2(G92), .ZN(n581) );
  NAND2_X1 U655 ( .A1(G66), .A2(n653), .ZN(n580) );
  NAND2_X1 U656 ( .A1(n581), .A2(n580), .ZN(n585) );
  NAND2_X1 U657 ( .A1(G79), .A2(n652), .ZN(n583) );
  NAND2_X1 U658 ( .A1(G54), .A2(n649), .ZN(n582) );
  NAND2_X1 U659 ( .A1(n583), .A2(n582), .ZN(n584) );
  NOR2_X1 U660 ( .A1(n585), .A2(n584), .ZN(n586) );
  XOR2_X1 U661 ( .A(KEYINPUT15), .B(n586), .Z(n980) );
  OR2_X1 U662 ( .A1(n980), .A2(G868), .ZN(n587) );
  NAND2_X1 U663 ( .A1(n588), .A2(n587), .ZN(G284) );
  NAND2_X1 U664 ( .A1(G91), .A2(n648), .ZN(n590) );
  NAND2_X1 U665 ( .A1(G78), .A2(n652), .ZN(n589) );
  NAND2_X1 U666 ( .A1(n590), .A2(n589), .ZN(n593) );
  NAND2_X1 U667 ( .A1(G65), .A2(n653), .ZN(n591) );
  XNOR2_X1 U668 ( .A(KEYINPUT73), .B(n591), .ZN(n592) );
  NOR2_X1 U669 ( .A1(n593), .A2(n592), .ZN(n595) );
  NAND2_X1 U670 ( .A1(n649), .A2(G53), .ZN(n594) );
  NAND2_X1 U671 ( .A1(n595), .A2(n594), .ZN(G299) );
  INV_X1 U672 ( .A(G868), .ZN(n669) );
  NOR2_X1 U673 ( .A1(G286), .A2(n669), .ZN(n596) );
  XNOR2_X1 U674 ( .A(n596), .B(KEYINPUT78), .ZN(n598) );
  NOR2_X1 U675 ( .A1(G299), .A2(G868), .ZN(n597) );
  NOR2_X1 U676 ( .A1(n598), .A2(n597), .ZN(G297) );
  NAND2_X1 U677 ( .A1(n599), .A2(G559), .ZN(n600) );
  NAND2_X1 U678 ( .A1(n600), .A2(n980), .ZN(n601) );
  XNOR2_X1 U679 ( .A(n601), .B(KEYINPUT79), .ZN(n602) );
  XOR2_X1 U680 ( .A(KEYINPUT16), .B(n602), .Z(G148) );
  NOR2_X1 U681 ( .A1(G868), .A2(n983), .ZN(n605) );
  NAND2_X1 U682 ( .A1(n980), .A2(G868), .ZN(n603) );
  NOR2_X1 U683 ( .A1(G559), .A2(n603), .ZN(n604) );
  NOR2_X1 U684 ( .A1(n605), .A2(n604), .ZN(G282) );
  NAND2_X1 U685 ( .A1(G123), .A2(n962), .ZN(n606) );
  XNOR2_X1 U686 ( .A(n606), .B(KEYINPUT18), .ZN(n608) );
  NAND2_X1 U687 ( .A1(G135), .A2(n965), .ZN(n607) );
  NAND2_X1 U688 ( .A1(n608), .A2(n607), .ZN(n609) );
  XOR2_X1 U689 ( .A(KEYINPUT80), .B(n609), .Z(n611) );
  NAND2_X1 U690 ( .A1(n961), .A2(G111), .ZN(n610) );
  NAND2_X1 U691 ( .A1(n611), .A2(n610), .ZN(n614) );
  NAND2_X1 U692 ( .A1(G99), .A2(n966), .ZN(n612) );
  XNOR2_X1 U693 ( .A(KEYINPUT81), .B(n612), .ZN(n613) );
  NOR2_X1 U694 ( .A1(n614), .A2(n613), .ZN(n950) );
  XOR2_X1 U695 ( .A(n950), .B(G2096), .Z(n616) );
  XNOR2_X1 U696 ( .A(G2100), .B(KEYINPUT82), .ZN(n615) );
  NOR2_X1 U697 ( .A1(n616), .A2(n615), .ZN(n617) );
  XNOR2_X1 U698 ( .A(KEYINPUT83), .B(n617), .ZN(G156) );
  NAND2_X1 U699 ( .A1(G559), .A2(n980), .ZN(n618) );
  XNOR2_X1 U700 ( .A(n618), .B(n983), .ZN(n665) );
  NOR2_X1 U701 ( .A1(n665), .A2(G860), .ZN(n626) );
  NAND2_X1 U702 ( .A1(n649), .A2(G55), .ZN(n620) );
  NAND2_X1 U703 ( .A1(G67), .A2(n653), .ZN(n619) );
  NAND2_X1 U704 ( .A1(n620), .A2(n619), .ZN(n621) );
  XNOR2_X1 U705 ( .A(KEYINPUT84), .B(n621), .ZN(n625) );
  NAND2_X1 U706 ( .A1(G93), .A2(n648), .ZN(n623) );
  NAND2_X1 U707 ( .A1(G80), .A2(n652), .ZN(n622) );
  NAND2_X1 U708 ( .A1(n623), .A2(n622), .ZN(n624) );
  OR2_X1 U709 ( .A1(n625), .A2(n624), .ZN(n668) );
  XOR2_X1 U710 ( .A(n626), .B(n668), .Z(G145) );
  NAND2_X1 U711 ( .A1(G74), .A2(G651), .ZN(n629) );
  NAND2_X1 U712 ( .A1(G87), .A2(n627), .ZN(n628) );
  NAND2_X1 U713 ( .A1(n629), .A2(n628), .ZN(n630) );
  NOR2_X1 U714 ( .A1(n653), .A2(n630), .ZN(n632) );
  NAND2_X1 U715 ( .A1(n649), .A2(G49), .ZN(n631) );
  NAND2_X1 U716 ( .A1(n632), .A2(n631), .ZN(G288) );
  NAND2_X1 U717 ( .A1(n648), .A2(G86), .ZN(n634) );
  NAND2_X1 U718 ( .A1(G61), .A2(n653), .ZN(n633) );
  NAND2_X1 U719 ( .A1(n634), .A2(n633), .ZN(n637) );
  NAND2_X1 U720 ( .A1(n652), .A2(G73), .ZN(n635) );
  XOR2_X1 U721 ( .A(KEYINPUT2), .B(n635), .Z(n636) );
  NOR2_X1 U722 ( .A1(n637), .A2(n636), .ZN(n638) );
  XOR2_X1 U723 ( .A(KEYINPUT85), .B(n638), .Z(n640) );
  NAND2_X1 U724 ( .A1(n649), .A2(G48), .ZN(n639) );
  NAND2_X1 U725 ( .A1(n640), .A2(n639), .ZN(n641) );
  XNOR2_X1 U726 ( .A(KEYINPUT86), .B(n641), .ZN(G305) );
  NAND2_X1 U727 ( .A1(G88), .A2(n648), .ZN(n643) );
  NAND2_X1 U728 ( .A1(G75), .A2(n652), .ZN(n642) );
  NAND2_X1 U729 ( .A1(n643), .A2(n642), .ZN(n647) );
  NAND2_X1 U730 ( .A1(n649), .A2(G50), .ZN(n645) );
  NAND2_X1 U731 ( .A1(G62), .A2(n653), .ZN(n644) );
  NAND2_X1 U732 ( .A1(n645), .A2(n644), .ZN(n646) );
  NOR2_X1 U733 ( .A1(n647), .A2(n646), .ZN(G166) );
  NAND2_X1 U734 ( .A1(G85), .A2(n648), .ZN(n651) );
  NAND2_X1 U735 ( .A1(G47), .A2(n649), .ZN(n650) );
  NAND2_X1 U736 ( .A1(n651), .A2(n650), .ZN(n657) );
  NAND2_X1 U737 ( .A1(n652), .A2(G72), .ZN(n655) );
  NAND2_X1 U738 ( .A1(G60), .A2(n653), .ZN(n654) );
  NAND2_X1 U739 ( .A1(n655), .A2(n654), .ZN(n656) );
  NOR2_X1 U740 ( .A1(n657), .A2(n656), .ZN(n658) );
  XNOR2_X1 U741 ( .A(n658), .B(KEYINPUT71), .ZN(G290) );
  XNOR2_X1 U742 ( .A(KEYINPUT87), .B(KEYINPUT19), .ZN(n660) );
  XOR2_X1 U743 ( .A(G288), .B(n668), .Z(n659) );
  XNOR2_X1 U744 ( .A(n660), .B(n659), .ZN(n661) );
  XOR2_X1 U745 ( .A(n661), .B(G305), .Z(n663) );
  XOR2_X1 U746 ( .A(G299), .B(G166), .Z(n662) );
  XNOR2_X1 U747 ( .A(n663), .B(n662), .ZN(n664) );
  XNOR2_X1 U748 ( .A(n664), .B(G290), .ZN(n979) );
  XNOR2_X1 U749 ( .A(KEYINPUT88), .B(n665), .ZN(n666) );
  XNOR2_X1 U750 ( .A(n979), .B(n666), .ZN(n667) );
  NAND2_X1 U751 ( .A1(n667), .A2(G868), .ZN(n671) );
  NAND2_X1 U752 ( .A1(n669), .A2(n668), .ZN(n670) );
  NAND2_X1 U753 ( .A1(n671), .A2(n670), .ZN(G295) );
  NAND2_X1 U754 ( .A1(G2078), .A2(G2084), .ZN(n672) );
  XNOR2_X1 U755 ( .A(n672), .B(KEYINPUT89), .ZN(n673) );
  XNOR2_X1 U756 ( .A(n673), .B(KEYINPUT20), .ZN(n674) );
  NAND2_X1 U757 ( .A1(n674), .A2(G2090), .ZN(n675) );
  XNOR2_X1 U758 ( .A(KEYINPUT21), .B(n675), .ZN(n676) );
  NAND2_X1 U759 ( .A1(n676), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U760 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  XOR2_X1 U761 ( .A(KEYINPUT74), .B(G132), .Z(G219) );
  NOR2_X1 U762 ( .A1(G219), .A2(G220), .ZN(n678) );
  XNOR2_X1 U763 ( .A(KEYINPUT90), .B(KEYINPUT22), .ZN(n677) );
  XNOR2_X1 U764 ( .A(n678), .B(n677), .ZN(n679) );
  NAND2_X1 U765 ( .A1(n679), .A2(G96), .ZN(n680) );
  NOR2_X1 U766 ( .A1(G218), .A2(n680), .ZN(n681) );
  XNOR2_X1 U767 ( .A(KEYINPUT91), .B(n681), .ZN(n948) );
  NAND2_X1 U768 ( .A1(G2106), .A2(n948), .ZN(n682) );
  XOR2_X1 U769 ( .A(KEYINPUT92), .B(n682), .Z(n687) );
  NOR2_X1 U770 ( .A1(G236), .A2(G238), .ZN(n684) );
  NOR2_X1 U771 ( .A1(G235), .A2(G237), .ZN(n683) );
  NAND2_X1 U772 ( .A1(n684), .A2(n683), .ZN(n685) );
  XOR2_X1 U773 ( .A(KEYINPUT93), .B(n685), .Z(n949) );
  AND2_X1 U774 ( .A1(n949), .A2(G567), .ZN(n686) );
  NOR2_X1 U775 ( .A1(n687), .A2(n686), .ZN(G319) );
  INV_X1 U776 ( .A(G319), .ZN(n689) );
  NAND2_X1 U777 ( .A1(G483), .A2(G661), .ZN(n688) );
  NOR2_X1 U778 ( .A1(n689), .A2(n688), .ZN(n829) );
  NAND2_X1 U779 ( .A1(n829), .A2(G36), .ZN(G176) );
  XOR2_X1 U780 ( .A(G166), .B(KEYINPUT96), .Z(G303) );
  XOR2_X1 U781 ( .A(G1981), .B(G305), .Z(n850) );
  NOR2_X1 U782 ( .A1(G164), .A2(G1384), .ZN(n776) );
  INV_X1 U783 ( .A(n776), .ZN(n690) );
  NAND2_X1 U784 ( .A1(G160), .A2(G40), .ZN(n777) );
  NAND2_X1 U785 ( .A1(G8), .A2(n738), .ZN(n772) );
  NOR2_X1 U786 ( .A1(G288), .A2(G1976), .ZN(n691) );
  XOR2_X1 U787 ( .A(n691), .B(KEYINPUT109), .Z(n757) );
  INV_X1 U788 ( .A(n757), .ZN(n692) );
  NOR2_X1 U789 ( .A1(n772), .A2(n692), .ZN(n693) );
  NAND2_X1 U790 ( .A1(KEYINPUT33), .A2(n693), .ZN(n694) );
  NAND2_X1 U791 ( .A1(n850), .A2(n694), .ZN(n763) );
  NAND2_X1 U792 ( .A1(G1961), .A2(n738), .ZN(n697) );
  XOR2_X1 U793 ( .A(G2078), .B(KEYINPUT25), .Z(n695) );
  XNOR2_X1 U794 ( .A(KEYINPUT104), .B(n695), .ZN(n922) );
  NAND2_X1 U795 ( .A1(n708), .A2(n922), .ZN(n696) );
  NAND2_X1 U796 ( .A1(n697), .A2(n696), .ZN(n730) );
  OR2_X1 U797 ( .A1(G301), .A2(n730), .ZN(n724) );
  INV_X1 U798 ( .A(G299), .ZN(n718) );
  NAND2_X1 U799 ( .A1(n708), .A2(G2072), .ZN(n698) );
  XNOR2_X1 U800 ( .A(n698), .B(KEYINPUT27), .ZN(n700) );
  INV_X1 U801 ( .A(G1956), .ZN(n992) );
  NOR2_X1 U802 ( .A1(n992), .A2(n708), .ZN(n699) );
  NAND2_X1 U803 ( .A1(n718), .A2(n717), .ZN(n716) );
  INV_X1 U804 ( .A(G1996), .ZN(n989) );
  XOR2_X1 U805 ( .A(KEYINPUT64), .B(KEYINPUT26), .Z(n701) );
  XNOR2_X1 U806 ( .A(n702), .B(n701), .ZN(n704) );
  NAND2_X1 U807 ( .A1(n738), .A2(G1341), .ZN(n703) );
  NAND2_X1 U808 ( .A1(n704), .A2(n703), .ZN(n705) );
  OR2_X1 U809 ( .A1(n980), .A2(n706), .ZN(n714) );
  NAND2_X1 U810 ( .A1(n980), .A2(n706), .ZN(n712) );
  NOR2_X1 U811 ( .A1(n708), .A2(n843), .ZN(n707) );
  XNOR2_X1 U812 ( .A(n707), .B(KEYINPUT105), .ZN(n710) );
  NAND2_X1 U813 ( .A1(n708), .A2(G2067), .ZN(n709) );
  NAND2_X1 U814 ( .A1(n710), .A2(n709), .ZN(n711) );
  NAND2_X1 U815 ( .A1(n712), .A2(n711), .ZN(n713) );
  NAND2_X1 U816 ( .A1(n714), .A2(n713), .ZN(n715) );
  NAND2_X1 U817 ( .A1(n716), .A2(n715), .ZN(n720) );
  NOR2_X1 U818 ( .A1(n718), .A2(n717), .ZN(n719) );
  NAND2_X1 U819 ( .A1(n720), .A2(n513), .ZN(n722) );
  NAND2_X1 U820 ( .A1(n724), .A2(n723), .ZN(n736) );
  NOR2_X1 U821 ( .A1(G1966), .A2(n772), .ZN(n751) );
  NOR2_X1 U822 ( .A1(G2084), .A2(n738), .ZN(n747) );
  NOR2_X1 U823 ( .A1(n751), .A2(n747), .ZN(n725) );
  NAND2_X1 U824 ( .A1(G8), .A2(n725), .ZN(n727) );
  NOR2_X1 U825 ( .A1(n728), .A2(G168), .ZN(n729) );
  XNOR2_X1 U826 ( .A(n729), .B(KEYINPUT107), .ZN(n733) );
  NAND2_X1 U827 ( .A1(G301), .A2(n730), .ZN(n731) );
  XNOR2_X1 U828 ( .A(KEYINPUT108), .B(n731), .ZN(n732) );
  NAND2_X1 U829 ( .A1(n733), .A2(n732), .ZN(n734) );
  XNOR2_X1 U830 ( .A(n734), .B(KEYINPUT31), .ZN(n735) );
  NAND2_X1 U831 ( .A1(n736), .A2(n735), .ZN(n749) );
  AND2_X1 U832 ( .A1(G286), .A2(G8), .ZN(n737) );
  NAND2_X1 U833 ( .A1(n749), .A2(n737), .ZN(n745) );
  INV_X1 U834 ( .A(G8), .ZN(n743) );
  NOR2_X1 U835 ( .A1(G1971), .A2(n772), .ZN(n740) );
  NOR2_X1 U836 ( .A1(G2090), .A2(n738), .ZN(n739) );
  NOR2_X1 U837 ( .A1(n740), .A2(n739), .ZN(n741) );
  NAND2_X1 U838 ( .A1(n741), .A2(G303), .ZN(n742) );
  OR2_X1 U839 ( .A1(n743), .A2(n742), .ZN(n744) );
  XNOR2_X1 U840 ( .A(n746), .B(KEYINPUT32), .ZN(n755) );
  NAND2_X1 U841 ( .A1(G8), .A2(n747), .ZN(n748) );
  XOR2_X1 U842 ( .A(KEYINPUT103), .B(n748), .Z(n753) );
  INV_X1 U843 ( .A(n749), .ZN(n750) );
  NOR2_X1 U844 ( .A1(n751), .A2(n750), .ZN(n752) );
  NAND2_X1 U845 ( .A1(n753), .A2(n752), .ZN(n754) );
  NAND2_X1 U846 ( .A1(n755), .A2(n754), .ZN(n771) );
  NOR2_X1 U847 ( .A1(G303), .A2(G1971), .ZN(n756) );
  NOR2_X1 U848 ( .A1(n757), .A2(n756), .ZN(n840) );
  NAND2_X1 U849 ( .A1(n771), .A2(n840), .ZN(n759) );
  NAND2_X1 U850 ( .A1(G1976), .A2(G288), .ZN(n839) );
  INV_X1 U851 ( .A(n839), .ZN(n758) );
  XNOR2_X1 U852 ( .A(n761), .B(KEYINPUT110), .ZN(n762) );
  NOR2_X1 U853 ( .A1(n763), .A2(n762), .ZN(n768) );
  NOR2_X1 U854 ( .A1(G1981), .A2(G305), .ZN(n764) );
  XOR2_X1 U855 ( .A(n764), .B(KEYINPUT24), .Z(n765) );
  XNOR2_X1 U856 ( .A(KEYINPUT102), .B(n765), .ZN(n766) );
  NOR2_X1 U857 ( .A1(n766), .A2(n772), .ZN(n767) );
  NOR2_X1 U858 ( .A1(n768), .A2(n767), .ZN(n775) );
  NOR2_X1 U859 ( .A1(G2090), .A2(G303), .ZN(n769) );
  NAND2_X1 U860 ( .A1(G8), .A2(n769), .ZN(n770) );
  NAND2_X1 U861 ( .A1(n771), .A2(n770), .ZN(n773) );
  NAND2_X1 U862 ( .A1(n773), .A2(n772), .ZN(n774) );
  NAND2_X1 U863 ( .A1(n775), .A2(n774), .ZN(n811) );
  XNOR2_X1 U864 ( .A(G1986), .B(G290), .ZN(n854) );
  NOR2_X1 U865 ( .A1(n776), .A2(n777), .ZN(n821) );
  NAND2_X1 U866 ( .A1(n854), .A2(n821), .ZN(n809) );
  NAND2_X1 U867 ( .A1(n961), .A2(G107), .ZN(n779) );
  NAND2_X1 U868 ( .A1(G119), .A2(n962), .ZN(n778) );
  NAND2_X1 U869 ( .A1(n779), .A2(n778), .ZN(n780) );
  XOR2_X1 U870 ( .A(KEYINPUT98), .B(n780), .Z(n784) );
  NAND2_X1 U871 ( .A1(G131), .A2(n965), .ZN(n782) );
  NAND2_X1 U872 ( .A1(G95), .A2(n966), .ZN(n781) );
  AND2_X1 U873 ( .A1(n782), .A2(n781), .ZN(n783) );
  NAND2_X1 U874 ( .A1(n784), .A2(n783), .ZN(n975) );
  NAND2_X1 U875 ( .A1(G1991), .A2(n975), .ZN(n795) );
  NAND2_X1 U876 ( .A1(n966), .A2(G105), .ZN(n786) );
  XNOR2_X1 U877 ( .A(KEYINPUT38), .B(KEYINPUT100), .ZN(n785) );
  XNOR2_X1 U878 ( .A(n786), .B(n785), .ZN(n793) );
  NAND2_X1 U879 ( .A1(G117), .A2(n961), .ZN(n788) );
  NAND2_X1 U880 ( .A1(G141), .A2(n965), .ZN(n787) );
  NAND2_X1 U881 ( .A1(n788), .A2(n787), .ZN(n791) );
  NAND2_X1 U882 ( .A1(G129), .A2(n962), .ZN(n789) );
  XNOR2_X1 U883 ( .A(KEYINPUT99), .B(n789), .ZN(n790) );
  NOR2_X1 U884 ( .A1(n791), .A2(n790), .ZN(n792) );
  NAND2_X1 U885 ( .A1(n793), .A2(n792), .ZN(n972) );
  NAND2_X1 U886 ( .A1(G1996), .A2(n972), .ZN(n794) );
  NAND2_X1 U887 ( .A1(n795), .A2(n794), .ZN(n891) );
  NAND2_X1 U888 ( .A1(n821), .A2(n891), .ZN(n796) );
  XNOR2_X1 U889 ( .A(KEYINPUT101), .B(n796), .ZN(n814) );
  INV_X1 U890 ( .A(n814), .ZN(n807) );
  NAND2_X1 U891 ( .A1(n966), .A2(G104), .ZN(n798) );
  NAND2_X1 U892 ( .A1(n965), .A2(G140), .ZN(n797) );
  NAND2_X1 U893 ( .A1(n798), .A2(n797), .ZN(n799) );
  XNOR2_X1 U894 ( .A(KEYINPUT34), .B(n799), .ZN(n804) );
  NAND2_X1 U895 ( .A1(n961), .A2(G116), .ZN(n801) );
  NAND2_X1 U896 ( .A1(G128), .A2(n962), .ZN(n800) );
  NAND2_X1 U897 ( .A1(n801), .A2(n800), .ZN(n802) );
  XOR2_X1 U898 ( .A(n802), .B(KEYINPUT35), .Z(n803) );
  NOR2_X1 U899 ( .A1(n804), .A2(n803), .ZN(n805) );
  XOR2_X1 U900 ( .A(KEYINPUT36), .B(n805), .Z(n806) );
  XNOR2_X1 U901 ( .A(KEYINPUT97), .B(n806), .ZN(n951) );
  XNOR2_X1 U902 ( .A(G2067), .B(KEYINPUT37), .ZN(n819) );
  NOR2_X1 U903 ( .A1(n951), .A2(n819), .ZN(n894) );
  NAND2_X1 U904 ( .A1(n894), .A2(n821), .ZN(n817) );
  AND2_X1 U905 ( .A1(n807), .A2(n817), .ZN(n808) );
  AND2_X1 U906 ( .A1(n809), .A2(n808), .ZN(n810) );
  NAND2_X1 U907 ( .A1(n811), .A2(n810), .ZN(n824) );
  NOR2_X1 U908 ( .A1(G1996), .A2(n972), .ZN(n887) );
  NOR2_X1 U909 ( .A1(G1986), .A2(G290), .ZN(n812) );
  NOR2_X1 U910 ( .A1(G1991), .A2(n975), .ZN(n890) );
  NOR2_X1 U911 ( .A1(n812), .A2(n890), .ZN(n813) );
  NOR2_X1 U912 ( .A1(n814), .A2(n813), .ZN(n815) );
  NOR2_X1 U913 ( .A1(n887), .A2(n815), .ZN(n816) );
  XNOR2_X1 U914 ( .A(KEYINPUT39), .B(n816), .ZN(n818) );
  NAND2_X1 U915 ( .A1(n818), .A2(n817), .ZN(n820) );
  NAND2_X1 U916 ( .A1(n951), .A2(n819), .ZN(n912) );
  NAND2_X1 U917 ( .A1(n820), .A2(n912), .ZN(n822) );
  NAND2_X1 U918 ( .A1(n822), .A2(n821), .ZN(n823) );
  NAND2_X1 U919 ( .A1(n824), .A2(n823), .ZN(n825) );
  XNOR2_X1 U920 ( .A(n825), .B(KEYINPUT40), .ZN(G329) );
  NAND2_X1 U921 ( .A1(G2106), .A2(n826), .ZN(G217) );
  AND2_X1 U922 ( .A1(G15), .A2(G2), .ZN(n827) );
  NAND2_X1 U923 ( .A1(G661), .A2(n827), .ZN(G259) );
  NAND2_X1 U924 ( .A1(G3), .A2(G1), .ZN(n828) );
  NAND2_X1 U925 ( .A1(n829), .A2(n828), .ZN(G188) );
  XOR2_X1 U927 ( .A(KEYINPUT44), .B(KEYINPUT112), .Z(n831) );
  NAND2_X1 U928 ( .A1(G124), .A2(n962), .ZN(n830) );
  XNOR2_X1 U929 ( .A(n831), .B(n830), .ZN(n838) );
  NAND2_X1 U930 ( .A1(G112), .A2(n961), .ZN(n833) );
  NAND2_X1 U931 ( .A1(G100), .A2(n966), .ZN(n832) );
  NAND2_X1 U932 ( .A1(n833), .A2(n832), .ZN(n834) );
  XNOR2_X1 U933 ( .A(n834), .B(KEYINPUT113), .ZN(n836) );
  NAND2_X1 U934 ( .A1(G136), .A2(n965), .ZN(n835) );
  NAND2_X1 U935 ( .A1(n836), .A2(n835), .ZN(n837) );
  NOR2_X1 U936 ( .A1(n838), .A2(n837), .ZN(G162) );
  NAND2_X1 U937 ( .A1(n840), .A2(n839), .ZN(n842) );
  XOR2_X1 U938 ( .A(n992), .B(G299), .Z(n841) );
  NOR2_X1 U939 ( .A1(n842), .A2(n841), .ZN(n849) );
  XOR2_X1 U940 ( .A(n980), .B(n843), .Z(n845) );
  NAND2_X1 U941 ( .A1(G1971), .A2(G303), .ZN(n844) );
  NAND2_X1 U942 ( .A1(n845), .A2(n844), .ZN(n847) );
  XNOR2_X1 U943 ( .A(G1341), .B(n983), .ZN(n846) );
  NOR2_X1 U944 ( .A1(n847), .A2(n846), .ZN(n848) );
  NAND2_X1 U945 ( .A1(n849), .A2(n848), .ZN(n858) );
  XNOR2_X1 U946 ( .A(G1966), .B(G168), .ZN(n851) );
  NAND2_X1 U947 ( .A1(n851), .A2(n850), .ZN(n852) );
  XNOR2_X1 U948 ( .A(n852), .B(KEYINPUT57), .ZN(n856) );
  XOR2_X1 U949 ( .A(G1961), .B(G171), .Z(n853) );
  NOR2_X1 U950 ( .A1(n854), .A2(n853), .ZN(n855) );
  NAND2_X1 U951 ( .A1(n856), .A2(n855), .ZN(n857) );
  NOR2_X1 U952 ( .A1(n858), .A2(n857), .ZN(n859) );
  XOR2_X1 U953 ( .A(KEYINPUT124), .B(n859), .Z(n861) );
  XNOR2_X1 U954 ( .A(G16), .B(KEYINPUT56), .ZN(n860) );
  NAND2_X1 U955 ( .A1(n861), .A2(n860), .ZN(n946) );
  XNOR2_X1 U956 ( .A(G1966), .B(G21), .ZN(n863) );
  XNOR2_X1 U957 ( .A(G1961), .B(G5), .ZN(n862) );
  NOR2_X1 U958 ( .A1(n863), .A2(n862), .ZN(n874) );
  XOR2_X1 U959 ( .A(G1341), .B(G19), .Z(n865) );
  XOR2_X1 U960 ( .A(G1956), .B(G20), .Z(n864) );
  NAND2_X1 U961 ( .A1(n865), .A2(n864), .ZN(n871) );
  XOR2_X1 U962 ( .A(G1981), .B(G6), .Z(n869) );
  XNOR2_X1 U963 ( .A(G4), .B(KEYINPUT125), .ZN(n866) );
  XOR2_X1 U964 ( .A(n866), .B(G1348), .Z(n867) );
  XNOR2_X1 U965 ( .A(n867), .B(KEYINPUT59), .ZN(n868) );
  NAND2_X1 U966 ( .A1(n869), .A2(n868), .ZN(n870) );
  NOR2_X1 U967 ( .A1(n871), .A2(n870), .ZN(n872) );
  XNOR2_X1 U968 ( .A(n872), .B(KEYINPUT60), .ZN(n873) );
  NAND2_X1 U969 ( .A1(n874), .A2(n873), .ZN(n881) );
  XNOR2_X1 U970 ( .A(G1971), .B(G22), .ZN(n876) );
  XNOR2_X1 U971 ( .A(G23), .B(G1976), .ZN(n875) );
  NOR2_X1 U972 ( .A1(n876), .A2(n875), .ZN(n878) );
  XOR2_X1 U973 ( .A(G1986), .B(G24), .Z(n877) );
  NAND2_X1 U974 ( .A1(n878), .A2(n877), .ZN(n879) );
  XNOR2_X1 U975 ( .A(KEYINPUT58), .B(n879), .ZN(n880) );
  NOR2_X1 U976 ( .A1(n881), .A2(n880), .ZN(n882) );
  XOR2_X1 U977 ( .A(KEYINPUT61), .B(n882), .Z(n883) );
  NOR2_X1 U978 ( .A1(G16), .A2(n883), .ZN(n884) );
  XOR2_X1 U979 ( .A(KEYINPUT126), .B(n884), .Z(n885) );
  NAND2_X1 U980 ( .A1(G11), .A2(n885), .ZN(n944) );
  INV_X1 U981 ( .A(G29), .ZN(n940) );
  XOR2_X1 U982 ( .A(G2090), .B(G162), .Z(n886) );
  NOR2_X1 U983 ( .A1(n887), .A2(n886), .ZN(n888) );
  XOR2_X1 U984 ( .A(KEYINPUT51), .B(n888), .Z(n898) );
  XOR2_X1 U985 ( .A(G2084), .B(G160), .Z(n889) );
  NOR2_X1 U986 ( .A1(n890), .A2(n889), .ZN(n893) );
  NOR2_X1 U987 ( .A1(n950), .A2(n891), .ZN(n892) );
  NAND2_X1 U988 ( .A1(n893), .A2(n892), .ZN(n895) );
  NOR2_X1 U989 ( .A1(n895), .A2(n894), .ZN(n896) );
  XOR2_X1 U990 ( .A(KEYINPUT117), .B(n896), .Z(n897) );
  NAND2_X1 U991 ( .A1(n898), .A2(n897), .ZN(n910) );
  NAND2_X1 U992 ( .A1(G139), .A2(n965), .ZN(n900) );
  NAND2_X1 U993 ( .A1(G103), .A2(n966), .ZN(n899) );
  NAND2_X1 U994 ( .A1(n900), .A2(n899), .ZN(n905) );
  NAND2_X1 U995 ( .A1(n961), .A2(G115), .ZN(n902) );
  NAND2_X1 U996 ( .A1(G127), .A2(n962), .ZN(n901) );
  NAND2_X1 U997 ( .A1(n902), .A2(n901), .ZN(n903) );
  XOR2_X1 U998 ( .A(KEYINPUT47), .B(n903), .Z(n904) );
  NOR2_X1 U999 ( .A1(n905), .A2(n904), .ZN(n958) );
  XOR2_X1 U1000 ( .A(G2072), .B(n958), .Z(n907) );
  XOR2_X1 U1001 ( .A(G164), .B(G2078), .Z(n906) );
  NOR2_X1 U1002 ( .A1(n907), .A2(n906), .ZN(n908) );
  XOR2_X1 U1003 ( .A(KEYINPUT50), .B(n908), .Z(n909) );
  NOR2_X1 U1004 ( .A1(n910), .A2(n909), .ZN(n911) );
  NAND2_X1 U1005 ( .A1(n912), .A2(n911), .ZN(n913) );
  XNOR2_X1 U1006 ( .A(n913), .B(KEYINPUT52), .ZN(n914) );
  XNOR2_X1 U1007 ( .A(n914), .B(KEYINPUT118), .ZN(n915) );
  NOR2_X1 U1008 ( .A1(KEYINPUT55), .A2(n915), .ZN(n916) );
  NOR2_X1 U1009 ( .A1(n940), .A2(n916), .ZN(n917) );
  XNOR2_X1 U1010 ( .A(n917), .B(KEYINPUT119), .ZN(n942) );
  XOR2_X1 U1011 ( .A(G2084), .B(G34), .Z(n918) );
  XNOR2_X1 U1012 ( .A(KEYINPUT54), .B(n918), .ZN(n936) );
  XNOR2_X1 U1013 ( .A(G2090), .B(G35), .ZN(n934) );
  XOR2_X1 U1014 ( .A(G1991), .B(G25), .Z(n919) );
  XNOR2_X1 U1015 ( .A(KEYINPUT120), .B(n919), .ZN(n920) );
  NAND2_X1 U1016 ( .A1(G28), .A2(n920), .ZN(n921) );
  XOR2_X1 U1017 ( .A(KEYINPUT121), .B(n921), .Z(n931) );
  XOR2_X1 U1018 ( .A(G32), .B(G1996), .Z(n926) );
  XNOR2_X1 U1019 ( .A(n922), .B(G27), .ZN(n924) );
  XNOR2_X1 U1020 ( .A(G26), .B(G2067), .ZN(n923) );
  NOR2_X1 U1021 ( .A1(n924), .A2(n923), .ZN(n925) );
  NAND2_X1 U1022 ( .A1(n926), .A2(n925), .ZN(n928) );
  XNOR2_X1 U1023 ( .A(G33), .B(G2072), .ZN(n927) );
  NOR2_X1 U1024 ( .A1(n928), .A2(n927), .ZN(n929) );
  XOR2_X1 U1025 ( .A(KEYINPUT122), .B(n929), .Z(n930) );
  NOR2_X1 U1026 ( .A1(n931), .A2(n930), .ZN(n932) );
  XNOR2_X1 U1027 ( .A(KEYINPUT53), .B(n932), .ZN(n933) );
  NOR2_X1 U1028 ( .A1(n934), .A2(n933), .ZN(n935) );
  NAND2_X1 U1029 ( .A1(n936), .A2(n935), .ZN(n938) );
  XNOR2_X1 U1030 ( .A(KEYINPUT123), .B(KEYINPUT55), .ZN(n937) );
  XNOR2_X1 U1031 ( .A(n938), .B(n937), .ZN(n939) );
  NAND2_X1 U1032 ( .A1(n940), .A2(n939), .ZN(n941) );
  NAND2_X1 U1033 ( .A1(n942), .A2(n941), .ZN(n943) );
  NOR2_X1 U1034 ( .A1(n944), .A2(n943), .ZN(n945) );
  NAND2_X1 U1035 ( .A1(n946), .A2(n945), .ZN(n947) );
  XOR2_X1 U1036 ( .A(KEYINPUT62), .B(n947), .Z(G311) );
  XNOR2_X1 U1037 ( .A(KEYINPUT127), .B(G311), .ZN(G150) );
  INV_X1 U1038 ( .A(G96), .ZN(G221) );
  NOR2_X1 U1039 ( .A1(n949), .A2(n948), .ZN(G325) );
  INV_X1 U1040 ( .A(G325), .ZN(G261) );
  XNOR2_X1 U1041 ( .A(n950), .B(G162), .ZN(n953) );
  XNOR2_X1 U1042 ( .A(n951), .B(G164), .ZN(n952) );
  XNOR2_X1 U1043 ( .A(n953), .B(n952), .ZN(n957) );
  XOR2_X1 U1044 ( .A(KEYINPUT114), .B(KEYINPUT115), .Z(n955) );
  XNOR2_X1 U1045 ( .A(KEYINPUT46), .B(KEYINPUT48), .ZN(n954) );
  XNOR2_X1 U1046 ( .A(n955), .B(n954), .ZN(n956) );
  XOR2_X1 U1047 ( .A(n957), .B(n956), .Z(n960) );
  XNOR2_X1 U1048 ( .A(G160), .B(n958), .ZN(n959) );
  XNOR2_X1 U1049 ( .A(n960), .B(n959), .ZN(n977) );
  NAND2_X1 U1050 ( .A1(n961), .A2(G118), .ZN(n964) );
  NAND2_X1 U1051 ( .A1(G130), .A2(n962), .ZN(n963) );
  NAND2_X1 U1052 ( .A1(n964), .A2(n963), .ZN(n971) );
  NAND2_X1 U1053 ( .A1(G142), .A2(n965), .ZN(n968) );
  NAND2_X1 U1054 ( .A1(G106), .A2(n966), .ZN(n967) );
  NAND2_X1 U1055 ( .A1(n968), .A2(n967), .ZN(n969) );
  XOR2_X1 U1056 ( .A(n969), .B(KEYINPUT45), .Z(n970) );
  NOR2_X1 U1057 ( .A1(n971), .A2(n970), .ZN(n973) );
  XNOR2_X1 U1058 ( .A(n973), .B(n972), .ZN(n974) );
  XOR2_X1 U1059 ( .A(n975), .B(n974), .Z(n976) );
  XNOR2_X1 U1060 ( .A(n977), .B(n976), .ZN(n978) );
  NOR2_X1 U1061 ( .A1(G37), .A2(n978), .ZN(G395) );
  XOR2_X1 U1062 ( .A(n979), .B(G286), .Z(n982) );
  XOR2_X1 U1063 ( .A(G301), .B(n980), .Z(n981) );
  XNOR2_X1 U1064 ( .A(n982), .B(n981), .ZN(n984) );
  XNOR2_X1 U1065 ( .A(n984), .B(n983), .ZN(n985) );
  NOR2_X1 U1066 ( .A1(G37), .A2(n985), .ZN(G397) );
  XOR2_X1 U1067 ( .A(G1971), .B(G1961), .Z(n987) );
  XNOR2_X1 U1068 ( .A(G1986), .B(G1966), .ZN(n986) );
  XNOR2_X1 U1069 ( .A(n987), .B(n986), .ZN(n988) );
  XOR2_X1 U1070 ( .A(n988), .B(KEYINPUT41), .Z(n991) );
  XOR2_X1 U1071 ( .A(n989), .B(G1976), .Z(n990) );
  XNOR2_X1 U1072 ( .A(n991), .B(n990), .ZN(n996) );
  XOR2_X1 U1073 ( .A(G2474), .B(G1981), .Z(n994) );
  XOR2_X1 U1074 ( .A(G1991), .B(n992), .Z(n993) );
  XNOR2_X1 U1075 ( .A(n994), .B(n993), .ZN(n995) );
  XNOR2_X1 U1076 ( .A(n996), .B(n995), .ZN(G229) );
  XOR2_X1 U1077 ( .A(G2100), .B(G2096), .Z(n998) );
  XNOR2_X1 U1078 ( .A(G2072), .B(G2090), .ZN(n997) );
  XNOR2_X1 U1079 ( .A(n998), .B(n997), .ZN(n1002) );
  XOR2_X1 U1080 ( .A(G2678), .B(KEYINPUT42), .Z(n1000) );
  XNOR2_X1 U1081 ( .A(G2067), .B(KEYINPUT43), .ZN(n999) );
  XNOR2_X1 U1082 ( .A(n1000), .B(n999), .ZN(n1001) );
  XOR2_X1 U1083 ( .A(n1002), .B(n1001), .Z(n1004) );
  XNOR2_X1 U1084 ( .A(G2078), .B(G2084), .ZN(n1003) );
  XNOR2_X1 U1085 ( .A(n1004), .B(n1003), .ZN(G227) );
  NOR2_X1 U1086 ( .A1(G395), .A2(G397), .ZN(n1005) );
  XNOR2_X1 U1087 ( .A(n1005), .B(KEYINPUT116), .ZN(n1006) );
  NAND2_X1 U1088 ( .A1(G319), .A2(n1006), .ZN(n1007) );
  NOR2_X1 U1089 ( .A1(G401), .A2(n1007), .ZN(n1010) );
  NOR2_X1 U1090 ( .A1(G229), .A2(G227), .ZN(n1008) );
  XOR2_X1 U1091 ( .A(KEYINPUT49), .B(n1008), .Z(n1009) );
  NAND2_X1 U1092 ( .A1(n1010), .A2(n1009), .ZN(G225) );
  INV_X1 U1093 ( .A(G225), .ZN(G308) );
endmodule

