//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 1 0 0 1 0 0 0 1 1 1 0 1 1 0 1 0 1 0 0 1 1 0 0 0 0 0 0 0 0 1 0 0 0 0 0 1 0 0 0 1 0 0 1 1 1 1 1 1 0 1 0 1 1 1 1 0 0 0 0 0 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:26:50 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n717,
    new_n718, new_n719, new_n720, new_n721, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n729, new_n731, new_n732, new_n733, new_n735,
    new_n736, new_n737, new_n738, new_n739, new_n740, new_n741, new_n742,
    new_n743, new_n744, new_n745, new_n746, new_n747, new_n748, new_n749,
    new_n750, new_n751, new_n752, new_n754, new_n755, new_n756, new_n757,
    new_n758, new_n759, new_n760, new_n761, new_n762, new_n763, new_n764,
    new_n765, new_n766, new_n767, new_n768, new_n769, new_n770, new_n771,
    new_n772, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n791, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n816, new_n817,
    new_n818, new_n819, new_n820, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n947, new_n948, new_n949, new_n950, new_n951, new_n952,
    new_n953, new_n954, new_n955, new_n956, new_n957, new_n958, new_n959,
    new_n960, new_n961, new_n962, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n976, new_n977, new_n978, new_n979, new_n981, new_n982, new_n983,
    new_n984, new_n985, new_n986, new_n987, new_n988, new_n989, new_n990,
    new_n991, new_n993, new_n994, new_n995, new_n996, new_n997, new_n998,
    new_n999, new_n1000, new_n1001, new_n1002, new_n1003, new_n1004,
    new_n1005, new_n1006, new_n1007, new_n1009, new_n1010, new_n1011,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1022, new_n1023, new_n1024,
    new_n1025, new_n1026, new_n1027, new_n1028, new_n1029, new_n1030,
    new_n1031, new_n1032, new_n1033, new_n1034, new_n1035, new_n1036,
    new_n1037, new_n1038, new_n1040, new_n1041, new_n1042, new_n1043,
    new_n1044, new_n1045, new_n1046, new_n1047, new_n1048, new_n1049,
    new_n1050, new_n1051, new_n1052, new_n1053;
  INV_X1    g000(.A(G221), .ZN(new_n187));
  XNOR2_X1  g001(.A(KEYINPUT9), .B(G234), .ZN(new_n188));
  INV_X1    g002(.A(new_n188), .ZN(new_n189));
  INV_X1    g003(.A(G902), .ZN(new_n190));
  AOI21_X1  g004(.A(new_n187), .B1(new_n189), .B2(new_n190), .ZN(new_n191));
  INV_X1    g005(.A(KEYINPUT11), .ZN(new_n192));
  INV_X1    g006(.A(G134), .ZN(new_n193));
  OAI21_X1  g007(.A(new_n192), .B1(new_n193), .B2(G137), .ZN(new_n194));
  AOI21_X1  g008(.A(G131), .B1(new_n193), .B2(G137), .ZN(new_n195));
  INV_X1    g009(.A(G137), .ZN(new_n196));
  NAND3_X1  g010(.A1(new_n196), .A2(KEYINPUT11), .A3(G134), .ZN(new_n197));
  NAND3_X1  g011(.A1(new_n194), .A2(new_n195), .A3(new_n197), .ZN(new_n198));
  INV_X1    g012(.A(KEYINPUT65), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n198), .A2(new_n199), .ZN(new_n200));
  NAND4_X1  g014(.A1(new_n194), .A2(new_n195), .A3(KEYINPUT65), .A4(new_n197), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n200), .A2(new_n201), .ZN(new_n202));
  OAI211_X1 g016(.A(new_n194), .B(new_n197), .C1(G134), .C2(new_n196), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n203), .A2(G131), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n202), .A2(new_n204), .ZN(new_n205));
  XNOR2_X1  g019(.A(G104), .B(G107), .ZN(new_n206));
  INV_X1    g020(.A(G101), .ZN(new_n207));
  OAI21_X1  g021(.A(KEYINPUT81), .B1(new_n206), .B2(new_n207), .ZN(new_n208));
  INV_X1    g022(.A(G104), .ZN(new_n209));
  OAI21_X1  g023(.A(KEYINPUT3), .B1(new_n209), .B2(G107), .ZN(new_n210));
  INV_X1    g024(.A(KEYINPUT3), .ZN(new_n211));
  INV_X1    g025(.A(G107), .ZN(new_n212));
  NAND3_X1  g026(.A1(new_n211), .A2(new_n212), .A3(G104), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n209), .A2(G107), .ZN(new_n214));
  NAND4_X1  g028(.A1(new_n210), .A2(new_n213), .A3(new_n207), .A4(new_n214), .ZN(new_n215));
  INV_X1    g029(.A(KEYINPUT81), .ZN(new_n216));
  NOR2_X1   g030(.A1(new_n209), .A2(G107), .ZN(new_n217));
  NOR2_X1   g031(.A1(new_n212), .A2(G104), .ZN(new_n218));
  OAI211_X1 g032(.A(new_n216), .B(G101), .C1(new_n217), .C2(new_n218), .ZN(new_n219));
  AND3_X1   g033(.A1(new_n208), .A2(new_n215), .A3(new_n219), .ZN(new_n220));
  INV_X1    g034(.A(G146), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n221), .A2(KEYINPUT64), .ZN(new_n222));
  INV_X1    g036(.A(KEYINPUT64), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n223), .A2(G146), .ZN(new_n224));
  NAND3_X1  g038(.A1(new_n222), .A2(new_n224), .A3(G143), .ZN(new_n225));
  NOR2_X1   g039(.A1(new_n221), .A2(G143), .ZN(new_n226));
  INV_X1    g040(.A(new_n226), .ZN(new_n227));
  INV_X1    g041(.A(G128), .ZN(new_n228));
  NOR2_X1   g042(.A1(new_n228), .A2(KEYINPUT1), .ZN(new_n229));
  NAND3_X1  g043(.A1(new_n225), .A2(new_n227), .A3(new_n229), .ZN(new_n230));
  XNOR2_X1  g044(.A(KEYINPUT64), .B(G146), .ZN(new_n231));
  AOI21_X1  g045(.A(new_n226), .B1(new_n231), .B2(G143), .ZN(new_n232));
  INV_X1    g046(.A(G143), .ZN(new_n233));
  NOR2_X1   g047(.A1(new_n233), .A2(G146), .ZN(new_n234));
  INV_X1    g048(.A(new_n234), .ZN(new_n235));
  AOI21_X1  g049(.A(new_n228), .B1(new_n235), .B2(KEYINPUT1), .ZN(new_n236));
  OAI21_X1  g050(.A(new_n230), .B1(new_n232), .B2(new_n236), .ZN(new_n237));
  AND2_X1   g051(.A1(new_n220), .A2(new_n237), .ZN(new_n238));
  AOI21_X1  g052(.A(new_n228), .B1(new_n225), .B2(KEYINPUT1), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n222), .A2(new_n224), .ZN(new_n240));
  AOI21_X1  g054(.A(new_n234), .B1(new_n240), .B2(new_n233), .ZN(new_n241));
  OAI21_X1  g055(.A(new_n230), .B1(new_n239), .B2(new_n241), .ZN(new_n242));
  NOR2_X1   g056(.A1(new_n242), .A2(new_n220), .ZN(new_n243));
  OAI21_X1  g057(.A(new_n205), .B1(new_n238), .B2(new_n243), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n244), .A2(KEYINPUT12), .ZN(new_n245));
  INV_X1    g059(.A(KEYINPUT12), .ZN(new_n246));
  OAI211_X1 g060(.A(new_n246), .B(new_n205), .C1(new_n238), .C2(new_n243), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n245), .A2(new_n247), .ZN(new_n248));
  INV_X1    g062(.A(KEYINPUT79), .ZN(new_n249));
  NAND3_X1  g063(.A1(new_n210), .A2(new_n213), .A3(new_n214), .ZN(new_n250));
  NAND3_X1  g064(.A1(new_n250), .A2(KEYINPUT78), .A3(G101), .ZN(new_n251));
  NAND3_X1  g065(.A1(new_n251), .A2(KEYINPUT4), .A3(new_n215), .ZN(new_n252));
  AOI21_X1  g066(.A(KEYINPUT78), .B1(new_n250), .B2(G101), .ZN(new_n253));
  OAI21_X1  g067(.A(new_n249), .B1(new_n252), .B2(new_n253), .ZN(new_n254));
  INV_X1    g068(.A(new_n253), .ZN(new_n255));
  AND2_X1   g069(.A1(new_n215), .A2(KEYINPUT4), .ZN(new_n256));
  NAND4_X1  g070(.A1(new_n255), .A2(new_n256), .A3(KEYINPUT79), .A4(new_n251), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n254), .A2(new_n257), .ZN(new_n258));
  AND2_X1   g072(.A1(KEYINPUT0), .A2(G128), .ZN(new_n259));
  NAND3_X1  g073(.A1(new_n225), .A2(new_n259), .A3(new_n227), .ZN(new_n260));
  NOR2_X1   g074(.A1(KEYINPUT0), .A2(G128), .ZN(new_n261));
  NOR2_X1   g075(.A1(new_n259), .A2(new_n261), .ZN(new_n262));
  INV_X1    g076(.A(new_n262), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n250), .A2(G101), .ZN(new_n264));
  INV_X1    g078(.A(KEYINPUT80), .ZN(new_n265));
  OR2_X1    g079(.A1(new_n265), .A2(KEYINPUT4), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n265), .A2(KEYINPUT4), .ZN(new_n267));
  AND2_X1   g081(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  OAI221_X1 g082(.A(new_n260), .B1(new_n241), .B2(new_n263), .C1(new_n264), .C2(new_n268), .ZN(new_n269));
  INV_X1    g083(.A(new_n269), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n258), .A2(new_n270), .ZN(new_n271));
  AOI22_X1  g085(.A1(new_n200), .A2(new_n201), .B1(G131), .B2(new_n203), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n242), .A2(new_n220), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n273), .A2(KEYINPUT10), .ZN(new_n274));
  INV_X1    g088(.A(KEYINPUT10), .ZN(new_n275));
  NAND3_X1  g089(.A1(new_n220), .A2(new_n237), .A3(new_n275), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n274), .A2(new_n276), .ZN(new_n277));
  NAND3_X1  g091(.A1(new_n271), .A2(new_n272), .A3(new_n277), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n278), .A2(KEYINPUT82), .ZN(new_n279));
  AOI22_X1  g093(.A1(new_n258), .A2(new_n270), .B1(new_n274), .B2(new_n276), .ZN(new_n280));
  INV_X1    g094(.A(KEYINPUT82), .ZN(new_n281));
  NAND3_X1  g095(.A1(new_n280), .A2(new_n281), .A3(new_n272), .ZN(new_n282));
  AOI21_X1  g096(.A(new_n248), .B1(new_n279), .B2(new_n282), .ZN(new_n283));
  INV_X1    g097(.A(KEYINPUT83), .ZN(new_n284));
  XOR2_X1   g098(.A(G110), .B(G140), .Z(new_n285));
  XNOR2_X1  g099(.A(new_n285), .B(KEYINPUT76), .ZN(new_n286));
  XOR2_X1   g100(.A(new_n286), .B(KEYINPUT77), .Z(new_n287));
  INV_X1    g101(.A(G953), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n288), .A2(G227), .ZN(new_n289));
  XOR2_X1   g103(.A(new_n287), .B(new_n289), .Z(new_n290));
  NAND3_X1  g104(.A1(new_n283), .A2(new_n284), .A3(new_n290), .ZN(new_n291));
  INV_X1    g105(.A(new_n280), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n292), .A2(new_n205), .ZN(new_n293));
  AOI21_X1  g107(.A(new_n281), .B1(new_n280), .B2(new_n272), .ZN(new_n294));
  AOI21_X1  g108(.A(new_n275), .B1(new_n242), .B2(new_n220), .ZN(new_n295));
  AOI21_X1  g109(.A(new_n295), .B1(new_n275), .B2(new_n238), .ZN(new_n296));
  AOI21_X1  g110(.A(new_n269), .B1(new_n254), .B2(new_n257), .ZN(new_n297));
  NOR4_X1   g111(.A1(new_n296), .A2(new_n297), .A3(KEYINPUT82), .A4(new_n205), .ZN(new_n298));
  OAI21_X1  g112(.A(new_n293), .B1(new_n294), .B2(new_n298), .ZN(new_n299));
  INV_X1    g113(.A(new_n290), .ZN(new_n300));
  AOI21_X1  g114(.A(KEYINPUT83), .B1(new_n299), .B2(new_n300), .ZN(new_n301));
  INV_X1    g115(.A(new_n248), .ZN(new_n302));
  OAI211_X1 g116(.A(new_n290), .B(new_n302), .C1(new_n294), .C2(new_n298), .ZN(new_n303));
  INV_X1    g117(.A(new_n303), .ZN(new_n304));
  OAI21_X1  g118(.A(new_n291), .B1(new_n301), .B2(new_n304), .ZN(new_n305));
  INV_X1    g119(.A(G469), .ZN(new_n306));
  NAND3_X1  g120(.A1(new_n305), .A2(new_n306), .A3(new_n190), .ZN(new_n307));
  OAI211_X1 g121(.A(new_n290), .B(new_n293), .C1(new_n294), .C2(new_n298), .ZN(new_n308));
  OAI211_X1 g122(.A(new_n308), .B(G469), .C1(new_n290), .C2(new_n283), .ZN(new_n309));
  INV_X1    g123(.A(new_n309), .ZN(new_n310));
  NOR2_X1   g124(.A1(new_n306), .A2(new_n190), .ZN(new_n311));
  NOR2_X1   g125(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  AOI21_X1  g126(.A(new_n191), .B1(new_n307), .B2(new_n312), .ZN(new_n313));
  INV_X1    g127(.A(KEYINPUT6), .ZN(new_n314));
  INV_X1    g128(.A(G116), .ZN(new_n315));
  NOR2_X1   g129(.A1(new_n315), .A2(G119), .ZN(new_n316));
  INV_X1    g130(.A(new_n316), .ZN(new_n317));
  OAI21_X1  g131(.A(G113), .B1(new_n317), .B2(KEYINPUT5), .ZN(new_n318));
  XNOR2_X1  g132(.A(KEYINPUT67), .B(G116), .ZN(new_n319));
  AOI21_X1  g133(.A(new_n316), .B1(new_n319), .B2(G119), .ZN(new_n320));
  AOI21_X1  g134(.A(new_n318), .B1(new_n320), .B2(KEYINPUT5), .ZN(new_n321));
  NAND3_X1  g135(.A1(new_n208), .A2(new_n215), .A3(new_n219), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n315), .A2(KEYINPUT67), .ZN(new_n323));
  INV_X1    g137(.A(KEYINPUT67), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n324), .A2(G116), .ZN(new_n325));
  NAND3_X1  g139(.A1(new_n323), .A2(new_n325), .A3(G119), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n326), .A2(new_n317), .ZN(new_n327));
  XOR2_X1   g141(.A(KEYINPUT2), .B(G113), .Z(new_n328));
  INV_X1    g142(.A(new_n328), .ZN(new_n329));
  NOR2_X1   g143(.A1(new_n327), .A2(new_n329), .ZN(new_n330));
  NOR3_X1   g144(.A1(new_n321), .A2(new_n322), .A3(new_n330), .ZN(new_n331));
  NOR2_X1   g145(.A1(new_n264), .A2(new_n268), .ZN(new_n332));
  INV_X1    g146(.A(KEYINPUT68), .ZN(new_n333));
  AOI21_X1  g147(.A(new_n328), .B1(new_n317), .B2(new_n326), .ZN(new_n334));
  OAI21_X1  g148(.A(new_n333), .B1(new_n330), .B2(new_n334), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n320), .A2(new_n328), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n327), .A2(new_n329), .ZN(new_n337));
  NAND3_X1  g151(.A1(new_n336), .A2(new_n337), .A3(KEYINPUT68), .ZN(new_n338));
  AOI21_X1  g152(.A(new_n332), .B1(new_n335), .B2(new_n338), .ZN(new_n339));
  AOI21_X1  g153(.A(new_n331), .B1(new_n258), .B2(new_n339), .ZN(new_n340));
  XNOR2_X1  g154(.A(G110), .B(G122), .ZN(new_n341));
  AOI21_X1  g155(.A(new_n314), .B1(new_n340), .B2(new_n341), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n258), .A2(new_n339), .ZN(new_n343));
  INV_X1    g157(.A(new_n331), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  INV_X1    g159(.A(new_n341), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n345), .A2(new_n346), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n342), .A2(new_n347), .ZN(new_n348));
  NAND3_X1  g162(.A1(new_n345), .A2(new_n314), .A3(new_n346), .ZN(new_n349));
  INV_X1    g163(.A(G125), .ZN(new_n350));
  OAI211_X1 g164(.A(new_n350), .B(new_n230), .C1(new_n239), .C2(new_n241), .ZN(new_n351));
  OAI21_X1  g165(.A(new_n235), .B1(new_n231), .B2(G143), .ZN(new_n352));
  AOI22_X1  g166(.A1(new_n352), .A2(new_n262), .B1(new_n232), .B2(new_n259), .ZN(new_n353));
  OAI21_X1  g167(.A(new_n351), .B1(new_n353), .B2(new_n350), .ZN(new_n354));
  INV_X1    g168(.A(G224), .ZN(new_n355));
  NOR2_X1   g169(.A1(new_n355), .A2(G953), .ZN(new_n356));
  XNOR2_X1  g170(.A(new_n354), .B(new_n356), .ZN(new_n357));
  NAND3_X1  g171(.A1(new_n348), .A2(new_n349), .A3(new_n357), .ZN(new_n358));
  XOR2_X1   g172(.A(new_n341), .B(KEYINPUT8), .Z(new_n359));
  OAI21_X1  g173(.A(new_n322), .B1(new_n321), .B2(new_n330), .ZN(new_n360));
  AOI21_X1  g174(.A(new_n359), .B1(new_n344), .B2(new_n360), .ZN(new_n361));
  INV_X1    g175(.A(KEYINPUT7), .ZN(new_n362));
  NOR2_X1   g176(.A1(new_n356), .A2(new_n362), .ZN(new_n363));
  OR2_X1    g177(.A1(new_n351), .A2(KEYINPUT84), .ZN(new_n364));
  OAI21_X1  g178(.A(new_n260), .B1(new_n241), .B2(new_n263), .ZN(new_n365));
  AOI22_X1  g179(.A1(new_n351), .A2(KEYINPUT84), .B1(new_n365), .B2(G125), .ZN(new_n366));
  AOI21_X1  g180(.A(new_n363), .B1(new_n364), .B2(new_n366), .ZN(new_n367));
  NOR3_X1   g181(.A1(new_n354), .A2(new_n362), .A3(new_n356), .ZN(new_n368));
  NOR3_X1   g182(.A1(new_n361), .A2(new_n367), .A3(new_n368), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n340), .A2(new_n341), .ZN(new_n370));
  AOI21_X1  g184(.A(G902), .B1(new_n369), .B2(new_n370), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n358), .A2(new_n371), .ZN(new_n372));
  OAI21_X1  g186(.A(G210), .B1(G237), .B2(G902), .ZN(new_n373));
  INV_X1    g187(.A(new_n373), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n372), .A2(new_n374), .ZN(new_n375));
  NAND3_X1  g189(.A1(new_n358), .A2(new_n371), .A3(new_n373), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n375), .A2(new_n376), .ZN(new_n377));
  OAI21_X1  g191(.A(G214), .B1(G237), .B2(G902), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n377), .A2(new_n378), .ZN(new_n379));
  INV_X1    g193(.A(KEYINPUT20), .ZN(new_n380));
  INV_X1    g194(.A(KEYINPUT16), .ZN(new_n381));
  INV_X1    g195(.A(G140), .ZN(new_n382));
  NAND3_X1  g196(.A1(new_n381), .A2(new_n382), .A3(G125), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n382), .A2(G125), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n350), .A2(G140), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n384), .A2(new_n385), .ZN(new_n386));
  OAI21_X1  g200(.A(new_n383), .B1(new_n386), .B2(new_n381), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n387), .A2(new_n221), .ZN(new_n388));
  OAI211_X1 g202(.A(G146), .B(new_n383), .C1(new_n386), .C2(new_n381), .ZN(new_n389));
  INV_X1    g203(.A(G237), .ZN(new_n390));
  NAND3_X1  g204(.A1(new_n390), .A2(new_n288), .A3(G214), .ZN(new_n391));
  NOR2_X1   g205(.A1(new_n391), .A2(new_n233), .ZN(new_n392));
  NOR2_X1   g206(.A1(G237), .A2(G953), .ZN(new_n393));
  AOI21_X1  g207(.A(G143), .B1(new_n393), .B2(G214), .ZN(new_n394));
  OAI211_X1 g208(.A(KEYINPUT17), .B(G131), .C1(new_n392), .C2(new_n394), .ZN(new_n395));
  NAND3_X1  g209(.A1(new_n388), .A2(new_n389), .A3(new_n395), .ZN(new_n396));
  INV_X1    g210(.A(KEYINPUT88), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n396), .A2(new_n397), .ZN(new_n398));
  NAND4_X1  g212(.A1(new_n388), .A2(new_n395), .A3(KEYINPUT88), .A4(new_n389), .ZN(new_n399));
  OAI21_X1  g213(.A(G131), .B1(new_n392), .B2(new_n394), .ZN(new_n400));
  INV_X1    g214(.A(KEYINPUT17), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n391), .A2(new_n233), .ZN(new_n402));
  INV_X1    g216(.A(G131), .ZN(new_n403));
  NAND3_X1  g217(.A1(new_n393), .A2(G143), .A3(G214), .ZN(new_n404));
  NAND3_X1  g218(.A1(new_n402), .A2(new_n403), .A3(new_n404), .ZN(new_n405));
  NAND3_X1  g219(.A1(new_n400), .A2(new_n401), .A3(new_n405), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n406), .A2(KEYINPUT89), .ZN(new_n407));
  INV_X1    g221(.A(KEYINPUT89), .ZN(new_n408));
  NAND4_X1  g222(.A1(new_n400), .A2(new_n408), .A3(new_n401), .A4(new_n405), .ZN(new_n409));
  NAND4_X1  g223(.A1(new_n398), .A2(new_n399), .A3(new_n407), .A4(new_n409), .ZN(new_n410));
  XNOR2_X1  g224(.A(G113), .B(G122), .ZN(new_n411));
  XNOR2_X1  g225(.A(new_n411), .B(new_n209), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n386), .A2(KEYINPUT75), .ZN(new_n413));
  XNOR2_X1  g227(.A(G125), .B(G140), .ZN(new_n414));
  INV_X1    g228(.A(KEYINPUT75), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n414), .A2(new_n415), .ZN(new_n416));
  NAND3_X1  g230(.A1(new_n413), .A2(new_n416), .A3(new_n231), .ZN(new_n417));
  OAI21_X1  g231(.A(new_n417), .B1(new_n221), .B2(new_n414), .ZN(new_n418));
  AOI21_X1  g232(.A(new_n403), .B1(new_n402), .B2(new_n404), .ZN(new_n419));
  NAND3_X1  g233(.A1(new_n419), .A2(KEYINPUT85), .A3(KEYINPUT18), .ZN(new_n420));
  NAND3_X1  g234(.A1(KEYINPUT85), .A2(KEYINPUT18), .A3(G131), .ZN(new_n421));
  NAND3_X1  g235(.A1(new_n402), .A2(new_n404), .A3(new_n421), .ZN(new_n422));
  NAND3_X1  g236(.A1(new_n418), .A2(new_n420), .A3(new_n422), .ZN(new_n423));
  NAND3_X1  g237(.A1(new_n410), .A2(new_n412), .A3(new_n423), .ZN(new_n424));
  INV_X1    g238(.A(KEYINPUT86), .ZN(new_n425));
  NOR3_X1   g239(.A1(new_n392), .A2(new_n394), .A3(G131), .ZN(new_n426));
  OAI21_X1  g240(.A(new_n425), .B1(new_n426), .B2(new_n419), .ZN(new_n427));
  NAND3_X1  g241(.A1(new_n400), .A2(KEYINPUT86), .A3(new_n405), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n427), .A2(new_n428), .ZN(new_n429));
  INV_X1    g243(.A(KEYINPUT87), .ZN(new_n430));
  AOI21_X1  g244(.A(new_n415), .B1(new_n430), .B2(KEYINPUT19), .ZN(new_n431));
  NOR2_X1   g245(.A1(new_n386), .A2(new_n431), .ZN(new_n432));
  OAI21_X1  g246(.A(new_n430), .B1(new_n414), .B2(new_n415), .ZN(new_n433));
  INV_X1    g247(.A(KEYINPUT19), .ZN(new_n434));
  AOI21_X1  g248(.A(new_n432), .B1(new_n433), .B2(new_n434), .ZN(new_n435));
  OAI21_X1  g249(.A(new_n389), .B1(new_n435), .B2(new_n240), .ZN(new_n436));
  OAI21_X1  g250(.A(new_n423), .B1(new_n429), .B2(new_n436), .ZN(new_n437));
  INV_X1    g251(.A(new_n412), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n437), .A2(new_n438), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n424), .A2(new_n439), .ZN(new_n440));
  NOR2_X1   g254(.A1(G475), .A2(G902), .ZN(new_n441));
  AOI21_X1  g255(.A(new_n380), .B1(new_n440), .B2(new_n441), .ZN(new_n442));
  INV_X1    g256(.A(new_n441), .ZN(new_n443));
  AOI211_X1 g257(.A(KEYINPUT20), .B(new_n443), .C1(new_n424), .C2(new_n439), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n410), .A2(new_n423), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n445), .A2(new_n438), .ZN(new_n446));
  AOI21_X1  g260(.A(G902), .B1(new_n446), .B2(new_n424), .ZN(new_n447));
  INV_X1    g261(.A(G475), .ZN(new_n448));
  OAI22_X1  g262(.A1(new_n442), .A2(new_n444), .B1(new_n447), .B2(new_n448), .ZN(new_n449));
  INV_X1    g263(.A(new_n449), .ZN(new_n450));
  INV_X1    g264(.A(G478), .ZN(new_n451));
  NOR2_X1   g265(.A1(KEYINPUT93), .A2(KEYINPUT15), .ZN(new_n452));
  INV_X1    g266(.A(new_n452), .ZN(new_n453));
  NAND2_X1  g267(.A1(KEYINPUT93), .A2(KEYINPUT15), .ZN(new_n454));
  AOI21_X1  g268(.A(new_n451), .B1(new_n453), .B2(new_n454), .ZN(new_n455));
  INV_X1    g269(.A(new_n455), .ZN(new_n456));
  NAND3_X1  g270(.A1(new_n323), .A2(new_n325), .A3(G122), .ZN(new_n457));
  INV_X1    g271(.A(KEYINPUT14), .ZN(new_n458));
  OR2_X1    g272(.A1(new_n315), .A2(G122), .ZN(new_n459));
  NAND3_X1  g273(.A1(new_n457), .A2(new_n458), .A3(new_n459), .ZN(new_n460));
  NAND3_X1  g274(.A1(new_n319), .A2(KEYINPUT14), .A3(G122), .ZN(new_n461));
  NAND3_X1  g275(.A1(new_n460), .A2(G107), .A3(new_n461), .ZN(new_n462));
  INV_X1    g276(.A(KEYINPUT92), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  NAND4_X1  g278(.A1(new_n460), .A2(KEYINPUT92), .A3(G107), .A4(new_n461), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  XNOR2_X1  g280(.A(G128), .B(G143), .ZN(new_n467));
  XNOR2_X1  g281(.A(new_n467), .B(new_n193), .ZN(new_n468));
  INV_X1    g282(.A(KEYINPUT91), .ZN(new_n469));
  NAND4_X1  g283(.A1(new_n457), .A2(new_n469), .A3(new_n212), .A4(new_n459), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n457), .A2(new_n459), .ZN(new_n471));
  OAI21_X1  g285(.A(KEYINPUT91), .B1(new_n471), .B2(G107), .ZN(new_n472));
  NAND4_X1  g286(.A1(new_n466), .A2(new_n468), .A3(new_n470), .A4(new_n472), .ZN(new_n473));
  OR2_X1    g287(.A1(new_n467), .A2(G134), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n467), .A2(G134), .ZN(new_n475));
  XNOR2_X1  g289(.A(KEYINPUT90), .B(KEYINPUT13), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n228), .A2(G143), .ZN(new_n477));
  NAND3_X1  g291(.A1(new_n476), .A2(G134), .A3(new_n477), .ZN(new_n478));
  NAND3_X1  g292(.A1(new_n474), .A2(new_n475), .A3(new_n478), .ZN(new_n479));
  NAND4_X1  g293(.A1(new_n467), .A2(new_n476), .A3(G134), .A4(new_n477), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  XNOR2_X1  g295(.A(new_n471), .B(new_n212), .ZN(new_n482));
  NOR2_X1   g296(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  INV_X1    g297(.A(new_n483), .ZN(new_n484));
  INV_X1    g298(.A(G217), .ZN(new_n485));
  NOR3_X1   g299(.A1(new_n188), .A2(new_n485), .A3(G953), .ZN(new_n486));
  NAND3_X1  g300(.A1(new_n473), .A2(new_n484), .A3(new_n486), .ZN(new_n487));
  INV_X1    g301(.A(new_n486), .ZN(new_n488));
  NAND3_X1  g302(.A1(new_n472), .A2(new_n468), .A3(new_n470), .ZN(new_n489));
  AOI21_X1  g303(.A(new_n489), .B1(new_n464), .B2(new_n465), .ZN(new_n490));
  OAI21_X1  g304(.A(new_n488), .B1(new_n490), .B2(new_n483), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n487), .A2(new_n491), .ZN(new_n492));
  AOI21_X1  g306(.A(new_n456), .B1(new_n492), .B2(new_n190), .ZN(new_n493));
  INV_X1    g307(.A(new_n493), .ZN(new_n494));
  NAND3_X1  g308(.A1(new_n492), .A2(new_n190), .A3(new_n456), .ZN(new_n495));
  NAND3_X1  g309(.A1(new_n494), .A2(KEYINPUT94), .A3(new_n495), .ZN(new_n496));
  INV_X1    g310(.A(KEYINPUT94), .ZN(new_n497));
  AOI211_X1 g311(.A(G902), .B(new_n455), .C1(new_n487), .C2(new_n491), .ZN(new_n498));
  OAI21_X1  g312(.A(new_n497), .B1(new_n493), .B2(new_n498), .ZN(new_n499));
  INV_X1    g313(.A(G952), .ZN(new_n500));
  NOR2_X1   g314(.A1(new_n500), .A2(G953), .ZN(new_n501));
  NAND2_X1  g315(.A1(G234), .A2(G237), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  XNOR2_X1  g317(.A(KEYINPUT21), .B(G898), .ZN(new_n504));
  INV_X1    g318(.A(new_n504), .ZN(new_n505));
  NAND3_X1  g319(.A1(new_n502), .A2(G902), .A3(G953), .ZN(new_n506));
  OAI21_X1  g320(.A(new_n503), .B1(new_n505), .B2(new_n506), .ZN(new_n507));
  NAND4_X1  g321(.A1(new_n450), .A2(new_n496), .A3(new_n499), .A4(new_n507), .ZN(new_n508));
  NOR2_X1   g322(.A1(new_n379), .A2(new_n508), .ZN(new_n509));
  AOI21_X1  g323(.A(new_n485), .B1(G234), .B2(new_n190), .ZN(new_n510));
  INV_X1    g324(.A(new_n510), .ZN(new_n511));
  XNOR2_X1  g325(.A(KEYINPUT24), .B(G110), .ZN(new_n512));
  INV_X1    g326(.A(KEYINPUT74), .ZN(new_n513));
  XNOR2_X1  g327(.A(new_n512), .B(new_n513), .ZN(new_n514));
  XNOR2_X1  g328(.A(G119), .B(G128), .ZN(new_n515));
  NOR2_X1   g329(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  INV_X1    g330(.A(KEYINPUT23), .ZN(new_n517));
  INV_X1    g331(.A(G119), .ZN(new_n518));
  OAI21_X1  g332(.A(new_n517), .B1(new_n518), .B2(G128), .ZN(new_n519));
  NAND3_X1  g333(.A1(new_n228), .A2(KEYINPUT23), .A3(G119), .ZN(new_n520));
  OAI211_X1 g334(.A(new_n519), .B(new_n520), .C1(G119), .C2(new_n228), .ZN(new_n521));
  NOR2_X1   g335(.A1(new_n521), .A2(G110), .ZN(new_n522));
  OAI211_X1 g336(.A(new_n417), .B(new_n389), .C1(new_n516), .C2(new_n522), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n388), .A2(new_n389), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n514), .A2(new_n515), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n521), .A2(G110), .ZN(new_n526));
  NAND3_X1  g340(.A1(new_n524), .A2(new_n525), .A3(new_n526), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n523), .A2(new_n527), .ZN(new_n528));
  XNOR2_X1  g342(.A(KEYINPUT22), .B(G137), .ZN(new_n529));
  NAND3_X1  g343(.A1(new_n288), .A2(G221), .A3(G234), .ZN(new_n530));
  XNOR2_X1  g344(.A(new_n529), .B(new_n530), .ZN(new_n531));
  INV_X1    g345(.A(new_n531), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n528), .A2(new_n532), .ZN(new_n533));
  NAND3_X1  g347(.A1(new_n523), .A2(new_n527), .A3(new_n531), .ZN(new_n534));
  NAND3_X1  g348(.A1(new_n533), .A2(new_n190), .A3(new_n534), .ZN(new_n535));
  INV_X1    g349(.A(KEYINPUT25), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  NAND4_X1  g351(.A1(new_n533), .A2(KEYINPUT25), .A3(new_n190), .A4(new_n534), .ZN(new_n538));
  AOI21_X1  g352(.A(new_n511), .B1(new_n537), .B2(new_n538), .ZN(new_n539));
  INV_X1    g353(.A(new_n533), .ZN(new_n540));
  INV_X1    g354(.A(new_n534), .ZN(new_n541));
  NOR2_X1   g355(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  NOR2_X1   g356(.A1(new_n510), .A2(G902), .ZN(new_n543));
  AOI21_X1  g357(.A(new_n539), .B1(new_n542), .B2(new_n543), .ZN(new_n544));
  INV_X1    g358(.A(new_n544), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n335), .A2(new_n338), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n205), .A2(new_n353), .ZN(new_n547));
  INV_X1    g361(.A(KEYINPUT30), .ZN(new_n548));
  XNOR2_X1  g362(.A(G134), .B(G137), .ZN(new_n549));
  OAI21_X1  g363(.A(KEYINPUT66), .B1(new_n549), .B2(new_n403), .ZN(new_n550));
  INV_X1    g364(.A(KEYINPUT66), .ZN(new_n551));
  NOR2_X1   g365(.A1(new_n193), .A2(G137), .ZN(new_n552));
  NOR2_X1   g366(.A1(new_n196), .A2(G134), .ZN(new_n553));
  OAI211_X1 g367(.A(new_n551), .B(G131), .C1(new_n552), .C2(new_n553), .ZN(new_n554));
  AOI22_X1  g368(.A1(new_n200), .A2(new_n201), .B1(new_n550), .B2(new_n554), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n555), .A2(new_n242), .ZN(new_n556));
  AND3_X1   g370(.A1(new_n547), .A2(new_n548), .A3(new_n556), .ZN(new_n557));
  AOI21_X1  g371(.A(new_n548), .B1(new_n547), .B2(new_n556), .ZN(new_n558));
  OAI21_X1  g372(.A(new_n546), .B1(new_n557), .B2(new_n558), .ZN(new_n559));
  XNOR2_X1  g373(.A(KEYINPUT26), .B(G101), .ZN(new_n560));
  XNOR2_X1  g374(.A(KEYINPUT69), .B(KEYINPUT27), .ZN(new_n561));
  XNOR2_X1  g375(.A(new_n560), .B(new_n561), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n393), .A2(G210), .ZN(new_n563));
  XNOR2_X1  g377(.A(new_n563), .B(KEYINPUT70), .ZN(new_n564));
  XOR2_X1   g378(.A(new_n562), .B(new_n564), .Z(new_n565));
  NAND4_X1  g379(.A1(new_n547), .A2(new_n556), .A3(new_n335), .A4(new_n338), .ZN(new_n566));
  NAND3_X1  g380(.A1(new_n559), .A2(new_n565), .A3(new_n566), .ZN(new_n567));
  INV_X1    g381(.A(KEYINPUT31), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  NAND4_X1  g383(.A1(new_n559), .A2(KEYINPUT31), .A3(new_n565), .A4(new_n566), .ZN(new_n570));
  INV_X1    g384(.A(KEYINPUT28), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n566), .A2(new_n571), .ZN(new_n572));
  AND2_X1   g386(.A1(new_n555), .A2(new_n242), .ZN(new_n573));
  NOR2_X1   g387(.A1(new_n272), .A2(new_n365), .ZN(new_n574));
  OAI21_X1  g388(.A(new_n546), .B1(new_n573), .B2(new_n574), .ZN(new_n575));
  INV_X1    g389(.A(KEYINPUT71), .ZN(new_n576));
  AND3_X1   g390(.A1(new_n575), .A2(new_n576), .A3(new_n566), .ZN(new_n577));
  OAI21_X1  g391(.A(KEYINPUT28), .B1(new_n575), .B2(new_n576), .ZN(new_n578));
  OAI21_X1  g392(.A(new_n572), .B1(new_n577), .B2(new_n578), .ZN(new_n579));
  INV_X1    g393(.A(new_n565), .ZN(new_n580));
  AOI22_X1  g394(.A1(new_n569), .A2(new_n570), .B1(new_n579), .B2(new_n580), .ZN(new_n581));
  NOR2_X1   g395(.A1(G472), .A2(G902), .ZN(new_n582));
  INV_X1    g396(.A(new_n582), .ZN(new_n583));
  OAI21_X1  g397(.A(KEYINPUT32), .B1(new_n581), .B2(new_n583), .ZN(new_n584));
  INV_X1    g398(.A(new_n566), .ZN(new_n585));
  OAI21_X1  g399(.A(KEYINPUT30), .B1(new_n573), .B2(new_n574), .ZN(new_n586));
  NAND3_X1  g400(.A1(new_n547), .A2(new_n548), .A3(new_n556), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  AOI21_X1  g402(.A(new_n585), .B1(new_n588), .B2(new_n546), .ZN(new_n589));
  AOI21_X1  g403(.A(KEYINPUT31), .B1(new_n589), .B2(new_n565), .ZN(new_n590));
  INV_X1    g404(.A(new_n546), .ZN(new_n591));
  AOI21_X1  g405(.A(new_n591), .B1(new_n586), .B2(new_n587), .ZN(new_n592));
  NOR4_X1   g406(.A1(new_n592), .A2(new_n568), .A3(new_n580), .A4(new_n585), .ZN(new_n593));
  AOI22_X1  g407(.A1(new_n547), .A2(new_n556), .B1(new_n335), .B2(new_n338), .ZN(new_n594));
  AOI21_X1  g408(.A(new_n571), .B1(new_n594), .B2(KEYINPUT71), .ZN(new_n595));
  NAND3_X1  g409(.A1(new_n575), .A2(new_n576), .A3(new_n566), .ZN(new_n596));
  AOI22_X1  g410(.A1(new_n595), .A2(new_n596), .B1(new_n571), .B2(new_n566), .ZN(new_n597));
  OAI22_X1  g411(.A1(new_n590), .A2(new_n593), .B1(new_n565), .B2(new_n597), .ZN(new_n598));
  INV_X1    g412(.A(KEYINPUT32), .ZN(new_n599));
  NAND3_X1  g413(.A1(new_n598), .A2(new_n599), .A3(new_n582), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n584), .A2(new_n600), .ZN(new_n601));
  INV_X1    g415(.A(KEYINPUT72), .ZN(new_n602));
  NAND3_X1  g416(.A1(new_n575), .A2(new_n602), .A3(new_n566), .ZN(new_n603));
  OAI211_X1 g417(.A(KEYINPUT72), .B(new_n546), .C1(new_n573), .C2(new_n574), .ZN(new_n604));
  NAND3_X1  g418(.A1(new_n603), .A2(KEYINPUT28), .A3(new_n604), .ZN(new_n605));
  AND2_X1   g419(.A1(new_n565), .A2(KEYINPUT29), .ZN(new_n606));
  NAND3_X1  g420(.A1(new_n605), .A2(new_n572), .A3(new_n606), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n607), .A2(KEYINPUT73), .ZN(new_n608));
  INV_X1    g422(.A(KEYINPUT73), .ZN(new_n609));
  NAND4_X1  g423(.A1(new_n605), .A2(new_n609), .A3(new_n572), .A4(new_n606), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n608), .A2(new_n610), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n559), .A2(new_n566), .ZN(new_n612));
  AOI21_X1  g426(.A(KEYINPUT29), .B1(new_n612), .B2(new_n580), .ZN(new_n613));
  OAI211_X1 g427(.A(new_n565), .B(new_n572), .C1(new_n577), .C2(new_n578), .ZN(new_n614));
  AOI21_X1  g428(.A(G902), .B1(new_n613), .B2(new_n614), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n611), .A2(new_n615), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n616), .A2(G472), .ZN(new_n617));
  AOI21_X1  g431(.A(new_n545), .B1(new_n601), .B2(new_n617), .ZN(new_n618));
  NAND3_X1  g432(.A1(new_n313), .A2(new_n509), .A3(new_n618), .ZN(new_n619));
  XNOR2_X1  g433(.A(new_n619), .B(G101), .ZN(G3));
  INV_X1    g434(.A(G472), .ZN(new_n621));
  AOI21_X1  g435(.A(new_n621), .B1(new_n598), .B2(new_n190), .ZN(new_n622));
  AOI21_X1  g436(.A(new_n622), .B1(new_n598), .B2(new_n582), .ZN(new_n623));
  NAND3_X1  g437(.A1(new_n313), .A2(new_n544), .A3(new_n623), .ZN(new_n624));
  OAI21_X1  g438(.A(new_n378), .B1(new_n376), .B2(KEYINPUT95), .ZN(new_n625));
  INV_X1    g439(.A(new_n625), .ZN(new_n626));
  NAND3_X1  g440(.A1(new_n375), .A2(KEYINPUT95), .A3(new_n376), .ZN(new_n627));
  AOI21_X1  g441(.A(G478), .B1(new_n492), .B2(new_n190), .ZN(new_n628));
  INV_X1    g442(.A(new_n628), .ZN(new_n629));
  NOR2_X1   g443(.A1(KEYINPUT96), .A2(KEYINPUT33), .ZN(new_n630));
  INV_X1    g444(.A(new_n630), .ZN(new_n631));
  INV_X1    g445(.A(KEYINPUT96), .ZN(new_n632));
  INV_X1    g446(.A(KEYINPUT33), .ZN(new_n633));
  NOR2_X1   g447(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  INV_X1    g448(.A(new_n634), .ZN(new_n635));
  NAND3_X1  g449(.A1(new_n492), .A2(new_n631), .A3(new_n635), .ZN(new_n636));
  NAND4_X1  g450(.A1(new_n487), .A2(new_n491), .A3(new_n632), .A4(new_n633), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  NOR2_X1   g452(.A1(new_n451), .A2(G902), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  INV_X1    g454(.A(new_n442), .ZN(new_n641));
  NAND3_X1  g455(.A1(new_n440), .A2(new_n380), .A3(new_n441), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  INV_X1    g457(.A(new_n447), .ZN(new_n644));
  NAND2_X1  g458(.A1(new_n644), .A2(G475), .ZN(new_n645));
  AOI22_X1  g459(.A1(new_n629), .A2(new_n640), .B1(new_n643), .B2(new_n645), .ZN(new_n646));
  AND4_X1   g460(.A1(new_n507), .A2(new_n626), .A3(new_n627), .A4(new_n646), .ZN(new_n647));
  INV_X1    g461(.A(new_n647), .ZN(new_n648));
  NOR2_X1   g462(.A1(new_n624), .A2(new_n648), .ZN(new_n649));
  XNOR2_X1  g463(.A(new_n649), .B(KEYINPUT97), .ZN(new_n650));
  XOR2_X1   g464(.A(KEYINPUT34), .B(G104), .Z(new_n651));
  XNOR2_X1  g465(.A(new_n650), .B(new_n651), .ZN(G6));
  NAND2_X1  g466(.A1(new_n496), .A2(new_n499), .ZN(new_n653));
  XOR2_X1   g467(.A(new_n507), .B(KEYINPUT99), .Z(new_n654));
  AND2_X1   g468(.A1(new_n645), .A2(new_n654), .ZN(new_n655));
  NAND3_X1  g469(.A1(new_n641), .A2(KEYINPUT98), .A3(new_n642), .ZN(new_n656));
  INV_X1    g470(.A(KEYINPUT98), .ZN(new_n657));
  OAI21_X1  g471(.A(new_n657), .B1(new_n442), .B2(new_n444), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n656), .A2(new_n658), .ZN(new_n659));
  AND3_X1   g473(.A1(new_n653), .A2(new_n655), .A3(new_n659), .ZN(new_n660));
  AND3_X1   g474(.A1(new_n660), .A2(new_n627), .A3(new_n626), .ZN(new_n661));
  INV_X1    g475(.A(new_n661), .ZN(new_n662));
  NOR2_X1   g476(.A1(new_n624), .A2(new_n662), .ZN(new_n663));
  XNOR2_X1  g477(.A(KEYINPUT35), .B(G107), .ZN(new_n664));
  XNOR2_X1  g478(.A(new_n663), .B(new_n664), .ZN(G9));
  INV_X1    g479(.A(new_n539), .ZN(new_n666));
  NAND2_X1  g480(.A1(new_n528), .A2(KEYINPUT100), .ZN(new_n667));
  INV_X1    g481(.A(KEYINPUT100), .ZN(new_n668));
  NAND3_X1  g482(.A1(new_n523), .A2(new_n668), .A3(new_n527), .ZN(new_n669));
  NAND2_X1  g483(.A1(new_n667), .A2(new_n669), .ZN(new_n670));
  OAI21_X1  g484(.A(new_n670), .B1(KEYINPUT36), .B2(new_n532), .ZN(new_n671));
  NOR2_X1   g485(.A1(new_n532), .A2(KEYINPUT36), .ZN(new_n672));
  NAND3_X1  g486(.A1(new_n667), .A2(new_n672), .A3(new_n669), .ZN(new_n673));
  NAND2_X1  g487(.A1(new_n671), .A2(new_n673), .ZN(new_n674));
  NAND2_X1  g488(.A1(new_n674), .A2(new_n543), .ZN(new_n675));
  NAND3_X1  g489(.A1(new_n666), .A2(new_n675), .A3(KEYINPUT101), .ZN(new_n676));
  INV_X1    g490(.A(KEYINPUT101), .ZN(new_n677));
  INV_X1    g491(.A(new_n543), .ZN(new_n678));
  AOI21_X1  g492(.A(new_n678), .B1(new_n671), .B2(new_n673), .ZN(new_n679));
  OAI21_X1  g493(.A(new_n677), .B1(new_n679), .B2(new_n539), .ZN(new_n680));
  NAND2_X1  g494(.A1(new_n676), .A2(new_n680), .ZN(new_n681));
  INV_X1    g495(.A(new_n681), .ZN(new_n682));
  NAND4_X1  g496(.A1(new_n313), .A2(new_n509), .A3(new_n623), .A4(new_n682), .ZN(new_n683));
  XOR2_X1   g497(.A(KEYINPUT37), .B(G110), .Z(new_n684));
  XNOR2_X1  g498(.A(new_n683), .B(new_n684), .ZN(G12));
  AND3_X1   g499(.A1(new_n358), .A2(new_n371), .A3(new_n373), .ZN(new_n686));
  AOI21_X1  g500(.A(new_n373), .B1(new_n358), .B2(new_n371), .ZN(new_n687));
  NOR2_X1   g501(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  AOI21_X1  g502(.A(new_n625), .B1(new_n688), .B2(KEYINPUT95), .ZN(new_n689));
  AOI21_X1  g503(.A(new_n681), .B1(new_n601), .B2(new_n617), .ZN(new_n690));
  OR2_X1    g504(.A1(new_n506), .A2(G900), .ZN(new_n691));
  NAND2_X1  g505(.A1(new_n691), .A2(new_n503), .ZN(new_n692));
  INV_X1    g506(.A(new_n692), .ZN(new_n693));
  AOI21_X1  g507(.A(new_n693), .B1(new_n644), .B2(G475), .ZN(new_n694));
  AND3_X1   g508(.A1(new_n653), .A2(new_n659), .A3(new_n694), .ZN(new_n695));
  NAND4_X1  g509(.A1(new_n313), .A2(new_n689), .A3(new_n690), .A4(new_n695), .ZN(new_n696));
  XNOR2_X1  g510(.A(new_n696), .B(G128), .ZN(G30));
  XNOR2_X1  g511(.A(KEYINPUT102), .B(KEYINPUT38), .ZN(new_n698));
  XNOR2_X1  g512(.A(new_n688), .B(new_n698), .ZN(new_n699));
  NOR2_X1   g513(.A1(new_n679), .A2(new_n539), .ZN(new_n700));
  INV_X1    g514(.A(new_n700), .ZN(new_n701));
  NAND2_X1  g515(.A1(new_n612), .A2(new_n565), .ZN(new_n702));
  AND2_X1   g516(.A1(new_n603), .A2(new_n604), .ZN(new_n703));
  OAI211_X1 g517(.A(new_n702), .B(new_n190), .C1(new_n565), .C2(new_n703), .ZN(new_n704));
  NAND2_X1  g518(.A1(new_n704), .A2(G472), .ZN(new_n705));
  AOI21_X1  g519(.A(new_n701), .B1(new_n601), .B2(new_n705), .ZN(new_n706));
  AOI21_X1  g520(.A(new_n450), .B1(new_n496), .B2(new_n499), .ZN(new_n707));
  NAND4_X1  g521(.A1(new_n699), .A2(new_n378), .A3(new_n706), .A4(new_n707), .ZN(new_n708));
  XOR2_X1   g522(.A(new_n708), .B(KEYINPUT103), .Z(new_n709));
  XNOR2_X1  g523(.A(new_n692), .B(KEYINPUT39), .ZN(new_n710));
  NAND2_X1  g524(.A1(new_n313), .A2(new_n710), .ZN(new_n711));
  XNOR2_X1  g525(.A(new_n711), .B(KEYINPUT40), .ZN(new_n712));
  OR3_X1    g526(.A1(new_n709), .A2(KEYINPUT104), .A3(new_n712), .ZN(new_n713));
  OAI21_X1  g527(.A(KEYINPUT104), .B1(new_n709), .B2(new_n712), .ZN(new_n714));
  NAND2_X1  g528(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  XNOR2_X1  g529(.A(new_n715), .B(new_n233), .ZN(G45));
  INV_X1    g530(.A(KEYINPUT105), .ZN(new_n717));
  NAND4_X1  g531(.A1(new_n689), .A2(new_n717), .A3(new_n646), .A4(new_n692), .ZN(new_n718));
  NAND4_X1  g532(.A1(new_n626), .A2(new_n627), .A3(new_n646), .A4(new_n692), .ZN(new_n719));
  NAND2_X1  g533(.A1(new_n719), .A2(KEYINPUT105), .ZN(new_n720));
  NAND4_X1  g534(.A1(new_n718), .A2(new_n720), .A3(new_n313), .A4(new_n690), .ZN(new_n721));
  XNOR2_X1  g535(.A(new_n721), .B(G146), .ZN(G48));
  AND3_X1   g536(.A1(new_n305), .A2(new_n306), .A3(new_n190), .ZN(new_n723));
  AOI21_X1  g537(.A(new_n306), .B1(new_n305), .B2(new_n190), .ZN(new_n724));
  NOR3_X1   g538(.A1(new_n723), .A2(new_n724), .A3(new_n191), .ZN(new_n725));
  NAND3_X1  g539(.A1(new_n725), .A2(new_n618), .A3(new_n647), .ZN(new_n726));
  XNOR2_X1  g540(.A(KEYINPUT41), .B(G113), .ZN(new_n727));
  XNOR2_X1  g541(.A(new_n726), .B(new_n727), .ZN(G15));
  NAND3_X1  g542(.A1(new_n725), .A2(new_n618), .A3(new_n661), .ZN(new_n729));
  XNOR2_X1  g543(.A(new_n729), .B(G116), .ZN(G18));
  AOI211_X1 g544(.A(new_n508), .B(new_n681), .C1(new_n601), .C2(new_n617), .ZN(new_n731));
  NAND3_X1  g545(.A1(new_n731), .A2(new_n725), .A3(new_n689), .ZN(new_n732));
  XOR2_X1   g546(.A(KEYINPUT106), .B(G119), .Z(new_n733));
  XNOR2_X1  g547(.A(new_n732), .B(new_n733), .ZN(G21));
  OAI21_X1  g548(.A(G472), .B1(new_n581), .B2(G902), .ZN(new_n735));
  NOR2_X1   g549(.A1(new_n590), .A2(new_n593), .ZN(new_n736));
  INV_X1    g550(.A(KEYINPUT107), .ZN(new_n737));
  NAND3_X1  g551(.A1(new_n605), .A2(new_n737), .A3(new_n572), .ZN(new_n738));
  NAND2_X1  g552(.A1(new_n605), .A2(new_n572), .ZN(new_n739));
  AOI21_X1  g553(.A(new_n565), .B1(new_n739), .B2(KEYINPUT107), .ZN(new_n740));
  AOI21_X1  g554(.A(new_n736), .B1(new_n738), .B2(new_n740), .ZN(new_n741));
  OAI211_X1 g555(.A(new_n735), .B(new_n544), .C1(new_n741), .C2(new_n583), .ZN(new_n742));
  INV_X1    g556(.A(KEYINPUT108), .ZN(new_n743));
  NAND2_X1  g557(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  NAND2_X1  g558(.A1(new_n740), .A2(new_n738), .ZN(new_n745));
  INV_X1    g559(.A(new_n736), .ZN(new_n746));
  NAND2_X1  g560(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  NAND2_X1  g561(.A1(new_n747), .A2(new_n582), .ZN(new_n748));
  NAND4_X1  g562(.A1(new_n748), .A2(KEYINPUT108), .A3(new_n544), .A4(new_n735), .ZN(new_n749));
  NAND2_X1  g563(.A1(new_n744), .A2(new_n749), .ZN(new_n750));
  AND4_X1   g564(.A1(new_n627), .A2(new_n626), .A3(new_n654), .A4(new_n707), .ZN(new_n751));
  NAND3_X1  g565(.A1(new_n750), .A2(new_n725), .A3(new_n751), .ZN(new_n752));
  XNOR2_X1  g566(.A(new_n752), .B(G122), .ZN(G24));
  NOR2_X1   g567(.A1(new_n303), .A2(KEYINPUT83), .ZN(new_n754));
  AOI22_X1  g568(.A1(new_n279), .A2(new_n282), .B1(new_n205), .B2(new_n292), .ZN(new_n755));
  OAI21_X1  g569(.A(new_n284), .B1(new_n755), .B2(new_n290), .ZN(new_n756));
  AOI21_X1  g570(.A(new_n754), .B1(new_n303), .B2(new_n756), .ZN(new_n757));
  OAI21_X1  g571(.A(G469), .B1(new_n757), .B2(G902), .ZN(new_n758));
  INV_X1    g572(.A(new_n191), .ZN(new_n759));
  NAND4_X1  g573(.A1(new_n689), .A2(new_n758), .A3(new_n759), .A4(new_n307), .ZN(new_n760));
  AOI21_X1  g574(.A(new_n583), .B1(new_n745), .B2(new_n746), .ZN(new_n761));
  NOR3_X1   g575(.A1(new_n761), .A2(new_n622), .A3(new_n700), .ZN(new_n762));
  INV_X1    g576(.A(new_n639), .ZN(new_n763));
  AOI21_X1  g577(.A(new_n763), .B1(new_n636), .B2(new_n637), .ZN(new_n764));
  OAI211_X1 g578(.A(new_n449), .B(new_n692), .C1(new_n628), .C2(new_n764), .ZN(new_n765));
  INV_X1    g579(.A(new_n765), .ZN(new_n766));
  NAND2_X1  g580(.A1(new_n762), .A2(new_n766), .ZN(new_n767));
  OAI21_X1  g581(.A(KEYINPUT109), .B1(new_n760), .B2(new_n767), .ZN(new_n768));
  INV_X1    g582(.A(KEYINPUT109), .ZN(new_n769));
  NOR4_X1   g583(.A1(new_n761), .A2(new_n622), .A3(new_n765), .A4(new_n700), .ZN(new_n770));
  NAND4_X1  g584(.A1(new_n725), .A2(new_n769), .A3(new_n689), .A4(new_n770), .ZN(new_n771));
  NAND2_X1  g585(.A1(new_n768), .A2(new_n771), .ZN(new_n772));
  XNOR2_X1  g586(.A(new_n772), .B(G125), .ZN(G27));
  INV_X1    g587(.A(KEYINPUT111), .ZN(new_n774));
  OAI21_X1  g588(.A(new_n774), .B1(new_n283), .B2(new_n290), .ZN(new_n775));
  OAI21_X1  g589(.A(new_n302), .B1(new_n294), .B2(new_n298), .ZN(new_n776));
  NAND3_X1  g590(.A1(new_n776), .A2(KEYINPUT111), .A3(new_n300), .ZN(new_n777));
  NAND4_X1  g591(.A1(new_n775), .A2(new_n777), .A3(G469), .A4(new_n308), .ZN(new_n778));
  XOR2_X1   g592(.A(new_n311), .B(KEYINPUT110), .Z(new_n779));
  AND2_X1   g593(.A1(new_n778), .A2(new_n779), .ZN(new_n780));
  NAND2_X1  g594(.A1(new_n780), .A2(new_n307), .ZN(new_n781));
  NAND4_X1  g595(.A1(new_n375), .A2(new_n759), .A3(new_n378), .A4(new_n376), .ZN(new_n782));
  INV_X1    g596(.A(new_n782), .ZN(new_n783));
  NAND4_X1  g597(.A1(new_n781), .A2(new_n618), .A3(new_n766), .A4(new_n783), .ZN(new_n784));
  INV_X1    g598(.A(KEYINPUT42), .ZN(new_n785));
  NAND2_X1  g599(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  AOI21_X1  g600(.A(new_n782), .B1(new_n780), .B2(new_n307), .ZN(new_n787));
  NAND4_X1  g601(.A1(new_n787), .A2(KEYINPUT42), .A3(new_n618), .A4(new_n766), .ZN(new_n788));
  NAND2_X1  g602(.A1(new_n786), .A2(new_n788), .ZN(new_n789));
  XNOR2_X1  g603(.A(new_n789), .B(G131), .ZN(G33));
  NAND4_X1  g604(.A1(new_n781), .A2(new_n618), .A3(new_n695), .A4(new_n783), .ZN(new_n791));
  XNOR2_X1  g605(.A(new_n791), .B(G134), .ZN(G36));
  INV_X1    g606(.A(new_n779), .ZN(new_n793));
  OAI21_X1  g607(.A(new_n308), .B1(new_n290), .B2(new_n283), .ZN(new_n794));
  INV_X1    g608(.A(KEYINPUT45), .ZN(new_n795));
  AOI21_X1  g609(.A(new_n306), .B1(new_n794), .B2(new_n795), .ZN(new_n796));
  NAND4_X1  g610(.A1(new_n775), .A2(new_n777), .A3(KEYINPUT45), .A4(new_n308), .ZN(new_n797));
  AOI21_X1  g611(.A(new_n793), .B1(new_n796), .B2(new_n797), .ZN(new_n798));
  AND2_X1   g612(.A1(new_n798), .A2(KEYINPUT46), .ZN(new_n799));
  OAI21_X1  g613(.A(new_n307), .B1(new_n798), .B2(KEYINPUT46), .ZN(new_n800));
  OAI211_X1 g614(.A(new_n759), .B(new_n710), .C1(new_n799), .C2(new_n800), .ZN(new_n801));
  INV_X1    g615(.A(new_n801), .ZN(new_n802));
  NOR2_X1   g616(.A1(new_n764), .A2(new_n628), .ZN(new_n803));
  NOR2_X1   g617(.A1(new_n803), .A2(new_n449), .ZN(new_n804));
  INV_X1    g618(.A(new_n804), .ZN(new_n805));
  NAND2_X1  g619(.A1(new_n805), .A2(KEYINPUT43), .ZN(new_n806));
  OR3_X1    g620(.A1(new_n803), .A2(KEYINPUT43), .A3(new_n449), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n806), .A2(new_n807), .ZN(new_n808));
  OR3_X1    g622(.A1(new_n808), .A2(new_n623), .A3(new_n700), .ZN(new_n809));
  INV_X1    g623(.A(KEYINPUT44), .ZN(new_n810));
  AND2_X1   g624(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  NAND3_X1  g625(.A1(new_n375), .A2(new_n378), .A3(new_n376), .ZN(new_n812));
  NOR2_X1   g626(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  OAI211_X1 g627(.A(new_n802), .B(new_n813), .C1(new_n810), .C2(new_n809), .ZN(new_n814));
  XNOR2_X1  g628(.A(new_n814), .B(G137), .ZN(G39));
  NAND2_X1  g629(.A1(new_n601), .A2(new_n617), .ZN(new_n816));
  OAI21_X1  g630(.A(new_n759), .B1(new_n799), .B2(new_n800), .ZN(new_n817));
  XNOR2_X1  g631(.A(new_n817), .B(KEYINPUT47), .ZN(new_n818));
  NAND2_X1  g632(.A1(new_n766), .A2(new_n545), .ZN(new_n819));
  OR4_X1    g633(.A1(new_n816), .A2(new_n818), .A3(new_n812), .A4(new_n819), .ZN(new_n820));
  XNOR2_X1  g634(.A(new_n820), .B(G140), .ZN(G42));
  NOR2_X1   g635(.A1(new_n493), .A2(new_n498), .ZN(new_n822));
  NOR2_X1   g636(.A1(new_n449), .A2(new_n822), .ZN(new_n823));
  OAI21_X1  g637(.A(new_n654), .B1(new_n646), .B2(new_n823), .ZN(new_n824));
  NOR2_X1   g638(.A1(new_n824), .A2(new_n379), .ZN(new_n825));
  NAND4_X1  g639(.A1(new_n825), .A2(new_n313), .A3(new_n544), .A4(new_n623), .ZN(new_n826));
  NAND3_X1  g640(.A1(new_n826), .A2(new_n683), .A3(new_n619), .ZN(new_n827));
  INV_X1    g641(.A(new_n827), .ZN(new_n828));
  OAI211_X1 g642(.A(new_n725), .B(new_n618), .C1(new_n647), .C2(new_n661), .ZN(new_n829));
  NAND4_X1  g643(.A1(new_n828), .A2(new_n732), .A3(new_n752), .A4(new_n829), .ZN(new_n830));
  NAND3_X1  g644(.A1(new_n770), .A2(new_n781), .A3(new_n783), .ZN(new_n831));
  NAND2_X1  g645(.A1(new_n307), .A2(new_n312), .ZN(new_n832));
  NAND3_X1  g646(.A1(new_n659), .A2(new_n694), .A3(new_n822), .ZN(new_n833));
  NOR2_X1   g647(.A1(new_n812), .A2(new_n833), .ZN(new_n834));
  NAND4_X1  g648(.A1(new_n690), .A2(new_n832), .A3(new_n834), .A4(new_n759), .ZN(new_n835));
  AND3_X1   g649(.A1(new_n791), .A2(new_n831), .A3(new_n835), .ZN(new_n836));
  NAND2_X1  g650(.A1(new_n789), .A2(new_n836), .ZN(new_n837));
  OAI21_X1  g651(.A(KEYINPUT112), .B1(new_n830), .B2(new_n837), .ZN(new_n838));
  INV_X1    g652(.A(KEYINPUT52), .ZN(new_n839));
  AND2_X1   g653(.A1(new_n768), .A2(new_n771), .ZN(new_n840));
  AND3_X1   g654(.A1(new_n626), .A2(new_n627), .A3(new_n707), .ZN(new_n841));
  NOR2_X1   g655(.A1(new_n693), .A2(new_n191), .ZN(new_n842));
  NAND4_X1  g656(.A1(new_n841), .A2(new_n781), .A3(new_n706), .A4(new_n842), .ZN(new_n843));
  OAI211_X1 g657(.A(new_n313), .B(new_n690), .C1(new_n719), .C2(KEYINPUT105), .ZN(new_n844));
  INV_X1    g658(.A(new_n720), .ZN(new_n845));
  OAI211_X1 g659(.A(new_n696), .B(new_n843), .C1(new_n844), .C2(new_n845), .ZN(new_n846));
  OAI21_X1  g660(.A(new_n839), .B1(new_n840), .B2(new_n846), .ZN(new_n847));
  AND2_X1   g661(.A1(new_n721), .A2(new_n696), .ZN(new_n848));
  AND2_X1   g662(.A1(new_n843), .A2(KEYINPUT52), .ZN(new_n849));
  NAND3_X1  g663(.A1(new_n848), .A2(new_n772), .A3(new_n849), .ZN(new_n850));
  NAND2_X1  g664(.A1(new_n847), .A2(new_n850), .ZN(new_n851));
  NAND3_X1  g665(.A1(new_n829), .A2(new_n732), .A3(new_n752), .ZN(new_n852));
  NOR2_X1   g666(.A1(new_n852), .A2(new_n827), .ZN(new_n853));
  INV_X1    g667(.A(KEYINPUT112), .ZN(new_n854));
  NAND4_X1  g668(.A1(new_n853), .A2(new_n854), .A3(new_n789), .A4(new_n836), .ZN(new_n855));
  INV_X1    g669(.A(KEYINPUT53), .ZN(new_n856));
  NAND4_X1  g670(.A1(new_n838), .A2(new_n851), .A3(new_n855), .A4(new_n856), .ZN(new_n857));
  NOR3_X1   g671(.A1(new_n837), .A2(new_n827), .A3(new_n852), .ZN(new_n858));
  INV_X1    g672(.A(new_n846), .ZN(new_n859));
  AOI21_X1  g673(.A(KEYINPUT52), .B1(new_n859), .B2(new_n772), .ZN(new_n860));
  NOR3_X1   g674(.A1(new_n840), .A2(new_n846), .A3(new_n839), .ZN(new_n861));
  OAI21_X1  g675(.A(new_n858), .B1(new_n860), .B2(new_n861), .ZN(new_n862));
  INV_X1    g676(.A(new_n862), .ZN(new_n863));
  OAI211_X1 g677(.A(new_n857), .B(KEYINPUT54), .C1(new_n863), .C2(new_n856), .ZN(new_n864));
  INV_X1    g678(.A(KEYINPUT51), .ZN(new_n865));
  INV_X1    g679(.A(new_n808), .ZN(new_n866));
  INV_X1    g680(.A(new_n503), .ZN(new_n867));
  NAND3_X1  g681(.A1(new_n866), .A2(new_n750), .A3(new_n867), .ZN(new_n868));
  NOR2_X1   g682(.A1(new_n868), .A2(new_n812), .ZN(new_n869));
  INV_X1    g683(.A(new_n869), .ZN(new_n870));
  NAND2_X1  g684(.A1(new_n758), .A2(new_n307), .ZN(new_n871));
  NAND2_X1  g685(.A1(new_n871), .A2(KEYINPUT114), .ZN(new_n872));
  INV_X1    g686(.A(KEYINPUT114), .ZN(new_n873));
  NAND3_X1  g687(.A1(new_n758), .A2(new_n873), .A3(new_n307), .ZN(new_n874));
  AOI21_X1  g688(.A(new_n759), .B1(new_n872), .B2(new_n874), .ZN(new_n875));
  INV_X1    g689(.A(KEYINPUT115), .ZN(new_n876));
  XNOR2_X1  g690(.A(new_n875), .B(new_n876), .ZN(new_n877));
  AOI21_X1  g691(.A(new_n870), .B1(new_n877), .B2(new_n818), .ZN(new_n878));
  INV_X1    g692(.A(new_n871), .ZN(new_n879));
  NOR2_X1   g693(.A1(new_n782), .A2(new_n503), .ZN(new_n880));
  NAND4_X1  g694(.A1(new_n866), .A2(new_n879), .A3(new_n762), .A4(new_n880), .ZN(new_n881));
  NAND2_X1  g695(.A1(new_n601), .A2(new_n705), .ZN(new_n882));
  NOR2_X1   g696(.A1(new_n882), .A2(new_n545), .ZN(new_n883));
  NOR3_X1   g697(.A1(new_n449), .A2(new_n764), .A3(new_n628), .ZN(new_n884));
  NAND4_X1  g698(.A1(new_n879), .A2(new_n880), .A3(new_n883), .A4(new_n884), .ZN(new_n885));
  NAND2_X1  g699(.A1(new_n881), .A2(new_n885), .ZN(new_n886));
  AND3_X1   g700(.A1(new_n866), .A2(new_n750), .A3(new_n867), .ZN(new_n887));
  INV_X1    g701(.A(new_n378), .ZN(new_n888));
  XNOR2_X1  g702(.A(new_n377), .B(new_n698), .ZN(new_n889));
  NAND3_X1  g703(.A1(new_n725), .A2(new_n888), .A3(new_n889), .ZN(new_n890));
  INV_X1    g704(.A(new_n890), .ZN(new_n891));
  NAND3_X1  g705(.A1(new_n887), .A2(new_n891), .A3(KEYINPUT50), .ZN(new_n892));
  INV_X1    g706(.A(KEYINPUT50), .ZN(new_n893));
  OAI21_X1  g707(.A(new_n893), .B1(new_n868), .B2(new_n890), .ZN(new_n894));
  AOI21_X1  g708(.A(new_n886), .B1(new_n892), .B2(new_n894), .ZN(new_n895));
  INV_X1    g709(.A(new_n895), .ZN(new_n896));
  OAI21_X1  g710(.A(new_n865), .B1(new_n878), .B2(new_n896), .ZN(new_n897));
  NAND2_X1  g711(.A1(new_n872), .A2(new_n874), .ZN(new_n898));
  NAND2_X1  g712(.A1(new_n898), .A2(new_n191), .ZN(new_n899));
  NAND2_X1  g713(.A1(new_n818), .A2(new_n899), .ZN(new_n900));
  NAND2_X1  g714(.A1(new_n900), .A2(new_n869), .ZN(new_n901));
  NAND3_X1  g715(.A1(new_n901), .A2(KEYINPUT51), .A3(new_n895), .ZN(new_n902));
  NAND4_X1  g716(.A1(new_n879), .A2(new_n646), .A3(new_n880), .A4(new_n883), .ZN(new_n903));
  OAI211_X1 g717(.A(new_n903), .B(new_n501), .C1(new_n868), .C2(new_n760), .ZN(new_n904));
  NAND3_X1  g718(.A1(new_n866), .A2(new_n879), .A3(new_n880), .ZN(new_n905));
  INV_X1    g719(.A(new_n618), .ZN(new_n906));
  OR3_X1    g720(.A1(new_n905), .A2(KEYINPUT48), .A3(new_n906), .ZN(new_n907));
  OAI21_X1  g721(.A(KEYINPUT48), .B1(new_n905), .B2(new_n906), .ZN(new_n908));
  AOI21_X1  g722(.A(new_n904), .B1(new_n907), .B2(new_n908), .ZN(new_n909));
  NAND4_X1  g723(.A1(new_n897), .A2(new_n902), .A3(KEYINPUT116), .A4(new_n909), .ZN(new_n910));
  INV_X1    g724(.A(KEYINPUT116), .ZN(new_n911));
  NAND2_X1  g725(.A1(new_n899), .A2(new_n876), .ZN(new_n912));
  INV_X1    g726(.A(KEYINPUT47), .ZN(new_n913));
  OR2_X1    g727(.A1(new_n817), .A2(new_n913), .ZN(new_n914));
  NAND2_X1  g728(.A1(new_n817), .A2(new_n913), .ZN(new_n915));
  NAND2_X1  g729(.A1(new_n875), .A2(KEYINPUT115), .ZN(new_n916));
  NAND4_X1  g730(.A1(new_n912), .A2(new_n914), .A3(new_n915), .A4(new_n916), .ZN(new_n917));
  NAND2_X1  g731(.A1(new_n917), .A2(new_n869), .ZN(new_n918));
  AOI21_X1  g732(.A(KEYINPUT51), .B1(new_n918), .B2(new_n895), .ZN(new_n919));
  AOI21_X1  g733(.A(new_n870), .B1(new_n818), .B2(new_n899), .ZN(new_n920));
  INV_X1    g734(.A(new_n886), .ZN(new_n921));
  AOI21_X1  g735(.A(KEYINPUT50), .B1(new_n887), .B2(new_n891), .ZN(new_n922));
  NOR3_X1   g736(.A1(new_n868), .A2(new_n890), .A3(new_n893), .ZN(new_n923));
  OAI211_X1 g737(.A(KEYINPUT51), .B(new_n921), .C1(new_n922), .C2(new_n923), .ZN(new_n924));
  OAI21_X1  g738(.A(new_n909), .B1(new_n920), .B2(new_n924), .ZN(new_n925));
  OAI21_X1  g739(.A(new_n911), .B1(new_n919), .B2(new_n925), .ZN(new_n926));
  NAND2_X1  g740(.A1(new_n862), .A2(new_n856), .ZN(new_n927));
  INV_X1    g741(.A(KEYINPUT54), .ZN(new_n928));
  INV_X1    g742(.A(KEYINPUT113), .ZN(new_n929));
  XNOR2_X1  g743(.A(new_n852), .B(new_n929), .ZN(new_n930));
  NOR3_X1   g744(.A1(new_n837), .A2(new_n856), .A3(new_n827), .ZN(new_n931));
  NAND3_X1  g745(.A1(new_n851), .A2(new_n930), .A3(new_n931), .ZN(new_n932));
  NAND3_X1  g746(.A1(new_n927), .A2(new_n928), .A3(new_n932), .ZN(new_n933));
  NAND4_X1  g747(.A1(new_n864), .A2(new_n910), .A3(new_n926), .A4(new_n933), .ZN(new_n934));
  NAND2_X1  g748(.A1(new_n500), .A2(new_n288), .ZN(new_n935));
  NAND2_X1  g749(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  OR2_X1    g750(.A1(new_n871), .A2(KEYINPUT49), .ZN(new_n937));
  NAND2_X1  g751(.A1(new_n871), .A2(KEYINPUT49), .ZN(new_n938));
  NAND3_X1  g752(.A1(new_n544), .A2(new_n759), .A3(new_n378), .ZN(new_n939));
  NOR3_X1   g753(.A1(new_n882), .A2(new_n805), .A3(new_n939), .ZN(new_n940));
  NAND4_X1  g754(.A1(new_n937), .A2(new_n889), .A3(new_n938), .A4(new_n940), .ZN(new_n941));
  NAND2_X1  g755(.A1(new_n936), .A2(new_n941), .ZN(new_n942));
  NAND2_X1  g756(.A1(new_n942), .A2(KEYINPUT117), .ZN(new_n943));
  INV_X1    g757(.A(KEYINPUT117), .ZN(new_n944));
  NAND3_X1  g758(.A1(new_n936), .A2(new_n944), .A3(new_n941), .ZN(new_n945));
  NAND2_X1  g759(.A1(new_n943), .A2(new_n945), .ZN(G75));
  AND3_X1   g760(.A1(new_n851), .A2(new_n930), .A3(new_n931), .ZN(new_n947));
  AND2_X1   g761(.A1(new_n843), .A2(new_n696), .ZN(new_n948));
  NAND4_X1  g762(.A1(new_n772), .A2(new_n948), .A3(KEYINPUT52), .A4(new_n721), .ZN(new_n949));
  NAND2_X1  g763(.A1(new_n847), .A2(new_n949), .ZN(new_n950));
  AOI21_X1  g764(.A(KEYINPUT53), .B1(new_n950), .B2(new_n858), .ZN(new_n951));
  NOR2_X1   g765(.A1(new_n947), .A2(new_n951), .ZN(new_n952));
  NOR2_X1   g766(.A1(new_n952), .A2(new_n190), .ZN(new_n953));
  NAND2_X1  g767(.A1(new_n953), .A2(G210), .ZN(new_n954));
  INV_X1    g768(.A(KEYINPUT56), .ZN(new_n955));
  NAND2_X1  g769(.A1(new_n348), .A2(new_n349), .ZN(new_n956));
  XNOR2_X1  g770(.A(new_n956), .B(KEYINPUT118), .ZN(new_n957));
  XNOR2_X1  g771(.A(new_n357), .B(KEYINPUT55), .ZN(new_n958));
  XNOR2_X1  g772(.A(new_n957), .B(new_n958), .ZN(new_n959));
  AND3_X1   g773(.A1(new_n954), .A2(new_n955), .A3(new_n959), .ZN(new_n960));
  AOI21_X1  g774(.A(new_n959), .B1(new_n954), .B2(new_n955), .ZN(new_n961));
  NOR2_X1   g775(.A1(new_n288), .A2(G952), .ZN(new_n962));
  NOR3_X1   g776(.A1(new_n960), .A2(new_n961), .A3(new_n962), .ZN(G51));
  NAND2_X1  g777(.A1(new_n796), .A2(new_n797), .ZN(new_n964));
  XNOR2_X1  g778(.A(new_n964), .B(KEYINPUT120), .ZN(new_n965));
  NOR3_X1   g779(.A1(new_n952), .A2(new_n190), .A3(new_n965), .ZN(new_n966));
  XOR2_X1   g780(.A(new_n779), .B(KEYINPUT57), .Z(new_n967));
  NOR3_X1   g781(.A1(new_n947), .A2(new_n951), .A3(KEYINPUT54), .ZN(new_n968));
  AOI21_X1  g782(.A(new_n928), .B1(new_n927), .B2(new_n932), .ZN(new_n969));
  OAI21_X1  g783(.A(new_n967), .B1(new_n968), .B2(new_n969), .ZN(new_n970));
  NAND2_X1  g784(.A1(new_n970), .A2(new_n305), .ZN(new_n971));
  INV_X1    g785(.A(KEYINPUT119), .ZN(new_n972));
  AOI21_X1  g786(.A(new_n966), .B1(new_n971), .B2(new_n972), .ZN(new_n973));
  NAND3_X1  g787(.A1(new_n970), .A2(KEYINPUT119), .A3(new_n305), .ZN(new_n974));
  AOI21_X1  g788(.A(new_n962), .B1(new_n973), .B2(new_n974), .ZN(G54));
  NAND3_X1  g789(.A1(new_n953), .A2(KEYINPUT58), .A3(G475), .ZN(new_n976));
  NAND3_X1  g790(.A1(new_n976), .A2(new_n424), .A3(new_n439), .ZN(new_n977));
  INV_X1    g791(.A(new_n962), .ZN(new_n978));
  NAND4_X1  g792(.A1(new_n953), .A2(KEYINPUT58), .A3(G475), .A4(new_n440), .ZN(new_n979));
  AND3_X1   g793(.A1(new_n977), .A2(new_n978), .A3(new_n979), .ZN(G60));
  XNOR2_X1  g794(.A(KEYINPUT121), .B(KEYINPUT59), .ZN(new_n981));
  NAND2_X1  g795(.A1(G478), .A2(G902), .ZN(new_n982));
  XNOR2_X1  g796(.A(new_n981), .B(new_n982), .ZN(new_n983));
  AOI21_X1  g797(.A(new_n983), .B1(new_n864), .B2(new_n933), .ZN(new_n984));
  OAI21_X1  g798(.A(new_n978), .B1(new_n984), .B2(new_n638), .ZN(new_n985));
  OR2_X1    g799(.A1(new_n968), .A2(new_n969), .ZN(new_n986));
  AOI21_X1  g800(.A(new_n983), .B1(new_n636), .B2(new_n637), .ZN(new_n987));
  NAND2_X1  g801(.A1(new_n986), .A2(new_n987), .ZN(new_n988));
  INV_X1    g802(.A(KEYINPUT122), .ZN(new_n989));
  NAND2_X1  g803(.A1(new_n988), .A2(new_n989), .ZN(new_n990));
  NAND3_X1  g804(.A1(new_n986), .A2(KEYINPUT122), .A3(new_n987), .ZN(new_n991));
  AOI21_X1  g805(.A(new_n985), .B1(new_n990), .B2(new_n991), .ZN(G63));
  NAND2_X1  g806(.A1(G217), .A2(G902), .ZN(new_n993));
  XOR2_X1   g807(.A(new_n993), .B(KEYINPUT123), .Z(new_n994));
  XNOR2_X1  g808(.A(new_n994), .B(KEYINPUT60), .ZN(new_n995));
  OAI22_X1  g809(.A1(new_n952), .A2(new_n995), .B1(new_n541), .B2(new_n540), .ZN(new_n996));
  OR2_X1    g810(.A1(new_n996), .A2(KEYINPUT125), .ZN(new_n997));
  AOI21_X1  g811(.A(new_n995), .B1(new_n927), .B2(new_n932), .ZN(new_n998));
  NAND2_X1  g812(.A1(new_n998), .A2(new_n674), .ZN(new_n999));
  NAND2_X1  g813(.A1(new_n996), .A2(KEYINPUT125), .ZN(new_n1000));
  INV_X1    g814(.A(KEYINPUT61), .ZN(new_n1001));
  NOR2_X1   g815(.A1(new_n962), .A2(new_n1001), .ZN(new_n1002));
  NAND4_X1  g816(.A1(new_n997), .A2(new_n999), .A3(new_n1000), .A4(new_n1002), .ZN(new_n1003));
  AOI21_X1  g817(.A(KEYINPUT124), .B1(new_n996), .B2(new_n978), .ZN(new_n1004));
  OAI211_X1 g818(.A(KEYINPUT124), .B(new_n978), .C1(new_n998), .C2(new_n542), .ZN(new_n1005));
  NAND2_X1  g819(.A1(new_n1005), .A2(new_n999), .ZN(new_n1006));
  OAI21_X1  g820(.A(new_n1001), .B1(new_n1004), .B2(new_n1006), .ZN(new_n1007));
  NAND2_X1  g821(.A1(new_n1003), .A2(new_n1007), .ZN(G66));
  OAI21_X1  g822(.A(G953), .B1(new_n504), .B2(new_n355), .ZN(new_n1009));
  OAI21_X1  g823(.A(new_n1009), .B1(new_n853), .B2(G953), .ZN(new_n1010));
  OAI21_X1  g824(.A(new_n957), .B1(G898), .B2(new_n288), .ZN(new_n1011));
  XNOR2_X1  g825(.A(new_n1010), .B(new_n1011), .ZN(G69));
  AOI21_X1  g826(.A(new_n288), .B1(G227), .B2(G900), .ZN(new_n1013));
  XOR2_X1   g827(.A(new_n588), .B(new_n435), .Z(new_n1014));
  AND2_X1   g828(.A1(new_n848), .A2(new_n772), .ZN(new_n1015));
  NAND3_X1  g829(.A1(new_n713), .A2(new_n714), .A3(new_n1015), .ZN(new_n1016));
  OR2_X1    g830(.A1(new_n1016), .A2(KEYINPUT62), .ZN(new_n1017));
  NAND2_X1  g831(.A1(new_n1016), .A2(KEYINPUT62), .ZN(new_n1018));
  NOR2_X1   g832(.A1(new_n646), .A2(new_n823), .ZN(new_n1019));
  OR4_X1    g833(.A1(new_n906), .A2(new_n711), .A3(new_n812), .A4(new_n1019), .ZN(new_n1020));
  NAND3_X1  g834(.A1(new_n820), .A2(new_n814), .A3(new_n1020), .ZN(new_n1021));
  INV_X1    g835(.A(new_n1021), .ZN(new_n1022));
  NAND3_X1  g836(.A1(new_n1017), .A2(new_n1018), .A3(new_n1022), .ZN(new_n1023));
  AOI21_X1  g837(.A(new_n1014), .B1(new_n1023), .B2(new_n288), .ZN(new_n1024));
  NAND3_X1  g838(.A1(new_n802), .A2(new_n618), .A3(new_n841), .ZN(new_n1025));
  AND2_X1   g839(.A1(new_n1015), .A2(new_n1025), .ZN(new_n1026));
  AND2_X1   g840(.A1(new_n789), .A2(new_n791), .ZN(new_n1027));
  NAND4_X1  g841(.A1(new_n820), .A2(new_n1026), .A3(new_n814), .A4(new_n1027), .ZN(new_n1028));
  NOR2_X1   g842(.A1(new_n1028), .A2(G953), .ZN(new_n1029));
  NAND2_X1  g843(.A1(G900), .A2(G953), .ZN(new_n1030));
  NAND2_X1  g844(.A1(new_n1014), .A2(new_n1030), .ZN(new_n1031));
  NOR2_X1   g845(.A1(new_n1029), .A2(new_n1031), .ZN(new_n1032));
  OAI21_X1  g846(.A(new_n1013), .B1(new_n1024), .B2(new_n1032), .ZN(new_n1033));
  INV_X1    g847(.A(new_n1032), .ZN(new_n1034));
  INV_X1    g848(.A(new_n1013), .ZN(new_n1035));
  AOI21_X1  g849(.A(new_n1021), .B1(KEYINPUT62), .B2(new_n1016), .ZN(new_n1036));
  AOI21_X1  g850(.A(G953), .B1(new_n1036), .B2(new_n1017), .ZN(new_n1037));
  OAI211_X1 g851(.A(new_n1034), .B(new_n1035), .C1(new_n1037), .C2(new_n1014), .ZN(new_n1038));
  NAND2_X1  g852(.A1(new_n1033), .A2(new_n1038), .ZN(G72));
  NAND3_X1  g853(.A1(new_n1036), .A2(new_n853), .A3(new_n1017), .ZN(new_n1040));
  XNOR2_X1  g854(.A(KEYINPUT126), .B(KEYINPUT63), .ZN(new_n1041));
  NOR2_X1   g855(.A1(new_n621), .A2(new_n190), .ZN(new_n1042));
  XOR2_X1   g856(.A(new_n1041), .B(new_n1042), .Z(new_n1043));
  INV_X1    g857(.A(new_n1043), .ZN(new_n1044));
  AOI21_X1  g858(.A(new_n702), .B1(new_n1040), .B2(new_n1044), .ZN(new_n1045));
  OAI21_X1  g859(.A(new_n1044), .B1(new_n1028), .B2(new_n830), .ZN(new_n1046));
  NAND3_X1  g860(.A1(new_n1046), .A2(new_n580), .A3(new_n589), .ZN(new_n1047));
  AOI21_X1  g861(.A(KEYINPUT127), .B1(new_n589), .B2(new_n565), .ZN(new_n1048));
  NAND2_X1  g862(.A1(new_n612), .A2(new_n580), .ZN(new_n1049));
  XNOR2_X1  g863(.A(new_n1048), .B(new_n1049), .ZN(new_n1050));
  NOR2_X1   g864(.A1(new_n1050), .A2(new_n1043), .ZN(new_n1051));
  OAI211_X1 g865(.A(new_n857), .B(new_n1051), .C1(new_n863), .C2(new_n856), .ZN(new_n1052));
  NAND3_X1  g866(.A1(new_n1047), .A2(new_n978), .A3(new_n1052), .ZN(new_n1053));
  NOR2_X1   g867(.A1(new_n1045), .A2(new_n1053), .ZN(G57));
endmodule


