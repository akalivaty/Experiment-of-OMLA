//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 0 0 1 0 1 0 1 0 1 1 1 1 0 1 0 0 1 1 0 1 1 1 0 1 0 1 0 0 1 0 0 1 1 0 0 1 0 0 0 0 0 1 0 0 0 0 0 0 0 0 0 1 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:17:47 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n677, new_n678, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n699, new_n700, new_n701, new_n702, new_n703,
    new_n704, new_n705, new_n706, new_n707, new_n708, new_n709, new_n710,
    new_n711, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n746, new_n747, new_n748, new_n749,
    new_n750, new_n751, new_n752, new_n754, new_n755, new_n756, new_n757,
    new_n758, new_n759, new_n760, new_n761, new_n762, new_n764, new_n765,
    new_n767, new_n768, new_n769, new_n770, new_n771, new_n772, new_n773,
    new_n774, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n790, new_n791, new_n792, new_n793, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n845, new_n846, new_n848, new_n849,
    new_n851, new_n852, new_n853, new_n854, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n893, new_n894, new_n896,
    new_n897, new_n898, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n908, new_n909, new_n910, new_n912, new_n913,
    new_n914, new_n916, new_n917, new_n918, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n934, new_n935, new_n936, new_n937, new_n938,
    new_n939, new_n941, new_n942, new_n943;
  INV_X1    g000(.A(KEYINPUT28), .ZN(new_n202));
  INV_X1    g001(.A(KEYINPUT68), .ZN(new_n203));
  INV_X1    g002(.A(G183gat), .ZN(new_n204));
  OAI21_X1  g003(.A(new_n203), .B1(new_n204), .B2(KEYINPUT27), .ZN(new_n205));
  INV_X1    g004(.A(KEYINPUT27), .ZN(new_n206));
  OAI21_X1  g005(.A(KEYINPUT67), .B1(new_n206), .B2(G183gat), .ZN(new_n207));
  INV_X1    g006(.A(KEYINPUT67), .ZN(new_n208));
  NAND3_X1  g007(.A1(new_n208), .A2(new_n204), .A3(KEYINPUT27), .ZN(new_n209));
  NAND3_X1  g008(.A1(new_n205), .A2(new_n207), .A3(new_n209), .ZN(new_n210));
  NAND3_X1  g009(.A1(new_n206), .A2(KEYINPUT68), .A3(G183gat), .ZN(new_n211));
  INV_X1    g010(.A(G190gat), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  OAI21_X1  g012(.A(new_n202), .B1(new_n210), .B2(new_n213), .ZN(new_n214));
  XNOR2_X1  g013(.A(KEYINPUT27), .B(G183gat), .ZN(new_n215));
  NAND3_X1  g014(.A1(new_n215), .A2(KEYINPUT28), .A3(new_n212), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n214), .A2(new_n216), .ZN(new_n217));
  INV_X1    g016(.A(G169gat), .ZN(new_n218));
  INV_X1    g017(.A(G176gat), .ZN(new_n219));
  NOR2_X1   g018(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  NOR2_X1   g019(.A1(G169gat), .A2(G176gat), .ZN(new_n221));
  NOR3_X1   g020(.A1(new_n220), .A2(KEYINPUT26), .A3(new_n221), .ZN(new_n222));
  NAND2_X1  g021(.A1(G183gat), .A2(G190gat), .ZN(new_n223));
  INV_X1    g022(.A(new_n221), .ZN(new_n224));
  INV_X1    g023(.A(KEYINPUT26), .ZN(new_n225));
  OAI21_X1  g024(.A(new_n223), .B1(new_n224), .B2(new_n225), .ZN(new_n226));
  NOR2_X1   g025(.A1(new_n222), .A2(new_n226), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n217), .A2(new_n227), .ZN(new_n228));
  INV_X1    g027(.A(KEYINPUT24), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n223), .A2(new_n229), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n204), .A2(new_n212), .ZN(new_n231));
  NAND3_X1  g030(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n232));
  NAND3_X1  g031(.A1(new_n230), .A2(new_n231), .A3(new_n232), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n233), .A2(KEYINPUT64), .ZN(new_n234));
  INV_X1    g033(.A(KEYINPUT23), .ZN(new_n235));
  NOR3_X1   g034(.A1(new_n235), .A2(G169gat), .A3(G176gat), .ZN(new_n236));
  OAI21_X1  g035(.A(KEYINPUT23), .B1(new_n218), .B2(new_n219), .ZN(new_n237));
  AOI21_X1  g036(.A(new_n236), .B1(new_n224), .B2(new_n237), .ZN(new_n238));
  INV_X1    g037(.A(KEYINPUT64), .ZN(new_n239));
  NAND4_X1  g038(.A1(new_n230), .A2(new_n231), .A3(new_n239), .A4(new_n232), .ZN(new_n240));
  NAND3_X1  g039(.A1(new_n234), .A2(new_n238), .A3(new_n240), .ZN(new_n241));
  INV_X1    g040(.A(KEYINPUT25), .ZN(new_n242));
  AND2_X1   g041(.A1(new_n241), .A2(new_n242), .ZN(new_n243));
  INV_X1    g042(.A(KEYINPUT66), .ZN(new_n244));
  NAND3_X1  g043(.A1(new_n204), .A2(new_n212), .A3(KEYINPUT65), .ZN(new_n245));
  INV_X1    g044(.A(KEYINPUT65), .ZN(new_n246));
  OAI21_X1  g045(.A(new_n246), .B1(G183gat), .B2(G190gat), .ZN(new_n247));
  AND4_X1   g046(.A1(new_n230), .A2(new_n245), .A3(new_n247), .A4(new_n232), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n221), .A2(KEYINPUT23), .ZN(new_n249));
  AOI21_X1  g048(.A(new_n235), .B1(G169gat), .B2(G176gat), .ZN(new_n250));
  OAI211_X1 g049(.A(KEYINPUT25), .B(new_n249), .C1(new_n250), .C2(new_n221), .ZN(new_n251));
  OAI21_X1  g050(.A(new_n244), .B1(new_n248), .B2(new_n251), .ZN(new_n252));
  NAND4_X1  g051(.A1(new_n230), .A2(new_n245), .A3(new_n247), .A4(new_n232), .ZN(new_n253));
  NAND4_X1  g052(.A1(new_n238), .A2(KEYINPUT66), .A3(new_n253), .A4(KEYINPUT25), .ZN(new_n254));
  NAND2_X1  g053(.A1(new_n252), .A2(new_n254), .ZN(new_n255));
  OAI21_X1  g054(.A(new_n228), .B1(new_n243), .B2(new_n255), .ZN(new_n256));
  INV_X1    g055(.A(KEYINPUT73), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  INV_X1    g057(.A(G113gat), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n259), .A2(KEYINPUT71), .ZN(new_n260));
  INV_X1    g059(.A(KEYINPUT71), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n261), .A2(G113gat), .ZN(new_n262));
  NAND3_X1  g061(.A1(new_n260), .A2(new_n262), .A3(G120gat), .ZN(new_n263));
  XNOR2_X1  g062(.A(KEYINPUT70), .B(G120gat), .ZN(new_n264));
  OAI21_X1  g063(.A(new_n263), .B1(new_n264), .B2(new_n259), .ZN(new_n265));
  INV_X1    g064(.A(G134gat), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n266), .A2(G127gat), .ZN(new_n267));
  INV_X1    g066(.A(G127gat), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n268), .A2(G134gat), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n267), .A2(new_n269), .ZN(new_n270));
  NOR2_X1   g069(.A1(new_n270), .A2(KEYINPUT1), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n265), .A2(new_n271), .ZN(new_n272));
  INV_X1    g071(.A(KEYINPUT72), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  OR2_X1    g073(.A1(KEYINPUT69), .A2(G120gat), .ZN(new_n275));
  NAND2_X1  g074(.A1(KEYINPUT69), .A2(G120gat), .ZN(new_n276));
  NAND3_X1  g075(.A1(new_n275), .A2(new_n259), .A3(new_n276), .ZN(new_n277));
  INV_X1    g076(.A(KEYINPUT1), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  AOI21_X1  g078(.A(new_n259), .B1(new_n275), .B2(new_n276), .ZN(new_n280));
  OAI21_X1  g079(.A(new_n270), .B1(new_n279), .B2(new_n280), .ZN(new_n281));
  NAND3_X1  g080(.A1(new_n265), .A2(new_n271), .A3(KEYINPUT72), .ZN(new_n282));
  NAND3_X1  g081(.A1(new_n274), .A2(new_n281), .A3(new_n282), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n241), .A2(new_n242), .ZN(new_n284));
  NAND3_X1  g083(.A1(new_n284), .A2(new_n252), .A3(new_n254), .ZN(new_n285));
  NAND3_X1  g084(.A1(new_n285), .A2(KEYINPUT73), .A3(new_n228), .ZN(new_n286));
  NAND3_X1  g085(.A1(new_n258), .A2(new_n283), .A3(new_n286), .ZN(new_n287));
  INV_X1    g086(.A(G227gat), .ZN(new_n288));
  INV_X1    g087(.A(G233gat), .ZN(new_n289));
  NOR2_X1   g088(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  AND3_X1   g089(.A1(new_n265), .A2(KEYINPUT72), .A3(new_n271), .ZN(new_n291));
  AOI21_X1  g090(.A(KEYINPUT72), .B1(new_n265), .B2(new_n271), .ZN(new_n292));
  NOR2_X1   g091(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  NAND4_X1  g092(.A1(new_n256), .A2(new_n257), .A3(new_n281), .A4(new_n293), .ZN(new_n294));
  NAND3_X1  g093(.A1(new_n287), .A2(new_n290), .A3(new_n294), .ZN(new_n295));
  INV_X1    g094(.A(KEYINPUT74), .ZN(new_n296));
  NAND2_X1  g095(.A1(new_n295), .A2(new_n296), .ZN(new_n297));
  NAND4_X1  g096(.A1(new_n287), .A2(KEYINPUT74), .A3(new_n290), .A4(new_n294), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n297), .A2(new_n298), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n299), .A2(KEYINPUT32), .ZN(new_n300));
  INV_X1    g099(.A(KEYINPUT75), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  INV_X1    g101(.A(KEYINPUT32), .ZN(new_n303));
  AOI21_X1  g102(.A(new_n303), .B1(new_n297), .B2(new_n298), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n304), .A2(KEYINPUT75), .ZN(new_n305));
  XNOR2_X1  g104(.A(G15gat), .B(G43gat), .ZN(new_n306));
  XNOR2_X1  g105(.A(G71gat), .B(G99gat), .ZN(new_n307));
  XNOR2_X1  g106(.A(new_n306), .B(new_n307), .ZN(new_n308));
  INV_X1    g107(.A(KEYINPUT33), .ZN(new_n309));
  AOI21_X1  g108(.A(new_n308), .B1(new_n299), .B2(new_n309), .ZN(new_n310));
  NAND3_X1  g109(.A1(new_n302), .A2(new_n305), .A3(new_n310), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n287), .A2(new_n294), .ZN(new_n312));
  OAI21_X1  g111(.A(new_n312), .B1(new_n288), .B2(new_n289), .ZN(new_n313));
  XOR2_X1   g112(.A(new_n313), .B(KEYINPUT34), .Z(new_n314));
  INV_X1    g113(.A(new_n308), .ZN(new_n315));
  AND2_X1   g114(.A1(new_n315), .A2(KEYINPUT76), .ZN(new_n316));
  OAI21_X1  g115(.A(KEYINPUT33), .B1(new_n315), .B2(KEYINPUT76), .ZN(new_n317));
  OAI21_X1  g116(.A(new_n304), .B1(new_n316), .B2(new_n317), .ZN(new_n318));
  AND3_X1   g117(.A1(new_n311), .A2(new_n314), .A3(new_n318), .ZN(new_n319));
  AOI21_X1  g118(.A(new_n314), .B1(new_n311), .B2(new_n318), .ZN(new_n320));
  AOI21_X1  g119(.A(new_n319), .B1(KEYINPUT77), .B2(new_n320), .ZN(new_n321));
  XNOR2_X1  g120(.A(G1gat), .B(G29gat), .ZN(new_n322));
  XNOR2_X1  g121(.A(new_n322), .B(KEYINPUT0), .ZN(new_n323));
  XNOR2_X1  g122(.A(G57gat), .B(G85gat), .ZN(new_n324));
  XOR2_X1   g123(.A(new_n323), .B(new_n324), .Z(new_n325));
  INV_X1    g124(.A(new_n325), .ZN(new_n326));
  INV_X1    g125(.A(KEYINPUT4), .ZN(new_n327));
  INV_X1    g126(.A(KEYINPUT82), .ZN(new_n328));
  NOR3_X1   g127(.A1(new_n328), .A2(G155gat), .A3(G162gat), .ZN(new_n329));
  INV_X1    g128(.A(G155gat), .ZN(new_n330));
  INV_X1    g129(.A(G162gat), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n330), .A2(new_n331), .ZN(new_n332));
  NAND2_X1  g131(.A1(G155gat), .A2(G162gat), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n333), .A2(KEYINPUT82), .ZN(new_n334));
  AOI21_X1  g133(.A(new_n329), .B1(new_n332), .B2(new_n334), .ZN(new_n335));
  OR2_X1    g134(.A1(KEYINPUT83), .A2(KEYINPUT2), .ZN(new_n336));
  INV_X1    g135(.A(G141gat), .ZN(new_n337));
  INV_X1    g136(.A(G148gat), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n337), .A2(new_n338), .ZN(new_n339));
  NAND2_X1  g138(.A1(G141gat), .A2(G148gat), .ZN(new_n340));
  NAND2_X1  g139(.A1(KEYINPUT83), .A2(KEYINPUT2), .ZN(new_n341));
  NAND4_X1  g140(.A1(new_n336), .A2(new_n339), .A3(new_n340), .A4(new_n341), .ZN(new_n342));
  OAI21_X1  g141(.A(new_n333), .B1(new_n332), .B2(KEYINPUT2), .ZN(new_n343));
  AND2_X1   g142(.A1(new_n339), .A2(new_n340), .ZN(new_n344));
  AOI22_X1  g143(.A1(new_n335), .A2(new_n342), .B1(new_n343), .B2(new_n344), .ZN(new_n345));
  NAND4_X1  g144(.A1(new_n293), .A2(new_n327), .A3(new_n281), .A4(new_n345), .ZN(new_n346));
  NAND4_X1  g145(.A1(new_n274), .A2(new_n281), .A3(new_n282), .A4(new_n345), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n347), .A2(KEYINPUT4), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n346), .A2(new_n348), .ZN(new_n349));
  INV_X1    g148(.A(KEYINPUT84), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n283), .A2(new_n350), .ZN(new_n351));
  NAND4_X1  g150(.A1(new_n274), .A2(KEYINPUT84), .A3(new_n281), .A4(new_n282), .ZN(new_n352));
  XNOR2_X1  g151(.A(new_n345), .B(KEYINPUT3), .ZN(new_n353));
  NAND3_X1  g152(.A1(new_n351), .A2(new_n352), .A3(new_n353), .ZN(new_n354));
  NAND2_X1  g153(.A1(G225gat), .A2(G233gat), .ZN(new_n355));
  AND3_X1   g154(.A1(new_n349), .A2(new_n354), .A3(new_n355), .ZN(new_n356));
  INV_X1    g155(.A(new_n345), .ZN(new_n357));
  NAND3_X1  g156(.A1(new_n351), .A2(new_n352), .A3(new_n357), .ZN(new_n358));
  AOI21_X1  g157(.A(new_n355), .B1(new_n358), .B2(new_n347), .ZN(new_n359));
  INV_X1    g158(.A(KEYINPUT5), .ZN(new_n360));
  NOR3_X1   g159(.A1(new_n356), .A2(new_n359), .A3(new_n360), .ZN(new_n361));
  OR3_X1    g160(.A1(new_n347), .A2(KEYINPUT85), .A3(KEYINPUT4), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n346), .A2(KEYINPUT85), .ZN(new_n363));
  NAND3_X1  g162(.A1(new_n362), .A2(new_n363), .A3(new_n348), .ZN(new_n364));
  INV_X1    g163(.A(new_n355), .ZN(new_n365));
  NOR2_X1   g164(.A1(new_n365), .A2(KEYINPUT5), .ZN(new_n366));
  NAND3_X1  g165(.A1(new_n364), .A2(new_n354), .A3(new_n366), .ZN(new_n367));
  INV_X1    g166(.A(new_n367), .ZN(new_n368));
  OAI21_X1  g167(.A(new_n326), .B1(new_n361), .B2(new_n368), .ZN(new_n369));
  INV_X1    g168(.A(KEYINPUT6), .ZN(new_n370));
  NAND3_X1  g169(.A1(new_n349), .A2(new_n354), .A3(new_n355), .ZN(new_n371));
  AND2_X1   g170(.A1(new_n358), .A2(new_n347), .ZN(new_n372));
  OAI211_X1 g171(.A(KEYINPUT5), .B(new_n371), .C1(new_n372), .C2(new_n355), .ZN(new_n373));
  NAND3_X1  g172(.A1(new_n373), .A2(new_n325), .A3(new_n367), .ZN(new_n374));
  NAND3_X1  g173(.A1(new_n369), .A2(new_n370), .A3(new_n374), .ZN(new_n375));
  OAI211_X1 g174(.A(KEYINPUT6), .B(new_n326), .C1(new_n361), .C2(new_n368), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n375), .A2(new_n376), .ZN(new_n377));
  AND2_X1   g176(.A1(G226gat), .A2(G233gat), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n256), .A2(new_n378), .ZN(new_n379));
  AOI21_X1  g178(.A(KEYINPUT29), .B1(new_n285), .B2(new_n228), .ZN(new_n380));
  OAI21_X1  g179(.A(new_n379), .B1(new_n380), .B2(new_n378), .ZN(new_n381));
  XNOR2_X1  g180(.A(G197gat), .B(G204gat), .ZN(new_n382));
  NAND2_X1  g181(.A1(G211gat), .A2(G218gat), .ZN(new_n383));
  OAI21_X1  g182(.A(new_n383), .B1(KEYINPUT79), .B2(KEYINPUT22), .ZN(new_n384));
  AND2_X1   g183(.A1(KEYINPUT79), .A2(KEYINPUT22), .ZN(new_n385));
  OAI21_X1  g184(.A(new_n382), .B1(new_n384), .B2(new_n385), .ZN(new_n386));
  XNOR2_X1  g185(.A(G211gat), .B(G218gat), .ZN(new_n387));
  XNOR2_X1  g186(.A(new_n386), .B(new_n387), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n381), .A2(new_n388), .ZN(new_n389));
  INV_X1    g188(.A(new_n388), .ZN(new_n390));
  OAI211_X1 g189(.A(new_n379), .B(new_n390), .C1(new_n378), .C2(new_n380), .ZN(new_n391));
  XNOR2_X1  g190(.A(G8gat), .B(G36gat), .ZN(new_n392));
  XNOR2_X1  g191(.A(G64gat), .B(G92gat), .ZN(new_n393));
  XOR2_X1   g192(.A(new_n392), .B(new_n393), .Z(new_n394));
  NAND3_X1  g193(.A1(new_n389), .A2(new_n391), .A3(new_n394), .ZN(new_n395));
  INV_X1    g194(.A(KEYINPUT81), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n395), .A2(new_n396), .ZN(new_n397));
  INV_X1    g196(.A(KEYINPUT30), .ZN(new_n398));
  NAND4_X1  g197(.A1(new_n389), .A2(KEYINPUT81), .A3(new_n391), .A4(new_n394), .ZN(new_n399));
  NAND3_X1  g198(.A1(new_n397), .A2(new_n398), .A3(new_n399), .ZN(new_n400));
  XOR2_X1   g199(.A(new_n394), .B(KEYINPUT80), .Z(new_n401));
  AOI21_X1  g200(.A(new_n401), .B1(new_n389), .B2(new_n391), .ZN(new_n402));
  INV_X1    g201(.A(new_n395), .ZN(new_n403));
  AOI21_X1  g202(.A(new_n402), .B1(new_n403), .B2(KEYINPUT30), .ZN(new_n404));
  AND2_X1   g203(.A1(new_n400), .A2(new_n404), .ZN(new_n405));
  AND3_X1   g204(.A1(new_n377), .A2(KEYINPUT86), .A3(new_n405), .ZN(new_n406));
  AOI21_X1  g205(.A(KEYINPUT86), .B1(new_n377), .B2(new_n405), .ZN(new_n407));
  OR2_X1    g206(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  INV_X1    g207(.A(KEYINPUT3), .ZN(new_n409));
  AOI21_X1  g208(.A(KEYINPUT29), .B1(new_n345), .B2(new_n409), .ZN(new_n410));
  NOR2_X1   g209(.A1(new_n390), .A2(new_n410), .ZN(new_n411));
  OAI21_X1  g210(.A(new_n409), .B1(new_n388), .B2(KEYINPUT29), .ZN(new_n412));
  AOI21_X1  g211(.A(new_n411), .B1(new_n357), .B2(new_n412), .ZN(new_n413));
  XNOR2_X1  g212(.A(new_n413), .B(G22gat), .ZN(new_n414));
  NAND2_X1  g213(.A1(G228gat), .A2(G233gat), .ZN(new_n415));
  XNOR2_X1  g214(.A(new_n414), .B(new_n415), .ZN(new_n416));
  INV_X1    g215(.A(new_n416), .ZN(new_n417));
  XNOR2_X1  g216(.A(G78gat), .B(G106gat), .ZN(new_n418));
  XNOR2_X1  g217(.A(KEYINPUT31), .B(G50gat), .ZN(new_n419));
  XOR2_X1   g218(.A(new_n418), .B(new_n419), .Z(new_n420));
  XNOR2_X1  g219(.A(new_n420), .B(KEYINPUT87), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n417), .A2(new_n421), .ZN(new_n422));
  INV_X1    g221(.A(KEYINPUT87), .ZN(new_n423));
  NAND3_X1  g222(.A1(new_n416), .A2(new_n423), .A3(new_n420), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n422), .A2(new_n424), .ZN(new_n425));
  INV_X1    g224(.A(new_n425), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n299), .A2(new_n309), .ZN(new_n427));
  OAI211_X1 g226(.A(new_n427), .B(new_n315), .C1(KEYINPUT75), .C2(new_n304), .ZN(new_n428));
  INV_X1    g227(.A(new_n305), .ZN(new_n429));
  OAI21_X1  g228(.A(new_n318), .B1(new_n428), .B2(new_n429), .ZN(new_n430));
  INV_X1    g229(.A(new_n314), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  INV_X1    g231(.A(KEYINPUT77), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n432), .A2(new_n433), .ZN(new_n434));
  NAND4_X1  g233(.A1(new_n321), .A2(new_n408), .A3(new_n426), .A4(new_n434), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n435), .A2(KEYINPUT35), .ZN(new_n436));
  NAND3_X1  g235(.A1(new_n311), .A2(new_n314), .A3(new_n318), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n432), .A2(new_n437), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n400), .A2(new_n404), .ZN(new_n439));
  NOR3_X1   g238(.A1(new_n438), .A2(new_n425), .A3(new_n439), .ZN(new_n440));
  INV_X1    g239(.A(new_n377), .ZN(new_n441));
  NOR2_X1   g240(.A1(new_n441), .A2(KEYINPUT35), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n440), .A2(new_n442), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n436), .A2(new_n443), .ZN(new_n444));
  NOR2_X1   g243(.A1(new_n406), .A2(new_n407), .ZN(new_n445));
  AOI21_X1  g244(.A(new_n325), .B1(new_n373), .B2(new_n367), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n364), .A2(new_n354), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n447), .A2(new_n365), .ZN(new_n448));
  INV_X1    g247(.A(KEYINPUT39), .ZN(new_n449));
  AOI21_X1  g248(.A(new_n449), .B1(new_n372), .B2(new_n355), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n448), .A2(new_n450), .ZN(new_n451));
  NAND3_X1  g250(.A1(new_n447), .A2(new_n449), .A3(new_n365), .ZN(new_n452));
  NAND3_X1  g251(.A1(new_n451), .A2(new_n325), .A3(new_n452), .ZN(new_n453));
  INV_X1    g252(.A(KEYINPUT40), .ZN(new_n454));
  AOI21_X1  g253(.A(new_n446), .B1(new_n453), .B2(new_n454), .ZN(new_n455));
  NAND4_X1  g254(.A1(new_n451), .A2(KEYINPUT40), .A3(new_n325), .A4(new_n452), .ZN(new_n456));
  NAND3_X1  g255(.A1(new_n455), .A2(new_n439), .A3(new_n456), .ZN(new_n457));
  INV_X1    g256(.A(KEYINPUT88), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  NAND4_X1  g258(.A1(new_n455), .A2(new_n439), .A3(KEYINPUT88), .A4(new_n456), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  INV_X1    g260(.A(KEYINPUT37), .ZN(new_n462));
  NAND3_X1  g261(.A1(new_n389), .A2(new_n462), .A3(new_n391), .ZN(new_n463));
  INV_X1    g262(.A(new_n394), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  AOI21_X1  g264(.A(new_n462), .B1(new_n389), .B2(new_n391), .ZN(new_n466));
  OAI21_X1  g265(.A(KEYINPUT38), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  NOR2_X1   g266(.A1(new_n401), .A2(KEYINPUT38), .ZN(new_n468));
  AND3_X1   g267(.A1(new_n389), .A2(KEYINPUT89), .A3(new_n391), .ZN(new_n469));
  OAI21_X1  g268(.A(KEYINPUT37), .B1(new_n389), .B2(KEYINPUT89), .ZN(new_n470));
  OAI211_X1 g269(.A(new_n463), .B(new_n468), .C1(new_n469), .C2(new_n470), .ZN(new_n471));
  AND4_X1   g270(.A1(new_n397), .A2(new_n467), .A3(new_n399), .A4(new_n471), .ZN(new_n472));
  AOI21_X1  g271(.A(new_n425), .B1(new_n441), .B2(new_n472), .ZN(new_n473));
  AOI22_X1  g272(.A1(new_n425), .A2(new_n445), .B1(new_n461), .B2(new_n473), .ZN(new_n474));
  INV_X1    g273(.A(KEYINPUT36), .ZN(new_n475));
  NAND3_X1  g274(.A1(new_n430), .A2(KEYINPUT77), .A3(new_n431), .ZN(new_n476));
  NAND3_X1  g275(.A1(new_n434), .A2(new_n476), .A3(new_n437), .ZN(new_n477));
  OAI21_X1  g276(.A(KEYINPUT78), .B1(new_n319), .B2(new_n320), .ZN(new_n478));
  AOI21_X1  g277(.A(new_n475), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  AOI211_X1 g278(.A(KEYINPUT78), .B(KEYINPUT36), .C1(new_n432), .C2(new_n437), .ZN(new_n480));
  OAI21_X1  g279(.A(new_n474), .B1(new_n479), .B2(new_n480), .ZN(new_n481));
  NAND2_X1  g280(.A1(new_n444), .A2(new_n481), .ZN(new_n482));
  XNOR2_X1  g281(.A(G15gat), .B(G22gat), .ZN(new_n483));
  OR3_X1    g282(.A1(new_n483), .A2(KEYINPUT95), .A3(G1gat), .ZN(new_n484));
  OAI21_X1  g283(.A(KEYINPUT95), .B1(new_n483), .B2(G1gat), .ZN(new_n485));
  AND2_X1   g284(.A1(KEYINPUT93), .A2(G1gat), .ZN(new_n486));
  OAI21_X1  g285(.A(KEYINPUT16), .B1(KEYINPUT93), .B2(G1gat), .ZN(new_n487));
  OAI21_X1  g286(.A(new_n483), .B1(new_n486), .B2(new_n487), .ZN(new_n488));
  INV_X1    g287(.A(KEYINPUT94), .ZN(new_n489));
  OAI211_X1 g288(.A(new_n484), .B(new_n485), .C1(new_n488), .C2(new_n489), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n490), .A2(G8gat), .ZN(new_n491));
  NAND2_X1  g290(.A1(KEYINPUT94), .A2(G8gat), .ZN(new_n492));
  AND2_X1   g291(.A1(new_n488), .A2(new_n492), .ZN(new_n493));
  OR3_X1    g292(.A1(new_n483), .A2(G1gat), .A3(G8gat), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n491), .A2(new_n495), .ZN(new_n496));
  XNOR2_X1  g295(.A(G57gat), .B(G64gat), .ZN(new_n497));
  INV_X1    g296(.A(new_n497), .ZN(new_n498));
  OR2_X1    g297(.A1(G71gat), .A2(G78gat), .ZN(new_n499));
  NAND2_X1  g298(.A1(G71gat), .A2(G78gat), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  INV_X1    g300(.A(KEYINPUT9), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n500), .A2(new_n502), .ZN(new_n503));
  NAND3_X1  g302(.A1(new_n498), .A2(new_n501), .A3(new_n503), .ZN(new_n504));
  OAI211_X1 g303(.A(new_n500), .B(new_n499), .C1(new_n497), .C2(new_n502), .ZN(new_n505));
  AND2_X1   g304(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  NAND2_X1  g305(.A1(new_n506), .A2(KEYINPUT97), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n504), .A2(new_n505), .ZN(new_n508));
  INV_X1    g307(.A(KEYINPUT97), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  AND2_X1   g309(.A1(new_n507), .A2(new_n510), .ZN(new_n511));
  AOI21_X1  g310(.A(new_n496), .B1(new_n511), .B2(KEYINPUT21), .ZN(new_n512));
  XNOR2_X1  g311(.A(new_n512), .B(KEYINPUT98), .ZN(new_n513));
  XNOR2_X1  g312(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n514));
  XNOR2_X1  g313(.A(new_n514), .B(new_n330), .ZN(new_n515));
  XNOR2_X1  g314(.A(new_n513), .B(new_n515), .ZN(new_n516));
  NOR2_X1   g315(.A1(new_n506), .A2(KEYINPUT21), .ZN(new_n517));
  NAND2_X1  g316(.A1(G231gat), .A2(G233gat), .ZN(new_n518));
  XNOR2_X1  g317(.A(new_n517), .B(new_n518), .ZN(new_n519));
  XNOR2_X1  g318(.A(new_n519), .B(new_n268), .ZN(new_n520));
  XOR2_X1   g319(.A(G183gat), .B(G211gat), .Z(new_n521));
  XNOR2_X1  g320(.A(new_n520), .B(new_n521), .ZN(new_n522));
  XNOR2_X1  g321(.A(new_n516), .B(new_n522), .ZN(new_n523));
  XNOR2_X1  g322(.A(G134gat), .B(G162gat), .ZN(new_n524));
  INV_X1    g323(.A(KEYINPUT99), .ZN(new_n525));
  INV_X1    g324(.A(G85gat), .ZN(new_n526));
  INV_X1    g325(.A(G92gat), .ZN(new_n527));
  OAI21_X1  g326(.A(new_n525), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  NAND3_X1  g327(.A1(KEYINPUT99), .A2(G85gat), .A3(G92gat), .ZN(new_n529));
  NAND3_X1  g328(.A1(new_n528), .A2(KEYINPUT7), .A3(new_n529), .ZN(new_n530));
  INV_X1    g329(.A(KEYINPUT7), .ZN(new_n531));
  OAI211_X1 g330(.A(new_n525), .B(new_n531), .C1(new_n526), .C2(new_n527), .ZN(new_n532));
  NAND2_X1  g331(.A1(G99gat), .A2(G106gat), .ZN(new_n533));
  AOI22_X1  g332(.A1(KEYINPUT8), .A2(new_n533), .B1(new_n526), .B2(new_n527), .ZN(new_n534));
  NAND3_X1  g333(.A1(new_n530), .A2(new_n532), .A3(new_n534), .ZN(new_n535));
  XOR2_X1   g334(.A(G99gat), .B(G106gat), .Z(new_n536));
  NAND2_X1  g335(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  INV_X1    g336(.A(new_n536), .ZN(new_n538));
  NAND4_X1  g337(.A1(new_n538), .A2(new_n530), .A3(new_n532), .A4(new_n534), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n537), .A2(new_n539), .ZN(new_n540));
  INV_X1    g339(.A(KEYINPUT100), .ZN(new_n541));
  XNOR2_X1  g340(.A(new_n540), .B(new_n541), .ZN(new_n542));
  INV_X1    g341(.A(KEYINPUT17), .ZN(new_n543));
  INV_X1    g342(.A(G29gat), .ZN(new_n544));
  INV_X1    g343(.A(G36gat), .ZN(new_n545));
  NAND3_X1  g344(.A1(new_n544), .A2(new_n545), .A3(KEYINPUT14), .ZN(new_n546));
  INV_X1    g345(.A(KEYINPUT14), .ZN(new_n547));
  OAI21_X1  g346(.A(new_n547), .B1(G29gat), .B2(G36gat), .ZN(new_n548));
  NAND2_X1  g347(.A1(new_n546), .A2(new_n548), .ZN(new_n549));
  INV_X1    g348(.A(KEYINPUT91), .ZN(new_n550));
  AOI22_X1  g349(.A1(new_n549), .A2(new_n550), .B1(G29gat), .B2(G36gat), .ZN(new_n551));
  NAND3_X1  g350(.A1(new_n546), .A2(new_n548), .A3(KEYINPUT91), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  INV_X1    g352(.A(G43gat), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n554), .A2(G50gat), .ZN(new_n555));
  INV_X1    g354(.A(G50gat), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n556), .A2(G43gat), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n555), .A2(new_n557), .ZN(new_n558));
  OR2_X1    g357(.A1(new_n558), .A2(KEYINPUT90), .ZN(new_n559));
  INV_X1    g358(.A(KEYINPUT15), .ZN(new_n560));
  AOI21_X1  g359(.A(new_n560), .B1(new_n558), .B2(KEYINPUT90), .ZN(new_n561));
  NAND3_X1  g360(.A1(new_n553), .A2(new_n559), .A3(new_n561), .ZN(new_n562));
  NAND2_X1  g361(.A1(new_n559), .A2(new_n561), .ZN(new_n563));
  OR2_X1    g362(.A1(KEYINPUT92), .A2(G43gat), .ZN(new_n564));
  NAND2_X1  g363(.A1(KEYINPUT92), .A2(G43gat), .ZN(new_n565));
  AOI21_X1  g364(.A(G50gat), .B1(new_n564), .B2(new_n565), .ZN(new_n566));
  INV_X1    g365(.A(new_n555), .ZN(new_n567));
  OAI21_X1  g366(.A(new_n560), .B1(new_n566), .B2(new_n567), .ZN(new_n568));
  AOI21_X1  g367(.A(new_n549), .B1(G29gat), .B2(G36gat), .ZN(new_n569));
  NAND3_X1  g368(.A1(new_n563), .A2(new_n568), .A3(new_n569), .ZN(new_n570));
  AOI21_X1  g369(.A(new_n543), .B1(new_n562), .B2(new_n570), .ZN(new_n571));
  AND3_X1   g370(.A1(new_n562), .A2(new_n570), .A3(new_n543), .ZN(new_n572));
  OAI21_X1  g371(.A(new_n542), .B1(new_n571), .B2(new_n572), .ZN(new_n573));
  INV_X1    g372(.A(KEYINPUT101), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n562), .A2(new_n570), .ZN(new_n575));
  AND2_X1   g374(.A1(new_n537), .A2(new_n539), .ZN(new_n576));
  AND2_X1   g375(.A1(G232gat), .A2(G233gat), .ZN(new_n577));
  AOI22_X1  g376(.A1(new_n575), .A2(new_n576), .B1(KEYINPUT41), .B2(new_n577), .ZN(new_n578));
  NAND3_X1  g377(.A1(new_n573), .A2(new_n574), .A3(new_n578), .ZN(new_n579));
  INV_X1    g378(.A(new_n579), .ZN(new_n580));
  AOI21_X1  g379(.A(new_n574), .B1(new_n573), .B2(new_n578), .ZN(new_n581));
  OAI21_X1  g380(.A(new_n524), .B1(new_n580), .B2(new_n581), .ZN(new_n582));
  NAND2_X1  g381(.A1(new_n573), .A2(new_n578), .ZN(new_n583));
  NAND2_X1  g382(.A1(new_n583), .A2(KEYINPUT101), .ZN(new_n584));
  INV_X1    g383(.A(new_n524), .ZN(new_n585));
  NAND3_X1  g384(.A1(new_n584), .A2(new_n579), .A3(new_n585), .ZN(new_n586));
  NOR2_X1   g385(.A1(new_n577), .A2(KEYINPUT41), .ZN(new_n587));
  XNOR2_X1  g386(.A(G190gat), .B(G218gat), .ZN(new_n588));
  XNOR2_X1  g387(.A(new_n587), .B(new_n588), .ZN(new_n589));
  AND3_X1   g388(.A1(new_n582), .A2(new_n586), .A3(new_n589), .ZN(new_n590));
  AOI21_X1  g389(.A(new_n589), .B1(new_n582), .B2(new_n586), .ZN(new_n591));
  NOR2_X1   g390(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  XNOR2_X1  g391(.A(G120gat), .B(G148gat), .ZN(new_n593));
  XNOR2_X1  g392(.A(G176gat), .B(G204gat), .ZN(new_n594));
  XOR2_X1   g393(.A(new_n593), .B(new_n594), .Z(new_n595));
  INV_X1    g394(.A(new_n595), .ZN(new_n596));
  NAND2_X1  g395(.A1(new_n536), .A2(KEYINPUT102), .ZN(new_n597));
  NAND3_X1  g396(.A1(new_n504), .A2(new_n505), .A3(new_n597), .ZN(new_n598));
  NAND2_X1  g397(.A1(new_n540), .A2(new_n598), .ZN(new_n599));
  NAND4_X1  g398(.A1(new_n506), .A2(new_n537), .A3(new_n539), .A4(new_n597), .ZN(new_n600));
  INV_X1    g399(.A(KEYINPUT10), .ZN(new_n601));
  NAND3_X1  g400(.A1(new_n599), .A2(new_n600), .A3(new_n601), .ZN(new_n602));
  NAND4_X1  g401(.A1(new_n576), .A2(new_n507), .A3(KEYINPUT10), .A4(new_n510), .ZN(new_n603));
  AND2_X1   g402(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  NAND2_X1  g403(.A1(G230gat), .A2(G233gat), .ZN(new_n605));
  INV_X1    g404(.A(new_n605), .ZN(new_n606));
  NOR2_X1   g405(.A1(new_n604), .A2(new_n606), .ZN(new_n607));
  AOI21_X1  g406(.A(new_n605), .B1(new_n599), .B2(new_n600), .ZN(new_n608));
  OAI21_X1  g407(.A(new_n596), .B1(new_n607), .B2(new_n608), .ZN(new_n609));
  NAND2_X1  g408(.A1(new_n602), .A2(new_n603), .ZN(new_n610));
  NAND2_X1  g409(.A1(new_n610), .A2(KEYINPUT103), .ZN(new_n611));
  INV_X1    g410(.A(KEYINPUT103), .ZN(new_n612));
  NAND3_X1  g411(.A1(new_n602), .A2(new_n603), .A3(new_n612), .ZN(new_n613));
  NAND3_X1  g412(.A1(new_n611), .A2(new_n605), .A3(new_n613), .ZN(new_n614));
  INV_X1    g413(.A(new_n614), .ZN(new_n615));
  AOI21_X1  g414(.A(new_n596), .B1(new_n608), .B2(KEYINPUT104), .ZN(new_n616));
  OAI21_X1  g415(.A(new_n616), .B1(KEYINPUT104), .B2(new_n608), .ZN(new_n617));
  OAI21_X1  g416(.A(new_n609), .B1(new_n615), .B2(new_n617), .ZN(new_n618));
  INV_X1    g417(.A(new_n618), .ZN(new_n619));
  NAND3_X1  g418(.A1(new_n523), .A2(new_n592), .A3(new_n619), .ZN(new_n620));
  INV_X1    g419(.A(KEYINPUT96), .ZN(new_n621));
  AOI22_X1  g420(.A1(new_n490), .A2(G8gat), .B1(new_n493), .B2(new_n494), .ZN(new_n622));
  OAI211_X1 g421(.A(new_n621), .B(new_n622), .C1(new_n572), .C2(new_n571), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n575), .A2(KEYINPUT17), .ZN(new_n624));
  NAND3_X1  g423(.A1(new_n562), .A2(new_n570), .A3(new_n543), .ZN(new_n625));
  AOI21_X1  g424(.A(new_n496), .B1(new_n624), .B2(new_n625), .ZN(new_n626));
  INV_X1    g425(.A(new_n575), .ZN(new_n627));
  OAI21_X1  g426(.A(KEYINPUT96), .B1(new_n627), .B2(new_n622), .ZN(new_n628));
  OAI21_X1  g427(.A(new_n623), .B1(new_n626), .B2(new_n628), .ZN(new_n629));
  NAND2_X1  g428(.A1(G229gat), .A2(G233gat), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  INV_X1    g430(.A(KEYINPUT18), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  XNOR2_X1  g432(.A(G113gat), .B(G141gat), .ZN(new_n634));
  XNOR2_X1  g433(.A(new_n634), .B(G197gat), .ZN(new_n635));
  XOR2_X1   g434(.A(KEYINPUT11), .B(G169gat), .Z(new_n636));
  XNOR2_X1  g435(.A(new_n635), .B(new_n636), .ZN(new_n637));
  XNOR2_X1  g436(.A(new_n637), .B(KEYINPUT12), .ZN(new_n638));
  NAND3_X1  g437(.A1(new_n629), .A2(KEYINPUT18), .A3(new_n630), .ZN(new_n639));
  XNOR2_X1  g438(.A(new_n622), .B(new_n575), .ZN(new_n640));
  XOR2_X1   g439(.A(new_n630), .B(KEYINPUT13), .Z(new_n641));
  INV_X1    g440(.A(new_n641), .ZN(new_n642));
  NOR2_X1   g441(.A1(new_n640), .A2(new_n642), .ZN(new_n643));
  INV_X1    g442(.A(new_n643), .ZN(new_n644));
  NAND4_X1  g443(.A1(new_n633), .A2(new_n638), .A3(new_n639), .A4(new_n644), .ZN(new_n645));
  INV_X1    g444(.A(new_n645), .ZN(new_n646));
  OAI21_X1  g445(.A(new_n622), .B1(new_n572), .B2(new_n571), .ZN(new_n647));
  AOI21_X1  g446(.A(new_n621), .B1(new_n496), .B2(new_n575), .ZN(new_n648));
  NAND2_X1  g447(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  AOI22_X1  g448(.A1(new_n649), .A2(new_n623), .B1(G229gat), .B2(G233gat), .ZN(new_n650));
  AOI21_X1  g449(.A(new_n643), .B1(new_n650), .B2(KEYINPUT18), .ZN(new_n651));
  AOI21_X1  g450(.A(new_n638), .B1(new_n651), .B2(new_n633), .ZN(new_n652));
  NOR2_X1   g451(.A1(new_n646), .A2(new_n652), .ZN(new_n653));
  NOR2_X1   g452(.A1(new_n620), .A2(new_n653), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n482), .A2(new_n654), .ZN(new_n655));
  NOR2_X1   g454(.A1(new_n655), .A2(new_n377), .ZN(new_n656));
  XOR2_X1   g455(.A(new_n656), .B(G1gat), .Z(G1324gat));
  NOR2_X1   g456(.A1(new_n655), .A2(new_n405), .ZN(new_n658));
  XNOR2_X1  g457(.A(KEYINPUT16), .B(G8gat), .ZN(new_n659));
  XOR2_X1   g458(.A(new_n659), .B(KEYINPUT106), .Z(new_n660));
  INV_X1    g459(.A(new_n660), .ZN(new_n661));
  NAND3_X1  g460(.A1(new_n658), .A2(KEYINPUT42), .A3(new_n661), .ZN(new_n662));
  INV_X1    g461(.A(KEYINPUT42), .ZN(new_n663));
  INV_X1    g462(.A(KEYINPUT105), .ZN(new_n664));
  XNOR2_X1  g463(.A(new_n658), .B(new_n664), .ZN(new_n665));
  AOI21_X1  g464(.A(new_n663), .B1(new_n665), .B2(G8gat), .ZN(new_n666));
  NOR2_X1   g465(.A1(new_n665), .A2(new_n660), .ZN(new_n667));
  OAI21_X1  g466(.A(new_n662), .B1(new_n666), .B2(new_n667), .ZN(G1325gat));
  NAND2_X1  g467(.A1(new_n476), .A2(new_n437), .ZN(new_n669));
  NOR2_X1   g468(.A1(new_n320), .A2(KEYINPUT77), .ZN(new_n670));
  OAI21_X1  g469(.A(new_n478), .B1(new_n669), .B2(new_n670), .ZN(new_n671));
  AOI21_X1  g470(.A(new_n480), .B1(new_n671), .B2(KEYINPUT36), .ZN(new_n672));
  INV_X1    g471(.A(new_n672), .ZN(new_n673));
  OAI21_X1  g472(.A(G15gat), .B1(new_n655), .B2(new_n673), .ZN(new_n674));
  OR2_X1    g473(.A1(new_n438), .A2(G15gat), .ZN(new_n675));
  OAI21_X1  g474(.A(new_n674), .B1(new_n655), .B2(new_n675), .ZN(G1326gat));
  NOR2_X1   g475(.A1(new_n655), .A2(new_n426), .ZN(new_n677));
  XOR2_X1   g476(.A(KEYINPUT43), .B(G22gat), .Z(new_n678));
  XNOR2_X1  g477(.A(new_n677), .B(new_n678), .ZN(G1327gat));
  INV_X1    g478(.A(new_n592), .ZN(new_n680));
  NOR3_X1   g479(.A1(new_n523), .A2(new_n653), .A3(new_n618), .ZN(new_n681));
  NAND3_X1  g480(.A1(new_n482), .A2(new_n680), .A3(new_n681), .ZN(new_n682));
  NAND2_X1  g481(.A1(new_n441), .A2(new_n544), .ZN(new_n683));
  OR3_X1    g482(.A1(new_n682), .A2(KEYINPUT45), .A3(new_n683), .ZN(new_n684));
  OAI21_X1  g483(.A(KEYINPUT45), .B1(new_n682), .B2(new_n683), .ZN(new_n685));
  NAND2_X1  g484(.A1(new_n461), .A2(new_n473), .ZN(new_n686));
  OAI21_X1  g485(.A(new_n686), .B1(new_n426), .B2(new_n408), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n671), .A2(KEYINPUT36), .ZN(new_n688));
  INV_X1    g487(.A(new_n480), .ZN(new_n689));
  AOI21_X1  g488(.A(new_n687), .B1(new_n688), .B2(new_n689), .ZN(new_n690));
  AOI22_X1  g489(.A1(new_n435), .A2(KEYINPUT35), .B1(new_n440), .B2(new_n442), .ZN(new_n691));
  OAI21_X1  g490(.A(new_n680), .B1(new_n690), .B2(new_n691), .ZN(new_n692));
  INV_X1    g491(.A(KEYINPUT44), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  OAI211_X1 g493(.A(KEYINPUT44), .B(new_n680), .C1(new_n690), .C2(new_n691), .ZN(new_n695));
  NAND4_X1  g494(.A1(new_n694), .A2(new_n441), .A3(new_n681), .A4(new_n695), .ZN(new_n696));
  AOI22_X1  g495(.A1(new_n684), .A2(new_n685), .B1(G29gat), .B2(new_n696), .ZN(new_n697));
  XNOR2_X1  g496(.A(new_n697), .B(KEYINPUT107), .ZN(G1328gat));
  NOR4_X1   g497(.A1(new_n682), .A2(KEYINPUT46), .A3(G36gat), .A4(new_n405), .ZN(new_n699));
  INV_X1    g498(.A(KEYINPUT46), .ZN(new_n700));
  INV_X1    g499(.A(new_n681), .ZN(new_n701));
  NOR2_X1   g500(.A1(new_n692), .A2(new_n701), .ZN(new_n702));
  NOR2_X1   g501(.A1(new_n405), .A2(G36gat), .ZN(new_n703));
  AOI21_X1  g502(.A(new_n700), .B1(new_n702), .B2(new_n703), .ZN(new_n704));
  NOR2_X1   g503(.A1(new_n699), .A2(new_n704), .ZN(new_n705));
  NAND3_X1  g504(.A1(new_n694), .A2(new_n681), .A3(new_n695), .ZN(new_n706));
  OAI21_X1  g505(.A(G36gat), .B1(new_n706), .B2(new_n405), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n705), .A2(new_n707), .ZN(new_n708));
  NAND2_X1  g507(.A1(new_n708), .A2(KEYINPUT108), .ZN(new_n709));
  INV_X1    g508(.A(KEYINPUT108), .ZN(new_n710));
  NAND3_X1  g509(.A1(new_n705), .A2(new_n710), .A3(new_n707), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n709), .A2(new_n711), .ZN(G1329gat));
  NAND2_X1  g511(.A1(new_n564), .A2(new_n565), .ZN(new_n713));
  NOR2_X1   g512(.A1(new_n438), .A2(new_n713), .ZN(new_n714));
  INV_X1    g513(.A(new_n714), .ZN(new_n715));
  NOR2_X1   g514(.A1(new_n682), .A2(new_n715), .ZN(new_n716));
  INV_X1    g515(.A(KEYINPUT47), .ZN(new_n717));
  NOR2_X1   g516(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  NAND4_X1  g517(.A1(new_n694), .A2(new_n672), .A3(new_n681), .A4(new_n695), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n719), .A2(KEYINPUT110), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n720), .A2(new_n713), .ZN(new_n721));
  NOR2_X1   g520(.A1(new_n719), .A2(KEYINPUT110), .ZN(new_n722));
  OAI21_X1  g521(.A(new_n718), .B1(new_n721), .B2(new_n722), .ZN(new_n723));
  NAND2_X1  g522(.A1(new_n719), .A2(new_n713), .ZN(new_n724));
  INV_X1    g523(.A(new_n716), .ZN(new_n725));
  NAND2_X1  g524(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  AOI21_X1  g525(.A(KEYINPUT109), .B1(new_n726), .B2(new_n717), .ZN(new_n727));
  AOI21_X1  g526(.A(new_n716), .B1(new_n719), .B2(new_n713), .ZN(new_n728));
  INV_X1    g527(.A(KEYINPUT109), .ZN(new_n729));
  NOR3_X1   g528(.A1(new_n728), .A2(new_n729), .A3(KEYINPUT47), .ZN(new_n730));
  OAI21_X1  g529(.A(new_n723), .B1(new_n727), .B2(new_n730), .ZN(G1330gat));
  OAI21_X1  g530(.A(G50gat), .B1(new_n706), .B2(new_n426), .ZN(new_n732));
  NOR2_X1   g531(.A1(new_n426), .A2(G50gat), .ZN(new_n733));
  INV_X1    g532(.A(KEYINPUT48), .ZN(new_n734));
  AOI22_X1  g533(.A1(new_n702), .A2(new_n733), .B1(KEYINPUT111), .B2(new_n734), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n732), .A2(new_n735), .ZN(new_n736));
  OR2_X1    g535(.A1(new_n734), .A2(KEYINPUT111), .ZN(new_n737));
  XNOR2_X1  g536(.A(new_n736), .B(new_n737), .ZN(G1331gat));
  INV_X1    g537(.A(new_n523), .ZN(new_n739));
  INV_X1    g538(.A(new_n653), .ZN(new_n740));
  NOR3_X1   g539(.A1(new_n739), .A2(new_n740), .A3(new_n680), .ZN(new_n741));
  NAND3_X1  g540(.A1(new_n482), .A2(new_n618), .A3(new_n741), .ZN(new_n742));
  INV_X1    g541(.A(new_n742), .ZN(new_n743));
  NAND2_X1  g542(.A1(new_n743), .A2(new_n441), .ZN(new_n744));
  XNOR2_X1  g543(.A(new_n744), .B(G57gat), .ZN(G1332gat));
  AND2_X1   g544(.A1(new_n482), .A2(new_n741), .ZN(new_n746));
  NOR2_X1   g545(.A1(new_n405), .A2(new_n619), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  OAI21_X1  g547(.A(new_n748), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n749));
  XOR2_X1   g548(.A(KEYINPUT49), .B(G64gat), .Z(new_n750));
  OAI21_X1  g549(.A(new_n749), .B1(new_n748), .B2(new_n750), .ZN(new_n751));
  INV_X1    g550(.A(KEYINPUT112), .ZN(new_n752));
  XNOR2_X1  g551(.A(new_n751), .B(new_n752), .ZN(G1333gat));
  OR3_X1    g552(.A1(new_n742), .A2(KEYINPUT113), .A3(new_n438), .ZN(new_n754));
  INV_X1    g553(.A(G71gat), .ZN(new_n755));
  OAI21_X1  g554(.A(KEYINPUT113), .B1(new_n742), .B2(new_n438), .ZN(new_n756));
  NAND3_X1  g555(.A1(new_n754), .A2(new_n755), .A3(new_n756), .ZN(new_n757));
  NAND3_X1  g556(.A1(new_n743), .A2(G71gat), .A3(new_n672), .ZN(new_n758));
  NAND2_X1  g557(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n759), .A2(KEYINPUT50), .ZN(new_n760));
  INV_X1    g559(.A(KEYINPUT50), .ZN(new_n761));
  NAND3_X1  g560(.A1(new_n757), .A2(new_n761), .A3(new_n758), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n760), .A2(new_n762), .ZN(G1334gat));
  NOR2_X1   g562(.A1(new_n742), .A2(new_n426), .ZN(new_n764));
  XOR2_X1   g563(.A(KEYINPUT114), .B(G78gat), .Z(new_n765));
  XNOR2_X1  g564(.A(new_n764), .B(new_n765), .ZN(G1335gat));
  NOR2_X1   g565(.A1(new_n740), .A2(new_n523), .ZN(new_n767));
  OAI211_X1 g566(.A(new_n680), .B(new_n767), .C1(new_n690), .C2(new_n691), .ZN(new_n768));
  INV_X1    g567(.A(KEYINPUT51), .ZN(new_n769));
  XNOR2_X1  g568(.A(new_n768), .B(new_n769), .ZN(new_n770));
  NAND4_X1  g569(.A1(new_n770), .A2(new_n526), .A3(new_n441), .A4(new_n618), .ZN(new_n771));
  NOR3_X1   g570(.A1(new_n740), .A2(new_n523), .A3(new_n619), .ZN(new_n772));
  NAND3_X1  g571(.A1(new_n694), .A2(new_n695), .A3(new_n772), .ZN(new_n773));
  OAI21_X1  g572(.A(G85gat), .B1(new_n773), .B2(new_n377), .ZN(new_n774));
  NAND2_X1  g573(.A1(new_n771), .A2(new_n774), .ZN(G1336gat));
  AND2_X1   g574(.A1(new_n768), .A2(new_n769), .ZN(new_n776));
  NOR2_X1   g575(.A1(new_n768), .A2(new_n769), .ZN(new_n777));
  OAI21_X1  g576(.A(new_n747), .B1(new_n776), .B2(new_n777), .ZN(new_n778));
  NAND2_X1  g577(.A1(new_n778), .A2(new_n527), .ZN(new_n779));
  INV_X1    g578(.A(KEYINPUT52), .ZN(new_n780));
  NOR2_X1   g579(.A1(new_n780), .A2(KEYINPUT115), .ZN(new_n781));
  INV_X1    g580(.A(new_n781), .ZN(new_n782));
  NOR2_X1   g581(.A1(new_n405), .A2(new_n527), .ZN(new_n783));
  NAND4_X1  g582(.A1(new_n694), .A2(new_n695), .A3(new_n772), .A4(new_n783), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n780), .A2(KEYINPUT115), .ZN(new_n785));
  AND2_X1   g584(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  AND3_X1   g585(.A1(new_n779), .A2(new_n782), .A3(new_n786), .ZN(new_n787));
  AOI21_X1  g586(.A(new_n782), .B1(new_n779), .B2(new_n786), .ZN(new_n788));
  NOR2_X1   g587(.A1(new_n787), .A2(new_n788), .ZN(G1337gat));
  NOR3_X1   g588(.A1(new_n438), .A2(G99gat), .A3(new_n619), .ZN(new_n790));
  XOR2_X1   g589(.A(new_n790), .B(KEYINPUT116), .Z(new_n791));
  NAND2_X1  g590(.A1(new_n770), .A2(new_n791), .ZN(new_n792));
  OAI21_X1  g591(.A(G99gat), .B1(new_n773), .B2(new_n673), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n792), .A2(new_n793), .ZN(G1338gat));
  NOR2_X1   g593(.A1(new_n426), .A2(G106gat), .ZN(new_n795));
  NAND3_X1  g594(.A1(new_n770), .A2(new_n618), .A3(new_n795), .ZN(new_n796));
  OAI21_X1  g595(.A(G106gat), .B1(new_n773), .B2(new_n426), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n798), .A2(KEYINPUT53), .ZN(new_n799));
  INV_X1    g598(.A(KEYINPUT53), .ZN(new_n800));
  NAND3_X1  g599(.A1(new_n796), .A2(new_n800), .A3(new_n797), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n799), .A2(new_n801), .ZN(G1339gat));
  OR2_X1    g601(.A1(new_n620), .A2(new_n740), .ZN(new_n803));
  NAND2_X1  g602(.A1(new_n640), .A2(new_n642), .ZN(new_n804));
  OAI21_X1  g603(.A(new_n804), .B1(new_n629), .B2(new_n630), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n805), .A2(new_n637), .ZN(new_n806));
  OAI211_X1 g605(.A(new_n645), .B(new_n806), .C1(new_n590), .C2(new_n591), .ZN(new_n807));
  INV_X1    g606(.A(KEYINPUT54), .ZN(new_n808));
  AOI21_X1  g607(.A(new_n808), .B1(new_n604), .B2(new_n606), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n614), .A2(new_n809), .ZN(new_n810));
  NAND3_X1  g609(.A1(new_n610), .A2(new_n808), .A3(new_n605), .ZN(new_n811));
  INV_X1    g610(.A(KEYINPUT117), .ZN(new_n812));
  AND3_X1   g611(.A1(new_n811), .A2(new_n812), .A3(new_n596), .ZN(new_n813));
  AOI21_X1  g612(.A(new_n812), .B1(new_n811), .B2(new_n596), .ZN(new_n814));
  OAI21_X1  g613(.A(new_n810), .B1(new_n813), .B2(new_n814), .ZN(new_n815));
  INV_X1    g614(.A(KEYINPUT55), .ZN(new_n816));
  OAI21_X1  g615(.A(KEYINPUT118), .B1(new_n815), .B2(new_n816), .ZN(new_n817));
  NOR2_X1   g616(.A1(new_n615), .A2(new_n617), .ZN(new_n818));
  AOI21_X1  g617(.A(new_n818), .B1(new_n815), .B2(new_n816), .ZN(new_n819));
  INV_X1    g618(.A(new_n814), .ZN(new_n820));
  NAND3_X1  g619(.A1(new_n811), .A2(new_n812), .A3(new_n596), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  INV_X1    g621(.A(KEYINPUT118), .ZN(new_n823));
  NAND4_X1  g622(.A1(new_n822), .A2(new_n823), .A3(KEYINPUT55), .A4(new_n810), .ZN(new_n824));
  NAND3_X1  g623(.A1(new_n817), .A2(new_n819), .A3(new_n824), .ZN(new_n825));
  NOR2_X1   g624(.A1(new_n807), .A2(new_n825), .ZN(new_n826));
  NAND3_X1  g625(.A1(new_n645), .A2(new_n618), .A3(new_n806), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n827), .A2(KEYINPUT119), .ZN(new_n828));
  INV_X1    g627(.A(KEYINPUT119), .ZN(new_n829));
  NAND4_X1  g628(.A1(new_n645), .A2(new_n829), .A3(new_n618), .A4(new_n806), .ZN(new_n830));
  OAI211_X1 g629(.A(new_n828), .B(new_n830), .C1(new_n825), .C2(new_n653), .ZN(new_n831));
  AOI21_X1  g630(.A(new_n826), .B1(new_n831), .B2(new_n592), .ZN(new_n832));
  INV_X1    g631(.A(KEYINPUT120), .ZN(new_n833));
  OAI21_X1  g632(.A(new_n739), .B1(new_n832), .B2(new_n833), .ZN(new_n834));
  AOI211_X1 g633(.A(KEYINPUT120), .B(new_n826), .C1(new_n592), .C2(new_n831), .ZN(new_n835));
  OAI21_X1  g634(.A(new_n803), .B1(new_n834), .B2(new_n835), .ZN(new_n836));
  AND2_X1   g635(.A1(new_n836), .A2(new_n441), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n837), .A2(new_n440), .ZN(new_n838));
  OAI21_X1  g637(.A(G113gat), .B1(new_n838), .B2(new_n653), .ZN(new_n839));
  NOR2_X1   g638(.A1(new_n477), .A2(new_n425), .ZN(new_n840));
  AND2_X1   g639(.A1(new_n837), .A2(new_n840), .ZN(new_n841));
  NAND2_X1  g640(.A1(new_n841), .A2(new_n405), .ZN(new_n842));
  NAND3_X1  g641(.A1(new_n740), .A2(new_n260), .A3(new_n262), .ZN(new_n843));
  OAI21_X1  g642(.A(new_n839), .B1(new_n842), .B2(new_n843), .ZN(G1340gat));
  OAI21_X1  g643(.A(G120gat), .B1(new_n838), .B2(new_n619), .ZN(new_n845));
  OR2_X1    g644(.A1(new_n619), .A2(new_n264), .ZN(new_n846));
  OAI21_X1  g645(.A(new_n845), .B1(new_n842), .B2(new_n846), .ZN(G1341gat));
  OAI21_X1  g646(.A(G127gat), .B1(new_n838), .B2(new_n739), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n523), .A2(new_n268), .ZN(new_n849));
  OAI21_X1  g648(.A(new_n848), .B1(new_n842), .B2(new_n849), .ZN(G1342gat));
  NOR2_X1   g649(.A1(new_n592), .A2(new_n439), .ZN(new_n851));
  NAND3_X1  g650(.A1(new_n841), .A2(new_n266), .A3(new_n851), .ZN(new_n852));
  XOR2_X1   g651(.A(new_n852), .B(KEYINPUT56), .Z(new_n853));
  OAI21_X1  g652(.A(G134gat), .B1(new_n838), .B2(new_n592), .ZN(new_n854));
  NAND2_X1  g653(.A1(new_n853), .A2(new_n854), .ZN(G1343gat));
  NOR3_X1   g654(.A1(new_n672), .A2(new_n377), .A3(new_n439), .ZN(new_n856));
  INV_X1    g655(.A(KEYINPUT57), .ZN(new_n857));
  NAND3_X1  g656(.A1(new_n836), .A2(new_n857), .A3(new_n425), .ZN(new_n858));
  OAI21_X1  g657(.A(new_n827), .B1(new_n825), .B2(new_n653), .ZN(new_n859));
  AOI21_X1  g658(.A(new_n826), .B1(new_n592), .B2(new_n859), .ZN(new_n860));
  OAI21_X1  g659(.A(new_n803), .B1(new_n860), .B2(new_n523), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n861), .A2(new_n425), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n862), .A2(KEYINPUT57), .ZN(new_n863));
  NAND3_X1  g662(.A1(new_n856), .A2(new_n858), .A3(new_n863), .ZN(new_n864));
  OAI21_X1  g663(.A(G141gat), .B1(new_n864), .B2(new_n653), .ZN(new_n865));
  AOI21_X1  g664(.A(KEYINPUT58), .B1(new_n865), .B2(KEYINPUT121), .ZN(new_n866));
  AND2_X1   g665(.A1(new_n836), .A2(new_n425), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n867), .A2(new_n856), .ZN(new_n868));
  NAND2_X1  g667(.A1(new_n740), .A2(new_n337), .ZN(new_n869));
  OAI21_X1  g668(.A(new_n865), .B1(new_n868), .B2(new_n869), .ZN(new_n870));
  XOR2_X1   g669(.A(new_n866), .B(new_n870), .Z(G1344gat));
  INV_X1    g670(.A(KEYINPUT123), .ZN(new_n872));
  INV_X1    g671(.A(KEYINPUT59), .ZN(new_n873));
  NAND3_X1  g672(.A1(new_n836), .A2(KEYINPUT57), .A3(new_n425), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n862), .A2(new_n857), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  NAND3_X1  g675(.A1(new_n876), .A2(new_n618), .A3(new_n856), .ZN(new_n877));
  AOI21_X1  g676(.A(new_n873), .B1(new_n877), .B2(G148gat), .ZN(new_n878));
  NAND4_X1  g677(.A1(new_n856), .A2(new_n858), .A3(new_n618), .A4(new_n863), .ZN(new_n879));
  INV_X1    g678(.A(KEYINPUT122), .ZN(new_n880));
  NOR2_X1   g679(.A1(new_n338), .A2(KEYINPUT59), .ZN(new_n881));
  NAND3_X1  g680(.A1(new_n879), .A2(new_n880), .A3(new_n881), .ZN(new_n882));
  INV_X1    g681(.A(new_n882), .ZN(new_n883));
  AOI21_X1  g682(.A(new_n880), .B1(new_n879), .B2(new_n881), .ZN(new_n884));
  NOR3_X1   g683(.A1(new_n878), .A2(new_n883), .A3(new_n884), .ZN(new_n885));
  NOR3_X1   g684(.A1(new_n868), .A2(G148gat), .A3(new_n619), .ZN(new_n886));
  OAI21_X1  g685(.A(new_n872), .B1(new_n885), .B2(new_n886), .ZN(new_n887));
  INV_X1    g686(.A(new_n886), .ZN(new_n888));
  INV_X1    g687(.A(new_n884), .ZN(new_n889));
  NAND2_X1  g688(.A1(new_n889), .A2(new_n882), .ZN(new_n890));
  OAI211_X1 g689(.A(KEYINPUT123), .B(new_n888), .C1(new_n890), .C2(new_n878), .ZN(new_n891));
  NAND2_X1  g690(.A1(new_n887), .A2(new_n891), .ZN(G1345gat));
  OAI21_X1  g691(.A(G155gat), .B1(new_n864), .B2(new_n739), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n523), .A2(new_n330), .ZN(new_n894));
  OAI21_X1  g693(.A(new_n893), .B1(new_n868), .B2(new_n894), .ZN(G1346gat));
  OAI21_X1  g694(.A(G162gat), .B1(new_n864), .B2(new_n592), .ZN(new_n896));
  NAND2_X1  g695(.A1(new_n673), .A2(new_n441), .ZN(new_n897));
  NAND3_X1  g696(.A1(new_n867), .A2(new_n331), .A3(new_n851), .ZN(new_n898));
  OAI21_X1  g697(.A(new_n896), .B1(new_n897), .B2(new_n898), .ZN(G1347gat));
  AND3_X1   g698(.A1(new_n836), .A2(new_n377), .A3(new_n439), .ZN(new_n900));
  AND2_X1   g699(.A1(new_n900), .A2(new_n840), .ZN(new_n901));
  NAND3_X1  g700(.A1(new_n901), .A2(new_n218), .A3(new_n740), .ZN(new_n902));
  NOR2_X1   g701(.A1(new_n438), .A2(new_n425), .ZN(new_n903));
  NAND2_X1  g702(.A1(new_n900), .A2(new_n903), .ZN(new_n904));
  OAI21_X1  g703(.A(G169gat), .B1(new_n904), .B2(new_n653), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n902), .A2(new_n905), .ZN(new_n906));
  XNOR2_X1  g705(.A(new_n906), .B(KEYINPUT124), .ZN(G1348gat));
  NOR3_X1   g706(.A1(new_n904), .A2(new_n219), .A3(new_n619), .ZN(new_n908));
  XNOR2_X1  g707(.A(new_n908), .B(KEYINPUT125), .ZN(new_n909));
  AOI21_X1  g708(.A(G176gat), .B1(new_n901), .B2(new_n618), .ZN(new_n910));
  NOR2_X1   g709(.A1(new_n909), .A2(new_n910), .ZN(G1349gat));
  NAND3_X1  g710(.A1(new_n901), .A2(new_n215), .A3(new_n523), .ZN(new_n912));
  OAI21_X1  g711(.A(G183gat), .B1(new_n904), .B2(new_n739), .ZN(new_n913));
  NAND2_X1  g712(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  XNOR2_X1  g713(.A(new_n914), .B(KEYINPUT60), .ZN(G1350gat));
  OAI21_X1  g714(.A(G190gat), .B1(new_n904), .B2(new_n592), .ZN(new_n916));
  XNOR2_X1  g715(.A(new_n916), .B(KEYINPUT61), .ZN(new_n917));
  NAND3_X1  g716(.A1(new_n901), .A2(new_n212), .A3(new_n680), .ZN(new_n918));
  NAND2_X1  g717(.A1(new_n917), .A2(new_n918), .ZN(G1351gat));
  NOR3_X1   g718(.A1(new_n672), .A2(new_n441), .A3(new_n405), .ZN(new_n920));
  NAND2_X1  g719(.A1(new_n867), .A2(new_n920), .ZN(new_n921));
  INV_X1    g720(.A(new_n921), .ZN(new_n922));
  AOI21_X1  g721(.A(G197gat), .B1(new_n922), .B2(new_n740), .ZN(new_n923));
  AND2_X1   g722(.A1(new_n876), .A2(new_n920), .ZN(new_n924));
  AND2_X1   g723(.A1(new_n740), .A2(G197gat), .ZN(new_n925));
  AOI21_X1  g724(.A(new_n923), .B1(new_n924), .B2(new_n925), .ZN(G1352gat));
  OR2_X1    g725(.A1(new_n619), .A2(G204gat), .ZN(new_n927));
  NOR3_X1   g726(.A1(new_n921), .A2(KEYINPUT62), .A3(new_n927), .ZN(new_n928));
  XOR2_X1   g727(.A(new_n928), .B(KEYINPUT126), .Z(new_n929));
  NAND3_X1  g728(.A1(new_n876), .A2(new_n618), .A3(new_n920), .ZN(new_n930));
  NAND2_X1  g729(.A1(new_n930), .A2(G204gat), .ZN(new_n931));
  OAI21_X1  g730(.A(KEYINPUT62), .B1(new_n921), .B2(new_n927), .ZN(new_n932));
  NAND3_X1  g731(.A1(new_n929), .A2(new_n931), .A3(new_n932), .ZN(G1353gat));
  NAND2_X1  g732(.A1(new_n924), .A2(new_n523), .ZN(new_n934));
  NAND2_X1  g733(.A1(new_n934), .A2(G211gat), .ZN(new_n935));
  OR2_X1    g734(.A1(new_n935), .A2(KEYINPUT63), .ZN(new_n936));
  NAND2_X1  g735(.A1(new_n935), .A2(KEYINPUT63), .ZN(new_n937));
  NOR3_X1   g736(.A1(new_n921), .A2(G211gat), .A3(new_n739), .ZN(new_n938));
  XNOR2_X1  g737(.A(new_n938), .B(KEYINPUT127), .ZN(new_n939));
  NAND3_X1  g738(.A1(new_n936), .A2(new_n937), .A3(new_n939), .ZN(G1354gat));
  INV_X1    g739(.A(G218gat), .ZN(new_n941));
  NAND3_X1  g740(.A1(new_n922), .A2(new_n941), .A3(new_n680), .ZN(new_n942));
  AND2_X1   g741(.A1(new_n924), .A2(new_n680), .ZN(new_n943));
  OAI21_X1  g742(.A(new_n942), .B1(new_n943), .B2(new_n941), .ZN(G1355gat));
endmodule


