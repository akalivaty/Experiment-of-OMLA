//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 1 0 0 0 0 1 1 0 0 1 0 1 0 1 1 1 0 1 1 1 0 0 0 0 0 0 1 0 0 0 1 0 0 0 0 1 0 0 1 0 0 0 0 1 0 0 0 1 0 0 0 0 1 1 0 1 1 1 0 1 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:22:57 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n735, new_n736, new_n737, new_n738,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n752, new_n754, new_n755,
    new_n756, new_n758, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n768, new_n769, new_n770, new_n771,
    new_n772, new_n773, new_n774, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n789, new_n790, new_n791, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n812, new_n813, new_n814, new_n815, new_n816, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n945,
    new_n946, new_n947, new_n948, new_n949, new_n950, new_n951, new_n952,
    new_n953, new_n954, new_n955, new_n956, new_n957, new_n958, new_n959,
    new_n960, new_n961, new_n962, new_n963, new_n964, new_n965, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n995, new_n996, new_n997, new_n998,
    new_n999, new_n1000, new_n1001, new_n1002, new_n1003, new_n1004,
    new_n1005, new_n1007, new_n1008, new_n1009, new_n1010, new_n1011,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1022, new_n1023, new_n1024,
    new_n1025, new_n1026, new_n1027, new_n1028, new_n1029, new_n1030,
    new_n1031, new_n1032, new_n1033, new_n1034, new_n1035, new_n1036,
    new_n1037, new_n1038, new_n1039, new_n1041, new_n1042, new_n1043,
    new_n1044, new_n1045, new_n1046, new_n1047, new_n1048, new_n1049,
    new_n1050, new_n1051, new_n1052, new_n1053, new_n1054, new_n1055,
    new_n1056, new_n1057;
  INV_X1    g000(.A(G217), .ZN(new_n187));
  XNOR2_X1  g001(.A(KEYINPUT69), .B(G902), .ZN(new_n188));
  AOI21_X1  g002(.A(new_n187), .B1(new_n188), .B2(G234), .ZN(new_n189));
  INV_X1    g003(.A(new_n189), .ZN(new_n190));
  XNOR2_X1  g004(.A(KEYINPUT22), .B(G137), .ZN(new_n191));
  INV_X1    g005(.A(G953), .ZN(new_n192));
  NAND3_X1  g006(.A1(new_n192), .A2(G221), .A3(G234), .ZN(new_n193));
  XNOR2_X1  g007(.A(new_n191), .B(new_n193), .ZN(new_n194));
  INV_X1    g008(.A(G140), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n195), .A2(G125), .ZN(new_n196));
  INV_X1    g010(.A(G125), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n197), .A2(G140), .ZN(new_n198));
  NAND3_X1  g012(.A1(new_n196), .A2(new_n198), .A3(KEYINPUT16), .ZN(new_n199));
  OR3_X1    g013(.A1(new_n197), .A2(KEYINPUT16), .A3(G140), .ZN(new_n200));
  NAND3_X1  g014(.A1(new_n199), .A2(new_n200), .A3(G146), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n201), .A2(KEYINPUT70), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n199), .A2(new_n200), .ZN(new_n203));
  INV_X1    g017(.A(G146), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  INV_X1    g019(.A(KEYINPUT70), .ZN(new_n206));
  NAND4_X1  g020(.A1(new_n199), .A2(new_n200), .A3(new_n206), .A4(G146), .ZN(new_n207));
  NAND3_X1  g021(.A1(new_n202), .A2(new_n205), .A3(new_n207), .ZN(new_n208));
  INV_X1    g022(.A(KEYINPUT23), .ZN(new_n209));
  INV_X1    g023(.A(G119), .ZN(new_n210));
  OAI21_X1  g024(.A(new_n209), .B1(new_n210), .B2(G128), .ZN(new_n211));
  INV_X1    g025(.A(G128), .ZN(new_n212));
  NAND3_X1  g026(.A1(new_n212), .A2(KEYINPUT23), .A3(G119), .ZN(new_n213));
  OAI211_X1 g027(.A(new_n211), .B(new_n213), .C1(G119), .C2(new_n212), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n214), .A2(G110), .ZN(new_n215));
  XOR2_X1   g029(.A(KEYINPUT24), .B(G110), .Z(new_n216));
  XNOR2_X1  g030(.A(G119), .B(G128), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  AND2_X1   g032(.A1(new_n215), .A2(new_n218), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n208), .A2(new_n219), .ZN(new_n220));
  XNOR2_X1  g034(.A(G125), .B(G140), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n221), .A2(new_n204), .ZN(new_n222));
  AND2_X1   g036(.A1(new_n201), .A2(new_n222), .ZN(new_n223));
  OAI22_X1  g037(.A1(new_n214), .A2(G110), .B1(new_n217), .B2(new_n216), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  AND3_X1   g039(.A1(new_n220), .A2(KEYINPUT71), .A3(new_n225), .ZN(new_n226));
  AOI21_X1  g040(.A(KEYINPUT71), .B1(new_n220), .B2(new_n225), .ZN(new_n227));
  OAI21_X1  g041(.A(new_n194), .B1(new_n226), .B2(new_n227), .ZN(new_n228));
  AOI22_X1  g042(.A1(new_n208), .A2(new_n219), .B1(new_n224), .B2(new_n223), .ZN(new_n229));
  AOI21_X1  g043(.A(new_n194), .B1(new_n229), .B2(KEYINPUT71), .ZN(new_n230));
  INV_X1    g044(.A(new_n230), .ZN(new_n231));
  NAND3_X1  g045(.A1(new_n228), .A2(new_n188), .A3(new_n231), .ZN(new_n232));
  INV_X1    g046(.A(KEYINPUT25), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n232), .A2(new_n233), .ZN(new_n234));
  NAND4_X1  g048(.A1(new_n228), .A2(KEYINPUT25), .A3(new_n188), .A4(new_n231), .ZN(new_n235));
  AOI21_X1  g049(.A(new_n190), .B1(new_n234), .B2(new_n235), .ZN(new_n236));
  INV_X1    g050(.A(KEYINPUT71), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n215), .A2(new_n218), .ZN(new_n238));
  AOI21_X1  g052(.A(G146), .B1(new_n199), .B2(new_n200), .ZN(new_n239));
  AND3_X1   g053(.A1(new_n199), .A2(G146), .A3(new_n200), .ZN(new_n240));
  AOI21_X1  g054(.A(new_n239), .B1(new_n240), .B2(new_n206), .ZN(new_n241));
  AOI21_X1  g055(.A(new_n238), .B1(new_n241), .B2(new_n202), .ZN(new_n242));
  INV_X1    g056(.A(new_n225), .ZN(new_n243));
  OAI21_X1  g057(.A(new_n237), .B1(new_n242), .B2(new_n243), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n229), .A2(KEYINPUT71), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n244), .A2(new_n245), .ZN(new_n246));
  AOI21_X1  g060(.A(new_n230), .B1(new_n246), .B2(new_n194), .ZN(new_n247));
  NOR2_X1   g061(.A1(new_n189), .A2(G902), .ZN(new_n248));
  AND2_X1   g062(.A1(new_n247), .A2(new_n248), .ZN(new_n249));
  OR2_X1    g063(.A1(new_n236), .A2(new_n249), .ZN(new_n250));
  INV_X1    g064(.A(KEYINPUT31), .ZN(new_n251));
  INV_X1    g065(.A(G116), .ZN(new_n252));
  NOR2_X1   g066(.A1(new_n252), .A2(G119), .ZN(new_n253));
  INV_X1    g067(.A(KEYINPUT67), .ZN(new_n254));
  OAI21_X1  g068(.A(new_n254), .B1(new_n210), .B2(G116), .ZN(new_n255));
  NAND3_X1  g069(.A1(new_n252), .A2(KEYINPUT67), .A3(G119), .ZN(new_n256));
  AOI21_X1  g070(.A(new_n253), .B1(new_n255), .B2(new_n256), .ZN(new_n257));
  XOR2_X1   g071(.A(KEYINPUT2), .B(G113), .Z(new_n258));
  AND2_X1   g072(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  NOR2_X1   g073(.A1(new_n257), .A2(new_n258), .ZN(new_n260));
  NOR2_X1   g074(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  INV_X1    g075(.A(new_n261), .ZN(new_n262));
  INV_X1    g076(.A(G134), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n263), .A2(KEYINPUT65), .ZN(new_n264));
  INV_X1    g078(.A(KEYINPUT65), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n265), .A2(G134), .ZN(new_n266));
  AOI21_X1  g080(.A(G137), .B1(new_n264), .B2(new_n266), .ZN(new_n267));
  INV_X1    g081(.A(G137), .ZN(new_n268));
  NOR2_X1   g082(.A1(new_n268), .A2(G134), .ZN(new_n269));
  OAI21_X1  g083(.A(G131), .B1(new_n267), .B2(new_n269), .ZN(new_n270));
  INV_X1    g084(.A(KEYINPUT66), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  OAI211_X1 g086(.A(KEYINPUT66), .B(G131), .C1(new_n267), .C2(new_n269), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n204), .A2(G143), .ZN(new_n275));
  INV_X1    g089(.A(G143), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n276), .A2(G146), .ZN(new_n277));
  OAI211_X1 g091(.A(new_n275), .B(new_n277), .C1(KEYINPUT1), .C2(new_n212), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n275), .A2(new_n277), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n275), .A2(KEYINPUT1), .ZN(new_n280));
  NAND3_X1  g094(.A1(new_n279), .A2(new_n280), .A3(G128), .ZN(new_n281));
  INV_X1    g095(.A(KEYINPUT11), .ZN(new_n282));
  AOI21_X1  g096(.A(new_n282), .B1(G134), .B2(new_n268), .ZN(new_n283));
  AOI21_X1  g097(.A(new_n283), .B1(new_n267), .B2(new_n282), .ZN(new_n284));
  INV_X1    g098(.A(G131), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n264), .A2(new_n266), .ZN(new_n286));
  OAI21_X1  g100(.A(new_n285), .B1(new_n286), .B2(new_n268), .ZN(new_n287));
  OAI211_X1 g101(.A(new_n278), .B(new_n281), .C1(new_n284), .C2(new_n287), .ZN(new_n288));
  OAI21_X1  g102(.A(KEYINPUT30), .B1(new_n274), .B2(new_n288), .ZN(new_n289));
  NAND2_X1  g103(.A1(KEYINPUT0), .A2(G128), .ZN(new_n290));
  OR2_X1    g104(.A1(KEYINPUT0), .A2(G128), .ZN(new_n291));
  NAND3_X1  g105(.A1(new_n279), .A2(new_n290), .A3(new_n291), .ZN(new_n292));
  NAND4_X1  g106(.A1(new_n275), .A2(new_n277), .A3(KEYINPUT0), .A4(G128), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  AND3_X1   g108(.A1(new_n264), .A2(new_n266), .A3(G137), .ZN(new_n295));
  OAI21_X1  g109(.A(G131), .B1(new_n284), .B2(new_n295), .ZN(new_n296));
  NOR2_X1   g110(.A1(new_n265), .A2(G134), .ZN(new_n297));
  NOR2_X1   g111(.A1(new_n263), .A2(KEYINPUT65), .ZN(new_n298));
  OAI211_X1 g112(.A(new_n282), .B(new_n268), .C1(new_n297), .C2(new_n298), .ZN(new_n299));
  INV_X1    g113(.A(new_n283), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n299), .A2(new_n300), .ZN(new_n301));
  INV_X1    g115(.A(new_n295), .ZN(new_n302));
  NAND3_X1  g116(.A1(new_n301), .A2(new_n285), .A3(new_n302), .ZN(new_n303));
  AOI21_X1  g117(.A(new_n294), .B1(new_n296), .B2(new_n303), .ZN(new_n304));
  OAI21_X1  g118(.A(new_n262), .B1(new_n289), .B2(new_n304), .ZN(new_n305));
  XOR2_X1   g119(.A(KEYINPUT64), .B(KEYINPUT30), .Z(new_n306));
  INV_X1    g120(.A(new_n294), .ZN(new_n307));
  AOI21_X1  g121(.A(new_n285), .B1(new_n301), .B2(new_n302), .ZN(new_n308));
  NOR2_X1   g122(.A1(new_n284), .A2(new_n287), .ZN(new_n309));
  OAI21_X1  g123(.A(new_n307), .B1(new_n308), .B2(new_n309), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n281), .A2(new_n278), .ZN(new_n311));
  INV_X1    g125(.A(new_n311), .ZN(new_n312));
  NAND4_X1  g126(.A1(new_n303), .A2(new_n272), .A3(new_n312), .A4(new_n273), .ZN(new_n313));
  AOI21_X1  g127(.A(new_n306), .B1(new_n310), .B2(new_n313), .ZN(new_n314));
  NOR2_X1   g128(.A1(new_n305), .A2(new_n314), .ZN(new_n315));
  NAND3_X1  g129(.A1(new_n310), .A2(new_n261), .A3(new_n313), .ZN(new_n316));
  NOR2_X1   g130(.A1(G237), .A2(G953), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n317), .A2(G210), .ZN(new_n318));
  XNOR2_X1  g132(.A(new_n318), .B(KEYINPUT27), .ZN(new_n319));
  XNOR2_X1  g133(.A(KEYINPUT26), .B(G101), .ZN(new_n320));
  XNOR2_X1  g134(.A(new_n319), .B(new_n320), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n316), .A2(new_n321), .ZN(new_n322));
  OAI21_X1  g136(.A(new_n251), .B1(new_n315), .B2(new_n322), .ZN(new_n323));
  NAND3_X1  g137(.A1(new_n310), .A2(KEYINPUT30), .A3(new_n313), .ZN(new_n324));
  INV_X1    g138(.A(new_n274), .ZN(new_n325));
  INV_X1    g139(.A(new_n288), .ZN(new_n326));
  AOI21_X1  g140(.A(new_n295), .B1(new_n299), .B2(new_n300), .ZN(new_n327));
  OAI22_X1  g141(.A1(new_n327), .A2(new_n285), .B1(new_n284), .B2(new_n287), .ZN(new_n328));
  AOI22_X1  g142(.A1(new_n325), .A2(new_n326), .B1(new_n328), .B2(new_n307), .ZN(new_n329));
  OAI211_X1 g143(.A(new_n324), .B(new_n262), .C1(new_n329), .C2(new_n306), .ZN(new_n330));
  INV_X1    g144(.A(new_n321), .ZN(new_n331));
  AOI21_X1  g145(.A(new_n331), .B1(new_n329), .B2(new_n261), .ZN(new_n332));
  NAND3_X1  g146(.A1(new_n330), .A2(new_n332), .A3(KEYINPUT31), .ZN(new_n333));
  XOR2_X1   g147(.A(KEYINPUT68), .B(KEYINPUT28), .Z(new_n334));
  AND3_X1   g148(.A1(new_n310), .A2(new_n261), .A3(new_n313), .ZN(new_n335));
  AOI21_X1  g149(.A(new_n261), .B1(new_n310), .B2(new_n313), .ZN(new_n336));
  OAI21_X1  g150(.A(new_n334), .B1(new_n335), .B2(new_n336), .ZN(new_n337));
  INV_X1    g151(.A(KEYINPUT28), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n316), .A2(new_n338), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n337), .A2(new_n339), .ZN(new_n340));
  AOI22_X1  g154(.A1(new_n323), .A2(new_n333), .B1(new_n340), .B2(new_n331), .ZN(new_n341));
  NOR2_X1   g155(.A1(G472), .A2(G902), .ZN(new_n342));
  INV_X1    g156(.A(new_n342), .ZN(new_n343));
  OAI21_X1  g157(.A(KEYINPUT32), .B1(new_n341), .B2(new_n343), .ZN(new_n344));
  INV_X1    g158(.A(new_n334), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n310), .A2(new_n313), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n346), .A2(new_n262), .ZN(new_n347));
  AOI21_X1  g161(.A(new_n345), .B1(new_n347), .B2(new_n316), .ZN(new_n348));
  AOI21_X1  g162(.A(KEYINPUT28), .B1(new_n329), .B2(new_n261), .ZN(new_n349));
  OAI21_X1  g163(.A(new_n331), .B1(new_n348), .B2(new_n349), .ZN(new_n350));
  NOR3_X1   g164(.A1(new_n315), .A2(new_n251), .A3(new_n322), .ZN(new_n351));
  AOI21_X1  g165(.A(KEYINPUT31), .B1(new_n330), .B2(new_n332), .ZN(new_n352));
  OAI21_X1  g166(.A(new_n350), .B1(new_n351), .B2(new_n352), .ZN(new_n353));
  INV_X1    g167(.A(KEYINPUT32), .ZN(new_n354));
  NAND3_X1  g168(.A1(new_n353), .A2(new_n354), .A3(new_n342), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n344), .A2(new_n355), .ZN(new_n356));
  INV_X1    g170(.A(new_n188), .ZN(new_n357));
  AOI21_X1  g171(.A(new_n338), .B1(new_n347), .B2(new_n316), .ZN(new_n358));
  NOR2_X1   g172(.A1(new_n358), .A2(new_n349), .ZN(new_n359));
  INV_X1    g173(.A(KEYINPUT29), .ZN(new_n360));
  NOR2_X1   g174(.A1(new_n331), .A2(new_n360), .ZN(new_n361));
  AOI21_X1  g175(.A(new_n357), .B1(new_n359), .B2(new_n361), .ZN(new_n362));
  OAI21_X1  g176(.A(new_n316), .B1(new_n305), .B2(new_n314), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n363), .A2(new_n331), .ZN(new_n364));
  OAI211_X1 g178(.A(new_n364), .B(new_n360), .C1(new_n340), .C2(new_n331), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n362), .A2(new_n365), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n366), .A2(G472), .ZN(new_n367));
  AOI21_X1  g181(.A(new_n250), .B1(new_n356), .B2(new_n367), .ZN(new_n368));
  XNOR2_X1  g182(.A(KEYINPUT9), .B(G234), .ZN(new_n369));
  OAI21_X1  g183(.A(G221), .B1(new_n369), .B2(G902), .ZN(new_n370));
  INV_X1    g184(.A(new_n370), .ZN(new_n371));
  INV_X1    g185(.A(G469), .ZN(new_n372));
  INV_X1    g186(.A(G902), .ZN(new_n373));
  NOR2_X1   g187(.A1(new_n372), .A2(new_n373), .ZN(new_n374));
  XNOR2_X1  g188(.A(G110), .B(G140), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n192), .A2(G227), .ZN(new_n376));
  XOR2_X1   g190(.A(new_n375), .B(new_n376), .Z(new_n377));
  INV_X1    g191(.A(new_n328), .ZN(new_n378));
  INV_X1    g192(.A(G107), .ZN(new_n379));
  NOR2_X1   g193(.A1(new_n379), .A2(G104), .ZN(new_n380));
  INV_X1    g194(.A(new_n380), .ZN(new_n381));
  AND3_X1   g195(.A1(new_n379), .A2(KEYINPUT3), .A3(G104), .ZN(new_n382));
  AOI21_X1  g196(.A(KEYINPUT3), .B1(new_n379), .B2(G104), .ZN(new_n383));
  OAI21_X1  g197(.A(new_n381), .B1(new_n382), .B2(new_n383), .ZN(new_n384));
  NAND3_X1  g198(.A1(new_n384), .A2(KEYINPUT72), .A3(G101), .ZN(new_n385));
  INV_X1    g199(.A(KEYINPUT72), .ZN(new_n386));
  INV_X1    g200(.A(KEYINPUT3), .ZN(new_n387));
  INV_X1    g201(.A(G104), .ZN(new_n388));
  OAI21_X1  g202(.A(new_n387), .B1(new_n388), .B2(G107), .ZN(new_n389));
  NAND3_X1  g203(.A1(new_n379), .A2(KEYINPUT3), .A3(G104), .ZN(new_n390));
  AOI21_X1  g204(.A(new_n380), .B1(new_n389), .B2(new_n390), .ZN(new_n391));
  INV_X1    g205(.A(G101), .ZN(new_n392));
  OAI21_X1  g206(.A(new_n386), .B1(new_n391), .B2(new_n392), .ZN(new_n393));
  INV_X1    g207(.A(KEYINPUT4), .ZN(new_n394));
  AOI21_X1  g208(.A(new_n394), .B1(new_n391), .B2(new_n392), .ZN(new_n395));
  NAND3_X1  g209(.A1(new_n385), .A2(new_n393), .A3(new_n395), .ZN(new_n396));
  INV_X1    g210(.A(KEYINPUT73), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n396), .A2(new_n397), .ZN(new_n398));
  NAND4_X1  g212(.A1(new_n385), .A2(new_n393), .A3(new_n395), .A4(KEYINPUT73), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n398), .A2(new_n399), .ZN(new_n400));
  NAND3_X1  g214(.A1(new_n384), .A2(new_n394), .A3(G101), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n307), .A2(new_n401), .ZN(new_n402));
  INV_X1    g216(.A(new_n402), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n400), .A2(new_n403), .ZN(new_n404));
  OAI21_X1  g218(.A(KEYINPUT74), .B1(new_n379), .B2(G104), .ZN(new_n405));
  INV_X1    g219(.A(KEYINPUT74), .ZN(new_n406));
  NAND3_X1  g220(.A1(new_n406), .A2(new_n388), .A3(G107), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n379), .A2(G104), .ZN(new_n408));
  NAND3_X1  g222(.A1(new_n405), .A2(new_n407), .A3(new_n408), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n409), .A2(G101), .ZN(new_n410));
  OAI211_X1 g224(.A(new_n381), .B(new_n392), .C1(new_n382), .C2(new_n383), .ZN(new_n411));
  NAND4_X1  g225(.A1(new_n410), .A2(new_n411), .A3(new_n281), .A4(new_n278), .ZN(new_n412));
  INV_X1    g226(.A(KEYINPUT10), .ZN(new_n413));
  XNOR2_X1  g227(.A(new_n412), .B(new_n413), .ZN(new_n414));
  INV_X1    g228(.A(new_n414), .ZN(new_n415));
  AOI21_X1  g229(.A(new_n378), .B1(new_n404), .B2(new_n415), .ZN(new_n416));
  AOI21_X1  g230(.A(new_n402), .B1(new_n398), .B2(new_n399), .ZN(new_n417));
  NOR3_X1   g231(.A1(new_n417), .A2(new_n328), .A3(new_n414), .ZN(new_n418));
  OAI21_X1  g232(.A(new_n377), .B1(new_n416), .B2(new_n418), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n410), .A2(new_n411), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n420), .A2(new_n311), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n421), .A2(new_n412), .ZN(new_n422));
  XNOR2_X1  g236(.A(KEYINPUT75), .B(KEYINPUT12), .ZN(new_n423));
  NAND3_X1  g237(.A1(new_n422), .A2(new_n328), .A3(new_n423), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n424), .A2(KEYINPUT76), .ZN(new_n425));
  INV_X1    g239(.A(KEYINPUT76), .ZN(new_n426));
  NAND4_X1  g240(.A1(new_n422), .A2(new_n426), .A3(new_n328), .A4(new_n423), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n422), .A2(new_n328), .ZN(new_n428));
  INV_X1    g242(.A(KEYINPUT12), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n428), .A2(new_n429), .ZN(new_n430));
  NAND3_X1  g244(.A1(new_n425), .A2(new_n427), .A3(new_n430), .ZN(new_n431));
  NAND3_X1  g245(.A1(new_n404), .A2(new_n378), .A3(new_n415), .ZN(new_n432));
  INV_X1    g246(.A(new_n377), .ZN(new_n433));
  NAND3_X1  g247(.A1(new_n431), .A2(new_n432), .A3(new_n433), .ZN(new_n434));
  AOI21_X1  g248(.A(new_n357), .B1(new_n419), .B2(new_n434), .ZN(new_n435));
  AOI21_X1  g249(.A(new_n374), .B1(new_n435), .B2(new_n372), .ZN(new_n436));
  INV_X1    g250(.A(KEYINPUT77), .ZN(new_n437));
  AND3_X1   g251(.A1(new_n431), .A2(new_n432), .A3(new_n437), .ZN(new_n438));
  AOI21_X1  g252(.A(new_n437), .B1(new_n431), .B2(new_n432), .ZN(new_n439));
  OAI21_X1  g253(.A(new_n377), .B1(new_n438), .B2(new_n439), .ZN(new_n440));
  NOR2_X1   g254(.A1(new_n417), .A2(new_n414), .ZN(new_n441));
  AOI21_X1  g255(.A(new_n377), .B1(new_n441), .B2(new_n378), .ZN(new_n442));
  OAI21_X1  g256(.A(new_n328), .B1(new_n417), .B2(new_n414), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  NAND3_X1  g258(.A1(new_n440), .A2(G469), .A3(new_n444), .ZN(new_n445));
  AOI21_X1  g259(.A(new_n371), .B1(new_n436), .B2(new_n445), .ZN(new_n446));
  OAI21_X1  g260(.A(G214), .B1(G237), .B2(G902), .ZN(new_n447));
  INV_X1    g261(.A(new_n447), .ZN(new_n448));
  OAI21_X1  g262(.A(new_n401), .B1(new_n259), .B2(new_n260), .ZN(new_n449));
  AOI21_X1  g263(.A(new_n449), .B1(new_n398), .B2(new_n399), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n210), .A2(G116), .ZN(new_n451));
  OAI21_X1  g265(.A(G113), .B1(new_n451), .B2(KEYINPUT5), .ZN(new_n452));
  AOI21_X1  g266(.A(new_n452), .B1(new_n257), .B2(KEYINPUT5), .ZN(new_n453));
  NOR3_X1   g267(.A1(new_n420), .A2(new_n259), .A3(new_n453), .ZN(new_n454));
  XNOR2_X1  g268(.A(G110), .B(G122), .ZN(new_n455));
  INV_X1    g269(.A(new_n455), .ZN(new_n456));
  NOR3_X1   g270(.A1(new_n450), .A2(new_n454), .A3(new_n456), .ZN(new_n457));
  XNOR2_X1  g271(.A(new_n455), .B(KEYINPUT8), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n255), .A2(new_n256), .ZN(new_n459));
  NAND3_X1  g273(.A1(new_n459), .A2(KEYINPUT5), .A3(new_n451), .ZN(new_n460));
  INV_X1    g274(.A(new_n452), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n257), .A2(new_n258), .ZN(new_n463));
  AOI22_X1  g277(.A1(new_n462), .A2(new_n463), .B1(new_n411), .B2(new_n410), .ZN(new_n464));
  OAI21_X1  g278(.A(new_n458), .B1(new_n454), .B2(new_n464), .ZN(new_n465));
  AOI21_X1  g279(.A(G125), .B1(new_n281), .B2(new_n278), .ZN(new_n466));
  AOI21_X1  g280(.A(new_n197), .B1(new_n292), .B2(new_n293), .ZN(new_n467));
  OAI21_X1  g281(.A(KEYINPUT79), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n294), .A2(G125), .ZN(new_n469));
  INV_X1    g283(.A(KEYINPUT79), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n192), .A2(G224), .ZN(new_n472));
  NAND4_X1  g286(.A1(new_n468), .A2(new_n471), .A3(KEYINPUT7), .A4(new_n472), .ZN(new_n473));
  INV_X1    g287(.A(KEYINPUT81), .ZN(new_n474));
  INV_X1    g288(.A(new_n466), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n475), .A2(new_n469), .ZN(new_n476));
  INV_X1    g290(.A(KEYINPUT7), .ZN(new_n477));
  AOI22_X1  g291(.A1(KEYINPUT80), .A2(new_n477), .B1(new_n192), .B2(G224), .ZN(new_n478));
  OAI21_X1  g292(.A(new_n478), .B1(KEYINPUT80), .B2(new_n477), .ZN(new_n479));
  AOI21_X1  g293(.A(new_n474), .B1(new_n476), .B2(new_n479), .ZN(new_n480));
  OAI211_X1 g294(.A(new_n474), .B(new_n479), .C1(new_n466), .C2(new_n467), .ZN(new_n481));
  INV_X1    g295(.A(new_n481), .ZN(new_n482));
  OAI211_X1 g296(.A(new_n465), .B(new_n473), .C1(new_n480), .C2(new_n482), .ZN(new_n483));
  OAI21_X1  g297(.A(new_n373), .B1(new_n457), .B2(new_n483), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n484), .A2(KEYINPUT82), .ZN(new_n485));
  INV_X1    g299(.A(KEYINPUT82), .ZN(new_n486));
  OAI211_X1 g300(.A(new_n486), .B(new_n373), .C1(new_n457), .C2(new_n483), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n485), .A2(new_n487), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n468), .A2(new_n471), .ZN(new_n489));
  XOR2_X1   g303(.A(new_n489), .B(new_n472), .Z(new_n490));
  INV_X1    g304(.A(new_n450), .ZN(new_n491));
  INV_X1    g305(.A(new_n454), .ZN(new_n492));
  NAND3_X1  g306(.A1(new_n491), .A2(new_n492), .A3(new_n455), .ZN(new_n493));
  OAI21_X1  g307(.A(new_n456), .B1(new_n450), .B2(new_n454), .ZN(new_n494));
  NAND3_X1  g308(.A1(new_n493), .A2(KEYINPUT6), .A3(new_n494), .ZN(new_n495));
  INV_X1    g309(.A(KEYINPUT6), .ZN(new_n496));
  OAI211_X1 g310(.A(new_n496), .B(new_n456), .C1(new_n450), .C2(new_n454), .ZN(new_n497));
  INV_X1    g311(.A(KEYINPUT78), .ZN(new_n498));
  AND2_X1   g312(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  NOR2_X1   g313(.A1(new_n497), .A2(new_n498), .ZN(new_n500));
  OAI211_X1 g314(.A(new_n490), .B(new_n495), .C1(new_n499), .C2(new_n500), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n488), .A2(new_n501), .ZN(new_n502));
  OAI21_X1  g316(.A(G210), .B1(G237), .B2(G902), .ZN(new_n503));
  INV_X1    g317(.A(new_n503), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n502), .A2(new_n504), .ZN(new_n505));
  NAND3_X1  g319(.A1(new_n488), .A2(new_n501), .A3(new_n503), .ZN(new_n506));
  AOI21_X1  g320(.A(new_n448), .B1(new_n505), .B2(new_n506), .ZN(new_n507));
  INV_X1    g321(.A(G237), .ZN(new_n508));
  NAND4_X1  g322(.A1(new_n508), .A2(new_n192), .A3(G143), .A4(G214), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n509), .A2(KEYINPUT83), .ZN(new_n510));
  INV_X1    g324(.A(KEYINPUT83), .ZN(new_n511));
  NAND4_X1  g325(.A1(new_n317), .A2(new_n511), .A3(G143), .A4(G214), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n510), .A2(new_n512), .ZN(new_n513));
  AOI21_X1  g327(.A(G143), .B1(new_n317), .B2(G214), .ZN(new_n514));
  INV_X1    g328(.A(new_n514), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n513), .A2(new_n515), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n516), .A2(G131), .ZN(new_n517));
  NOR2_X1   g331(.A1(new_n514), .A2(G131), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n513), .A2(new_n518), .ZN(new_n519));
  INV_X1    g333(.A(KEYINPUT85), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  INV_X1    g335(.A(KEYINPUT17), .ZN(new_n522));
  NAND3_X1  g336(.A1(new_n513), .A2(KEYINPUT85), .A3(new_n518), .ZN(new_n523));
  NAND4_X1  g337(.A1(new_n517), .A2(new_n521), .A3(new_n522), .A4(new_n523), .ZN(new_n524));
  AOI21_X1  g338(.A(new_n514), .B1(new_n510), .B2(new_n512), .ZN(new_n525));
  NOR3_X1   g339(.A1(new_n525), .A2(new_n522), .A3(new_n285), .ZN(new_n526));
  NOR2_X1   g340(.A1(new_n208), .A2(new_n526), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n524), .A2(new_n527), .ZN(new_n528));
  NAND4_X1  g342(.A1(new_n516), .A2(KEYINPUT84), .A3(KEYINPUT18), .A4(G131), .ZN(new_n529));
  INV_X1    g343(.A(KEYINPUT84), .ZN(new_n530));
  NAND2_X1  g344(.A1(KEYINPUT18), .A2(G131), .ZN(new_n531));
  OAI21_X1  g345(.A(new_n530), .B1(new_n525), .B2(new_n531), .ZN(new_n532));
  OR2_X1    g346(.A1(new_n221), .A2(new_n204), .ZN(new_n533));
  AOI22_X1  g347(.A1(new_n525), .A2(new_n531), .B1(new_n533), .B2(new_n222), .ZN(new_n534));
  NAND3_X1  g348(.A1(new_n529), .A2(new_n532), .A3(new_n534), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n528), .A2(new_n535), .ZN(new_n536));
  XNOR2_X1  g350(.A(G113), .B(G122), .ZN(new_n537));
  XNOR2_X1  g351(.A(new_n537), .B(new_n388), .ZN(new_n538));
  INV_X1    g352(.A(new_n538), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n536), .A2(new_n539), .ZN(new_n540));
  NAND3_X1  g354(.A1(new_n528), .A2(new_n538), .A3(new_n535), .ZN(new_n541));
  AOI21_X1  g355(.A(G902), .B1(new_n540), .B2(new_n541), .ZN(new_n542));
  INV_X1    g356(.A(KEYINPUT86), .ZN(new_n543));
  OAI21_X1  g357(.A(G475), .B1(new_n542), .B2(new_n543), .ZN(new_n544));
  AND3_X1   g358(.A1(new_n528), .A2(new_n538), .A3(new_n535), .ZN(new_n545));
  AOI21_X1  g359(.A(new_n538), .B1(new_n528), .B2(new_n535), .ZN(new_n546));
  OAI211_X1 g360(.A(new_n543), .B(new_n373), .C1(new_n545), .C2(new_n546), .ZN(new_n547));
  INV_X1    g361(.A(new_n547), .ZN(new_n548));
  INV_X1    g362(.A(KEYINPUT20), .ZN(new_n549));
  INV_X1    g363(.A(KEYINPUT19), .ZN(new_n550));
  XNOR2_X1  g364(.A(new_n221), .B(new_n550), .ZN(new_n551));
  OAI21_X1  g365(.A(new_n201), .B1(new_n551), .B2(G146), .ZN(new_n552));
  AOI22_X1  g366(.A1(new_n520), .A2(new_n519), .B1(new_n516), .B2(G131), .ZN(new_n553));
  AOI21_X1  g367(.A(new_n552), .B1(new_n553), .B2(new_n523), .ZN(new_n554));
  INV_X1    g368(.A(new_n535), .ZN(new_n555));
  OAI21_X1  g369(.A(new_n539), .B1(new_n554), .B2(new_n555), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n556), .A2(new_n541), .ZN(new_n557));
  NOR2_X1   g371(.A1(G475), .A2(G902), .ZN(new_n558));
  AOI21_X1  g372(.A(new_n549), .B1(new_n557), .B2(new_n558), .ZN(new_n559));
  INV_X1    g373(.A(new_n558), .ZN(new_n560));
  AOI211_X1 g374(.A(KEYINPUT20), .B(new_n560), .C1(new_n556), .C2(new_n541), .ZN(new_n561));
  OAI22_X1  g375(.A1(new_n544), .A2(new_n548), .B1(new_n559), .B2(new_n561), .ZN(new_n562));
  AND2_X1   g376(.A1(new_n192), .A2(G952), .ZN(new_n563));
  INV_X1    g377(.A(G234), .ZN(new_n564));
  OAI21_X1  g378(.A(new_n563), .B1(new_n564), .B2(new_n508), .ZN(new_n565));
  INV_X1    g379(.A(new_n565), .ZN(new_n566));
  AOI211_X1 g380(.A(new_n192), .B(new_n188), .C1(G234), .C2(G237), .ZN(new_n567));
  XNOR2_X1  g381(.A(KEYINPUT21), .B(G898), .ZN(new_n568));
  AOI21_X1  g382(.A(new_n566), .B1(new_n567), .B2(new_n568), .ZN(new_n569));
  INV_X1    g383(.A(KEYINPUT90), .ZN(new_n570));
  INV_X1    g384(.A(KEYINPUT87), .ZN(new_n571));
  OAI21_X1  g385(.A(new_n571), .B1(new_n212), .B2(G143), .ZN(new_n572));
  NAND3_X1  g386(.A1(new_n276), .A2(KEYINPUT87), .A3(G128), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  INV_X1    g388(.A(KEYINPUT88), .ZN(new_n575));
  OAI21_X1  g389(.A(new_n575), .B1(new_n276), .B2(G128), .ZN(new_n576));
  NAND3_X1  g390(.A1(new_n212), .A2(KEYINPUT88), .A3(G143), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  XNOR2_X1  g392(.A(KEYINPUT65), .B(G134), .ZN(new_n579));
  AND3_X1   g393(.A1(new_n574), .A2(new_n578), .A3(new_n579), .ZN(new_n580));
  AOI21_X1  g394(.A(new_n579), .B1(new_n574), .B2(new_n578), .ZN(new_n581));
  NOR2_X1   g395(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  INV_X1    g396(.A(G122), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n583), .A2(G116), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n252), .A2(G122), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n586), .A2(new_n379), .ZN(new_n587));
  NAND3_X1  g401(.A1(new_n584), .A2(new_n585), .A3(G107), .ZN(new_n588));
  NAND3_X1  g402(.A1(new_n584), .A2(KEYINPUT14), .A3(G107), .ZN(new_n589));
  NAND3_X1  g403(.A1(new_n587), .A2(new_n588), .A3(new_n589), .ZN(new_n590));
  NAND4_X1  g404(.A1(new_n584), .A2(new_n585), .A3(KEYINPUT14), .A4(G107), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  OAI21_X1  g406(.A(new_n570), .B1(new_n582), .B2(new_n592), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n574), .A2(new_n578), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n594), .A2(new_n286), .ZN(new_n595));
  NAND3_X1  g409(.A1(new_n574), .A2(new_n578), .A3(new_n579), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  NAND4_X1  g411(.A1(new_n597), .A2(KEYINPUT90), .A3(new_n590), .A4(new_n591), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n593), .A2(new_n598), .ZN(new_n599));
  AND3_X1   g413(.A1(new_n596), .A2(new_n587), .A3(new_n588), .ZN(new_n600));
  NAND3_X1  g414(.A1(new_n572), .A2(KEYINPUT13), .A3(new_n573), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n601), .A2(new_n578), .ZN(new_n602));
  AOI21_X1  g416(.A(KEYINPUT13), .B1(new_n572), .B2(new_n573), .ZN(new_n603));
  OAI211_X1 g417(.A(KEYINPUT89), .B(G134), .C1(new_n602), .C2(new_n603), .ZN(new_n604));
  INV_X1    g418(.A(new_n604), .ZN(new_n605));
  INV_X1    g419(.A(KEYINPUT13), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n574), .A2(new_n606), .ZN(new_n607));
  NAND3_X1  g421(.A1(new_n607), .A2(new_n578), .A3(new_n601), .ZN(new_n608));
  AOI21_X1  g422(.A(KEYINPUT89), .B1(new_n608), .B2(G134), .ZN(new_n609));
  OAI21_X1  g423(.A(new_n600), .B1(new_n605), .B2(new_n609), .ZN(new_n610));
  NOR3_X1   g424(.A1(new_n369), .A2(new_n187), .A3(G953), .ZN(new_n611));
  AND3_X1   g425(.A1(new_n599), .A2(new_n610), .A3(new_n611), .ZN(new_n612));
  AOI21_X1  g426(.A(new_n611), .B1(new_n599), .B2(new_n610), .ZN(new_n613));
  OAI21_X1  g427(.A(new_n188), .B1(new_n612), .B2(new_n613), .ZN(new_n614));
  INV_X1    g428(.A(G478), .ZN(new_n615));
  NOR2_X1   g429(.A1(KEYINPUT91), .A2(KEYINPUT15), .ZN(new_n616));
  INV_X1    g430(.A(new_n616), .ZN(new_n617));
  NAND2_X1  g431(.A1(KEYINPUT91), .A2(KEYINPUT15), .ZN(new_n618));
  AOI21_X1  g432(.A(new_n615), .B1(new_n617), .B2(new_n618), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n614), .A2(new_n619), .ZN(new_n620));
  INV_X1    g434(.A(new_n619), .ZN(new_n621));
  OAI211_X1 g435(.A(new_n188), .B(new_n621), .C1(new_n612), .C2(new_n613), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n620), .A2(new_n622), .ZN(new_n623));
  NOR3_X1   g437(.A1(new_n562), .A2(new_n569), .A3(new_n623), .ZN(new_n624));
  NAND4_X1  g438(.A1(new_n368), .A2(new_n446), .A3(new_n507), .A4(new_n624), .ZN(new_n625));
  XNOR2_X1  g439(.A(new_n625), .B(G101), .ZN(G3));
  INV_X1    g440(.A(KEYINPUT33), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n627), .A2(KEYINPUT92), .ZN(new_n628));
  OR2_X1    g442(.A1(new_n627), .A2(KEYINPUT92), .ZN(new_n629));
  OAI211_X1 g443(.A(new_n628), .B(new_n629), .C1(new_n612), .C2(new_n613), .ZN(new_n630));
  NAND2_X1  g444(.A1(new_n599), .A2(new_n610), .ZN(new_n631));
  INV_X1    g445(.A(new_n611), .ZN(new_n632));
  NAND2_X1  g446(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  NAND3_X1  g447(.A1(new_n599), .A2(new_n610), .A3(new_n611), .ZN(new_n634));
  NAND4_X1  g448(.A1(new_n633), .A2(KEYINPUT92), .A3(new_n627), .A4(new_n634), .ZN(new_n635));
  NAND2_X1  g449(.A1(new_n630), .A2(new_n635), .ZN(new_n636));
  NOR2_X1   g450(.A1(new_n357), .A2(new_n615), .ZN(new_n637));
  AOI22_X1  g451(.A1(new_n636), .A2(new_n637), .B1(new_n615), .B2(new_n614), .ZN(new_n638));
  INV_X1    g452(.A(new_n638), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n639), .A2(new_n562), .ZN(new_n640));
  INV_X1    g454(.A(new_n640), .ZN(new_n641));
  INV_X1    g455(.A(new_n569), .ZN(new_n642));
  NAND3_X1  g456(.A1(new_n507), .A2(new_n641), .A3(new_n642), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n323), .A2(new_n333), .ZN(new_n644));
  AOI21_X1  g458(.A(new_n357), .B1(new_n644), .B2(new_n350), .ZN(new_n645));
  INV_X1    g459(.A(G472), .ZN(new_n646));
  OAI22_X1  g460(.A1(new_n645), .A2(new_n646), .B1(new_n343), .B2(new_n341), .ZN(new_n647));
  NOR2_X1   g461(.A1(new_n647), .A2(new_n250), .ZN(new_n648));
  NAND2_X1  g462(.A1(new_n648), .A2(new_n446), .ZN(new_n649));
  NOR2_X1   g463(.A1(new_n643), .A2(new_n649), .ZN(new_n650));
  XNOR2_X1  g464(.A(KEYINPUT34), .B(G104), .ZN(new_n651));
  XNOR2_X1  g465(.A(new_n650), .B(new_n651), .ZN(G6));
  AND3_X1   g466(.A1(new_n488), .A2(new_n501), .A3(new_n503), .ZN(new_n653));
  AOI21_X1  g467(.A(new_n503), .B1(new_n488), .B2(new_n501), .ZN(new_n654));
  OAI211_X1 g468(.A(new_n447), .B(new_n642), .C1(new_n653), .C2(new_n654), .ZN(new_n655));
  OAI21_X1  g469(.A(KEYINPUT93), .B1(new_n544), .B2(new_n548), .ZN(new_n656));
  INV_X1    g470(.A(G475), .ZN(new_n657));
  OAI21_X1  g471(.A(new_n373), .B1(new_n545), .B2(new_n546), .ZN(new_n658));
  AOI21_X1  g472(.A(new_n657), .B1(new_n658), .B2(KEYINPUT86), .ZN(new_n659));
  INV_X1    g473(.A(KEYINPUT93), .ZN(new_n660));
  NAND3_X1  g474(.A1(new_n659), .A2(new_n660), .A3(new_n547), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n557), .A2(new_n558), .ZN(new_n662));
  NAND2_X1  g476(.A1(new_n662), .A2(KEYINPUT20), .ZN(new_n663));
  NAND3_X1  g477(.A1(new_n557), .A2(new_n549), .A3(new_n558), .ZN(new_n664));
  AOI22_X1  g478(.A1(new_n663), .A2(new_n664), .B1(new_n620), .B2(new_n622), .ZN(new_n665));
  NAND3_X1  g479(.A1(new_n656), .A2(new_n661), .A3(new_n665), .ZN(new_n666));
  NOR2_X1   g480(.A1(new_n655), .A2(new_n666), .ZN(new_n667));
  NAND3_X1  g481(.A1(new_n667), .A2(new_n446), .A3(new_n648), .ZN(new_n668));
  XOR2_X1   g482(.A(KEYINPUT35), .B(G107), .Z(new_n669));
  XNOR2_X1  g483(.A(new_n668), .B(new_n669), .ZN(G9));
  INV_X1    g484(.A(KEYINPUT36), .ZN(new_n671));
  NAND2_X1  g485(.A1(new_n194), .A2(new_n671), .ZN(new_n672));
  XNOR2_X1  g486(.A(new_n229), .B(new_n672), .ZN(new_n673));
  NAND2_X1  g487(.A1(new_n673), .A2(new_n248), .ZN(new_n674));
  INV_X1    g488(.A(new_n674), .ZN(new_n675));
  NOR2_X1   g489(.A1(new_n236), .A2(new_n675), .ZN(new_n676));
  NOR2_X1   g490(.A1(new_n647), .A2(new_n676), .ZN(new_n677));
  NAND4_X1  g491(.A1(new_n677), .A2(new_n507), .A3(new_n446), .A4(new_n624), .ZN(new_n678));
  XNOR2_X1  g492(.A(new_n678), .B(KEYINPUT94), .ZN(new_n679));
  XNOR2_X1  g493(.A(KEYINPUT37), .B(G110), .ZN(new_n680));
  XNOR2_X1  g494(.A(new_n679), .B(new_n680), .ZN(G12));
  AOI22_X1  g495(.A1(new_n344), .A2(new_n355), .B1(G472), .B2(new_n366), .ZN(new_n682));
  INV_X1    g496(.A(G900), .ZN(new_n683));
  AOI21_X1  g497(.A(new_n566), .B1(new_n567), .B2(new_n683), .ZN(new_n684));
  INV_X1    g498(.A(new_n684), .ZN(new_n685));
  NAND4_X1  g499(.A1(new_n656), .A2(new_n661), .A3(new_n665), .A4(new_n685), .ZN(new_n686));
  NOR3_X1   g500(.A1(new_n682), .A2(new_n686), .A3(new_n676), .ZN(new_n687));
  AND3_X1   g501(.A1(new_n440), .A2(G469), .A3(new_n444), .ZN(new_n688));
  NAND2_X1  g502(.A1(new_n419), .A2(new_n434), .ZN(new_n689));
  NAND3_X1  g503(.A1(new_n689), .A2(new_n372), .A3(new_n188), .ZN(new_n690));
  INV_X1    g504(.A(new_n374), .ZN(new_n691));
  NAND2_X1  g505(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  OAI21_X1  g506(.A(new_n370), .B1(new_n688), .B2(new_n692), .ZN(new_n693));
  OAI21_X1  g507(.A(new_n447), .B1(new_n653), .B2(new_n654), .ZN(new_n694));
  NOR2_X1   g508(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  NAND3_X1  g509(.A1(new_n687), .A2(new_n695), .A3(KEYINPUT95), .ZN(new_n696));
  INV_X1    g510(.A(KEYINPUT95), .ZN(new_n697));
  AND4_X1   g511(.A1(new_n656), .A2(new_n661), .A3(new_n665), .A4(new_n685), .ZN(new_n698));
  NOR3_X1   g512(.A1(new_n341), .A2(KEYINPUT32), .A3(new_n343), .ZN(new_n699));
  AOI21_X1  g513(.A(new_n354), .B1(new_n353), .B2(new_n342), .ZN(new_n700));
  OAI21_X1  g514(.A(new_n367), .B1(new_n699), .B2(new_n700), .ZN(new_n701));
  AOI21_X1  g515(.A(KEYINPUT25), .B1(new_n247), .B2(new_n188), .ZN(new_n702));
  INV_X1    g516(.A(new_n235), .ZN(new_n703));
  OAI21_X1  g517(.A(new_n189), .B1(new_n702), .B2(new_n703), .ZN(new_n704));
  NAND2_X1  g518(.A1(new_n704), .A2(new_n674), .ZN(new_n705));
  NAND3_X1  g519(.A1(new_n698), .A2(new_n701), .A3(new_n705), .ZN(new_n706));
  NAND2_X1  g520(.A1(new_n505), .A2(new_n506), .ZN(new_n707));
  NAND3_X1  g521(.A1(new_n707), .A2(new_n446), .A3(new_n447), .ZN(new_n708));
  OAI21_X1  g522(.A(new_n697), .B1(new_n706), .B2(new_n708), .ZN(new_n709));
  NAND2_X1  g523(.A1(new_n696), .A2(new_n709), .ZN(new_n710));
  XNOR2_X1  g524(.A(new_n710), .B(G128), .ZN(G30));
  XOR2_X1   g525(.A(new_n684), .B(KEYINPUT39), .Z(new_n712));
  NAND2_X1  g526(.A1(new_n446), .A2(new_n712), .ZN(new_n713));
  XOR2_X1   g527(.A(new_n713), .B(KEYINPUT100), .Z(new_n714));
  OR2_X1    g528(.A1(new_n714), .A2(KEYINPUT40), .ZN(new_n715));
  XOR2_X1   g529(.A(new_n707), .B(KEYINPUT96), .Z(new_n716));
  XNOR2_X1  g530(.A(KEYINPUT97), .B(KEYINPUT38), .ZN(new_n717));
  XNOR2_X1  g531(.A(new_n716), .B(new_n717), .ZN(new_n718));
  NAND2_X1  g532(.A1(new_n714), .A2(KEYINPUT40), .ZN(new_n719));
  NAND3_X1  g533(.A1(new_n562), .A2(new_n447), .A3(new_n623), .ZN(new_n720));
  INV_X1    g534(.A(new_n720), .ZN(new_n721));
  NAND2_X1  g535(.A1(new_n721), .A2(new_n676), .ZN(new_n722));
  XNOR2_X1  g536(.A(new_n722), .B(KEYINPUT99), .ZN(new_n723));
  NAND2_X1  g537(.A1(new_n330), .A2(new_n332), .ZN(new_n724));
  AOI21_X1  g538(.A(new_n321), .B1(new_n347), .B2(new_n316), .ZN(new_n725));
  INV_X1    g539(.A(KEYINPUT98), .ZN(new_n726));
  OAI21_X1  g540(.A(new_n724), .B1(new_n725), .B2(new_n726), .ZN(new_n727));
  AND2_X1   g541(.A1(new_n725), .A2(new_n726), .ZN(new_n728));
  OAI21_X1  g542(.A(new_n373), .B1(new_n727), .B2(new_n728), .ZN(new_n729));
  NAND2_X1  g543(.A1(new_n729), .A2(G472), .ZN(new_n730));
  NAND2_X1  g544(.A1(new_n356), .A2(new_n730), .ZN(new_n731));
  AND2_X1   g545(.A1(new_n723), .A2(new_n731), .ZN(new_n732));
  NAND4_X1  g546(.A1(new_n715), .A2(new_n718), .A3(new_n719), .A4(new_n732), .ZN(new_n733));
  XNOR2_X1  g547(.A(new_n733), .B(G143), .ZN(G45));
  NAND3_X1  g548(.A1(new_n639), .A2(new_n562), .A3(new_n685), .ZN(new_n735));
  NOR3_X1   g549(.A1(new_n682), .A2(new_n735), .A3(new_n676), .ZN(new_n736));
  NAND2_X1  g550(.A1(new_n736), .A2(new_n695), .ZN(new_n737));
  XNOR2_X1  g551(.A(KEYINPUT101), .B(G146), .ZN(new_n738));
  XNOR2_X1  g552(.A(new_n737), .B(new_n738), .ZN(G48));
  NAND2_X1  g553(.A1(new_n432), .A2(new_n443), .ZN(new_n740));
  AOI22_X1  g554(.A1(new_n377), .A2(new_n740), .B1(new_n442), .B2(new_n431), .ZN(new_n741));
  OAI21_X1  g555(.A(G469), .B1(new_n741), .B2(new_n357), .ZN(new_n742));
  NAND3_X1  g556(.A1(new_n742), .A2(new_n370), .A3(new_n690), .ZN(new_n743));
  INV_X1    g557(.A(KEYINPUT102), .ZN(new_n744));
  NAND2_X1  g558(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  NAND4_X1  g559(.A1(new_n742), .A2(KEYINPUT102), .A3(new_n370), .A4(new_n690), .ZN(new_n746));
  AND2_X1   g560(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  INV_X1    g561(.A(new_n655), .ZN(new_n748));
  NAND4_X1  g562(.A1(new_n747), .A2(new_n368), .A3(new_n641), .A4(new_n748), .ZN(new_n749));
  XNOR2_X1  g563(.A(KEYINPUT41), .B(G113), .ZN(new_n750));
  XNOR2_X1  g564(.A(new_n749), .B(new_n750), .ZN(G15));
  NAND3_X1  g565(.A1(new_n747), .A2(new_n667), .A3(new_n368), .ZN(new_n752));
  XNOR2_X1  g566(.A(new_n752), .B(G116), .ZN(G18));
  NOR2_X1   g567(.A1(new_n694), .A2(new_n743), .ZN(new_n754));
  AOI21_X1  g568(.A(new_n676), .B1(new_n356), .B2(new_n367), .ZN(new_n755));
  NAND3_X1  g569(.A1(new_n754), .A2(new_n624), .A3(new_n755), .ZN(new_n756));
  XNOR2_X1  g570(.A(new_n756), .B(G119), .ZN(G21));
  AOI21_X1  g571(.A(new_n720), .B1(new_n505), .B2(new_n506), .ZN(new_n758));
  OAI21_X1  g572(.A(new_n331), .B1(new_n358), .B2(new_n349), .ZN(new_n759));
  OAI21_X1  g573(.A(new_n759), .B1(new_n351), .B2(new_n352), .ZN(new_n760));
  NAND2_X1  g574(.A1(new_n760), .A2(new_n342), .ZN(new_n761));
  XOR2_X1   g575(.A(KEYINPUT103), .B(G472), .Z(new_n762));
  INV_X1    g576(.A(new_n762), .ZN(new_n763));
  OAI21_X1  g577(.A(new_n761), .B1(new_n645), .B2(new_n763), .ZN(new_n764));
  NOR3_X1   g578(.A1(new_n764), .A2(new_n250), .A3(new_n569), .ZN(new_n765));
  NAND3_X1  g579(.A1(new_n747), .A2(new_n758), .A3(new_n765), .ZN(new_n766));
  XNOR2_X1  g580(.A(new_n766), .B(G122), .ZN(G24));
  INV_X1    g581(.A(KEYINPUT104), .ZN(new_n768));
  OAI21_X1  g582(.A(new_n768), .B1(new_n764), .B2(new_n676), .ZN(new_n769));
  OAI21_X1  g583(.A(new_n762), .B1(new_n341), .B2(new_n357), .ZN(new_n770));
  NAND4_X1  g584(.A1(new_n705), .A2(new_n770), .A3(KEYINPUT104), .A4(new_n761), .ZN(new_n771));
  NAND2_X1  g585(.A1(new_n769), .A2(new_n771), .ZN(new_n772));
  INV_X1    g586(.A(new_n735), .ZN(new_n773));
  NAND3_X1  g587(.A1(new_n772), .A2(new_n754), .A3(new_n773), .ZN(new_n774));
  XNOR2_X1  g588(.A(new_n774), .B(G125), .ZN(G27));
  NOR3_X1   g589(.A1(new_n653), .A2(new_n654), .A3(new_n448), .ZN(new_n776));
  AOI22_X1  g590(.A1(new_n659), .A2(new_n547), .B1(new_n663), .B2(new_n664), .ZN(new_n777));
  NOR4_X1   g591(.A1(new_n777), .A2(new_n638), .A3(KEYINPUT42), .A4(new_n684), .ZN(new_n778));
  AND4_X1   g592(.A1(new_n368), .A2(new_n446), .A3(new_n776), .A4(new_n778), .ZN(new_n779));
  NAND3_X1  g593(.A1(new_n505), .A2(new_n447), .A3(new_n506), .ZN(new_n780));
  NOR2_X1   g594(.A1(new_n693), .A2(new_n780), .ZN(new_n781));
  INV_X1    g595(.A(KEYINPUT105), .ZN(new_n782));
  OAI21_X1  g596(.A(new_n782), .B1(new_n682), .B2(new_n250), .ZN(new_n783));
  INV_X1    g597(.A(new_n250), .ZN(new_n784));
  NAND3_X1  g598(.A1(new_n701), .A2(KEYINPUT105), .A3(new_n784), .ZN(new_n785));
  NAND4_X1  g599(.A1(new_n781), .A2(new_n783), .A3(new_n785), .A4(new_n773), .ZN(new_n786));
  AOI21_X1  g600(.A(new_n779), .B1(new_n786), .B2(KEYINPUT42), .ZN(new_n787));
  XNOR2_X1  g601(.A(new_n787), .B(G131), .ZN(G33));
  NAND2_X1  g602(.A1(new_n776), .A2(new_n446), .ZN(new_n789));
  NAND2_X1  g603(.A1(new_n701), .A2(new_n784), .ZN(new_n790));
  NOR3_X1   g604(.A1(new_n789), .A2(new_n790), .A3(new_n686), .ZN(new_n791));
  XNOR2_X1  g605(.A(new_n791), .B(new_n263), .ZN(G36));
  AOI21_X1  g606(.A(KEYINPUT45), .B1(new_n440), .B2(new_n444), .ZN(new_n793));
  NOR2_X1   g607(.A1(new_n793), .A2(new_n372), .ZN(new_n794));
  NAND3_X1  g608(.A1(new_n440), .A2(KEYINPUT45), .A3(new_n444), .ZN(new_n795));
  NAND2_X1  g609(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  AOI21_X1  g610(.A(KEYINPUT46), .B1(new_n796), .B2(new_n691), .ZN(new_n797));
  AOI21_X1  g611(.A(new_n797), .B1(new_n372), .B2(new_n435), .ZN(new_n798));
  NAND3_X1  g612(.A1(new_n796), .A2(KEYINPUT46), .A3(new_n691), .ZN(new_n799));
  AOI21_X1  g613(.A(new_n371), .B1(new_n798), .B2(new_n799), .ZN(new_n800));
  NAND2_X1  g614(.A1(new_n800), .A2(new_n712), .ZN(new_n801));
  NOR2_X1   g615(.A1(new_n562), .A2(new_n638), .ZN(new_n802));
  OAI21_X1  g616(.A(new_n802), .B1(KEYINPUT106), .B2(KEYINPUT43), .ZN(new_n803));
  XOR2_X1   g617(.A(KEYINPUT106), .B(KEYINPUT43), .Z(new_n804));
  OAI21_X1  g618(.A(new_n803), .B1(new_n802), .B2(new_n804), .ZN(new_n805));
  NAND3_X1  g619(.A1(new_n805), .A2(new_n647), .A3(new_n705), .ZN(new_n806));
  INV_X1    g620(.A(KEYINPUT44), .ZN(new_n807));
  AOI21_X1  g621(.A(new_n780), .B1(new_n806), .B2(new_n807), .ZN(new_n808));
  OAI21_X1  g622(.A(new_n808), .B1(new_n807), .B2(new_n806), .ZN(new_n809));
  NOR2_X1   g623(.A1(new_n801), .A2(new_n809), .ZN(new_n810));
  XNOR2_X1  g624(.A(new_n810), .B(new_n268), .ZN(G39));
  INV_X1    g625(.A(KEYINPUT47), .ZN(new_n812));
  XNOR2_X1  g626(.A(new_n800), .B(new_n812), .ZN(new_n813));
  NOR4_X1   g627(.A1(new_n780), .A2(new_n701), .A3(new_n735), .A4(new_n784), .ZN(new_n814));
  INV_X1    g628(.A(new_n814), .ZN(new_n815));
  NOR2_X1   g629(.A1(new_n813), .A2(new_n815), .ZN(new_n816));
  XNOR2_X1  g630(.A(new_n816), .B(new_n195), .ZN(G42));
  INV_X1    g631(.A(new_n623), .ZN(new_n818));
  OAI21_X1  g632(.A(new_n640), .B1(new_n562), .B2(new_n818), .ZN(new_n819));
  NAND4_X1  g633(.A1(new_n748), .A2(new_n446), .A3(new_n648), .A4(new_n819), .ZN(new_n820));
  AND3_X1   g634(.A1(new_n820), .A2(new_n625), .A3(new_n678), .ZN(new_n821));
  INV_X1    g635(.A(new_n791), .ZN(new_n822));
  NAND3_X1  g636(.A1(new_n620), .A2(new_n622), .A3(new_n685), .ZN(new_n823));
  NOR2_X1   g637(.A1(new_n559), .A2(new_n561), .ZN(new_n824));
  NOR2_X1   g638(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  NAND4_X1  g639(.A1(new_n825), .A2(new_n656), .A3(KEYINPUT108), .A4(new_n661), .ZN(new_n826));
  NAND3_X1  g640(.A1(new_n825), .A2(new_n656), .A3(new_n661), .ZN(new_n827));
  INV_X1    g641(.A(KEYINPUT108), .ZN(new_n828));
  NAND2_X1  g642(.A1(new_n827), .A2(new_n828), .ZN(new_n829));
  AND3_X1   g643(.A1(new_n755), .A2(new_n826), .A3(new_n829), .ZN(new_n830));
  AOI21_X1  g644(.A(new_n735), .B1(new_n769), .B2(new_n771), .ZN(new_n831));
  OAI21_X1  g645(.A(new_n781), .B1(new_n830), .B2(new_n831), .ZN(new_n832));
  NAND3_X1  g646(.A1(new_n821), .A2(new_n822), .A3(new_n832), .ZN(new_n833));
  NAND2_X1  g647(.A1(new_n786), .A2(KEYINPUT42), .ZN(new_n834));
  INV_X1    g648(.A(new_n779), .ZN(new_n835));
  NAND2_X1  g649(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  NAND4_X1  g650(.A1(new_n749), .A2(new_n752), .A3(new_n766), .A4(new_n756), .ZN(new_n837));
  NOR3_X1   g651(.A1(new_n833), .A2(new_n836), .A3(new_n837), .ZN(new_n838));
  INV_X1    g652(.A(KEYINPUT52), .ZN(new_n839));
  AND2_X1   g653(.A1(new_n696), .A2(new_n709), .ZN(new_n840));
  NOR3_X1   g654(.A1(new_n236), .A2(new_n675), .A3(new_n684), .ZN(new_n841));
  OAI211_X1 g655(.A(new_n841), .B(new_n370), .C1(new_n688), .C2(new_n692), .ZN(new_n842));
  NAND2_X1  g656(.A1(new_n842), .A2(KEYINPUT109), .ZN(new_n843));
  INV_X1    g657(.A(KEYINPUT109), .ZN(new_n844));
  NAND3_X1  g658(.A1(new_n446), .A2(new_n844), .A3(new_n841), .ZN(new_n845));
  NAND4_X1  g659(.A1(new_n843), .A2(new_n731), .A3(new_n758), .A4(new_n845), .ZN(new_n846));
  NAND3_X1  g660(.A1(new_n846), .A2(new_n774), .A3(new_n737), .ZN(new_n847));
  OAI21_X1  g661(.A(new_n839), .B1(new_n840), .B2(new_n847), .ZN(new_n848));
  AND2_X1   g662(.A1(new_n774), .A2(new_n737), .ZN(new_n849));
  NAND4_X1  g663(.A1(new_n849), .A2(new_n710), .A3(KEYINPUT52), .A4(new_n846), .ZN(new_n850));
  NAND2_X1  g664(.A1(new_n848), .A2(new_n850), .ZN(new_n851));
  AOI21_X1  g665(.A(KEYINPUT53), .B1(new_n838), .B2(new_n851), .ZN(new_n852));
  INV_X1    g666(.A(KEYINPUT53), .ZN(new_n853));
  NOR3_X1   g667(.A1(new_n836), .A2(new_n837), .A3(new_n853), .ZN(new_n854));
  INV_X1    g668(.A(KEYINPUT110), .ZN(new_n855));
  NAND2_X1  g669(.A1(new_n833), .A2(new_n855), .ZN(new_n856));
  NAND2_X1  g670(.A1(new_n353), .A2(new_n188), .ZN(new_n857));
  AOI22_X1  g671(.A1(new_n857), .A2(new_n762), .B1(new_n342), .B2(new_n760), .ZN(new_n858));
  AOI21_X1  g672(.A(KEYINPUT104), .B1(new_n858), .B2(new_n705), .ZN(new_n859));
  AND4_X1   g673(.A1(KEYINPUT104), .A2(new_n705), .A3(new_n770), .A4(new_n761), .ZN(new_n860));
  OAI21_X1  g674(.A(new_n773), .B1(new_n859), .B2(new_n860), .ZN(new_n861));
  NAND3_X1  g675(.A1(new_n755), .A2(new_n829), .A3(new_n826), .ZN(new_n862));
  NAND2_X1  g676(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  AOI21_X1  g677(.A(new_n791), .B1(new_n863), .B2(new_n781), .ZN(new_n864));
  NAND3_X1  g678(.A1(new_n864), .A2(KEYINPUT110), .A3(new_n821), .ZN(new_n865));
  NAND4_X1  g679(.A1(new_n851), .A2(new_n854), .A3(new_n856), .A4(new_n865), .ZN(new_n866));
  INV_X1    g680(.A(KEYINPUT111), .ZN(new_n867));
  NAND2_X1  g681(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  NOR2_X1   g682(.A1(new_n764), .A2(new_n250), .ZN(new_n869));
  NAND4_X1  g683(.A1(new_n869), .A2(new_n745), .A3(new_n642), .A4(new_n746), .ZN(new_n870));
  NAND2_X1  g684(.A1(new_n721), .A2(new_n707), .ZN(new_n871));
  INV_X1    g685(.A(new_n743), .ZN(new_n872));
  NAND2_X1  g686(.A1(new_n507), .A2(new_n872), .ZN(new_n873));
  NAND3_X1  g687(.A1(new_n701), .A2(new_n624), .A3(new_n705), .ZN(new_n874));
  OAI22_X1  g688(.A1(new_n870), .A2(new_n871), .B1(new_n873), .B2(new_n874), .ZN(new_n875));
  NAND3_X1  g689(.A1(new_n368), .A2(new_n745), .A3(new_n746), .ZN(new_n876));
  NOR2_X1   g690(.A1(new_n876), .A2(new_n643), .ZN(new_n877));
  NOR2_X1   g691(.A1(new_n875), .A2(new_n877), .ZN(new_n878));
  NAND4_X1  g692(.A1(new_n878), .A2(new_n787), .A3(KEYINPUT53), .A4(new_n752), .ZN(new_n879));
  AOI21_X1  g693(.A(new_n879), .B1(new_n848), .B2(new_n850), .ZN(new_n880));
  NAND3_X1  g694(.A1(new_n820), .A2(new_n625), .A3(new_n678), .ZN(new_n881));
  AOI21_X1  g695(.A(new_n789), .B1(new_n861), .B2(new_n862), .ZN(new_n882));
  NOR4_X1   g696(.A1(new_n881), .A2(new_n882), .A3(new_n855), .A4(new_n791), .ZN(new_n883));
  AOI21_X1  g697(.A(KEYINPUT110), .B1(new_n864), .B2(new_n821), .ZN(new_n884));
  NOR2_X1   g698(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  NAND3_X1  g699(.A1(new_n880), .A2(KEYINPUT111), .A3(new_n885), .ZN(new_n886));
  AOI21_X1  g700(.A(new_n852), .B1(new_n868), .B2(new_n886), .ZN(new_n887));
  INV_X1    g701(.A(KEYINPUT54), .ZN(new_n888));
  NAND2_X1  g702(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  NAND2_X1  g703(.A1(new_n838), .A2(new_n851), .ZN(new_n890));
  XNOR2_X1  g704(.A(new_n890), .B(new_n853), .ZN(new_n891));
  NAND2_X1  g705(.A1(new_n891), .A2(KEYINPUT54), .ZN(new_n892));
  AND2_X1   g706(.A1(new_n889), .A2(new_n892), .ZN(new_n893));
  NAND3_X1  g707(.A1(new_n742), .A2(new_n371), .A3(new_n690), .ZN(new_n894));
  NAND2_X1  g708(.A1(new_n813), .A2(new_n894), .ZN(new_n895));
  NAND2_X1  g709(.A1(new_n805), .A2(new_n566), .ZN(new_n896));
  NOR3_X1   g710(.A1(new_n896), .A2(new_n250), .A3(new_n764), .ZN(new_n897));
  AND2_X1   g711(.A1(new_n897), .A2(new_n776), .ZN(new_n898));
  AND2_X1   g712(.A1(new_n895), .A2(new_n898), .ZN(new_n899));
  INV_X1    g713(.A(KEYINPUT51), .ZN(new_n900));
  NAND2_X1  g714(.A1(new_n776), .A2(new_n872), .ZN(new_n901));
  NOR2_X1   g715(.A1(new_n896), .A2(new_n901), .ZN(new_n902));
  OR2_X1    g716(.A1(new_n902), .A2(KEYINPUT113), .ZN(new_n903));
  NAND2_X1  g717(.A1(new_n902), .A2(KEYINPUT113), .ZN(new_n904));
  NAND2_X1  g718(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  NAND2_X1  g719(.A1(new_n905), .A2(new_n772), .ZN(new_n906));
  NOR4_X1   g720(.A1(new_n901), .A2(new_n250), .A3(new_n565), .A4(new_n731), .ZN(new_n907));
  NAND3_X1  g721(.A1(new_n907), .A2(new_n777), .A3(new_n638), .ZN(new_n908));
  XOR2_X1   g722(.A(new_n908), .B(KEYINPUT114), .Z(new_n909));
  INV_X1    g723(.A(new_n718), .ZN(new_n910));
  NOR2_X1   g724(.A1(KEYINPUT112), .A2(KEYINPUT50), .ZN(new_n911));
  NOR2_X1   g725(.A1(new_n743), .A2(new_n447), .ZN(new_n912));
  NAND4_X1  g726(.A1(new_n910), .A2(new_n897), .A3(new_n911), .A4(new_n912), .ZN(new_n913));
  XOR2_X1   g727(.A(KEYINPUT112), .B(KEYINPUT50), .Z(new_n914));
  NAND2_X1  g728(.A1(new_n897), .A2(new_n912), .ZN(new_n915));
  OAI21_X1  g729(.A(new_n914), .B1(new_n915), .B2(new_n718), .ZN(new_n916));
  NAND4_X1  g730(.A1(new_n906), .A2(new_n909), .A3(new_n913), .A4(new_n916), .ZN(new_n917));
  NOR3_X1   g731(.A1(new_n899), .A2(new_n900), .A3(new_n917), .ZN(new_n918));
  INV_X1    g732(.A(new_n897), .ZN(new_n919));
  OAI21_X1  g733(.A(new_n563), .B1(new_n919), .B2(new_n873), .ZN(new_n920));
  AOI21_X1  g734(.A(new_n920), .B1(new_n641), .B2(new_n907), .ZN(new_n921));
  NAND2_X1  g735(.A1(new_n783), .A2(new_n785), .ZN(new_n922));
  AOI21_X1  g736(.A(new_n922), .B1(new_n903), .B2(new_n904), .ZN(new_n923));
  XOR2_X1   g737(.A(KEYINPUT116), .B(KEYINPUT48), .Z(new_n924));
  OAI21_X1  g738(.A(new_n921), .B1(new_n923), .B2(new_n924), .ZN(new_n925));
  INV_X1    g739(.A(KEYINPUT48), .ZN(new_n926));
  NOR2_X1   g740(.A1(new_n926), .A2(KEYINPUT116), .ZN(new_n927));
  AND2_X1   g741(.A1(new_n923), .A2(new_n927), .ZN(new_n928));
  OR2_X1    g742(.A1(new_n925), .A2(new_n928), .ZN(new_n929));
  NOR2_X1   g743(.A1(new_n918), .A2(new_n929), .ZN(new_n930));
  OAI21_X1  g744(.A(new_n900), .B1(new_n899), .B2(new_n917), .ZN(new_n931));
  INV_X1    g745(.A(KEYINPUT115), .ZN(new_n932));
  AND2_X1   g746(.A1(new_n931), .A2(new_n932), .ZN(new_n933));
  NOR2_X1   g747(.A1(new_n931), .A2(new_n932), .ZN(new_n934));
  OAI211_X1 g748(.A(new_n893), .B(new_n930), .C1(new_n933), .C2(new_n934), .ZN(new_n935));
  OAI21_X1  g749(.A(new_n935), .B1(G952), .B2(G953), .ZN(new_n936));
  NAND2_X1  g750(.A1(new_n742), .A2(new_n690), .ZN(new_n937));
  AOI21_X1  g751(.A(new_n731), .B1(KEYINPUT49), .B2(new_n937), .ZN(new_n938));
  OAI21_X1  g752(.A(new_n938), .B1(KEYINPUT49), .B2(new_n937), .ZN(new_n939));
  INV_X1    g753(.A(KEYINPUT107), .ZN(new_n940));
  NAND4_X1  g754(.A1(new_n784), .A2(new_n802), .A3(new_n370), .A4(new_n447), .ZN(new_n941));
  AOI21_X1  g755(.A(new_n939), .B1(new_n940), .B2(new_n941), .ZN(new_n942));
  OAI211_X1 g756(.A(new_n910), .B(new_n942), .C1(new_n940), .C2(new_n941), .ZN(new_n943));
  NAND2_X1  g757(.A1(new_n936), .A2(new_n943), .ZN(G75));
  OAI21_X1  g758(.A(new_n495), .B1(new_n499), .B2(new_n500), .ZN(new_n945));
  XNOR2_X1  g759(.A(new_n945), .B(new_n490), .ZN(new_n946));
  XOR2_X1   g760(.A(new_n946), .B(KEYINPUT55), .Z(new_n947));
  NOR3_X1   g761(.A1(new_n887), .A2(new_n188), .A3(new_n503), .ZN(new_n948));
  OAI21_X1  g762(.A(new_n947), .B1(new_n948), .B2(KEYINPUT56), .ZN(new_n949));
  INV_X1    g763(.A(new_n852), .ZN(new_n950));
  NAND2_X1  g764(.A1(new_n851), .A2(new_n854), .ZN(new_n951));
  NAND2_X1  g765(.A1(new_n856), .A2(new_n865), .ZN(new_n952));
  NOR3_X1   g766(.A1(new_n951), .A2(new_n952), .A3(new_n867), .ZN(new_n953));
  AOI21_X1  g767(.A(KEYINPUT111), .B1(new_n880), .B2(new_n885), .ZN(new_n954));
  OAI21_X1  g768(.A(new_n950), .B1(new_n953), .B2(new_n954), .ZN(new_n955));
  NAND3_X1  g769(.A1(new_n955), .A2(new_n357), .A3(new_n504), .ZN(new_n956));
  INV_X1    g770(.A(KEYINPUT56), .ZN(new_n957));
  INV_X1    g771(.A(new_n947), .ZN(new_n958));
  NAND3_X1  g772(.A1(new_n956), .A2(new_n957), .A3(new_n958), .ZN(new_n959));
  NOR2_X1   g773(.A1(new_n192), .A2(G952), .ZN(new_n960));
  INV_X1    g774(.A(new_n960), .ZN(new_n961));
  NAND3_X1  g775(.A1(new_n949), .A2(new_n959), .A3(new_n961), .ZN(new_n962));
  NAND2_X1  g776(.A1(new_n962), .A2(KEYINPUT117), .ZN(new_n963));
  INV_X1    g777(.A(KEYINPUT117), .ZN(new_n964));
  NAND4_X1  g778(.A1(new_n949), .A2(new_n964), .A3(new_n959), .A4(new_n961), .ZN(new_n965));
  NAND2_X1  g779(.A1(new_n963), .A2(new_n965), .ZN(G51));
  INV_X1    g780(.A(KEYINPUT118), .ZN(new_n967));
  NOR3_X1   g781(.A1(new_n887), .A2(new_n188), .A3(new_n796), .ZN(new_n968));
  XNOR2_X1  g782(.A(new_n374), .B(KEYINPUT57), .ZN(new_n969));
  NAND2_X1  g783(.A1(new_n868), .A2(new_n886), .ZN(new_n970));
  AOI21_X1  g784(.A(new_n888), .B1(new_n970), .B2(new_n950), .ZN(new_n971));
  AOI211_X1 g785(.A(KEYINPUT54), .B(new_n852), .C1(new_n868), .C2(new_n886), .ZN(new_n972));
  OAI21_X1  g786(.A(new_n969), .B1(new_n971), .B2(new_n972), .ZN(new_n973));
  AOI21_X1  g787(.A(new_n968), .B1(new_n973), .B2(new_n689), .ZN(new_n974));
  OAI21_X1  g788(.A(new_n967), .B1(new_n974), .B2(new_n960), .ZN(new_n975));
  NAND2_X1  g789(.A1(new_n955), .A2(KEYINPUT54), .ZN(new_n976));
  NAND2_X1  g790(.A1(new_n976), .A2(new_n889), .ZN(new_n977));
  AOI21_X1  g791(.A(new_n741), .B1(new_n977), .B2(new_n969), .ZN(new_n978));
  OAI211_X1 g792(.A(KEYINPUT118), .B(new_n961), .C1(new_n978), .C2(new_n968), .ZN(new_n979));
  NAND2_X1  g793(.A1(new_n975), .A2(new_n979), .ZN(G54));
  NOR2_X1   g794(.A1(new_n887), .A2(new_n188), .ZN(new_n981));
  INV_X1    g795(.A(KEYINPUT58), .ZN(new_n982));
  OR3_X1    g796(.A1(new_n982), .A2(new_n657), .A3(KEYINPUT119), .ZN(new_n983));
  OAI21_X1  g797(.A(KEYINPUT119), .B1(new_n982), .B2(new_n657), .ZN(new_n984));
  AND2_X1   g798(.A1(new_n983), .A2(new_n984), .ZN(new_n985));
  AND3_X1   g799(.A1(new_n981), .A2(new_n557), .A3(new_n985), .ZN(new_n986));
  AOI21_X1  g800(.A(new_n557), .B1(new_n981), .B2(new_n985), .ZN(new_n987));
  NOR3_X1   g801(.A1(new_n986), .A2(new_n987), .A3(new_n960), .ZN(G60));
  NAND2_X1  g802(.A1(G478), .A2(G902), .ZN(new_n989));
  XOR2_X1   g803(.A(new_n989), .B(KEYINPUT59), .Z(new_n990));
  OAI211_X1 g804(.A(new_n635), .B(new_n630), .C1(new_n893), .C2(new_n990), .ZN(new_n991));
  INV_X1    g805(.A(new_n990), .ZN(new_n992));
  NAND3_X1  g806(.A1(new_n977), .A2(new_n636), .A3(new_n992), .ZN(new_n993));
  AND3_X1   g807(.A1(new_n991), .A2(new_n961), .A3(new_n993), .ZN(G63));
  INV_X1    g808(.A(new_n247), .ZN(new_n995));
  XNOR2_X1  g809(.A(KEYINPUT121), .B(KEYINPUT60), .ZN(new_n996));
  NAND2_X1  g810(.A1(G217), .A2(G902), .ZN(new_n997));
  XNOR2_X1  g811(.A(new_n996), .B(new_n997), .ZN(new_n998));
  OAI21_X1  g812(.A(new_n995), .B1(new_n887), .B2(new_n998), .ZN(new_n999));
  OR2_X1    g813(.A1(new_n887), .A2(new_n998), .ZN(new_n1000));
  INV_X1    g814(.A(new_n673), .ZN(new_n1001));
  OAI211_X1 g815(.A(new_n961), .B(new_n999), .C1(new_n1000), .C2(new_n1001), .ZN(new_n1002));
  INV_X1    g816(.A(KEYINPUT120), .ZN(new_n1003));
  AND3_X1   g817(.A1(new_n1002), .A2(new_n1003), .A3(KEYINPUT61), .ZN(new_n1004));
  AOI21_X1  g818(.A(KEYINPUT61), .B1(new_n1002), .B2(new_n1003), .ZN(new_n1005));
  NOR2_X1   g819(.A1(new_n1004), .A2(new_n1005), .ZN(G66));
  INV_X1    g820(.A(G224), .ZN(new_n1007));
  OAI21_X1  g821(.A(G953), .B1(new_n568), .B2(new_n1007), .ZN(new_n1008));
  NOR2_X1   g822(.A1(new_n837), .A2(new_n881), .ZN(new_n1009));
  OAI21_X1  g823(.A(new_n1008), .B1(new_n1009), .B2(G953), .ZN(new_n1010));
  OAI21_X1  g824(.A(new_n945), .B1(G898), .B2(new_n192), .ZN(new_n1011));
  XNOR2_X1  g825(.A(new_n1010), .B(new_n1011), .ZN(G69));
  AOI21_X1  g826(.A(new_n192), .B1(G227), .B2(G900), .ZN(new_n1013));
  NOR3_X1   g827(.A1(new_n801), .A2(new_n871), .A3(new_n922), .ZN(new_n1014));
  NAND2_X1  g828(.A1(new_n787), .A2(new_n822), .ZN(new_n1015));
  NOR3_X1   g829(.A1(new_n816), .A2(new_n1014), .A3(new_n1015), .ZN(new_n1016));
  NAND2_X1  g830(.A1(new_n849), .A2(new_n710), .ZN(new_n1017));
  INV_X1    g831(.A(new_n1017), .ZN(new_n1018));
  OAI21_X1  g832(.A(new_n1018), .B1(new_n801), .B2(new_n809), .ZN(new_n1019));
  INV_X1    g833(.A(KEYINPUT125), .ZN(new_n1020));
  XNOR2_X1  g834(.A(new_n1019), .B(new_n1020), .ZN(new_n1021));
  NAND3_X1  g835(.A1(new_n1016), .A2(new_n192), .A3(new_n1021), .ZN(new_n1022));
  OAI21_X1  g836(.A(new_n324), .B1(new_n329), .B2(new_n306), .ZN(new_n1023));
  XNOR2_X1  g837(.A(new_n1023), .B(new_n551), .ZN(new_n1024));
  NAND2_X1  g838(.A1(G900), .A2(G953), .ZN(new_n1025));
  NAND3_X1  g839(.A1(new_n1022), .A2(new_n1024), .A3(new_n1025), .ZN(new_n1026));
  AOI21_X1  g840(.A(new_n1013), .B1(new_n1026), .B2(KEYINPUT124), .ZN(new_n1027));
  INV_X1    g841(.A(KEYINPUT62), .ZN(new_n1028));
  AOI21_X1  g842(.A(new_n1028), .B1(new_n733), .B2(new_n1018), .ZN(new_n1029));
  NAND3_X1  g843(.A1(new_n819), .A2(new_n368), .A3(new_n776), .ZN(new_n1030));
  NOR2_X1   g844(.A1(new_n714), .A2(new_n1030), .ZN(new_n1031));
  XNOR2_X1  g845(.A(new_n1031), .B(KEYINPUT123), .ZN(new_n1032));
  NOR4_X1   g846(.A1(new_n816), .A2(new_n1029), .A3(new_n810), .A4(new_n1032), .ZN(new_n1033));
  NAND3_X1  g847(.A1(new_n733), .A2(new_n1028), .A3(new_n1018), .ZN(new_n1034));
  XNOR2_X1  g848(.A(new_n1034), .B(KEYINPUT122), .ZN(new_n1035));
  AOI21_X1  g849(.A(G953), .B1(new_n1033), .B2(new_n1035), .ZN(new_n1036));
  OAI21_X1  g850(.A(new_n1026), .B1(new_n1036), .B2(new_n1024), .ZN(new_n1037));
  AND2_X1   g851(.A1(new_n1027), .A2(new_n1037), .ZN(new_n1038));
  NOR2_X1   g852(.A1(new_n1027), .A2(new_n1037), .ZN(new_n1039));
  NOR2_X1   g853(.A1(new_n1038), .A2(new_n1039), .ZN(G72));
  NAND3_X1  g854(.A1(new_n1016), .A2(new_n1009), .A3(new_n1021), .ZN(new_n1041));
  XNOR2_X1  g855(.A(KEYINPUT126), .B(KEYINPUT63), .ZN(new_n1042));
  NOR2_X1   g856(.A1(new_n646), .A2(new_n373), .ZN(new_n1043));
  XNOR2_X1  g857(.A(new_n1042), .B(new_n1043), .ZN(new_n1044));
  NAND2_X1  g858(.A1(new_n1041), .A2(new_n1044), .ZN(new_n1045));
  INV_X1    g859(.A(new_n363), .ZN(new_n1046));
  NAND3_X1  g860(.A1(new_n1045), .A2(new_n331), .A3(new_n1046), .ZN(new_n1047));
  NAND2_X1  g861(.A1(new_n364), .A2(new_n724), .ZN(new_n1048));
  NAND3_X1  g862(.A1(new_n891), .A2(new_n1044), .A3(new_n1048), .ZN(new_n1049));
  NAND3_X1  g863(.A1(new_n1047), .A2(new_n961), .A3(new_n1049), .ZN(new_n1050));
  NAND3_X1  g864(.A1(new_n1033), .A2(new_n1009), .A3(new_n1035), .ZN(new_n1051));
  NAND2_X1  g865(.A1(new_n1051), .A2(new_n1044), .ZN(new_n1052));
  NOR2_X1   g866(.A1(new_n1046), .A2(new_n331), .ZN(new_n1053));
  NAND2_X1  g867(.A1(new_n1052), .A2(new_n1053), .ZN(new_n1054));
  NAND2_X1  g868(.A1(new_n1054), .A2(KEYINPUT127), .ZN(new_n1055));
  INV_X1    g869(.A(KEYINPUT127), .ZN(new_n1056));
  NAND3_X1  g870(.A1(new_n1052), .A2(new_n1056), .A3(new_n1053), .ZN(new_n1057));
  AOI21_X1  g871(.A(new_n1050), .B1(new_n1055), .B2(new_n1057), .ZN(G57));
endmodule


