//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 0 0 0 1 1 0 1 0 0 1 0 1 0 1 0 1 1 0 1 0 1 0 1 1 1 1 1 0 1 0 0 1 1 1 1 0 0 1 0 1 1 0 0 0 1 1 0 1 1 1 0 0 0 0 0 0 1 0 1 0 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:39:24 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n236, new_n237,
    new_n238, new_n240, new_n241, new_n242, new_n243, new_n244, new_n245,
    new_n246, new_n248, new_n249, new_n250, new_n251, new_n252, new_n253,
    new_n254, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n822, new_n823, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1192, new_n1193,
    new_n1194, new_n1195, new_n1196, new_n1197, new_n1198, new_n1199,
    new_n1200, new_n1201, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1214, new_n1215, new_n1216, new_n1217, new_n1218,
    new_n1219, new_n1220, new_n1221, new_n1222, new_n1224, new_n1225,
    new_n1226, new_n1227, new_n1228, new_n1229, new_n1230, new_n1231,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1293,
    new_n1294, new_n1295, new_n1296, new_n1297, new_n1298, new_n1299,
    new_n1300, new_n1301, new_n1302, new_n1303, new_n1304, new_n1305,
    new_n1306, new_n1307, new_n1308, new_n1309, new_n1310, new_n1311,
    new_n1312, new_n1313;
  INV_X1    g0000(.A(KEYINPUT64), .ZN(new_n201));
  INV_X1    g0001(.A(G58), .ZN(new_n202));
  INV_X1    g0002(.A(G68), .ZN(new_n203));
  NAND3_X1  g0003(.A1(new_n201), .A2(new_n202), .A3(new_n203), .ZN(new_n204));
  OAI21_X1  g0004(.A(KEYINPUT64), .B1(G58), .B2(G68), .ZN(new_n205));
  NAND2_X1  g0005(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  INV_X1    g0006(.A(new_n206), .ZN(new_n207));
  NOR3_X1   g0007(.A1(new_n207), .A2(G50), .A3(G77), .ZN(G353));
  OAI21_X1  g0008(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0009(.A1(G1), .A2(G20), .ZN(new_n210));
  INV_X1    g0010(.A(G238), .ZN(new_n211));
  NOR2_X1   g0011(.A1(new_n203), .A2(new_n211), .ZN(new_n212));
  NAND2_X1  g0012(.A1(G97), .A2(G257), .ZN(new_n213));
  INV_X1    g0013(.A(G87), .ZN(new_n214));
  INV_X1    g0014(.A(G250), .ZN(new_n215));
  OAI21_X1  g0015(.A(new_n213), .B1(new_n214), .B2(new_n215), .ZN(new_n216));
  AOI211_X1 g0016(.A(new_n212), .B(new_n216), .C1(G107), .C2(G264), .ZN(new_n217));
  NAND2_X1  g0017(.A1(G116), .A2(G270), .ZN(new_n218));
  AND2_X1   g0018(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  INV_X1    g0019(.A(G50), .ZN(new_n220));
  INV_X1    g0020(.A(G226), .ZN(new_n221));
  INV_X1    g0021(.A(G77), .ZN(new_n222));
  INV_X1    g0022(.A(G244), .ZN(new_n223));
  OAI221_X1 g0023(.A(new_n219), .B1(new_n220), .B2(new_n221), .C1(new_n222), .C2(new_n223), .ZN(new_n224));
  INV_X1    g0024(.A(G232), .ZN(new_n225));
  NOR2_X1   g0025(.A1(new_n202), .A2(new_n225), .ZN(new_n226));
  OAI21_X1  g0026(.A(new_n210), .B1(new_n224), .B2(new_n226), .ZN(new_n227));
  XNOR2_X1  g0027(.A(new_n227), .B(KEYINPUT1), .ZN(new_n228));
  NOR2_X1   g0028(.A1(new_n206), .A2(new_n220), .ZN(new_n229));
  NAND2_X1  g0029(.A1(G1), .A2(G13), .ZN(new_n230));
  INV_X1    g0030(.A(G20), .ZN(new_n231));
  NOR2_X1   g0031(.A1(new_n230), .A2(new_n231), .ZN(new_n232));
  NOR2_X1   g0032(.A1(new_n210), .A2(G13), .ZN(new_n233));
  OAI211_X1 g0033(.A(new_n233), .B(G250), .C1(G257), .C2(G264), .ZN(new_n234));
  INV_X1    g0034(.A(KEYINPUT0), .ZN(new_n235));
  AOI22_X1  g0035(.A1(new_n229), .A2(new_n232), .B1(new_n234), .B2(new_n235), .ZN(new_n236));
  OAI21_X1  g0036(.A(new_n236), .B1(new_n235), .B2(new_n234), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n237), .B(KEYINPUT65), .ZN(new_n238));
  NOR2_X1   g0038(.A1(new_n228), .A2(new_n238), .ZN(G361));
  XNOR2_X1  g0039(.A(G250), .B(G257), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n240), .B(G264), .ZN(new_n241));
  XOR2_X1   g0041(.A(new_n241), .B(G270), .Z(new_n242));
  XNOR2_X1  g0042(.A(KEYINPUT2), .B(G226), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n243), .B(new_n225), .ZN(new_n244));
  XNOR2_X1  g0044(.A(G238), .B(G244), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XOR2_X1   g0046(.A(new_n242), .B(new_n246), .Z(G358));
  XNOR2_X1  g0047(.A(G50), .B(G58), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n248), .B(KEYINPUT66), .ZN(new_n249));
  XNOR2_X1  g0049(.A(G68), .B(G77), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n249), .B(new_n250), .ZN(new_n251));
  XOR2_X1   g0051(.A(G107), .B(G116), .Z(new_n252));
  XNOR2_X1  g0052(.A(G87), .B(G97), .ZN(new_n253));
  XNOR2_X1  g0053(.A(new_n252), .B(new_n253), .ZN(new_n254));
  XNOR2_X1  g0054(.A(new_n251), .B(new_n254), .ZN(G351));
  NAND3_X1  g0055(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n256));
  AND2_X1   g0056(.A1(new_n256), .A2(new_n230), .ZN(new_n257));
  OAI21_X1  g0057(.A(G20), .B1(new_n207), .B2(G50), .ZN(new_n258));
  XOR2_X1   g0058(.A(KEYINPUT8), .B(G58), .Z(new_n259));
  INV_X1    g0059(.A(G33), .ZN(new_n260));
  NOR2_X1   g0060(.A1(new_n260), .A2(G20), .ZN(new_n261));
  NOR2_X1   g0061(.A1(G20), .A2(G33), .ZN(new_n262));
  AOI22_X1  g0062(.A1(new_n259), .A2(new_n261), .B1(G150), .B2(new_n262), .ZN(new_n263));
  AOI21_X1  g0063(.A(new_n257), .B1(new_n258), .B2(new_n263), .ZN(new_n264));
  INV_X1    g0064(.A(G1), .ZN(new_n265));
  NAND3_X1  g0065(.A1(new_n265), .A2(G13), .A3(G20), .ZN(new_n266));
  INV_X1    g0066(.A(new_n266), .ZN(new_n267));
  AOI21_X1  g0067(.A(new_n264), .B1(new_n220), .B2(new_n267), .ZN(new_n268));
  OAI21_X1  g0068(.A(new_n257), .B1(G1), .B2(new_n231), .ZN(new_n269));
  INV_X1    g0069(.A(new_n269), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n270), .A2(G50), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n268), .A2(new_n271), .ZN(new_n272));
  XNOR2_X1  g0072(.A(new_n272), .B(KEYINPUT9), .ZN(new_n273));
  NAND2_X1  g0073(.A1(G33), .A2(G41), .ZN(new_n274));
  NAND3_X1  g0074(.A1(new_n274), .A2(G1), .A3(G13), .ZN(new_n275));
  INV_X1    g0075(.A(new_n275), .ZN(new_n276));
  AND2_X1   g0076(.A1(KEYINPUT3), .A2(G33), .ZN(new_n277));
  NOR2_X1   g0077(.A1(KEYINPUT3), .A2(G33), .ZN(new_n278));
  NOR2_X1   g0078(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  NOR2_X1   g0079(.A1(new_n279), .A2(G1698), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n280), .A2(G222), .ZN(new_n281));
  XNOR2_X1  g0081(.A(new_n281), .B(KEYINPUT67), .ZN(new_n282));
  INV_X1    g0082(.A(KEYINPUT3), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n283), .A2(new_n260), .ZN(new_n284));
  NAND2_X1  g0084(.A1(KEYINPUT3), .A2(G33), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n286), .A2(G1698), .ZN(new_n287));
  INV_X1    g0087(.A(G223), .ZN(new_n288));
  OAI22_X1  g0088(.A1(new_n287), .A2(new_n288), .B1(new_n222), .B2(new_n286), .ZN(new_n289));
  OAI21_X1  g0089(.A(new_n276), .B1(new_n282), .B2(new_n289), .ZN(new_n290));
  OAI21_X1  g0090(.A(new_n265), .B1(G41), .B2(G45), .ZN(new_n291));
  INV_X1    g0091(.A(G274), .ZN(new_n292));
  NOR2_X1   g0092(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  INV_X1    g0093(.A(new_n293), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n275), .A2(new_n291), .ZN(new_n295));
  INV_X1    g0095(.A(new_n295), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n296), .A2(G226), .ZN(new_n297));
  AND3_X1   g0097(.A1(new_n290), .A2(new_n294), .A3(new_n297), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n298), .A2(G190), .ZN(new_n299));
  INV_X1    g0099(.A(G200), .ZN(new_n300));
  OAI211_X1 g0100(.A(new_n273), .B(new_n299), .C1(new_n300), .C2(new_n298), .ZN(new_n301));
  INV_X1    g0101(.A(new_n301), .ZN(new_n302));
  INV_X1    g0102(.A(KEYINPUT69), .ZN(new_n303));
  NAND3_X1  g0103(.A1(new_n273), .A2(new_n299), .A3(new_n303), .ZN(new_n304));
  INV_X1    g0104(.A(KEYINPUT10), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n302), .A2(new_n306), .ZN(new_n307));
  NAND3_X1  g0107(.A1(new_n301), .A2(new_n304), .A3(new_n305), .ZN(new_n308));
  INV_X1    g0108(.A(G179), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n298), .A2(new_n309), .ZN(new_n310));
  OAI211_X1 g0110(.A(new_n310), .B(new_n272), .C1(G169), .C2(new_n298), .ZN(new_n311));
  NAND3_X1  g0111(.A1(new_n307), .A2(new_n308), .A3(new_n311), .ZN(new_n312));
  INV_X1    g0112(.A(G1698), .ZN(new_n313));
  NAND3_X1  g0113(.A1(new_n286), .A2(G226), .A3(new_n313), .ZN(new_n314));
  NAND2_X1  g0114(.A1(G33), .A2(G97), .ZN(new_n315));
  OAI211_X1 g0115(.A(new_n314), .B(new_n315), .C1(new_n287), .C2(new_n225), .ZN(new_n316));
  AOI21_X1  g0116(.A(new_n293), .B1(new_n316), .B2(new_n276), .ZN(new_n317));
  INV_X1    g0117(.A(KEYINPUT13), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n296), .A2(G238), .ZN(new_n319));
  AND3_X1   g0119(.A1(new_n317), .A2(new_n318), .A3(new_n319), .ZN(new_n320));
  AOI21_X1  g0120(.A(new_n318), .B1(new_n317), .B2(new_n319), .ZN(new_n321));
  NOR2_X1   g0121(.A1(new_n320), .A2(new_n321), .ZN(new_n322));
  INV_X1    g0122(.A(new_n322), .ZN(new_n323));
  INV_X1    g0123(.A(KEYINPUT73), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n324), .A2(KEYINPUT14), .ZN(new_n325));
  NAND3_X1  g0125(.A1(new_n323), .A2(G169), .A3(new_n325), .ZN(new_n326));
  INV_X1    g0126(.A(G169), .ZN(new_n327));
  OAI211_X1 g0127(.A(new_n324), .B(KEYINPUT14), .C1(new_n322), .C2(new_n327), .ZN(new_n328));
  NOR2_X1   g0128(.A1(new_n324), .A2(KEYINPUT14), .ZN(new_n329));
  AOI21_X1  g0129(.A(new_n329), .B1(new_n322), .B2(G179), .ZN(new_n330));
  NAND3_X1  g0130(.A1(new_n326), .A2(new_n328), .A3(new_n330), .ZN(new_n331));
  AOI22_X1  g0131(.A1(new_n261), .A2(G77), .B1(G20), .B2(new_n203), .ZN(new_n332));
  XNOR2_X1  g0132(.A(new_n332), .B(KEYINPUT70), .ZN(new_n333));
  INV_X1    g0133(.A(new_n262), .ZN(new_n334));
  OAI21_X1  g0134(.A(new_n333), .B1(new_n220), .B2(new_n334), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n256), .A2(new_n230), .ZN(new_n336));
  XOR2_X1   g0136(.A(KEYINPUT71), .B(KEYINPUT11), .Z(new_n337));
  AND3_X1   g0137(.A1(new_n335), .A2(new_n336), .A3(new_n337), .ZN(new_n338));
  INV_X1    g0138(.A(G13), .ZN(new_n339));
  NOR2_X1   g0139(.A1(new_n339), .A2(G1), .ZN(new_n340));
  NAND3_X1  g0140(.A1(new_n340), .A2(G20), .A3(new_n203), .ZN(new_n341));
  INV_X1    g0141(.A(KEYINPUT12), .ZN(new_n342));
  OR2_X1    g0142(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n341), .A2(new_n342), .ZN(new_n344));
  OAI211_X1 g0144(.A(new_n343), .B(new_n344), .C1(new_n203), .C2(new_n269), .ZN(new_n345));
  XNOR2_X1  g0145(.A(new_n345), .B(KEYINPUT72), .ZN(new_n346));
  AOI21_X1  g0146(.A(new_n337), .B1(new_n335), .B2(new_n336), .ZN(new_n347));
  NOR3_X1   g0147(.A1(new_n338), .A2(new_n346), .A3(new_n347), .ZN(new_n348));
  INV_X1    g0148(.A(new_n348), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n323), .A2(G200), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n322), .A2(G190), .ZN(new_n351));
  AND2_X1   g0151(.A1(new_n351), .A2(new_n348), .ZN(new_n352));
  AOI22_X1  g0152(.A1(new_n331), .A2(new_n349), .B1(new_n350), .B2(new_n352), .ZN(new_n353));
  AOI22_X1  g0153(.A1(new_n280), .A2(G232), .B1(G107), .B2(new_n279), .ZN(new_n354));
  OAI21_X1  g0154(.A(new_n354), .B1(new_n211), .B2(new_n287), .ZN(new_n355));
  AOI21_X1  g0155(.A(new_n293), .B1(new_n355), .B2(new_n276), .ZN(new_n356));
  OAI21_X1  g0156(.A(new_n356), .B1(new_n223), .B2(new_n295), .ZN(new_n357));
  NOR2_X1   g0157(.A1(new_n357), .A2(G179), .ZN(new_n358));
  AOI21_X1  g0158(.A(new_n358), .B1(new_n327), .B2(new_n357), .ZN(new_n359));
  OR2_X1    g0159(.A1(KEYINPUT15), .A2(G87), .ZN(new_n360));
  NAND2_X1  g0160(.A1(KEYINPUT15), .A2(G87), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  INV_X1    g0162(.A(new_n362), .ZN(new_n363));
  AOI22_X1  g0163(.A1(new_n363), .A2(new_n261), .B1(G20), .B2(G77), .ZN(new_n364));
  XNOR2_X1  g0164(.A(new_n259), .B(KEYINPUT68), .ZN(new_n365));
  OAI21_X1  g0165(.A(new_n364), .B1(new_n365), .B2(new_n334), .ZN(new_n366));
  AOI22_X1  g0166(.A1(new_n366), .A2(new_n336), .B1(new_n222), .B2(new_n267), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n270), .A2(G77), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n359), .A2(new_n369), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n353), .A2(new_n370), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n221), .A2(G1698), .ZN(new_n372));
  OAI221_X1 g0172(.A(new_n372), .B1(G223), .B2(G1698), .C1(new_n277), .C2(new_n278), .ZN(new_n373));
  NAND2_X1  g0173(.A1(G33), .A2(G87), .ZN(new_n374));
  AOI21_X1  g0174(.A(new_n275), .B1(new_n373), .B2(new_n374), .ZN(new_n375));
  NOR2_X1   g0175(.A1(new_n295), .A2(new_n225), .ZN(new_n376));
  OR3_X1    g0176(.A1(new_n375), .A2(new_n293), .A3(new_n376), .ZN(new_n377));
  OAI21_X1  g0177(.A(KEYINPUT76), .B1(new_n377), .B2(G190), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n377), .A2(new_n300), .ZN(new_n379));
  NOR3_X1   g0179(.A1(new_n375), .A2(new_n376), .A3(new_n293), .ZN(new_n380));
  INV_X1    g0180(.A(KEYINPUT76), .ZN(new_n381));
  INV_X1    g0181(.A(G190), .ZN(new_n382));
  NAND3_X1  g0182(.A1(new_n380), .A2(new_n381), .A3(new_n382), .ZN(new_n383));
  NAND3_X1  g0183(.A1(new_n378), .A2(new_n379), .A3(new_n383), .ZN(new_n384));
  NAND3_X1  g0184(.A1(new_n284), .A2(new_n231), .A3(new_n285), .ZN(new_n385));
  INV_X1    g0185(.A(KEYINPUT7), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n385), .A2(new_n386), .ZN(new_n387));
  INV_X1    g0187(.A(KEYINPUT74), .ZN(new_n388));
  NAND4_X1  g0188(.A1(new_n284), .A2(KEYINPUT7), .A3(new_n231), .A4(new_n285), .ZN(new_n389));
  NAND3_X1  g0189(.A1(new_n387), .A2(new_n388), .A3(new_n389), .ZN(new_n390));
  OAI211_X1 g0190(.A(new_n390), .B(G68), .C1(new_n388), .C2(new_n389), .ZN(new_n391));
  NOR2_X1   g0191(.A1(new_n202), .A2(new_n203), .ZN(new_n392));
  OAI21_X1  g0192(.A(G20), .B1(new_n206), .B2(new_n392), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n262), .A2(G159), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n393), .A2(new_n394), .ZN(new_n395));
  INV_X1    g0195(.A(new_n395), .ZN(new_n396));
  NAND3_X1  g0196(.A1(new_n391), .A2(KEYINPUT16), .A3(new_n396), .ZN(new_n397));
  INV_X1    g0197(.A(KEYINPUT16), .ZN(new_n398));
  AOI21_X1  g0198(.A(new_n203), .B1(new_n387), .B2(new_n389), .ZN(new_n399));
  OAI21_X1  g0199(.A(new_n398), .B1(new_n395), .B2(new_n399), .ZN(new_n400));
  NAND3_X1  g0200(.A1(new_n397), .A2(new_n336), .A3(new_n400), .ZN(new_n401));
  NOR2_X1   g0201(.A1(new_n259), .A2(new_n267), .ZN(new_n402));
  AOI21_X1  g0202(.A(new_n402), .B1(new_n269), .B2(new_n259), .ZN(new_n403));
  INV_X1    g0203(.A(new_n403), .ZN(new_n404));
  NAND3_X1  g0204(.A1(new_n384), .A2(new_n401), .A3(new_n404), .ZN(new_n405));
  INV_X1    g0205(.A(KEYINPUT17), .ZN(new_n406));
  XNOR2_X1  g0206(.A(new_n405), .B(new_n406), .ZN(new_n407));
  INV_X1    g0207(.A(new_n407), .ZN(new_n408));
  NAND3_X1  g0208(.A1(new_n380), .A2(KEYINPUT75), .A3(new_n309), .ZN(new_n409));
  INV_X1    g0209(.A(new_n409), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n380), .A2(new_n309), .ZN(new_n411));
  OAI21_X1  g0211(.A(KEYINPUT75), .B1(new_n380), .B2(G169), .ZN(new_n412));
  AOI21_X1  g0212(.A(new_n410), .B1(new_n411), .B2(new_n412), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n401), .A2(new_n404), .ZN(new_n414));
  AND3_X1   g0214(.A1(new_n413), .A2(KEYINPUT18), .A3(new_n414), .ZN(new_n415));
  AOI21_X1  g0215(.A(KEYINPUT18), .B1(new_n413), .B2(new_n414), .ZN(new_n416));
  NOR2_X1   g0216(.A1(new_n415), .A2(new_n416), .ZN(new_n417));
  INV_X1    g0217(.A(new_n417), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n408), .A2(new_n418), .ZN(new_n419));
  INV_X1    g0219(.A(new_n369), .ZN(new_n420));
  OAI21_X1  g0220(.A(new_n420), .B1(new_n382), .B2(new_n357), .ZN(new_n421));
  AND2_X1   g0221(.A1(new_n357), .A2(G200), .ZN(new_n422));
  OR2_X1    g0222(.A1(new_n421), .A2(new_n422), .ZN(new_n423));
  INV_X1    g0223(.A(new_n423), .ZN(new_n424));
  NOR4_X1   g0224(.A1(new_n312), .A2(new_n371), .A3(new_n419), .A4(new_n424), .ZN(new_n425));
  INV_X1    g0225(.A(G45), .ZN(new_n426));
  NOR2_X1   g0226(.A1(new_n426), .A2(G1), .ZN(new_n427));
  AND2_X1   g0227(.A1(KEYINPUT5), .A2(G41), .ZN(new_n428));
  NOR2_X1   g0228(.A1(KEYINPUT5), .A2(G41), .ZN(new_n429));
  OAI21_X1  g0229(.A(new_n427), .B1(new_n428), .B2(new_n429), .ZN(new_n430));
  AND3_X1   g0230(.A1(new_n430), .A2(G257), .A3(new_n275), .ZN(new_n431));
  OAI21_X1  g0231(.A(G244), .B1(new_n277), .B2(new_n278), .ZN(new_n432));
  INV_X1    g0232(.A(KEYINPUT4), .ZN(new_n433));
  AOI22_X1  g0233(.A1(new_n432), .A2(new_n433), .B1(G33), .B2(G283), .ZN(new_n434));
  NAND4_X1  g0234(.A1(new_n286), .A2(KEYINPUT4), .A3(G244), .A4(new_n313), .ZN(new_n435));
  AOI21_X1  g0235(.A(new_n433), .B1(new_n286), .B2(G250), .ZN(new_n436));
  OAI211_X1 g0236(.A(new_n434), .B(new_n435), .C1(new_n313), .C2(new_n436), .ZN(new_n437));
  AOI21_X1  g0237(.A(new_n431), .B1(new_n437), .B2(new_n276), .ZN(new_n438));
  OAI211_X1 g0238(.A(new_n427), .B(G274), .C1(new_n429), .C2(new_n428), .ZN(new_n439));
  NAND3_X1  g0239(.A1(new_n438), .A2(G190), .A3(new_n439), .ZN(new_n440));
  INV_X1    g0240(.A(new_n439), .ZN(new_n441));
  AOI211_X1 g0241(.A(new_n441), .B(new_n431), .C1(new_n437), .C2(new_n276), .ZN(new_n442));
  OAI21_X1  g0242(.A(new_n440), .B1(new_n300), .B2(new_n442), .ZN(new_n443));
  NOR2_X1   g0243(.A1(new_n266), .A2(G97), .ZN(new_n444));
  INV_X1    g0244(.A(new_n444), .ZN(new_n445));
  OAI211_X1 g0245(.A(new_n257), .B(new_n266), .C1(G1), .C2(new_n260), .ZN(new_n446));
  INV_X1    g0246(.A(G97), .ZN(new_n447));
  NOR2_X1   g0247(.A1(new_n446), .A2(new_n447), .ZN(new_n448));
  INV_X1    g0248(.A(new_n448), .ZN(new_n449));
  INV_X1    g0249(.A(KEYINPUT77), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n387), .A2(new_n389), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n451), .A2(G107), .ZN(new_n452));
  INV_X1    g0252(.A(KEYINPUT6), .ZN(new_n453));
  AND2_X1   g0253(.A1(G97), .A2(G107), .ZN(new_n454));
  NOR2_X1   g0254(.A1(G97), .A2(G107), .ZN(new_n455));
  OAI21_X1  g0255(.A(new_n453), .B1(new_n454), .B2(new_n455), .ZN(new_n456));
  INV_X1    g0256(.A(G107), .ZN(new_n457));
  NAND3_X1  g0257(.A1(new_n457), .A2(KEYINPUT6), .A3(G97), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n456), .A2(new_n458), .ZN(new_n459));
  AOI22_X1  g0259(.A1(new_n459), .A2(G20), .B1(G77), .B2(new_n262), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n452), .A2(new_n460), .ZN(new_n461));
  AOI21_X1  g0261(.A(new_n450), .B1(new_n461), .B2(new_n336), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n262), .A2(G77), .ZN(new_n463));
  AND3_X1   g0263(.A1(new_n457), .A2(KEYINPUT6), .A3(G97), .ZN(new_n464));
  XNOR2_X1  g0264(.A(G97), .B(G107), .ZN(new_n465));
  AOI21_X1  g0265(.A(new_n464), .B1(new_n465), .B2(new_n453), .ZN(new_n466));
  OAI21_X1  g0266(.A(new_n463), .B1(new_n466), .B2(new_n231), .ZN(new_n467));
  AOI21_X1  g0267(.A(new_n457), .B1(new_n387), .B2(new_n389), .ZN(new_n468));
  OAI211_X1 g0268(.A(new_n450), .B(new_n336), .C1(new_n467), .C2(new_n468), .ZN(new_n469));
  INV_X1    g0269(.A(new_n469), .ZN(new_n470));
  OAI211_X1 g0270(.A(new_n445), .B(new_n449), .C1(new_n462), .C2(new_n470), .ZN(new_n471));
  NOR2_X1   g0271(.A1(new_n443), .A2(new_n471), .ZN(new_n472));
  OAI21_X1  g0272(.A(KEYINPUT23), .B1(new_n231), .B2(G107), .ZN(new_n473));
  INV_X1    g0273(.A(KEYINPUT23), .ZN(new_n474));
  NAND3_X1  g0274(.A1(new_n474), .A2(new_n457), .A3(G20), .ZN(new_n475));
  NAND3_X1  g0275(.A1(new_n231), .A2(G33), .A3(G116), .ZN(new_n476));
  NAND3_X1  g0276(.A1(new_n473), .A2(new_n475), .A3(new_n476), .ZN(new_n477));
  INV_X1    g0277(.A(KEYINPUT84), .ZN(new_n478));
  XNOR2_X1  g0278(.A(new_n477), .B(new_n478), .ZN(new_n479));
  OAI211_X1 g0279(.A(new_n231), .B(G87), .C1(new_n277), .C2(new_n278), .ZN(new_n480));
  XNOR2_X1  g0280(.A(new_n480), .B(KEYINPUT22), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n479), .A2(new_n481), .ZN(new_n482));
  INV_X1    g0282(.A(KEYINPUT24), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  NAND3_X1  g0284(.A1(new_n479), .A2(new_n481), .A3(KEYINPUT24), .ZN(new_n485));
  NAND3_X1  g0285(.A1(new_n484), .A2(new_n336), .A3(new_n485), .ZN(new_n486));
  NAND3_X1  g0286(.A1(new_n286), .A2(G257), .A3(G1698), .ZN(new_n487));
  INV_X1    g0287(.A(G294), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n286), .A2(new_n313), .ZN(new_n489));
  OAI221_X1 g0289(.A(new_n487), .B1(new_n260), .B2(new_n488), .C1(new_n489), .C2(new_n215), .ZN(new_n490));
  AND2_X1   g0290(.A1(new_n430), .A2(new_n275), .ZN(new_n491));
  AOI22_X1  g0291(.A1(new_n490), .A2(new_n276), .B1(G264), .B2(new_n491), .ZN(new_n492));
  NAND3_X1  g0292(.A1(new_n492), .A2(G190), .A3(new_n439), .ZN(new_n493));
  INV_X1    g0293(.A(new_n446), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n494), .A2(G107), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n267), .A2(new_n457), .ZN(new_n496));
  XNOR2_X1  g0296(.A(new_n496), .B(KEYINPUT85), .ZN(new_n497));
  XNOR2_X1  g0297(.A(new_n497), .B(KEYINPUT25), .ZN(new_n498));
  NAND4_X1  g0298(.A1(new_n486), .A2(new_n493), .A3(new_n495), .A4(new_n498), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n490), .A2(new_n276), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n491), .A2(G264), .ZN(new_n501));
  NAND3_X1  g0301(.A1(new_n500), .A2(new_n439), .A3(new_n501), .ZN(new_n502));
  INV_X1    g0302(.A(new_n502), .ZN(new_n503));
  NOR2_X1   g0303(.A1(new_n503), .A2(new_n300), .ZN(new_n504));
  NOR2_X1   g0304(.A1(new_n499), .A2(new_n504), .ZN(new_n505));
  INV_X1    g0305(.A(KEYINPUT78), .ZN(new_n506));
  OAI21_X1  g0306(.A(new_n336), .B1(new_n467), .B2(new_n468), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n507), .A2(KEYINPUT77), .ZN(new_n508));
  AOI211_X1 g0308(.A(new_n444), .B(new_n448), .C1(new_n508), .C2(new_n469), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n437), .A2(new_n276), .ZN(new_n510));
  INV_X1    g0310(.A(new_n431), .ZN(new_n511));
  NAND4_X1  g0311(.A1(new_n510), .A2(new_n309), .A3(new_n439), .A4(new_n511), .ZN(new_n512));
  OAI21_X1  g0312(.A(new_n512), .B1(new_n442), .B2(G169), .ZN(new_n513));
  OAI21_X1  g0313(.A(new_n506), .B1(new_n509), .B2(new_n513), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n438), .A2(new_n439), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n515), .A2(new_n327), .ZN(new_n516));
  NAND4_X1  g0316(.A1(new_n471), .A2(KEYINPUT78), .A3(new_n516), .A4(new_n512), .ZN(new_n517));
  AOI211_X1 g0317(.A(new_n472), .B(new_n505), .C1(new_n514), .C2(new_n517), .ZN(new_n518));
  NOR2_X1   g0318(.A1(new_n502), .A2(G179), .ZN(new_n519));
  AOI21_X1  g0319(.A(G169), .B1(new_n492), .B2(new_n439), .ZN(new_n520));
  NOR2_X1   g0320(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  NAND3_X1  g0321(.A1(new_n486), .A2(new_n495), .A3(new_n498), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  INV_X1    g0323(.A(KEYINPUT83), .ZN(new_n524));
  NOR2_X1   g0324(.A1(new_n266), .A2(G116), .ZN(new_n525));
  INV_X1    g0325(.A(G116), .ZN(new_n526));
  NOR2_X1   g0326(.A1(new_n446), .A2(new_n526), .ZN(new_n527));
  AOI21_X1  g0327(.A(G20), .B1(new_n260), .B2(G97), .ZN(new_n528));
  NAND2_X1  g0328(.A1(G33), .A2(G283), .ZN(new_n529));
  NAND3_X1  g0329(.A1(new_n528), .A2(KEYINPUT81), .A3(new_n529), .ZN(new_n530));
  AND2_X1   g0330(.A1(new_n530), .A2(new_n336), .ZN(new_n531));
  AOI21_X1  g0331(.A(KEYINPUT81), .B1(new_n528), .B2(new_n529), .ZN(new_n532));
  INV_X1    g0332(.A(new_n532), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n526), .A2(G20), .ZN(new_n534));
  NAND4_X1  g0334(.A1(new_n531), .A2(KEYINPUT20), .A3(new_n533), .A4(new_n534), .ZN(new_n535));
  INV_X1    g0335(.A(KEYINPUT20), .ZN(new_n536));
  NAND3_X1  g0336(.A1(new_n530), .A2(new_n336), .A3(new_n534), .ZN(new_n537));
  OAI21_X1  g0337(.A(new_n536), .B1(new_n537), .B2(new_n532), .ZN(new_n538));
  AOI211_X1 g0338(.A(new_n525), .B(new_n527), .C1(new_n535), .C2(new_n538), .ZN(new_n539));
  NOR2_X1   g0339(.A1(new_n279), .A2(new_n313), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n279), .A2(G303), .ZN(new_n541));
  INV_X1    g0341(.A(KEYINPUT80), .ZN(new_n542));
  AOI22_X1  g0342(.A1(G264), .A2(new_n540), .B1(new_n541), .B2(new_n542), .ZN(new_n543));
  NAND3_X1  g0343(.A1(new_n286), .A2(G264), .A3(G1698), .ZN(new_n544));
  INV_X1    g0344(.A(G257), .ZN(new_n545));
  OAI22_X1  g0345(.A1(new_n544), .A2(KEYINPUT80), .B1(new_n489), .B2(new_n545), .ZN(new_n546));
  OAI21_X1  g0346(.A(new_n276), .B1(new_n543), .B2(new_n546), .ZN(new_n547));
  AOI21_X1  g0347(.A(new_n441), .B1(new_n491), .B2(G270), .ZN(new_n548));
  NAND3_X1  g0348(.A1(new_n547), .A2(G190), .A3(new_n548), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n539), .A2(new_n549), .ZN(new_n550));
  AOI21_X1  g0350(.A(new_n300), .B1(new_n547), .B2(new_n548), .ZN(new_n551));
  OAI21_X1  g0351(.A(new_n524), .B1(new_n550), .B2(new_n551), .ZN(new_n552));
  INV_X1    g0352(.A(new_n551), .ZN(new_n553));
  NAND4_X1  g0353(.A1(new_n553), .A2(new_n539), .A3(KEYINPUT83), .A4(new_n549), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n552), .A2(new_n554), .ZN(new_n555));
  NAND3_X1  g0355(.A1(new_n214), .A2(new_n447), .A3(new_n457), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n315), .A2(new_n231), .ZN(new_n557));
  NAND3_X1  g0357(.A1(new_n556), .A2(new_n557), .A3(KEYINPUT19), .ZN(new_n558));
  OAI211_X1 g0358(.A(new_n231), .B(G68), .C1(new_n277), .C2(new_n278), .ZN(new_n559));
  INV_X1    g0359(.A(KEYINPUT19), .ZN(new_n560));
  OAI21_X1  g0360(.A(new_n560), .B1(new_n315), .B2(G20), .ZN(new_n561));
  NAND3_X1  g0361(.A1(new_n558), .A2(new_n559), .A3(new_n561), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n562), .A2(new_n336), .ZN(new_n563));
  AOI21_X1  g0363(.A(new_n266), .B1(new_n360), .B2(new_n361), .ZN(new_n564));
  INV_X1    g0364(.A(new_n564), .ZN(new_n565));
  AOI21_X1  g0365(.A(KEYINPUT79), .B1(new_n563), .B2(new_n565), .ZN(new_n566));
  INV_X1    g0366(.A(KEYINPUT79), .ZN(new_n567));
  AOI211_X1 g0367(.A(new_n567), .B(new_n564), .C1(new_n562), .C2(new_n336), .ZN(new_n568));
  OAI22_X1  g0368(.A1(new_n566), .A2(new_n568), .B1(new_n362), .B2(new_n446), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n211), .A2(new_n313), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n223), .A2(G1698), .ZN(new_n571));
  OAI211_X1 g0371(.A(new_n570), .B(new_n571), .C1(new_n277), .C2(new_n278), .ZN(new_n572));
  NAND2_X1  g0372(.A1(G33), .A2(G116), .ZN(new_n573));
  AOI21_X1  g0373(.A(new_n275), .B1(new_n572), .B2(new_n573), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n427), .A2(new_n292), .ZN(new_n575));
  OAI21_X1  g0375(.A(new_n215), .B1(new_n426), .B2(G1), .ZN(new_n576));
  AND3_X1   g0376(.A1(new_n575), .A2(new_n275), .A3(new_n576), .ZN(new_n577));
  NOR2_X1   g0377(.A1(new_n574), .A2(new_n577), .ZN(new_n578));
  INV_X1    g0378(.A(new_n578), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n579), .A2(new_n327), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n578), .A2(new_n309), .ZN(new_n581));
  NAND3_X1  g0381(.A1(new_n569), .A2(new_n580), .A3(new_n581), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n563), .A2(new_n565), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n583), .A2(new_n567), .ZN(new_n584));
  NAND3_X1  g0384(.A1(new_n563), .A2(KEYINPUT79), .A3(new_n565), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n578), .A2(G190), .ZN(new_n587));
  OAI21_X1  g0387(.A(G200), .B1(new_n574), .B2(new_n577), .ZN(new_n588));
  AND2_X1   g0388(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n494), .A2(G87), .ZN(new_n590));
  NAND3_X1  g0390(.A1(new_n586), .A2(new_n589), .A3(new_n590), .ZN(new_n591));
  AND2_X1   g0391(.A1(new_n582), .A2(new_n591), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n535), .A2(new_n538), .ZN(new_n593));
  INV_X1    g0393(.A(new_n527), .ZN(new_n594));
  INV_X1    g0394(.A(new_n525), .ZN(new_n595));
  NAND3_X1  g0395(.A1(new_n593), .A2(new_n594), .A3(new_n595), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n547), .A2(new_n548), .ZN(new_n597));
  NAND3_X1  g0397(.A1(new_n596), .A2(G169), .A3(new_n597), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n598), .A2(KEYINPUT21), .ZN(new_n599));
  INV_X1    g0399(.A(KEYINPUT21), .ZN(new_n600));
  NAND4_X1  g0400(.A1(new_n596), .A2(new_n597), .A3(new_n600), .A4(G169), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n599), .A2(new_n601), .ZN(new_n602));
  INV_X1    g0402(.A(new_n597), .ZN(new_n603));
  INV_X1    g0403(.A(KEYINPUT82), .ZN(new_n604));
  NAND4_X1  g0404(.A1(new_n603), .A2(new_n596), .A3(new_n604), .A4(G179), .ZN(new_n605));
  NAND3_X1  g0405(.A1(new_n547), .A2(G179), .A3(new_n548), .ZN(new_n606));
  OAI21_X1  g0406(.A(KEYINPUT82), .B1(new_n539), .B2(new_n606), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n605), .A2(new_n607), .ZN(new_n608));
  NAND4_X1  g0408(.A1(new_n555), .A2(new_n592), .A3(new_n602), .A4(new_n608), .ZN(new_n609));
  INV_X1    g0409(.A(new_n609), .ZN(new_n610));
  AND4_X1   g0410(.A1(new_n425), .A2(new_n518), .A3(new_n523), .A4(new_n610), .ZN(G372));
  NAND2_X1  g0411(.A1(new_n307), .A2(new_n308), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n352), .A2(new_n350), .ZN(new_n613));
  NAND3_X1  g0413(.A1(new_n371), .A2(new_n613), .A3(new_n408), .ZN(new_n614));
  AOI21_X1  g0414(.A(new_n612), .B1(new_n614), .B2(new_n418), .ZN(new_n615));
  INV_X1    g0415(.A(new_n311), .ZN(new_n616));
  NOR2_X1   g0416(.A1(new_n615), .A2(new_n616), .ZN(new_n617));
  INV_X1    g0417(.A(new_n589), .ZN(new_n618));
  OAI21_X1  g0418(.A(new_n590), .B1(new_n566), .B2(new_n568), .ZN(new_n619));
  INV_X1    g0419(.A(KEYINPUT86), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  OAI211_X1 g0421(.A(KEYINPUT86), .B(new_n590), .C1(new_n566), .C2(new_n568), .ZN(new_n622));
  AOI21_X1  g0422(.A(new_n618), .B1(new_n621), .B2(new_n622), .ZN(new_n623));
  AND3_X1   g0423(.A1(new_n569), .A2(new_n581), .A3(new_n580), .ZN(new_n624));
  NOR3_X1   g0424(.A1(new_n623), .A2(KEYINPUT87), .A3(new_n624), .ZN(new_n625));
  INV_X1    g0425(.A(new_n625), .ZN(new_n626));
  OAI21_X1  g0426(.A(KEYINPUT87), .B1(new_n623), .B2(new_n624), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n602), .A2(new_n608), .ZN(new_n629));
  INV_X1    g0429(.A(KEYINPUT88), .ZN(new_n630));
  XNOR2_X1  g0430(.A(new_n523), .B(new_n630), .ZN(new_n631));
  OAI211_X1 g0431(.A(new_n518), .B(new_n628), .C1(new_n629), .C2(new_n631), .ZN(new_n632));
  INV_X1    g0432(.A(KEYINPUT26), .ZN(new_n633));
  NOR2_X1   g0433(.A1(new_n509), .A2(new_n513), .ZN(new_n634));
  INV_X1    g0434(.A(KEYINPUT87), .ZN(new_n635));
  AOI21_X1  g0435(.A(KEYINPUT86), .B1(new_n586), .B2(new_n590), .ZN(new_n636));
  INV_X1    g0436(.A(new_n622), .ZN(new_n637));
  OAI21_X1  g0437(.A(new_n589), .B1(new_n636), .B2(new_n637), .ZN(new_n638));
  AOI21_X1  g0438(.A(new_n635), .B1(new_n638), .B2(new_n582), .ZN(new_n639));
  OAI211_X1 g0439(.A(new_n633), .B(new_n634), .C1(new_n639), .C2(new_n625), .ZN(new_n640));
  NAND3_X1  g0440(.A1(new_n514), .A2(new_n517), .A3(new_n592), .ZN(new_n641));
  AOI21_X1  g0441(.A(new_n624), .B1(new_n641), .B2(KEYINPUT26), .ZN(new_n642));
  AND3_X1   g0442(.A1(new_n640), .A2(new_n642), .A3(KEYINPUT89), .ZN(new_n643));
  AOI21_X1  g0443(.A(KEYINPUT89), .B1(new_n640), .B2(new_n642), .ZN(new_n644));
  OAI21_X1  g0444(.A(new_n632), .B1(new_n643), .B2(new_n644), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n425), .A2(new_n645), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n617), .A2(new_n646), .ZN(new_n647));
  XNOR2_X1  g0447(.A(new_n647), .B(KEYINPUT90), .ZN(G369));
  NAND2_X1  g0448(.A1(new_n340), .A2(new_n231), .ZN(new_n649));
  OR2_X1    g0449(.A1(new_n649), .A2(KEYINPUT27), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n649), .A2(KEYINPUT27), .ZN(new_n651));
  NAND3_X1  g0451(.A1(new_n650), .A2(new_n651), .A3(G213), .ZN(new_n652));
  INV_X1    g0452(.A(G343), .ZN(new_n653));
  NOR2_X1   g0453(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n596), .A2(new_n654), .ZN(new_n655));
  INV_X1    g0455(.A(new_n655), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n629), .A2(new_n656), .ZN(new_n657));
  NAND4_X1  g0457(.A1(new_n555), .A2(new_n608), .A3(new_n602), .A4(new_n655), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n659), .A2(G330), .ZN(new_n660));
  NAND3_X1  g0460(.A1(new_n521), .A2(new_n522), .A3(new_n654), .ZN(new_n661));
  AND3_X1   g0461(.A1(new_n486), .A2(new_n495), .A3(new_n498), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n502), .A2(new_n327), .ZN(new_n663));
  OAI21_X1  g0463(.A(new_n663), .B1(G179), .B2(new_n502), .ZN(new_n664));
  OAI22_X1  g0464(.A1(new_n662), .A2(new_n664), .B1(new_n499), .B2(new_n504), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n522), .A2(new_n654), .ZN(new_n666));
  INV_X1    g0466(.A(new_n666), .ZN(new_n667));
  OAI21_X1  g0467(.A(new_n661), .B1(new_n665), .B2(new_n667), .ZN(new_n668));
  INV_X1    g0468(.A(new_n668), .ZN(new_n669));
  NOR2_X1   g0469(.A1(new_n660), .A2(new_n669), .ZN(new_n670));
  INV_X1    g0470(.A(new_n670), .ZN(new_n671));
  INV_X1    g0471(.A(new_n654), .ZN(new_n672));
  INV_X1    g0472(.A(new_n665), .ZN(new_n673));
  AOI21_X1  g0473(.A(new_n654), .B1(new_n602), .B2(new_n608), .ZN(new_n674));
  AOI22_X1  g0474(.A1(new_n631), .A2(new_n672), .B1(new_n673), .B2(new_n674), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n671), .A2(new_n675), .ZN(G399));
  INV_X1    g0476(.A(new_n233), .ZN(new_n677));
  NOR2_X1   g0477(.A1(new_n677), .A2(G41), .ZN(new_n678));
  INV_X1    g0478(.A(new_n678), .ZN(new_n679));
  NOR2_X1   g0479(.A1(new_n556), .A2(G116), .ZN(new_n680));
  NAND3_X1  g0480(.A1(new_n679), .A2(G1), .A3(new_n680), .ZN(new_n681));
  INV_X1    g0481(.A(new_n229), .ZN(new_n682));
  OAI21_X1  g0482(.A(new_n681), .B1(new_n682), .B2(new_n679), .ZN(new_n683));
  XNOR2_X1  g0483(.A(new_n683), .B(KEYINPUT28), .ZN(new_n684));
  INV_X1    g0484(.A(KEYINPUT29), .ZN(new_n685));
  NAND3_X1  g0485(.A1(new_n602), .A2(new_n523), .A3(new_n608), .ZN(new_n686));
  NAND3_X1  g0486(.A1(new_n518), .A2(new_n628), .A3(new_n686), .ZN(new_n687));
  OAI21_X1  g0487(.A(new_n634), .B1(new_n639), .B2(new_n625), .ZN(new_n688));
  AOI21_X1  g0488(.A(new_n624), .B1(new_n688), .B2(KEYINPUT26), .ZN(new_n689));
  AND2_X1   g0489(.A1(new_n514), .A2(new_n517), .ZN(new_n690));
  NAND3_X1  g0490(.A1(new_n690), .A2(new_n633), .A3(new_n592), .ZN(new_n691));
  NAND3_X1  g0491(.A1(new_n687), .A2(new_n689), .A3(new_n691), .ZN(new_n692));
  AOI21_X1  g0492(.A(new_n685), .B1(new_n692), .B2(new_n672), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n640), .A2(new_n642), .ZN(new_n694));
  INV_X1    g0494(.A(KEYINPUT89), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  NAND3_X1  g0496(.A1(new_n640), .A2(new_n642), .A3(KEYINPUT89), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  AOI21_X1  g0498(.A(new_n654), .B1(new_n698), .B2(new_n632), .ZN(new_n699));
  AOI21_X1  g0499(.A(new_n693), .B1(new_n699), .B2(new_n685), .ZN(new_n700));
  NAND3_X1  g0500(.A1(new_n503), .A2(new_n438), .A3(new_n578), .ZN(new_n701));
  INV_X1    g0501(.A(KEYINPUT30), .ZN(new_n702));
  OR3_X1    g0502(.A1(new_n701), .A2(new_n702), .A3(new_n606), .ZN(new_n703));
  OAI21_X1  g0503(.A(new_n702), .B1(new_n701), .B2(new_n606), .ZN(new_n704));
  NOR3_X1   g0504(.A1(new_n503), .A2(new_n603), .A3(G179), .ZN(new_n705));
  NAND3_X1  g0505(.A1(new_n705), .A2(new_n515), .A3(new_n579), .ZN(new_n706));
  NAND3_X1  g0506(.A1(new_n703), .A2(new_n704), .A3(new_n706), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n707), .A2(new_n654), .ZN(new_n708));
  INV_X1    g0508(.A(new_n708), .ZN(new_n709));
  NAND4_X1  g0509(.A1(new_n518), .A2(new_n523), .A3(new_n610), .A4(new_n672), .ZN(new_n710));
  AOI21_X1  g0510(.A(new_n709), .B1(new_n710), .B2(KEYINPUT31), .ZN(new_n711));
  NAND3_X1  g0511(.A1(new_n707), .A2(KEYINPUT31), .A3(new_n654), .ZN(new_n712));
  INV_X1    g0512(.A(new_n712), .ZN(new_n713));
  OAI21_X1  g0513(.A(G330), .B1(new_n711), .B2(new_n713), .ZN(new_n714));
  AND2_X1   g0514(.A1(new_n700), .A2(new_n714), .ZN(new_n715));
  OAI21_X1  g0515(.A(new_n684), .B1(new_n715), .B2(G1), .ZN(new_n716));
  XNOR2_X1  g0516(.A(new_n716), .B(KEYINPUT91), .ZN(G364));
  AOI21_X1  g0517(.A(new_n230), .B1(G20), .B2(new_n327), .ZN(new_n718));
  NOR2_X1   g0518(.A1(new_n231), .A2(new_n309), .ZN(new_n719));
  INV_X1    g0519(.A(new_n719), .ZN(new_n720));
  NOR3_X1   g0520(.A1(new_n720), .A2(new_n300), .A3(G190), .ZN(new_n721));
  INV_X1    g0521(.A(G317), .ZN(new_n722));
  NAND2_X1  g0522(.A1(new_n722), .A2(KEYINPUT33), .ZN(new_n723));
  OR2_X1    g0523(.A1(new_n722), .A2(KEYINPUT33), .ZN(new_n724));
  NAND3_X1  g0524(.A1(new_n721), .A2(new_n723), .A3(new_n724), .ZN(new_n725));
  NOR2_X1   g0525(.A1(new_n300), .A2(G179), .ZN(new_n726));
  XNOR2_X1  g0526(.A(new_n726), .B(KEYINPUT94), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n727), .A2(G20), .ZN(new_n728));
  NOR2_X1   g0528(.A1(new_n728), .A2(G190), .ZN(new_n729));
  INV_X1    g0529(.A(new_n729), .ZN(new_n730));
  INV_X1    g0530(.A(G283), .ZN(new_n731));
  INV_X1    g0531(.A(G303), .ZN(new_n732));
  NOR2_X1   g0532(.A1(new_n728), .A2(new_n382), .ZN(new_n733));
  INV_X1    g0533(.A(new_n733), .ZN(new_n734));
  OAI221_X1 g0534(.A(new_n725), .B1(new_n730), .B2(new_n731), .C1(new_n732), .C2(new_n734), .ZN(new_n735));
  NAND2_X1  g0535(.A1(new_n719), .A2(G190), .ZN(new_n736));
  NOR2_X1   g0536(.A1(new_n736), .A2(G200), .ZN(new_n737));
  INV_X1    g0537(.A(new_n737), .ZN(new_n738));
  INV_X1    g0538(.A(G322), .ZN(new_n739));
  NOR2_X1   g0539(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  NOR3_X1   g0540(.A1(new_n720), .A2(G190), .A3(G200), .ZN(new_n741));
  INV_X1    g0541(.A(new_n741), .ZN(new_n742));
  INV_X1    g0542(.A(G311), .ZN(new_n743));
  NOR2_X1   g0543(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  NOR2_X1   g0544(.A1(G179), .A2(G200), .ZN(new_n745));
  NAND3_X1  g0545(.A1(new_n745), .A2(G20), .A3(new_n382), .ZN(new_n746));
  INV_X1    g0546(.A(new_n746), .ZN(new_n747));
  AOI21_X1  g0547(.A(new_n286), .B1(new_n747), .B2(G329), .ZN(new_n748));
  NAND2_X1  g0548(.A1(new_n745), .A2(G190), .ZN(new_n749));
  NAND2_X1  g0549(.A1(new_n749), .A2(G20), .ZN(new_n750));
  INV_X1    g0550(.A(new_n750), .ZN(new_n751));
  NOR2_X1   g0551(.A1(new_n736), .A2(new_n300), .ZN(new_n752));
  INV_X1    g0552(.A(new_n752), .ZN(new_n753));
  INV_X1    g0553(.A(G326), .ZN(new_n754));
  OAI221_X1 g0554(.A(new_n748), .B1(new_n488), .B2(new_n751), .C1(new_n753), .C2(new_n754), .ZN(new_n755));
  NOR4_X1   g0555(.A1(new_n735), .A2(new_n740), .A3(new_n744), .A4(new_n755), .ZN(new_n756));
  AOI22_X1  g0556(.A1(new_n721), .A2(G68), .B1(G97), .B2(new_n750), .ZN(new_n757));
  AOI22_X1  g0557(.A1(G77), .A2(new_n741), .B1(new_n737), .B2(G58), .ZN(new_n758));
  OAI221_X1 g0558(.A(new_n757), .B1(KEYINPUT93), .B2(new_n758), .C1(new_n734), .C2(new_n214), .ZN(new_n759));
  NAND2_X1  g0559(.A1(new_n758), .A2(KEYINPUT93), .ZN(new_n760));
  OAI211_X1 g0560(.A(new_n760), .B(new_n286), .C1(new_n730), .C2(new_n457), .ZN(new_n761));
  NOR2_X1   g0561(.A1(new_n753), .A2(new_n220), .ZN(new_n762));
  NAND2_X1  g0562(.A1(new_n747), .A2(G159), .ZN(new_n763));
  XNOR2_X1  g0563(.A(new_n763), .B(KEYINPUT32), .ZN(new_n764));
  NOR4_X1   g0564(.A1(new_n759), .A2(new_n761), .A3(new_n762), .A4(new_n764), .ZN(new_n765));
  OAI21_X1  g0565(.A(new_n718), .B1(new_n756), .B2(new_n765), .ZN(new_n766));
  NOR2_X1   g0566(.A1(new_n339), .A2(G20), .ZN(new_n767));
  NAND2_X1  g0567(.A1(new_n767), .A2(G45), .ZN(new_n768));
  NAND3_X1  g0568(.A1(new_n679), .A2(G1), .A3(new_n768), .ZN(new_n769));
  XOR2_X1   g0569(.A(new_n769), .B(KEYINPUT92), .Z(new_n770));
  INV_X1    g0570(.A(new_n770), .ZN(new_n771));
  NAND3_X1  g0571(.A1(new_n286), .A2(G355), .A3(new_n233), .ZN(new_n772));
  NOR2_X1   g0572(.A1(new_n251), .A2(new_n426), .ZN(new_n773));
  NOR2_X1   g0573(.A1(new_n677), .A2(new_n286), .ZN(new_n774));
  OAI21_X1  g0574(.A(new_n774), .B1(new_n682), .B2(G45), .ZN(new_n775));
  OAI221_X1 g0575(.A(new_n772), .B1(G116), .B2(new_n233), .C1(new_n773), .C2(new_n775), .ZN(new_n776));
  NOR2_X1   g0576(.A1(G13), .A2(G33), .ZN(new_n777));
  INV_X1    g0577(.A(new_n777), .ZN(new_n778));
  NOR2_X1   g0578(.A1(new_n778), .A2(G20), .ZN(new_n779));
  NOR2_X1   g0579(.A1(new_n779), .A2(new_n718), .ZN(new_n780));
  AOI21_X1  g0580(.A(new_n771), .B1(new_n776), .B2(new_n780), .ZN(new_n781));
  INV_X1    g0581(.A(new_n779), .ZN(new_n782));
  OAI211_X1 g0582(.A(new_n766), .B(new_n781), .C1(new_n659), .C2(new_n782), .ZN(new_n783));
  NAND2_X1  g0583(.A1(new_n660), .A2(new_n771), .ZN(new_n784));
  NOR2_X1   g0584(.A1(new_n659), .A2(G330), .ZN(new_n785));
  OAI21_X1  g0585(.A(new_n783), .B1(new_n784), .B2(new_n785), .ZN(G396));
  OAI22_X1  g0586(.A1(new_n421), .A2(new_n422), .B1(new_n420), .B2(new_n672), .ZN(new_n787));
  NAND2_X1  g0587(.A1(new_n370), .A2(new_n787), .ZN(new_n788));
  NAND3_X1  g0588(.A1(new_n359), .A2(new_n369), .A3(new_n672), .ZN(new_n789));
  NAND2_X1  g0589(.A1(new_n788), .A2(new_n789), .ZN(new_n790));
  INV_X1    g0590(.A(new_n790), .ZN(new_n791));
  NOR2_X1   g0591(.A1(new_n699), .A2(new_n791), .ZN(new_n792));
  NAND3_X1  g0592(.A1(new_n645), .A2(new_n672), .A3(new_n791), .ZN(new_n793));
  INV_X1    g0593(.A(new_n793), .ZN(new_n794));
  OR3_X1    g0594(.A1(new_n792), .A2(new_n794), .A3(new_n714), .ZN(new_n795));
  OAI21_X1  g0595(.A(new_n714), .B1(new_n792), .B2(new_n794), .ZN(new_n796));
  NAND3_X1  g0596(.A1(new_n795), .A2(new_n771), .A3(new_n796), .ZN(new_n797));
  NOR2_X1   g0597(.A1(new_n718), .A2(new_n777), .ZN(new_n798));
  NAND2_X1  g0598(.A1(new_n798), .A2(new_n222), .ZN(new_n799));
  OAI22_X1  g0599(.A1(new_n734), .A2(new_n457), .B1(new_n732), .B2(new_n753), .ZN(new_n800));
  NOR2_X1   g0600(.A1(new_n730), .A2(new_n214), .ZN(new_n801));
  OAI22_X1  g0601(.A1(new_n751), .A2(new_n447), .B1(new_n743), .B2(new_n746), .ZN(new_n802));
  OAI21_X1  g0602(.A(new_n279), .B1(new_n738), .B2(new_n488), .ZN(new_n803));
  NOR4_X1   g0603(.A1(new_n800), .A2(new_n801), .A3(new_n802), .A4(new_n803), .ZN(new_n804));
  INV_X1    g0604(.A(new_n721), .ZN(new_n805));
  OAI221_X1 g0605(.A(new_n804), .B1(new_n526), .B2(new_n742), .C1(new_n731), .C2(new_n805), .ZN(new_n806));
  AOI22_X1  g0606(.A1(G150), .A2(new_n721), .B1(new_n737), .B2(G143), .ZN(new_n807));
  INV_X1    g0607(.A(G137), .ZN(new_n808));
  INV_X1    g0608(.A(G159), .ZN(new_n809));
  OAI221_X1 g0609(.A(new_n807), .B1(new_n808), .B2(new_n753), .C1(new_n809), .C2(new_n742), .ZN(new_n810));
  XOR2_X1   g0610(.A(new_n810), .B(KEYINPUT34), .Z(new_n811));
  OAI22_X1  g0611(.A1(new_n220), .A2(new_n734), .B1(new_n730), .B2(new_n203), .ZN(new_n812));
  INV_X1    g0612(.A(KEYINPUT95), .ZN(new_n813));
  OR2_X1    g0613(.A1(new_n812), .A2(new_n813), .ZN(new_n814));
  AOI22_X1  g0614(.A1(new_n812), .A2(new_n813), .B1(G132), .B2(new_n747), .ZN(new_n815));
  NAND2_X1  g0615(.A1(new_n750), .A2(G58), .ZN(new_n816));
  NAND4_X1  g0616(.A1(new_n814), .A2(new_n815), .A3(new_n286), .A4(new_n816), .ZN(new_n817));
  OAI21_X1  g0617(.A(new_n806), .B1(new_n811), .B2(new_n817), .ZN(new_n818));
  AOI21_X1  g0618(.A(new_n771), .B1(new_n818), .B2(new_n718), .ZN(new_n819));
  OAI211_X1 g0619(.A(new_n799), .B(new_n819), .C1(new_n791), .C2(new_n778), .ZN(new_n820));
  NAND2_X1  g0620(.A1(new_n797), .A2(new_n820), .ZN(G384));
  NAND2_X1  g0621(.A1(new_n710), .A2(KEYINPUT31), .ZN(new_n822));
  NAND2_X1  g0622(.A1(new_n822), .A2(new_n708), .ZN(new_n823));
  XNOR2_X1  g0623(.A(new_n712), .B(KEYINPUT100), .ZN(new_n824));
  NAND2_X1  g0624(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  INV_X1    g0625(.A(new_n652), .ZN(new_n826));
  NAND2_X1  g0626(.A1(new_n391), .A2(new_n396), .ZN(new_n827));
  NAND2_X1  g0627(.A1(new_n827), .A2(new_n398), .ZN(new_n828));
  NAND3_X1  g0628(.A1(new_n828), .A2(new_n336), .A3(new_n397), .ZN(new_n829));
  NAND2_X1  g0629(.A1(new_n829), .A2(new_n404), .ZN(new_n830));
  OAI211_X1 g0630(.A(new_n826), .B(new_n830), .C1(new_n407), .C2(new_n417), .ZN(new_n831));
  OAI21_X1  g0631(.A(new_n414), .B1(new_n413), .B2(new_n826), .ZN(new_n832));
  NAND2_X1  g0632(.A1(new_n832), .A2(new_n405), .ZN(new_n833));
  INV_X1    g0633(.A(KEYINPUT37), .ZN(new_n834));
  NAND2_X1  g0634(.A1(new_n833), .A2(new_n834), .ZN(new_n835));
  OAI21_X1  g0635(.A(new_n830), .B1(new_n413), .B2(new_n826), .ZN(new_n836));
  NAND3_X1  g0636(.A1(new_n836), .A2(KEYINPUT37), .A3(new_n405), .ZN(new_n837));
  NAND3_X1  g0637(.A1(new_n831), .A2(new_n835), .A3(new_n837), .ZN(new_n838));
  INV_X1    g0638(.A(KEYINPUT38), .ZN(new_n839));
  NAND2_X1  g0639(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  NAND4_X1  g0640(.A1(new_n831), .A2(KEYINPUT38), .A3(new_n835), .A4(new_n837), .ZN(new_n841));
  NAND2_X1  g0641(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  NAND3_X1  g0642(.A1(new_n331), .A2(new_n349), .A3(new_n654), .ZN(new_n843));
  NAND2_X1  g0643(.A1(new_n843), .A2(KEYINPUT97), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n331), .A2(new_n349), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n349), .A2(new_n654), .ZN(new_n846));
  NAND3_X1  g0646(.A1(new_n845), .A2(new_n613), .A3(new_n846), .ZN(new_n847));
  NAND2_X1  g0647(.A1(new_n844), .A2(new_n847), .ZN(new_n848));
  NAND3_X1  g0648(.A1(new_n353), .A2(KEYINPUT97), .A3(new_n846), .ZN(new_n849));
  AOI21_X1  g0649(.A(new_n790), .B1(new_n848), .B2(new_n849), .ZN(new_n850));
  NAND3_X1  g0650(.A1(new_n825), .A2(new_n842), .A3(new_n850), .ZN(new_n851));
  INV_X1    g0651(.A(KEYINPUT40), .ZN(new_n852));
  INV_X1    g0652(.A(KEYINPUT100), .ZN(new_n853));
  XNOR2_X1  g0653(.A(new_n712), .B(new_n853), .ZN(new_n854));
  OAI21_X1  g0654(.A(new_n850), .B1(new_n711), .B2(new_n854), .ZN(new_n855));
  INV_X1    g0655(.A(new_n855), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n414), .A2(new_n826), .ZN(new_n857));
  INV_X1    g0657(.A(KEYINPUT98), .ZN(new_n858));
  AOI21_X1  g0658(.A(new_n834), .B1(new_n857), .B2(new_n858), .ZN(new_n859));
  INV_X1    g0659(.A(new_n405), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n412), .A2(new_n411), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n861), .A2(new_n409), .ZN(new_n862));
  AOI22_X1  g0662(.A1(new_n862), .A2(new_n652), .B1(new_n401), .B2(new_n404), .ZN(new_n863));
  OAI21_X1  g0663(.A(KEYINPUT99), .B1(new_n860), .B2(new_n863), .ZN(new_n864));
  INV_X1    g0664(.A(KEYINPUT99), .ZN(new_n865));
  NAND3_X1  g0665(.A1(new_n832), .A2(new_n865), .A3(new_n405), .ZN(new_n866));
  AOI21_X1  g0666(.A(new_n859), .B1(new_n864), .B2(new_n866), .ZN(new_n867));
  INV_X1    g0667(.A(new_n867), .ZN(new_n868));
  INV_X1    g0668(.A(new_n857), .ZN(new_n869));
  OAI21_X1  g0669(.A(new_n869), .B1(new_n407), .B2(new_n417), .ZN(new_n870));
  NAND3_X1  g0670(.A1(new_n864), .A2(new_n866), .A3(new_n859), .ZN(new_n871));
  NAND3_X1  g0671(.A1(new_n868), .A2(new_n870), .A3(new_n871), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n872), .A2(new_n839), .ZN(new_n873));
  AOI21_X1  g0673(.A(new_n852), .B1(new_n873), .B2(new_n841), .ZN(new_n874));
  AOI22_X1  g0674(.A1(new_n851), .A2(new_n852), .B1(new_n856), .B2(new_n874), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n825), .A2(new_n425), .ZN(new_n876));
  XNOR2_X1  g0676(.A(new_n875), .B(new_n876), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n877), .A2(G330), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n417), .A2(new_n652), .ZN(new_n879));
  INV_X1    g0679(.A(KEYINPUT39), .ZN(new_n880));
  INV_X1    g0680(.A(new_n871), .ZN(new_n881));
  NOR2_X1   g0681(.A1(new_n881), .A2(new_n867), .ZN(new_n882));
  AOI21_X1  g0682(.A(KEYINPUT38), .B1(new_n882), .B2(new_n870), .ZN(new_n883));
  INV_X1    g0683(.A(new_n841), .ZN(new_n884));
  OAI21_X1  g0684(.A(new_n880), .B1(new_n883), .B2(new_n884), .ZN(new_n885));
  NOR2_X1   g0685(.A1(new_n845), .A2(new_n654), .ZN(new_n886));
  NAND3_X1  g0686(.A1(new_n840), .A2(KEYINPUT39), .A3(new_n841), .ZN(new_n887));
  NAND3_X1  g0687(.A1(new_n885), .A2(new_n886), .A3(new_n887), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n793), .A2(new_n789), .ZN(new_n889));
  INV_X1    g0689(.A(new_n849), .ZN(new_n890));
  AOI22_X1  g0690(.A1(new_n353), .A2(new_n846), .B1(new_n843), .B2(KEYINPUT97), .ZN(new_n891));
  NOR2_X1   g0691(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  INV_X1    g0692(.A(new_n892), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n889), .A2(new_n893), .ZN(new_n894));
  INV_X1    g0694(.A(new_n842), .ZN(new_n895));
  OAI211_X1 g0695(.A(new_n879), .B(new_n888), .C1(new_n894), .C2(new_n895), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n692), .A2(new_n672), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n897), .A2(KEYINPUT29), .ZN(new_n898));
  NAND3_X1  g0698(.A1(new_n645), .A2(new_n685), .A3(new_n672), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  AOI211_X1 g0700(.A(new_n616), .B(new_n615), .C1(new_n900), .C2(new_n425), .ZN(new_n901));
  XNOR2_X1  g0701(.A(new_n896), .B(new_n901), .ZN(new_n902));
  XNOR2_X1  g0702(.A(new_n878), .B(new_n902), .ZN(new_n903));
  OAI21_X1  g0703(.A(new_n903), .B1(new_n265), .B2(new_n767), .ZN(new_n904));
  AOI21_X1  g0704(.A(new_n526), .B1(new_n459), .B2(KEYINPUT35), .ZN(new_n905));
  OAI211_X1 g0705(.A(new_n905), .B(new_n232), .C1(KEYINPUT35), .C2(new_n459), .ZN(new_n906));
  XNOR2_X1  g0706(.A(new_n906), .B(KEYINPUT36), .ZN(new_n907));
  NOR3_X1   g0707(.A1(new_n682), .A2(new_n222), .A3(new_n392), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n220), .A2(G68), .ZN(new_n909));
  XNOR2_X1  g0709(.A(new_n909), .B(KEYINPUT96), .ZN(new_n910));
  OAI211_X1 g0710(.A(G1), .B(new_n339), .C1(new_n908), .C2(new_n910), .ZN(new_n911));
  NAND3_X1  g0711(.A1(new_n904), .A2(new_n907), .A3(new_n911), .ZN(G367));
  NAND3_X1  g0712(.A1(new_n621), .A2(new_n622), .A3(new_n654), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n628), .A2(new_n913), .ZN(new_n914));
  OR2_X1    g0714(.A1(new_n913), .A2(new_n582), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n916), .A2(KEYINPUT43), .ZN(new_n917));
  INV_X1    g0717(.A(new_n916), .ZN(new_n918));
  INV_X1    g0718(.A(KEYINPUT102), .ZN(new_n919));
  INV_X1    g0719(.A(KEYINPUT43), .ZN(new_n920));
  NAND3_X1  g0720(.A1(new_n918), .A2(new_n919), .A3(new_n920), .ZN(new_n921));
  OAI21_X1  g0721(.A(KEYINPUT102), .B1(new_n916), .B2(KEYINPUT43), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  AOI21_X1  g0723(.A(new_n472), .B1(new_n514), .B2(new_n517), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n471), .A2(new_n654), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n634), .A2(new_n654), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  AND2_X1   g0728(.A1(new_n928), .A2(KEYINPUT101), .ZN(new_n929));
  NOR2_X1   g0729(.A1(new_n928), .A2(KEYINPUT101), .ZN(new_n930));
  NOR2_X1   g0730(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n931), .A2(new_n670), .ZN(new_n932));
  OR2_X1    g0732(.A1(new_n923), .A2(new_n932), .ZN(new_n933));
  NOR3_X1   g0733(.A1(new_n929), .A2(new_n930), .A3(new_n523), .ZN(new_n934));
  OAI21_X1  g0734(.A(new_n672), .B1(new_n934), .B2(new_n690), .ZN(new_n935));
  AND2_X1   g0735(.A1(new_n926), .A2(new_n927), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n673), .A2(new_n674), .ZN(new_n937));
  NOR2_X1   g0737(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  XNOR2_X1  g0738(.A(new_n938), .B(KEYINPUT42), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n935), .A2(new_n939), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n923), .A2(new_n932), .ZN(new_n941));
  AND4_X1   g0741(.A1(new_n917), .A2(new_n933), .A3(new_n940), .A4(new_n941), .ZN(new_n942));
  AOI22_X1  g0742(.A1(new_n941), .A2(new_n933), .B1(new_n940), .B2(new_n917), .ZN(new_n943));
  NOR2_X1   g0743(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  XNOR2_X1  g0744(.A(new_n678), .B(KEYINPUT41), .ZN(new_n945));
  INV_X1    g0745(.A(new_n945), .ZN(new_n946));
  INV_X1    g0746(.A(KEYINPUT105), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n629), .A2(new_n672), .ZN(new_n948));
  OAI211_X1 g0748(.A(new_n523), .B(new_n666), .C1(new_n504), .C2(new_n499), .ZN(new_n949));
  NAND4_X1  g0749(.A1(new_n948), .A2(KEYINPUT103), .A3(new_n949), .A4(new_n661), .ZN(new_n950));
  AND2_X1   g0750(.A1(new_n950), .A2(new_n937), .ZN(new_n951));
  INV_X1    g0751(.A(KEYINPUT104), .ZN(new_n952));
  INV_X1    g0752(.A(KEYINPUT103), .ZN(new_n953));
  OAI21_X1  g0753(.A(new_n953), .B1(new_n668), .B2(new_n674), .ZN(new_n954));
  NAND4_X1  g0754(.A1(new_n951), .A2(new_n952), .A3(new_n660), .A4(new_n954), .ZN(new_n955));
  NAND3_X1  g0755(.A1(new_n954), .A2(new_n937), .A3(new_n950), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n660), .A2(new_n952), .ZN(new_n957));
  NAND3_X1  g0757(.A1(new_n659), .A2(KEYINPUT104), .A3(G330), .ZN(new_n958));
  NAND3_X1  g0758(.A1(new_n956), .A2(new_n957), .A3(new_n958), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n955), .A2(new_n959), .ZN(new_n960));
  NAND4_X1  g0760(.A1(new_n700), .A2(new_n947), .A3(new_n714), .A4(new_n960), .ZN(new_n961));
  NAND4_X1  g0761(.A1(new_n898), .A2(new_n899), .A3(new_n960), .A4(new_n714), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n962), .A2(KEYINPUT105), .ZN(new_n963));
  INV_X1    g0763(.A(KEYINPUT45), .ZN(new_n964));
  XNOR2_X1  g0764(.A(new_n523), .B(KEYINPUT88), .ZN(new_n965));
  OAI21_X1  g0765(.A(new_n937), .B1(new_n965), .B2(new_n654), .ZN(new_n966));
  OAI21_X1  g0766(.A(new_n964), .B1(new_n936), .B2(new_n966), .ZN(new_n967));
  NAND3_X1  g0767(.A1(new_n675), .A2(KEYINPUT45), .A3(new_n928), .ZN(new_n968));
  AND2_X1   g0768(.A1(new_n967), .A2(new_n968), .ZN(new_n969));
  OAI21_X1  g0769(.A(KEYINPUT44), .B1(new_n675), .B2(new_n928), .ZN(new_n970));
  INV_X1    g0770(.A(KEYINPUT44), .ZN(new_n971));
  NAND3_X1  g0771(.A1(new_n936), .A2(new_n966), .A3(new_n971), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n970), .A2(new_n972), .ZN(new_n973));
  NOR3_X1   g0773(.A1(new_n969), .A2(new_n670), .A3(new_n973), .ZN(new_n974));
  AND2_X1   g0774(.A1(new_n970), .A2(new_n972), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n967), .A2(new_n968), .ZN(new_n976));
  AOI21_X1  g0776(.A(new_n671), .B1(new_n975), .B2(new_n976), .ZN(new_n977));
  NOR2_X1   g0777(.A1(new_n974), .A2(new_n977), .ZN(new_n978));
  NAND3_X1  g0778(.A1(new_n961), .A2(new_n963), .A3(new_n978), .ZN(new_n979));
  AOI21_X1  g0779(.A(new_n946), .B1(new_n979), .B2(new_n715), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n768), .A2(G1), .ZN(new_n981));
  OAI21_X1  g0781(.A(new_n944), .B1(new_n980), .B2(new_n981), .ZN(new_n982));
  INV_X1    g0782(.A(KEYINPUT106), .ZN(new_n983));
  AOI21_X1  g0783(.A(new_n771), .B1(new_n918), .B2(new_n779), .ZN(new_n984));
  INV_X1    g0784(.A(new_n774), .ZN(new_n985));
  OAI221_X1 g0785(.A(new_n780), .B1(new_n233), .B2(new_n362), .C1(new_n242), .C2(new_n985), .ZN(new_n986));
  OAI221_X1 g0786(.A(new_n279), .B1(new_n738), .B2(new_n732), .C1(new_n743), .C2(new_n753), .ZN(new_n987));
  OAI22_X1  g0787(.A1(new_n730), .A2(new_n447), .B1(new_n457), .B2(new_n751), .ZN(new_n988));
  AOI211_X1 g0788(.A(new_n987), .B(new_n988), .C1(G317), .C2(new_n747), .ZN(new_n989));
  NOR2_X1   g0789(.A1(new_n734), .A2(new_n526), .ZN(new_n990));
  AOI22_X1  g0790(.A1(new_n990), .A2(KEYINPUT46), .B1(G283), .B2(new_n741), .ZN(new_n991));
  AND2_X1   g0791(.A1(new_n989), .A2(new_n991), .ZN(new_n992));
  OAI221_X1 g0792(.A(new_n992), .B1(KEYINPUT46), .B2(new_n990), .C1(new_n488), .C2(new_n805), .ZN(new_n993));
  AOI22_X1  g0793(.A1(new_n752), .A2(G143), .B1(G68), .B2(new_n750), .ZN(new_n994));
  OAI221_X1 g0794(.A(new_n994), .B1(new_n808), .B2(new_n746), .C1(new_n730), .C2(new_n222), .ZN(new_n995));
  AOI211_X1 g0795(.A(new_n279), .B(new_n995), .C1(G58), .C2(new_n733), .ZN(new_n996));
  OAI221_X1 g0796(.A(new_n996), .B1(new_n220), .B2(new_n742), .C1(new_n809), .C2(new_n805), .ZN(new_n997));
  INV_X1    g0797(.A(G150), .ZN(new_n998));
  NOR2_X1   g0798(.A1(new_n738), .A2(new_n998), .ZN(new_n999));
  OAI21_X1  g0799(.A(new_n993), .B1(new_n997), .B2(new_n999), .ZN(new_n1000));
  XOR2_X1   g0800(.A(new_n1000), .B(KEYINPUT47), .Z(new_n1001));
  INV_X1    g0801(.A(new_n718), .ZN(new_n1002));
  OAI211_X1 g0802(.A(new_n984), .B(new_n986), .C1(new_n1001), .C2(new_n1002), .ZN(new_n1003));
  AND3_X1   g0803(.A1(new_n982), .A2(new_n983), .A3(new_n1003), .ZN(new_n1004));
  AOI21_X1  g0804(.A(new_n983), .B1(new_n982), .B2(new_n1003), .ZN(new_n1005));
  NOR2_X1   g0805(.A1(new_n1004), .A2(new_n1005), .ZN(new_n1006));
  INV_X1    g0806(.A(new_n1006), .ZN(G387));
  OAI22_X1  g0807(.A1(new_n730), .A2(new_n447), .B1(new_n203), .B2(new_n742), .ZN(new_n1008));
  NOR2_X1   g0808(.A1(new_n734), .A2(new_n222), .ZN(new_n1009));
  OAI21_X1  g0809(.A(new_n286), .B1(new_n753), .B2(new_n809), .ZN(new_n1010));
  NOR2_X1   g0810(.A1(new_n746), .A2(new_n998), .ZN(new_n1011));
  NOR4_X1   g0811(.A1(new_n1008), .A2(new_n1009), .A3(new_n1010), .A4(new_n1011), .ZN(new_n1012));
  NAND2_X1  g0812(.A1(new_n721), .A2(new_n259), .ZN(new_n1013));
  NOR2_X1   g0813(.A1(new_n751), .A2(new_n362), .ZN(new_n1014));
  INV_X1    g0814(.A(new_n1014), .ZN(new_n1015));
  NAND2_X1  g0815(.A1(new_n737), .A2(G50), .ZN(new_n1016));
  NAND4_X1  g0816(.A1(new_n1012), .A2(new_n1013), .A3(new_n1015), .A4(new_n1016), .ZN(new_n1017));
  AOI22_X1  g0817(.A1(G311), .A2(new_n721), .B1(new_n737), .B2(G317), .ZN(new_n1018));
  OAI221_X1 g0818(.A(new_n1018), .B1(new_n732), .B2(new_n742), .C1(new_n739), .C2(new_n753), .ZN(new_n1019));
  XNOR2_X1  g0819(.A(new_n1019), .B(KEYINPUT48), .ZN(new_n1020));
  OAI221_X1 g0820(.A(new_n1020), .B1(new_n731), .B2(new_n751), .C1(new_n488), .C2(new_n734), .ZN(new_n1021));
  XOR2_X1   g0821(.A(new_n1021), .B(KEYINPUT49), .Z(new_n1022));
  OAI221_X1 g0822(.A(new_n279), .B1(new_n754), .B2(new_n746), .C1(new_n730), .C2(new_n526), .ZN(new_n1023));
  OAI21_X1  g0823(.A(new_n1017), .B1(new_n1022), .B2(new_n1023), .ZN(new_n1024));
  AOI21_X1  g0824(.A(new_n771), .B1(new_n1024), .B2(new_n718), .ZN(new_n1025));
  OAI21_X1  g0825(.A(new_n1025), .B1(new_n668), .B2(new_n782), .ZN(new_n1026));
  AOI21_X1  g0826(.A(new_n985), .B1(new_n246), .B2(G45), .ZN(new_n1027));
  OR3_X1    g0827(.A1(new_n365), .A2(KEYINPUT50), .A3(G50), .ZN(new_n1028));
  OAI21_X1  g0828(.A(KEYINPUT50), .B1(new_n365), .B2(G50), .ZN(new_n1029));
  NAND4_X1  g0829(.A1(new_n1028), .A2(new_n1029), .A3(new_n426), .A4(new_n680), .ZN(new_n1030));
  NOR2_X1   g0830(.A1(new_n203), .A2(new_n222), .ZN(new_n1031));
  OAI21_X1  g0831(.A(new_n1027), .B1(new_n1030), .B2(new_n1031), .ZN(new_n1032));
  NAND2_X1  g0832(.A1(new_n286), .A2(new_n233), .ZN(new_n1033));
  OAI221_X1 g0833(.A(new_n1032), .B1(G107), .B2(new_n233), .C1(new_n680), .C2(new_n1033), .ZN(new_n1034));
  XOR2_X1   g0834(.A(new_n1034), .B(KEYINPUT107), .Z(new_n1035));
  AOI21_X1  g0835(.A(new_n1026), .B1(new_n780), .B2(new_n1035), .ZN(new_n1036));
  AOI21_X1  g0836(.A(new_n1036), .B1(new_n981), .B2(new_n960), .ZN(new_n1037));
  NAND2_X1  g0837(.A1(new_n961), .A2(new_n963), .ZN(new_n1038));
  OAI21_X1  g0838(.A(new_n1038), .B1(new_n715), .B2(new_n960), .ZN(new_n1039));
  OAI21_X1  g0839(.A(new_n1037), .B1(new_n1039), .B2(new_n679), .ZN(G393));
  OAI21_X1  g0840(.A(new_n780), .B1(new_n254), .B2(new_n985), .ZN(new_n1041));
  AOI21_X1  g0841(.A(new_n1041), .B1(G97), .B2(new_n677), .ZN(new_n1042));
  OAI22_X1  g0842(.A1(new_n730), .A2(new_n457), .B1(new_n488), .B2(new_n742), .ZN(new_n1043));
  AOI22_X1  g0843(.A1(G311), .A2(new_n737), .B1(new_n752), .B2(G317), .ZN(new_n1044));
  AOI21_X1  g0844(.A(new_n1043), .B1(KEYINPUT52), .B2(new_n1044), .ZN(new_n1045));
  OAI21_X1  g0845(.A(new_n1045), .B1(new_n732), .B2(new_n805), .ZN(new_n1046));
  OAI221_X1 g0846(.A(new_n279), .B1(KEYINPUT52), .B2(new_n1044), .C1(new_n734), .C2(new_n731), .ZN(new_n1047));
  NOR2_X1   g0847(.A1(new_n1046), .A2(new_n1047), .ZN(new_n1048));
  OAI221_X1 g0848(.A(new_n1048), .B1(new_n526), .B2(new_n751), .C1(new_n739), .C2(new_n746), .ZN(new_n1049));
  NOR2_X1   g0849(.A1(new_n751), .A2(new_n222), .ZN(new_n1050));
  OAI21_X1  g0850(.A(new_n286), .B1(new_n365), .B2(new_n742), .ZN(new_n1051));
  AOI22_X1  g0851(.A1(G150), .A2(new_n752), .B1(new_n737), .B2(G159), .ZN(new_n1052));
  OAI22_X1  g0852(.A1(new_n1052), .A2(KEYINPUT51), .B1(new_n220), .B2(new_n805), .ZN(new_n1053));
  AOI211_X1 g0853(.A(new_n1051), .B(new_n1053), .C1(G143), .C2(new_n747), .ZN(new_n1054));
  AOI21_X1  g0854(.A(new_n801), .B1(KEYINPUT51), .B2(new_n1052), .ZN(new_n1055));
  OAI211_X1 g0855(.A(new_n1054), .B(new_n1055), .C1(new_n203), .C2(new_n734), .ZN(new_n1056));
  OAI21_X1  g0856(.A(new_n1049), .B1(new_n1050), .B2(new_n1056), .ZN(new_n1057));
  AOI211_X1 g0857(.A(new_n771), .B(new_n1042), .C1(new_n1057), .C2(new_n718), .ZN(new_n1058));
  OAI21_X1  g0858(.A(new_n1058), .B1(new_n931), .B2(new_n782), .ZN(new_n1059));
  OAI21_X1  g0859(.A(new_n670), .B1(new_n969), .B2(new_n973), .ZN(new_n1060));
  NAND3_X1  g0860(.A1(new_n975), .A2(new_n671), .A3(new_n976), .ZN(new_n1061));
  NAND2_X1  g0861(.A1(new_n1060), .A2(new_n1061), .ZN(new_n1062));
  INV_X1    g0862(.A(new_n981), .ZN(new_n1063));
  OAI21_X1  g0863(.A(new_n1059), .B1(new_n1062), .B2(new_n1063), .ZN(new_n1064));
  XNOR2_X1  g0864(.A(new_n1064), .B(KEYINPUT108), .ZN(new_n1065));
  NAND2_X1  g0865(.A1(new_n1038), .A2(new_n1062), .ZN(new_n1066));
  NAND3_X1  g0866(.A1(new_n1066), .A2(new_n678), .A3(new_n979), .ZN(new_n1067));
  NAND2_X1  g0867(.A1(new_n1065), .A2(new_n1067), .ZN(G390));
  INV_X1    g0868(.A(KEYINPUT112), .ZN(new_n1069));
  INV_X1    g0869(.A(KEYINPUT109), .ZN(new_n1070));
  INV_X1    g0870(.A(new_n886), .ZN(new_n1071));
  NAND3_X1  g0871(.A1(new_n894), .A2(new_n1070), .A3(new_n1071), .ZN(new_n1072));
  NAND2_X1  g0872(.A1(new_n885), .A2(new_n887), .ZN(new_n1073));
  AOI21_X1  g0873(.A(new_n892), .B1(new_n793), .B2(new_n789), .ZN(new_n1074));
  OAI21_X1  g0874(.A(KEYINPUT109), .B1(new_n1074), .B2(new_n886), .ZN(new_n1075));
  NAND3_X1  g0875(.A1(new_n1072), .A2(new_n1073), .A3(new_n1075), .ZN(new_n1076));
  NAND3_X1  g0876(.A1(new_n692), .A2(new_n672), .A3(new_n788), .ZN(new_n1077));
  NAND2_X1  g0877(.A1(new_n1077), .A2(new_n789), .ZN(new_n1078));
  NAND2_X1  g0878(.A1(new_n1078), .A2(new_n893), .ZN(new_n1079));
  OAI211_X1 g0879(.A(new_n1079), .B(new_n1071), .C1(new_n884), .C2(new_n883), .ZN(new_n1080));
  NAND2_X1  g0880(.A1(new_n1076), .A2(new_n1080), .ZN(new_n1081));
  NAND3_X1  g0881(.A1(new_n825), .A2(G330), .A3(new_n850), .ZN(new_n1082));
  NAND2_X1  g0882(.A1(new_n1081), .A2(new_n1082), .ZN(new_n1083));
  NOR3_X1   g0883(.A1(new_n714), .A2(new_n790), .A3(new_n892), .ZN(new_n1084));
  NAND3_X1  g0884(.A1(new_n1076), .A2(new_n1080), .A3(new_n1084), .ZN(new_n1085));
  AOI21_X1  g0885(.A(new_n1063), .B1(new_n1083), .B2(new_n1085), .ZN(new_n1086));
  NAND2_X1  g0886(.A1(new_n1073), .A2(new_n777), .ZN(new_n1087));
  XOR2_X1   g0887(.A(KEYINPUT54), .B(G143), .Z(new_n1088));
  INV_X1    g0888(.A(new_n1088), .ZN(new_n1089));
  OAI22_X1  g0889(.A1(new_n730), .A2(new_n220), .B1(new_n742), .B2(new_n1089), .ZN(new_n1090));
  INV_X1    g0890(.A(G128), .ZN(new_n1091));
  NOR2_X1   g0891(.A1(new_n753), .A2(new_n1091), .ZN(new_n1092));
  NAND2_X1  g0892(.A1(new_n733), .A2(G150), .ZN(new_n1093));
  XNOR2_X1  g0893(.A(KEYINPUT111), .B(KEYINPUT53), .ZN(new_n1094));
  NOR2_X1   g0894(.A1(new_n1093), .A2(new_n1094), .ZN(new_n1095));
  AND2_X1   g0895(.A1(new_n747), .A2(G125), .ZN(new_n1096));
  OAI21_X1  g0896(.A(new_n286), .B1(new_n751), .B2(new_n809), .ZN(new_n1097));
  OR4_X1    g0897(.A1(new_n1092), .A2(new_n1095), .A3(new_n1096), .A4(new_n1097), .ZN(new_n1098));
  AOI211_X1 g0898(.A(new_n1090), .B(new_n1098), .C1(new_n1093), .C2(new_n1094), .ZN(new_n1099));
  INV_X1    g0899(.A(G132), .ZN(new_n1100));
  OAI221_X1 g0900(.A(new_n1099), .B1(new_n1100), .B2(new_n738), .C1(new_n808), .C2(new_n805), .ZN(new_n1101));
  NOR2_X1   g0901(.A1(new_n730), .A2(new_n203), .ZN(new_n1102));
  OAI22_X1  g0902(.A1(new_n734), .A2(new_n214), .B1(new_n457), .B2(new_n805), .ZN(new_n1103));
  AOI211_X1 g0903(.A(new_n1102), .B(new_n1103), .C1(G283), .C2(new_n752), .ZN(new_n1104));
  AOI211_X1 g0904(.A(new_n286), .B(new_n1050), .C1(G294), .C2(new_n747), .ZN(new_n1105));
  AND2_X1   g0905(.A1(new_n1104), .A2(new_n1105), .ZN(new_n1106));
  OAI221_X1 g0906(.A(new_n1106), .B1(new_n447), .B2(new_n742), .C1(new_n526), .C2(new_n738), .ZN(new_n1107));
  AOI21_X1  g0907(.A(new_n1002), .B1(new_n1101), .B2(new_n1107), .ZN(new_n1108));
  INV_X1    g0908(.A(new_n259), .ZN(new_n1109));
  AOI211_X1 g0909(.A(new_n771), .B(new_n1108), .C1(new_n1109), .C2(new_n798), .ZN(new_n1110));
  NAND2_X1  g0910(.A1(new_n1087), .A2(new_n1110), .ZN(new_n1111));
  INV_X1    g0911(.A(new_n1111), .ZN(new_n1112));
  OAI21_X1  g0912(.A(new_n1069), .B1(new_n1086), .B2(new_n1112), .ZN(new_n1113));
  AND3_X1   g0913(.A1(new_n1076), .A2(new_n1080), .A3(new_n1084), .ZN(new_n1114));
  INV_X1    g0914(.A(new_n1082), .ZN(new_n1115));
  AOI21_X1  g0915(.A(new_n1115), .B1(new_n1076), .B2(new_n1080), .ZN(new_n1116));
  OAI21_X1  g0916(.A(new_n981), .B1(new_n1114), .B2(new_n1116), .ZN(new_n1117));
  NAND3_X1  g0917(.A1(new_n1117), .A2(KEYINPUT112), .A3(new_n1111), .ZN(new_n1118));
  NAND3_X1  g0918(.A1(new_n825), .A2(G330), .A3(new_n425), .ZN(new_n1119));
  XNOR2_X1  g0919(.A(new_n1119), .B(KEYINPUT110), .ZN(new_n1120));
  OAI211_X1 g0920(.A(G330), .B(new_n791), .C1(new_n711), .C2(new_n854), .ZN(new_n1121));
  AND2_X1   g0921(.A1(new_n1121), .A2(new_n892), .ZN(new_n1122));
  NOR3_X1   g0922(.A1(new_n1122), .A2(new_n1084), .A3(new_n1078), .ZN(new_n1123));
  OAI21_X1  g0923(.A(new_n892), .B1(new_n714), .B2(new_n790), .ZN(new_n1124));
  AOI22_X1  g0924(.A1(new_n1124), .A2(new_n1082), .B1(new_n789), .B2(new_n793), .ZN(new_n1125));
  OAI211_X1 g0925(.A(new_n1120), .B(new_n901), .C1(new_n1123), .C2(new_n1125), .ZN(new_n1126));
  INV_X1    g0926(.A(new_n1126), .ZN(new_n1127));
  OAI21_X1  g0927(.A(new_n1127), .B1(new_n1114), .B2(new_n1116), .ZN(new_n1128));
  NAND3_X1  g0928(.A1(new_n1083), .A2(new_n1085), .A3(new_n1126), .ZN(new_n1129));
  NAND3_X1  g0929(.A1(new_n1128), .A2(new_n1129), .A3(new_n678), .ZN(new_n1130));
  NAND3_X1  g0930(.A1(new_n1113), .A2(new_n1118), .A3(new_n1130), .ZN(G378));
  INV_X1    g0931(.A(new_n896), .ZN(new_n1132));
  XOR2_X1   g0932(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1133));
  XNOR2_X1  g0933(.A(new_n312), .B(new_n1133), .ZN(new_n1134));
  NAND2_X1  g0934(.A1(new_n272), .A2(new_n826), .ZN(new_n1135));
  NAND2_X1  g0935(.A1(new_n1134), .A2(new_n1135), .ZN(new_n1136));
  OR2_X1    g0936(.A1(new_n312), .A2(new_n1133), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n312), .A2(new_n1133), .ZN(new_n1138));
  NAND4_X1  g0938(.A1(new_n1137), .A2(new_n272), .A3(new_n826), .A4(new_n1138), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n1136), .A2(new_n1139), .ZN(new_n1140));
  AOI21_X1  g0940(.A(new_n1140), .B1(new_n875), .B2(G330), .ZN(new_n1141));
  OAI21_X1  g0941(.A(new_n852), .B1(new_n895), .B2(new_n855), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n856), .A2(new_n874), .ZN(new_n1143));
  AND4_X1   g0943(.A1(G330), .A2(new_n1142), .A3(new_n1143), .A4(new_n1140), .ZN(new_n1144));
  OAI21_X1  g0944(.A(new_n1132), .B1(new_n1141), .B2(new_n1144), .ZN(new_n1145));
  NAND3_X1  g0945(.A1(new_n1143), .A2(new_n1142), .A3(G330), .ZN(new_n1146));
  INV_X1    g0946(.A(new_n1140), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n1146), .A2(new_n1147), .ZN(new_n1148));
  NAND3_X1  g0948(.A1(new_n875), .A2(G330), .A3(new_n1140), .ZN(new_n1149));
  NAND3_X1  g0949(.A1(new_n1148), .A2(new_n1149), .A3(new_n896), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n1145), .A2(new_n1150), .ZN(new_n1151));
  NAND2_X1  g0951(.A1(new_n1151), .A2(new_n981), .ZN(new_n1152));
  AOI21_X1  g0952(.A(new_n771), .B1(new_n220), .B2(new_n798), .ZN(new_n1153));
  INV_X1    g0953(.A(G124), .ZN(new_n1154));
  OAI21_X1  g0954(.A(new_n260), .B1(new_n746), .B2(new_n1154), .ZN(new_n1155));
  NOR2_X1   g0955(.A1(new_n738), .A2(new_n1091), .ZN(new_n1156));
  AOI22_X1  g0956(.A1(G132), .A2(new_n721), .B1(new_n741), .B2(G137), .ZN(new_n1157));
  XOR2_X1   g0957(.A(new_n1157), .B(KEYINPUT115), .Z(new_n1158));
  AOI211_X1 g0958(.A(new_n1156), .B(new_n1158), .C1(G125), .C2(new_n752), .ZN(new_n1159));
  OAI221_X1 g0959(.A(new_n1159), .B1(new_n998), .B2(new_n751), .C1(new_n734), .C2(new_n1089), .ZN(new_n1160));
  XOR2_X1   g0960(.A(KEYINPUT116), .B(KEYINPUT59), .Z(new_n1161));
  AOI211_X1 g0961(.A(G41), .B(new_n1155), .C1(new_n1160), .C2(new_n1161), .ZN(new_n1162));
  OAI221_X1 g0962(.A(new_n1162), .B1(new_n809), .B2(new_n730), .C1(new_n1161), .C2(new_n1160), .ZN(new_n1163));
  INV_X1    g0963(.A(KEYINPUT114), .ZN(new_n1164));
  AOI22_X1  g0964(.A1(new_n363), .A2(new_n741), .B1(new_n721), .B2(G97), .ZN(new_n1165));
  AOI21_X1  g0965(.A(new_n1009), .B1(new_n1164), .B2(new_n1165), .ZN(new_n1166));
  OAI221_X1 g0966(.A(new_n1166), .B1(new_n457), .B2(new_n738), .C1(new_n731), .C2(new_n746), .ZN(new_n1167));
  OR2_X1    g0967(.A1(new_n1165), .A2(new_n1164), .ZN(new_n1168));
  NAND2_X1  g0968(.A1(new_n729), .A2(G58), .ZN(new_n1169));
  AOI22_X1  g0969(.A1(new_n752), .A2(G116), .B1(G68), .B2(new_n750), .ZN(new_n1170));
  NAND4_X1  g0970(.A1(new_n1168), .A2(new_n279), .A3(new_n1169), .A4(new_n1170), .ZN(new_n1171));
  NOR3_X1   g0971(.A1(new_n1167), .A2(G41), .A3(new_n1171), .ZN(new_n1172));
  XOR2_X1   g0972(.A(new_n1172), .B(KEYINPUT58), .Z(new_n1173));
  OAI21_X1  g0973(.A(new_n220), .B1(new_n277), .B2(G41), .ZN(new_n1174));
  XNOR2_X1  g0974(.A(new_n1174), .B(KEYINPUT113), .ZN(new_n1175));
  AND3_X1   g0975(.A1(new_n1163), .A2(new_n1173), .A3(new_n1175), .ZN(new_n1176));
  OAI221_X1 g0976(.A(new_n1153), .B1(new_n1002), .B2(new_n1176), .C1(new_n1147), .C2(new_n778), .ZN(new_n1177));
  NAND2_X1  g0977(.A1(new_n1152), .A2(new_n1177), .ZN(new_n1178));
  INV_X1    g0978(.A(new_n1178), .ZN(new_n1179));
  NAND2_X1  g0979(.A1(new_n1120), .A2(new_n901), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n1083), .A2(new_n1085), .ZN(new_n1181));
  AOI21_X1  g0981(.A(new_n1180), .B1(new_n1181), .B2(new_n1127), .ZN(new_n1182));
  INV_X1    g0982(.A(KEYINPUT117), .ZN(new_n1183));
  NAND3_X1  g0983(.A1(new_n1145), .A2(new_n1183), .A3(new_n1150), .ZN(new_n1184));
  OAI211_X1 g0984(.A(KEYINPUT117), .B(new_n1132), .C1(new_n1141), .C2(new_n1144), .ZN(new_n1185));
  NAND3_X1  g0985(.A1(new_n1184), .A2(KEYINPUT57), .A3(new_n1185), .ZN(new_n1186));
  OAI21_X1  g0986(.A(new_n678), .B1(new_n1182), .B2(new_n1186), .ZN(new_n1187));
  INV_X1    g0987(.A(new_n1180), .ZN(new_n1188));
  NAND2_X1  g0988(.A1(new_n1128), .A2(new_n1188), .ZN(new_n1189));
  AOI21_X1  g0989(.A(KEYINPUT57), .B1(new_n1189), .B2(new_n1151), .ZN(new_n1190));
  OAI21_X1  g0990(.A(new_n1179), .B1(new_n1187), .B2(new_n1190), .ZN(G375));
  NOR2_X1   g0991(.A1(new_n1123), .A2(new_n1125), .ZN(new_n1192));
  NAND2_X1  g0992(.A1(new_n1192), .A2(new_n1180), .ZN(new_n1193));
  NAND3_X1  g0993(.A1(new_n1193), .A2(new_n945), .A3(new_n1126), .ZN(new_n1194));
  XOR2_X1   g0994(.A(new_n1194), .B(KEYINPUT118), .Z(new_n1195));
  OAI22_X1  g0995(.A1(new_n730), .A2(new_n222), .B1(new_n488), .B2(new_n753), .ZN(new_n1196));
  NOR2_X1   g0996(.A1(new_n734), .A2(new_n447), .ZN(new_n1197));
  NOR2_X1   g0997(.A1(new_n805), .A2(new_n526), .ZN(new_n1198));
  OAI211_X1 g0998(.A(new_n1015), .B(new_n279), .C1(new_n731), .C2(new_n738), .ZN(new_n1199));
  NOR4_X1   g0999(.A1(new_n1196), .A2(new_n1197), .A3(new_n1198), .A4(new_n1199), .ZN(new_n1200));
  OAI221_X1 g1000(.A(new_n1200), .B1(new_n457), .B2(new_n742), .C1(new_n732), .C2(new_n746), .ZN(new_n1201));
  OAI21_X1  g1001(.A(new_n1169), .B1(new_n1100), .B2(new_n753), .ZN(new_n1202));
  NOR2_X1   g1002(.A1(new_n734), .A2(new_n809), .ZN(new_n1203));
  NOR2_X1   g1003(.A1(new_n751), .A2(new_n220), .ZN(new_n1204));
  OAI221_X1 g1004(.A(new_n286), .B1(new_n746), .B2(new_n1091), .C1(new_n738), .C2(new_n808), .ZN(new_n1205));
  NOR4_X1   g1005(.A1(new_n1202), .A2(new_n1203), .A3(new_n1204), .A4(new_n1205), .ZN(new_n1206));
  OAI221_X1 g1006(.A(new_n1206), .B1(new_n998), .B2(new_n742), .C1(new_n805), .C2(new_n1089), .ZN(new_n1207));
  AOI21_X1  g1007(.A(new_n1002), .B1(new_n1201), .B2(new_n1207), .ZN(new_n1208));
  AOI211_X1 g1008(.A(new_n771), .B(new_n1208), .C1(new_n203), .C2(new_n798), .ZN(new_n1209));
  OAI21_X1  g1009(.A(new_n1209), .B1(new_n893), .B2(new_n778), .ZN(new_n1210));
  OAI21_X1  g1010(.A(new_n1210), .B1(new_n1192), .B2(new_n1063), .ZN(new_n1211));
  INV_X1    g1011(.A(new_n1211), .ZN(new_n1212));
  NAND2_X1  g1012(.A1(new_n1195), .A2(new_n1212), .ZN(G381));
  INV_X1    g1013(.A(G384), .ZN(new_n1214));
  NOR2_X1   g1014(.A1(G393), .A2(G396), .ZN(new_n1215));
  NAND4_X1  g1015(.A1(new_n1195), .A2(new_n1214), .A3(new_n1212), .A4(new_n1215), .ZN(new_n1216));
  INV_X1    g1016(.A(G390), .ZN(new_n1217));
  NAND2_X1  g1017(.A1(new_n1006), .A2(new_n1217), .ZN(new_n1218));
  NOR2_X1   g1018(.A1(new_n1216), .A2(new_n1218), .ZN(new_n1219));
  OR2_X1    g1019(.A1(new_n1219), .A2(KEYINPUT119), .ZN(new_n1220));
  NOR2_X1   g1020(.A1(G375), .A2(G378), .ZN(new_n1221));
  NAND2_X1  g1021(.A1(new_n1219), .A2(KEYINPUT119), .ZN(new_n1222));
  NAND3_X1  g1022(.A1(new_n1220), .A2(new_n1221), .A3(new_n1222), .ZN(G407));
  NAND2_X1  g1023(.A1(new_n653), .A2(G213), .ZN(new_n1224));
  XOR2_X1   g1024(.A(new_n1224), .B(KEYINPUT120), .Z(new_n1225));
  INV_X1    g1025(.A(new_n1225), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n1221), .A2(new_n1226), .ZN(new_n1227));
  NAND3_X1  g1027(.A1(G407), .A2(G213), .A3(new_n1227), .ZN(new_n1228));
  INV_X1    g1028(.A(KEYINPUT121), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n1228), .A2(new_n1229), .ZN(new_n1230));
  NAND4_X1  g1030(.A1(G407), .A2(KEYINPUT121), .A3(G213), .A4(new_n1227), .ZN(new_n1231));
  NAND2_X1  g1031(.A1(new_n1230), .A2(new_n1231), .ZN(G409));
  OAI211_X1 g1032(.A(G378), .B(new_n1179), .C1(new_n1187), .C2(new_n1190), .ZN(new_n1233));
  AND3_X1   g1033(.A1(new_n1113), .A2(new_n1118), .A3(new_n1130), .ZN(new_n1234));
  AOI21_X1  g1034(.A(new_n1126), .B1(new_n1083), .B2(new_n1085), .ZN(new_n1235));
  OAI211_X1 g1035(.A(new_n945), .B(new_n1151), .C1(new_n1235), .C2(new_n1180), .ZN(new_n1236));
  NAND3_X1  g1036(.A1(new_n1184), .A2(new_n981), .A3(new_n1185), .ZN(new_n1237));
  NAND3_X1  g1037(.A1(new_n1236), .A2(new_n1177), .A3(new_n1237), .ZN(new_n1238));
  NAND2_X1  g1038(.A1(new_n1234), .A2(new_n1238), .ZN(new_n1239));
  NAND2_X1  g1039(.A1(new_n1233), .A2(new_n1239), .ZN(new_n1240));
  NAND2_X1  g1040(.A1(new_n1240), .A2(new_n1224), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(new_n1241), .A2(KEYINPUT123), .ZN(new_n1242));
  INV_X1    g1042(.A(KEYINPUT60), .ZN(new_n1243));
  AOI21_X1  g1043(.A(new_n1243), .B1(new_n1193), .B2(new_n1126), .ZN(new_n1244));
  AOI21_X1  g1044(.A(KEYINPUT60), .B1(new_n1192), .B2(new_n1180), .ZN(new_n1245));
  NOR3_X1   g1045(.A1(new_n1244), .A2(new_n679), .A3(new_n1245), .ZN(new_n1246));
  INV_X1    g1046(.A(new_n1246), .ZN(new_n1247));
  OR2_X1    g1047(.A1(G384), .A2(KEYINPUT122), .ZN(new_n1248));
  NAND2_X1  g1048(.A1(G384), .A2(KEYINPUT122), .ZN(new_n1249));
  NAND4_X1  g1049(.A1(new_n1247), .A2(new_n1212), .A3(new_n1248), .A4(new_n1249), .ZN(new_n1250));
  OAI211_X1 g1050(.A(KEYINPUT122), .B(G384), .C1(new_n1246), .C2(new_n1211), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n1250), .A2(new_n1251), .ZN(new_n1252));
  INV_X1    g1052(.A(G2897), .ZN(new_n1253));
  OAI21_X1  g1053(.A(new_n1252), .B1(new_n1253), .B2(new_n1224), .ZN(new_n1254));
  NAND4_X1  g1054(.A1(new_n1250), .A2(new_n1251), .A3(G2897), .A4(new_n1226), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(new_n1254), .A2(new_n1255), .ZN(new_n1256));
  INV_X1    g1056(.A(new_n1256), .ZN(new_n1257));
  INV_X1    g1057(.A(KEYINPUT123), .ZN(new_n1258));
  NAND3_X1  g1058(.A1(new_n1240), .A2(new_n1258), .A3(new_n1224), .ZN(new_n1259));
  NAND3_X1  g1059(.A1(new_n1242), .A2(new_n1257), .A3(new_n1259), .ZN(new_n1260));
  OAI211_X1 g1060(.A(KEYINPUT124), .B(new_n1217), .C1(new_n1004), .C2(new_n1005), .ZN(new_n1261));
  XOR2_X1   g1061(.A(G393), .B(G396), .Z(new_n1262));
  INV_X1    g1062(.A(new_n1262), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n982), .A2(new_n1003), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(new_n1264), .A2(KEYINPUT106), .ZN(new_n1265));
  NAND3_X1  g1065(.A1(new_n982), .A2(new_n983), .A3(new_n1003), .ZN(new_n1266));
  AOI21_X1  g1066(.A(G390), .B1(new_n1265), .B2(new_n1266), .ZN(new_n1267));
  NAND3_X1  g1067(.A1(G390), .A2(new_n982), .A3(new_n1003), .ZN(new_n1268));
  AND2_X1   g1068(.A1(new_n1268), .A2(KEYINPUT124), .ZN(new_n1269));
  OAI211_X1 g1069(.A(new_n1261), .B(new_n1263), .C1(new_n1267), .C2(new_n1269), .ZN(new_n1270));
  INV_X1    g1070(.A(new_n1268), .ZN(new_n1271));
  AOI21_X1  g1071(.A(G390), .B1(new_n1003), .B2(new_n982), .ZN(new_n1272));
  OAI21_X1  g1072(.A(new_n1262), .B1(new_n1271), .B2(new_n1272), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(new_n1270), .A2(new_n1273), .ZN(new_n1274));
  INV_X1    g1074(.A(KEYINPUT61), .ZN(new_n1275));
  AND3_X1   g1075(.A1(new_n1274), .A2(KEYINPUT125), .A3(new_n1275), .ZN(new_n1276));
  AOI21_X1  g1076(.A(KEYINPUT125), .B1(new_n1274), .B2(new_n1275), .ZN(new_n1277));
  NOR2_X1   g1077(.A1(new_n1276), .A2(new_n1277), .ZN(new_n1278));
  AOI21_X1  g1078(.A(new_n1226), .B1(new_n1233), .B2(new_n1239), .ZN(new_n1279));
  NAND3_X1  g1079(.A1(new_n1279), .A2(KEYINPUT63), .A3(new_n1252), .ZN(new_n1280));
  INV_X1    g1080(.A(KEYINPUT63), .ZN(new_n1281));
  INV_X1    g1081(.A(new_n1252), .ZN(new_n1282));
  OAI21_X1  g1082(.A(new_n1281), .B1(new_n1241), .B2(new_n1282), .ZN(new_n1283));
  NAND4_X1  g1083(.A1(new_n1260), .A2(new_n1278), .A3(new_n1280), .A4(new_n1283), .ZN(new_n1284));
  INV_X1    g1084(.A(new_n1274), .ZN(new_n1285));
  INV_X1    g1085(.A(KEYINPUT62), .ZN(new_n1286));
  NAND4_X1  g1086(.A1(new_n1240), .A2(new_n1286), .A3(new_n1224), .A4(new_n1252), .ZN(new_n1287));
  XOR2_X1   g1087(.A(KEYINPUT126), .B(KEYINPUT61), .Z(new_n1288));
  OAI211_X1 g1088(.A(new_n1287), .B(new_n1288), .C1(new_n1256), .C2(new_n1279), .ZN(new_n1289));
  AOI21_X1  g1089(.A(new_n1286), .B1(new_n1279), .B2(new_n1252), .ZN(new_n1290));
  OAI21_X1  g1090(.A(new_n1285), .B1(new_n1289), .B2(new_n1290), .ZN(new_n1291));
  NAND2_X1  g1091(.A1(new_n1284), .A2(new_n1291), .ZN(G405));
  AND3_X1   g1092(.A1(new_n1184), .A2(KEYINPUT57), .A3(new_n1185), .ZN(new_n1293));
  AOI21_X1  g1093(.A(new_n679), .B1(new_n1293), .B2(new_n1189), .ZN(new_n1294));
  OAI21_X1  g1094(.A(new_n1151), .B1(new_n1235), .B2(new_n1180), .ZN(new_n1295));
  INV_X1    g1095(.A(KEYINPUT57), .ZN(new_n1296));
  NAND2_X1  g1096(.A1(new_n1295), .A2(new_n1296), .ZN(new_n1297));
  NAND2_X1  g1097(.A1(new_n1294), .A2(new_n1297), .ZN(new_n1298));
  AOI21_X1  g1098(.A(G378), .B1(new_n1298), .B2(new_n1179), .ZN(new_n1299));
  NAND2_X1  g1099(.A1(new_n1274), .A2(new_n1299), .ZN(new_n1300));
  AOI21_X1  g1100(.A(new_n1178), .B1(new_n1294), .B2(new_n1297), .ZN(new_n1301));
  OAI211_X1 g1101(.A(new_n1270), .B(new_n1273), .C1(new_n1301), .C2(G378), .ZN(new_n1302));
  NAND2_X1  g1102(.A1(new_n1233), .A2(KEYINPUT127), .ZN(new_n1303));
  AND3_X1   g1103(.A1(new_n1300), .A2(new_n1302), .A3(new_n1303), .ZN(new_n1304));
  AOI21_X1  g1104(.A(new_n1303), .B1(new_n1300), .B2(new_n1302), .ZN(new_n1305));
  OAI21_X1  g1105(.A(new_n1252), .B1(new_n1304), .B2(new_n1305), .ZN(new_n1306));
  INV_X1    g1106(.A(new_n1303), .ZN(new_n1307));
  NAND2_X1  g1107(.A1(G375), .A2(new_n1234), .ZN(new_n1308));
  AOI21_X1  g1108(.A(new_n1308), .B1(new_n1273), .B2(new_n1270), .ZN(new_n1309));
  NOR2_X1   g1109(.A1(new_n1274), .A2(new_n1299), .ZN(new_n1310));
  OAI21_X1  g1110(.A(new_n1307), .B1(new_n1309), .B2(new_n1310), .ZN(new_n1311));
  NAND3_X1  g1111(.A1(new_n1300), .A2(new_n1302), .A3(new_n1303), .ZN(new_n1312));
  NAND3_X1  g1112(.A1(new_n1311), .A2(new_n1282), .A3(new_n1312), .ZN(new_n1313));
  AND2_X1   g1113(.A1(new_n1306), .A2(new_n1313), .ZN(G402));
endmodule


