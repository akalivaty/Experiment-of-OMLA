//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 0 1 1 0 1 0 0 0 0 1 0 0 1 1 0 0 0 0 1 1 1 0 1 1 1 1 0 1 1 1 1 1 1 0 0 0 0 0 0 1 1 0 1 1 1 1 0 1 1 1 0 0 1 1 1 1 0 1 0 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:17:02 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n677, new_n678, new_n679,
    new_n681, new_n682, new_n683, new_n684, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n719, new_n720, new_n721, new_n722, new_n723, new_n724,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n750, new_n751, new_n752, new_n753, new_n755, new_n756,
    new_n757, new_n758, new_n759, new_n760, new_n762, new_n763, new_n764,
    new_n766, new_n767, new_n769, new_n770, new_n771, new_n772, new_n773,
    new_n774, new_n775, new_n776, new_n777, new_n778, new_n779, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n792, new_n793, new_n794, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n863,
    new_n864, new_n865, new_n867, new_n868, new_n869, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n917, new_n918, new_n919, new_n921, new_n922, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n931, new_n932, new_n933,
    new_n935, new_n936, new_n937, new_n938, new_n939, new_n940, new_n942,
    new_n943, new_n944, new_n945, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n952, new_n953, new_n954, new_n955, new_n956, new_n957,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n968, new_n969, new_n970, new_n971, new_n972, new_n974,
    new_n975, new_n976, new_n977;
  INV_X1    g000(.A(G134gat), .ZN(new_n202));
  NAND2_X1  g001(.A1(new_n202), .A2(G127gat), .ZN(new_n203));
  INV_X1    g002(.A(KEYINPUT67), .ZN(new_n204));
  NAND2_X1  g003(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  INV_X1    g004(.A(KEYINPUT68), .ZN(new_n206));
  OAI21_X1  g005(.A(new_n206), .B1(new_n202), .B2(G127gat), .ZN(new_n207));
  NAND3_X1  g006(.A1(new_n202), .A2(KEYINPUT67), .A3(G127gat), .ZN(new_n208));
  INV_X1    g007(.A(G127gat), .ZN(new_n209));
  NAND3_X1  g008(.A1(new_n209), .A2(KEYINPUT68), .A3(G134gat), .ZN(new_n210));
  NAND4_X1  g009(.A1(new_n205), .A2(new_n207), .A3(new_n208), .A4(new_n210), .ZN(new_n211));
  INV_X1    g010(.A(KEYINPUT1), .ZN(new_n212));
  INV_X1    g011(.A(G120gat), .ZN(new_n213));
  AND2_X1   g012(.A1(new_n213), .A2(G113gat), .ZN(new_n214));
  NOR2_X1   g013(.A1(new_n213), .A2(G113gat), .ZN(new_n215));
  OAI21_X1  g014(.A(new_n212), .B1(new_n214), .B2(new_n215), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n211), .A2(new_n216), .ZN(new_n217));
  XNOR2_X1  g016(.A(G127gat), .B(G134gat), .ZN(new_n218));
  OAI211_X1 g017(.A(new_n218), .B(new_n212), .C1(new_n214), .C2(new_n215), .ZN(new_n219));
  INV_X1    g018(.A(KEYINPUT69), .ZN(new_n220));
  NAND3_X1  g019(.A1(new_n217), .A2(new_n219), .A3(new_n220), .ZN(new_n221));
  INV_X1    g020(.A(new_n221), .ZN(new_n222));
  AOI21_X1  g021(.A(new_n220), .B1(new_n217), .B2(new_n219), .ZN(new_n223));
  NOR2_X1   g022(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  AND2_X1   g023(.A1(G183gat), .A2(G190gat), .ZN(new_n225));
  NOR2_X1   g024(.A1(G169gat), .A2(G176gat), .ZN(new_n226));
  INV_X1    g025(.A(new_n226), .ZN(new_n227));
  OR2_X1    g026(.A1(new_n227), .A2(KEYINPUT26), .ZN(new_n228));
  NAND2_X1  g027(.A1(G169gat), .A2(G176gat), .ZN(new_n229));
  INV_X1    g028(.A(new_n229), .ZN(new_n230));
  AOI21_X1  g029(.A(new_n230), .B1(new_n227), .B2(KEYINPUT26), .ZN(new_n231));
  AOI21_X1  g030(.A(new_n225), .B1(new_n228), .B2(new_n231), .ZN(new_n232));
  INV_X1    g031(.A(new_n232), .ZN(new_n233));
  INV_X1    g032(.A(KEYINPUT66), .ZN(new_n234));
  INV_X1    g033(.A(KEYINPUT65), .ZN(new_n235));
  NAND2_X1  g034(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n236));
  INV_X1    g035(.A(new_n236), .ZN(new_n237));
  NOR2_X1   g036(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n238));
  OAI21_X1  g037(.A(new_n235), .B1(new_n237), .B2(new_n238), .ZN(new_n239));
  INV_X1    g038(.A(KEYINPUT27), .ZN(new_n240));
  INV_X1    g039(.A(G183gat), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n240), .A2(new_n241), .ZN(new_n242));
  NAND3_X1  g041(.A1(new_n242), .A2(KEYINPUT65), .A3(new_n236), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n239), .A2(new_n243), .ZN(new_n244));
  INV_X1    g043(.A(KEYINPUT28), .ZN(new_n245));
  NOR2_X1   g044(.A1(new_n245), .A2(G190gat), .ZN(new_n246));
  AOI21_X1  g045(.A(new_n234), .B1(new_n244), .B2(new_n246), .ZN(new_n247));
  INV_X1    g046(.A(new_n246), .ZN(new_n248));
  AOI211_X1 g047(.A(KEYINPUT66), .B(new_n248), .C1(new_n239), .C2(new_n243), .ZN(new_n249));
  NOR2_X1   g048(.A1(new_n247), .A2(new_n249), .ZN(new_n250));
  INV_X1    g049(.A(G190gat), .ZN(new_n251));
  OAI21_X1  g050(.A(new_n251), .B1(new_n237), .B2(new_n238), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n252), .A2(new_n245), .ZN(new_n253));
  AOI21_X1  g052(.A(new_n233), .B1(new_n250), .B2(new_n253), .ZN(new_n254));
  NAND2_X1  g053(.A1(new_n241), .A2(new_n251), .ZN(new_n255));
  INV_X1    g054(.A(KEYINPUT24), .ZN(new_n256));
  NAND2_X1  g055(.A1(new_n256), .A2(KEYINPUT64), .ZN(new_n257));
  NAND2_X1  g056(.A1(G183gat), .A2(G190gat), .ZN(new_n258));
  NAND3_X1  g057(.A1(new_n255), .A2(new_n257), .A3(new_n258), .ZN(new_n259));
  OAI21_X1  g058(.A(new_n259), .B1(new_n257), .B2(new_n258), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n229), .A2(KEYINPUT23), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n227), .A2(new_n261), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n226), .A2(KEYINPUT23), .ZN(new_n263));
  NAND2_X1  g062(.A1(new_n262), .A2(new_n263), .ZN(new_n264));
  OAI21_X1  g063(.A(KEYINPUT25), .B1(new_n260), .B2(new_n264), .ZN(new_n265));
  NOR2_X1   g064(.A1(G183gat), .A2(G190gat), .ZN(new_n266));
  NOR2_X1   g065(.A1(new_n225), .A2(new_n266), .ZN(new_n267));
  AOI21_X1  g066(.A(KEYINPUT25), .B1(new_n267), .B2(KEYINPUT24), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n225), .A2(new_n256), .ZN(new_n269));
  NAND4_X1  g068(.A1(new_n268), .A2(new_n263), .A3(new_n262), .A4(new_n269), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n265), .A2(new_n270), .ZN(new_n271));
  OAI211_X1 g070(.A(KEYINPUT70), .B(new_n224), .C1(new_n254), .C2(new_n271), .ZN(new_n272));
  INV_X1    g071(.A(KEYINPUT70), .ZN(new_n273));
  NOR3_X1   g072(.A1(new_n237), .A2(new_n238), .A3(new_n235), .ZN(new_n274));
  AOI21_X1  g073(.A(KEYINPUT65), .B1(new_n242), .B2(new_n236), .ZN(new_n275));
  OAI21_X1  g074(.A(new_n246), .B1(new_n274), .B2(new_n275), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n276), .A2(KEYINPUT66), .ZN(new_n277));
  NAND3_X1  g076(.A1(new_n244), .A2(new_n234), .A3(new_n246), .ZN(new_n278));
  NAND3_X1  g077(.A1(new_n277), .A2(new_n253), .A3(new_n278), .ZN(new_n279));
  AOI21_X1  g078(.A(new_n271), .B1(new_n279), .B2(new_n232), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n217), .A2(new_n219), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n281), .A2(KEYINPUT69), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n282), .A2(new_n221), .ZN(new_n283));
  OAI21_X1  g082(.A(new_n273), .B1(new_n280), .B2(new_n283), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n280), .A2(new_n283), .ZN(new_n285));
  NAND3_X1  g084(.A1(new_n272), .A2(new_n284), .A3(new_n285), .ZN(new_n286));
  NAND2_X1  g085(.A1(G227gat), .A2(G233gat), .ZN(new_n287));
  INV_X1    g086(.A(new_n287), .ZN(new_n288));
  AND3_X1   g087(.A1(new_n286), .A2(KEYINPUT71), .A3(new_n288), .ZN(new_n289));
  AOI21_X1  g088(.A(KEYINPUT71), .B1(new_n286), .B2(new_n288), .ZN(new_n290));
  OAI21_X1  g089(.A(KEYINPUT32), .B1(new_n289), .B2(new_n290), .ZN(new_n291));
  INV_X1    g090(.A(KEYINPUT33), .ZN(new_n292));
  OAI21_X1  g091(.A(new_n292), .B1(new_n289), .B2(new_n290), .ZN(new_n293));
  XNOR2_X1  g092(.A(G15gat), .B(G43gat), .ZN(new_n294));
  XNOR2_X1  g093(.A(new_n294), .B(G71gat), .ZN(new_n295));
  INV_X1    g094(.A(G99gat), .ZN(new_n296));
  XNOR2_X1  g095(.A(new_n295), .B(new_n296), .ZN(new_n297));
  NAND3_X1  g096(.A1(new_n291), .A2(new_n293), .A3(new_n297), .ZN(new_n298));
  INV_X1    g097(.A(new_n297), .ZN(new_n299));
  OAI221_X1 g098(.A(KEYINPUT32), .B1(new_n292), .B2(new_n299), .C1(new_n289), .C2(new_n290), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n298), .A2(new_n300), .ZN(new_n301));
  NAND4_X1  g100(.A1(new_n272), .A2(new_n284), .A3(new_n287), .A4(new_n285), .ZN(new_n302));
  OR3_X1    g101(.A1(new_n302), .A2(KEYINPUT72), .A3(KEYINPUT73), .ZN(new_n303));
  AOI21_X1  g102(.A(KEYINPUT34), .B1(new_n302), .B2(KEYINPUT72), .ZN(new_n304));
  OAI21_X1  g103(.A(KEYINPUT73), .B1(new_n302), .B2(KEYINPUT72), .ZN(new_n305));
  AND3_X1   g104(.A1(new_n303), .A2(new_n304), .A3(new_n305), .ZN(new_n306));
  AOI21_X1  g105(.A(new_n304), .B1(new_n303), .B2(new_n305), .ZN(new_n307));
  NOR2_X1   g106(.A1(new_n306), .A2(new_n307), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n301), .A2(new_n308), .ZN(new_n309));
  INV_X1    g108(.A(KEYINPUT74), .ZN(new_n310));
  OAI211_X1 g109(.A(new_n298), .B(new_n300), .C1(new_n306), .C2(new_n307), .ZN(new_n311));
  NAND3_X1  g110(.A1(new_n309), .A2(new_n310), .A3(new_n311), .ZN(new_n312));
  NAND3_X1  g111(.A1(new_n301), .A2(new_n308), .A3(KEYINPUT74), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  NAND2_X1  g113(.A1(G228gat), .A2(G233gat), .ZN(new_n315));
  INV_X1    g114(.A(new_n315), .ZN(new_n316));
  XNOR2_X1  g115(.A(G141gat), .B(G148gat), .ZN(new_n317));
  INV_X1    g116(.A(new_n317), .ZN(new_n318));
  INV_X1    g117(.A(G162gat), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n319), .A2(G155gat), .ZN(new_n320));
  INV_X1    g119(.A(G155gat), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n321), .A2(G162gat), .ZN(new_n322));
  AND2_X1   g121(.A1(new_n320), .A2(new_n322), .ZN(new_n323));
  AND2_X1   g122(.A1(KEYINPUT80), .A2(G155gat), .ZN(new_n324));
  NOR2_X1   g123(.A1(KEYINPUT80), .A2(G155gat), .ZN(new_n325));
  NOR3_X1   g124(.A1(new_n324), .A2(new_n325), .A3(new_n319), .ZN(new_n326));
  INV_X1    g125(.A(KEYINPUT2), .ZN(new_n327));
  OAI211_X1 g126(.A(new_n318), .B(new_n323), .C1(new_n326), .C2(new_n327), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n328), .A2(KEYINPUT81), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n320), .A2(new_n322), .ZN(new_n330));
  XNOR2_X1  g129(.A(KEYINPUT79), .B(KEYINPUT2), .ZN(new_n331));
  OAI21_X1  g130(.A(new_n330), .B1(new_n317), .B2(new_n331), .ZN(new_n332));
  OR2_X1    g131(.A1(KEYINPUT80), .A2(G155gat), .ZN(new_n333));
  NAND2_X1  g132(.A1(KEYINPUT80), .A2(G155gat), .ZN(new_n334));
  NAND3_X1  g133(.A1(new_n333), .A2(G162gat), .A3(new_n334), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n335), .A2(KEYINPUT2), .ZN(new_n336));
  INV_X1    g135(.A(KEYINPUT81), .ZN(new_n337));
  NAND4_X1  g136(.A1(new_n336), .A2(new_n337), .A3(new_n323), .A4(new_n318), .ZN(new_n338));
  NAND3_X1  g137(.A1(new_n329), .A2(new_n332), .A3(new_n338), .ZN(new_n339));
  OR2_X1    g138(.A1(KEYINPUT75), .A2(KEYINPUT22), .ZN(new_n340));
  NAND2_X1  g139(.A1(G211gat), .A2(G218gat), .ZN(new_n341));
  NAND2_X1  g140(.A1(KEYINPUT75), .A2(KEYINPUT22), .ZN(new_n342));
  NAND3_X1  g141(.A1(new_n340), .A2(new_n341), .A3(new_n342), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n343), .A2(KEYINPUT76), .ZN(new_n344));
  XNOR2_X1  g143(.A(G197gat), .B(G204gat), .ZN(new_n345));
  INV_X1    g144(.A(KEYINPUT76), .ZN(new_n346));
  NAND4_X1  g145(.A1(new_n340), .A2(new_n346), .A3(new_n341), .A4(new_n342), .ZN(new_n347));
  NAND3_X1  g146(.A1(new_n344), .A2(new_n345), .A3(new_n347), .ZN(new_n348));
  XNOR2_X1  g147(.A(G211gat), .B(G218gat), .ZN(new_n349));
  INV_X1    g148(.A(new_n349), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n348), .A2(new_n350), .ZN(new_n351));
  NAND4_X1  g150(.A1(new_n344), .A2(new_n349), .A3(new_n345), .A4(new_n347), .ZN(new_n352));
  AOI21_X1  g151(.A(KEYINPUT29), .B1(new_n351), .B2(new_n352), .ZN(new_n353));
  OAI21_X1  g152(.A(new_n339), .B1(new_n353), .B2(KEYINPUT3), .ZN(new_n354));
  XOR2_X1   g153(.A(KEYINPUT77), .B(KEYINPUT29), .Z(new_n355));
  INV_X1    g154(.A(new_n338), .ZN(new_n356));
  AOI21_X1  g155(.A(new_n330), .B1(new_n335), .B2(KEYINPUT2), .ZN(new_n357));
  AOI21_X1  g156(.A(new_n337), .B1(new_n357), .B2(new_n318), .ZN(new_n358));
  NOR2_X1   g157(.A1(new_n356), .A2(new_n358), .ZN(new_n359));
  INV_X1    g158(.A(KEYINPUT3), .ZN(new_n360));
  NAND4_X1  g159(.A1(new_n359), .A2(KEYINPUT82), .A3(new_n360), .A4(new_n332), .ZN(new_n361));
  NAND4_X1  g160(.A1(new_n329), .A2(new_n360), .A3(new_n332), .A4(new_n338), .ZN(new_n362));
  INV_X1    g161(.A(KEYINPUT82), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n362), .A2(new_n363), .ZN(new_n364));
  AOI21_X1  g163(.A(new_n355), .B1(new_n361), .B2(new_n364), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n351), .A2(new_n352), .ZN(new_n366));
  OAI211_X1 g165(.A(new_n316), .B(new_n354), .C1(new_n365), .C2(new_n366), .ZN(new_n367));
  AND3_X1   g166(.A1(new_n329), .A2(new_n332), .A3(new_n338), .ZN(new_n368));
  INV_X1    g167(.A(new_n355), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n366), .A2(new_n369), .ZN(new_n370));
  AOI21_X1  g169(.A(new_n368), .B1(new_n370), .B2(new_n360), .ZN(new_n371));
  AND2_X1   g170(.A1(new_n362), .A2(new_n363), .ZN(new_n372));
  NOR2_X1   g171(.A1(new_n362), .A2(new_n363), .ZN(new_n373));
  OAI21_X1  g172(.A(new_n369), .B1(new_n372), .B2(new_n373), .ZN(new_n374));
  INV_X1    g173(.A(new_n366), .ZN(new_n375));
  AOI21_X1  g174(.A(new_n371), .B1(new_n374), .B2(new_n375), .ZN(new_n376));
  OAI21_X1  g175(.A(new_n367), .B1(new_n376), .B2(new_n316), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n377), .A2(G22gat), .ZN(new_n378));
  INV_X1    g177(.A(G22gat), .ZN(new_n379));
  OAI211_X1 g178(.A(new_n367), .B(new_n379), .C1(new_n376), .C2(new_n316), .ZN(new_n380));
  NAND3_X1  g179(.A1(new_n378), .A2(KEYINPUT85), .A3(new_n380), .ZN(new_n381));
  OR2_X1    g180(.A1(new_n380), .A2(KEYINPUT85), .ZN(new_n382));
  XNOR2_X1  g181(.A(G78gat), .B(G106gat), .ZN(new_n383));
  XNOR2_X1  g182(.A(KEYINPUT31), .B(G50gat), .ZN(new_n384));
  XNOR2_X1  g183(.A(new_n383), .B(new_n384), .ZN(new_n385));
  INV_X1    g184(.A(new_n385), .ZN(new_n386));
  NAND3_X1  g185(.A1(new_n381), .A2(new_n382), .A3(new_n386), .ZN(new_n387));
  INV_X1    g186(.A(KEYINPUT88), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n378), .A2(KEYINPUT86), .ZN(new_n389));
  INV_X1    g188(.A(KEYINPUT86), .ZN(new_n390));
  NAND3_X1  g189(.A1(new_n377), .A2(new_n390), .A3(G22gat), .ZN(new_n391));
  AOI21_X1  g190(.A(new_n386), .B1(new_n389), .B2(new_n391), .ZN(new_n392));
  XOR2_X1   g191(.A(new_n380), .B(KEYINPUT87), .Z(new_n393));
  AOI21_X1  g192(.A(new_n388), .B1(new_n392), .B2(new_n393), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n361), .A2(new_n364), .ZN(new_n395));
  AOI21_X1  g194(.A(new_n366), .B1(new_n395), .B2(new_n369), .ZN(new_n396));
  OAI21_X1  g195(.A(new_n315), .B1(new_n396), .B2(new_n371), .ZN(new_n397));
  AOI211_X1 g196(.A(KEYINPUT86), .B(new_n379), .C1(new_n397), .C2(new_n367), .ZN(new_n398));
  AOI21_X1  g197(.A(new_n390), .B1(new_n377), .B2(G22gat), .ZN(new_n399));
  OAI21_X1  g198(.A(new_n385), .B1(new_n398), .B2(new_n399), .ZN(new_n400));
  XNOR2_X1  g199(.A(new_n380), .B(KEYINPUT87), .ZN(new_n401));
  NOR3_X1   g200(.A1(new_n400), .A2(new_n401), .A3(KEYINPUT88), .ZN(new_n402));
  OAI21_X1  g201(.A(new_n387), .B1(new_n394), .B2(new_n402), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n314), .A2(new_n403), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n404), .A2(KEYINPUT93), .ZN(new_n405));
  INV_X1    g204(.A(KEYINPUT93), .ZN(new_n406));
  NAND3_X1  g205(.A1(new_n314), .A2(new_n406), .A3(new_n403), .ZN(new_n407));
  INV_X1    g206(.A(G226gat), .ZN(new_n408));
  INV_X1    g207(.A(G233gat), .ZN(new_n409));
  NOR2_X1   g208(.A1(new_n408), .A2(new_n409), .ZN(new_n410));
  INV_X1    g209(.A(new_n410), .ZN(new_n411));
  OAI21_X1  g210(.A(new_n411), .B1(new_n280), .B2(KEYINPUT29), .ZN(new_n412));
  OAI21_X1  g211(.A(new_n410), .B1(new_n254), .B2(new_n271), .ZN(new_n413));
  NAND3_X1  g212(.A1(new_n412), .A2(new_n413), .A3(KEYINPUT78), .ZN(new_n414));
  OR3_X1    g213(.A1(new_n280), .A2(KEYINPUT78), .A3(new_n411), .ZN(new_n415));
  NAND3_X1  g214(.A1(new_n414), .A2(new_n415), .A3(new_n366), .ZN(new_n416));
  OAI21_X1  g215(.A(new_n411), .B1(new_n280), .B2(new_n355), .ZN(new_n417));
  NAND3_X1  g216(.A1(new_n417), .A2(new_n413), .A3(new_n375), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n416), .A2(new_n418), .ZN(new_n419));
  XNOR2_X1  g218(.A(G8gat), .B(G36gat), .ZN(new_n420));
  XNOR2_X1  g219(.A(G64gat), .B(G92gat), .ZN(new_n421));
  XNOR2_X1  g220(.A(new_n420), .B(new_n421), .ZN(new_n422));
  INV_X1    g221(.A(new_n422), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n419), .A2(new_n423), .ZN(new_n424));
  INV_X1    g223(.A(new_n424), .ZN(new_n425));
  OAI21_X1  g224(.A(KEYINPUT30), .B1(new_n419), .B2(new_n423), .ZN(new_n426));
  XNOR2_X1  g225(.A(new_n425), .B(new_n426), .ZN(new_n427));
  XNOR2_X1  g226(.A(G1gat), .B(G29gat), .ZN(new_n428));
  XNOR2_X1  g227(.A(new_n428), .B(G85gat), .ZN(new_n429));
  XNOR2_X1  g228(.A(KEYINPUT0), .B(G57gat), .ZN(new_n430));
  XOR2_X1   g229(.A(new_n429), .B(new_n430), .Z(new_n431));
  NAND2_X1  g230(.A1(G225gat), .A2(G233gat), .ZN(new_n432));
  XNOR2_X1  g231(.A(new_n432), .B(KEYINPUT83), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n339), .A2(KEYINPUT3), .ZN(new_n434));
  OAI211_X1 g233(.A(new_n434), .B(new_n281), .C1(new_n372), .C2(new_n373), .ZN(new_n435));
  INV_X1    g234(.A(KEYINPUT4), .ZN(new_n436));
  NOR3_X1   g235(.A1(new_n339), .A2(new_n436), .A3(new_n281), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n283), .A2(new_n368), .ZN(new_n438));
  AOI21_X1  g237(.A(new_n437), .B1(new_n436), .B2(new_n438), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n435), .A2(new_n439), .ZN(new_n440));
  INV_X1    g239(.A(KEYINPUT5), .ZN(new_n441));
  AOI21_X1  g240(.A(new_n433), .B1(new_n440), .B2(new_n441), .ZN(new_n442));
  OAI21_X1  g241(.A(KEYINPUT4), .B1(new_n224), .B2(new_n339), .ZN(new_n443));
  INV_X1    g242(.A(KEYINPUT84), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n443), .A2(new_n444), .ZN(new_n445));
  NAND3_X1  g244(.A1(new_n438), .A2(KEYINPUT84), .A3(KEYINPUT4), .ZN(new_n446));
  NAND4_X1  g245(.A1(new_n368), .A2(new_n436), .A3(new_n217), .A4(new_n219), .ZN(new_n447));
  NAND3_X1  g246(.A1(new_n445), .A2(new_n446), .A3(new_n447), .ZN(new_n448));
  NAND3_X1  g247(.A1(new_n448), .A2(KEYINPUT5), .A3(new_n435), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n442), .A2(new_n449), .ZN(new_n450));
  XNOR2_X1  g249(.A(new_n339), .B(new_n281), .ZN(new_n451));
  INV_X1    g250(.A(new_n433), .ZN(new_n452));
  NOR3_X1   g251(.A1(new_n451), .A2(new_n441), .A3(new_n452), .ZN(new_n453));
  INV_X1    g252(.A(new_n453), .ZN(new_n454));
  AOI21_X1  g253(.A(new_n431), .B1(new_n450), .B2(new_n454), .ZN(new_n455));
  INV_X1    g254(.A(new_n455), .ZN(new_n456));
  AOI21_X1  g255(.A(new_n453), .B1(new_n442), .B2(new_n449), .ZN(new_n457));
  AOI21_X1  g256(.A(KEYINPUT6), .B1(new_n457), .B2(new_n431), .ZN(new_n458));
  AND2_X1   g257(.A1(new_n456), .A2(new_n458), .ZN(new_n459));
  NOR2_X1   g258(.A1(new_n456), .A2(new_n458), .ZN(new_n460));
  OAI21_X1  g259(.A(new_n427), .B1(new_n459), .B2(new_n460), .ZN(new_n461));
  INV_X1    g260(.A(new_n461), .ZN(new_n462));
  NAND3_X1  g261(.A1(new_n405), .A2(new_n407), .A3(new_n462), .ZN(new_n463));
  INV_X1    g262(.A(new_n431), .ZN(new_n464));
  INV_X1    g263(.A(KEYINPUT90), .ZN(new_n465));
  NOR2_X1   g264(.A1(new_n457), .A2(new_n465), .ZN(new_n466));
  AOI211_X1 g265(.A(KEYINPUT90), .B(new_n453), .C1(new_n442), .C2(new_n449), .ZN(new_n467));
  OAI21_X1  g266(.A(new_n464), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n468), .A2(new_n458), .ZN(new_n469));
  AOI21_X1  g268(.A(KEYINPUT91), .B1(new_n455), .B2(KEYINPUT6), .ZN(new_n470));
  INV_X1    g269(.A(KEYINPUT91), .ZN(new_n471));
  INV_X1    g270(.A(KEYINPUT6), .ZN(new_n472));
  NOR4_X1   g271(.A1(new_n457), .A2(new_n471), .A3(new_n472), .A4(new_n431), .ZN(new_n473));
  NOR2_X1   g272(.A1(new_n470), .A2(new_n473), .ZN(new_n474));
  AOI21_X1  g273(.A(KEYINPUT35), .B1(new_n469), .B2(new_n474), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n309), .A2(new_n311), .ZN(new_n476));
  INV_X1    g275(.A(new_n476), .ZN(new_n477));
  NAND4_X1  g276(.A1(new_n475), .A2(new_n403), .A3(new_n477), .A4(new_n427), .ZN(new_n478));
  INV_X1    g277(.A(KEYINPUT92), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  INV_X1    g279(.A(new_n387), .ZN(new_n481));
  NAND3_X1  g280(.A1(new_n392), .A2(new_n393), .A3(new_n388), .ZN(new_n482));
  OAI21_X1  g281(.A(KEYINPUT88), .B1(new_n400), .B2(new_n401), .ZN(new_n483));
  AOI21_X1  g282(.A(new_n481), .B1(new_n482), .B2(new_n483), .ZN(new_n484));
  NOR2_X1   g283(.A1(new_n484), .A2(new_n476), .ZN(new_n485));
  NAND4_X1  g284(.A1(new_n485), .A2(KEYINPUT92), .A3(new_n475), .A4(new_n427), .ZN(new_n486));
  AOI22_X1  g285(.A1(new_n463), .A2(KEYINPUT35), .B1(new_n480), .B2(new_n486), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n484), .A2(new_n461), .ZN(new_n488));
  NAND3_X1  g287(.A1(new_n312), .A2(KEYINPUT36), .A3(new_n313), .ZN(new_n489));
  INV_X1    g288(.A(KEYINPUT36), .ZN(new_n490));
  NAND3_X1  g289(.A1(new_n309), .A2(new_n490), .A3(new_n311), .ZN(new_n491));
  NAND3_X1  g290(.A1(new_n488), .A2(new_n489), .A3(new_n491), .ZN(new_n492));
  AOI21_X1  g291(.A(new_n375), .B1(new_n417), .B2(new_n413), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n414), .A2(new_n415), .ZN(new_n494));
  AOI21_X1  g293(.A(new_n493), .B1(new_n494), .B2(new_n375), .ZN(new_n495));
  AOI21_X1  g294(.A(KEYINPUT38), .B1(new_n495), .B2(KEYINPUT37), .ZN(new_n496));
  INV_X1    g295(.A(KEYINPUT37), .ZN(new_n497));
  AOI21_X1  g296(.A(new_n423), .B1(new_n419), .B2(new_n497), .ZN(new_n498));
  AOI21_X1  g297(.A(new_n425), .B1(new_n496), .B2(new_n498), .ZN(new_n499));
  NAND3_X1  g298(.A1(new_n416), .A2(KEYINPUT37), .A3(new_n418), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n498), .A2(new_n500), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n501), .A2(KEYINPUT38), .ZN(new_n502));
  AND2_X1   g301(.A1(new_n499), .A2(new_n502), .ZN(new_n503));
  NAND3_X1  g302(.A1(new_n503), .A2(new_n469), .A3(new_n474), .ZN(new_n504));
  NAND3_X1  g303(.A1(new_n451), .A2(KEYINPUT39), .A3(new_n452), .ZN(new_n505));
  XNOR2_X1  g304(.A(new_n440), .B(KEYINPUT39), .ZN(new_n506));
  OAI211_X1 g305(.A(new_n431), .B(new_n505), .C1(new_n506), .C2(new_n452), .ZN(new_n507));
  INV_X1    g306(.A(KEYINPUT40), .ZN(new_n508));
  OAI21_X1  g307(.A(new_n507), .B1(KEYINPUT89), .B2(new_n508), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n508), .A2(KEYINPUT89), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  XNOR2_X1  g310(.A(new_n426), .B(new_n424), .ZN(new_n512));
  NAND3_X1  g311(.A1(new_n507), .A2(KEYINPUT89), .A3(new_n508), .ZN(new_n513));
  NAND4_X1  g312(.A1(new_n511), .A2(new_n512), .A3(new_n468), .A4(new_n513), .ZN(new_n514));
  AND3_X1   g313(.A1(new_n403), .A2(new_n504), .A3(new_n514), .ZN(new_n515));
  NOR2_X1   g314(.A1(new_n492), .A2(new_n515), .ZN(new_n516));
  NOR2_X1   g315(.A1(new_n487), .A2(new_n516), .ZN(new_n517));
  XNOR2_X1  g316(.A(G15gat), .B(G22gat), .ZN(new_n518));
  INV_X1    g317(.A(KEYINPUT16), .ZN(new_n519));
  AOI21_X1  g318(.A(G1gat), .B1(new_n518), .B2(new_n519), .ZN(new_n520));
  INV_X1    g319(.A(G8gat), .ZN(new_n521));
  XNOR2_X1  g320(.A(new_n520), .B(new_n521), .ZN(new_n522));
  AND2_X1   g321(.A1(new_n518), .A2(KEYINPUT96), .ZN(new_n523));
  XNOR2_X1  g322(.A(new_n522), .B(new_n523), .ZN(new_n524));
  INV_X1    g323(.A(new_n524), .ZN(new_n525));
  OR2_X1    g324(.A1(G29gat), .A2(G36gat), .ZN(new_n526));
  XNOR2_X1  g325(.A(new_n526), .B(KEYINPUT14), .ZN(new_n527));
  INV_X1    g326(.A(G29gat), .ZN(new_n528));
  XOR2_X1   g327(.A(KEYINPUT95), .B(G36gat), .Z(new_n529));
  OAI21_X1  g328(.A(new_n527), .B1(new_n528), .B2(new_n529), .ZN(new_n530));
  XNOR2_X1  g329(.A(G43gat), .B(G50gat), .ZN(new_n531));
  AND2_X1   g330(.A1(new_n531), .A2(KEYINPUT15), .ZN(new_n532));
  NOR2_X1   g331(.A1(new_n531), .A2(KEYINPUT15), .ZN(new_n533));
  OR3_X1    g332(.A1(new_n530), .A2(new_n532), .A3(new_n533), .ZN(new_n534));
  NAND3_X1  g333(.A1(new_n530), .A2(KEYINPUT15), .A3(new_n531), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  NOR2_X1   g335(.A1(KEYINPUT97), .A2(KEYINPUT17), .ZN(new_n537));
  AND2_X1   g336(.A1(KEYINPUT97), .A2(KEYINPUT17), .ZN(new_n538));
  NOR3_X1   g337(.A1(new_n536), .A2(new_n537), .A3(new_n538), .ZN(new_n539));
  AND2_X1   g338(.A1(new_n536), .A2(new_n538), .ZN(new_n540));
  OAI21_X1  g339(.A(new_n525), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n524), .A2(new_n536), .ZN(new_n542));
  NAND2_X1  g341(.A1(G229gat), .A2(G233gat), .ZN(new_n543));
  NAND3_X1  g342(.A1(new_n541), .A2(new_n542), .A3(new_n543), .ZN(new_n544));
  INV_X1    g343(.A(KEYINPUT18), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  XNOR2_X1  g345(.A(new_n524), .B(new_n536), .ZN(new_n547));
  XOR2_X1   g346(.A(new_n543), .B(KEYINPUT13), .Z(new_n548));
  NAND2_X1  g347(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  NAND4_X1  g348(.A1(new_n541), .A2(KEYINPUT18), .A3(new_n542), .A4(new_n543), .ZN(new_n550));
  NAND3_X1  g349(.A1(new_n546), .A2(new_n549), .A3(new_n550), .ZN(new_n551));
  XNOR2_X1  g350(.A(G113gat), .B(G141gat), .ZN(new_n552));
  XNOR2_X1  g351(.A(new_n552), .B(G197gat), .ZN(new_n553));
  XOR2_X1   g352(.A(KEYINPUT11), .B(G169gat), .Z(new_n554));
  XNOR2_X1  g353(.A(new_n553), .B(new_n554), .ZN(new_n555));
  XOR2_X1   g354(.A(new_n555), .B(KEYINPUT94), .Z(new_n556));
  XOR2_X1   g355(.A(new_n556), .B(KEYINPUT12), .Z(new_n557));
  INV_X1    g356(.A(new_n557), .ZN(new_n558));
  NAND2_X1  g357(.A1(new_n551), .A2(new_n558), .ZN(new_n559));
  NAND4_X1  g358(.A1(new_n546), .A2(new_n557), .A3(new_n549), .A4(new_n550), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  INV_X1    g360(.A(new_n561), .ZN(new_n562));
  NOR2_X1   g361(.A1(new_n517), .A2(new_n562), .ZN(new_n563));
  XOR2_X1   g362(.A(G71gat), .B(G78gat), .Z(new_n564));
  NAND2_X1  g363(.A1(new_n564), .A2(KEYINPUT98), .ZN(new_n565));
  XOR2_X1   g364(.A(G57gat), .B(G64gat), .Z(new_n566));
  INV_X1    g365(.A(KEYINPUT9), .ZN(new_n567));
  INV_X1    g366(.A(G71gat), .ZN(new_n568));
  INV_X1    g367(.A(G78gat), .ZN(new_n569));
  OAI21_X1  g368(.A(new_n567), .B1(new_n568), .B2(new_n569), .ZN(new_n570));
  XNOR2_X1  g369(.A(G71gat), .B(G78gat), .ZN(new_n571));
  INV_X1    g370(.A(KEYINPUT98), .ZN(new_n572));
  NAND2_X1  g371(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  NAND4_X1  g372(.A1(new_n565), .A2(new_n566), .A3(new_n570), .A4(new_n573), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n566), .A2(KEYINPUT9), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n575), .A2(new_n564), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n574), .A2(new_n576), .ZN(new_n577));
  NOR2_X1   g376(.A1(new_n577), .A2(KEYINPUT99), .ZN(new_n578));
  INV_X1    g377(.A(KEYINPUT99), .ZN(new_n579));
  AOI21_X1  g378(.A(new_n579), .B1(new_n574), .B2(new_n576), .ZN(new_n580));
  OR2_X1    g379(.A1(new_n578), .A2(new_n580), .ZN(new_n581));
  AOI21_X1  g380(.A(new_n524), .B1(new_n581), .B2(KEYINPUT21), .ZN(new_n582));
  XNOR2_X1  g381(.A(new_n582), .B(KEYINPUT100), .ZN(new_n583));
  XNOR2_X1  g382(.A(new_n583), .B(G127gat), .ZN(new_n584));
  INV_X1    g383(.A(new_n584), .ZN(new_n585));
  NOR2_X1   g384(.A1(new_n581), .A2(KEYINPUT21), .ZN(new_n586));
  XOR2_X1   g385(.A(G183gat), .B(G211gat), .Z(new_n587));
  XNOR2_X1  g386(.A(new_n586), .B(new_n587), .ZN(new_n588));
  NAND2_X1  g387(.A1(G231gat), .A2(G233gat), .ZN(new_n589));
  XNOR2_X1  g388(.A(new_n588), .B(new_n589), .ZN(new_n590));
  NAND2_X1  g389(.A1(new_n585), .A2(new_n590), .ZN(new_n591));
  INV_X1    g390(.A(new_n590), .ZN(new_n592));
  NAND2_X1  g391(.A1(new_n592), .A2(new_n584), .ZN(new_n593));
  NAND2_X1  g392(.A1(new_n591), .A2(new_n593), .ZN(new_n594));
  XNOR2_X1  g393(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n595));
  XNOR2_X1  g394(.A(new_n595), .B(G155gat), .ZN(new_n596));
  INV_X1    g395(.A(new_n596), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n594), .A2(new_n597), .ZN(new_n598));
  INV_X1    g397(.A(KEYINPUT101), .ZN(new_n599));
  INV_X1    g398(.A(KEYINPUT7), .ZN(new_n600));
  NAND2_X1  g399(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  NAND2_X1  g400(.A1(KEYINPUT101), .A2(KEYINPUT7), .ZN(new_n602));
  NAND4_X1  g401(.A1(new_n601), .A2(G85gat), .A3(G92gat), .A4(new_n602), .ZN(new_n603));
  NAND2_X1  g402(.A1(G99gat), .A2(G106gat), .ZN(new_n604));
  INV_X1    g403(.A(G85gat), .ZN(new_n605));
  INV_X1    g404(.A(G92gat), .ZN(new_n606));
  AOI22_X1  g405(.A1(KEYINPUT8), .A2(new_n604), .B1(new_n605), .B2(new_n606), .ZN(new_n607));
  OAI211_X1 g406(.A(new_n599), .B(new_n600), .C1(new_n605), .C2(new_n606), .ZN(new_n608));
  NAND3_X1  g407(.A1(new_n603), .A2(new_n607), .A3(new_n608), .ZN(new_n609));
  XNOR2_X1  g408(.A(G99gat), .B(G106gat), .ZN(new_n610));
  INV_X1    g409(.A(new_n610), .ZN(new_n611));
  OR2_X1    g410(.A1(new_n609), .A2(new_n611), .ZN(new_n612));
  NAND2_X1  g411(.A1(new_n609), .A2(new_n611), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  OAI21_X1  g413(.A(new_n614), .B1(new_n539), .B2(new_n540), .ZN(new_n615));
  NAND3_X1  g414(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n616));
  INV_X1    g415(.A(new_n614), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n536), .A2(new_n617), .ZN(new_n618));
  NAND3_X1  g417(.A1(new_n615), .A2(new_n616), .A3(new_n618), .ZN(new_n619));
  XNOR2_X1  g418(.A(G190gat), .B(G218gat), .ZN(new_n620));
  AND2_X1   g419(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  NOR2_X1   g420(.A1(new_n619), .A2(new_n620), .ZN(new_n622));
  XNOR2_X1  g421(.A(G134gat), .B(G162gat), .ZN(new_n623));
  AOI21_X1  g422(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n624));
  XOR2_X1   g423(.A(new_n623), .B(new_n624), .Z(new_n625));
  INV_X1    g424(.A(new_n625), .ZN(new_n626));
  OR3_X1    g425(.A1(new_n621), .A2(new_n622), .A3(new_n626), .ZN(new_n627));
  OAI21_X1  g426(.A(new_n626), .B1(new_n621), .B2(new_n622), .ZN(new_n628));
  NAND2_X1  g427(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  NAND3_X1  g428(.A1(new_n591), .A2(new_n596), .A3(new_n593), .ZN(new_n630));
  NAND3_X1  g429(.A1(new_n598), .A2(new_n629), .A3(new_n630), .ZN(new_n631));
  INV_X1    g430(.A(KEYINPUT102), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  NAND4_X1  g432(.A1(new_n598), .A2(new_n629), .A3(KEYINPUT102), .A4(new_n630), .ZN(new_n634));
  AND2_X1   g433(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  NAND3_X1  g434(.A1(new_n581), .A2(KEYINPUT10), .A3(new_n617), .ZN(new_n636));
  OAI21_X1  g435(.A(new_n614), .B1(new_n578), .B2(new_n580), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n617), .A2(new_n577), .ZN(new_n638));
  NAND2_X1  g437(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  INV_X1    g438(.A(KEYINPUT10), .ZN(new_n640));
  AOI21_X1  g439(.A(KEYINPUT103), .B1(new_n639), .B2(new_n640), .ZN(new_n641));
  INV_X1    g440(.A(KEYINPUT103), .ZN(new_n642));
  AOI211_X1 g441(.A(new_n642), .B(KEYINPUT10), .C1(new_n637), .C2(new_n638), .ZN(new_n643));
  OAI21_X1  g442(.A(new_n636), .B1(new_n641), .B2(new_n643), .ZN(new_n644));
  NAND2_X1  g443(.A1(G230gat), .A2(G233gat), .ZN(new_n645));
  NAND2_X1  g444(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  INV_X1    g445(.A(KEYINPUT104), .ZN(new_n647));
  NAND2_X1  g446(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  NAND3_X1  g447(.A1(new_n644), .A2(KEYINPUT104), .A3(new_n645), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  XNOR2_X1  g449(.A(G120gat), .B(G148gat), .ZN(new_n651));
  XNOR2_X1  g450(.A(G176gat), .B(G204gat), .ZN(new_n652));
  XNOR2_X1  g451(.A(new_n651), .B(new_n652), .ZN(new_n653));
  INV_X1    g452(.A(new_n653), .ZN(new_n654));
  OAI211_X1 g453(.A(new_n650), .B(new_n654), .C1(new_n645), .C2(new_n639), .ZN(new_n655));
  XNOR2_X1  g454(.A(new_n645), .B(KEYINPUT105), .ZN(new_n656));
  AND2_X1   g455(.A1(new_n644), .A2(new_n656), .ZN(new_n657));
  NOR2_X1   g456(.A1(new_n639), .A2(new_n645), .ZN(new_n658));
  OAI21_X1  g457(.A(new_n653), .B1(new_n657), .B2(new_n658), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n655), .A2(new_n659), .ZN(new_n660));
  INV_X1    g459(.A(new_n660), .ZN(new_n661));
  AND2_X1   g460(.A1(new_n635), .A2(new_n661), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n563), .A2(new_n662), .ZN(new_n663));
  INV_X1    g462(.A(new_n663), .ZN(new_n664));
  NOR2_X1   g463(.A1(new_n459), .A2(new_n460), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  XNOR2_X1  g465(.A(new_n666), .B(G1gat), .ZN(G1324gat));
  NOR2_X1   g466(.A1(new_n663), .A2(new_n427), .ZN(new_n668));
  NOR2_X1   g467(.A1(new_n519), .A2(new_n521), .ZN(new_n669));
  INV_X1    g468(.A(new_n669), .ZN(new_n670));
  NAND2_X1  g469(.A1(new_n519), .A2(new_n521), .ZN(new_n671));
  NAND3_X1  g470(.A1(new_n668), .A2(new_n670), .A3(new_n671), .ZN(new_n672));
  INV_X1    g471(.A(KEYINPUT42), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  NAND4_X1  g473(.A1(new_n668), .A2(KEYINPUT42), .A3(new_n670), .A4(new_n671), .ZN(new_n675));
  OAI211_X1 g474(.A(new_n674), .B(new_n675), .C1(new_n521), .C2(new_n668), .ZN(G1325gat));
  NAND2_X1  g475(.A1(new_n489), .A2(new_n491), .ZN(new_n677));
  AND3_X1   g476(.A1(new_n664), .A2(G15gat), .A3(new_n677), .ZN(new_n678));
  AOI21_X1  g477(.A(G15gat), .B1(new_n664), .B2(new_n477), .ZN(new_n679));
  NOR2_X1   g478(.A1(new_n678), .A2(new_n679), .ZN(G1326gat));
  NOR2_X1   g479(.A1(new_n663), .A2(new_n403), .ZN(new_n681));
  XNOR2_X1  g480(.A(KEYINPUT43), .B(G22gat), .ZN(new_n682));
  XNOR2_X1  g481(.A(KEYINPUT106), .B(KEYINPUT107), .ZN(new_n683));
  XNOR2_X1  g482(.A(new_n682), .B(new_n683), .ZN(new_n684));
  XNOR2_X1  g483(.A(new_n681), .B(new_n684), .ZN(G1327gat));
  INV_X1    g484(.A(new_n629), .ZN(new_n686));
  OAI211_X1 g485(.A(KEYINPUT44), .B(new_n686), .C1(new_n487), .C2(new_n516), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n598), .A2(new_n630), .ZN(new_n688));
  INV_X1    g487(.A(new_n688), .ZN(new_n689));
  NOR2_X1   g488(.A1(new_n689), .A2(new_n660), .ZN(new_n690));
  INV_X1    g489(.A(new_n690), .ZN(new_n691));
  AND3_X1   g490(.A1(new_n559), .A2(KEYINPUT108), .A3(new_n560), .ZN(new_n692));
  AOI21_X1  g491(.A(KEYINPUT108), .B1(new_n559), .B2(new_n560), .ZN(new_n693));
  NOR2_X1   g492(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  INV_X1    g493(.A(new_n694), .ZN(new_n695));
  NOR2_X1   g494(.A1(new_n691), .A2(new_n695), .ZN(new_n696));
  NAND2_X1  g495(.A1(new_n480), .A2(new_n486), .ZN(new_n697));
  AND3_X1   g496(.A1(new_n314), .A2(new_n406), .A3(new_n403), .ZN(new_n698));
  AOI21_X1  g497(.A(new_n406), .B1(new_n314), .B2(new_n403), .ZN(new_n699));
  NOR3_X1   g498(.A1(new_n698), .A2(new_n699), .A3(new_n461), .ZN(new_n700));
  INV_X1    g499(.A(KEYINPUT35), .ZN(new_n701));
  OAI21_X1  g500(.A(new_n697), .B1(new_n700), .B2(new_n701), .ZN(new_n702));
  AND2_X1   g501(.A1(new_n489), .A2(new_n491), .ZN(new_n703));
  NAND3_X1  g502(.A1(new_n403), .A2(new_n504), .A3(new_n514), .ZN(new_n704));
  NAND4_X1  g503(.A1(new_n703), .A2(KEYINPUT109), .A3(new_n488), .A4(new_n704), .ZN(new_n705));
  INV_X1    g504(.A(KEYINPUT109), .ZN(new_n706));
  OAI21_X1  g505(.A(new_n706), .B1(new_n492), .B2(new_n515), .ZN(new_n707));
  AND2_X1   g506(.A1(new_n705), .A2(new_n707), .ZN(new_n708));
  AOI21_X1  g507(.A(new_n629), .B1(new_n702), .B2(new_n708), .ZN(new_n709));
  OAI211_X1 g508(.A(new_n687), .B(new_n696), .C1(new_n709), .C2(KEYINPUT44), .ZN(new_n710));
  INV_X1    g509(.A(new_n665), .ZN(new_n711));
  OAI21_X1  g510(.A(G29gat), .B1(new_n710), .B2(new_n711), .ZN(new_n712));
  OAI211_X1 g511(.A(new_n686), .B(new_n561), .C1(new_n487), .C2(new_n516), .ZN(new_n713));
  NOR2_X1   g512(.A1(new_n713), .A2(new_n691), .ZN(new_n714));
  NAND3_X1  g513(.A1(new_n714), .A2(new_n528), .A3(new_n665), .ZN(new_n715));
  AND2_X1   g514(.A1(new_n715), .A2(KEYINPUT45), .ZN(new_n716));
  NOR2_X1   g515(.A1(new_n715), .A2(KEYINPUT45), .ZN(new_n717));
  OAI21_X1  g516(.A(new_n712), .B1(new_n716), .B2(new_n717), .ZN(G1328gat));
  NAND3_X1  g517(.A1(new_n714), .A2(new_n529), .A3(new_n512), .ZN(new_n719));
  XOR2_X1   g518(.A(KEYINPUT110), .B(KEYINPUT46), .Z(new_n720));
  INV_X1    g519(.A(new_n720), .ZN(new_n721));
  OR2_X1    g520(.A1(new_n719), .A2(new_n721), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n719), .A2(new_n721), .ZN(new_n723));
  NOR2_X1   g522(.A1(new_n710), .A2(new_n427), .ZN(new_n724));
  OAI211_X1 g523(.A(new_n722), .B(new_n723), .C1(new_n529), .C2(new_n724), .ZN(G1329gat));
  OAI21_X1  g524(.A(G43gat), .B1(new_n710), .B2(new_n703), .ZN(new_n726));
  NOR2_X1   g525(.A1(new_n476), .A2(G43gat), .ZN(new_n727));
  INV_X1    g526(.A(new_n727), .ZN(new_n728));
  NOR3_X1   g527(.A1(new_n713), .A2(new_n691), .A3(new_n728), .ZN(new_n729));
  INV_X1    g528(.A(new_n729), .ZN(new_n730));
  NAND2_X1  g529(.A1(new_n726), .A2(new_n730), .ZN(new_n731));
  AOI21_X1  g530(.A(KEYINPUT47), .B1(new_n731), .B2(KEYINPUT111), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n705), .A2(new_n707), .ZN(new_n733));
  OAI21_X1  g532(.A(new_n686), .B1(new_n487), .B2(new_n733), .ZN(new_n734));
  INV_X1    g533(.A(KEYINPUT44), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  NAND4_X1  g535(.A1(new_n736), .A2(new_n677), .A3(new_n696), .A4(new_n687), .ZN(new_n737));
  AOI21_X1  g536(.A(new_n729), .B1(new_n737), .B2(G43gat), .ZN(new_n738));
  INV_X1    g537(.A(KEYINPUT111), .ZN(new_n739));
  INV_X1    g538(.A(KEYINPUT47), .ZN(new_n740));
  NOR3_X1   g539(.A1(new_n738), .A2(new_n739), .A3(new_n740), .ZN(new_n741));
  NOR2_X1   g540(.A1(new_n732), .A2(new_n741), .ZN(G1330gat));
  INV_X1    g541(.A(new_n710), .ZN(new_n743));
  NAND3_X1  g542(.A1(new_n743), .A2(G50gat), .A3(new_n484), .ZN(new_n744));
  NOR3_X1   g543(.A1(new_n713), .A2(new_n403), .A3(new_n691), .ZN(new_n745));
  OR2_X1    g544(.A1(new_n745), .A2(G50gat), .ZN(new_n746));
  AND3_X1   g545(.A1(new_n744), .A2(new_n746), .A3(KEYINPUT48), .ZN(new_n747));
  AOI21_X1  g546(.A(KEYINPUT48), .B1(new_n744), .B2(new_n746), .ZN(new_n748));
  NOR2_X1   g547(.A1(new_n747), .A2(new_n748), .ZN(G1331gat));
  NAND2_X1  g548(.A1(new_n702), .A2(new_n708), .ZN(new_n750));
  NOR2_X1   g549(.A1(new_n661), .A2(new_n694), .ZN(new_n751));
  NAND3_X1  g550(.A1(new_n750), .A2(new_n635), .A3(new_n751), .ZN(new_n752));
  NOR2_X1   g551(.A1(new_n752), .A2(new_n711), .ZN(new_n753));
  XOR2_X1   g552(.A(new_n753), .B(G57gat), .Z(G1332gat));
  NAND4_X1  g553(.A1(new_n750), .A2(new_n635), .A3(new_n512), .A4(new_n751), .ZN(new_n755));
  AND2_X1   g554(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n756));
  OR3_X1    g555(.A1(new_n755), .A2(KEYINPUT112), .A3(new_n756), .ZN(new_n757));
  OAI21_X1  g556(.A(KEYINPUT112), .B1(new_n755), .B2(new_n756), .ZN(new_n758));
  NAND2_X1  g557(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  NOR2_X1   g558(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n760));
  XNOR2_X1  g559(.A(new_n759), .B(new_n760), .ZN(G1333gat));
  OAI21_X1  g560(.A(G71gat), .B1(new_n752), .B2(new_n703), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n477), .A2(new_n568), .ZN(new_n763));
  OAI21_X1  g562(.A(new_n762), .B1(new_n752), .B2(new_n763), .ZN(new_n764));
  XOR2_X1   g563(.A(new_n764), .B(KEYINPUT50), .Z(G1334gat));
  NOR2_X1   g564(.A1(new_n752), .A2(new_n403), .ZN(new_n766));
  XOR2_X1   g565(.A(KEYINPUT113), .B(G78gat), .Z(new_n767));
  XNOR2_X1  g566(.A(new_n766), .B(new_n767), .ZN(G1335gat));
  NAND4_X1  g567(.A1(new_n736), .A2(new_n688), .A3(new_n687), .A4(new_n751), .ZN(new_n769));
  OAI21_X1  g568(.A(G85gat), .B1(new_n769), .B2(new_n711), .ZN(new_n770));
  NOR2_X1   g569(.A1(new_n689), .A2(new_n694), .ZN(new_n771));
  OAI211_X1 g570(.A(new_n686), .B(new_n771), .C1(new_n487), .C2(new_n733), .ZN(new_n772));
  INV_X1    g571(.A(KEYINPUT51), .ZN(new_n773));
  NAND2_X1  g572(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  NAND4_X1  g573(.A1(new_n750), .A2(KEYINPUT51), .A3(new_n686), .A4(new_n771), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  NAND3_X1  g575(.A1(new_n665), .A2(new_n660), .A3(new_n605), .ZN(new_n777));
  XOR2_X1   g576(.A(new_n777), .B(KEYINPUT114), .Z(new_n778));
  NAND2_X1  g577(.A1(new_n776), .A2(new_n778), .ZN(new_n779));
  NAND2_X1  g578(.A1(new_n770), .A2(new_n779), .ZN(G1336gat));
  OAI21_X1  g579(.A(G92gat), .B1(new_n769), .B2(new_n427), .ZN(new_n781));
  NAND3_X1  g580(.A1(new_n774), .A2(new_n775), .A3(KEYINPUT115), .ZN(new_n782));
  INV_X1    g581(.A(KEYINPUT115), .ZN(new_n783));
  NAND3_X1  g582(.A1(new_n772), .A2(new_n783), .A3(new_n773), .ZN(new_n784));
  NOR3_X1   g583(.A1(new_n661), .A2(G92gat), .A3(new_n427), .ZN(new_n785));
  NAND3_X1  g584(.A1(new_n782), .A2(new_n784), .A3(new_n785), .ZN(new_n786));
  NAND2_X1  g585(.A1(new_n781), .A2(new_n786), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n787), .A2(KEYINPUT52), .ZN(new_n788));
  AOI21_X1  g587(.A(KEYINPUT52), .B1(new_n776), .B2(new_n785), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n781), .A2(new_n789), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n788), .A2(new_n790), .ZN(G1337gat));
  OAI21_X1  g590(.A(G99gat), .B1(new_n769), .B2(new_n703), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n776), .A2(new_n660), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n477), .A2(new_n296), .ZN(new_n794));
  OAI21_X1  g593(.A(new_n792), .B1(new_n793), .B2(new_n794), .ZN(G1338gat));
  OAI21_X1  g594(.A(G106gat), .B1(new_n769), .B2(new_n403), .ZN(new_n796));
  INV_X1    g595(.A(KEYINPUT53), .ZN(new_n797));
  NOR2_X1   g596(.A1(new_n403), .A2(G106gat), .ZN(new_n798));
  INV_X1    g597(.A(new_n798), .ZN(new_n799));
  OAI211_X1 g598(.A(new_n796), .B(new_n797), .C1(new_n793), .C2(new_n799), .ZN(new_n800));
  NOR2_X1   g599(.A1(new_n799), .A2(new_n661), .ZN(new_n801));
  NAND3_X1  g600(.A1(new_n782), .A2(new_n784), .A3(new_n801), .ZN(new_n802));
  AND2_X1   g601(.A1(new_n796), .A2(new_n802), .ZN(new_n803));
  OAI21_X1  g602(.A(new_n800), .B1(new_n803), .B2(new_n797), .ZN(G1339gat));
  AOI21_X1  g603(.A(new_n543), .B1(new_n541), .B2(new_n542), .ZN(new_n805));
  NOR2_X1   g604(.A1(new_n547), .A2(new_n548), .ZN(new_n806));
  OAI21_X1  g605(.A(new_n555), .B1(new_n805), .B2(new_n806), .ZN(new_n807));
  AND2_X1   g606(.A1(new_n560), .A2(new_n807), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n660), .A2(new_n808), .ZN(new_n809));
  XNOR2_X1  g608(.A(KEYINPUT117), .B(KEYINPUT54), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n657), .A2(new_n810), .ZN(new_n811));
  INV_X1    g610(.A(new_n656), .ZN(new_n812));
  OAI211_X1 g611(.A(new_n812), .B(new_n636), .C1(new_n641), .C2(new_n643), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n813), .A2(KEYINPUT116), .ZN(new_n814));
  AND3_X1   g613(.A1(new_n644), .A2(KEYINPUT104), .A3(new_n645), .ZN(new_n815));
  AOI21_X1  g614(.A(KEYINPUT104), .B1(new_n644), .B2(new_n645), .ZN(new_n816));
  OAI21_X1  g615(.A(new_n814), .B1(new_n815), .B2(new_n816), .ZN(new_n817));
  OAI21_X1  g616(.A(KEYINPUT54), .B1(new_n813), .B2(KEYINPUT116), .ZN(new_n818));
  OAI211_X1 g617(.A(new_n653), .B(new_n811), .C1(new_n817), .C2(new_n818), .ZN(new_n819));
  INV_X1    g618(.A(KEYINPUT55), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  INV_X1    g620(.A(new_n818), .ZN(new_n822));
  NAND3_X1  g621(.A1(new_n650), .A2(new_n822), .A3(new_n814), .ZN(new_n823));
  NAND4_X1  g622(.A1(new_n823), .A2(KEYINPUT55), .A3(new_n653), .A4(new_n811), .ZN(new_n824));
  NAND3_X1  g623(.A1(new_n821), .A2(new_n655), .A3(new_n824), .ZN(new_n825));
  OAI21_X1  g624(.A(new_n809), .B1(new_n825), .B2(new_n695), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n826), .A2(new_n629), .ZN(new_n827));
  NAND4_X1  g626(.A1(new_n821), .A2(new_n655), .A3(new_n824), .A4(new_n808), .ZN(new_n828));
  NOR2_X1   g627(.A1(new_n828), .A2(new_n629), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n829), .A2(KEYINPUT118), .ZN(new_n830));
  INV_X1    g629(.A(KEYINPUT118), .ZN(new_n831));
  OAI21_X1  g630(.A(new_n831), .B1(new_n828), .B2(new_n629), .ZN(new_n832));
  NAND3_X1  g631(.A1(new_n827), .A2(new_n830), .A3(new_n832), .ZN(new_n833));
  NAND2_X1  g632(.A1(new_n833), .A2(new_n688), .ZN(new_n834));
  AND4_X1   g633(.A1(new_n633), .A2(new_n634), .A3(new_n661), .A4(new_n695), .ZN(new_n835));
  INV_X1    g634(.A(new_n835), .ZN(new_n836));
  NAND2_X1  g635(.A1(new_n834), .A2(new_n836), .ZN(new_n837));
  NOR2_X1   g636(.A1(new_n711), .A2(new_n512), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n837), .A2(new_n838), .ZN(new_n839));
  NOR2_X1   g638(.A1(new_n698), .A2(new_n699), .ZN(new_n840));
  INV_X1    g639(.A(new_n840), .ZN(new_n841));
  NOR3_X1   g640(.A1(new_n839), .A2(KEYINPUT119), .A3(new_n841), .ZN(new_n842));
  INV_X1    g641(.A(KEYINPUT119), .ZN(new_n843));
  AOI21_X1  g642(.A(new_n835), .B1(new_n833), .B2(new_n688), .ZN(new_n844));
  INV_X1    g643(.A(new_n838), .ZN(new_n845));
  NOR2_X1   g644(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  AOI21_X1  g645(.A(new_n843), .B1(new_n846), .B2(new_n840), .ZN(new_n847));
  OR4_X1    g646(.A1(G113gat), .A2(new_n842), .A3(new_n695), .A4(new_n847), .ZN(new_n848));
  INV_X1    g647(.A(new_n485), .ZN(new_n849));
  NOR2_X1   g648(.A1(new_n839), .A2(new_n849), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n850), .A2(new_n561), .ZN(new_n851));
  NAND2_X1  g650(.A1(new_n851), .A2(G113gat), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n848), .A2(new_n852), .ZN(G1340gat));
  NAND2_X1  g652(.A1(new_n660), .A2(new_n213), .ZN(new_n854));
  NOR3_X1   g653(.A1(new_n842), .A2(new_n847), .A3(new_n854), .ZN(new_n855));
  INV_X1    g654(.A(new_n855), .ZN(new_n856));
  INV_X1    g655(.A(KEYINPUT120), .ZN(new_n857));
  AOI21_X1  g656(.A(new_n213), .B1(new_n850), .B2(new_n660), .ZN(new_n858));
  INV_X1    g657(.A(new_n858), .ZN(new_n859));
  NAND3_X1  g658(.A1(new_n856), .A2(new_n857), .A3(new_n859), .ZN(new_n860));
  OAI21_X1  g659(.A(KEYINPUT120), .B1(new_n855), .B2(new_n858), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n860), .A2(new_n861), .ZN(G1341gat));
  NOR2_X1   g661(.A1(new_n839), .A2(new_n841), .ZN(new_n863));
  AOI21_X1  g662(.A(G127gat), .B1(new_n863), .B2(new_n689), .ZN(new_n864));
  NOR2_X1   g663(.A1(new_n688), .A2(new_n209), .ZN(new_n865));
  AOI21_X1  g664(.A(new_n864), .B1(new_n850), .B2(new_n865), .ZN(G1342gat));
  NOR4_X1   g665(.A1(new_n839), .A2(G134gat), .A3(new_n629), .A4(new_n841), .ZN(new_n867));
  XNOR2_X1  g666(.A(new_n867), .B(KEYINPUT56), .ZN(new_n868));
  NOR3_X1   g667(.A1(new_n839), .A2(new_n629), .A3(new_n849), .ZN(new_n869));
  OAI21_X1  g668(.A(new_n868), .B1(new_n202), .B2(new_n869), .ZN(G1343gat));
  INV_X1    g669(.A(G141gat), .ZN(new_n871));
  INV_X1    g670(.A(KEYINPUT57), .ZN(new_n872));
  NAND3_X1  g671(.A1(new_n837), .A2(new_n872), .A3(new_n484), .ZN(new_n873));
  NOR2_X1   g672(.A1(new_n845), .A2(new_n677), .ZN(new_n874));
  NAND4_X1  g673(.A1(new_n821), .A2(new_n655), .A3(new_n824), .A4(new_n561), .ZN(new_n875));
  AOI21_X1  g674(.A(new_n686), .B1(new_n875), .B2(new_n809), .ZN(new_n876));
  INV_X1    g675(.A(new_n876), .ZN(new_n877));
  NAND3_X1  g676(.A1(new_n877), .A2(new_n830), .A3(new_n832), .ZN(new_n878));
  AOI21_X1  g677(.A(new_n835), .B1(new_n878), .B2(new_n688), .ZN(new_n879));
  OAI21_X1  g678(.A(KEYINPUT57), .B1(new_n879), .B2(new_n403), .ZN(new_n880));
  AND3_X1   g679(.A1(new_n873), .A2(new_n874), .A3(new_n880), .ZN(new_n881));
  AOI21_X1  g680(.A(new_n871), .B1(new_n881), .B2(new_n694), .ZN(new_n882));
  NOR2_X1   g681(.A1(new_n677), .A2(new_n403), .ZN(new_n883));
  XNOR2_X1  g682(.A(new_n883), .B(KEYINPUT121), .ZN(new_n884));
  AND3_X1   g683(.A1(new_n837), .A2(new_n838), .A3(new_n884), .ZN(new_n885));
  INV_X1    g684(.A(KEYINPUT122), .ZN(new_n886));
  NAND4_X1  g685(.A1(new_n885), .A2(new_n886), .A3(new_n871), .A4(new_n561), .ZN(new_n887));
  NAND4_X1  g686(.A1(new_n846), .A2(new_n871), .A3(new_n561), .A4(new_n884), .ZN(new_n888));
  NAND2_X1  g687(.A1(new_n888), .A2(KEYINPUT122), .ZN(new_n889));
  NAND2_X1  g688(.A1(new_n887), .A2(new_n889), .ZN(new_n890));
  OAI21_X1  g689(.A(KEYINPUT58), .B1(new_n882), .B2(new_n890), .ZN(new_n891));
  AOI21_X1  g690(.A(new_n871), .B1(new_n881), .B2(new_n561), .ZN(new_n892));
  INV_X1    g691(.A(KEYINPUT58), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n888), .A2(new_n893), .ZN(new_n894));
  OAI21_X1  g693(.A(new_n891), .B1(new_n892), .B2(new_n894), .ZN(G1344gat));
  INV_X1    g694(.A(G148gat), .ZN(new_n896));
  NAND3_X1  g695(.A1(new_n885), .A2(new_n896), .A3(new_n660), .ZN(new_n897));
  NAND4_X1  g696(.A1(new_n873), .A2(new_n880), .A3(new_n660), .A4(new_n874), .ZN(new_n898));
  INV_X1    g697(.A(KEYINPUT123), .ZN(new_n899));
  INV_X1    g698(.A(KEYINPUT59), .ZN(new_n900));
  AND2_X1   g699(.A1(new_n900), .A2(G148gat), .ZN(new_n901));
  AND3_X1   g700(.A1(new_n898), .A2(new_n899), .A3(new_n901), .ZN(new_n902));
  AOI21_X1  g701(.A(new_n899), .B1(new_n898), .B2(new_n901), .ZN(new_n903));
  NOR2_X1   g702(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  INV_X1    g703(.A(KEYINPUT124), .ZN(new_n905));
  OAI21_X1  g704(.A(new_n688), .B1(new_n876), .B2(new_n829), .ZN(new_n906));
  NAND4_X1  g705(.A1(new_n633), .A2(new_n634), .A3(new_n661), .A4(new_n562), .ZN(new_n907));
  AND2_X1   g706(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  OAI211_X1 g707(.A(new_n905), .B(new_n872), .C1(new_n908), .C2(new_n403), .ZN(new_n909));
  AOI21_X1  g708(.A(new_n403), .B1(new_n906), .B2(new_n907), .ZN(new_n910));
  OAI21_X1  g709(.A(KEYINPUT124), .B1(new_n910), .B2(KEYINPUT57), .ZN(new_n911));
  NAND2_X1  g710(.A1(new_n909), .A2(new_n911), .ZN(new_n912));
  NOR3_X1   g711(.A1(new_n844), .A2(new_n872), .A3(new_n403), .ZN(new_n913));
  OAI211_X1 g712(.A(new_n660), .B(new_n874), .C1(new_n912), .C2(new_n913), .ZN(new_n914));
  AOI21_X1  g713(.A(new_n900), .B1(new_n914), .B2(G148gat), .ZN(new_n915));
  OAI21_X1  g714(.A(new_n897), .B1(new_n904), .B2(new_n915), .ZN(G1345gat));
  NAND2_X1  g715(.A1(new_n333), .A2(new_n334), .ZN(new_n917));
  NOR2_X1   g716(.A1(new_n688), .A2(new_n917), .ZN(new_n918));
  NAND2_X1  g717(.A1(new_n885), .A2(new_n689), .ZN(new_n919));
  AOI22_X1  g718(.A1(new_n881), .A2(new_n918), .B1(new_n919), .B2(new_n917), .ZN(G1346gat));
  AOI21_X1  g719(.A(G162gat), .B1(new_n885), .B2(new_n686), .ZN(new_n921));
  NOR2_X1   g720(.A1(new_n629), .A2(new_n319), .ZN(new_n922));
  AOI21_X1  g721(.A(new_n921), .B1(new_n881), .B2(new_n922), .ZN(G1347gat));
  NOR4_X1   g722(.A1(new_n844), .A2(new_n665), .A3(new_n849), .A4(new_n427), .ZN(new_n924));
  INV_X1    g723(.A(new_n924), .ZN(new_n925));
  OAI21_X1  g724(.A(G169gat), .B1(new_n925), .B2(new_n562), .ZN(new_n926));
  NOR3_X1   g725(.A1(new_n844), .A2(new_n665), .A3(new_n841), .ZN(new_n927));
  NAND2_X1  g726(.A1(new_n927), .A2(new_n512), .ZN(new_n928));
  OR2_X1    g727(.A1(new_n695), .A2(G169gat), .ZN(new_n929));
  OAI21_X1  g728(.A(new_n926), .B1(new_n928), .B2(new_n929), .ZN(G1348gat));
  INV_X1    g729(.A(new_n928), .ZN(new_n931));
  AOI21_X1  g730(.A(G176gat), .B1(new_n931), .B2(new_n660), .ZN(new_n932));
  AND2_X1   g731(.A1(new_n660), .A2(G176gat), .ZN(new_n933));
  AOI21_X1  g732(.A(new_n932), .B1(new_n924), .B2(new_n933), .ZN(G1349gat));
  NAND3_X1  g733(.A1(new_n931), .A2(new_n689), .A3(new_n244), .ZN(new_n935));
  OAI21_X1  g734(.A(G183gat), .B1(new_n925), .B2(new_n688), .ZN(new_n936));
  NAND2_X1  g735(.A1(new_n935), .A2(new_n936), .ZN(new_n937));
  NAND2_X1  g736(.A1(new_n937), .A2(KEYINPUT60), .ZN(new_n938));
  INV_X1    g737(.A(KEYINPUT60), .ZN(new_n939));
  NAND3_X1  g738(.A1(new_n935), .A2(new_n939), .A3(new_n936), .ZN(new_n940));
  NAND2_X1  g739(.A1(new_n938), .A2(new_n940), .ZN(G1350gat));
  NAND3_X1  g740(.A1(new_n931), .A2(new_n251), .A3(new_n686), .ZN(new_n942));
  OAI21_X1  g741(.A(G190gat), .B1(new_n925), .B2(new_n629), .ZN(new_n943));
  AND2_X1   g742(.A1(new_n943), .A2(KEYINPUT61), .ZN(new_n944));
  NOR2_X1   g743(.A1(new_n943), .A2(KEYINPUT61), .ZN(new_n945));
  OAI21_X1  g744(.A(new_n942), .B1(new_n944), .B2(new_n945), .ZN(G1351gat));
  NOR3_X1   g745(.A1(new_n677), .A2(new_n665), .A3(new_n427), .ZN(new_n947));
  XOR2_X1   g746(.A(new_n947), .B(KEYINPUT125), .Z(new_n948));
  OAI211_X1 g747(.A(new_n561), .B(new_n948), .C1(new_n912), .C2(new_n913), .ZN(new_n949));
  NAND2_X1  g748(.A1(new_n949), .A2(G197gat), .ZN(new_n950));
  AND3_X1   g749(.A1(new_n837), .A2(new_n484), .A3(new_n947), .ZN(new_n951));
  INV_X1    g750(.A(G197gat), .ZN(new_n952));
  NAND3_X1  g751(.A1(new_n951), .A2(new_n952), .A3(new_n694), .ZN(new_n953));
  NAND2_X1  g752(.A1(new_n950), .A2(new_n953), .ZN(new_n954));
  NAND2_X1  g753(.A1(new_n954), .A2(KEYINPUT126), .ZN(new_n955));
  INV_X1    g754(.A(KEYINPUT126), .ZN(new_n956));
  NAND3_X1  g755(.A1(new_n950), .A2(new_n956), .A3(new_n953), .ZN(new_n957));
  NAND2_X1  g756(.A1(new_n955), .A2(new_n957), .ZN(G1352gat));
  OAI211_X1 g757(.A(new_n660), .B(new_n948), .C1(new_n912), .C2(new_n913), .ZN(new_n959));
  INV_X1    g758(.A(KEYINPUT127), .ZN(new_n960));
  OR2_X1    g759(.A1(new_n959), .A2(new_n960), .ZN(new_n961));
  NAND2_X1  g760(.A1(new_n959), .A2(new_n960), .ZN(new_n962));
  NAND3_X1  g761(.A1(new_n961), .A2(G204gat), .A3(new_n962), .ZN(new_n963));
  INV_X1    g762(.A(G204gat), .ZN(new_n964));
  NAND3_X1  g763(.A1(new_n951), .A2(new_n964), .A3(new_n660), .ZN(new_n965));
  XOR2_X1   g764(.A(new_n965), .B(KEYINPUT62), .Z(new_n966));
  NAND2_X1  g765(.A1(new_n963), .A2(new_n966), .ZN(G1353gat));
  INV_X1    g766(.A(G211gat), .ZN(new_n968));
  NAND3_X1  g767(.A1(new_n951), .A2(new_n968), .A3(new_n689), .ZN(new_n969));
  OAI211_X1 g768(.A(new_n689), .B(new_n947), .C1(new_n912), .C2(new_n913), .ZN(new_n970));
  AND3_X1   g769(.A1(new_n970), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n971));
  AOI21_X1  g770(.A(KEYINPUT63), .B1(new_n970), .B2(G211gat), .ZN(new_n972));
  OAI21_X1  g771(.A(new_n969), .B1(new_n971), .B2(new_n972), .ZN(G1354gat));
  OAI211_X1 g772(.A(new_n686), .B(new_n948), .C1(new_n912), .C2(new_n913), .ZN(new_n974));
  NAND2_X1  g773(.A1(new_n974), .A2(G218gat), .ZN(new_n975));
  INV_X1    g774(.A(G218gat), .ZN(new_n976));
  NAND3_X1  g775(.A1(new_n951), .A2(new_n976), .A3(new_n686), .ZN(new_n977));
  NAND2_X1  g776(.A1(new_n975), .A2(new_n977), .ZN(G1355gat));
endmodule


