

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601,
         n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612,
         n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623,
         n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634,
         n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645,
         n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656,
         n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667,
         n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678,
         n679, n680, n681, n682, n683, n684, n685, n687, n688, n689, n690,
         n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701,
         n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712,
         n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723,
         n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734,
         n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745,
         n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756,
         n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n767,
         n768, n769, n770, n771, n772, n773, n774, n775, n776, n777, n778,
         n779, n780, n781, n782, n783, n784, n785, n786, n787, n788, n789,
         n790, n791, n792, n793, n794, n795, n796, n797, n798, n799, n800,
         n801, n802, n803, n804, n805, n806, n807, n808, n809, n810, n811,
         n812, n813, n814, n815, n816, n817, n818, n819, n820, n821, n822,
         n823, n824, n825, n826, n827, n828, n829, n830, n831, n832, n833,
         n834, n835, n836, n837, n838, n839, n840, n841, n842, n843, n844,
         n845, n846, n847, n848, n849, n850, n851, n852, n853, n854, n855,
         n856, n857, n858, n859, n860, n861, n862, n863, n864, n865, n866,
         n867, n868, n869, n870, n871, n872, n873, n874, n875, n876, n877,
         n878, n879, n880, n881, n882, n883, n884, n885, n886, n887, n888,
         n889, n890, n891, n892, n893, n894, n895, n896, n897, n898, n899,
         n900, n901, n902, n903, n904, n905, n906, n907, n908, n909, n910,
         n911, n912, n913, n914, n915, n916, n917, n918, n919, n920, n921,
         n922, n923, n924, n925, n926, n927, n928, n929, n930, n931, n932,
         n933, n934, n935, n936, n937, n938, n939, n940, n941, n942, n943,
         n944, n945, n946, n947, n948, n949, n950, n951, n952, n953, n954,
         n955, n956, n957, n958, n959, n960, n961, n962, n963, n964, n965,
         n966, n967, n968, n969, n970, n971, n972, n973, n974, n975, n976,
         n977, n978, n979, n980, n981, n982, n983, n984, n985, n986, n987,
         n988, n989, n990, n991, n992, n993, n994, n995, n996, n997, n998,
         n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008,
         n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018,
         n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028,
         n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038,
         n1039, n1040, n1041;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  XOR2_X1 U554 ( .A(KEYINPUT15), .B(n584), .Z(n1021) );
  XNOR2_X2 U555 ( .A(n774), .B(n773), .ZN(n805) );
  OR2_X2 U556 ( .A1(n772), .A2(n771), .ZN(n774) );
  XNOR2_X2 U557 ( .A(G2104), .B(KEYINPUT67), .ZN(n523) );
  OR2_X1 U558 ( .A1(n778), .A2(n770), .ZN(n768) );
  XNOR2_X1 U559 ( .A(n723), .B(KEYINPUT30), .ZN(n724) );
  INV_X1 U560 ( .A(KEYINPUT64), .ZN(n790) );
  INV_X1 U561 ( .A(KEYINPUT68), .ZN(n524) );
  NOR2_X1 U562 ( .A1(n761), .A2(n760), .ZN(n762) );
  BUF_X1 U563 ( .A(n736), .Z(n763) );
  INV_X1 U564 ( .A(n746), .ZN(n736) );
  INV_X1 U565 ( .A(KEYINPUT97), .ZN(n719) );
  XNOR2_X1 U566 ( .A(n720), .B(n719), .ZN(n811) );
  NOR2_X1 U567 ( .A1(n684), .A2(G1384), .ZN(n685) );
  XNOR2_X1 U568 ( .A(n685), .B(KEYINPUT65), .ZN(n717) );
  NOR2_X1 U569 ( .A1(G2105), .A2(n523), .ZN(n521) );
  NOR2_X1 U570 ( .A1(G651), .A2(n653), .ZN(n647) );
  AND2_X1 U571 ( .A1(n533), .A2(n532), .ZN(G160) );
  XOR2_X2 U572 ( .A(KEYINPUT69), .B(n521), .Z(n888) );
  NAND2_X1 U573 ( .A1(n888), .A2(G101), .ZN(n522) );
  XOR2_X1 U574 ( .A(KEYINPUT23), .B(n522), .Z(n533) );
  NAND2_X1 U575 ( .A1(n523), .A2(G2105), .ZN(n525) );
  XNOR2_X2 U576 ( .A(n525), .B(n524), .ZN(n885) );
  AND2_X1 U577 ( .A1(G125), .A2(n885), .ZN(n531) );
  AND2_X1 U578 ( .A1(G2105), .A2(G2104), .ZN(n884) );
  NAND2_X1 U579 ( .A1(G113), .A2(n884), .ZN(n528) );
  NOR2_X1 U580 ( .A1(G2105), .A2(G2104), .ZN(n526) );
  XOR2_X1 U581 ( .A(KEYINPUT17), .B(n526), .Z(n604) );
  NAND2_X1 U582 ( .A1(G137), .A2(n604), .ZN(n527) );
  NAND2_X1 U583 ( .A1(n528), .A2(n527), .ZN(n529) );
  XNOR2_X1 U584 ( .A(KEYINPUT70), .B(n529), .ZN(n530) );
  NOR2_X1 U585 ( .A1(n531), .A2(n530), .ZN(n532) );
  NOR2_X1 U586 ( .A1(G651), .A2(G543), .ZN(n638) );
  NAND2_X1 U587 ( .A1(G89), .A2(n638), .ZN(n534) );
  XNOR2_X1 U588 ( .A(n534), .B(KEYINPUT4), .ZN(n535) );
  XNOR2_X1 U589 ( .A(n535), .B(KEYINPUT78), .ZN(n538) );
  INV_X1 U590 ( .A(G651), .ZN(n540) );
  XOR2_X1 U591 ( .A(KEYINPUT0), .B(G543), .Z(n653) );
  OR2_X1 U592 ( .A1(n540), .A2(n653), .ZN(n536) );
  XNOR2_X1 U593 ( .A(KEYINPUT71), .B(n536), .ZN(n636) );
  NAND2_X1 U594 ( .A1(G76), .A2(n636), .ZN(n537) );
  NAND2_X1 U595 ( .A1(n538), .A2(n537), .ZN(n539) );
  XNOR2_X1 U596 ( .A(n539), .B(KEYINPUT5), .ZN(n548) );
  NAND2_X1 U597 ( .A1(n647), .A2(G51), .ZN(n545) );
  NOR2_X1 U598 ( .A1(G543), .A2(n540), .ZN(n542) );
  XNOR2_X1 U599 ( .A(KEYINPUT73), .B(KEYINPUT1), .ZN(n541) );
  XNOR2_X1 U600 ( .A(n542), .B(n541), .ZN(n543) );
  XNOR2_X2 U601 ( .A(KEYINPUT72), .B(n543), .ZN(n652) );
  NAND2_X1 U602 ( .A1(G63), .A2(n652), .ZN(n544) );
  NAND2_X1 U603 ( .A1(n545), .A2(n544), .ZN(n546) );
  XOR2_X1 U604 ( .A(KEYINPUT6), .B(n546), .Z(n547) );
  NAND2_X1 U605 ( .A1(n548), .A2(n547), .ZN(n549) );
  XNOR2_X1 U606 ( .A(n549), .B(KEYINPUT7), .ZN(G168) );
  NAND2_X1 U607 ( .A1(G90), .A2(n638), .ZN(n551) );
  NAND2_X1 U608 ( .A1(G77), .A2(n636), .ZN(n550) );
  NAND2_X1 U609 ( .A1(n551), .A2(n550), .ZN(n552) );
  XNOR2_X1 U610 ( .A(n552), .B(KEYINPUT9), .ZN(n554) );
  NAND2_X1 U611 ( .A1(G52), .A2(n647), .ZN(n553) );
  NAND2_X1 U612 ( .A1(n554), .A2(n553), .ZN(n557) );
  NAND2_X1 U613 ( .A1(n652), .A2(G64), .ZN(n555) );
  XOR2_X1 U614 ( .A(KEYINPUT74), .B(n555), .Z(n556) );
  NOR2_X1 U615 ( .A1(n557), .A2(n556), .ZN(G171) );
  INV_X1 U616 ( .A(G171), .ZN(G301) );
  AND2_X1 U617 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U618 ( .A(G132), .ZN(G219) );
  INV_X1 U619 ( .A(G82), .ZN(G220) );
  INV_X1 U620 ( .A(G57), .ZN(G237) );
  INV_X1 U621 ( .A(G69), .ZN(G235) );
  INV_X1 U622 ( .A(G108), .ZN(G238) );
  INV_X1 U623 ( .A(G120), .ZN(G236) );
  NAND2_X1 U624 ( .A1(n885), .A2(G126), .ZN(n559) );
  NAND2_X1 U625 ( .A1(n884), .A2(G114), .ZN(n558) );
  NAND2_X1 U626 ( .A1(n559), .A2(n558), .ZN(n560) );
  XNOR2_X1 U627 ( .A(n560), .B(KEYINPUT92), .ZN(n564) );
  NAND2_X1 U628 ( .A1(n604), .A2(G138), .ZN(n562) );
  NAND2_X1 U629 ( .A1(n888), .A2(G102), .ZN(n561) );
  NAND2_X1 U630 ( .A1(n562), .A2(n561), .ZN(n563) );
  NOR2_X1 U631 ( .A1(n564), .A2(n563), .ZN(n684) );
  BUF_X1 U632 ( .A(n684), .Z(G164) );
  XOR2_X1 U633 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  XOR2_X1 U634 ( .A(KEYINPUT11), .B(KEYINPUT76), .Z(n567) );
  NAND2_X1 U635 ( .A1(G7), .A2(G661), .ZN(n565) );
  XOR2_X1 U636 ( .A(n565), .B(KEYINPUT10), .Z(n930) );
  NAND2_X1 U637 ( .A1(G567), .A2(n930), .ZN(n566) );
  XNOR2_X1 U638 ( .A(n567), .B(n566), .ZN(G234) );
  NAND2_X1 U639 ( .A1(n652), .A2(G56), .ZN(n568) );
  XOR2_X1 U640 ( .A(KEYINPUT14), .B(n568), .Z(n574) );
  NAND2_X1 U641 ( .A1(n638), .A2(G81), .ZN(n569) );
  XNOR2_X1 U642 ( .A(n569), .B(KEYINPUT12), .ZN(n571) );
  NAND2_X1 U643 ( .A1(G68), .A2(n636), .ZN(n570) );
  NAND2_X1 U644 ( .A1(n571), .A2(n570), .ZN(n572) );
  XOR2_X1 U645 ( .A(KEYINPUT13), .B(n572), .Z(n573) );
  NOR2_X1 U646 ( .A1(n574), .A2(n573), .ZN(n576) );
  NAND2_X1 U647 ( .A1(n647), .A2(G43), .ZN(n575) );
  NAND2_X1 U648 ( .A1(n576), .A2(n575), .ZN(n1012) );
  INV_X1 U649 ( .A(G860), .ZN(n618) );
  OR2_X1 U650 ( .A1(n1012), .A2(n618), .ZN(G153) );
  NAND2_X1 U651 ( .A1(G868), .A2(G301), .ZN(n586) );
  NAND2_X1 U652 ( .A1(G79), .A2(n636), .ZN(n578) );
  NAND2_X1 U653 ( .A1(G54), .A2(n647), .ZN(n577) );
  NAND2_X1 U654 ( .A1(n578), .A2(n577), .ZN(n583) );
  NAND2_X1 U655 ( .A1(n638), .A2(G92), .ZN(n580) );
  NAND2_X1 U656 ( .A1(G66), .A2(n652), .ZN(n579) );
  NAND2_X1 U657 ( .A1(n580), .A2(n579), .ZN(n581) );
  XOR2_X1 U658 ( .A(KEYINPUT77), .B(n581), .Z(n582) );
  NOR2_X1 U659 ( .A1(n583), .A2(n582), .ZN(n584) );
  INV_X1 U660 ( .A(n1021), .ZN(n905) );
  INV_X1 U661 ( .A(G868), .ZN(n667) );
  NAND2_X1 U662 ( .A1(n905), .A2(n667), .ZN(n585) );
  NAND2_X1 U663 ( .A1(n586), .A2(n585), .ZN(G284) );
  NAND2_X1 U664 ( .A1(n638), .A2(G91), .ZN(n588) );
  NAND2_X1 U665 ( .A1(G65), .A2(n652), .ZN(n587) );
  NAND2_X1 U666 ( .A1(n588), .A2(n587), .ZN(n591) );
  NAND2_X1 U667 ( .A1(G53), .A2(n647), .ZN(n589) );
  XNOR2_X1 U668 ( .A(KEYINPUT75), .B(n589), .ZN(n590) );
  NOR2_X1 U669 ( .A1(n591), .A2(n590), .ZN(n593) );
  NAND2_X1 U670 ( .A1(n636), .A2(G78), .ZN(n592) );
  NAND2_X1 U671 ( .A1(n593), .A2(n592), .ZN(G299) );
  NOR2_X1 U672 ( .A1(G868), .A2(G299), .ZN(n595) );
  NOR2_X1 U673 ( .A1(G286), .A2(n667), .ZN(n594) );
  NOR2_X1 U674 ( .A1(n595), .A2(n594), .ZN(G297) );
  NAND2_X1 U675 ( .A1(n618), .A2(G559), .ZN(n596) );
  NAND2_X1 U676 ( .A1(n596), .A2(n1021), .ZN(n597) );
  XNOR2_X1 U677 ( .A(n597), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U678 ( .A1(G868), .A2(n1012), .ZN(n600) );
  NAND2_X1 U679 ( .A1(n1021), .A2(G868), .ZN(n598) );
  NOR2_X1 U680 ( .A1(G559), .A2(n598), .ZN(n599) );
  NOR2_X1 U681 ( .A1(n600), .A2(n599), .ZN(G282) );
  NAND2_X1 U682 ( .A1(G111), .A2(n884), .ZN(n602) );
  NAND2_X1 U683 ( .A1(G99), .A2(n888), .ZN(n601) );
  NAND2_X1 U684 ( .A1(n602), .A2(n601), .ZN(n603) );
  XNOR2_X1 U685 ( .A(n603), .B(KEYINPUT79), .ZN(n606) );
  BUF_X1 U686 ( .A(n604), .Z(n889) );
  NAND2_X1 U687 ( .A1(G135), .A2(n889), .ZN(n605) );
  NAND2_X1 U688 ( .A1(n606), .A2(n605), .ZN(n609) );
  NAND2_X1 U689 ( .A1(n885), .A2(G123), .ZN(n607) );
  XOR2_X1 U690 ( .A(KEYINPUT18), .B(n607), .Z(n608) );
  NOR2_X1 U691 ( .A1(n609), .A2(n608), .ZN(n985) );
  XNOR2_X1 U692 ( .A(G2096), .B(n985), .ZN(n610) );
  INV_X1 U693 ( .A(G2100), .ZN(n856) );
  NAND2_X1 U694 ( .A1(n610), .A2(n856), .ZN(G156) );
  NAND2_X1 U695 ( .A1(n638), .A2(G93), .ZN(n612) );
  NAND2_X1 U696 ( .A1(G67), .A2(n652), .ZN(n611) );
  NAND2_X1 U697 ( .A1(n612), .A2(n611), .ZN(n616) );
  NAND2_X1 U698 ( .A1(G80), .A2(n636), .ZN(n614) );
  NAND2_X1 U699 ( .A1(G55), .A2(n647), .ZN(n613) );
  NAND2_X1 U700 ( .A1(n614), .A2(n613), .ZN(n615) );
  OR2_X1 U701 ( .A1(n616), .A2(n615), .ZN(n666) );
  XNOR2_X1 U702 ( .A(n666), .B(KEYINPUT80), .ZN(n620) );
  NAND2_X1 U703 ( .A1(G559), .A2(n1021), .ZN(n617) );
  XOR2_X1 U704 ( .A(n1012), .B(n617), .Z(n664) );
  NAND2_X1 U705 ( .A1(n664), .A2(n618), .ZN(n619) );
  XNOR2_X1 U706 ( .A(n620), .B(n619), .ZN(G145) );
  AND2_X1 U707 ( .A1(n638), .A2(G85), .ZN(n624) );
  NAND2_X1 U708 ( .A1(n647), .A2(G47), .ZN(n622) );
  NAND2_X1 U709 ( .A1(G60), .A2(n652), .ZN(n621) );
  NAND2_X1 U710 ( .A1(n622), .A2(n621), .ZN(n623) );
  NOR2_X1 U711 ( .A1(n624), .A2(n623), .ZN(n626) );
  NAND2_X1 U712 ( .A1(n636), .A2(G72), .ZN(n625) );
  NAND2_X1 U713 ( .A1(n626), .A2(n625), .ZN(G290) );
  NAND2_X1 U714 ( .A1(G50), .A2(n647), .ZN(n633) );
  NAND2_X1 U715 ( .A1(G88), .A2(n638), .ZN(n628) );
  NAND2_X1 U716 ( .A1(G75), .A2(n636), .ZN(n627) );
  NAND2_X1 U717 ( .A1(n628), .A2(n627), .ZN(n631) );
  NAND2_X1 U718 ( .A1(G62), .A2(n652), .ZN(n629) );
  XNOR2_X1 U719 ( .A(KEYINPUT85), .B(n629), .ZN(n630) );
  NOR2_X1 U720 ( .A1(n631), .A2(n630), .ZN(n632) );
  NAND2_X1 U721 ( .A1(n633), .A2(n632), .ZN(n634) );
  XOR2_X1 U722 ( .A(n634), .B(KEYINPUT86), .Z(G166) );
  NAND2_X1 U723 ( .A1(G48), .A2(n647), .ZN(n635) );
  XNOR2_X1 U724 ( .A(n635), .B(KEYINPUT84), .ZN(n645) );
  NAND2_X1 U725 ( .A1(G73), .A2(n636), .ZN(n637) );
  XNOR2_X1 U726 ( .A(n637), .B(KEYINPUT2), .ZN(n640) );
  NAND2_X1 U727 ( .A1(n638), .A2(G86), .ZN(n639) );
  NAND2_X1 U728 ( .A1(n640), .A2(n639), .ZN(n643) );
  NAND2_X1 U729 ( .A1(G61), .A2(n652), .ZN(n641) );
  XNOR2_X1 U730 ( .A(KEYINPUT83), .B(n641), .ZN(n642) );
  NOR2_X1 U731 ( .A1(n643), .A2(n642), .ZN(n644) );
  NAND2_X1 U732 ( .A1(n645), .A2(n644), .ZN(G305) );
  NAND2_X1 U733 ( .A1(G651), .A2(G74), .ZN(n646) );
  XOR2_X1 U734 ( .A(KEYINPUT81), .B(n646), .Z(n649) );
  NAND2_X1 U735 ( .A1(n647), .A2(G49), .ZN(n648) );
  NAND2_X1 U736 ( .A1(n649), .A2(n648), .ZN(n650) );
  XNOR2_X1 U737 ( .A(KEYINPUT82), .B(n650), .ZN(n651) );
  NOR2_X1 U738 ( .A1(n652), .A2(n651), .ZN(n655) );
  NAND2_X1 U739 ( .A1(n653), .A2(G87), .ZN(n654) );
  NAND2_X1 U740 ( .A1(n655), .A2(n654), .ZN(G288) );
  XOR2_X1 U741 ( .A(KEYINPUT19), .B(KEYINPUT88), .Z(n657) );
  XOR2_X1 U742 ( .A(G299), .B(KEYINPUT87), .Z(n656) );
  XNOR2_X1 U743 ( .A(n657), .B(n656), .ZN(n658) );
  XOR2_X1 U744 ( .A(n666), .B(n658), .Z(n660) );
  XOR2_X1 U745 ( .A(G290), .B(G166), .Z(n659) );
  XNOR2_X1 U746 ( .A(n660), .B(n659), .ZN(n661) );
  XNOR2_X1 U747 ( .A(n661), .B(G305), .ZN(n662) );
  XNOR2_X1 U748 ( .A(n662), .B(G288), .ZN(n907) );
  XOR2_X1 U749 ( .A(n907), .B(KEYINPUT89), .Z(n663) );
  XNOR2_X1 U750 ( .A(n664), .B(n663), .ZN(n665) );
  NAND2_X1 U751 ( .A1(n665), .A2(G868), .ZN(n669) );
  NAND2_X1 U752 ( .A1(n667), .A2(n666), .ZN(n668) );
  NAND2_X1 U753 ( .A1(n669), .A2(n668), .ZN(G295) );
  NAND2_X1 U754 ( .A1(G2078), .A2(G2084), .ZN(n670) );
  XOR2_X1 U755 ( .A(KEYINPUT20), .B(n670), .Z(n671) );
  NAND2_X1 U756 ( .A1(G2090), .A2(n671), .ZN(n672) );
  XNOR2_X1 U757 ( .A(KEYINPUT21), .B(n672), .ZN(n673) );
  NAND2_X1 U758 ( .A1(n673), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U759 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U760 ( .A1(G236), .A2(G238), .ZN(n675) );
  NOR2_X1 U761 ( .A1(G235), .A2(G237), .ZN(n674) );
  NAND2_X1 U762 ( .A1(n675), .A2(n674), .ZN(n676) );
  XNOR2_X1 U763 ( .A(KEYINPUT90), .B(n676), .ZN(n838) );
  NAND2_X1 U764 ( .A1(G567), .A2(n838), .ZN(n681) );
  NOR2_X1 U765 ( .A1(G220), .A2(G219), .ZN(n677) );
  XOR2_X1 U766 ( .A(KEYINPUT22), .B(n677), .Z(n678) );
  NOR2_X1 U767 ( .A1(G218), .A2(n678), .ZN(n679) );
  NAND2_X1 U768 ( .A1(G96), .A2(n679), .ZN(n837) );
  NAND2_X1 U769 ( .A1(G2106), .A2(n837), .ZN(n680) );
  NAND2_X1 U770 ( .A1(n681), .A2(n680), .ZN(n682) );
  XOR2_X1 U771 ( .A(KEYINPUT91), .B(n682), .Z(n861) );
  NAND2_X1 U772 ( .A1(G661), .A2(G483), .ZN(n683) );
  NOR2_X1 U773 ( .A1(n861), .A2(n683), .ZN(n836) );
  NAND2_X1 U774 ( .A1(n836), .A2(G36), .ZN(G176) );
  INV_X1 U775 ( .A(G166), .ZN(G303) );
  NAND2_X1 U776 ( .A1(G160), .A2(G40), .ZN(n718) );
  INV_X1 U777 ( .A(n718), .ZN(n687) );
  NAND2_X1 U778 ( .A1(n717), .A2(n687), .ZN(n715) );
  INV_X1 U779 ( .A(n715), .ZN(n829) );
  NAND2_X1 U780 ( .A1(G104), .A2(n888), .ZN(n689) );
  NAND2_X1 U781 ( .A1(G140), .A2(n889), .ZN(n688) );
  NAND2_X1 U782 ( .A1(n689), .A2(n688), .ZN(n690) );
  XNOR2_X1 U783 ( .A(KEYINPUT34), .B(n690), .ZN(n695) );
  NAND2_X1 U784 ( .A1(G116), .A2(n884), .ZN(n692) );
  NAND2_X1 U785 ( .A1(G128), .A2(n885), .ZN(n691) );
  NAND2_X1 U786 ( .A1(n692), .A2(n691), .ZN(n693) );
  XOR2_X1 U787 ( .A(KEYINPUT35), .B(n693), .Z(n694) );
  NOR2_X1 U788 ( .A1(n695), .A2(n694), .ZN(n696) );
  XNOR2_X1 U789 ( .A(KEYINPUT36), .B(n696), .ZN(n883) );
  XOR2_X1 U790 ( .A(G2067), .B(KEYINPUT37), .Z(n697) );
  XNOR2_X1 U791 ( .A(KEYINPUT93), .B(n697), .ZN(n820) );
  NOR2_X1 U792 ( .A1(n883), .A2(n820), .ZN(n997) );
  NAND2_X1 U793 ( .A1(n829), .A2(n997), .ZN(n826) );
  XOR2_X1 U794 ( .A(KEYINPUT96), .B(G1991), .Z(n961) );
  NAND2_X1 U795 ( .A1(G107), .A2(n884), .ZN(n699) );
  NAND2_X1 U796 ( .A1(G119), .A2(n885), .ZN(n698) );
  NAND2_X1 U797 ( .A1(n699), .A2(n698), .ZN(n704) );
  NAND2_X1 U798 ( .A1(G95), .A2(n888), .ZN(n701) );
  NAND2_X1 U799 ( .A1(G131), .A2(n889), .ZN(n700) );
  NAND2_X1 U800 ( .A1(n701), .A2(n700), .ZN(n702) );
  XNOR2_X1 U801 ( .A(KEYINPUT94), .B(n702), .ZN(n703) );
  NOR2_X1 U802 ( .A1(n704), .A2(n703), .ZN(n705) );
  XOR2_X1 U803 ( .A(n705), .B(KEYINPUT95), .Z(n898) );
  NOR2_X1 U804 ( .A1(n961), .A2(n898), .ZN(n714) );
  NAND2_X1 U805 ( .A1(G117), .A2(n884), .ZN(n707) );
  NAND2_X1 U806 ( .A1(G141), .A2(n889), .ZN(n706) );
  NAND2_X1 U807 ( .A1(n707), .A2(n706), .ZN(n710) );
  NAND2_X1 U808 ( .A1(n888), .A2(G105), .ZN(n708) );
  XOR2_X1 U809 ( .A(KEYINPUT38), .B(n708), .Z(n709) );
  NOR2_X1 U810 ( .A1(n710), .A2(n709), .ZN(n712) );
  NAND2_X1 U811 ( .A1(G129), .A2(n885), .ZN(n711) );
  NAND2_X1 U812 ( .A1(n712), .A2(n711), .ZN(n873) );
  AND2_X1 U813 ( .A1(n873), .A2(G1996), .ZN(n713) );
  NOR2_X1 U814 ( .A1(n714), .A2(n713), .ZN(n1000) );
  NOR2_X1 U815 ( .A1(n1000), .A2(n715), .ZN(n823) );
  INV_X1 U816 ( .A(n823), .ZN(n716) );
  NAND2_X1 U817 ( .A1(n826), .A2(n716), .ZN(n817) );
  NOR2_X2 U818 ( .A1(n718), .A2(n717), .ZN(n746) );
  NAND2_X1 U819 ( .A1(n736), .A2(G8), .ZN(n720) );
  NOR2_X1 U820 ( .A1(n811), .A2(G1966), .ZN(n780) );
  INV_X1 U821 ( .A(G8), .ZN(n721) );
  NOR2_X1 U822 ( .A1(G2084), .A2(n763), .ZN(n777) );
  OR2_X1 U823 ( .A1(n721), .A2(n777), .ZN(n722) );
  OR2_X1 U824 ( .A1(n780), .A2(n722), .ZN(n723) );
  NOR2_X1 U825 ( .A1(n724), .A2(G168), .ZN(n728) );
  NAND2_X1 U826 ( .A1(G1961), .A2(n763), .ZN(n726) );
  XOR2_X1 U827 ( .A(KEYINPUT25), .B(G2078), .Z(n960) );
  NAND2_X1 U828 ( .A1(n746), .A2(n960), .ZN(n725) );
  NAND2_X1 U829 ( .A1(n726), .A2(n725), .ZN(n759) );
  AND2_X1 U830 ( .A1(G301), .A2(n759), .ZN(n727) );
  NOR2_X1 U831 ( .A1(n728), .A2(n727), .ZN(n729) );
  XNOR2_X1 U832 ( .A(n729), .B(KEYINPUT31), .ZN(n779) );
  XNOR2_X1 U833 ( .A(KEYINPUT66), .B(KEYINPUT26), .ZN(n737) );
  NOR2_X1 U834 ( .A1(G1996), .A2(n737), .ZN(n730) );
  NOR2_X1 U835 ( .A1(n730), .A2(n1012), .ZN(n734) );
  NAND2_X1 U836 ( .A1(G1348), .A2(n736), .ZN(n732) );
  NAND2_X1 U837 ( .A1(G2067), .A2(n746), .ZN(n731) );
  NAND2_X1 U838 ( .A1(n732), .A2(n731), .ZN(n743) );
  NAND2_X1 U839 ( .A1(n743), .A2(n905), .ZN(n733) );
  NAND2_X1 U840 ( .A1(n734), .A2(n733), .ZN(n742) );
  INV_X1 U841 ( .A(G1341), .ZN(n917) );
  NAND2_X1 U842 ( .A1(n917), .A2(n737), .ZN(n735) );
  NAND2_X1 U843 ( .A1(n735), .A2(n763), .ZN(n740) );
  INV_X1 U844 ( .A(G1996), .ZN(n840) );
  NOR2_X1 U845 ( .A1(n840), .A2(n736), .ZN(n738) );
  NAND2_X1 U846 ( .A1(n738), .A2(n737), .ZN(n739) );
  NAND2_X1 U847 ( .A1(n740), .A2(n739), .ZN(n741) );
  NOR2_X1 U848 ( .A1(n742), .A2(n741), .ZN(n745) );
  NOR2_X1 U849 ( .A1(n743), .A2(n905), .ZN(n744) );
  NOR2_X1 U850 ( .A1(n745), .A2(n744), .ZN(n751) );
  INV_X1 U851 ( .A(G299), .ZN(n753) );
  NAND2_X1 U852 ( .A1(n746), .A2(G2072), .ZN(n747) );
  XNOR2_X1 U853 ( .A(n747), .B(KEYINPUT27), .ZN(n749) );
  INV_X1 U854 ( .A(G1956), .ZN(n839) );
  NOR2_X1 U855 ( .A1(n839), .A2(n746), .ZN(n748) );
  NOR2_X1 U856 ( .A1(n749), .A2(n748), .ZN(n752) );
  NAND2_X1 U857 ( .A1(n753), .A2(n752), .ZN(n750) );
  NAND2_X1 U858 ( .A1(n751), .A2(n750), .ZN(n757) );
  NOR2_X1 U859 ( .A1(n753), .A2(n752), .ZN(n755) );
  XNOR2_X1 U860 ( .A(KEYINPUT28), .B(KEYINPUT99), .ZN(n754) );
  XNOR2_X1 U861 ( .A(n755), .B(n754), .ZN(n756) );
  NAND2_X1 U862 ( .A1(n757), .A2(n756), .ZN(n758) );
  XNOR2_X1 U863 ( .A(n758), .B(KEYINPUT29), .ZN(n761) );
  NOR2_X1 U864 ( .A1(G301), .A2(n759), .ZN(n760) );
  XNOR2_X1 U865 ( .A(n762), .B(KEYINPUT100), .ZN(n778) );
  NOR2_X1 U866 ( .A1(G1971), .A2(n811), .ZN(n765) );
  NOR2_X1 U867 ( .A1(G2090), .A2(n763), .ZN(n764) );
  NOR2_X1 U868 ( .A1(n765), .A2(n764), .ZN(n766) );
  NAND2_X1 U869 ( .A1(G303), .A2(n766), .ZN(n767) );
  NOR2_X1 U870 ( .A1(n721), .A2(n767), .ZN(n770) );
  NOR2_X1 U871 ( .A1(n779), .A2(n768), .ZN(n772) );
  AND2_X1 U872 ( .A1(G286), .A2(G8), .ZN(n769) );
  NOR2_X1 U873 ( .A1(n770), .A2(n769), .ZN(n771) );
  XNOR2_X1 U874 ( .A(KEYINPUT32), .B(KEYINPUT102), .ZN(n773) );
  NAND2_X1 U875 ( .A1(G1976), .A2(G288), .ZN(n1019) );
  INV_X1 U876 ( .A(n1019), .ZN(n775) );
  OR2_X1 U877 ( .A1(n811), .A2(n775), .ZN(n787) );
  INV_X1 U878 ( .A(n787), .ZN(n776) );
  AND2_X1 U879 ( .A1(n805), .A2(n776), .ZN(n785) );
  AND2_X1 U880 ( .A1(n777), .A2(G8), .ZN(n784) );
  NOR2_X1 U881 ( .A1(n779), .A2(n778), .ZN(n781) );
  NOR2_X1 U882 ( .A1(n781), .A2(n780), .ZN(n782) );
  XNOR2_X1 U883 ( .A(n782), .B(KEYINPUT101), .ZN(n783) );
  OR2_X1 U884 ( .A1(n784), .A2(n783), .ZN(n806) );
  NAND2_X1 U885 ( .A1(n785), .A2(n806), .ZN(n789) );
  NOR2_X1 U886 ( .A1(G1976), .A2(G288), .ZN(n793) );
  NOR2_X1 U887 ( .A1(G303), .A2(G1971), .ZN(n786) );
  NOR2_X1 U888 ( .A1(n793), .A2(n786), .ZN(n1015) );
  OR2_X1 U889 ( .A1(n787), .A2(n1015), .ZN(n788) );
  NAND2_X1 U890 ( .A1(n789), .A2(n788), .ZN(n791) );
  XNOR2_X1 U891 ( .A(n791), .B(n790), .ZN(n792) );
  INV_X1 U892 ( .A(KEYINPUT33), .ZN(n795) );
  NAND2_X1 U893 ( .A1(n792), .A2(n795), .ZN(n800) );
  INV_X1 U894 ( .A(n811), .ZN(n803) );
  NAND2_X1 U895 ( .A1(n803), .A2(n793), .ZN(n794) );
  NOR2_X1 U896 ( .A1(n795), .A2(n794), .ZN(n796) );
  XNOR2_X1 U897 ( .A(n796), .B(KEYINPUT103), .ZN(n798) );
  XNOR2_X1 U898 ( .A(G1981), .B(G305), .ZN(n1030) );
  INV_X1 U899 ( .A(n1030), .ZN(n797) );
  AND2_X1 U900 ( .A1(n798), .A2(n797), .ZN(n799) );
  AND2_X1 U901 ( .A1(n800), .A2(n799), .ZN(n815) );
  NOR2_X1 U902 ( .A1(G1981), .A2(G305), .ZN(n801) );
  XNOR2_X1 U903 ( .A(n801), .B(KEYINPUT98), .ZN(n802) );
  XNOR2_X1 U904 ( .A(n802), .B(KEYINPUT24), .ZN(n804) );
  NAND2_X1 U905 ( .A1(n804), .A2(n803), .ZN(n813) );
  NAND2_X1 U906 ( .A1(n806), .A2(n805), .ZN(n809) );
  NOR2_X1 U907 ( .A1(G2090), .A2(G303), .ZN(n807) );
  NAND2_X1 U908 ( .A1(G8), .A2(n807), .ZN(n808) );
  NAND2_X1 U909 ( .A1(n809), .A2(n808), .ZN(n810) );
  NAND2_X1 U910 ( .A1(n811), .A2(n810), .ZN(n812) );
  NAND2_X1 U911 ( .A1(n813), .A2(n812), .ZN(n814) );
  NOR2_X1 U912 ( .A1(n815), .A2(n814), .ZN(n816) );
  NOR2_X1 U913 ( .A1(n817), .A2(n816), .ZN(n819) );
  XNOR2_X1 U914 ( .A(G1986), .B(G290), .ZN(n1018) );
  NAND2_X1 U915 ( .A1(n1018), .A2(n829), .ZN(n818) );
  NAND2_X1 U916 ( .A1(n819), .A2(n818), .ZN(n832) );
  NAND2_X1 U917 ( .A1(n883), .A2(n820), .ZN(n996) );
  NOR2_X1 U918 ( .A1(G1996), .A2(n873), .ZN(n991) );
  NOR2_X1 U919 ( .A1(G1986), .A2(G290), .ZN(n821) );
  AND2_X1 U920 ( .A1(n961), .A2(n898), .ZN(n986) );
  NOR2_X1 U921 ( .A1(n821), .A2(n986), .ZN(n822) );
  NOR2_X1 U922 ( .A1(n823), .A2(n822), .ZN(n824) );
  NOR2_X1 U923 ( .A1(n991), .A2(n824), .ZN(n825) );
  XNOR2_X1 U924 ( .A(n825), .B(KEYINPUT39), .ZN(n827) );
  NAND2_X1 U925 ( .A1(n827), .A2(n826), .ZN(n828) );
  NAND2_X1 U926 ( .A1(n996), .A2(n828), .ZN(n830) );
  NAND2_X1 U927 ( .A1(n830), .A2(n829), .ZN(n831) );
  NAND2_X1 U928 ( .A1(n832), .A2(n831), .ZN(n833) );
  XNOR2_X1 U929 ( .A(n833), .B(KEYINPUT40), .ZN(G329) );
  NAND2_X1 U930 ( .A1(G2106), .A2(n930), .ZN(G217) );
  AND2_X1 U931 ( .A1(G15), .A2(G2), .ZN(n834) );
  NAND2_X1 U932 ( .A1(G661), .A2(n834), .ZN(G259) );
  NAND2_X1 U933 ( .A1(G3), .A2(G1), .ZN(n835) );
  NAND2_X1 U934 ( .A1(n836), .A2(n835), .ZN(G188) );
  INV_X1 U936 ( .A(G96), .ZN(G221) );
  NOR2_X1 U937 ( .A1(n838), .A2(n837), .ZN(G325) );
  INV_X1 U938 ( .A(G325), .ZN(G261) );
  XNOR2_X1 U939 ( .A(G1991), .B(G2474), .ZN(n850) );
  XNOR2_X1 U940 ( .A(n839), .B(G1961), .ZN(n842) );
  XOR2_X1 U941 ( .A(n840), .B(G1986), .Z(n841) );
  XNOR2_X1 U942 ( .A(n842), .B(n841), .ZN(n846) );
  XOR2_X1 U943 ( .A(G1976), .B(G1981), .Z(n844) );
  XNOR2_X1 U944 ( .A(G1971), .B(G1966), .ZN(n843) );
  XNOR2_X1 U945 ( .A(n844), .B(n843), .ZN(n845) );
  XOR2_X1 U946 ( .A(n846), .B(n845), .Z(n848) );
  XNOR2_X1 U947 ( .A(KEYINPUT106), .B(KEYINPUT41), .ZN(n847) );
  XNOR2_X1 U948 ( .A(n848), .B(n847), .ZN(n849) );
  XNOR2_X1 U949 ( .A(n850), .B(n849), .ZN(G229) );
  XOR2_X1 U950 ( .A(KEYINPUT42), .B(G2084), .Z(n852) );
  XNOR2_X1 U951 ( .A(G2067), .B(G2090), .ZN(n851) );
  XNOR2_X1 U952 ( .A(n852), .B(n851), .ZN(n853) );
  XOR2_X1 U953 ( .A(n853), .B(G2096), .Z(n855) );
  XNOR2_X1 U954 ( .A(G2078), .B(G2072), .ZN(n854) );
  XNOR2_X1 U955 ( .A(n855), .B(n854), .ZN(n860) );
  XOR2_X1 U956 ( .A(KEYINPUT43), .B(KEYINPUT105), .Z(n858) );
  XOR2_X1 U957 ( .A(G2678), .B(n856), .Z(n857) );
  XNOR2_X1 U958 ( .A(n858), .B(n857), .ZN(n859) );
  XOR2_X1 U959 ( .A(n860), .B(n859), .Z(G227) );
  INV_X1 U960 ( .A(n861), .ZN(G319) );
  NAND2_X1 U961 ( .A1(G112), .A2(n884), .ZN(n863) );
  NAND2_X1 U962 ( .A1(G100), .A2(n888), .ZN(n862) );
  NAND2_X1 U963 ( .A1(n863), .A2(n862), .ZN(n869) );
  NAND2_X1 U964 ( .A1(G124), .A2(n885), .ZN(n864) );
  XNOR2_X1 U965 ( .A(n864), .B(KEYINPUT44), .ZN(n866) );
  NAND2_X1 U966 ( .A1(G136), .A2(n889), .ZN(n865) );
  NAND2_X1 U967 ( .A1(n866), .A2(n865), .ZN(n867) );
  XOR2_X1 U968 ( .A(KEYINPUT107), .B(n867), .Z(n868) );
  NOR2_X1 U969 ( .A1(n869), .A2(n868), .ZN(G162) );
  XOR2_X1 U970 ( .A(KEYINPUT109), .B(KEYINPUT46), .Z(n871) );
  XNOR2_X1 U971 ( .A(n985), .B(KEYINPUT48), .ZN(n870) );
  XNOR2_X1 U972 ( .A(n871), .B(n870), .ZN(n872) );
  XOR2_X1 U973 ( .A(n873), .B(n872), .Z(n902) );
  NAND2_X1 U974 ( .A1(G115), .A2(n884), .ZN(n875) );
  NAND2_X1 U975 ( .A1(G127), .A2(n885), .ZN(n874) );
  NAND2_X1 U976 ( .A1(n875), .A2(n874), .ZN(n876) );
  XNOR2_X1 U977 ( .A(n876), .B(KEYINPUT47), .ZN(n878) );
  NAND2_X1 U978 ( .A1(G139), .A2(n889), .ZN(n877) );
  NAND2_X1 U979 ( .A1(n878), .A2(n877), .ZN(n881) );
  NAND2_X1 U980 ( .A1(n888), .A2(G103), .ZN(n879) );
  XOR2_X1 U981 ( .A(KEYINPUT110), .B(n879), .Z(n880) );
  NOR2_X1 U982 ( .A1(n881), .A2(n880), .ZN(n981) );
  XOR2_X1 U983 ( .A(G164), .B(n981), .Z(n882) );
  XNOR2_X1 U984 ( .A(n883), .B(n882), .ZN(n897) );
  NAND2_X1 U985 ( .A1(G118), .A2(n884), .ZN(n887) );
  NAND2_X1 U986 ( .A1(G130), .A2(n885), .ZN(n886) );
  NAND2_X1 U987 ( .A1(n887), .A2(n886), .ZN(n895) );
  NAND2_X1 U988 ( .A1(G106), .A2(n888), .ZN(n891) );
  NAND2_X1 U989 ( .A1(G142), .A2(n889), .ZN(n890) );
  NAND2_X1 U990 ( .A1(n891), .A2(n890), .ZN(n892) );
  XOR2_X1 U991 ( .A(KEYINPUT45), .B(n892), .Z(n893) );
  XNOR2_X1 U992 ( .A(KEYINPUT108), .B(n893), .ZN(n894) );
  NOR2_X1 U993 ( .A1(n895), .A2(n894), .ZN(n896) );
  XOR2_X1 U994 ( .A(n897), .B(n896), .Z(n900) );
  XNOR2_X1 U995 ( .A(G160), .B(n898), .ZN(n899) );
  XNOR2_X1 U996 ( .A(n900), .B(n899), .ZN(n901) );
  XNOR2_X1 U997 ( .A(n902), .B(n901), .ZN(n903) );
  XNOR2_X1 U998 ( .A(n903), .B(G162), .ZN(n904) );
  NOR2_X1 U999 ( .A1(G37), .A2(n904), .ZN(G395) );
  XOR2_X1 U1000 ( .A(G301), .B(n905), .Z(n906) );
  XNOR2_X1 U1001 ( .A(KEYINPUT111), .B(n906), .ZN(n909) );
  XNOR2_X1 U1002 ( .A(n1012), .B(n907), .ZN(n908) );
  XNOR2_X1 U1003 ( .A(n909), .B(n908), .ZN(n910) );
  XNOR2_X1 U1004 ( .A(n910), .B(G286), .ZN(n911) );
  NOR2_X1 U1005 ( .A1(G37), .A2(n911), .ZN(G397) );
  XNOR2_X1 U1006 ( .A(KEYINPUT49), .B(KEYINPUT112), .ZN(n913) );
  NOR2_X1 U1007 ( .A1(G229), .A2(G227), .ZN(n912) );
  XNOR2_X1 U1008 ( .A(n913), .B(n912), .ZN(n926) );
  XOR2_X1 U1009 ( .A(G2438), .B(G2435), .Z(n915) );
  XNOR2_X1 U1010 ( .A(G2443), .B(G2430), .ZN(n914) );
  XNOR2_X1 U1011 ( .A(n915), .B(n914), .ZN(n916) );
  XOR2_X1 U1012 ( .A(n916), .B(G2454), .Z(n919) );
  XOR2_X1 U1013 ( .A(n917), .B(G1348), .Z(n918) );
  XNOR2_X1 U1014 ( .A(n919), .B(n918), .ZN(n923) );
  XOR2_X1 U1015 ( .A(G2451), .B(G2427), .Z(n921) );
  XNOR2_X1 U1016 ( .A(KEYINPUT104), .B(G2446), .ZN(n920) );
  XNOR2_X1 U1017 ( .A(n921), .B(n920), .ZN(n922) );
  XOR2_X1 U1018 ( .A(n923), .B(n922), .Z(n924) );
  NAND2_X1 U1019 ( .A1(G14), .A2(n924), .ZN(n929) );
  NAND2_X1 U1020 ( .A1(G319), .A2(n929), .ZN(n925) );
  NOR2_X1 U1021 ( .A1(n926), .A2(n925), .ZN(n928) );
  NOR2_X1 U1022 ( .A1(G395), .A2(G397), .ZN(n927) );
  NAND2_X1 U1023 ( .A1(n928), .A2(n927), .ZN(G225) );
  INV_X1 U1024 ( .A(G225), .ZN(G308) );
  INV_X1 U1025 ( .A(n929), .ZN(G401) );
  INV_X1 U1026 ( .A(n930), .ZN(G223) );
  XOR2_X1 U1027 ( .A(G1986), .B(G24), .Z(n934) );
  XNOR2_X1 U1028 ( .A(G1971), .B(G22), .ZN(n932) );
  XNOR2_X1 U1029 ( .A(G23), .B(G1976), .ZN(n931) );
  NOR2_X1 U1030 ( .A1(n932), .A2(n931), .ZN(n933) );
  NAND2_X1 U1031 ( .A1(n934), .A2(n933), .ZN(n936) );
  XOR2_X1 U1032 ( .A(KEYINPUT126), .B(KEYINPUT58), .Z(n935) );
  XNOR2_X1 U1033 ( .A(n936), .B(n935), .ZN(n953) );
  XNOR2_X1 U1034 ( .A(G1961), .B(G5), .ZN(n951) );
  XNOR2_X1 U1035 ( .A(KEYINPUT124), .B(KEYINPUT60), .ZN(n946) );
  XNOR2_X1 U1036 ( .A(KEYINPUT123), .B(G1981), .ZN(n937) );
  XNOR2_X1 U1037 ( .A(n937), .B(G6), .ZN(n944) );
  XOR2_X1 U1038 ( .A(G1348), .B(KEYINPUT59), .Z(n938) );
  XNOR2_X1 U1039 ( .A(G4), .B(n938), .ZN(n942) );
  XOR2_X1 U1040 ( .A(G1956), .B(G20), .Z(n940) );
  XOR2_X1 U1041 ( .A(G1341), .B(G19), .Z(n939) );
  NAND2_X1 U1042 ( .A1(n940), .A2(n939), .ZN(n941) );
  NOR2_X1 U1043 ( .A1(n942), .A2(n941), .ZN(n943) );
  NAND2_X1 U1044 ( .A1(n944), .A2(n943), .ZN(n945) );
  XNOR2_X1 U1045 ( .A(n946), .B(n945), .ZN(n948) );
  XNOR2_X1 U1046 ( .A(G21), .B(G1966), .ZN(n947) );
  NOR2_X1 U1047 ( .A1(n948), .A2(n947), .ZN(n949) );
  XNOR2_X1 U1048 ( .A(KEYINPUT125), .B(n949), .ZN(n950) );
  NOR2_X1 U1049 ( .A1(n951), .A2(n950), .ZN(n952) );
  NAND2_X1 U1050 ( .A1(n953), .A2(n952), .ZN(n954) );
  XNOR2_X1 U1051 ( .A(n954), .B(KEYINPUT127), .ZN(n955) );
  XOR2_X1 U1052 ( .A(KEYINPUT61), .B(n955), .Z(n956) );
  NOR2_X1 U1053 ( .A1(G16), .A2(n956), .ZN(n980) );
  XOR2_X1 U1054 ( .A(KEYINPUT55), .B(KEYINPUT116), .Z(n1007) );
  XNOR2_X1 U1055 ( .A(G2067), .B(G26), .ZN(n958) );
  XNOR2_X1 U1056 ( .A(G33), .B(G2072), .ZN(n957) );
  NOR2_X1 U1057 ( .A1(n958), .A2(n957), .ZN(n967) );
  XOR2_X1 U1058 ( .A(G32), .B(G1996), .Z(n959) );
  NAND2_X1 U1059 ( .A1(n959), .A2(G28), .ZN(n965) );
  XOR2_X1 U1060 ( .A(n960), .B(G27), .Z(n963) );
  XNOR2_X1 U1061 ( .A(n961), .B(G25), .ZN(n962) );
  NAND2_X1 U1062 ( .A1(n963), .A2(n962), .ZN(n964) );
  NOR2_X1 U1063 ( .A1(n965), .A2(n964), .ZN(n966) );
  NAND2_X1 U1064 ( .A1(n967), .A2(n966), .ZN(n968) );
  XNOR2_X1 U1065 ( .A(n968), .B(KEYINPUT53), .ZN(n971) );
  XOR2_X1 U1066 ( .A(G2084), .B(G34), .Z(n969) );
  XNOR2_X1 U1067 ( .A(KEYINPUT54), .B(n969), .ZN(n970) );
  NAND2_X1 U1068 ( .A1(n971), .A2(n970), .ZN(n973) );
  XNOR2_X1 U1069 ( .A(G35), .B(G2090), .ZN(n972) );
  NOR2_X1 U1070 ( .A1(n973), .A2(n972), .ZN(n974) );
  XNOR2_X1 U1071 ( .A(n1007), .B(n974), .ZN(n975) );
  NOR2_X1 U1072 ( .A1(G29), .A2(n975), .ZN(n976) );
  XNOR2_X1 U1073 ( .A(KEYINPUT117), .B(n976), .ZN(n977) );
  NAND2_X1 U1074 ( .A1(n977), .A2(G11), .ZN(n978) );
  XNOR2_X1 U1075 ( .A(n978), .B(KEYINPUT118), .ZN(n979) );
  NOR2_X1 U1076 ( .A1(n980), .A2(n979), .ZN(n1011) );
  XOR2_X1 U1077 ( .A(G2072), .B(n981), .Z(n983) );
  XOR2_X1 U1078 ( .A(G164), .B(G2078), .Z(n982) );
  NOR2_X1 U1079 ( .A1(n983), .A2(n982), .ZN(n984) );
  XOR2_X1 U1080 ( .A(KEYINPUT50), .B(n984), .Z(n1005) );
  XNOR2_X1 U1081 ( .A(G160), .B(G2084), .ZN(n988) );
  NOR2_X1 U1082 ( .A1(n986), .A2(n985), .ZN(n987) );
  NAND2_X1 U1083 ( .A1(n988), .A2(n987), .ZN(n989) );
  XNOR2_X1 U1084 ( .A(KEYINPUT113), .B(n989), .ZN(n995) );
  XOR2_X1 U1085 ( .A(G2090), .B(G162), .Z(n990) );
  XNOR2_X1 U1086 ( .A(KEYINPUT114), .B(n990), .ZN(n992) );
  NOR2_X1 U1087 ( .A1(n992), .A2(n991), .ZN(n993) );
  XOR2_X1 U1088 ( .A(KEYINPUT51), .B(n993), .Z(n994) );
  NAND2_X1 U1089 ( .A1(n995), .A2(n994), .ZN(n1002) );
  INV_X1 U1090 ( .A(n996), .ZN(n998) );
  NOR2_X1 U1091 ( .A1(n998), .A2(n997), .ZN(n999) );
  NAND2_X1 U1092 ( .A1(n1000), .A2(n999), .ZN(n1001) );
  NOR2_X1 U1093 ( .A1(n1002), .A2(n1001), .ZN(n1003) );
  XNOR2_X1 U1094 ( .A(KEYINPUT115), .B(n1003), .ZN(n1004) );
  NOR2_X1 U1095 ( .A1(n1005), .A2(n1004), .ZN(n1006) );
  XNOR2_X1 U1096 ( .A(KEYINPUT52), .B(n1006), .ZN(n1008) );
  NAND2_X1 U1097 ( .A1(n1008), .A2(n1007), .ZN(n1009) );
  NAND2_X1 U1098 ( .A1(n1009), .A2(G29), .ZN(n1010) );
  NAND2_X1 U1099 ( .A1(n1011), .A2(n1010), .ZN(n1040) );
  XOR2_X1 U1100 ( .A(KEYINPUT56), .B(G16), .Z(n1038) );
  XOR2_X1 U1101 ( .A(n1012), .B(G1341), .Z(n1014) );
  NAND2_X1 U1102 ( .A1(G1971), .A2(G303), .ZN(n1013) );
  NAND2_X1 U1103 ( .A1(n1014), .A2(n1013), .ZN(n1035) );
  XOR2_X1 U1104 ( .A(G299), .B(G1956), .Z(n1016) );
  NAND2_X1 U1105 ( .A1(n1016), .A2(n1015), .ZN(n1017) );
  NOR2_X1 U1106 ( .A1(n1018), .A2(n1017), .ZN(n1020) );
  NAND2_X1 U1107 ( .A1(n1020), .A2(n1019), .ZN(n1027) );
  XNOR2_X1 U1108 ( .A(G1348), .B(KEYINPUT120), .ZN(n1022) );
  XOR2_X1 U1109 ( .A(n1022), .B(n1021), .Z(n1024) );
  XOR2_X1 U1110 ( .A(G1961), .B(G171), .Z(n1023) );
  NOR2_X1 U1111 ( .A1(n1024), .A2(n1023), .ZN(n1025) );
  XNOR2_X1 U1112 ( .A(n1025), .B(KEYINPUT121), .ZN(n1026) );
  NOR2_X1 U1113 ( .A1(n1027), .A2(n1026), .ZN(n1033) );
  XNOR2_X1 U1114 ( .A(G168), .B(G1966), .ZN(n1028) );
  XNOR2_X1 U1115 ( .A(n1028), .B(KEYINPUT119), .ZN(n1029) );
  NOR2_X1 U1116 ( .A1(n1030), .A2(n1029), .ZN(n1031) );
  XOR2_X1 U1117 ( .A(KEYINPUT57), .B(n1031), .Z(n1032) );
  NAND2_X1 U1118 ( .A1(n1033), .A2(n1032), .ZN(n1034) );
  NOR2_X1 U1119 ( .A1(n1035), .A2(n1034), .ZN(n1036) );
  XNOR2_X1 U1120 ( .A(KEYINPUT122), .B(n1036), .ZN(n1037) );
  NOR2_X1 U1121 ( .A1(n1038), .A2(n1037), .ZN(n1039) );
  NOR2_X1 U1122 ( .A1(n1040), .A2(n1039), .ZN(n1041) );
  XOR2_X1 U1123 ( .A(n1041), .B(KEYINPUT62), .Z(G150) );
  INV_X1 U1124 ( .A(G150), .ZN(G311) );
endmodule

