

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361,
         n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372,
         n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383,
         n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394,
         n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405,
         n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416,
         n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427,
         n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438,
         n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449,
         n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460,
         n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471,
         n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482,
         n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493,
         n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504,
         n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515,
         n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526,
         n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537,
         n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
         n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559,
         n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570,
         n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581,
         n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592,
         n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603,
         n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614,
         n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625,
         n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636,
         n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647,
         n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658,
         n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669,
         n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680,
         n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691,
         n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702,
         n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713,
         n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724,
         n725, n726, n727, n728, n729, n730, n731;

  XNOR2_X1 U372 ( .A(n539), .B(n538), .ZN(n574) );
  XOR2_X1 U373 ( .A(n617), .B(n616), .Z(n351) );
  AND2_X2 U374 ( .A1(n389), .A2(n685), .ZN(n700) );
  XNOR2_X2 U375 ( .A(n527), .B(n526), .ZN(n730) );
  NOR2_X2 U376 ( .A1(n540), .A2(n676), .ZN(n527) );
  XOR2_X2 U377 ( .A(G113), .B(G104), .Z(n499) );
  OR2_X2 U378 ( .A1(n393), .A2(n726), .ZN(n392) );
  XOR2_X2 U379 ( .A(G107), .B(G122), .Z(n511) );
  NOR2_X2 U380 ( .A1(n528), .A2(n490), .ZN(n370) );
  XNOR2_X2 U381 ( .A(n419), .B(G472), .ZN(n650) );
  INV_X2 U382 ( .A(G953), .ZN(n612) );
  XNOR2_X1 U383 ( .A(n559), .B(KEYINPUT87), .ZN(n415) );
  NAND2_X1 U384 ( .A1(n728), .A2(n730), .ZN(n364) );
  XNOR2_X1 U385 ( .A(KEYINPUT10), .B(KEYINPUT67), .ZN(n369) );
  XOR2_X1 U386 ( .A(KEYINPUT4), .B(G146), .Z(n443) );
  XNOR2_X1 U387 ( .A(n565), .B(KEYINPUT75), .ZN(n593) );
  NAND2_X1 U388 ( .A1(n652), .A2(n651), .ZN(n565) );
  XNOR2_X1 U389 ( .A(n557), .B(n377), .ZN(n661) );
  XNOR2_X1 U390 ( .A(n483), .B(KEYINPUT66), .ZN(n564) );
  OR2_X2 U391 ( .A1(n383), .A2(n380), .ZN(n548) );
  XNOR2_X1 U392 ( .A(n440), .B(n359), .ZN(n537) );
  NOR2_X1 U393 ( .A1(n617), .A2(G902), .ZN(n419) );
  XNOR2_X1 U394 ( .A(n420), .B(n448), .ZN(n617) );
  XNOR2_X1 U395 ( .A(n717), .B(n456), .ZN(n416) );
  XNOR2_X1 U396 ( .A(n469), .B(n468), .ZN(n470) );
  XNOR2_X2 U397 ( .A(n502), .B(n461), .ZN(n716) );
  XNOR2_X1 U398 ( .A(n443), .B(n358), .ZN(n378) );
  XNOR2_X1 U399 ( .A(n435), .B(n434), .ZN(n447) );
  INV_X1 U400 ( .A(n369), .ZN(n460) );
  AND2_X2 U401 ( .A1(n389), .A2(n685), .ZN(n352) );
  XNOR2_X1 U402 ( .A(n479), .B(n478), .ZN(n353) );
  XNOR2_X1 U403 ( .A(n479), .B(n478), .ZN(n646) );
  XNOR2_X1 U404 ( .A(n471), .B(n470), .ZN(n702) );
  XNOR2_X1 U405 ( .A(n716), .B(n464), .ZN(n471) );
  NAND2_X1 U406 ( .A1(n608), .A2(n386), .ZN(n385) );
  XNOR2_X2 U407 ( .A(n418), .B(G134), .ZN(n514) );
  XOR2_X1 U408 ( .A(KEYINPUT69), .B(n524), .Z(n544) );
  NAND2_X1 U409 ( .A1(n385), .A2(n384), .ZN(n383) );
  NAND2_X1 U410 ( .A1(n458), .A2(n382), .ZN(n381) );
  XNOR2_X1 U411 ( .A(n373), .B(n447), .ZN(n448) );
  XNOR2_X1 U412 ( .A(n446), .B(n357), .ZN(n373) );
  INV_X1 U413 ( .A(KEYINPUT45), .ZN(n394) );
  XOR2_X1 U414 ( .A(KEYINPUT94), .B(KEYINPUT95), .Z(n475) );
  XNOR2_X1 U415 ( .A(n443), .B(G131), .ZN(n417) );
  XNOR2_X1 U416 ( .A(n392), .B(n424), .ZN(n396) );
  INV_X1 U417 ( .A(KEYINPUT44), .ZN(n424) );
  NAND2_X1 U418 ( .A1(n627), .A2(n731), .ZN(n393) );
  NAND2_X1 U419 ( .A1(n661), .A2(n660), .ZN(n664) );
  XNOR2_X1 U420 ( .A(n482), .B(n481), .ZN(n647) );
  XOR2_X1 U421 ( .A(KEYINPUT77), .B(G110), .Z(n450) );
  XOR2_X1 U422 ( .A(G116), .B(KEYINPUT3), .Z(n435) );
  XOR2_X1 U423 ( .A(KEYINPUT9), .B(KEYINPUT7), .Z(n509) );
  XNOR2_X1 U424 ( .A(n705), .B(n426), .ZN(n690) );
  XNOR2_X1 U425 ( .A(n438), .B(n378), .ZN(n439) );
  XNOR2_X1 U426 ( .A(n370), .B(n491), .ZN(n561) );
  XNOR2_X1 U427 ( .A(n594), .B(KEYINPUT97), .ZN(n657) );
  INV_X1 U428 ( .A(KEYINPUT28), .ZN(n374) );
  XNOR2_X1 U429 ( .A(KEYINPUT0), .B(KEYINPUT88), .ZN(n428) );
  NOR2_X1 U430 ( .A1(n687), .A2(n686), .ZN(n413) );
  INV_X1 U431 ( .A(KEYINPUT86), .ZN(n412) );
  INV_X1 U432 ( .A(KEYINPUT46), .ZN(n408) );
  NOR2_X1 U433 ( .A1(G953), .A2(G237), .ZN(n492) );
  OR2_X1 U434 ( .A1(G237), .A2(G902), .ZN(n441) );
  INV_X1 U435 ( .A(G902), .ZN(n382) );
  NAND2_X1 U436 ( .A1(n386), .A2(G902), .ZN(n384) );
  XNOR2_X1 U437 ( .A(G137), .B(KEYINPUT76), .ZN(n444) );
  XNOR2_X1 U438 ( .A(G902), .B(KEYINPUT15), .ZN(n472) );
  XNOR2_X1 U439 ( .A(G146), .B(G122), .ZN(n495) );
  XNOR2_X1 U440 ( .A(G137), .B(KEYINPUT68), .ZN(n461) );
  XNOR2_X1 U441 ( .A(G101), .B(G104), .ZN(n455) );
  XOR2_X1 U442 ( .A(KEYINPUT18), .B(KEYINPUT80), .Z(n437) );
  XNOR2_X1 U443 ( .A(G125), .B(KEYINPUT17), .ZN(n436) );
  INV_X1 U444 ( .A(G143), .ZN(n431) );
  NAND2_X1 U445 ( .A1(G234), .A2(G237), .ZN(n485) );
  INV_X1 U446 ( .A(KEYINPUT38), .ZN(n377) );
  XNOR2_X1 U447 ( .A(n477), .B(n476), .ZN(n478) );
  XNOR2_X1 U448 ( .A(G146), .B(G110), .ZN(n466) );
  XNOR2_X1 U449 ( .A(G128), .B(G119), .ZN(n463) );
  INV_X1 U450 ( .A(n472), .ZN(n606) );
  NAND2_X1 U451 ( .A1(n388), .A2(n387), .ZN(n685) );
  NOR2_X1 U452 ( .A1(n679), .A2(n682), .ZN(n388) );
  BUF_X1 U453 ( .A(n652), .Z(n371) );
  NOR2_X1 U454 ( .A1(n544), .A2(n422), .ZN(n421) );
  OR2_X1 U455 ( .A1(n620), .A2(n423), .ZN(n422) );
  INV_X1 U456 ( .A(n660), .ZN(n423) );
  XNOR2_X1 U457 ( .A(n427), .B(KEYINPUT22), .ZN(n584) );
  NAND2_X1 U458 ( .A1(n597), .A2(n581), .ZN(n427) );
  NOR2_X1 U459 ( .A1(n484), .A2(n367), .ZN(n366) );
  INV_X1 U460 ( .A(n521), .ZN(n367) );
  INV_X1 U461 ( .A(n650), .ZN(n600) );
  NOR2_X1 U462 ( .A1(n584), .A2(n371), .ZN(n590) );
  XNOR2_X1 U463 ( .A(n425), .B(n355), .ZN(n705) );
  XNOR2_X1 U464 ( .A(n513), .B(n376), .ZN(n698) );
  XNOR2_X1 U465 ( .A(n515), .B(n512), .ZN(n376) );
  NAND2_X1 U466 ( .A1(n700), .A2(G475), .ZN(n694) );
  XNOR2_X1 U467 ( .A(n579), .B(KEYINPUT35), .ZN(n726) );
  XNOR2_X1 U468 ( .A(n596), .B(n595), .ZN(n639) );
  AND2_X1 U469 ( .A1(n411), .A2(n410), .ZN(n689) );
  AND2_X1 U470 ( .A1(n688), .A2(n612), .ZN(n410) );
  XNOR2_X1 U471 ( .A(n413), .B(n412), .ZN(n411) );
  AND2_X1 U472 ( .A1(n650), .A2(n592), .ZN(n354) );
  XNOR2_X1 U473 ( .A(KEYINPUT16), .B(n450), .ZN(n355) );
  BUF_X1 U474 ( .A(n353), .Z(n379) );
  AND2_X1 U475 ( .A1(n729), .A2(n606), .ZN(n356) );
  AND2_X1 U476 ( .A1(n492), .A2(G210), .ZN(n357) );
  AND2_X1 U477 ( .A1(G224), .A2(n612), .ZN(n358) );
  AND2_X1 U478 ( .A1(G210), .A2(n441), .ZN(n359) );
  XOR2_X1 U479 ( .A(n690), .B(n430), .Z(n360) );
  XOR2_X1 U480 ( .A(n693), .B(n692), .Z(n361) );
  NOR2_X1 U481 ( .A1(G952), .A2(n612), .ZN(n704) );
  INV_X1 U482 ( .A(n704), .ZN(n401) );
  XOR2_X1 U483 ( .A(n618), .B(KEYINPUT114), .Z(n362) );
  XOR2_X1 U484 ( .A(KEYINPUT56), .B(KEYINPUT122), .Z(n363) );
  XNOR2_X1 U485 ( .A(n364), .B(n408), .ZN(n407) );
  XNOR2_X2 U486 ( .A(n548), .B(n547), .ZN(n652) );
  NOR2_X1 U487 ( .A1(n414), .A2(n681), .ZN(n391) );
  XNOR2_X1 U488 ( .A(n576), .B(n577), .ZN(n372) );
  XNOR2_X1 U489 ( .A(n598), .B(KEYINPUT108), .ZN(n365) );
  NAND2_X1 U490 ( .A1(n404), .A2(n727), .ZN(n559) );
  NAND2_X1 U491 ( .A1(n366), .A2(n365), .ZN(n528) );
  NOR2_X1 U492 ( .A1(n695), .A2(n704), .ZN(n696) );
  NAND2_X1 U493 ( .A1(n523), .A2(n592), .ZN(n524) );
  XNOR2_X1 U494 ( .A(n375), .B(n374), .ZN(n525) );
  AND2_X1 U495 ( .A1(n553), .A2(n429), .ZN(n409) );
  NAND2_X1 U496 ( .A1(n368), .A2(n557), .ZN(n529) );
  INV_X1 U497 ( .A(n528), .ZN(n368) );
  XNOR2_X1 U498 ( .A(n391), .B(KEYINPUT85), .ZN(n390) );
  XNOR2_X1 U499 ( .A(n433), .B(n447), .ZN(n425) );
  NAND2_X1 U500 ( .A1(n372), .A2(n578), .ZN(n579) );
  NOR2_X1 U501 ( .A1(n544), .A2(n650), .ZN(n375) );
  NAND2_X1 U502 ( .A1(n585), .A2(n421), .ZN(n554) );
  NOR2_X2 U503 ( .A1(n564), .A2(n548), .ZN(n598) );
  NOR2_X1 U504 ( .A1(n608), .A2(n381), .ZN(n380) );
  INV_X1 U505 ( .A(n458), .ZN(n386) );
  INV_X1 U506 ( .A(n681), .ZN(n387) );
  NAND2_X1 U507 ( .A1(n415), .A2(n729), .ZN(n679) );
  NAND2_X1 U508 ( .A1(n390), .A2(n607), .ZN(n389) );
  NAND2_X1 U509 ( .A1(n582), .A2(n354), .ZN(n627) );
  XNOR2_X2 U510 ( .A(n395), .B(n394), .ZN(n681) );
  NAND2_X1 U511 ( .A1(n396), .A2(n605), .ZN(n395) );
  XNOR2_X1 U512 ( .A(n397), .B(n363), .ZN(G51) );
  NAND2_X1 U513 ( .A1(n398), .A2(n401), .ZN(n397) );
  XNOR2_X1 U514 ( .A(n399), .B(n360), .ZN(n398) );
  NAND2_X1 U515 ( .A1(n352), .A2(G210), .ZN(n399) );
  XNOR2_X1 U516 ( .A(n400), .B(n362), .ZN(G57) );
  NAND2_X1 U517 ( .A1(n402), .A2(n401), .ZN(n400) );
  XNOR2_X1 U518 ( .A(n403), .B(n351), .ZN(n402) );
  NAND2_X1 U519 ( .A1(n352), .A2(G472), .ZN(n403) );
  XNOR2_X1 U520 ( .A(n406), .B(n405), .ZN(n404) );
  INV_X1 U521 ( .A(KEYINPUT48), .ZN(n405) );
  NAND2_X1 U522 ( .A1(n409), .A2(n407), .ZN(n406) );
  NAND2_X1 U523 ( .A1(n415), .A2(n356), .ZN(n414) );
  OR2_X2 U524 ( .A1(n548), .A2(n525), .ZN(n540) );
  XNOR2_X2 U525 ( .A(G125), .B(G140), .ZN(n459) );
  NOR2_X2 U526 ( .A1(n561), .A2(n620), .ZN(n517) );
  XNOR2_X2 U527 ( .A(n517), .B(n518), .ZN(n728) );
  XNOR2_X2 U528 ( .A(n416), .B(n453), .ZN(n608) );
  XNOR2_X2 U529 ( .A(n514), .B(n417), .ZN(n717) );
  XNOR2_X1 U530 ( .A(n418), .B(n439), .ZN(n426) );
  XNOR2_X2 U531 ( .A(n432), .B(n431), .ZN(n418) );
  INV_X1 U532 ( .A(n717), .ZN(n420) );
  NOR2_X1 U533 ( .A1(n554), .A2(n545), .ZN(n546) );
  XNOR2_X2 U534 ( .A(n588), .B(KEYINPUT32), .ZN(n731) );
  XNOR2_X2 U535 ( .A(n575), .B(n428), .ZN(n597) );
  NOR2_X1 U536 ( .A1(n613), .A2(n704), .ZN(n615) );
  NOR2_X2 U537 ( .A1(G902), .A2(n702), .ZN(n479) );
  XNOR2_X1 U538 ( .A(n694), .B(n361), .ZN(n695) );
  XNOR2_X2 U539 ( .A(n460), .B(n459), .ZN(n502) );
  NOR2_X2 U540 ( .A1(n540), .A2(n574), .ZN(n633) );
  NOR2_X2 U541 ( .A1(n574), .A2(n573), .ZN(n575) );
  AND2_X1 U542 ( .A1(n645), .A2(n552), .ZN(n429) );
  XNOR2_X1 U543 ( .A(KEYINPUT54), .B(KEYINPUT55), .ZN(n430) );
  XNOR2_X1 U544 ( .A(n451), .B(G107), .ZN(n452) );
  INV_X1 U545 ( .A(KEYINPUT103), .ZN(n603) );
  XNOR2_X1 U546 ( .A(n452), .B(n461), .ZN(n453) );
  XNOR2_X1 U547 ( .A(n604), .B(n603), .ZN(n605) );
  XNOR2_X1 U548 ( .A(n455), .B(n454), .ZN(n456) );
  INV_X1 U549 ( .A(KEYINPUT79), .ZN(n462) );
  INV_X1 U550 ( .A(KEYINPUT19), .ZN(n538) );
  XNOR2_X1 U551 ( .A(n463), .B(n462), .ZN(n464) );
  XNOR2_X1 U552 ( .A(n608), .B(n609), .ZN(n610) );
  XNOR2_X1 U553 ( .A(KEYINPUT31), .B(KEYINPUT98), .ZN(n595) );
  INV_X1 U554 ( .A(KEYINPUT40), .ZN(n518) );
  XNOR2_X2 U555 ( .A(G128), .B(KEYINPUT64), .ZN(n432) );
  XNOR2_X1 U556 ( .A(n499), .B(n511), .ZN(n433) );
  XNOR2_X1 U557 ( .A(G119), .B(G101), .ZN(n434) );
  XNOR2_X1 U558 ( .A(n437), .B(n436), .ZN(n438) );
  NAND2_X1 U559 ( .A1(n690), .A2(n472), .ZN(n440) );
  BUF_X2 U560 ( .A(n537), .Z(n557) );
  INV_X1 U561 ( .A(n661), .ZN(n490) );
  NAND2_X1 U562 ( .A1(n441), .A2(G214), .ZN(n442) );
  XOR2_X1 U563 ( .A(KEYINPUT91), .B(n442), .Z(n660) );
  XOR2_X1 U564 ( .A(G113), .B(KEYINPUT5), .Z(n445) );
  XNOR2_X1 U565 ( .A(n445), .B(n444), .ZN(n446) );
  NAND2_X1 U566 ( .A1(n660), .A2(n600), .ZN(n449) );
  XNOR2_X1 U567 ( .A(n449), .B(KEYINPUT30), .ZN(n484) );
  XOR2_X1 U568 ( .A(n450), .B(G140), .Z(n451) );
  NAND2_X1 U569 ( .A1(G227), .A2(n612), .ZN(n454) );
  XOR2_X1 U570 ( .A(G469), .B(KEYINPUT71), .Z(n457) );
  XNOR2_X1 U571 ( .A(KEYINPUT72), .B(n457), .ZN(n458) );
  NAND2_X1 U572 ( .A1(G234), .A2(n612), .ZN(n465) );
  XOR2_X1 U573 ( .A(KEYINPUT8), .B(n465), .Z(n507) );
  AND2_X1 U574 ( .A1(G221), .A2(n507), .ZN(n469) );
  XOR2_X1 U575 ( .A(KEYINPUT24), .B(KEYINPUT23), .Z(n467) );
  XNOR2_X1 U576 ( .A(n467), .B(n466), .ZN(n468) );
  NAND2_X1 U577 ( .A1(n472), .A2(G234), .ZN(n473) );
  XNOR2_X1 U578 ( .A(n473), .B(KEYINPUT20), .ZN(n480) );
  NAND2_X1 U579 ( .A1(G217), .A2(n480), .ZN(n477) );
  XNOR2_X1 U580 ( .A(KEYINPUT25), .B(KEYINPUT78), .ZN(n474) );
  XNOR2_X1 U581 ( .A(n475), .B(n474), .ZN(n476) );
  XOR2_X1 U582 ( .A(KEYINPUT96), .B(KEYINPUT21), .Z(n482) );
  NAND2_X1 U583 ( .A1(n480), .A2(G221), .ZN(n481) );
  NAND2_X1 U584 ( .A1(n646), .A2(n647), .ZN(n483) );
  XNOR2_X1 U585 ( .A(n485), .B(KEYINPUT14), .ZN(n487) );
  NAND2_X1 U586 ( .A1(G952), .A2(n487), .ZN(n674) );
  NOR2_X1 U587 ( .A1(G953), .A2(n674), .ZN(n486) );
  XOR2_X1 U588 ( .A(KEYINPUT92), .B(n486), .Z(n569) );
  NAND2_X1 U589 ( .A1(G902), .A2(n487), .ZN(n570) );
  NOR2_X1 U590 ( .A1(G900), .A2(n570), .ZN(n488) );
  NAND2_X1 U591 ( .A1(G953), .A2(n488), .ZN(n489) );
  NAND2_X1 U592 ( .A1(n569), .A2(n489), .ZN(n521) );
  XNOR2_X1 U593 ( .A(KEYINPUT74), .B(KEYINPUT39), .ZN(n491) );
  XNOR2_X1 U594 ( .A(KEYINPUT13), .B(G475), .ZN(n506) );
  XOR2_X1 U595 ( .A(KEYINPUT100), .B(KEYINPUT11), .Z(n494) );
  NAND2_X1 U596 ( .A1(G214), .A2(n492), .ZN(n493) );
  XNOR2_X1 U597 ( .A(n494), .B(n493), .ZN(n498) );
  XOR2_X1 U598 ( .A(KEYINPUT12), .B(KEYINPUT99), .Z(n496) );
  XNOR2_X1 U599 ( .A(n496), .B(n495), .ZN(n497) );
  XOR2_X1 U600 ( .A(n498), .B(n497), .Z(n504) );
  XNOR2_X1 U601 ( .A(G143), .B(G131), .ZN(n500) );
  XNOR2_X1 U602 ( .A(n500), .B(n499), .ZN(n501) );
  XNOR2_X1 U603 ( .A(n502), .B(n501), .ZN(n503) );
  XNOR2_X1 U604 ( .A(n504), .B(n503), .ZN(n691) );
  NOR2_X1 U605 ( .A1(G902), .A2(n691), .ZN(n505) );
  XNOR2_X1 U606 ( .A(n506), .B(n505), .ZN(n534) );
  NAND2_X1 U607 ( .A1(G217), .A2(n507), .ZN(n508) );
  XNOR2_X1 U608 ( .A(n509), .B(n508), .ZN(n510) );
  XOR2_X1 U609 ( .A(n510), .B(KEYINPUT101), .Z(n513) );
  XNOR2_X1 U610 ( .A(n511), .B(G116), .ZN(n512) );
  INV_X1 U611 ( .A(n514), .ZN(n515) );
  NOR2_X1 U612 ( .A1(n698), .A2(G902), .ZN(n516) );
  XNOR2_X1 U613 ( .A(n516), .B(G478), .ZN(n533) );
  NAND2_X1 U614 ( .A1(n534), .A2(n533), .ZN(n620) );
  INV_X1 U615 ( .A(n534), .ZN(n530) );
  NAND2_X1 U616 ( .A1(n530), .A2(n533), .ZN(n663) );
  NOR2_X1 U617 ( .A1(n663), .A2(n664), .ZN(n520) );
  XNOR2_X1 U618 ( .A(KEYINPUT110), .B(KEYINPUT41), .ZN(n519) );
  XNOR2_X1 U619 ( .A(n520), .B(n519), .ZN(n676) );
  INV_X1 U620 ( .A(n353), .ZN(n592) );
  NAND2_X1 U621 ( .A1(n647), .A2(n521), .ZN(n522) );
  XOR2_X1 U622 ( .A(KEYINPUT70), .B(n522), .Z(n523) );
  XNOR2_X1 U623 ( .A(KEYINPUT111), .B(KEYINPUT42), .ZN(n526) );
  XNOR2_X1 U624 ( .A(n529), .B(KEYINPUT109), .ZN(n532) );
  OR2_X1 U625 ( .A1(n530), .A2(n533), .ZN(n531) );
  XOR2_X1 U626 ( .A(KEYINPUT106), .B(n531), .Z(n563) );
  NAND2_X1 U627 ( .A1(n532), .A2(n563), .ZN(n632) );
  NOR2_X1 U628 ( .A1(n534), .A2(n533), .ZN(n640) );
  XOR2_X1 U629 ( .A(KEYINPUT102), .B(n640), .Z(n560) );
  AND2_X1 U630 ( .A1(n620), .A2(n560), .ZN(n665) );
  NAND2_X1 U631 ( .A1(KEYINPUT47), .A2(n665), .ZN(n535) );
  NAND2_X1 U632 ( .A1(n632), .A2(n535), .ZN(n536) );
  XNOR2_X1 U633 ( .A(n536), .B(KEYINPUT83), .ZN(n543) );
  NAND2_X1 U634 ( .A1(n537), .A2(n660), .ZN(n539) );
  NOR2_X1 U635 ( .A1(KEYINPUT47), .A2(n665), .ZN(n541) );
  NAND2_X1 U636 ( .A1(n633), .A2(n541), .ZN(n542) );
  AND2_X1 U637 ( .A1(n543), .A2(n542), .ZN(n553) );
  INV_X1 U638 ( .A(n557), .ZN(n545) );
  XOR2_X1 U639 ( .A(KEYINPUT6), .B(n650), .Z(n589) );
  XNOR2_X1 U640 ( .A(KEYINPUT36), .B(n546), .ZN(n550) );
  INV_X1 U641 ( .A(KEYINPUT1), .ZN(n547) );
  XNOR2_X1 U642 ( .A(KEYINPUT89), .B(n371), .ZN(n583) );
  INV_X1 U643 ( .A(n583), .ZN(n549) );
  NAND2_X1 U644 ( .A1(n550), .A2(n549), .ZN(n645) );
  INV_X1 U645 ( .A(n633), .ZN(n551) );
  NAND2_X1 U646 ( .A1(KEYINPUT47), .A2(n551), .ZN(n552) );
  NOR2_X1 U647 ( .A1(n371), .A2(n554), .ZN(n555) );
  XNOR2_X1 U648 ( .A(n555), .B(KEYINPUT43), .ZN(n556) );
  NOR2_X1 U649 ( .A1(n557), .A2(n556), .ZN(n558) );
  XNOR2_X1 U650 ( .A(KEYINPUT107), .B(n558), .ZN(n727) );
  NOR2_X1 U651 ( .A1(n561), .A2(n560), .ZN(n562) );
  XOR2_X1 U652 ( .A(KEYINPUT112), .B(n562), .Z(n729) );
  XOR2_X1 U653 ( .A(n563), .B(KEYINPUT81), .Z(n578) );
  XOR2_X1 U654 ( .A(KEYINPUT34), .B(KEYINPUT82), .Z(n577) );
  INV_X1 U655 ( .A(n564), .ZN(n651) );
  INV_X1 U656 ( .A(n589), .ZN(n585) );
  NAND2_X1 U657 ( .A1(n593), .A2(n585), .ZN(n568) );
  XNOR2_X1 U658 ( .A(KEYINPUT105), .B(KEYINPUT33), .ZN(n566) );
  XNOR2_X1 U659 ( .A(n566), .B(KEYINPUT73), .ZN(n567) );
  XNOR2_X1 U660 ( .A(n568), .B(n567), .ZN(n668) );
  INV_X1 U661 ( .A(n569), .ZN(n572) );
  XNOR2_X1 U662 ( .A(G898), .B(KEYINPUT93), .ZN(n711) );
  NAND2_X1 U663 ( .A1(G953), .A2(n711), .ZN(n706) );
  NOR2_X1 U664 ( .A1(n570), .A2(n706), .ZN(n571) );
  NOR2_X1 U665 ( .A1(n572), .A2(n571), .ZN(n573) );
  NAND2_X1 U666 ( .A1(n668), .A2(n597), .ZN(n576) );
  INV_X1 U667 ( .A(n647), .ZN(n580) );
  NOR2_X1 U668 ( .A1(n580), .A2(n663), .ZN(n581) );
  XNOR2_X1 U669 ( .A(n590), .B(KEYINPUT104), .ZN(n582) );
  NOR2_X1 U670 ( .A1(n584), .A2(n583), .ZN(n587) );
  NOR2_X1 U671 ( .A1(n379), .A2(n585), .ZN(n586) );
  NAND2_X1 U672 ( .A1(n587), .A2(n586), .ZN(n588) );
  NAND2_X1 U673 ( .A1(n590), .A2(n589), .ZN(n591) );
  NOR2_X1 U674 ( .A1(n592), .A2(n591), .ZN(n619) );
  NAND2_X1 U675 ( .A1(n593), .A2(n600), .ZN(n594) );
  NAND2_X1 U676 ( .A1(n657), .A2(n597), .ZN(n596) );
  NAND2_X1 U677 ( .A1(n598), .A2(n597), .ZN(n599) );
  NOR2_X1 U678 ( .A1(n600), .A2(n599), .ZN(n623) );
  NOR2_X1 U679 ( .A1(n639), .A2(n623), .ZN(n601) );
  NOR2_X1 U680 ( .A1(n665), .A2(n601), .ZN(n602) );
  NOR2_X1 U681 ( .A1(n619), .A2(n602), .ZN(n604) );
  NAND2_X1 U682 ( .A1(KEYINPUT2), .A2(n606), .ZN(n607) );
  NAND2_X1 U683 ( .A1(n700), .A2(G469), .ZN(n611) );
  XOR2_X1 U684 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n609) );
  XNOR2_X1 U685 ( .A(n611), .B(n610), .ZN(n613) );
  INV_X1 U686 ( .A(KEYINPUT123), .ZN(n614) );
  XNOR2_X1 U687 ( .A(n615), .B(n614), .ZN(G54) );
  XOR2_X1 U688 ( .A(KEYINPUT62), .B(KEYINPUT113), .Z(n616) );
  INV_X1 U689 ( .A(KEYINPUT63), .ZN(n618) );
  XOR2_X1 U690 ( .A(G101), .B(n619), .Z(G3) );
  XOR2_X1 U691 ( .A(G104), .B(KEYINPUT115), .Z(n622) );
  INV_X1 U692 ( .A(n620), .ZN(n636) );
  NAND2_X1 U693 ( .A1(n623), .A2(n636), .ZN(n621) );
  XNOR2_X1 U694 ( .A(n622), .B(n621), .ZN(G6) );
  XOR2_X1 U695 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n625) );
  NAND2_X1 U696 ( .A1(n623), .A2(n640), .ZN(n624) );
  XNOR2_X1 U697 ( .A(n625), .B(n624), .ZN(n626) );
  XNOR2_X1 U698 ( .A(G107), .B(n626), .ZN(G9) );
  XNOR2_X1 U699 ( .A(n627), .B(G110), .ZN(G12) );
  XOR2_X1 U700 ( .A(KEYINPUT116), .B(KEYINPUT29), .Z(n629) );
  NAND2_X1 U701 ( .A1(n633), .A2(n640), .ZN(n628) );
  XNOR2_X1 U702 ( .A(n629), .B(n628), .ZN(n630) );
  XNOR2_X1 U703 ( .A(G128), .B(n630), .ZN(G30) );
  XOR2_X1 U704 ( .A(G143), .B(KEYINPUT117), .Z(n631) );
  XNOR2_X1 U705 ( .A(n632), .B(n631), .ZN(G45) );
  NAND2_X1 U706 ( .A1(n633), .A2(n636), .ZN(n634) );
  XNOR2_X1 U707 ( .A(n634), .B(KEYINPUT118), .ZN(n635) );
  XNOR2_X1 U708 ( .A(G146), .B(n635), .ZN(G48) );
  XOR2_X1 U709 ( .A(G113), .B(KEYINPUT119), .Z(n638) );
  NAND2_X1 U710 ( .A1(n636), .A2(n639), .ZN(n637) );
  XNOR2_X1 U711 ( .A(n638), .B(n637), .ZN(G15) );
  XOR2_X1 U712 ( .A(KEYINPUT120), .B(KEYINPUT121), .Z(n642) );
  NAND2_X1 U713 ( .A1(n640), .A2(n639), .ZN(n641) );
  XNOR2_X1 U714 ( .A(n642), .B(n641), .ZN(n643) );
  XNOR2_X1 U715 ( .A(G116), .B(n643), .ZN(G18) );
  XOR2_X1 U716 ( .A(G125), .B(KEYINPUT37), .Z(n644) );
  XNOR2_X1 U717 ( .A(n645), .B(n644), .ZN(G27) );
  NOR2_X1 U718 ( .A1(n647), .A2(n379), .ZN(n648) );
  XNOR2_X1 U719 ( .A(n648), .B(KEYINPUT49), .ZN(n649) );
  NAND2_X1 U720 ( .A1(n650), .A2(n649), .ZN(n655) );
  NOR2_X1 U721 ( .A1(n371), .A2(n651), .ZN(n653) );
  XNOR2_X1 U722 ( .A(n653), .B(KEYINPUT50), .ZN(n654) );
  NOR2_X1 U723 ( .A1(n655), .A2(n654), .ZN(n656) );
  NOR2_X1 U724 ( .A1(n657), .A2(n656), .ZN(n658) );
  XOR2_X1 U725 ( .A(KEYINPUT51), .B(n658), .Z(n659) );
  NOR2_X1 U726 ( .A1(n676), .A2(n659), .ZN(n671) );
  NOR2_X1 U727 ( .A1(n661), .A2(n660), .ZN(n662) );
  NOR2_X1 U728 ( .A1(n663), .A2(n662), .ZN(n667) );
  NOR2_X1 U729 ( .A1(n665), .A2(n664), .ZN(n666) );
  NOR2_X1 U730 ( .A1(n667), .A2(n666), .ZN(n669) );
  INV_X1 U731 ( .A(n668), .ZN(n675) );
  NOR2_X1 U732 ( .A1(n669), .A2(n675), .ZN(n670) );
  NOR2_X1 U733 ( .A1(n671), .A2(n670), .ZN(n672) );
  XNOR2_X1 U734 ( .A(n672), .B(KEYINPUT52), .ZN(n673) );
  NOR2_X1 U735 ( .A1(n674), .A2(n673), .ZN(n678) );
  NOR2_X1 U736 ( .A1(n676), .A2(n675), .ZN(n677) );
  NOR2_X1 U737 ( .A1(n678), .A2(n677), .ZN(n688) );
  INV_X1 U738 ( .A(KEYINPUT2), .ZN(n682) );
  NAND2_X1 U739 ( .A1(n679), .A2(n682), .ZN(n680) );
  XNOR2_X1 U740 ( .A(n680), .B(KEYINPUT84), .ZN(n684) );
  NAND2_X1 U741 ( .A1(n681), .A2(n682), .ZN(n683) );
  NAND2_X1 U742 ( .A1(n684), .A2(n683), .ZN(n687) );
  INV_X1 U743 ( .A(n685), .ZN(n686) );
  XNOR2_X1 U744 ( .A(n689), .B(KEYINPUT53), .ZN(G75) );
  XOR2_X1 U745 ( .A(KEYINPUT65), .B(KEYINPUT59), .Z(n693) );
  XNOR2_X1 U746 ( .A(n691), .B(KEYINPUT90), .ZN(n692) );
  XNOR2_X1 U747 ( .A(KEYINPUT60), .B(n696), .ZN(G60) );
  NAND2_X1 U748 ( .A1(G478), .A2(n352), .ZN(n697) );
  XNOR2_X1 U749 ( .A(n698), .B(n697), .ZN(n699) );
  NOR2_X1 U750 ( .A1(n704), .A2(n699), .ZN(G63) );
  NAND2_X1 U751 ( .A1(G217), .A2(n352), .ZN(n701) );
  XNOR2_X1 U752 ( .A(n702), .B(n701), .ZN(n703) );
  NOR2_X1 U753 ( .A1(n704), .A2(n703), .ZN(G66) );
  NAND2_X1 U754 ( .A1(n706), .A2(n705), .ZN(n715) );
  XOR2_X1 U755 ( .A(KEYINPUT61), .B(KEYINPUT125), .Z(n708) );
  NAND2_X1 U756 ( .A1(G224), .A2(G953), .ZN(n707) );
  XNOR2_X1 U757 ( .A(n708), .B(n707), .ZN(n709) );
  XOR2_X1 U758 ( .A(KEYINPUT124), .B(n709), .Z(n710) );
  NOR2_X1 U759 ( .A1(n711), .A2(n710), .ZN(n713) );
  NOR2_X1 U760 ( .A1(G953), .A2(n681), .ZN(n712) );
  NOR2_X1 U761 ( .A1(n713), .A2(n712), .ZN(n714) );
  XNOR2_X1 U762 ( .A(n715), .B(n714), .ZN(G69) );
  XOR2_X1 U763 ( .A(n717), .B(n716), .Z(n719) );
  XOR2_X1 U764 ( .A(n719), .B(n679), .Z(n718) );
  NOR2_X1 U765 ( .A1(G953), .A2(n718), .ZN(n724) );
  XNOR2_X1 U766 ( .A(G227), .B(n719), .ZN(n720) );
  NAND2_X1 U767 ( .A1(n720), .A2(G900), .ZN(n721) );
  NAND2_X1 U768 ( .A1(n721), .A2(G953), .ZN(n722) );
  XOR2_X1 U769 ( .A(KEYINPUT126), .B(n722), .Z(n723) );
  NOR2_X1 U770 ( .A1(n724), .A2(n723), .ZN(n725) );
  XNOR2_X1 U771 ( .A(KEYINPUT127), .B(n725), .ZN(G72) );
  XOR2_X1 U772 ( .A(n726), .B(G122), .Z(G24) );
  XNOR2_X1 U773 ( .A(G140), .B(n727), .ZN(G42) );
  XNOR2_X1 U774 ( .A(n728), .B(G131), .ZN(G33) );
  XNOR2_X1 U775 ( .A(G134), .B(n729), .ZN(G36) );
  XNOR2_X1 U776 ( .A(n730), .B(G137), .ZN(G39) );
  XNOR2_X1 U777 ( .A(n731), .B(G119), .ZN(G21) );
endmodule

