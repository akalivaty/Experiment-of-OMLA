//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 0 1 1 1 1 1 0 1 1 1 0 0 1 0 1 0 0 1 0 1 0 1 0 0 0 0 0 1 0 0 0 1 1 0 1 1 0 1 0 1 0 0 1 1 1 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:17:09 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n658,
    new_n659, new_n660, new_n662, new_n663, new_n664, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n684, new_n685, new_n686, new_n687, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n717, new_n718, new_n719, new_n720,
    new_n722, new_n723, new_n724, new_n725, new_n726, new_n727, new_n729,
    new_n730, new_n731, new_n733, new_n734, new_n736, new_n737, new_n738,
    new_n739, new_n740, new_n741, new_n742, new_n743, new_n744, new_n745,
    new_n746, new_n747, new_n748, new_n749, new_n750, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n764, new_n765, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n819, new_n820,
    new_n821, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n830, new_n831, new_n832, new_n833, new_n834, new_n835, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n875,
    new_n876, new_n877, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n886, new_n887, new_n889, new_n890, new_n891, new_n892,
    new_n893, new_n894, new_n895, new_n896, new_n897, new_n898, new_n899,
    new_n900, new_n901, new_n902, new_n904, new_n905, new_n906, new_n907,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n924,
    new_n925, new_n926, new_n927, new_n928, new_n929, new_n931, new_n932;
  XNOR2_X1  g000(.A(G113gat), .B(G141gat), .ZN(new_n202));
  XNOR2_X1  g001(.A(KEYINPUT87), .B(KEYINPUT11), .ZN(new_n203));
  XNOR2_X1  g002(.A(new_n202), .B(new_n203), .ZN(new_n204));
  XOR2_X1   g003(.A(G169gat), .B(G197gat), .Z(new_n205));
  XNOR2_X1  g004(.A(new_n204), .B(new_n205), .ZN(new_n206));
  XNOR2_X1  g005(.A(new_n206), .B(KEYINPUT12), .ZN(new_n207));
  INV_X1    g006(.A(new_n207), .ZN(new_n208));
  XNOR2_X1  g007(.A(G15gat), .B(G22gat), .ZN(new_n209));
  INV_X1    g008(.A(KEYINPUT88), .ZN(new_n210));
  NAND2_X1  g009(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  INV_X1    g010(.A(G8gat), .ZN(new_n212));
  XNOR2_X1  g011(.A(new_n211), .B(new_n212), .ZN(new_n213));
  INV_X1    g012(.A(KEYINPUT16), .ZN(new_n214));
  AOI21_X1  g013(.A(G1gat), .B1(new_n209), .B2(new_n214), .ZN(new_n215));
  XNOR2_X1  g014(.A(new_n213), .B(new_n215), .ZN(new_n216));
  OR2_X1    g015(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n217));
  NAND2_X1  g016(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n218));
  AOI21_X1  g017(.A(G36gat), .B1(new_n217), .B2(new_n218), .ZN(new_n219));
  INV_X1    g018(.A(G29gat), .ZN(new_n220));
  AND3_X1   g019(.A1(new_n220), .A2(KEYINPUT14), .A3(G36gat), .ZN(new_n221));
  OR3_X1    g020(.A1(new_n219), .A2(KEYINPUT15), .A3(new_n221), .ZN(new_n222));
  OAI21_X1  g021(.A(KEYINPUT15), .B1(new_n219), .B2(new_n221), .ZN(new_n223));
  XNOR2_X1  g022(.A(G43gat), .B(G50gat), .ZN(new_n224));
  NAND3_X1  g023(.A1(new_n222), .A2(new_n223), .A3(new_n224), .ZN(new_n225));
  OR2_X1    g024(.A1(new_n223), .A2(new_n224), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  NOR2_X1   g026(.A1(new_n227), .A2(KEYINPUT17), .ZN(new_n228));
  INV_X1    g027(.A(KEYINPUT17), .ZN(new_n229));
  AOI21_X1  g028(.A(new_n229), .B1(new_n225), .B2(new_n226), .ZN(new_n230));
  OAI21_X1  g029(.A(new_n216), .B1(new_n228), .B2(new_n230), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n231), .A2(KEYINPUT89), .ZN(new_n232));
  AND2_X1   g031(.A1(new_n213), .A2(new_n215), .ZN(new_n233));
  NOR2_X1   g032(.A1(new_n213), .A2(new_n215), .ZN(new_n234));
  NOR2_X1   g033(.A1(new_n233), .A2(new_n234), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n235), .A2(new_n227), .ZN(new_n236));
  INV_X1    g035(.A(KEYINPUT89), .ZN(new_n237));
  OAI211_X1 g036(.A(new_n237), .B(new_n216), .C1(new_n228), .C2(new_n230), .ZN(new_n238));
  AND3_X1   g037(.A1(new_n232), .A2(new_n236), .A3(new_n238), .ZN(new_n239));
  INV_X1    g038(.A(KEYINPUT92), .ZN(new_n240));
  NAND2_X1  g039(.A1(G229gat), .A2(G233gat), .ZN(new_n241));
  NAND4_X1  g040(.A1(new_n239), .A2(new_n240), .A3(KEYINPUT18), .A4(new_n241), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n236), .A2(KEYINPUT93), .ZN(new_n243));
  INV_X1    g042(.A(new_n227), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n216), .A2(new_n244), .ZN(new_n245));
  XNOR2_X1  g044(.A(new_n243), .B(new_n245), .ZN(new_n246));
  XOR2_X1   g045(.A(new_n241), .B(KEYINPUT13), .Z(new_n247));
  NAND2_X1  g046(.A1(new_n246), .A2(new_n247), .ZN(new_n248));
  NAND4_X1  g047(.A1(new_n232), .A2(new_n241), .A3(new_n236), .A4(new_n238), .ZN(new_n249));
  INV_X1    g048(.A(KEYINPUT18), .ZN(new_n250));
  OAI21_X1  g049(.A(KEYINPUT92), .B1(new_n249), .B2(new_n250), .ZN(new_n251));
  NAND3_X1  g050(.A1(new_n242), .A2(new_n248), .A3(new_n251), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n249), .A2(KEYINPUT90), .ZN(new_n253));
  AND2_X1   g052(.A1(new_n238), .A2(new_n236), .ZN(new_n254));
  INV_X1    g053(.A(KEYINPUT90), .ZN(new_n255));
  NAND4_X1  g054(.A1(new_n254), .A2(new_n255), .A3(new_n241), .A4(new_n232), .ZN(new_n256));
  XNOR2_X1  g055(.A(KEYINPUT91), .B(KEYINPUT18), .ZN(new_n257));
  AND3_X1   g056(.A1(new_n253), .A2(new_n256), .A3(new_n257), .ZN(new_n258));
  OAI21_X1  g057(.A(new_n208), .B1(new_n252), .B2(new_n258), .ZN(new_n259));
  NAND4_X1  g058(.A1(new_n254), .A2(KEYINPUT18), .A3(new_n241), .A4(new_n232), .ZN(new_n260));
  AOI22_X1  g059(.A1(new_n260), .A2(KEYINPUT92), .B1(new_n246), .B2(new_n247), .ZN(new_n261));
  NAND3_X1  g060(.A1(new_n253), .A2(new_n256), .A3(new_n257), .ZN(new_n262));
  NAND4_X1  g061(.A1(new_n261), .A2(new_n262), .A3(new_n242), .A4(new_n207), .ZN(new_n263));
  NAND2_X1  g062(.A1(new_n259), .A2(new_n263), .ZN(new_n264));
  INV_X1    g063(.A(new_n264), .ZN(new_n265));
  INV_X1    g064(.A(KEYINPUT36), .ZN(new_n266));
  XOR2_X1   g065(.A(KEYINPUT67), .B(G190gat), .Z(new_n267));
  XNOR2_X1  g066(.A(KEYINPUT27), .B(G183gat), .ZN(new_n268));
  NAND3_X1  g067(.A1(new_n267), .A2(KEYINPUT28), .A3(new_n268), .ZN(new_n269));
  INV_X1    g068(.A(KEYINPUT69), .ZN(new_n270));
  INV_X1    g069(.A(G183gat), .ZN(new_n271));
  OAI21_X1  g070(.A(new_n270), .B1(new_n271), .B2(KEYINPUT27), .ZN(new_n272));
  OAI211_X1 g071(.A(new_n267), .B(new_n272), .C1(new_n270), .C2(new_n268), .ZN(new_n273));
  INV_X1    g072(.A(KEYINPUT70), .ZN(new_n274));
  AND2_X1   g073(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  INV_X1    g074(.A(KEYINPUT28), .ZN(new_n276));
  OAI21_X1  g075(.A(new_n276), .B1(new_n273), .B2(new_n274), .ZN(new_n277));
  OAI21_X1  g076(.A(new_n269), .B1(new_n275), .B2(new_n277), .ZN(new_n278));
  NOR2_X1   g077(.A1(G169gat), .A2(G176gat), .ZN(new_n279));
  AOI22_X1  g078(.A1(new_n279), .A2(KEYINPUT26), .B1(G183gat), .B2(G190gat), .ZN(new_n280));
  OR2_X1    g079(.A1(new_n279), .A2(KEYINPUT26), .ZN(new_n281));
  INV_X1    g080(.A(G169gat), .ZN(new_n282));
  INV_X1    g081(.A(G176gat), .ZN(new_n283));
  NOR2_X1   g082(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  OAI21_X1  g083(.A(new_n280), .B1(new_n281), .B2(new_n284), .ZN(new_n285));
  XOR2_X1   g084(.A(new_n285), .B(KEYINPUT71), .Z(new_n286));
  NAND2_X1  g085(.A1(new_n278), .A2(new_n286), .ZN(new_n287));
  INV_X1    g086(.A(new_n287), .ZN(new_n288));
  INV_X1    g087(.A(KEYINPUT25), .ZN(new_n289));
  NAND3_X1  g088(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n290));
  AOI21_X1  g089(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n291));
  OAI221_X1 g090(.A(new_n290), .B1(G183gat), .B2(G190gat), .C1(new_n291), .C2(KEYINPUT64), .ZN(new_n292));
  AOI21_X1  g091(.A(new_n292), .B1(KEYINPUT64), .B2(new_n291), .ZN(new_n293));
  XOR2_X1   g092(.A(KEYINPUT65), .B(G169gat), .Z(new_n294));
  INV_X1    g093(.A(KEYINPUT23), .ZN(new_n295));
  NOR2_X1   g094(.A1(new_n295), .A2(G176gat), .ZN(new_n296));
  NAND2_X1  g095(.A1(new_n294), .A2(new_n296), .ZN(new_n297));
  INV_X1    g096(.A(new_n279), .ZN(new_n298));
  OAI21_X1  g097(.A(new_n298), .B1(new_n284), .B2(new_n295), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n297), .A2(new_n299), .ZN(new_n300));
  OAI21_X1  g099(.A(new_n289), .B1(new_n293), .B2(new_n300), .ZN(new_n301));
  INV_X1    g100(.A(KEYINPUT66), .ZN(new_n302));
  XNOR2_X1  g101(.A(new_n301), .B(new_n302), .ZN(new_n303));
  AOI21_X1  g102(.A(new_n289), .B1(new_n296), .B2(new_n282), .ZN(new_n304));
  INV_X1    g103(.A(new_n267), .ZN(new_n305));
  NOR2_X1   g104(.A1(new_n305), .A2(G183gat), .ZN(new_n306));
  INV_X1    g105(.A(new_n291), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n307), .A2(new_n290), .ZN(new_n308));
  OAI211_X1 g107(.A(new_n299), .B(new_n304), .C1(new_n306), .C2(new_n308), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n303), .A2(new_n309), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n310), .A2(KEYINPUT68), .ZN(new_n311));
  INV_X1    g110(.A(KEYINPUT68), .ZN(new_n312));
  NAND3_X1  g111(.A1(new_n303), .A2(new_n312), .A3(new_n309), .ZN(new_n313));
  AOI21_X1  g112(.A(new_n288), .B1(new_n311), .B2(new_n313), .ZN(new_n314));
  XNOR2_X1  g113(.A(G113gat), .B(G120gat), .ZN(new_n315));
  INV_X1    g114(.A(KEYINPUT72), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n315), .A2(new_n316), .ZN(new_n317));
  INV_X1    g116(.A(KEYINPUT1), .ZN(new_n318));
  INV_X1    g117(.A(G120gat), .ZN(new_n319));
  OR3_X1    g118(.A1(new_n316), .A2(new_n319), .A3(G113gat), .ZN(new_n320));
  XNOR2_X1  g119(.A(G127gat), .B(G134gat), .ZN(new_n321));
  NAND4_X1  g120(.A1(new_n317), .A2(new_n318), .A3(new_n320), .A4(new_n321), .ZN(new_n322));
  XNOR2_X1  g121(.A(new_n322), .B(KEYINPUT73), .ZN(new_n323));
  INV_X1    g122(.A(new_n321), .ZN(new_n324));
  OAI21_X1  g123(.A(new_n324), .B1(new_n315), .B2(KEYINPUT1), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n323), .A2(new_n325), .ZN(new_n326));
  NOR2_X1   g125(.A1(new_n314), .A2(new_n326), .ZN(new_n327));
  AND2_X1   g126(.A1(new_n323), .A2(new_n325), .ZN(new_n328));
  AOI211_X1 g127(.A(new_n328), .B(new_n288), .C1(new_n311), .C2(new_n313), .ZN(new_n329));
  NOR2_X1   g128(.A1(new_n327), .A2(new_n329), .ZN(new_n330));
  INV_X1    g129(.A(G227gat), .ZN(new_n331));
  INV_X1    g130(.A(G233gat), .ZN(new_n332));
  NOR2_X1   g131(.A1(new_n331), .A2(new_n332), .ZN(new_n333));
  OAI21_X1  g132(.A(KEYINPUT34), .B1(new_n330), .B2(new_n333), .ZN(new_n334));
  NAND2_X1  g133(.A1(new_n311), .A2(new_n313), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n335), .A2(new_n287), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n336), .A2(new_n328), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n314), .A2(new_n326), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n337), .A2(new_n338), .ZN(new_n339));
  INV_X1    g138(.A(KEYINPUT34), .ZN(new_n340));
  INV_X1    g139(.A(new_n333), .ZN(new_n341));
  NAND3_X1  g140(.A1(new_n339), .A2(new_n340), .A3(new_n341), .ZN(new_n342));
  AOI21_X1  g141(.A(KEYINPUT33), .B1(new_n330), .B2(new_n333), .ZN(new_n343));
  XNOR2_X1  g142(.A(G15gat), .B(G43gat), .ZN(new_n344));
  XNOR2_X1  g143(.A(new_n344), .B(KEYINPUT74), .ZN(new_n345));
  XNOR2_X1  g144(.A(G71gat), .B(G99gat), .ZN(new_n346));
  XNOR2_X1  g145(.A(new_n346), .B(KEYINPUT75), .ZN(new_n347));
  XNOR2_X1  g146(.A(new_n345), .B(new_n347), .ZN(new_n348));
  OAI211_X1 g147(.A(new_n334), .B(new_n342), .C1(new_n343), .C2(new_n348), .ZN(new_n349));
  NAND3_X1  g148(.A1(new_n337), .A2(new_n333), .A3(new_n338), .ZN(new_n350));
  INV_X1    g149(.A(KEYINPUT33), .ZN(new_n351));
  AOI21_X1  g150(.A(new_n348), .B1(new_n350), .B2(new_n351), .ZN(new_n352));
  AOI21_X1  g151(.A(new_n340), .B1(new_n339), .B2(new_n341), .ZN(new_n353));
  AOI211_X1 g152(.A(KEYINPUT34), .B(new_n333), .C1(new_n337), .C2(new_n338), .ZN(new_n354));
  OAI21_X1  g153(.A(new_n352), .B1(new_n353), .B2(new_n354), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n350), .A2(KEYINPUT32), .ZN(new_n356));
  INV_X1    g155(.A(new_n356), .ZN(new_n357));
  AND3_X1   g156(.A1(new_n349), .A2(new_n355), .A3(new_n357), .ZN(new_n358));
  AOI21_X1  g157(.A(new_n357), .B1(new_n349), .B2(new_n355), .ZN(new_n359));
  OAI21_X1  g158(.A(new_n266), .B1(new_n358), .B2(new_n359), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n349), .A2(new_n355), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n361), .A2(new_n356), .ZN(new_n362));
  NAND3_X1  g161(.A1(new_n349), .A2(new_n355), .A3(new_n357), .ZN(new_n363));
  NAND3_X1  g162(.A1(new_n362), .A2(KEYINPUT36), .A3(new_n363), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n360), .A2(new_n364), .ZN(new_n365));
  XOR2_X1   g164(.A(G141gat), .B(G148gat), .Z(new_n366));
  INV_X1    g165(.A(G155gat), .ZN(new_n367));
  INV_X1    g166(.A(G162gat), .ZN(new_n368));
  OAI21_X1  g167(.A(KEYINPUT2), .B1(new_n367), .B2(new_n368), .ZN(new_n369));
  NAND3_X1  g168(.A1(new_n366), .A2(KEYINPUT78), .A3(new_n369), .ZN(new_n370));
  XNOR2_X1  g169(.A(G155gat), .B(G162gat), .ZN(new_n371));
  XNOR2_X1  g170(.A(new_n370), .B(new_n371), .ZN(new_n372));
  INV_X1    g171(.A(new_n372), .ZN(new_n373));
  OAI21_X1  g172(.A(KEYINPUT4), .B1(new_n326), .B2(new_n373), .ZN(new_n374));
  INV_X1    g173(.A(KEYINPUT4), .ZN(new_n375));
  NAND3_X1  g174(.A1(new_n328), .A2(new_n375), .A3(new_n372), .ZN(new_n376));
  INV_X1    g175(.A(KEYINPUT81), .ZN(new_n377));
  AND3_X1   g176(.A1(new_n376), .A2(KEYINPUT80), .A3(new_n377), .ZN(new_n378));
  AOI21_X1  g177(.A(new_n377), .B1(new_n376), .B2(KEYINPUT80), .ZN(new_n379));
  OAI21_X1  g178(.A(new_n374), .B1(new_n378), .B2(new_n379), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n376), .A2(KEYINPUT80), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n381), .A2(KEYINPUT81), .ZN(new_n382));
  INV_X1    g181(.A(new_n374), .ZN(new_n383));
  NAND3_X1  g182(.A1(new_n376), .A2(KEYINPUT80), .A3(new_n377), .ZN(new_n384));
  NAND3_X1  g183(.A1(new_n382), .A2(new_n383), .A3(new_n384), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n373), .A2(KEYINPUT3), .ZN(new_n386));
  INV_X1    g185(.A(KEYINPUT3), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n372), .A2(new_n387), .ZN(new_n388));
  NAND3_X1  g187(.A1(new_n386), .A2(new_n326), .A3(new_n388), .ZN(new_n389));
  NAND3_X1  g188(.A1(new_n380), .A2(new_n385), .A3(new_n389), .ZN(new_n390));
  NAND2_X1  g189(.A1(G225gat), .A2(G233gat), .ZN(new_n391));
  INV_X1    g190(.A(new_n391), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n390), .A2(new_n392), .ZN(new_n393));
  INV_X1    g192(.A(KEYINPUT39), .ZN(new_n394));
  XNOR2_X1  g193(.A(new_n326), .B(new_n373), .ZN(new_n395));
  INV_X1    g194(.A(new_n395), .ZN(new_n396));
  AOI21_X1  g195(.A(new_n394), .B1(new_n396), .B2(new_n391), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n393), .A2(new_n397), .ZN(new_n398));
  XNOR2_X1  g197(.A(G1gat), .B(G29gat), .ZN(new_n399));
  XNOR2_X1  g198(.A(new_n399), .B(KEYINPUT0), .ZN(new_n400));
  XNOR2_X1  g199(.A(G57gat), .B(G85gat), .ZN(new_n401));
  XOR2_X1   g200(.A(new_n400), .B(new_n401), .Z(new_n402));
  XOR2_X1   g201(.A(KEYINPUT85), .B(KEYINPUT39), .Z(new_n403));
  NAND3_X1  g202(.A1(new_n390), .A2(new_n392), .A3(new_n403), .ZN(new_n404));
  NAND3_X1  g203(.A1(new_n398), .A2(new_n402), .A3(new_n404), .ZN(new_n405));
  INV_X1    g204(.A(KEYINPUT40), .ZN(new_n406));
  INV_X1    g205(.A(new_n402), .ZN(new_n407));
  INV_X1    g206(.A(KEYINPUT5), .ZN(new_n408));
  NAND3_X1  g207(.A1(new_n389), .A2(new_n408), .A3(new_n391), .ZN(new_n409));
  INV_X1    g208(.A(new_n409), .ZN(new_n410));
  NAND3_X1  g209(.A1(new_n380), .A2(new_n385), .A3(new_n410), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n376), .A2(new_n374), .ZN(new_n412));
  NAND3_X1  g211(.A1(new_n412), .A2(new_n391), .A3(new_n389), .ZN(new_n413));
  AOI21_X1  g212(.A(new_n408), .B1(new_n395), .B2(new_n392), .ZN(new_n414));
  AND3_X1   g213(.A1(new_n413), .A2(new_n414), .A3(KEYINPUT79), .ZN(new_n415));
  AOI21_X1  g214(.A(KEYINPUT79), .B1(new_n413), .B2(new_n414), .ZN(new_n416));
  OAI21_X1  g215(.A(new_n411), .B1(new_n415), .B2(new_n416), .ZN(new_n417));
  AOI22_X1  g216(.A1(new_n405), .A2(new_n406), .B1(new_n407), .B2(new_n417), .ZN(new_n418));
  AND2_X1   g217(.A1(G226gat), .A2(G233gat), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n314), .A2(new_n419), .ZN(new_n420));
  AOI21_X1  g219(.A(new_n288), .B1(new_n309), .B2(new_n303), .ZN(new_n421));
  NOR2_X1   g220(.A1(new_n419), .A2(KEYINPUT29), .ZN(new_n422));
  INV_X1    g221(.A(new_n422), .ZN(new_n423));
  NOR2_X1   g222(.A1(new_n421), .A2(new_n423), .ZN(new_n424));
  INV_X1    g223(.A(new_n424), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n420), .A2(new_n425), .ZN(new_n426));
  INV_X1    g225(.A(KEYINPUT22), .ZN(new_n427));
  AOI22_X1  g226(.A1(new_n427), .A2(KEYINPUT76), .B1(G211gat), .B2(G218gat), .ZN(new_n428));
  OAI21_X1  g227(.A(new_n428), .B1(KEYINPUT76), .B2(new_n427), .ZN(new_n429));
  XNOR2_X1  g228(.A(G197gat), .B(G204gat), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n429), .A2(new_n430), .ZN(new_n431));
  XNOR2_X1  g230(.A(G211gat), .B(G218gat), .ZN(new_n432));
  XNOR2_X1  g231(.A(new_n431), .B(new_n432), .ZN(new_n433));
  INV_X1    g232(.A(new_n433), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n426), .A2(new_n434), .ZN(new_n435));
  INV_X1    g234(.A(KEYINPUT30), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n421), .A2(new_n419), .ZN(new_n437));
  XOR2_X1   g236(.A(new_n433), .B(KEYINPUT77), .Z(new_n438));
  OAI211_X1 g237(.A(new_n437), .B(new_n438), .C1(new_n314), .C2(new_n423), .ZN(new_n439));
  XNOR2_X1  g238(.A(G8gat), .B(G36gat), .ZN(new_n440));
  XNOR2_X1  g239(.A(G64gat), .B(G92gat), .ZN(new_n441));
  XOR2_X1   g240(.A(new_n440), .B(new_n441), .Z(new_n442));
  NAND4_X1  g241(.A1(new_n435), .A2(new_n436), .A3(new_n439), .A4(new_n442), .ZN(new_n443));
  INV_X1    g242(.A(new_n442), .ZN(new_n444));
  INV_X1    g243(.A(new_n439), .ZN(new_n445));
  AOI21_X1  g244(.A(new_n433), .B1(new_n420), .B2(new_n425), .ZN(new_n446));
  OAI21_X1  g245(.A(new_n444), .B1(new_n445), .B2(new_n446), .ZN(new_n447));
  AOI21_X1  g246(.A(new_n424), .B1(new_n314), .B2(new_n419), .ZN(new_n448));
  OAI211_X1 g247(.A(new_n439), .B(new_n442), .C1(new_n448), .C2(new_n433), .ZN(new_n449));
  NAND3_X1  g248(.A1(new_n447), .A2(KEYINPUT30), .A3(new_n449), .ZN(new_n450));
  NAND4_X1  g249(.A1(new_n398), .A2(KEYINPUT40), .A3(new_n402), .A4(new_n404), .ZN(new_n451));
  NAND4_X1  g250(.A1(new_n418), .A2(new_n443), .A3(new_n450), .A4(new_n451), .ZN(new_n452));
  INV_X1    g251(.A(KEYINPUT29), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n434), .A2(new_n453), .ZN(new_n454));
  AOI21_X1  g253(.A(new_n372), .B1(new_n454), .B2(new_n387), .ZN(new_n455));
  AOI21_X1  g254(.A(new_n434), .B1(new_n388), .B2(new_n453), .ZN(new_n456));
  INV_X1    g255(.A(G228gat), .ZN(new_n457));
  OAI22_X1  g256(.A1(new_n455), .A2(new_n456), .B1(new_n457), .B2(new_n332), .ZN(new_n458));
  OR2_X1    g257(.A1(new_n458), .A2(KEYINPUT83), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n458), .A2(KEYINPUT83), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  NOR3_X1   g260(.A1(new_n455), .A2(new_n457), .A3(new_n332), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n388), .A2(new_n453), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n438), .A2(new_n463), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n462), .A2(new_n464), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n461), .A2(new_n465), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n466), .A2(G22gat), .ZN(new_n467));
  AOI22_X1  g266(.A1(new_n459), .A2(new_n460), .B1(new_n464), .B2(new_n462), .ZN(new_n468));
  INV_X1    g267(.A(G22gat), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n467), .A2(new_n470), .ZN(new_n471));
  INV_X1    g270(.A(KEYINPUT84), .ZN(new_n472));
  AOI21_X1  g271(.A(new_n472), .B1(new_n468), .B2(new_n469), .ZN(new_n473));
  XNOR2_X1  g272(.A(KEYINPUT31), .B(G50gat), .ZN(new_n474));
  XNOR2_X1  g273(.A(new_n474), .B(KEYINPUT82), .ZN(new_n475));
  XOR2_X1   g274(.A(G78gat), .B(G106gat), .Z(new_n476));
  XOR2_X1   g275(.A(new_n475), .B(new_n476), .Z(new_n477));
  INV_X1    g276(.A(new_n477), .ZN(new_n478));
  OAI21_X1  g277(.A(new_n471), .B1(new_n473), .B2(new_n478), .ZN(new_n479));
  NAND4_X1  g278(.A1(new_n467), .A2(new_n470), .A3(new_n472), .A4(new_n477), .ZN(new_n480));
  AND2_X1   g279(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  INV_X1    g280(.A(KEYINPUT37), .ZN(new_n482));
  NAND4_X1  g281(.A1(new_n435), .A2(KEYINPUT86), .A3(new_n482), .A4(new_n439), .ZN(new_n483));
  OAI211_X1 g282(.A(new_n439), .B(new_n482), .C1(new_n448), .C2(new_n433), .ZN(new_n484));
  INV_X1    g283(.A(KEYINPUT86), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n483), .A2(new_n486), .ZN(new_n487));
  INV_X1    g286(.A(KEYINPUT38), .ZN(new_n488));
  NAND2_X1  g287(.A1(new_n444), .A2(new_n488), .ZN(new_n489));
  AOI22_X1  g288(.A1(new_n336), .A2(new_n422), .B1(new_n419), .B2(new_n421), .ZN(new_n490));
  OAI22_X1  g289(.A1(new_n490), .A2(new_n438), .B1(new_n426), .B2(new_n434), .ZN(new_n491));
  AOI21_X1  g290(.A(new_n489), .B1(new_n491), .B2(KEYINPUT37), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n487), .A2(new_n492), .ZN(new_n493));
  NAND3_X1  g292(.A1(new_n417), .A2(KEYINPUT6), .A3(new_n407), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n417), .A2(new_n407), .ZN(new_n495));
  INV_X1    g294(.A(KEYINPUT6), .ZN(new_n496));
  OAI211_X1 g295(.A(new_n411), .B(new_n402), .C1(new_n416), .C2(new_n415), .ZN(new_n497));
  NAND3_X1  g296(.A1(new_n495), .A2(new_n496), .A3(new_n497), .ZN(new_n498));
  NAND4_X1  g297(.A1(new_n493), .A2(new_n494), .A3(new_n498), .A4(new_n449), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n435), .A2(new_n439), .ZN(new_n500));
  AOI21_X1  g299(.A(new_n442), .B1(new_n500), .B2(KEYINPUT37), .ZN(new_n501));
  AOI21_X1  g300(.A(new_n488), .B1(new_n487), .B2(new_n501), .ZN(new_n502));
  OAI211_X1 g301(.A(new_n452), .B(new_n481), .C1(new_n499), .C2(new_n502), .ZN(new_n503));
  AOI22_X1  g302(.A1(new_n494), .A2(new_n498), .B1(new_n450), .B2(new_n443), .ZN(new_n504));
  OR2_X1    g303(.A1(new_n504), .A2(new_n481), .ZN(new_n505));
  NAND3_X1  g304(.A1(new_n365), .A2(new_n503), .A3(new_n505), .ZN(new_n506));
  NOR2_X1   g305(.A1(new_n358), .A2(new_n359), .ZN(new_n507));
  INV_X1    g306(.A(KEYINPUT35), .ZN(new_n508));
  NAND4_X1  g307(.A1(new_n507), .A2(new_n508), .A3(new_n481), .A4(new_n504), .ZN(new_n509));
  NAND4_X1  g308(.A1(new_n362), .A2(new_n504), .A3(new_n481), .A4(new_n363), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n510), .A2(KEYINPUT35), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n509), .A2(new_n511), .ZN(new_n512));
  AOI21_X1  g311(.A(new_n265), .B1(new_n506), .B2(new_n512), .ZN(new_n513));
  NAND2_X1  g312(.A1(G71gat), .A2(G78gat), .ZN(new_n514));
  INV_X1    g313(.A(KEYINPUT9), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  OR2_X1    g315(.A1(G57gat), .A2(G64gat), .ZN(new_n517));
  NAND2_X1  g316(.A1(G57gat), .A2(G64gat), .ZN(new_n518));
  NAND3_X1  g317(.A1(new_n516), .A2(new_n517), .A3(new_n518), .ZN(new_n519));
  NAND3_X1  g318(.A1(new_n517), .A2(KEYINPUT94), .A3(new_n518), .ZN(new_n520));
  XNOR2_X1  g319(.A(G71gat), .B(G78gat), .ZN(new_n521));
  NAND3_X1  g320(.A1(new_n519), .A2(new_n520), .A3(new_n521), .ZN(new_n522));
  AND2_X1   g321(.A1(G57gat), .A2(G64gat), .ZN(new_n523));
  NOR2_X1   g322(.A1(G57gat), .A2(G64gat), .ZN(new_n524));
  NOR2_X1   g323(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  AND2_X1   g324(.A1(G71gat), .A2(G78gat), .ZN(new_n526));
  NOR2_X1   g325(.A1(G71gat), .A2(G78gat), .ZN(new_n527));
  NOR2_X1   g326(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  OAI211_X1 g327(.A(new_n516), .B(new_n525), .C1(new_n528), .C2(KEYINPUT94), .ZN(new_n529));
  NAND2_X1  g328(.A1(new_n522), .A2(new_n529), .ZN(new_n530));
  AOI21_X1  g329(.A(new_n235), .B1(KEYINPUT21), .B2(new_n530), .ZN(new_n531));
  XNOR2_X1  g330(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n532));
  XNOR2_X1  g331(.A(new_n532), .B(new_n367), .ZN(new_n533));
  INV_X1    g332(.A(new_n533), .ZN(new_n534));
  OR2_X1    g333(.A1(new_n530), .A2(KEYINPUT21), .ZN(new_n535));
  AND2_X1   g334(.A1(G231gat), .A2(G233gat), .ZN(new_n536));
  OR2_X1    g335(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n535), .A2(new_n536), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n539), .A2(G127gat), .ZN(new_n540));
  XOR2_X1   g339(.A(G183gat), .B(G211gat), .Z(new_n541));
  INV_X1    g340(.A(new_n541), .ZN(new_n542));
  INV_X1    g341(.A(G127gat), .ZN(new_n543));
  NAND3_X1  g342(.A1(new_n537), .A2(new_n543), .A3(new_n538), .ZN(new_n544));
  NAND3_X1  g343(.A1(new_n540), .A2(new_n542), .A3(new_n544), .ZN(new_n545));
  INV_X1    g344(.A(new_n545), .ZN(new_n546));
  AOI21_X1  g345(.A(new_n542), .B1(new_n540), .B2(new_n544), .ZN(new_n547));
  OAI21_X1  g346(.A(new_n534), .B1(new_n546), .B2(new_n547), .ZN(new_n548));
  INV_X1    g347(.A(new_n548), .ZN(new_n549));
  NOR3_X1   g348(.A1(new_n546), .A2(new_n534), .A3(new_n547), .ZN(new_n550));
  OAI21_X1  g349(.A(new_n531), .B1(new_n549), .B2(new_n550), .ZN(new_n551));
  INV_X1    g350(.A(new_n550), .ZN(new_n552));
  INV_X1    g351(.A(new_n531), .ZN(new_n553));
  NAND3_X1  g352(.A1(new_n552), .A2(new_n553), .A3(new_n548), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n551), .A2(new_n554), .ZN(new_n555));
  XNOR2_X1  g354(.A(KEYINPUT95), .B(KEYINPUT96), .ZN(new_n556));
  INV_X1    g355(.A(new_n556), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n555), .A2(new_n557), .ZN(new_n558));
  NAND3_X1  g357(.A1(new_n551), .A2(new_n554), .A3(new_n556), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  OR2_X1    g359(.A1(new_n228), .A2(new_n230), .ZN(new_n561));
  NAND2_X1  g360(.A1(G85gat), .A2(G92gat), .ZN(new_n562));
  NAND2_X1  g361(.A1(KEYINPUT97), .A2(KEYINPUT7), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  NAND2_X1  g363(.A1(G99gat), .A2(G106gat), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n565), .A2(KEYINPUT8), .ZN(new_n566));
  INV_X1    g365(.A(G85gat), .ZN(new_n567));
  INV_X1    g366(.A(G92gat), .ZN(new_n568));
  NAND2_X1  g367(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  NAND4_X1  g368(.A1(KEYINPUT97), .A2(KEYINPUT7), .A3(G85gat), .A4(G92gat), .ZN(new_n570));
  NAND4_X1  g369(.A1(new_n564), .A2(new_n566), .A3(new_n569), .A4(new_n570), .ZN(new_n571));
  XNOR2_X1  g370(.A(G99gat), .B(G106gat), .ZN(new_n572));
  INV_X1    g371(.A(new_n572), .ZN(new_n573));
  NAND2_X1  g372(.A1(new_n571), .A2(new_n573), .ZN(new_n574));
  AOI22_X1  g373(.A1(KEYINPUT8), .A2(new_n565), .B1(new_n567), .B2(new_n568), .ZN(new_n575));
  NAND4_X1  g374(.A1(new_n575), .A2(new_n572), .A3(new_n564), .A4(new_n570), .ZN(new_n576));
  NAND3_X1  g375(.A1(new_n574), .A2(KEYINPUT98), .A3(new_n576), .ZN(new_n577));
  AND2_X1   g376(.A1(new_n564), .A2(new_n570), .ZN(new_n578));
  INV_X1    g377(.A(KEYINPUT98), .ZN(new_n579));
  NAND4_X1  g378(.A1(new_n578), .A2(new_n579), .A3(new_n572), .A4(new_n575), .ZN(new_n580));
  NAND2_X1  g379(.A1(new_n577), .A2(new_n580), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n581), .A2(KEYINPUT99), .ZN(new_n582));
  INV_X1    g381(.A(KEYINPUT99), .ZN(new_n583));
  NAND3_X1  g382(.A1(new_n577), .A2(new_n583), .A3(new_n580), .ZN(new_n584));
  NAND2_X1  g383(.A1(new_n582), .A2(new_n584), .ZN(new_n585));
  NAND2_X1  g384(.A1(new_n561), .A2(new_n585), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n586), .A2(KEYINPUT100), .ZN(new_n587));
  INV_X1    g386(.A(KEYINPUT100), .ZN(new_n588));
  NAND3_X1  g387(.A1(new_n561), .A2(new_n588), .A3(new_n585), .ZN(new_n589));
  NAND2_X1  g388(.A1(new_n587), .A2(new_n589), .ZN(new_n590));
  AND2_X1   g389(.A1(G232gat), .A2(G233gat), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n591), .A2(KEYINPUT41), .ZN(new_n592));
  OAI21_X1  g391(.A(new_n592), .B1(new_n585), .B2(new_n244), .ZN(new_n593));
  INV_X1    g392(.A(new_n593), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n590), .A2(new_n594), .ZN(new_n595));
  XOR2_X1   g394(.A(G190gat), .B(G218gat), .Z(new_n596));
  NAND2_X1  g395(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  NOR2_X1   g396(.A1(new_n591), .A2(KEYINPUT41), .ZN(new_n598));
  XNOR2_X1  g397(.A(G134gat), .B(G162gat), .ZN(new_n599));
  XNOR2_X1  g398(.A(new_n598), .B(new_n599), .ZN(new_n600));
  INV_X1    g399(.A(new_n596), .ZN(new_n601));
  NAND3_X1  g400(.A1(new_n590), .A2(new_n601), .A3(new_n594), .ZN(new_n602));
  NAND3_X1  g401(.A1(new_n597), .A2(new_n600), .A3(new_n602), .ZN(new_n603));
  INV_X1    g402(.A(new_n600), .ZN(new_n604));
  AOI21_X1  g403(.A(new_n601), .B1(new_n590), .B2(new_n594), .ZN(new_n605));
  AOI211_X1 g404(.A(new_n596), .B(new_n593), .C1(new_n587), .C2(new_n589), .ZN(new_n606));
  OAI21_X1  g405(.A(new_n604), .B1(new_n605), .B2(new_n606), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n603), .A2(new_n607), .ZN(new_n608));
  INV_X1    g407(.A(new_n608), .ZN(new_n609));
  XOR2_X1   g408(.A(G120gat), .B(G148gat), .Z(new_n610));
  XNOR2_X1  g409(.A(G176gat), .B(G204gat), .ZN(new_n611));
  XNOR2_X1  g410(.A(new_n610), .B(new_n611), .ZN(new_n612));
  XNOR2_X1  g411(.A(KEYINPUT103), .B(KEYINPUT104), .ZN(new_n613));
  XOR2_X1   g412(.A(new_n612), .B(new_n613), .Z(new_n614));
  INV_X1    g413(.A(new_n614), .ZN(new_n615));
  INV_X1    g414(.A(KEYINPUT10), .ZN(new_n616));
  AOI21_X1  g415(.A(new_n616), .B1(new_n522), .B2(new_n529), .ZN(new_n617));
  NAND3_X1  g416(.A1(new_n582), .A2(new_n584), .A3(new_n617), .ZN(new_n618));
  INV_X1    g417(.A(KEYINPUT102), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  NAND4_X1  g419(.A1(new_n582), .A2(KEYINPUT102), .A3(new_n584), .A4(new_n617), .ZN(new_n621));
  AOI21_X1  g420(.A(new_n530), .B1(new_n577), .B2(new_n580), .ZN(new_n622));
  AOI22_X1  g421(.A1(new_n576), .A2(new_n574), .B1(new_n522), .B2(new_n529), .ZN(new_n623));
  OAI21_X1  g422(.A(new_n616), .B1(new_n622), .B2(new_n623), .ZN(new_n624));
  NAND2_X1  g423(.A1(new_n624), .A2(KEYINPUT101), .ZN(new_n625));
  INV_X1    g424(.A(KEYINPUT101), .ZN(new_n626));
  OAI211_X1 g425(.A(new_n626), .B(new_n616), .C1(new_n622), .C2(new_n623), .ZN(new_n627));
  AOI22_X1  g426(.A1(new_n620), .A2(new_n621), .B1(new_n625), .B2(new_n627), .ZN(new_n628));
  NAND2_X1  g427(.A1(G230gat), .A2(G233gat), .ZN(new_n629));
  XOR2_X1   g428(.A(new_n629), .B(KEYINPUT105), .Z(new_n630));
  NOR2_X1   g429(.A1(new_n628), .A2(new_n630), .ZN(new_n631));
  NOR3_X1   g430(.A1(new_n622), .A2(new_n623), .A3(new_n629), .ZN(new_n632));
  OAI21_X1  g431(.A(new_n615), .B1(new_n631), .B2(new_n632), .ZN(new_n633));
  NAND2_X1  g432(.A1(new_n620), .A2(new_n621), .ZN(new_n634));
  NAND2_X1  g433(.A1(new_n625), .A2(new_n627), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n636), .A2(new_n629), .ZN(new_n637));
  NOR2_X1   g436(.A1(new_n615), .A2(new_n632), .ZN(new_n638));
  NAND2_X1  g437(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n633), .A2(new_n639), .ZN(new_n640));
  NOR3_X1   g439(.A1(new_n560), .A2(new_n609), .A3(new_n640), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n513), .A2(new_n641), .ZN(new_n642));
  INV_X1    g441(.A(new_n642), .ZN(new_n643));
  NAND2_X1  g442(.A1(new_n498), .A2(new_n494), .ZN(new_n644));
  INV_X1    g443(.A(new_n644), .ZN(new_n645));
  NAND2_X1  g444(.A1(new_n643), .A2(new_n645), .ZN(new_n646));
  XNOR2_X1  g445(.A(new_n646), .B(G1gat), .ZN(G1324gat));
  NAND2_X1  g446(.A1(new_n450), .A2(new_n443), .ZN(new_n648));
  NOR2_X1   g447(.A1(new_n642), .A2(new_n648), .ZN(new_n649));
  XOR2_X1   g448(.A(KEYINPUT16), .B(G8gat), .Z(new_n650));
  AND2_X1   g449(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  AND3_X1   g450(.A1(new_n651), .A2(KEYINPUT106), .A3(KEYINPUT42), .ZN(new_n652));
  INV_X1    g451(.A(new_n651), .ZN(new_n653));
  OAI21_X1  g452(.A(KEYINPUT42), .B1(new_n649), .B2(new_n212), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  AOI21_X1  g454(.A(KEYINPUT106), .B1(new_n651), .B2(KEYINPUT42), .ZN(new_n656));
  AOI21_X1  g455(.A(new_n652), .B1(new_n655), .B2(new_n656), .ZN(G1325gat));
  OAI21_X1  g456(.A(G15gat), .B1(new_n642), .B2(new_n365), .ZN(new_n658));
  INV_X1    g457(.A(new_n507), .ZN(new_n659));
  OR2_X1    g458(.A1(new_n659), .A2(G15gat), .ZN(new_n660));
  OAI21_X1  g459(.A(new_n658), .B1(new_n642), .B2(new_n660), .ZN(G1326gat));
  NOR2_X1   g460(.A1(new_n642), .A2(new_n481), .ZN(new_n662));
  XNOR2_X1  g461(.A(new_n662), .B(KEYINPUT107), .ZN(new_n663));
  XNOR2_X1  g462(.A(KEYINPUT43), .B(G22gat), .ZN(new_n664));
  XNOR2_X1  g463(.A(new_n663), .B(new_n664), .ZN(G1327gat));
  NAND2_X1  g464(.A1(new_n506), .A2(new_n512), .ZN(new_n666));
  INV_X1    g465(.A(new_n640), .ZN(new_n667));
  NAND3_X1  g466(.A1(new_n560), .A2(new_n609), .A3(new_n667), .ZN(new_n668));
  XOR2_X1   g467(.A(new_n668), .B(KEYINPUT108), .Z(new_n669));
  AND3_X1   g468(.A1(new_n666), .A2(new_n264), .A3(new_n669), .ZN(new_n670));
  NAND3_X1  g469(.A1(new_n670), .A2(new_n220), .A3(new_n645), .ZN(new_n671));
  XNOR2_X1  g470(.A(new_n671), .B(KEYINPUT45), .ZN(new_n672));
  AOI21_X1  g471(.A(new_n608), .B1(new_n506), .B2(new_n512), .ZN(new_n673));
  INV_X1    g472(.A(KEYINPUT44), .ZN(new_n674));
  XNOR2_X1  g473(.A(new_n673), .B(new_n674), .ZN(new_n675));
  AND3_X1   g474(.A1(new_n558), .A2(KEYINPUT109), .A3(new_n559), .ZN(new_n676));
  AOI21_X1  g475(.A(KEYINPUT109), .B1(new_n558), .B2(new_n559), .ZN(new_n677));
  XOR2_X1   g476(.A(new_n640), .B(KEYINPUT110), .Z(new_n678));
  INV_X1    g477(.A(new_n678), .ZN(new_n679));
  NOR4_X1   g478(.A1(new_n676), .A2(new_n677), .A3(new_n265), .A4(new_n679), .ZN(new_n680));
  NAND2_X1  g479(.A1(new_n675), .A2(new_n680), .ZN(new_n681));
  OAI21_X1  g480(.A(G29gat), .B1(new_n681), .B2(new_n644), .ZN(new_n682));
  NAND2_X1  g481(.A1(new_n672), .A2(new_n682), .ZN(G1328gat));
  INV_X1    g482(.A(new_n670), .ZN(new_n684));
  NOR3_X1   g483(.A1(new_n684), .A2(G36gat), .A3(new_n648), .ZN(new_n685));
  XNOR2_X1  g484(.A(new_n685), .B(KEYINPUT46), .ZN(new_n686));
  OAI21_X1  g485(.A(G36gat), .B1(new_n681), .B2(new_n648), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n686), .A2(new_n687), .ZN(G1329gat));
  INV_X1    g487(.A(G43gat), .ZN(new_n689));
  OAI21_X1  g488(.A(new_n689), .B1(new_n684), .B2(new_n659), .ZN(new_n690));
  INV_X1    g489(.A(new_n365), .ZN(new_n691));
  NAND2_X1  g490(.A1(new_n691), .A2(G43gat), .ZN(new_n692));
  OAI21_X1  g491(.A(new_n690), .B1(new_n681), .B2(new_n692), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n693), .A2(KEYINPUT47), .ZN(new_n694));
  INV_X1    g493(.A(KEYINPUT47), .ZN(new_n695));
  OAI211_X1 g494(.A(new_n695), .B(new_n690), .C1(new_n681), .C2(new_n692), .ZN(new_n696));
  NAND2_X1  g495(.A1(new_n694), .A2(new_n696), .ZN(G1330gat));
  NAND2_X1  g496(.A1(new_n670), .A2(KEYINPUT112), .ZN(new_n698));
  NOR2_X1   g497(.A1(new_n481), .A2(G50gat), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  NOR2_X1   g499(.A1(new_n670), .A2(KEYINPUT112), .ZN(new_n701));
  OAI21_X1  g500(.A(KEYINPUT113), .B1(new_n700), .B2(new_n701), .ZN(new_n702));
  OR2_X1    g501(.A1(new_n673), .A2(KEYINPUT44), .ZN(new_n703));
  INV_X1    g502(.A(new_n481), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n673), .A2(KEYINPUT44), .ZN(new_n705));
  NAND4_X1  g504(.A1(new_n703), .A2(new_n704), .A3(new_n705), .A4(new_n680), .ZN(new_n706));
  NAND2_X1  g505(.A1(new_n706), .A2(G50gat), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n702), .A2(new_n707), .ZN(new_n708));
  OR2_X1    g507(.A1(new_n670), .A2(KEYINPUT112), .ZN(new_n709));
  INV_X1    g508(.A(KEYINPUT113), .ZN(new_n710));
  NAND4_X1  g509(.A1(new_n709), .A2(new_n710), .A3(new_n698), .A4(new_n699), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n711), .A2(KEYINPUT48), .ZN(new_n712));
  AND2_X1   g511(.A1(new_n698), .A2(new_n699), .ZN(new_n713));
  AOI22_X1  g512(.A1(new_n713), .A2(new_n709), .B1(new_n706), .B2(G50gat), .ZN(new_n714));
  XNOR2_X1  g513(.A(KEYINPUT111), .B(KEYINPUT48), .ZN(new_n715));
  OAI22_X1  g514(.A1(new_n708), .A2(new_n712), .B1(new_n714), .B2(new_n715), .ZN(G1331gat));
  INV_X1    g515(.A(new_n560), .ZN(new_n717));
  NAND4_X1  g516(.A1(new_n717), .A2(new_n265), .A3(new_n608), .A4(new_n679), .ZN(new_n718));
  AOI21_X1  g517(.A(new_n718), .B1(new_n506), .B2(new_n512), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n719), .A2(new_n645), .ZN(new_n720));
  XNOR2_X1  g519(.A(new_n720), .B(G57gat), .ZN(G1332gat));
  INV_X1    g520(.A(new_n648), .ZN(new_n722));
  AND2_X1   g521(.A1(new_n719), .A2(new_n722), .ZN(new_n723));
  NOR2_X1   g522(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n724));
  AND2_X1   g523(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n725));
  OAI21_X1  g524(.A(new_n723), .B1(new_n724), .B2(new_n725), .ZN(new_n726));
  OAI21_X1  g525(.A(new_n726), .B1(new_n723), .B2(new_n724), .ZN(new_n727));
  XNOR2_X1  g526(.A(new_n727), .B(KEYINPUT114), .ZN(G1333gat));
  NAND2_X1  g527(.A1(new_n719), .A2(new_n691), .ZN(new_n729));
  NOR2_X1   g528(.A1(new_n659), .A2(G71gat), .ZN(new_n730));
  AOI22_X1  g529(.A1(new_n729), .A2(G71gat), .B1(new_n719), .B2(new_n730), .ZN(new_n731));
  XNOR2_X1  g530(.A(new_n731), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g531(.A1(new_n719), .A2(new_n704), .ZN(new_n733));
  XNOR2_X1  g532(.A(KEYINPUT115), .B(G78gat), .ZN(new_n734));
  XNOR2_X1  g533(.A(new_n733), .B(new_n734), .ZN(G1335gat));
  NOR2_X1   g534(.A1(new_n717), .A2(new_n264), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n736), .A2(new_n640), .ZN(new_n737));
  XOR2_X1   g536(.A(new_n737), .B(KEYINPUT116), .Z(new_n738));
  NAND2_X1  g537(.A1(new_n675), .A2(new_n738), .ZN(new_n739));
  OAI21_X1  g538(.A(G85gat), .B1(new_n739), .B2(new_n644), .ZN(new_n740));
  NAND4_X1  g539(.A1(new_n666), .A2(KEYINPUT51), .A3(new_n609), .A4(new_n736), .ZN(new_n741));
  INV_X1    g540(.A(KEYINPUT117), .ZN(new_n742));
  NAND2_X1  g541(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  NAND3_X1  g542(.A1(new_n666), .A2(new_n609), .A3(new_n736), .ZN(new_n744));
  INV_X1    g543(.A(KEYINPUT51), .ZN(new_n745));
  NAND2_X1  g544(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  NAND4_X1  g545(.A1(new_n673), .A2(KEYINPUT117), .A3(KEYINPUT51), .A4(new_n736), .ZN(new_n747));
  NAND3_X1  g546(.A1(new_n743), .A2(new_n746), .A3(new_n747), .ZN(new_n748));
  INV_X1    g547(.A(new_n748), .ZN(new_n749));
  NAND3_X1  g548(.A1(new_n645), .A2(new_n567), .A3(new_n640), .ZN(new_n750));
  OAI21_X1  g549(.A(new_n740), .B1(new_n749), .B2(new_n750), .ZN(G1336gat));
  NAND4_X1  g550(.A1(new_n703), .A2(new_n722), .A3(new_n705), .A4(new_n738), .ZN(new_n752));
  AOI21_X1  g551(.A(KEYINPUT52), .B1(new_n752), .B2(G92gat), .ZN(new_n753));
  INV_X1    g552(.A(KEYINPUT118), .ZN(new_n754));
  NOR3_X1   g553(.A1(new_n648), .A2(G92gat), .A3(new_n678), .ZN(new_n755));
  AND3_X1   g554(.A1(new_n748), .A2(new_n754), .A3(new_n755), .ZN(new_n756));
  AOI21_X1  g555(.A(new_n754), .B1(new_n748), .B2(new_n755), .ZN(new_n757));
  OAI21_X1  g556(.A(new_n753), .B1(new_n756), .B2(new_n757), .ZN(new_n758));
  AND2_X1   g557(.A1(new_n752), .A2(G92gat), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n746), .A2(new_n741), .ZN(new_n760));
  AND2_X1   g559(.A1(new_n760), .A2(new_n755), .ZN(new_n761));
  OAI21_X1  g560(.A(KEYINPUT52), .B1(new_n759), .B2(new_n761), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n758), .A2(new_n762), .ZN(G1337gat));
  OAI21_X1  g562(.A(G99gat), .B1(new_n739), .B2(new_n365), .ZN(new_n764));
  OR3_X1    g563(.A1(new_n659), .A2(G99gat), .A3(new_n667), .ZN(new_n765));
  OAI21_X1  g564(.A(new_n764), .B1(new_n749), .B2(new_n765), .ZN(G1338gat));
  NAND3_X1  g565(.A1(new_n675), .A2(new_n704), .A3(new_n738), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n767), .A2(G106gat), .ZN(new_n768));
  INV_X1    g567(.A(KEYINPUT53), .ZN(new_n769));
  NAND2_X1  g568(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  NOR3_X1   g569(.A1(new_n481), .A2(G106gat), .A3(new_n678), .ZN(new_n771));
  AND2_X1   g570(.A1(new_n748), .A2(new_n771), .ZN(new_n772));
  AOI22_X1  g571(.A1(new_n767), .A2(G106gat), .B1(new_n760), .B2(new_n771), .ZN(new_n773));
  OAI22_X1  g572(.A1(new_n770), .A2(new_n772), .B1(new_n773), .B2(new_n769), .ZN(G1339gat));
  NOR2_X1   g573(.A1(new_n676), .A2(new_n677), .ZN(new_n775));
  INV_X1    g574(.A(KEYINPUT55), .ZN(new_n776));
  INV_X1    g575(.A(KEYINPUT54), .ZN(new_n777));
  INV_X1    g576(.A(new_n630), .ZN(new_n778));
  NAND3_X1  g577(.A1(new_n636), .A2(new_n777), .A3(new_n778), .ZN(new_n779));
  NAND2_X1  g578(.A1(new_n779), .A2(new_n615), .ZN(new_n780));
  INV_X1    g579(.A(new_n629), .ZN(new_n781));
  OAI21_X1  g580(.A(KEYINPUT54), .B1(new_n628), .B2(new_n781), .ZN(new_n782));
  AND3_X1   g581(.A1(new_n634), .A2(new_n630), .A3(new_n635), .ZN(new_n783));
  OAI21_X1  g582(.A(KEYINPUT119), .B1(new_n782), .B2(new_n783), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n628), .A2(new_n630), .ZN(new_n785));
  INV_X1    g584(.A(KEYINPUT119), .ZN(new_n786));
  NAND4_X1  g585(.A1(new_n637), .A2(new_n785), .A3(new_n786), .A4(KEYINPUT54), .ZN(new_n787));
  AOI211_X1 g586(.A(new_n776), .B(new_n780), .C1(new_n784), .C2(new_n787), .ZN(new_n788));
  INV_X1    g587(.A(new_n639), .ZN(new_n789));
  OAI21_X1  g588(.A(KEYINPUT120), .B1(new_n788), .B2(new_n789), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n784), .A2(new_n787), .ZN(new_n791));
  INV_X1    g590(.A(new_n780), .ZN(new_n792));
  NAND3_X1  g591(.A1(new_n791), .A2(KEYINPUT55), .A3(new_n792), .ZN(new_n793));
  INV_X1    g592(.A(KEYINPUT120), .ZN(new_n794));
  NAND3_X1  g593(.A1(new_n793), .A2(new_n794), .A3(new_n639), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n791), .A2(new_n792), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n796), .A2(new_n776), .ZN(new_n797));
  NAND4_X1  g596(.A1(new_n790), .A2(new_n264), .A3(new_n795), .A4(new_n797), .ZN(new_n798));
  NOR2_X1   g597(.A1(new_n246), .A2(new_n247), .ZN(new_n799));
  NOR2_X1   g598(.A1(new_n239), .A2(new_n241), .ZN(new_n800));
  OAI21_X1  g599(.A(new_n206), .B1(new_n799), .B2(new_n800), .ZN(new_n801));
  NAND3_X1  g600(.A1(new_n263), .A2(new_n640), .A3(new_n801), .ZN(new_n802));
  AOI21_X1  g601(.A(new_n609), .B1(new_n798), .B2(new_n802), .ZN(new_n803));
  NAND3_X1  g602(.A1(new_n790), .A2(new_n795), .A3(new_n797), .ZN(new_n804));
  NAND3_X1  g603(.A1(new_n609), .A2(new_n263), .A3(new_n801), .ZN(new_n805));
  NOR2_X1   g604(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  OAI21_X1  g605(.A(new_n775), .B1(new_n803), .B2(new_n806), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n641), .A2(new_n265), .ZN(new_n808));
  NAND3_X1  g607(.A1(new_n807), .A2(KEYINPUT121), .A3(new_n808), .ZN(new_n809));
  INV_X1    g608(.A(new_n809), .ZN(new_n810));
  AOI21_X1  g609(.A(KEYINPUT121), .B1(new_n807), .B2(new_n808), .ZN(new_n811));
  NOR2_X1   g610(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  NOR2_X1   g611(.A1(new_n659), .A2(new_n704), .ZN(new_n813));
  AND2_X1   g612(.A1(new_n812), .A2(new_n813), .ZN(new_n814));
  NOR2_X1   g613(.A1(new_n722), .A2(new_n644), .ZN(new_n815));
  AND2_X1   g614(.A1(new_n814), .A2(new_n815), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n816), .A2(new_n264), .ZN(new_n817));
  XNOR2_X1  g616(.A(new_n817), .B(G113gat), .ZN(G1340gat));
  AOI21_X1  g617(.A(G120gat), .B1(new_n816), .B2(new_n640), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n814), .A2(new_n815), .ZN(new_n820));
  NOR3_X1   g619(.A1(new_n820), .A2(new_n319), .A3(new_n678), .ZN(new_n821));
  NOR2_X1   g620(.A1(new_n819), .A2(new_n821), .ZN(G1341gat));
  OAI21_X1  g621(.A(G127gat), .B1(new_n820), .B2(new_n775), .ZN(new_n823));
  NAND4_X1  g622(.A1(new_n814), .A2(new_n543), .A3(new_n717), .A4(new_n815), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  INV_X1    g624(.A(KEYINPUT122), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n825), .A2(new_n826), .ZN(new_n827));
  NAND3_X1  g626(.A1(new_n823), .A2(KEYINPUT122), .A3(new_n824), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n827), .A2(new_n828), .ZN(G1342gat));
  XOR2_X1   g628(.A(KEYINPUT123), .B(KEYINPUT56), .Z(new_n830));
  INV_X1    g629(.A(new_n830), .ZN(new_n831));
  OR4_X1    g630(.A1(G134gat), .A2(new_n820), .A3(new_n608), .A4(new_n831), .ZN(new_n832));
  NAND2_X1  g631(.A1(new_n816), .A2(new_n609), .ZN(new_n833));
  OAI21_X1  g632(.A(new_n831), .B1(new_n833), .B2(G134gat), .ZN(new_n834));
  NAND2_X1  g633(.A1(new_n833), .A2(G134gat), .ZN(new_n835));
  NAND3_X1  g634(.A1(new_n832), .A2(new_n834), .A3(new_n835), .ZN(G1343gat));
  NAND3_X1  g635(.A1(new_n365), .A2(new_n645), .A3(new_n648), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n264), .A2(new_n797), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n793), .A2(new_n639), .ZN(new_n839));
  OAI21_X1  g638(.A(new_n802), .B1(new_n838), .B2(new_n839), .ZN(new_n840));
  AOI21_X1  g639(.A(new_n806), .B1(new_n608), .B2(new_n840), .ZN(new_n841));
  OAI21_X1  g640(.A(new_n808), .B1(new_n841), .B2(new_n717), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n842), .A2(new_n704), .ZN(new_n843));
  AOI21_X1  g642(.A(new_n837), .B1(new_n843), .B2(KEYINPUT57), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n812), .A2(new_n704), .ZN(new_n845));
  OAI21_X1  g644(.A(new_n844), .B1(new_n845), .B2(KEYINPUT57), .ZN(new_n846));
  OAI21_X1  g645(.A(G141gat), .B1(new_n846), .B2(new_n265), .ZN(new_n847));
  NOR2_X1   g646(.A1(new_n845), .A2(new_n837), .ZN(new_n848));
  NOR2_X1   g647(.A1(new_n265), .A2(G141gat), .ZN(new_n849));
  AOI22_X1  g648(.A1(new_n848), .A2(new_n849), .B1(KEYINPUT124), .B2(KEYINPUT58), .ZN(new_n850));
  OR2_X1    g649(.A1(KEYINPUT124), .A2(KEYINPUT58), .ZN(new_n851));
  AND3_X1   g650(.A1(new_n847), .A2(new_n850), .A3(new_n851), .ZN(new_n852));
  AOI21_X1  g651(.A(new_n851), .B1(new_n847), .B2(new_n850), .ZN(new_n853));
  NOR2_X1   g652(.A1(new_n852), .A2(new_n853), .ZN(G1344gat));
  INV_X1    g653(.A(KEYINPUT59), .ZN(new_n855));
  OAI211_X1 g654(.A(new_n855), .B(G148gat), .C1(new_n846), .C2(new_n667), .ZN(new_n856));
  INV_X1    g655(.A(G148gat), .ZN(new_n857));
  NOR3_X1   g656(.A1(new_n810), .A2(new_n811), .A3(new_n481), .ZN(new_n858));
  NAND2_X1  g657(.A1(new_n858), .A2(KEYINPUT57), .ZN(new_n859));
  INV_X1    g658(.A(KEYINPUT57), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n843), .A2(new_n860), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n859), .A2(new_n861), .ZN(new_n862));
  NOR2_X1   g661(.A1(new_n837), .A2(new_n667), .ZN(new_n863));
  AOI21_X1  g662(.A(new_n857), .B1(new_n862), .B2(new_n863), .ZN(new_n864));
  OAI21_X1  g663(.A(new_n856), .B1(new_n864), .B2(new_n855), .ZN(new_n865));
  NAND3_X1  g664(.A1(new_n848), .A2(new_n857), .A3(new_n640), .ZN(new_n866));
  NAND2_X1  g665(.A1(new_n865), .A2(new_n866), .ZN(G1345gat));
  OAI21_X1  g666(.A(G155gat), .B1(new_n846), .B2(new_n775), .ZN(new_n868));
  NAND3_X1  g667(.A1(new_n848), .A2(new_n367), .A3(new_n717), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  NAND2_X1  g669(.A1(new_n870), .A2(KEYINPUT125), .ZN(new_n871));
  INV_X1    g670(.A(KEYINPUT125), .ZN(new_n872));
  NAND3_X1  g671(.A1(new_n868), .A2(new_n872), .A3(new_n869), .ZN(new_n873));
  NAND2_X1  g672(.A1(new_n871), .A2(new_n873), .ZN(G1346gat));
  OAI21_X1  g673(.A(G162gat), .B1(new_n846), .B2(new_n608), .ZN(new_n875));
  NOR2_X1   g674(.A1(new_n608), .A2(G162gat), .ZN(new_n876));
  NAND4_X1  g675(.A1(new_n365), .A2(new_n645), .A3(new_n648), .A4(new_n876), .ZN(new_n877));
  OAI21_X1  g676(.A(new_n875), .B1(new_n845), .B2(new_n877), .ZN(G1347gat));
  NAND2_X1  g677(.A1(new_n807), .A2(new_n808), .ZN(new_n879));
  INV_X1    g678(.A(KEYINPUT121), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  NOR2_X1   g680(.A1(new_n645), .A2(new_n648), .ZN(new_n882));
  NAND4_X1  g681(.A1(new_n881), .A2(new_n813), .A3(new_n809), .A4(new_n882), .ZN(new_n883));
  NOR2_X1   g682(.A1(new_n883), .A2(new_n265), .ZN(new_n884));
  MUX2_X1   g683(.A(G169gat), .B(new_n294), .S(new_n884), .Z(G1348gat));
  OAI21_X1  g684(.A(G176gat), .B1(new_n883), .B2(new_n678), .ZN(new_n886));
  NAND2_X1  g685(.A1(new_n640), .A2(new_n283), .ZN(new_n887));
  OAI21_X1  g686(.A(new_n886), .B1(new_n883), .B2(new_n887), .ZN(G1349gat));
  INV_X1    g687(.A(KEYINPUT127), .ZN(new_n889));
  OAI21_X1  g688(.A(G183gat), .B1(new_n883), .B2(new_n775), .ZN(new_n890));
  AND2_X1   g689(.A1(new_n717), .A2(new_n268), .ZN(new_n891));
  NAND4_X1  g690(.A1(new_n812), .A2(new_n813), .A3(new_n882), .A4(new_n891), .ZN(new_n892));
  NAND2_X1  g691(.A1(new_n890), .A2(new_n892), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n893), .A2(KEYINPUT126), .ZN(new_n894));
  INV_X1    g693(.A(KEYINPUT126), .ZN(new_n895));
  NAND3_X1  g694(.A1(new_n890), .A2(new_n895), .A3(new_n892), .ZN(new_n896));
  AND4_X1   g695(.A1(new_n889), .A2(new_n894), .A3(KEYINPUT60), .A4(new_n896), .ZN(new_n897));
  INV_X1    g696(.A(KEYINPUT60), .ZN(new_n898));
  NAND3_X1  g697(.A1(new_n890), .A2(new_n898), .A3(new_n892), .ZN(new_n899));
  NAND2_X1  g698(.A1(new_n899), .A2(KEYINPUT127), .ZN(new_n900));
  AOI21_X1  g699(.A(new_n898), .B1(new_n893), .B2(KEYINPUT126), .ZN(new_n901));
  AOI21_X1  g700(.A(new_n900), .B1(new_n901), .B2(new_n896), .ZN(new_n902));
  NOR2_X1   g701(.A1(new_n897), .A2(new_n902), .ZN(G1350gat));
  OR2_X1    g702(.A1(new_n883), .A2(new_n608), .ZN(new_n904));
  AND2_X1   g703(.A1(new_n904), .A2(G190gat), .ZN(new_n905));
  OR2_X1    g704(.A1(new_n905), .A2(KEYINPUT61), .ZN(new_n906));
  NAND2_X1  g705(.A1(new_n905), .A2(KEYINPUT61), .ZN(new_n907));
  OAI211_X1 g706(.A(new_n906), .B(new_n907), .C1(new_n305), .C2(new_n904), .ZN(G1351gat));
  NAND2_X1  g707(.A1(new_n365), .A2(new_n882), .ZN(new_n909));
  INV_X1    g708(.A(new_n909), .ZN(new_n910));
  NAND2_X1  g709(.A1(new_n858), .A2(new_n910), .ZN(new_n911));
  INV_X1    g710(.A(new_n911), .ZN(new_n912));
  AOI21_X1  g711(.A(G197gat), .B1(new_n912), .B2(new_n264), .ZN(new_n913));
  AOI21_X1  g712(.A(new_n909), .B1(new_n859), .B2(new_n861), .ZN(new_n914));
  AND2_X1   g713(.A1(new_n264), .A2(G197gat), .ZN(new_n915));
  AOI21_X1  g714(.A(new_n913), .B1(new_n914), .B2(new_n915), .ZN(G1352gat));
  INV_X1    g715(.A(new_n914), .ZN(new_n917));
  OAI21_X1  g716(.A(G204gat), .B1(new_n917), .B2(new_n678), .ZN(new_n918));
  NOR3_X1   g717(.A1(new_n911), .A2(G204gat), .A3(new_n667), .ZN(new_n919));
  INV_X1    g718(.A(KEYINPUT62), .ZN(new_n920));
  OR2_X1    g719(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  NAND2_X1  g720(.A1(new_n919), .A2(new_n920), .ZN(new_n922));
  NAND3_X1  g721(.A1(new_n918), .A2(new_n921), .A3(new_n922), .ZN(G1353gat));
  INV_X1    g722(.A(G211gat), .ZN(new_n924));
  NAND3_X1  g723(.A1(new_n912), .A2(new_n924), .A3(new_n717), .ZN(new_n925));
  NAND2_X1  g724(.A1(new_n914), .A2(new_n717), .ZN(new_n926));
  AOI21_X1  g725(.A(KEYINPUT63), .B1(new_n926), .B2(G211gat), .ZN(new_n927));
  INV_X1    g726(.A(KEYINPUT63), .ZN(new_n928));
  AOI211_X1 g727(.A(new_n928), .B(new_n924), .C1(new_n914), .C2(new_n717), .ZN(new_n929));
  OAI21_X1  g728(.A(new_n925), .B1(new_n927), .B2(new_n929), .ZN(G1354gat));
  OAI21_X1  g729(.A(G218gat), .B1(new_n917), .B2(new_n608), .ZN(new_n931));
  OR3_X1    g730(.A1(new_n911), .A2(G218gat), .A3(new_n608), .ZN(new_n932));
  NAND2_X1  g731(.A1(new_n931), .A2(new_n932), .ZN(G1355gat));
endmodule


