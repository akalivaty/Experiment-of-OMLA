//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 0 1 0 1 1 0 1 1 0 0 0 0 1 0 1 0 1 0 1 0 0 1 1 0 0 0 1 0 1 1 0 0 0 1 1 1 0 0 0 0 1 1 1 1 0 1 1 1 1 1 1 0 0 0 1 1 0 0 0 0 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:23:46 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n713, new_n714, new_n715, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n729, new_n731, new_n732, new_n733, new_n735,
    new_n736, new_n737, new_n738, new_n739, new_n740, new_n741, new_n742,
    new_n743, new_n744, new_n745, new_n746, new_n747, new_n748, new_n749,
    new_n751, new_n752, new_n753, new_n754, new_n755, new_n756, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n772, new_n773,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n806, new_n807, new_n808, new_n809, new_n810,
    new_n811, new_n812, new_n813, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n934, new_n935, new_n936, new_n937, new_n938,
    new_n939, new_n940, new_n941, new_n942, new_n943, new_n944, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n953, new_n954,
    new_n955, new_n957, new_n958, new_n959, new_n960, new_n961, new_n963,
    new_n964, new_n965, new_n966, new_n967, new_n968, new_n969, new_n970,
    new_n971, new_n972, new_n973, new_n974, new_n975, new_n976, new_n978,
    new_n979, new_n980, new_n981, new_n982, new_n983, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1021, new_n1022, new_n1023, new_n1024;
  INV_X1    g000(.A(KEYINPUT94), .ZN(new_n187));
  XNOR2_X1  g001(.A(KEYINPUT9), .B(G234), .ZN(new_n188));
  INV_X1    g002(.A(G217), .ZN(new_n189));
  NOR3_X1   g003(.A1(new_n188), .A2(new_n189), .A3(G953), .ZN(new_n190));
  INV_X1    g004(.A(new_n190), .ZN(new_n191));
  INV_X1    g005(.A(G107), .ZN(new_n192));
  INV_X1    g006(.A(KEYINPUT88), .ZN(new_n193));
  NOR2_X1   g007(.A1(new_n193), .A2(G122), .ZN(new_n194));
  INV_X1    g008(.A(G122), .ZN(new_n195));
  NOR2_X1   g009(.A1(new_n195), .A2(KEYINPUT88), .ZN(new_n196));
  OAI21_X1  g010(.A(G116), .B1(new_n194), .B2(new_n196), .ZN(new_n197));
  INV_X1    g011(.A(KEYINPUT90), .ZN(new_n198));
  INV_X1    g012(.A(KEYINPUT89), .ZN(new_n199));
  OAI21_X1  g013(.A(new_n199), .B1(new_n195), .B2(G116), .ZN(new_n200));
  INV_X1    g014(.A(G116), .ZN(new_n201));
  NAND3_X1  g015(.A1(new_n201), .A2(KEYINPUT89), .A3(G122), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n200), .A2(new_n202), .ZN(new_n203));
  AND3_X1   g017(.A1(new_n197), .A2(new_n198), .A3(new_n203), .ZN(new_n204));
  AOI21_X1  g018(.A(new_n198), .B1(new_n197), .B2(new_n203), .ZN(new_n205));
  OAI21_X1  g019(.A(new_n192), .B1(new_n204), .B2(new_n205), .ZN(new_n206));
  INV_X1    g020(.A(G143), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n207), .A2(G128), .ZN(new_n208));
  INV_X1    g022(.A(G128), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n209), .A2(G143), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n208), .A2(new_n210), .ZN(new_n211));
  XNOR2_X1  g025(.A(KEYINPUT91), .B(G134), .ZN(new_n212));
  XNOR2_X1  g026(.A(new_n211), .B(new_n212), .ZN(new_n213));
  INV_X1    g027(.A(new_n213), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n206), .A2(new_n214), .ZN(new_n215));
  INV_X1    g029(.A(KEYINPUT93), .ZN(new_n216));
  INV_X1    g030(.A(KEYINPUT14), .ZN(new_n217));
  NAND3_X1  g031(.A1(new_n200), .A2(new_n217), .A3(new_n202), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n197), .A2(new_n218), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n203), .A2(KEYINPUT14), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n220), .A2(KEYINPUT92), .ZN(new_n221));
  INV_X1    g035(.A(KEYINPUT92), .ZN(new_n222));
  NAND3_X1  g036(.A1(new_n203), .A2(new_n222), .A3(KEYINPUT14), .ZN(new_n223));
  AOI21_X1  g037(.A(new_n219), .B1(new_n221), .B2(new_n223), .ZN(new_n224));
  OAI21_X1  g038(.A(new_n216), .B1(new_n224), .B2(new_n192), .ZN(new_n225));
  AOI21_X1  g039(.A(new_n222), .B1(new_n203), .B2(KEYINPUT14), .ZN(new_n226));
  AOI211_X1 g040(.A(KEYINPUT92), .B(new_n217), .C1(new_n200), .C2(new_n202), .ZN(new_n227));
  OAI211_X1 g041(.A(new_n197), .B(new_n218), .C1(new_n226), .C2(new_n227), .ZN(new_n228));
  NAND3_X1  g042(.A1(new_n228), .A2(KEYINPUT93), .A3(G107), .ZN(new_n229));
  AOI21_X1  g043(.A(new_n215), .B1(new_n225), .B2(new_n229), .ZN(new_n230));
  INV_X1    g044(.A(G134), .ZN(new_n231));
  INV_X1    g045(.A(KEYINPUT13), .ZN(new_n232));
  AOI21_X1  g046(.A(new_n231), .B1(new_n210), .B2(new_n232), .ZN(new_n233));
  XNOR2_X1  g047(.A(new_n233), .B(new_n211), .ZN(new_n234));
  INV_X1    g048(.A(new_n205), .ZN(new_n235));
  NAND3_X1  g049(.A1(new_n197), .A2(new_n198), .A3(new_n203), .ZN(new_n236));
  NAND3_X1  g050(.A1(new_n235), .A2(G107), .A3(new_n236), .ZN(new_n237));
  AOI21_X1  g051(.A(new_n234), .B1(new_n237), .B2(new_n206), .ZN(new_n238));
  OAI21_X1  g052(.A(new_n191), .B1(new_n230), .B2(new_n238), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n235), .A2(new_n236), .ZN(new_n240));
  AOI21_X1  g054(.A(new_n213), .B1(new_n240), .B2(new_n192), .ZN(new_n241));
  NOR3_X1   g055(.A1(new_n224), .A2(new_n216), .A3(new_n192), .ZN(new_n242));
  AOI21_X1  g056(.A(KEYINPUT93), .B1(new_n228), .B2(G107), .ZN(new_n243));
  OAI21_X1  g057(.A(new_n241), .B1(new_n242), .B2(new_n243), .ZN(new_n244));
  INV_X1    g058(.A(new_n238), .ZN(new_n245));
  NAND3_X1  g059(.A1(new_n244), .A2(new_n245), .A3(new_n190), .ZN(new_n246));
  AOI21_X1  g060(.A(G902), .B1(new_n239), .B2(new_n246), .ZN(new_n247));
  INV_X1    g061(.A(G478), .ZN(new_n248));
  NOR2_X1   g062(.A1(new_n248), .A2(KEYINPUT15), .ZN(new_n249));
  INV_X1    g063(.A(new_n249), .ZN(new_n250));
  NOR2_X1   g064(.A1(new_n247), .A2(new_n250), .ZN(new_n251));
  AOI211_X1 g065(.A(G902), .B(new_n249), .C1(new_n239), .C2(new_n246), .ZN(new_n252));
  OAI21_X1  g066(.A(new_n187), .B1(new_n251), .B2(new_n252), .ZN(new_n253));
  INV_X1    g067(.A(G902), .ZN(new_n254));
  NOR3_X1   g068(.A1(new_n230), .A2(new_n238), .A3(new_n191), .ZN(new_n255));
  AOI21_X1  g069(.A(new_n190), .B1(new_n244), .B2(new_n245), .ZN(new_n256));
  OAI21_X1  g070(.A(new_n254), .B1(new_n255), .B2(new_n256), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n257), .A2(new_n249), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n247), .A2(new_n250), .ZN(new_n259));
  NAND3_X1  g073(.A1(new_n258), .A2(KEYINPUT94), .A3(new_n259), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n253), .A2(new_n260), .ZN(new_n261));
  INV_X1    g075(.A(G237), .ZN(new_n262));
  INV_X1    g076(.A(G953), .ZN(new_n263));
  NAND3_X1  g077(.A1(new_n262), .A2(new_n263), .A3(G214), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n264), .A2(new_n207), .ZN(new_n265));
  NOR2_X1   g079(.A1(G237), .A2(G953), .ZN(new_n266));
  NAND3_X1  g080(.A1(new_n266), .A2(G143), .A3(G214), .ZN(new_n267));
  NAND3_X1  g081(.A1(new_n265), .A2(KEYINPUT84), .A3(new_n267), .ZN(new_n268));
  NAND2_X1  g082(.A1(KEYINPUT18), .A2(G131), .ZN(new_n269));
  INV_X1    g083(.A(new_n269), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n268), .A2(new_n270), .ZN(new_n271));
  NAND4_X1  g085(.A1(new_n265), .A2(KEYINPUT84), .A3(new_n269), .A4(new_n267), .ZN(new_n272));
  INV_X1    g086(.A(G140), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n273), .A2(G125), .ZN(new_n274));
  INV_X1    g088(.A(G125), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n275), .A2(G140), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n274), .A2(new_n276), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n277), .A2(G146), .ZN(new_n278));
  INV_X1    g092(.A(G146), .ZN(new_n279));
  NAND3_X1  g093(.A1(new_n274), .A2(new_n276), .A3(new_n279), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n278), .A2(new_n280), .ZN(new_n281));
  NAND3_X1  g095(.A1(new_n271), .A2(new_n272), .A3(new_n281), .ZN(new_n282));
  XNOR2_X1  g096(.A(G113), .B(G122), .ZN(new_n283));
  XNOR2_X1  g097(.A(new_n283), .B(G104), .ZN(new_n284));
  XNOR2_X1  g098(.A(new_n284), .B(KEYINPUT86), .ZN(new_n285));
  NAND3_X1  g099(.A1(new_n274), .A2(new_n276), .A3(KEYINPUT16), .ZN(new_n286));
  OR3_X1    g100(.A1(new_n275), .A2(KEYINPUT16), .A3(G140), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n288), .A2(new_n279), .ZN(new_n289));
  NAND3_X1  g103(.A1(new_n286), .A2(new_n287), .A3(G146), .ZN(new_n290));
  NAND3_X1  g104(.A1(new_n289), .A2(KEYINPUT72), .A3(new_n290), .ZN(new_n291));
  INV_X1    g105(.A(KEYINPUT72), .ZN(new_n292));
  NAND3_X1  g106(.A1(new_n288), .A2(new_n292), .A3(new_n279), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n291), .A2(new_n293), .ZN(new_n294));
  INV_X1    g108(.A(new_n294), .ZN(new_n295));
  INV_X1    g109(.A(new_n267), .ZN(new_n296));
  AOI21_X1  g110(.A(G143), .B1(new_n266), .B2(G214), .ZN(new_n297));
  OAI21_X1  g111(.A(G131), .B1(new_n296), .B2(new_n297), .ZN(new_n298));
  INV_X1    g112(.A(KEYINPUT17), .ZN(new_n299));
  INV_X1    g113(.A(G131), .ZN(new_n300));
  NAND3_X1  g114(.A1(new_n265), .A2(new_n300), .A3(new_n267), .ZN(new_n301));
  NAND3_X1  g115(.A1(new_n298), .A2(new_n299), .A3(new_n301), .ZN(new_n302));
  AOI21_X1  g116(.A(new_n300), .B1(new_n265), .B2(new_n267), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n303), .A2(KEYINPUT17), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n302), .A2(new_n304), .ZN(new_n305));
  OAI211_X1 g119(.A(new_n282), .B(new_n285), .C1(new_n295), .C2(new_n305), .ZN(new_n306));
  INV_X1    g120(.A(new_n284), .ZN(new_n307));
  INV_X1    g121(.A(new_n282), .ZN(new_n308));
  AND2_X1   g122(.A1(new_n302), .A2(new_n304), .ZN(new_n309));
  AOI21_X1  g123(.A(new_n308), .B1(new_n309), .B2(new_n294), .ZN(new_n310));
  OAI21_X1  g124(.A(new_n306), .B1(new_n307), .B2(new_n310), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n311), .A2(new_n254), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n312), .A2(G475), .ZN(new_n313));
  AND3_X1   g127(.A1(new_n274), .A2(new_n276), .A3(KEYINPUT19), .ZN(new_n314));
  AOI21_X1  g128(.A(KEYINPUT19), .B1(new_n274), .B2(new_n276), .ZN(new_n315));
  OAI21_X1  g129(.A(new_n279), .B1(new_n314), .B2(new_n315), .ZN(new_n316));
  NOR3_X1   g130(.A1(new_n296), .A2(new_n297), .A3(G131), .ZN(new_n317));
  OAI211_X1 g131(.A(new_n316), .B(new_n290), .C1(new_n317), .C2(new_n303), .ZN(new_n318));
  INV_X1    g132(.A(KEYINPUT85), .ZN(new_n319));
  NAND3_X1  g133(.A1(new_n318), .A2(new_n282), .A3(new_n319), .ZN(new_n320));
  AND2_X1   g134(.A1(new_n320), .A2(new_n284), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n318), .A2(new_n282), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n322), .A2(KEYINPUT85), .ZN(new_n323));
  AOI22_X1  g137(.A1(new_n321), .A2(new_n323), .B1(new_n310), .B2(new_n285), .ZN(new_n324));
  NOR2_X1   g138(.A1(G475), .A2(G902), .ZN(new_n325));
  INV_X1    g139(.A(new_n325), .ZN(new_n326));
  OAI21_X1  g140(.A(KEYINPUT20), .B1(new_n324), .B2(new_n326), .ZN(new_n327));
  NAND3_X1  g141(.A1(new_n323), .A2(new_n284), .A3(new_n320), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n328), .A2(new_n306), .ZN(new_n329));
  INV_X1    g143(.A(KEYINPUT20), .ZN(new_n330));
  NAND4_X1  g144(.A1(new_n329), .A2(KEYINPUT87), .A3(new_n330), .A4(new_n325), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n327), .A2(new_n331), .ZN(new_n332));
  AOI21_X1  g146(.A(new_n326), .B1(new_n328), .B2(new_n306), .ZN(new_n333));
  AOI21_X1  g147(.A(KEYINPUT87), .B1(new_n333), .B2(new_n330), .ZN(new_n334));
  OAI21_X1  g148(.A(new_n313), .B1(new_n332), .B2(new_n334), .ZN(new_n335));
  INV_X1    g149(.A(new_n335), .ZN(new_n336));
  NAND2_X1  g150(.A1(G234), .A2(G237), .ZN(new_n337));
  NAND3_X1  g151(.A1(new_n337), .A2(G952), .A3(new_n263), .ZN(new_n338));
  INV_X1    g152(.A(new_n338), .ZN(new_n339));
  NAND3_X1  g153(.A1(new_n337), .A2(G902), .A3(G953), .ZN(new_n340));
  INV_X1    g154(.A(new_n340), .ZN(new_n341));
  XNOR2_X1  g155(.A(KEYINPUT21), .B(G898), .ZN(new_n342));
  AOI21_X1  g156(.A(new_n339), .B1(new_n341), .B2(new_n342), .ZN(new_n343));
  INV_X1    g157(.A(new_n343), .ZN(new_n344));
  NAND3_X1  g158(.A1(new_n261), .A2(new_n336), .A3(new_n344), .ZN(new_n345));
  INV_X1    g159(.A(G469), .ZN(new_n346));
  INV_X1    g160(.A(G104), .ZN(new_n347));
  OAI21_X1  g161(.A(KEYINPUT3), .B1(new_n347), .B2(G107), .ZN(new_n348));
  INV_X1    g162(.A(KEYINPUT74), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n348), .A2(new_n349), .ZN(new_n350));
  OAI211_X1 g164(.A(KEYINPUT74), .B(KEYINPUT3), .C1(new_n347), .C2(G107), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  INV_X1    g166(.A(KEYINPUT3), .ZN(new_n353));
  NAND3_X1  g167(.A1(new_n353), .A2(new_n192), .A3(G104), .ZN(new_n354));
  INV_X1    g168(.A(KEYINPUT75), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  NAND4_X1  g170(.A1(new_n353), .A2(new_n192), .A3(KEYINPUT75), .A4(G104), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  INV_X1    g172(.A(G101), .ZN(new_n359));
  NOR2_X1   g173(.A1(new_n192), .A2(G104), .ZN(new_n360));
  INV_X1    g174(.A(new_n360), .ZN(new_n361));
  NAND4_X1  g175(.A1(new_n352), .A2(new_n358), .A3(new_n359), .A4(new_n361), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n192), .A2(G104), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n361), .A2(new_n363), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n364), .A2(G101), .ZN(new_n365));
  AND2_X1   g179(.A1(new_n362), .A2(new_n365), .ZN(new_n366));
  INV_X1    g180(.A(KEYINPUT10), .ZN(new_n367));
  INV_X1    g181(.A(KEYINPUT1), .ZN(new_n368));
  AOI21_X1  g182(.A(new_n368), .B1(G143), .B2(new_n279), .ZN(new_n369));
  NOR2_X1   g183(.A1(new_n207), .A2(G146), .ZN(new_n370));
  NOR2_X1   g184(.A1(new_n279), .A2(G143), .ZN(new_n371));
  OAI22_X1  g185(.A1(new_n369), .A2(new_n209), .B1(new_n370), .B2(new_n371), .ZN(new_n372));
  OAI21_X1  g186(.A(KEYINPUT64), .B1(new_n207), .B2(G146), .ZN(new_n373));
  INV_X1    g187(.A(KEYINPUT64), .ZN(new_n374));
  NAND3_X1  g188(.A1(new_n374), .A2(new_n279), .A3(G143), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n207), .A2(G146), .ZN(new_n376));
  NOR2_X1   g190(.A1(new_n209), .A2(KEYINPUT1), .ZN(new_n377));
  NAND4_X1  g191(.A1(new_n373), .A2(new_n375), .A3(new_n376), .A4(new_n377), .ZN(new_n378));
  AOI21_X1  g192(.A(new_n367), .B1(new_n372), .B2(new_n378), .ZN(new_n379));
  AND3_X1   g193(.A1(new_n373), .A2(new_n375), .A3(new_n376), .ZN(new_n380));
  NOR2_X1   g194(.A1(new_n369), .A2(new_n209), .ZN(new_n381));
  OAI21_X1  g195(.A(new_n378), .B1(new_n380), .B2(new_n381), .ZN(new_n382));
  NAND3_X1  g196(.A1(new_n362), .A2(new_n365), .A3(new_n382), .ZN(new_n383));
  AOI22_X1  g197(.A1(new_n366), .A2(new_n379), .B1(new_n383), .B2(new_n367), .ZN(new_n384));
  INV_X1    g198(.A(new_n351), .ZN(new_n385));
  AOI21_X1  g199(.A(KEYINPUT74), .B1(new_n363), .B2(KEYINPUT3), .ZN(new_n386));
  OAI21_X1  g200(.A(new_n361), .B1(new_n385), .B2(new_n386), .ZN(new_n387));
  AND2_X1   g201(.A1(new_n356), .A2(new_n357), .ZN(new_n388));
  OAI21_X1  g202(.A(G101), .B1(new_n387), .B2(new_n388), .ZN(new_n389));
  NAND3_X1  g203(.A1(new_n389), .A2(KEYINPUT4), .A3(new_n362), .ZN(new_n390));
  NAND2_X1  g204(.A1(KEYINPUT0), .A2(G128), .ZN(new_n391));
  OR2_X1    g205(.A1(KEYINPUT0), .A2(G128), .ZN(new_n392));
  OAI211_X1 g206(.A(new_n391), .B(new_n392), .C1(new_n370), .C2(new_n371), .ZN(new_n393));
  INV_X1    g207(.A(new_n391), .ZN(new_n394));
  NAND4_X1  g208(.A1(new_n373), .A2(new_n375), .A3(new_n394), .A4(new_n376), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n393), .A2(new_n395), .ZN(new_n396));
  AOI21_X1  g210(.A(new_n360), .B1(new_n350), .B2(new_n351), .ZN(new_n397));
  AOI21_X1  g211(.A(new_n359), .B1(new_n397), .B2(new_n358), .ZN(new_n398));
  INV_X1    g212(.A(KEYINPUT4), .ZN(new_n399));
  AOI21_X1  g213(.A(new_n396), .B1(new_n398), .B2(new_n399), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n390), .A2(new_n400), .ZN(new_n401));
  INV_X1    g215(.A(KEYINPUT11), .ZN(new_n402));
  NOR2_X1   g216(.A1(new_n402), .A2(KEYINPUT65), .ZN(new_n403));
  NOR2_X1   g217(.A1(new_n231), .A2(G137), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n402), .A2(KEYINPUT65), .ZN(new_n405));
  AOI21_X1  g219(.A(new_n403), .B1(new_n404), .B2(new_n405), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n231), .A2(G137), .ZN(new_n407));
  INV_X1    g221(.A(KEYINPUT65), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n408), .A2(KEYINPUT11), .ZN(new_n409));
  INV_X1    g223(.A(G137), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n410), .A2(G134), .ZN(new_n411));
  OAI21_X1  g225(.A(new_n407), .B1(new_n409), .B2(new_n411), .ZN(new_n412));
  NOR3_X1   g226(.A1(new_n406), .A2(new_n412), .A3(G131), .ZN(new_n413));
  NOR2_X1   g227(.A1(new_n410), .A2(G134), .ZN(new_n414));
  AOI21_X1  g228(.A(new_n414), .B1(new_n403), .B2(new_n404), .ZN(new_n415));
  NOR2_X1   g229(.A1(new_n408), .A2(KEYINPUT11), .ZN(new_n416));
  OAI21_X1  g230(.A(new_n409), .B1(new_n416), .B2(new_n411), .ZN(new_n417));
  AOI21_X1  g231(.A(new_n300), .B1(new_n415), .B2(new_n417), .ZN(new_n418));
  NOR2_X1   g232(.A1(new_n413), .A2(new_n418), .ZN(new_n419));
  NAND3_X1  g233(.A1(new_n384), .A2(new_n401), .A3(new_n419), .ZN(new_n420));
  NOR2_X1   g234(.A1(new_n419), .A2(KEYINPUT76), .ZN(new_n421));
  INV_X1    g235(.A(new_n383), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n372), .A2(new_n378), .ZN(new_n423));
  AOI21_X1  g237(.A(new_n423), .B1(new_n362), .B2(new_n365), .ZN(new_n424));
  OAI21_X1  g238(.A(new_n421), .B1(new_n422), .B2(new_n424), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n425), .A2(KEYINPUT12), .ZN(new_n426));
  INV_X1    g240(.A(KEYINPUT12), .ZN(new_n427));
  OAI211_X1 g241(.A(new_n421), .B(new_n427), .C1(new_n422), .C2(new_n424), .ZN(new_n428));
  XNOR2_X1  g242(.A(G110), .B(G140), .ZN(new_n429));
  AND2_X1   g243(.A1(new_n263), .A2(G227), .ZN(new_n430));
  XNOR2_X1  g244(.A(new_n429), .B(new_n430), .ZN(new_n431));
  INV_X1    g245(.A(new_n431), .ZN(new_n432));
  NAND4_X1  g246(.A1(new_n420), .A2(new_n426), .A3(new_n428), .A4(new_n432), .ZN(new_n433));
  INV_X1    g247(.A(new_n433), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n384), .A2(new_n401), .ZN(new_n435));
  INV_X1    g249(.A(new_n419), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n435), .A2(new_n436), .ZN(new_n437));
  AOI21_X1  g251(.A(new_n432), .B1(new_n437), .B2(new_n420), .ZN(new_n438));
  OAI211_X1 g252(.A(new_n346), .B(new_n254), .C1(new_n434), .C2(new_n438), .ZN(new_n439));
  NOR2_X1   g253(.A1(new_n346), .A2(new_n254), .ZN(new_n440));
  INV_X1    g254(.A(new_n440), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n426), .A2(new_n428), .ZN(new_n442));
  INV_X1    g256(.A(new_n420), .ZN(new_n443));
  OAI21_X1  g257(.A(new_n431), .B1(new_n442), .B2(new_n443), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n420), .A2(new_n432), .ZN(new_n445));
  INV_X1    g259(.A(KEYINPUT77), .ZN(new_n446));
  OAI21_X1  g260(.A(new_n437), .B1(new_n445), .B2(new_n446), .ZN(new_n447));
  AOI21_X1  g261(.A(KEYINPUT77), .B1(new_n420), .B2(new_n432), .ZN(new_n448));
  OAI21_X1  g262(.A(new_n444), .B1(new_n447), .B2(new_n448), .ZN(new_n449));
  OAI211_X1 g263(.A(new_n439), .B(new_n441), .C1(new_n449), .C2(new_n346), .ZN(new_n450));
  OAI21_X1  g264(.A(G221), .B1(new_n188), .B2(G902), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  NOR2_X1   g266(.A1(new_n345), .A2(new_n452), .ZN(new_n453));
  XOR2_X1   g267(.A(G119), .B(G128), .Z(new_n454));
  XNOR2_X1  g268(.A(KEYINPUT24), .B(G110), .ZN(new_n455));
  NOR2_X1   g269(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  INV_X1    g270(.A(KEYINPUT23), .ZN(new_n457));
  INV_X1    g271(.A(G119), .ZN(new_n458));
  OAI21_X1  g272(.A(new_n457), .B1(new_n458), .B2(G128), .ZN(new_n459));
  NAND3_X1  g273(.A1(new_n209), .A2(KEYINPUT23), .A3(G119), .ZN(new_n460));
  OAI211_X1 g274(.A(new_n459), .B(new_n460), .C1(G119), .C2(new_n209), .ZN(new_n461));
  AOI21_X1  g275(.A(new_n456), .B1(G110), .B2(new_n461), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n295), .A2(new_n462), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n454), .A2(new_n455), .ZN(new_n464));
  OAI21_X1  g278(.A(new_n464), .B1(new_n461), .B2(G110), .ZN(new_n465));
  AND2_X1   g279(.A1(new_n465), .A2(KEYINPUT73), .ZN(new_n466));
  NOR2_X1   g280(.A1(new_n465), .A2(KEYINPUT73), .ZN(new_n467));
  OAI211_X1 g281(.A(new_n290), .B(new_n280), .C1(new_n466), .C2(new_n467), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n463), .A2(new_n468), .ZN(new_n469));
  XNOR2_X1  g283(.A(KEYINPUT22), .B(G137), .ZN(new_n470));
  NAND3_X1  g284(.A1(new_n263), .A2(G221), .A3(G234), .ZN(new_n471));
  XNOR2_X1  g285(.A(new_n470), .B(new_n471), .ZN(new_n472));
  INV_X1    g286(.A(new_n472), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n469), .A2(new_n473), .ZN(new_n474));
  NAND3_X1  g288(.A1(new_n463), .A2(new_n468), .A3(new_n472), .ZN(new_n475));
  NAND3_X1  g289(.A1(new_n474), .A2(new_n254), .A3(new_n475), .ZN(new_n476));
  INV_X1    g290(.A(KEYINPUT25), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  NAND4_X1  g292(.A1(new_n474), .A2(KEYINPUT25), .A3(new_n254), .A4(new_n475), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  AOI21_X1  g294(.A(new_n189), .B1(G234), .B2(new_n254), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  AND2_X1   g296(.A1(new_n474), .A2(new_n475), .ZN(new_n483));
  NOR2_X1   g297(.A1(new_n481), .A2(G902), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n482), .A2(new_n485), .ZN(new_n486));
  INV_X1    g300(.A(KEYINPUT28), .ZN(new_n487));
  INV_X1    g301(.A(KEYINPUT67), .ZN(new_n488));
  OAI21_X1  g302(.A(new_n488), .B1(new_n201), .B2(G119), .ZN(new_n489));
  NAND3_X1  g303(.A1(new_n458), .A2(KEYINPUT67), .A3(G116), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n201), .A2(G119), .ZN(new_n491));
  AND3_X1   g305(.A1(new_n489), .A2(new_n490), .A3(new_n491), .ZN(new_n492));
  XOR2_X1   g306(.A(KEYINPUT2), .B(G113), .Z(new_n493));
  XNOR2_X1  g307(.A(new_n492), .B(new_n493), .ZN(new_n494));
  NAND3_X1  g308(.A1(new_n415), .A2(new_n300), .A3(new_n417), .ZN(new_n495));
  OAI21_X1  g309(.A(G131), .B1(new_n404), .B2(new_n414), .ZN(new_n496));
  AND3_X1   g310(.A1(new_n423), .A2(new_n495), .A3(new_n496), .ZN(new_n497));
  OAI21_X1  g311(.A(G131), .B1(new_n406), .B2(new_n412), .ZN(new_n498));
  AOI21_X1  g312(.A(new_n396), .B1(new_n498), .B2(new_n495), .ZN(new_n499));
  OAI21_X1  g313(.A(new_n494), .B1(new_n497), .B2(new_n499), .ZN(new_n500));
  INV_X1    g314(.A(new_n396), .ZN(new_n501));
  OAI21_X1  g315(.A(new_n501), .B1(new_n413), .B2(new_n418), .ZN(new_n502));
  NAND3_X1  g316(.A1(new_n489), .A2(new_n490), .A3(new_n491), .ZN(new_n503));
  XNOR2_X1  g317(.A(new_n503), .B(new_n493), .ZN(new_n504));
  NAND3_X1  g318(.A1(new_n423), .A2(new_n495), .A3(new_n496), .ZN(new_n505));
  NAND3_X1  g319(.A1(new_n502), .A2(new_n504), .A3(new_n505), .ZN(new_n506));
  AOI21_X1  g320(.A(new_n487), .B1(new_n500), .B2(new_n506), .ZN(new_n507));
  NOR2_X1   g321(.A1(new_n497), .A2(new_n499), .ZN(new_n508));
  AOI21_X1  g322(.A(KEYINPUT28), .B1(new_n508), .B2(new_n504), .ZN(new_n509));
  XOR2_X1   g323(.A(KEYINPUT26), .B(G101), .Z(new_n510));
  NAND2_X1  g324(.A1(new_n266), .A2(G210), .ZN(new_n511));
  XNOR2_X1  g325(.A(new_n510), .B(new_n511), .ZN(new_n512));
  XNOR2_X1  g326(.A(KEYINPUT68), .B(KEYINPUT27), .ZN(new_n513));
  AND2_X1   g327(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  NOR2_X1   g328(.A1(new_n512), .A2(new_n513), .ZN(new_n515));
  OAI21_X1  g329(.A(KEYINPUT29), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  NOR3_X1   g330(.A1(new_n507), .A2(new_n509), .A3(new_n516), .ZN(new_n517));
  OAI21_X1  g331(.A(KEYINPUT70), .B1(new_n517), .B2(G902), .ZN(new_n518));
  NOR2_X1   g332(.A1(new_n514), .A2(new_n515), .ZN(new_n519));
  NAND2_X1  g333(.A1(KEYINPUT66), .A2(KEYINPUT30), .ZN(new_n520));
  INV_X1    g334(.A(KEYINPUT66), .ZN(new_n521));
  INV_X1    g335(.A(KEYINPUT30), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  OAI211_X1 g337(.A(new_n520), .B(new_n523), .C1(new_n497), .C2(new_n499), .ZN(new_n524));
  NAND4_X1  g338(.A1(new_n502), .A2(new_n521), .A3(new_n522), .A4(new_n505), .ZN(new_n525));
  AOI21_X1  g339(.A(new_n504), .B1(new_n524), .B2(new_n525), .ZN(new_n526));
  NOR3_X1   g340(.A1(new_n497), .A2(new_n499), .A3(new_n494), .ZN(new_n527));
  OAI21_X1  g341(.A(new_n519), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  XNOR2_X1  g342(.A(KEYINPUT69), .B(KEYINPUT28), .ZN(new_n529));
  AOI21_X1  g343(.A(new_n504), .B1(new_n502), .B2(new_n505), .ZN(new_n530));
  OAI21_X1  g344(.A(new_n529), .B1(new_n527), .B2(new_n530), .ZN(new_n531));
  INV_X1    g345(.A(new_n519), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n506), .A2(new_n487), .ZN(new_n533));
  NAND3_X1  g347(.A1(new_n531), .A2(new_n532), .A3(new_n533), .ZN(new_n534));
  INV_X1    g348(.A(KEYINPUT29), .ZN(new_n535));
  NAND3_X1  g349(.A1(new_n528), .A2(new_n534), .A3(new_n535), .ZN(new_n536));
  OAI21_X1  g350(.A(KEYINPUT28), .B1(new_n527), .B2(new_n530), .ZN(new_n537));
  INV_X1    g351(.A(new_n516), .ZN(new_n538));
  NAND3_X1  g352(.A1(new_n537), .A2(new_n533), .A3(new_n538), .ZN(new_n539));
  INV_X1    g353(.A(KEYINPUT70), .ZN(new_n540));
  NAND3_X1  g354(.A1(new_n539), .A2(new_n540), .A3(new_n254), .ZN(new_n541));
  NAND3_X1  g355(.A1(new_n518), .A2(new_n536), .A3(new_n541), .ZN(new_n542));
  INV_X1    g356(.A(KEYINPUT71), .ZN(new_n543));
  AND3_X1   g357(.A1(new_n542), .A2(new_n543), .A3(G472), .ZN(new_n544));
  AOI21_X1  g358(.A(new_n543), .B1(new_n542), .B2(G472), .ZN(new_n545));
  NOR2_X1   g359(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  AOI21_X1  g360(.A(new_n532), .B1(new_n531), .B2(new_n533), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n524), .A2(new_n525), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n548), .A2(new_n494), .ZN(new_n549));
  NAND3_X1  g363(.A1(new_n549), .A2(new_n532), .A3(new_n506), .ZN(new_n550));
  INV_X1    g364(.A(KEYINPUT31), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  AOI21_X1  g366(.A(new_n527), .B1(new_n548), .B2(new_n494), .ZN(new_n553));
  NAND3_X1  g367(.A1(new_n553), .A2(KEYINPUT31), .A3(new_n532), .ZN(new_n554));
  AOI21_X1  g368(.A(new_n547), .B1(new_n552), .B2(new_n554), .ZN(new_n555));
  NOR2_X1   g369(.A1(G472), .A2(G902), .ZN(new_n556));
  INV_X1    g370(.A(new_n556), .ZN(new_n557));
  OAI21_X1  g371(.A(KEYINPUT32), .B1(new_n555), .B2(new_n557), .ZN(new_n558));
  INV_X1    g372(.A(new_n547), .ZN(new_n559));
  AOI21_X1  g373(.A(KEYINPUT31), .B1(new_n553), .B2(new_n532), .ZN(new_n560));
  NOR4_X1   g374(.A1(new_n526), .A2(new_n551), .A3(new_n519), .A4(new_n527), .ZN(new_n561));
  OAI21_X1  g375(.A(new_n559), .B1(new_n560), .B2(new_n561), .ZN(new_n562));
  INV_X1    g376(.A(KEYINPUT32), .ZN(new_n563));
  NAND3_X1  g377(.A1(new_n562), .A2(new_n563), .A3(new_n556), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n558), .A2(new_n564), .ZN(new_n565));
  AOI21_X1  g379(.A(new_n486), .B1(new_n546), .B2(new_n565), .ZN(new_n566));
  OAI21_X1  g380(.A(G214), .B1(G237), .B2(G902), .ZN(new_n567));
  OAI21_X1  g381(.A(G210), .B1(G237), .B2(G902), .ZN(new_n568));
  XNOR2_X1  g382(.A(new_n568), .B(KEYINPUT81), .ZN(new_n569));
  INV_X1    g383(.A(new_n569), .ZN(new_n570));
  MUX2_X1   g384(.A(new_n423), .B(new_n501), .S(G125), .Z(new_n571));
  INV_X1    g385(.A(G224), .ZN(new_n572));
  OAI21_X1  g386(.A(KEYINPUT7), .B1(new_n572), .B2(G953), .ZN(new_n573));
  XNOR2_X1  g387(.A(new_n571), .B(new_n573), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n492), .A2(KEYINPUT5), .ZN(new_n575));
  NOR3_X1   g389(.A1(new_n201), .A2(KEYINPUT5), .A3(G119), .ZN(new_n576));
  INV_X1    g390(.A(G113), .ZN(new_n577));
  NOR2_X1   g391(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  AOI22_X1  g392(.A1(new_n575), .A2(new_n578), .B1(new_n493), .B2(new_n492), .ZN(new_n579));
  XOR2_X1   g393(.A(new_n366), .B(new_n579), .Z(new_n580));
  XNOR2_X1  g394(.A(G110), .B(G122), .ZN(new_n581));
  XOR2_X1   g395(.A(new_n581), .B(KEYINPUT8), .Z(new_n582));
  OAI21_X1  g396(.A(new_n574), .B1(new_n580), .B2(new_n582), .ZN(new_n583));
  AOI21_X1  g397(.A(new_n504), .B1(new_n398), .B2(new_n399), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n584), .A2(new_n390), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n366), .A2(new_n579), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  INV_X1    g401(.A(new_n581), .ZN(new_n588));
  NOR2_X1   g402(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  OAI21_X1  g403(.A(new_n254), .B1(new_n583), .B2(new_n589), .ZN(new_n590));
  INV_X1    g404(.A(new_n590), .ZN(new_n591));
  INV_X1    g405(.A(KEYINPUT80), .ZN(new_n592));
  INV_X1    g406(.A(KEYINPUT78), .ZN(new_n593));
  NOR2_X1   g407(.A1(new_n581), .A2(KEYINPUT6), .ZN(new_n594));
  NAND3_X1  g408(.A1(new_n587), .A2(new_n593), .A3(new_n594), .ZN(new_n595));
  AOI22_X1  g409(.A1(new_n584), .A2(new_n390), .B1(new_n366), .B2(new_n579), .ZN(new_n596));
  INV_X1    g410(.A(new_n594), .ZN(new_n597));
  OAI21_X1  g411(.A(KEYINPUT78), .B1(new_n596), .B2(new_n597), .ZN(new_n598));
  INV_X1    g412(.A(KEYINPUT6), .ZN(new_n599));
  AOI21_X1  g413(.A(new_n599), .B1(new_n596), .B2(new_n581), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n587), .A2(new_n588), .ZN(new_n601));
  AOI22_X1  g415(.A1(new_n595), .A2(new_n598), .B1(new_n600), .B2(new_n601), .ZN(new_n602));
  NOR2_X1   g416(.A1(new_n572), .A2(G953), .ZN(new_n603));
  XNOR2_X1  g417(.A(new_n603), .B(KEYINPUT79), .ZN(new_n604));
  XNOR2_X1  g418(.A(new_n571), .B(new_n604), .ZN(new_n605));
  AOI21_X1  g419(.A(new_n592), .B1(new_n602), .B2(new_n605), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n595), .A2(new_n598), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n600), .A2(new_n601), .ZN(new_n608));
  AND4_X1   g422(.A1(new_n592), .A2(new_n607), .A3(new_n608), .A4(new_n605), .ZN(new_n609));
  OAI211_X1 g423(.A(new_n570), .B(new_n591), .C1(new_n606), .C2(new_n609), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n610), .A2(KEYINPUT83), .ZN(new_n611));
  NAND3_X1  g425(.A1(new_n607), .A2(new_n608), .A3(new_n605), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n612), .A2(KEYINPUT80), .ZN(new_n613));
  NAND3_X1  g427(.A1(new_n602), .A2(new_n592), .A3(new_n605), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  INV_X1    g429(.A(KEYINPUT83), .ZN(new_n616));
  NAND4_X1  g430(.A1(new_n615), .A2(new_n616), .A3(new_n570), .A4(new_n591), .ZN(new_n617));
  OAI21_X1  g431(.A(new_n591), .B1(new_n606), .B2(new_n609), .ZN(new_n618));
  XNOR2_X1  g432(.A(new_n569), .B(KEYINPUT82), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  NAND3_X1  g434(.A1(new_n611), .A2(new_n617), .A3(new_n620), .ZN(new_n621));
  NAND4_X1  g435(.A1(new_n453), .A2(new_n566), .A3(new_n567), .A4(new_n621), .ZN(new_n622));
  XNOR2_X1  g436(.A(new_n622), .B(G101), .ZN(G3));
  INV_X1    g437(.A(new_n481), .ZN(new_n624));
  AOI21_X1  g438(.A(new_n624), .B1(new_n478), .B2(new_n479), .ZN(new_n625));
  AOI21_X1  g439(.A(new_n625), .B1(new_n483), .B2(new_n484), .ZN(new_n626));
  NOR2_X1   g440(.A1(new_n555), .A2(new_n557), .ZN(new_n627));
  INV_X1    g441(.A(new_n627), .ZN(new_n628));
  OAI21_X1  g442(.A(G472), .B1(new_n555), .B2(G902), .ZN(new_n629));
  NAND3_X1  g443(.A1(new_n626), .A2(new_n628), .A3(new_n629), .ZN(new_n630));
  NOR2_X1   g444(.A1(new_n630), .A2(new_n452), .ZN(new_n631));
  INV_X1    g445(.A(new_n567), .ZN(new_n632));
  NAND2_X1  g446(.A1(new_n618), .A2(new_n569), .ZN(new_n633));
  AOI21_X1  g447(.A(new_n632), .B1(new_n633), .B2(new_n610), .ZN(new_n634));
  OAI21_X1  g448(.A(KEYINPUT33), .B1(new_n190), .B2(KEYINPUT95), .ZN(new_n635));
  NOR3_X1   g449(.A1(new_n255), .A2(new_n256), .A3(new_n635), .ZN(new_n636));
  INV_X1    g450(.A(new_n635), .ZN(new_n637));
  AOI21_X1  g451(.A(new_n637), .B1(new_n239), .B2(new_n246), .ZN(new_n638));
  OAI21_X1  g452(.A(G478), .B1(new_n636), .B2(new_n638), .ZN(new_n639));
  NOR2_X1   g453(.A1(new_n248), .A2(new_n254), .ZN(new_n640));
  AOI21_X1  g454(.A(new_n640), .B1(new_n247), .B2(new_n248), .ZN(new_n641));
  AND4_X1   g455(.A1(new_n335), .A2(new_n344), .A3(new_n639), .A4(new_n641), .ZN(new_n642));
  NAND3_X1  g456(.A1(new_n631), .A2(new_n634), .A3(new_n642), .ZN(new_n643));
  XNOR2_X1  g457(.A(new_n643), .B(KEYINPUT96), .ZN(new_n644));
  XNOR2_X1  g458(.A(KEYINPUT34), .B(G104), .ZN(new_n645));
  XNOR2_X1  g459(.A(new_n644), .B(new_n645), .ZN(G6));
  XNOR2_X1  g460(.A(new_n343), .B(KEYINPUT98), .ZN(new_n647));
  INV_X1    g461(.A(new_n647), .ZN(new_n648));
  AOI211_X1 g462(.A(new_n632), .B(new_n648), .C1(new_n633), .C2(new_n610), .ZN(new_n649));
  AND2_X1   g463(.A1(new_n312), .A2(G475), .ZN(new_n650));
  INV_X1    g464(.A(KEYINPUT97), .ZN(new_n651));
  AOI21_X1  g465(.A(new_n330), .B1(new_n329), .B2(new_n325), .ZN(new_n652));
  AOI211_X1 g466(.A(KEYINPUT20), .B(new_n326), .C1(new_n328), .C2(new_n306), .ZN(new_n653));
  OAI21_X1  g467(.A(new_n651), .B1(new_n652), .B2(new_n653), .ZN(new_n654));
  NAND2_X1  g468(.A1(new_n333), .A2(new_n330), .ZN(new_n655));
  NAND3_X1  g469(.A1(new_n327), .A2(new_n655), .A3(KEYINPUT97), .ZN(new_n656));
  AOI21_X1  g470(.A(new_n650), .B1(new_n654), .B2(new_n656), .ZN(new_n657));
  NAND3_X1  g471(.A1(new_n657), .A2(new_n253), .A3(new_n260), .ZN(new_n658));
  INV_X1    g472(.A(new_n658), .ZN(new_n659));
  NAND3_X1  g473(.A1(new_n649), .A2(new_n631), .A3(new_n659), .ZN(new_n660));
  XOR2_X1   g474(.A(KEYINPUT35), .B(G107), .Z(new_n661));
  XNOR2_X1  g475(.A(new_n660), .B(new_n661), .ZN(G9));
  NOR2_X1   g476(.A1(new_n473), .A2(KEYINPUT36), .ZN(new_n663));
  XNOR2_X1  g477(.A(new_n663), .B(KEYINPUT99), .ZN(new_n664));
  XNOR2_X1  g478(.A(new_n469), .B(new_n664), .ZN(new_n665));
  AOI21_X1  g479(.A(new_n625), .B1(new_n484), .B2(new_n665), .ZN(new_n666));
  INV_X1    g480(.A(G472), .ZN(new_n667));
  AOI21_X1  g481(.A(new_n667), .B1(new_n562), .B2(new_n254), .ZN(new_n668));
  NOR3_X1   g482(.A1(new_n666), .A2(new_n627), .A3(new_n668), .ZN(new_n669));
  NAND4_X1  g483(.A1(new_n453), .A2(new_n621), .A3(new_n567), .A4(new_n669), .ZN(new_n670));
  XOR2_X1   g484(.A(KEYINPUT37), .B(G110), .Z(new_n671));
  XNOR2_X1  g485(.A(new_n670), .B(new_n671), .ZN(G12));
  NAND2_X1  g486(.A1(new_n542), .A2(G472), .ZN(new_n673));
  NAND2_X1  g487(.A1(new_n673), .A2(KEYINPUT71), .ZN(new_n674));
  NAND3_X1  g488(.A1(new_n542), .A2(new_n543), .A3(G472), .ZN(new_n675));
  AOI21_X1  g489(.A(new_n563), .B1(new_n562), .B2(new_n556), .ZN(new_n676));
  AND3_X1   g490(.A1(new_n562), .A2(new_n563), .A3(new_n556), .ZN(new_n677));
  OAI211_X1 g491(.A(new_n674), .B(new_n675), .C1(new_n676), .C2(new_n677), .ZN(new_n678));
  NAND2_X1  g492(.A1(new_n665), .A2(new_n484), .ZN(new_n679));
  NAND2_X1  g493(.A1(new_n482), .A2(new_n679), .ZN(new_n680));
  AND3_X1   g494(.A1(new_n680), .A2(new_n450), .A3(new_n451), .ZN(new_n681));
  OR2_X1    g495(.A1(new_n340), .A2(G900), .ZN(new_n682));
  NAND2_X1  g496(.A1(new_n682), .A2(new_n338), .ZN(new_n683));
  AND4_X1   g497(.A1(new_n260), .A2(new_n657), .A3(new_n253), .A4(new_n683), .ZN(new_n684));
  NAND4_X1  g498(.A1(new_n634), .A2(new_n678), .A3(new_n681), .A4(new_n684), .ZN(new_n685));
  XNOR2_X1  g499(.A(new_n685), .B(G128), .ZN(G30));
  INV_X1    g500(.A(KEYINPUT38), .ZN(new_n687));
  XNOR2_X1  g501(.A(new_n621), .B(new_n687), .ZN(new_n688));
  INV_X1    g502(.A(new_n553), .ZN(new_n689));
  NAND2_X1  g503(.A1(new_n689), .A2(new_n532), .ZN(new_n690));
  NAND2_X1  g504(.A1(new_n500), .A2(new_n506), .ZN(new_n691));
  OAI211_X1 g505(.A(new_n690), .B(new_n254), .C1(new_n532), .C2(new_n691), .ZN(new_n692));
  NAND2_X1  g506(.A1(new_n692), .A2(G472), .ZN(new_n693));
  NAND2_X1  g507(.A1(new_n565), .A2(new_n693), .ZN(new_n694));
  INV_X1    g508(.A(new_n694), .ZN(new_n695));
  NAND3_X1  g509(.A1(new_n253), .A2(new_n260), .A3(new_n335), .ZN(new_n696));
  OR3_X1    g510(.A1(new_n696), .A2(new_n680), .A3(new_n632), .ZN(new_n697));
  NOR3_X1   g511(.A1(new_n688), .A2(new_n695), .A3(new_n697), .ZN(new_n698));
  INV_X1    g512(.A(KEYINPUT40), .ZN(new_n699));
  AND2_X1   g513(.A1(new_n450), .A2(new_n451), .ZN(new_n700));
  INV_X1    g514(.A(KEYINPUT101), .ZN(new_n701));
  XNOR2_X1  g515(.A(new_n683), .B(KEYINPUT100), .ZN(new_n702));
  XNOR2_X1  g516(.A(new_n702), .B(KEYINPUT39), .ZN(new_n703));
  NAND3_X1  g517(.A1(new_n700), .A2(new_n701), .A3(new_n703), .ZN(new_n704));
  INV_X1    g518(.A(new_n704), .ZN(new_n705));
  AOI21_X1  g519(.A(new_n701), .B1(new_n700), .B2(new_n703), .ZN(new_n706));
  OAI21_X1  g520(.A(new_n699), .B1(new_n705), .B2(new_n706), .ZN(new_n707));
  INV_X1    g521(.A(new_n706), .ZN(new_n708));
  NAND3_X1  g522(.A1(new_n708), .A2(KEYINPUT40), .A3(new_n704), .ZN(new_n709));
  NAND2_X1  g523(.A1(new_n707), .A2(new_n709), .ZN(new_n710));
  NAND2_X1  g524(.A1(new_n698), .A2(new_n710), .ZN(new_n711));
  XNOR2_X1  g525(.A(new_n711), .B(G143), .ZN(G45));
  NAND4_X1  g526(.A1(new_n335), .A2(new_n639), .A3(new_n641), .A4(new_n683), .ZN(new_n713));
  INV_X1    g527(.A(new_n713), .ZN(new_n714));
  NAND4_X1  g528(.A1(new_n634), .A2(new_n678), .A3(new_n681), .A4(new_n714), .ZN(new_n715));
  XNOR2_X1  g529(.A(new_n715), .B(G146), .ZN(G48));
  OAI21_X1  g530(.A(new_n254), .B1(new_n434), .B2(new_n438), .ZN(new_n717));
  NOR2_X1   g531(.A1(new_n346), .A2(KEYINPUT102), .ZN(new_n718));
  AND2_X1   g532(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  NAND2_X1  g533(.A1(new_n437), .A2(new_n420), .ZN(new_n720));
  NAND2_X1  g534(.A1(new_n720), .A2(new_n431), .ZN(new_n721));
  AOI211_X1 g535(.A(G902), .B(new_n718), .C1(new_n721), .C2(new_n433), .ZN(new_n722));
  INV_X1    g536(.A(new_n451), .ZN(new_n723));
  NOR3_X1   g537(.A1(new_n719), .A2(new_n722), .A3(new_n723), .ZN(new_n724));
  NAND4_X1  g538(.A1(new_n566), .A2(new_n634), .A3(new_n642), .A4(new_n724), .ZN(new_n725));
  XOR2_X1   g539(.A(KEYINPUT41), .B(G113), .Z(new_n726));
  XNOR2_X1  g540(.A(new_n726), .B(KEYINPUT103), .ZN(new_n727));
  XNOR2_X1  g541(.A(new_n725), .B(new_n727), .ZN(G15));
  NAND4_X1  g542(.A1(new_n649), .A2(new_n566), .A3(new_n659), .A4(new_n724), .ZN(new_n729));
  XNOR2_X1  g543(.A(new_n729), .B(G116), .ZN(G18));
  AOI21_X1  g544(.A(new_n666), .B1(new_n546), .B2(new_n565), .ZN(new_n731));
  AOI211_X1 g545(.A(new_n343), .B(new_n335), .C1(new_n260), .C2(new_n253), .ZN(new_n732));
  NAND4_X1  g546(.A1(new_n731), .A2(new_n732), .A3(new_n634), .A4(new_n724), .ZN(new_n733));
  XNOR2_X1  g547(.A(new_n733), .B(G119), .ZN(G21));
  NAND2_X1  g548(.A1(new_n696), .A2(KEYINPUT106), .ZN(new_n735));
  INV_X1    g549(.A(KEYINPUT106), .ZN(new_n736));
  NAND4_X1  g550(.A1(new_n253), .A2(new_n260), .A3(new_n335), .A4(new_n736), .ZN(new_n737));
  AND3_X1   g551(.A1(new_n735), .A2(new_n724), .A3(new_n737), .ZN(new_n738));
  NAND2_X1  g552(.A1(new_n537), .A2(new_n533), .ZN(new_n739));
  AOI21_X1  g553(.A(new_n532), .B1(new_n739), .B2(KEYINPUT104), .ZN(new_n740));
  OAI21_X1  g554(.A(new_n740), .B1(KEYINPUT104), .B2(new_n739), .ZN(new_n741));
  NAND2_X1  g555(.A1(new_n552), .A2(new_n554), .ZN(new_n742));
  AOI21_X1  g556(.A(new_n557), .B1(new_n741), .B2(new_n742), .ZN(new_n743));
  INV_X1    g557(.A(KEYINPUT105), .ZN(new_n744));
  NAND2_X1  g558(.A1(new_n629), .A2(new_n744), .ZN(new_n745));
  NAND2_X1  g559(.A1(new_n668), .A2(KEYINPUT105), .ZN(new_n746));
  AOI211_X1 g560(.A(new_n743), .B(new_n486), .C1(new_n745), .C2(new_n746), .ZN(new_n747));
  NAND3_X1  g561(.A1(new_n738), .A2(new_n649), .A3(new_n747), .ZN(new_n748));
  XNOR2_X1  g562(.A(KEYINPUT107), .B(G122), .ZN(new_n749));
  XNOR2_X1  g563(.A(new_n748), .B(new_n749), .ZN(G24));
  NAND2_X1  g564(.A1(new_n745), .A2(new_n746), .ZN(new_n751));
  INV_X1    g565(.A(new_n743), .ZN(new_n752));
  NAND4_X1  g566(.A1(new_n751), .A2(new_n680), .A3(new_n714), .A4(new_n752), .ZN(new_n753));
  NAND2_X1  g567(.A1(new_n633), .A2(new_n610), .ZN(new_n754));
  NAND3_X1  g568(.A1(new_n754), .A2(new_n567), .A3(new_n724), .ZN(new_n755));
  OR2_X1    g569(.A1(new_n753), .A2(new_n755), .ZN(new_n756));
  XNOR2_X1  g570(.A(new_n756), .B(G125), .ZN(G27));
  NAND4_X1  g571(.A1(new_n611), .A2(new_n620), .A3(new_n567), .A4(new_n617), .ZN(new_n758));
  NOR2_X1   g572(.A1(new_n758), .A2(new_n452), .ZN(new_n759));
  AOI211_X1 g573(.A(new_n486), .B(new_n713), .C1(new_n546), .C2(new_n565), .ZN(new_n760));
  INV_X1    g574(.A(KEYINPUT108), .ZN(new_n761));
  NOR2_X1   g575(.A1(new_n761), .A2(KEYINPUT42), .ZN(new_n762));
  INV_X1    g576(.A(new_n762), .ZN(new_n763));
  NAND3_X1  g577(.A1(new_n759), .A2(new_n760), .A3(new_n763), .ZN(new_n764));
  AOI22_X1  g578(.A1(new_n610), .A2(KEYINPUT83), .B1(new_n618), .B2(new_n619), .ZN(new_n765));
  NAND4_X1  g579(.A1(new_n765), .A2(new_n700), .A3(new_n567), .A4(new_n617), .ZN(new_n766));
  NAND3_X1  g580(.A1(new_n678), .A2(new_n626), .A3(new_n714), .ZN(new_n767));
  OAI21_X1  g581(.A(new_n762), .B1(new_n766), .B2(new_n767), .ZN(new_n768));
  NAND2_X1  g582(.A1(new_n764), .A2(new_n768), .ZN(new_n769));
  XNOR2_X1  g583(.A(KEYINPUT109), .B(G131), .ZN(new_n770));
  XNOR2_X1  g584(.A(new_n769), .B(new_n770), .ZN(G33));
  AND2_X1   g585(.A1(new_n678), .A2(new_n684), .ZN(new_n772));
  NAND3_X1  g586(.A1(new_n759), .A2(new_n626), .A3(new_n772), .ZN(new_n773));
  XNOR2_X1  g587(.A(new_n773), .B(G134), .ZN(G36));
  INV_X1    g588(.A(new_n758), .ZN(new_n775));
  NAND2_X1  g589(.A1(new_n639), .A2(new_n641), .ZN(new_n776));
  NOR2_X1   g590(.A1(new_n776), .A2(new_n335), .ZN(new_n777));
  INV_X1    g591(.A(KEYINPUT43), .ZN(new_n778));
  XNOR2_X1  g592(.A(new_n777), .B(new_n778), .ZN(new_n779));
  OAI21_X1  g593(.A(new_n680), .B1(new_n627), .B2(new_n668), .ZN(new_n780));
  OR2_X1    g594(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  INV_X1    g595(.A(KEYINPUT44), .ZN(new_n782));
  OAI21_X1  g596(.A(new_n775), .B1(new_n781), .B2(new_n782), .ZN(new_n783));
  OAI21_X1  g597(.A(new_n782), .B1(new_n779), .B2(new_n780), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n784), .A2(KEYINPUT112), .ZN(new_n785));
  OR2_X1    g599(.A1(new_n784), .A2(KEYINPUT112), .ZN(new_n786));
  AOI21_X1  g600(.A(new_n783), .B1(new_n785), .B2(new_n786), .ZN(new_n787));
  INV_X1    g601(.A(KEYINPUT45), .ZN(new_n788));
  OR2_X1    g602(.A1(new_n449), .A2(new_n788), .ZN(new_n789));
  AOI21_X1  g603(.A(new_n346), .B1(new_n449), .B2(new_n788), .ZN(new_n790));
  AND3_X1   g604(.A1(new_n789), .A2(KEYINPUT110), .A3(new_n790), .ZN(new_n791));
  AOI21_X1  g605(.A(KEYINPUT110), .B1(new_n789), .B2(new_n790), .ZN(new_n792));
  OAI211_X1 g606(.A(KEYINPUT46), .B(new_n441), .C1(new_n791), .C2(new_n792), .ZN(new_n793));
  NAND2_X1  g607(.A1(new_n793), .A2(new_n439), .ZN(new_n794));
  INV_X1    g608(.A(new_n794), .ZN(new_n795));
  OAI21_X1  g609(.A(new_n441), .B1(new_n791), .B2(new_n792), .ZN(new_n796));
  INV_X1    g610(.A(KEYINPUT46), .ZN(new_n797));
  NAND2_X1  g611(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  NAND2_X1  g612(.A1(new_n795), .A2(new_n798), .ZN(new_n799));
  AND2_X1   g613(.A1(new_n703), .A2(new_n451), .ZN(new_n800));
  AOI21_X1  g614(.A(KEYINPUT111), .B1(new_n799), .B2(new_n800), .ZN(new_n801));
  AND3_X1   g615(.A1(new_n799), .A2(KEYINPUT111), .A3(new_n800), .ZN(new_n802));
  OAI21_X1  g616(.A(new_n787), .B1(new_n801), .B2(new_n802), .ZN(new_n803));
  XNOR2_X1  g617(.A(KEYINPUT113), .B(G137), .ZN(new_n804));
  XNOR2_X1  g618(.A(new_n803), .B(new_n804), .ZN(G39));
  INV_X1    g619(.A(KEYINPUT114), .ZN(new_n806));
  AND2_X1   g620(.A1(new_n806), .A2(KEYINPUT47), .ZN(new_n807));
  NOR2_X1   g621(.A1(new_n806), .A2(KEYINPUT47), .ZN(new_n808));
  INV_X1    g622(.A(new_n798), .ZN(new_n809));
  OAI221_X1 g623(.A(new_n451), .B1(new_n807), .B2(new_n808), .C1(new_n809), .C2(new_n794), .ZN(new_n810));
  NOR4_X1   g624(.A1(new_n758), .A2(new_n678), .A3(new_n626), .A4(new_n713), .ZN(new_n811));
  AOI21_X1  g625(.A(new_n723), .B1(new_n795), .B2(new_n798), .ZN(new_n812));
  OAI211_X1 g626(.A(new_n810), .B(new_n811), .C1(new_n812), .C2(new_n808), .ZN(new_n813));
  XNOR2_X1  g627(.A(new_n813), .B(G140), .ZN(G42));
  NAND2_X1  g628(.A1(new_n775), .A2(new_n724), .ZN(new_n815));
  INV_X1    g629(.A(KEYINPUT118), .ZN(new_n816));
  AOI21_X1  g630(.A(new_n338), .B1(new_n815), .B2(new_n816), .ZN(new_n817));
  INV_X1    g631(.A(new_n779), .ZN(new_n818));
  NAND3_X1  g632(.A1(new_n775), .A2(KEYINPUT118), .A3(new_n724), .ZN(new_n819));
  NAND4_X1  g633(.A1(new_n817), .A2(new_n566), .A3(new_n818), .A4(new_n819), .ZN(new_n820));
  OR2_X1    g634(.A1(new_n820), .A2(KEYINPUT120), .ZN(new_n821));
  NAND2_X1  g635(.A1(new_n820), .A2(KEYINPUT120), .ZN(new_n822));
  XNOR2_X1  g636(.A(KEYINPUT121), .B(KEYINPUT48), .ZN(new_n823));
  NAND3_X1  g637(.A1(new_n821), .A2(new_n822), .A3(new_n823), .ZN(new_n824));
  AND2_X1   g638(.A1(new_n817), .A2(new_n819), .ZN(new_n825));
  NAND3_X1  g639(.A1(new_n335), .A2(new_n639), .A3(new_n641), .ZN(new_n826));
  INV_X1    g640(.A(new_n826), .ZN(new_n827));
  NOR2_X1   g641(.A1(new_n694), .A2(new_n486), .ZN(new_n828));
  NAND3_X1  g642(.A1(new_n825), .A2(new_n827), .A3(new_n828), .ZN(new_n829));
  NAND2_X1  g643(.A1(new_n263), .A2(G952), .ZN(new_n830));
  AND3_X1   g644(.A1(new_n818), .A2(new_n339), .A3(new_n747), .ZN(new_n831));
  INV_X1    g645(.A(new_n755), .ZN(new_n832));
  AOI21_X1  g646(.A(new_n830), .B1(new_n831), .B2(new_n832), .ZN(new_n833));
  NAND3_X1  g647(.A1(new_n824), .A2(new_n829), .A3(new_n833), .ZN(new_n834));
  INV_X1    g648(.A(KEYINPUT121), .ZN(new_n835));
  AOI211_X1 g649(.A(new_n835), .B(KEYINPUT48), .C1(new_n821), .C2(new_n822), .ZN(new_n836));
  NOR2_X1   g650(.A1(new_n834), .A2(new_n836), .ZN(new_n837));
  INV_X1    g651(.A(KEYINPUT51), .ZN(new_n838));
  AOI21_X1  g652(.A(new_n743), .B1(new_n745), .B2(new_n746), .ZN(new_n839));
  NAND4_X1  g653(.A1(new_n825), .A2(new_n680), .A3(new_n839), .A4(new_n818), .ZN(new_n840));
  NAND4_X1  g654(.A1(new_n825), .A2(new_n336), .A3(new_n776), .A4(new_n828), .ZN(new_n841));
  AND2_X1   g655(.A1(new_n724), .A2(new_n632), .ZN(new_n842));
  NAND4_X1  g656(.A1(new_n831), .A2(new_n688), .A3(KEYINPUT50), .A4(new_n842), .ZN(new_n843));
  INV_X1    g657(.A(KEYINPUT50), .ZN(new_n844));
  NAND4_X1  g658(.A1(new_n818), .A2(new_n339), .A3(new_n747), .A4(new_n842), .ZN(new_n845));
  INV_X1    g659(.A(new_n688), .ZN(new_n846));
  OAI21_X1  g660(.A(new_n844), .B1(new_n845), .B2(new_n846), .ZN(new_n847));
  NAND2_X1  g661(.A1(new_n843), .A2(new_n847), .ZN(new_n848));
  NAND3_X1  g662(.A1(new_n840), .A2(new_n841), .A3(new_n848), .ZN(new_n849));
  NAND2_X1  g663(.A1(new_n831), .A2(new_n775), .ZN(new_n850));
  OAI21_X1  g664(.A(new_n810), .B1(new_n812), .B2(new_n808), .ZN(new_n851));
  NOR2_X1   g665(.A1(new_n719), .A2(new_n722), .ZN(new_n852));
  NAND2_X1  g666(.A1(new_n852), .A2(new_n723), .ZN(new_n853));
  AOI21_X1  g667(.A(new_n850), .B1(new_n851), .B2(new_n853), .ZN(new_n854));
  OAI21_X1  g668(.A(new_n838), .B1(new_n849), .B2(new_n854), .ZN(new_n855));
  NAND2_X1  g669(.A1(new_n855), .A2(KEYINPUT119), .ZN(new_n856));
  OR3_X1    g670(.A1(new_n849), .A2(new_n854), .A3(new_n838), .ZN(new_n857));
  INV_X1    g671(.A(KEYINPUT119), .ZN(new_n858));
  OAI211_X1 g672(.A(new_n858), .B(new_n838), .C1(new_n849), .C2(new_n854), .ZN(new_n859));
  NAND4_X1  g673(.A1(new_n837), .A2(new_n856), .A3(new_n857), .A4(new_n859), .ZN(new_n860));
  NAND3_X1  g674(.A1(new_n732), .A2(new_n678), .A3(new_n680), .ZN(new_n861));
  NAND2_X1  g675(.A1(new_n674), .A2(new_n675), .ZN(new_n862));
  NOR2_X1   g676(.A1(new_n677), .A2(new_n676), .ZN(new_n863));
  OAI211_X1 g677(.A(new_n724), .B(new_n626), .C1(new_n862), .C2(new_n863), .ZN(new_n864));
  AOI211_X1 g678(.A(new_n569), .B(new_n590), .C1(new_n613), .C2(new_n614), .ZN(new_n865));
  AOI21_X1  g679(.A(new_n570), .B1(new_n615), .B2(new_n591), .ZN(new_n866));
  OAI211_X1 g680(.A(new_n642), .B(new_n567), .C1(new_n865), .C2(new_n866), .ZN(new_n867));
  OAI22_X1  g681(.A1(new_n861), .A2(new_n755), .B1(new_n864), .B2(new_n867), .ZN(new_n868));
  OAI211_X1 g682(.A(new_n567), .B(new_n647), .C1(new_n866), .C2(new_n865), .ZN(new_n869));
  NOR3_X1   g683(.A1(new_n864), .A2(new_n869), .A3(new_n658), .ZN(new_n870));
  NOR2_X1   g684(.A1(new_n868), .A2(new_n870), .ZN(new_n871));
  OAI21_X1  g685(.A(new_n336), .B1(new_n251), .B2(new_n252), .ZN(new_n872));
  NOR2_X1   g686(.A1(new_n872), .A2(new_n648), .ZN(new_n873));
  NAND3_X1  g687(.A1(new_n873), .A2(new_n621), .A3(new_n567), .ZN(new_n874));
  NAND2_X1  g688(.A1(new_n874), .A2(KEYINPUT115), .ZN(new_n875));
  INV_X1    g689(.A(KEYINPUT115), .ZN(new_n876));
  NAND4_X1  g690(.A1(new_n873), .A2(new_n621), .A3(new_n876), .A4(new_n567), .ZN(new_n877));
  NAND3_X1  g691(.A1(new_n875), .A2(new_n631), .A3(new_n877), .ZN(new_n878));
  NAND3_X1  g692(.A1(new_n735), .A2(new_n724), .A3(new_n737), .ZN(new_n879));
  NOR2_X1   g693(.A1(new_n879), .A2(new_n869), .ZN(new_n880));
  NOR4_X1   g694(.A1(new_n630), .A2(new_n452), .A3(new_n826), .A4(new_n648), .ZN(new_n881));
  AOI21_X1  g695(.A(new_n632), .B1(new_n765), .B2(new_n617), .ZN(new_n882));
  AOI22_X1  g696(.A1(new_n880), .A2(new_n747), .B1(new_n881), .B2(new_n882), .ZN(new_n883));
  OAI211_X1 g697(.A(new_n882), .B(new_n453), .C1(new_n566), .C2(new_n669), .ZN(new_n884));
  NAND4_X1  g698(.A1(new_n871), .A2(new_n878), .A3(new_n883), .A4(new_n884), .ZN(new_n885));
  NAND3_X1  g699(.A1(new_n678), .A2(new_n684), .A3(new_n626), .ZN(new_n886));
  AOI21_X1  g700(.A(new_n452), .B1(new_n753), .B2(new_n886), .ZN(new_n887));
  INV_X1    g701(.A(new_n683), .ZN(new_n888));
  NOR3_X1   g702(.A1(new_n251), .A2(new_n252), .A3(new_n888), .ZN(new_n889));
  AND4_X1   g703(.A1(new_n678), .A2(new_n681), .A3(new_n657), .A4(new_n889), .ZN(new_n890));
  OAI21_X1  g704(.A(new_n775), .B1(new_n887), .B2(new_n890), .ZN(new_n891));
  NAND2_X1  g705(.A1(new_n891), .A2(new_n769), .ZN(new_n892));
  NOR2_X1   g706(.A1(new_n885), .A2(new_n892), .ZN(new_n893));
  INV_X1    g707(.A(KEYINPUT116), .ZN(new_n894));
  INV_X1    g708(.A(KEYINPUT52), .ZN(new_n895));
  OAI211_X1 g709(.A(new_n685), .B(new_n715), .C1(new_n755), .C2(new_n753), .ZN(new_n896));
  NAND3_X1  g710(.A1(new_n634), .A2(new_n735), .A3(new_n737), .ZN(new_n897));
  NOR2_X1   g711(.A1(new_n680), .A2(new_n888), .ZN(new_n898));
  NAND3_X1  g712(.A1(new_n694), .A2(new_n700), .A3(new_n898), .ZN(new_n899));
  NOR2_X1   g713(.A1(new_n897), .A2(new_n899), .ZN(new_n900));
  OAI21_X1  g714(.A(new_n895), .B1(new_n896), .B2(new_n900), .ZN(new_n901));
  AOI21_X1  g715(.A(new_n713), .B1(new_n546), .B2(new_n565), .ZN(new_n902));
  OAI211_X1 g716(.A(new_n634), .B(new_n681), .C1(new_n772), .C2(new_n902), .ZN(new_n903));
  AND3_X1   g717(.A1(new_n694), .A2(new_n700), .A3(new_n898), .ZN(new_n904));
  NAND4_X1  g718(.A1(new_n904), .A2(new_n634), .A3(new_n735), .A4(new_n737), .ZN(new_n905));
  NAND4_X1  g719(.A1(new_n903), .A2(new_n905), .A3(new_n756), .A4(KEYINPUT52), .ZN(new_n906));
  AOI21_X1  g720(.A(new_n894), .B1(new_n901), .B2(new_n906), .ZN(new_n907));
  AND2_X1   g721(.A1(new_n906), .A2(new_n894), .ZN(new_n908));
  OAI211_X1 g722(.A(new_n893), .B(KEYINPUT53), .C1(new_n907), .C2(new_n908), .ZN(new_n909));
  NAND2_X1  g723(.A1(new_n901), .A2(new_n906), .ZN(new_n910));
  AND2_X1   g724(.A1(new_n891), .A2(new_n769), .ZN(new_n911));
  NAND3_X1  g725(.A1(new_n729), .A2(new_n725), .A3(new_n733), .ZN(new_n912));
  NOR2_X1   g726(.A1(new_n826), .A2(new_n648), .ZN(new_n913));
  NAND4_X1  g727(.A1(new_n631), .A2(new_n567), .A3(new_n621), .A4(new_n913), .ZN(new_n914));
  NAND2_X1  g728(.A1(new_n748), .A2(new_n914), .ZN(new_n915));
  NAND2_X1  g729(.A1(new_n622), .A2(new_n670), .ZN(new_n916));
  NOR3_X1   g730(.A1(new_n912), .A2(new_n915), .A3(new_n916), .ZN(new_n917));
  NAND4_X1  g731(.A1(new_n910), .A2(new_n911), .A3(new_n878), .A4(new_n917), .ZN(new_n918));
  XNOR2_X1  g732(.A(KEYINPUT117), .B(KEYINPUT53), .ZN(new_n919));
  NAND2_X1  g733(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  INV_X1    g734(.A(KEYINPUT54), .ZN(new_n921));
  NAND3_X1  g735(.A1(new_n909), .A2(new_n920), .A3(new_n921), .ZN(new_n922));
  NOR2_X1   g736(.A1(new_n918), .A2(new_n919), .ZN(new_n923));
  INV_X1    g737(.A(KEYINPUT53), .ZN(new_n924));
  OAI21_X1  g738(.A(new_n893), .B1(new_n907), .B2(new_n908), .ZN(new_n925));
  AOI21_X1  g739(.A(new_n923), .B1(new_n924), .B2(new_n925), .ZN(new_n926));
  OAI21_X1  g740(.A(new_n922), .B1(new_n926), .B2(new_n921), .ZN(new_n927));
  NOR2_X1   g741(.A1(new_n860), .A2(new_n927), .ZN(new_n928));
  NOR2_X1   g742(.A1(G952), .A2(G953), .ZN(new_n929));
  XNOR2_X1  g743(.A(new_n852), .B(KEYINPUT49), .ZN(new_n930));
  NOR3_X1   g744(.A1(new_n486), .A2(new_n632), .A3(new_n723), .ZN(new_n931));
  NAND4_X1  g745(.A1(new_n930), .A2(new_n695), .A3(new_n777), .A4(new_n931), .ZN(new_n932));
  OAI22_X1  g746(.A1(new_n928), .A2(new_n929), .B1(new_n846), .B2(new_n932), .ZN(G75));
  NOR2_X1   g747(.A1(new_n263), .A2(G952), .ZN(new_n934));
  XNOR2_X1  g748(.A(new_n934), .B(KEYINPUT122), .ZN(new_n935));
  AOI21_X1  g749(.A(new_n254), .B1(new_n909), .B2(new_n920), .ZN(new_n936));
  AND2_X1   g750(.A1(new_n936), .A2(new_n619), .ZN(new_n937));
  XOR2_X1   g751(.A(new_n602), .B(new_n605), .Z(new_n938));
  XNOR2_X1  g752(.A(new_n938), .B(KEYINPUT55), .ZN(new_n939));
  INV_X1    g753(.A(KEYINPUT56), .ZN(new_n940));
  NAND2_X1  g754(.A1(new_n939), .A2(new_n940), .ZN(new_n941));
  OAI21_X1  g755(.A(new_n935), .B1(new_n937), .B2(new_n941), .ZN(new_n942));
  NAND2_X1  g756(.A1(new_n936), .A2(new_n569), .ZN(new_n943));
  AOI21_X1  g757(.A(new_n939), .B1(new_n943), .B2(new_n940), .ZN(new_n944));
  NOR2_X1   g758(.A1(new_n942), .A2(new_n944), .ZN(G51));
  NAND2_X1  g759(.A1(new_n909), .A2(new_n920), .ZN(new_n946));
  XNOR2_X1  g760(.A(new_n946), .B(new_n921), .ZN(new_n947));
  XOR2_X1   g761(.A(new_n440), .B(KEYINPUT57), .Z(new_n948));
  OAI22_X1  g762(.A1(new_n947), .A2(new_n948), .B1(new_n438), .B2(new_n434), .ZN(new_n949));
  INV_X1    g763(.A(new_n936), .ZN(new_n950));
  OR3_X1    g764(.A1(new_n950), .A2(new_n792), .A3(new_n791), .ZN(new_n951));
  AOI21_X1  g765(.A(new_n934), .B1(new_n949), .B2(new_n951), .ZN(G54));
  AND2_X1   g766(.A1(KEYINPUT58), .A2(G475), .ZN(new_n953));
  AND3_X1   g767(.A1(new_n936), .A2(new_n329), .A3(new_n953), .ZN(new_n954));
  AOI21_X1  g768(.A(new_n329), .B1(new_n936), .B2(new_n953), .ZN(new_n955));
  NOR3_X1   g769(.A1(new_n954), .A2(new_n955), .A3(new_n934), .ZN(G60));
  NOR2_X1   g770(.A1(new_n636), .A2(new_n638), .ZN(new_n957));
  XOR2_X1   g771(.A(new_n640), .B(KEYINPUT59), .Z(new_n958));
  NAND2_X1  g772(.A1(new_n957), .A2(new_n958), .ZN(new_n959));
  OAI21_X1  g773(.A(new_n935), .B1(new_n947), .B2(new_n959), .ZN(new_n960));
  AOI21_X1  g774(.A(new_n957), .B1(new_n927), .B2(new_n958), .ZN(new_n961));
  NOR2_X1   g775(.A1(new_n960), .A2(new_n961), .ZN(G63));
  NAND2_X1  g776(.A1(G217), .A2(G902), .ZN(new_n963));
  XOR2_X1   g777(.A(new_n963), .B(KEYINPUT123), .Z(new_n964));
  XOR2_X1   g778(.A(new_n964), .B(KEYINPUT60), .Z(new_n965));
  NAND3_X1  g779(.A1(new_n946), .A2(new_n665), .A3(new_n965), .ZN(new_n966));
  INV_X1    g780(.A(new_n965), .ZN(new_n967));
  AOI21_X1  g781(.A(new_n967), .B1(new_n909), .B2(new_n920), .ZN(new_n968));
  OAI211_X1 g782(.A(new_n966), .B(new_n935), .C1(new_n483), .C2(new_n968), .ZN(new_n969));
  NAND3_X1  g783(.A1(new_n966), .A2(KEYINPUT124), .A3(new_n935), .ZN(new_n970));
  NAND3_X1  g784(.A1(new_n969), .A2(KEYINPUT61), .A3(new_n970), .ZN(new_n971));
  OR2_X1    g785(.A1(new_n968), .A2(new_n483), .ZN(new_n972));
  INV_X1    g786(.A(new_n935), .ZN(new_n973));
  AOI21_X1  g787(.A(new_n973), .B1(new_n968), .B2(new_n665), .ZN(new_n974));
  INV_X1    g788(.A(KEYINPUT61), .ZN(new_n975));
  OAI211_X1 g789(.A(new_n972), .B(new_n974), .C1(KEYINPUT124), .C2(new_n975), .ZN(new_n976));
  AND2_X1   g790(.A1(new_n971), .A2(new_n976), .ZN(G66));
  OAI21_X1  g791(.A(G953), .B1(new_n342), .B2(new_n572), .ZN(new_n978));
  INV_X1    g792(.A(new_n885), .ZN(new_n979));
  OAI21_X1  g793(.A(new_n978), .B1(new_n979), .B2(G953), .ZN(new_n980));
  INV_X1    g794(.A(G898), .ZN(new_n981));
  AOI21_X1  g795(.A(new_n602), .B1(new_n981), .B2(G953), .ZN(new_n982));
  XNOR2_X1  g796(.A(new_n982), .B(KEYINPUT125), .ZN(new_n983));
  XNOR2_X1  g797(.A(new_n980), .B(new_n983), .ZN(G69));
  AOI21_X1  g798(.A(new_n263), .B1(G227), .B2(G900), .ZN(new_n985));
  INV_X1    g799(.A(KEYINPUT126), .ZN(new_n986));
  NAND2_X1  g800(.A1(new_n985), .A2(new_n986), .ZN(new_n987));
  XOR2_X1   g801(.A(new_n987), .B(KEYINPUT127), .Z(new_n988));
  INV_X1    g802(.A(new_n566), .ZN(new_n989));
  AOI21_X1  g803(.A(new_n989), .B1(new_n826), .B2(new_n872), .ZN(new_n990));
  NOR2_X1   g804(.A1(new_n705), .A2(new_n706), .ZN(new_n991));
  NAND3_X1  g805(.A1(new_n990), .A2(new_n991), .A3(new_n775), .ZN(new_n992));
  NAND2_X1  g806(.A1(new_n803), .A2(new_n992), .ZN(new_n993));
  INV_X1    g807(.A(new_n896), .ZN(new_n994));
  AOI21_X1  g808(.A(KEYINPUT62), .B1(new_n711), .B2(new_n994), .ZN(new_n995));
  INV_X1    g809(.A(KEYINPUT62), .ZN(new_n996));
  AOI211_X1 g810(.A(new_n996), .B(new_n896), .C1(new_n698), .C2(new_n710), .ZN(new_n997));
  OAI21_X1  g811(.A(new_n813), .B1(new_n995), .B2(new_n997), .ZN(new_n998));
  OAI21_X1  g812(.A(new_n263), .B1(new_n993), .B2(new_n998), .ZN(new_n999));
  NOR2_X1   g813(.A1(new_n314), .A2(new_n315), .ZN(new_n1000));
  XNOR2_X1  g814(.A(new_n548), .B(new_n1000), .ZN(new_n1001));
  NAND2_X1  g815(.A1(new_n999), .A2(new_n1001), .ZN(new_n1002));
  AOI21_X1  g816(.A(new_n1001), .B1(G900), .B2(G953), .ZN(new_n1003));
  NOR2_X1   g817(.A1(new_n897), .A2(new_n989), .ZN(new_n1004));
  OAI21_X1  g818(.A(new_n1004), .B1(new_n802), .B2(new_n801), .ZN(new_n1005));
  AND3_X1   g819(.A1(new_n994), .A2(new_n769), .A3(new_n773), .ZN(new_n1006));
  NAND4_X1  g820(.A1(new_n803), .A2(new_n1005), .A3(new_n1006), .A4(new_n813), .ZN(new_n1007));
  OAI21_X1  g821(.A(new_n1003), .B1(new_n1007), .B2(G953), .ZN(new_n1008));
  NAND2_X1  g822(.A1(new_n1002), .A2(new_n1008), .ZN(new_n1009));
  NOR2_X1   g823(.A1(new_n985), .A2(new_n986), .ZN(new_n1010));
  INV_X1    g824(.A(new_n1010), .ZN(new_n1011));
  AOI21_X1  g825(.A(new_n988), .B1(new_n1009), .B2(new_n1011), .ZN(new_n1012));
  INV_X1    g826(.A(new_n988), .ZN(new_n1013));
  AOI211_X1 g827(.A(new_n1010), .B(new_n1013), .C1(new_n1002), .C2(new_n1008), .ZN(new_n1014));
  NOR2_X1   g828(.A1(new_n1012), .A2(new_n1014), .ZN(G72));
  OR3_X1    g829(.A1(new_n993), .A2(new_n998), .A3(new_n885), .ZN(new_n1016));
  NAND2_X1  g830(.A1(G472), .A2(G902), .ZN(new_n1017));
  XOR2_X1   g831(.A(new_n1017), .B(KEYINPUT63), .Z(new_n1018));
  AOI21_X1  g832(.A(new_n690), .B1(new_n1016), .B2(new_n1018), .ZN(new_n1019));
  OAI21_X1  g833(.A(new_n1018), .B1(new_n1007), .B2(new_n885), .ZN(new_n1020));
  AND3_X1   g834(.A1(new_n1020), .A2(new_n519), .A3(new_n553), .ZN(new_n1021));
  INV_X1    g835(.A(new_n1018), .ZN(new_n1022));
  AND2_X1   g836(.A1(new_n550), .A2(new_n528), .ZN(new_n1023));
  NOR3_X1   g837(.A1(new_n926), .A2(new_n1022), .A3(new_n1023), .ZN(new_n1024));
  NOR4_X1   g838(.A1(new_n1019), .A2(new_n1021), .A3(new_n1024), .A4(new_n934), .ZN(G57));
endmodule


