//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 0 1 0 1 0 0 1 0 1 0 0 1 1 1 1 0 0 0 0 1 1 0 1 1 0 0 1 1 1 1 0 1 0 1 1 0 0 1 0 0 0 1 1 1 1 0 0 1 1 0 0 1 0 0 1 0 0 0 1 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:42:49 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n817, new_n818, new_n819, new_n820,
    new_n821, new_n822, new_n823, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1196, new_n1197, new_n1198, new_n1199,
    new_n1200, new_n1201, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1219, new_n1220, new_n1221, new_n1222, new_n1223, new_n1225,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1294, new_n1295, new_n1296, new_n1297, new_n1298, new_n1299,
    new_n1300, new_n1301, new_n1302, new_n1303, new_n1304;
  INV_X1    g0000(.A(G50), .ZN(new_n201));
  INV_X1    g0001(.A(G58), .ZN(new_n202));
  INV_X1    g0002(.A(G68), .ZN(new_n203));
  NAND3_X1  g0003(.A1(new_n201), .A2(new_n202), .A3(new_n203), .ZN(new_n204));
  NOR2_X1   g0004(.A1(new_n204), .A2(G77), .ZN(G353));
  OAI21_X1  g0005(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0006(.A(G1), .ZN(new_n207));
  INV_X1    g0007(.A(G20), .ZN(new_n208));
  NOR2_X1   g0008(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  INV_X1    g0009(.A(new_n209), .ZN(new_n210));
  NOR2_X1   g0010(.A1(new_n210), .A2(G13), .ZN(new_n211));
  OAI211_X1 g0011(.A(new_n211), .B(G250), .C1(G257), .C2(G264), .ZN(new_n212));
  XNOR2_X1  g0012(.A(new_n212), .B(KEYINPUT0), .ZN(new_n213));
  NAND2_X1  g0013(.A1(G1), .A2(G13), .ZN(new_n214));
  INV_X1    g0014(.A(new_n214), .ZN(new_n215));
  NAND2_X1  g0015(.A1(new_n215), .A2(G20), .ZN(new_n216));
  XNOR2_X1  g0016(.A(new_n216), .B(KEYINPUT64), .ZN(new_n217));
  OAI21_X1  g0017(.A(G50), .B1(G58), .B2(G68), .ZN(new_n218));
  AOI22_X1  g0018(.A1(G107), .A2(G264), .B1(G116), .B2(G270), .ZN(new_n219));
  INV_X1    g0019(.A(G77), .ZN(new_n220));
  INV_X1    g0020(.A(G244), .ZN(new_n221));
  INV_X1    g0021(.A(G87), .ZN(new_n222));
  INV_X1    g0022(.A(G250), .ZN(new_n223));
  OAI221_X1 g0023(.A(new_n219), .B1(new_n220), .B2(new_n221), .C1(new_n222), .C2(new_n223), .ZN(new_n224));
  AOI22_X1  g0024(.A1(G50), .A2(G226), .B1(G97), .B2(G257), .ZN(new_n225));
  INV_X1    g0025(.A(G232), .ZN(new_n226));
  INV_X1    g0026(.A(G238), .ZN(new_n227));
  OAI221_X1 g0027(.A(new_n225), .B1(new_n202), .B2(new_n226), .C1(new_n203), .C2(new_n227), .ZN(new_n228));
  OAI21_X1  g0028(.A(new_n210), .B1(new_n224), .B2(new_n228), .ZN(new_n229));
  OAI221_X1 g0029(.A(new_n213), .B1(new_n217), .B2(new_n218), .C1(KEYINPUT1), .C2(new_n229), .ZN(new_n230));
  AOI21_X1  g0030(.A(new_n230), .B1(KEYINPUT1), .B2(new_n229), .ZN(G361));
  XNOR2_X1  g0031(.A(G238), .B(G244), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n232), .B(KEYINPUT66), .ZN(new_n233));
  XNOR2_X1  g0033(.A(G226), .B(G232), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XNOR2_X1  g0035(.A(KEYINPUT65), .B(KEYINPUT2), .ZN(new_n236));
  XOR2_X1   g0036(.A(new_n235), .B(new_n236), .Z(new_n237));
  XNOR2_X1  g0037(.A(G264), .B(G270), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n238), .B(KEYINPUT67), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n239), .B(new_n223), .ZN(new_n240));
  INV_X1    g0040(.A(G257), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n237), .B(new_n242), .ZN(G358));
  XOR2_X1   g0043(.A(G68), .B(G77), .Z(new_n244));
  XNOR2_X1  g0044(.A(G50), .B(G58), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XOR2_X1   g0046(.A(G87), .B(G97), .Z(new_n247));
  XNOR2_X1  g0047(.A(G107), .B(G116), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n247), .B(new_n248), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n246), .B(new_n249), .ZN(G351));
  INV_X1    g0050(.A(G33), .ZN(new_n251));
  INV_X1    g0051(.A(G41), .ZN(new_n252));
  OAI21_X1  g0052(.A(new_n215), .B1(new_n251), .B2(new_n252), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n251), .A2(KEYINPUT3), .ZN(new_n254));
  INV_X1    g0054(.A(KEYINPUT3), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n255), .A2(G33), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n254), .A2(new_n256), .ZN(new_n257));
  INV_X1    g0057(.A(new_n257), .ZN(new_n258));
  INV_X1    g0058(.A(G1698), .ZN(new_n259));
  NAND3_X1  g0059(.A1(new_n258), .A2(G222), .A3(new_n259), .ZN(new_n260));
  XOR2_X1   g0060(.A(new_n260), .B(KEYINPUT70), .Z(new_n261));
  NOR2_X1   g0061(.A1(new_n257), .A2(new_n259), .ZN(new_n262));
  AOI22_X1  g0062(.A1(new_n262), .A2(G223), .B1(G77), .B2(new_n257), .ZN(new_n263));
  AOI21_X1  g0063(.A(new_n253), .B1(new_n261), .B2(new_n263), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n252), .A2(KEYINPUT68), .ZN(new_n265));
  INV_X1    g0065(.A(KEYINPUT68), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n266), .A2(G41), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n265), .A2(new_n267), .ZN(new_n268));
  OAI211_X1 g0068(.A(new_n207), .B(G274), .C1(new_n268), .C2(G45), .ZN(new_n269));
  OAI21_X1  g0069(.A(new_n207), .B1(G41), .B2(G45), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n253), .A2(new_n270), .ZN(new_n271));
  XNOR2_X1  g0071(.A(new_n271), .B(KEYINPUT69), .ZN(new_n272));
  INV_X1    g0072(.A(G226), .ZN(new_n273));
  OAI21_X1  g0073(.A(new_n269), .B1(new_n272), .B2(new_n273), .ZN(new_n274));
  OR2_X1    g0074(.A1(new_n264), .A2(new_n274), .ZN(new_n275));
  XOR2_X1   g0075(.A(KEYINPUT77), .B(G200), .Z(new_n276));
  INV_X1    g0076(.A(new_n276), .ZN(new_n277));
  INV_X1    g0077(.A(KEYINPUT79), .ZN(new_n278));
  AOI22_X1  g0078(.A1(new_n275), .A2(new_n277), .B1(new_n278), .B2(KEYINPUT10), .ZN(new_n279));
  AOI21_X1  g0079(.A(new_n215), .B1(new_n209), .B2(G33), .ZN(new_n280));
  XNOR2_X1  g0080(.A(KEYINPUT8), .B(G58), .ZN(new_n281));
  INV_X1    g0081(.A(KEYINPUT71), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  OR3_X1    g0083(.A1(new_n282), .A2(new_n202), .A3(KEYINPUT8), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  INV_X1    g0085(.A(new_n285), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n208), .A2(G33), .ZN(new_n287));
  XOR2_X1   g0087(.A(new_n287), .B(KEYINPUT72), .Z(new_n288));
  NAND2_X1  g0088(.A1(new_n286), .A2(new_n288), .ZN(new_n289));
  NOR2_X1   g0089(.A1(G20), .A2(G33), .ZN(new_n290));
  AOI22_X1  g0090(.A1(new_n204), .A2(G20), .B1(G150), .B2(new_n290), .ZN(new_n291));
  AOI21_X1  g0091(.A(new_n280), .B1(new_n289), .B2(new_n291), .ZN(new_n292));
  NAND3_X1  g0092(.A1(new_n207), .A2(G13), .A3(G20), .ZN(new_n293));
  INV_X1    g0093(.A(new_n293), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n294), .A2(new_n201), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n207), .A2(G20), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n280), .A2(new_n296), .ZN(new_n297));
  OAI21_X1  g0097(.A(new_n295), .B1(new_n297), .B2(new_n201), .ZN(new_n298));
  OR2_X1    g0098(.A1(new_n292), .A2(new_n298), .ZN(new_n299));
  INV_X1    g0099(.A(KEYINPUT9), .ZN(new_n300));
  NOR2_X1   g0100(.A1(new_n299), .A2(new_n300), .ZN(new_n301));
  NOR2_X1   g0101(.A1(new_n264), .A2(new_n274), .ZN(new_n302));
  AOI21_X1  g0102(.A(new_n301), .B1(G190), .B2(new_n302), .ZN(new_n303));
  INV_X1    g0103(.A(KEYINPUT78), .ZN(new_n304));
  AOI21_X1  g0104(.A(new_n304), .B1(new_n299), .B2(new_n300), .ZN(new_n305));
  NAND3_X1  g0105(.A1(new_n299), .A2(new_n304), .A3(new_n300), .ZN(new_n306));
  INV_X1    g0106(.A(new_n306), .ZN(new_n307));
  OAI211_X1 g0107(.A(new_n279), .B(new_n303), .C1(new_n305), .C2(new_n307), .ZN(new_n308));
  NOR2_X1   g0108(.A1(new_n278), .A2(KEYINPUT10), .ZN(new_n309));
  INV_X1    g0109(.A(new_n309), .ZN(new_n310));
  XNOR2_X1  g0110(.A(new_n308), .B(new_n310), .ZN(new_n311));
  INV_X1    g0111(.A(G169), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n275), .A2(new_n312), .ZN(new_n313));
  INV_X1    g0113(.A(G179), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n302), .A2(new_n314), .ZN(new_n315));
  NAND3_X1  g0115(.A1(new_n313), .A2(new_n299), .A3(new_n315), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n311), .A2(new_n316), .ZN(new_n317));
  OR2_X1    g0117(.A1(new_n293), .A2(KEYINPUT74), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n293), .A2(KEYINPUT74), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n318), .A2(new_n319), .ZN(new_n320));
  INV_X1    g0120(.A(new_n320), .ZN(new_n321));
  INV_X1    g0121(.A(new_n280), .ZN(new_n322));
  NOR2_X1   g0122(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  NAND3_X1  g0123(.A1(new_n323), .A2(G68), .A3(new_n296), .ZN(new_n324));
  XNOR2_X1  g0124(.A(new_n324), .B(KEYINPUT80), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n288), .A2(G77), .ZN(new_n326));
  AOI22_X1  g0126(.A1(new_n290), .A2(G50), .B1(G20), .B2(new_n203), .ZN(new_n327));
  AOI21_X1  g0127(.A(new_n280), .B1(new_n326), .B2(new_n327), .ZN(new_n328));
  OR2_X1    g0128(.A1(new_n328), .A2(KEYINPUT11), .ZN(new_n329));
  NAND3_X1  g0129(.A1(new_n321), .A2(KEYINPUT12), .A3(new_n203), .ZN(new_n330));
  NOR2_X1   g0130(.A1(new_n293), .A2(G68), .ZN(new_n331));
  OAI21_X1  g0131(.A(new_n330), .B1(KEYINPUT12), .B2(new_n331), .ZN(new_n332));
  AOI21_X1  g0132(.A(new_n332), .B1(new_n328), .B2(KEYINPUT11), .ZN(new_n333));
  NAND3_X1  g0133(.A1(new_n325), .A2(new_n329), .A3(new_n333), .ZN(new_n334));
  INV_X1    g0134(.A(KEYINPUT14), .ZN(new_n335));
  XOR2_X1   g0135(.A(new_n271), .B(KEYINPUT69), .Z(new_n336));
  NAND2_X1  g0136(.A1(new_n336), .A2(G238), .ZN(new_n337));
  INV_X1    g0137(.A(KEYINPUT13), .ZN(new_n338));
  INV_X1    g0138(.A(new_n269), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n226), .A2(G1698), .ZN(new_n340));
  OAI21_X1  g0140(.A(new_n340), .B1(G226), .B2(G1698), .ZN(new_n341));
  INV_X1    g0141(.A(G97), .ZN(new_n342));
  OAI22_X1  g0142(.A1(new_n341), .A2(new_n257), .B1(new_n251), .B2(new_n342), .ZN(new_n343));
  AOI21_X1  g0143(.A(new_n214), .B1(G33), .B2(G41), .ZN(new_n344));
  AOI21_X1  g0144(.A(new_n339), .B1(new_n343), .B2(new_n344), .ZN(new_n345));
  NAND3_X1  g0145(.A1(new_n337), .A2(new_n338), .A3(new_n345), .ZN(new_n346));
  INV_X1    g0146(.A(new_n346), .ZN(new_n347));
  AOI21_X1  g0147(.A(new_n338), .B1(new_n337), .B2(new_n345), .ZN(new_n348));
  OAI211_X1 g0148(.A(new_n335), .B(G169), .C1(new_n347), .C2(new_n348), .ZN(new_n349));
  INV_X1    g0149(.A(new_n348), .ZN(new_n350));
  NAND3_X1  g0150(.A1(new_n350), .A2(G179), .A3(new_n346), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n349), .A2(new_n351), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n350), .A2(new_n346), .ZN(new_n353));
  AOI21_X1  g0153(.A(new_n335), .B1(new_n353), .B2(G169), .ZN(new_n354));
  OAI21_X1  g0154(.A(new_n334), .B1(new_n352), .B2(new_n354), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n353), .A2(G200), .ZN(new_n356));
  INV_X1    g0156(.A(new_n334), .ZN(new_n357));
  INV_X1    g0157(.A(G190), .ZN(new_n358));
  OAI211_X1 g0158(.A(new_n356), .B(new_n357), .C1(new_n358), .C2(new_n353), .ZN(new_n359));
  NAND3_X1  g0159(.A1(new_n323), .A2(G77), .A3(new_n296), .ZN(new_n360));
  XNOR2_X1  g0160(.A(new_n360), .B(KEYINPUT75), .ZN(new_n361));
  INV_X1    g0161(.A(KEYINPUT76), .ZN(new_n362));
  NAND2_X1  g0162(.A1(G20), .A2(G77), .ZN(new_n363));
  INV_X1    g0163(.A(new_n290), .ZN(new_n364));
  XNOR2_X1  g0164(.A(KEYINPUT15), .B(G87), .ZN(new_n365));
  OAI221_X1 g0165(.A(new_n363), .B1(new_n281), .B2(new_n364), .C1(new_n287), .C2(new_n365), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n366), .A2(new_n322), .ZN(new_n367));
  OAI21_X1  g0167(.A(new_n367), .B1(G77), .B2(new_n320), .ZN(new_n368));
  OR3_X1    g0168(.A1(new_n361), .A2(new_n362), .A3(new_n368), .ZN(new_n369));
  OAI21_X1  g0169(.A(new_n269), .B1(new_n272), .B2(new_n221), .ZN(new_n370));
  INV_X1    g0170(.A(KEYINPUT73), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  OAI211_X1 g0172(.A(KEYINPUT73), .B(new_n269), .C1(new_n272), .C2(new_n221), .ZN(new_n373));
  NAND3_X1  g0173(.A1(new_n258), .A2(G232), .A3(new_n259), .ZN(new_n374));
  INV_X1    g0174(.A(G107), .ZN(new_n375));
  OAI21_X1  g0175(.A(new_n374), .B1(new_n375), .B2(new_n258), .ZN(new_n376));
  AOI21_X1  g0176(.A(new_n376), .B1(G238), .B2(new_n262), .ZN(new_n377));
  OAI211_X1 g0177(.A(new_n372), .B(new_n373), .C1(new_n253), .C2(new_n377), .ZN(new_n378));
  OR2_X1    g0178(.A1(new_n378), .A2(new_n358), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n378), .A2(new_n277), .ZN(new_n380));
  OAI21_X1  g0180(.A(new_n362), .B1(new_n361), .B2(new_n368), .ZN(new_n381));
  NAND4_X1  g0181(.A1(new_n369), .A2(new_n379), .A3(new_n380), .A4(new_n381), .ZN(new_n382));
  OR2_X1    g0182(.A1(new_n378), .A2(G179), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n378), .A2(new_n312), .ZN(new_n384));
  OR2_X1    g0184(.A1(new_n361), .A2(new_n368), .ZN(new_n385));
  NAND3_X1  g0185(.A1(new_n383), .A2(new_n384), .A3(new_n385), .ZN(new_n386));
  NAND4_X1  g0186(.A1(new_n355), .A2(new_n359), .A3(new_n382), .A4(new_n386), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n285), .A2(new_n294), .ZN(new_n388));
  OAI21_X1  g0188(.A(new_n388), .B1(new_n285), .B2(new_n297), .ZN(new_n389));
  INV_X1    g0189(.A(new_n389), .ZN(new_n390));
  NOR2_X1   g0190(.A1(new_n202), .A2(new_n203), .ZN(new_n391));
  NOR2_X1   g0191(.A1(G58), .A2(G68), .ZN(new_n392));
  OAI21_X1  g0192(.A(G20), .B1(new_n391), .B2(new_n392), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n290), .A2(G159), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n393), .A2(new_n394), .ZN(new_n395));
  INV_X1    g0195(.A(KEYINPUT16), .ZN(new_n396));
  NOR2_X1   g0196(.A1(new_n395), .A2(new_n396), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n251), .A2(KEYINPUT81), .ZN(new_n398));
  INV_X1    g0198(.A(KEYINPUT81), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n399), .A2(G33), .ZN(new_n400));
  NAND3_X1  g0200(.A1(new_n398), .A2(new_n400), .A3(KEYINPUT3), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n255), .A2(KEYINPUT82), .ZN(new_n402));
  INV_X1    g0202(.A(KEYINPUT82), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n403), .A2(KEYINPUT3), .ZN(new_n404));
  NAND3_X1  g0204(.A1(new_n402), .A2(new_n404), .A3(G33), .ZN(new_n405));
  AOI21_X1  g0205(.A(G20), .B1(new_n401), .B2(new_n405), .ZN(new_n406));
  INV_X1    g0206(.A(KEYINPUT7), .ZN(new_n407));
  OAI21_X1  g0207(.A(G68), .B1(new_n406), .B2(new_n407), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n407), .A2(KEYINPUT83), .ZN(new_n409));
  INV_X1    g0209(.A(KEYINPUT83), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n410), .A2(KEYINPUT7), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n409), .A2(new_n411), .ZN(new_n412));
  AOI211_X1 g0212(.A(G20), .B(new_n412), .C1(new_n401), .C2(new_n405), .ZN(new_n413));
  OAI21_X1  g0213(.A(new_n397), .B1(new_n408), .B2(new_n413), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n414), .A2(new_n322), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n208), .A2(KEYINPUT7), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n402), .A2(new_n404), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n417), .A2(new_n251), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n398), .A2(new_n400), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n419), .A2(new_n255), .ZN(new_n420));
  AOI21_X1  g0220(.A(new_n416), .B1(new_n418), .B2(new_n420), .ZN(new_n421));
  AOI21_X1  g0221(.A(new_n412), .B1(new_n208), .B2(new_n257), .ZN(new_n422));
  OAI21_X1  g0222(.A(G68), .B1(new_n421), .B2(new_n422), .ZN(new_n423));
  INV_X1    g0223(.A(new_n395), .ZN(new_n424));
  AOI21_X1  g0224(.A(KEYINPUT16), .B1(new_n423), .B2(new_n424), .ZN(new_n425));
  OAI21_X1  g0225(.A(new_n390), .B1(new_n415), .B2(new_n425), .ZN(new_n426));
  NOR2_X1   g0226(.A1(G223), .A2(G1698), .ZN(new_n427));
  AOI21_X1  g0227(.A(new_n427), .B1(new_n273), .B2(G1698), .ZN(new_n428));
  NAND3_X1  g0228(.A1(new_n401), .A2(new_n428), .A3(new_n405), .ZN(new_n429));
  NAND2_X1  g0229(.A1(G33), .A2(G87), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n429), .A2(new_n430), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n431), .A2(new_n344), .ZN(new_n432));
  NAND3_X1  g0232(.A1(new_n253), .A2(G232), .A3(new_n270), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n269), .A2(new_n433), .ZN(new_n434));
  INV_X1    g0234(.A(new_n434), .ZN(new_n435));
  NAND3_X1  g0235(.A1(new_n432), .A2(G179), .A3(new_n435), .ZN(new_n436));
  AOI21_X1  g0236(.A(new_n253), .B1(new_n429), .B2(new_n430), .ZN(new_n437));
  OAI21_X1  g0237(.A(G169), .B1(new_n437), .B2(new_n434), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n436), .A2(new_n438), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n426), .A2(new_n439), .ZN(new_n440));
  INV_X1    g0240(.A(KEYINPUT18), .ZN(new_n441));
  XNOR2_X1  g0241(.A(new_n440), .B(new_n441), .ZN(new_n442));
  NAND3_X1  g0242(.A1(new_n432), .A2(new_n358), .A3(new_n435), .ZN(new_n443));
  INV_X1    g0243(.A(G200), .ZN(new_n444));
  OAI21_X1  g0244(.A(new_n444), .B1(new_n437), .B2(new_n434), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n443), .A2(new_n445), .ZN(new_n446));
  OAI211_X1 g0246(.A(new_n446), .B(new_n390), .C1(new_n415), .C2(new_n425), .ZN(new_n447));
  XNOR2_X1  g0247(.A(KEYINPUT84), .B(KEYINPUT17), .ZN(new_n448));
  INV_X1    g0248(.A(new_n448), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n447), .A2(new_n449), .ZN(new_n450));
  INV_X1    g0250(.A(KEYINPUT17), .ZN(new_n451));
  NOR2_X1   g0251(.A1(new_n451), .A2(KEYINPUT84), .ZN(new_n452));
  OAI21_X1  g0252(.A(new_n450), .B1(new_n447), .B2(new_n452), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n442), .A2(new_n453), .ZN(new_n454));
  NOR3_X1   g0254(.A1(new_n317), .A2(new_n387), .A3(new_n454), .ZN(new_n455));
  AND2_X1   g0255(.A1(new_n401), .A2(new_n405), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n241), .A2(new_n259), .ZN(new_n457));
  OAI211_X1 g0257(.A(new_n456), .B(new_n457), .C1(G264), .C2(new_n259), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n257), .A2(G303), .ZN(new_n459));
  AOI21_X1  g0259(.A(new_n253), .B1(new_n458), .B2(new_n459), .ZN(new_n460));
  AOI21_X1  g0260(.A(KEYINPUT5), .B1(new_n265), .B2(new_n267), .ZN(new_n461));
  INV_X1    g0261(.A(KEYINPUT5), .ZN(new_n462));
  OAI211_X1 g0262(.A(new_n207), .B(G45), .C1(new_n462), .C2(G41), .ZN(new_n463));
  INV_X1    g0263(.A(G274), .ZN(new_n464));
  NOR4_X1   g0264(.A1(new_n461), .A2(new_n344), .A3(new_n463), .A4(new_n464), .ZN(new_n465));
  INV_X1    g0265(.A(new_n465), .ZN(new_n466));
  INV_X1    g0266(.A(G270), .ZN(new_n467));
  OAI21_X1  g0267(.A(new_n253), .B1(new_n461), .B2(new_n463), .ZN(new_n468));
  OAI21_X1  g0268(.A(new_n466), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  NOR2_X1   g0269(.A1(new_n460), .A2(new_n469), .ZN(new_n470));
  NOR2_X1   g0270(.A1(new_n470), .A2(new_n444), .ZN(new_n471));
  INV_X1    g0271(.A(G116), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n321), .A2(new_n472), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n207), .A2(G33), .ZN(new_n474));
  NAND4_X1  g0274(.A1(new_n320), .A2(G116), .A3(new_n280), .A4(new_n474), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n473), .A2(new_n475), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n209), .A2(G33), .ZN(new_n477));
  AOI22_X1  g0277(.A1(new_n477), .A2(new_n214), .B1(G20), .B2(new_n472), .ZN(new_n478));
  AOI21_X1  g0278(.A(G20), .B1(new_n251), .B2(G97), .ZN(new_n479));
  INV_X1    g0279(.A(G283), .ZN(new_n480));
  OAI21_X1  g0280(.A(new_n479), .B1(new_n251), .B2(new_n480), .ZN(new_n481));
  AOI21_X1  g0281(.A(KEYINPUT20), .B1(new_n478), .B2(new_n481), .ZN(new_n482));
  NAND3_X1  g0282(.A1(new_n478), .A2(KEYINPUT20), .A3(new_n481), .ZN(new_n483));
  AOI21_X1  g0283(.A(new_n482), .B1(new_n483), .B2(KEYINPUT90), .ZN(new_n484));
  OR2_X1    g0284(.A1(new_n483), .A2(KEYINPUT90), .ZN(new_n485));
  AOI21_X1  g0285(.A(new_n476), .B1(new_n484), .B2(new_n485), .ZN(new_n486));
  INV_X1    g0286(.A(new_n486), .ZN(new_n487));
  NOR3_X1   g0287(.A1(new_n460), .A2(new_n469), .A3(new_n358), .ZN(new_n488));
  NOR3_X1   g0288(.A1(new_n471), .A2(new_n487), .A3(new_n488), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n223), .A2(new_n259), .ZN(new_n490));
  OAI211_X1 g0290(.A(new_n456), .B(new_n490), .C1(G257), .C2(new_n259), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n419), .A2(G294), .ZN(new_n492));
  AOI21_X1  g0292(.A(new_n253), .B1(new_n491), .B2(new_n492), .ZN(new_n493));
  INV_X1    g0293(.A(new_n468), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n494), .A2(G264), .ZN(new_n495));
  INV_X1    g0295(.A(new_n495), .ZN(new_n496));
  NOR4_X1   g0296(.A1(new_n493), .A2(new_n496), .A3(new_n358), .A4(new_n465), .ZN(new_n497));
  NOR3_X1   g0297(.A1(new_n493), .A2(new_n465), .A3(new_n496), .ZN(new_n498));
  INV_X1    g0298(.A(new_n498), .ZN(new_n499));
  AOI21_X1  g0299(.A(new_n497), .B1(new_n499), .B2(G200), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n294), .A2(new_n375), .ZN(new_n501));
  OR2_X1    g0301(.A1(new_n501), .A2(KEYINPUT25), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n501), .A2(KEYINPUT25), .ZN(new_n503));
  NAND3_X1  g0303(.A1(new_n280), .A2(new_n293), .A3(new_n474), .ZN(new_n504));
  OAI211_X1 g0304(.A(new_n502), .B(new_n503), .C1(new_n504), .C2(new_n375), .ZN(new_n505));
  INV_X1    g0305(.A(KEYINPUT23), .ZN(new_n506));
  NAND3_X1  g0306(.A1(new_n506), .A2(new_n375), .A3(G20), .ZN(new_n507));
  XNOR2_X1  g0307(.A(new_n507), .B(KEYINPUT92), .ZN(new_n508));
  INV_X1    g0308(.A(KEYINPUT22), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n208), .A2(G87), .ZN(new_n510));
  OAI21_X1  g0310(.A(new_n509), .B1(new_n257), .B2(new_n510), .ZN(new_n511));
  NAND2_X1  g0311(.A1(KEYINPUT23), .A2(G107), .ZN(new_n512));
  AND3_X1   g0312(.A1(new_n508), .A2(new_n511), .A3(new_n512), .ZN(new_n513));
  NAND4_X1  g0313(.A1(new_n456), .A2(KEYINPUT22), .A3(new_n208), .A4(G87), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n419), .A2(G116), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n515), .A2(new_n506), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n516), .A2(new_n208), .ZN(new_n517));
  NAND3_X1  g0317(.A1(new_n513), .A2(new_n514), .A3(new_n517), .ZN(new_n518));
  XNOR2_X1  g0318(.A(new_n518), .B(KEYINPUT24), .ZN(new_n519));
  AOI21_X1  g0319(.A(new_n505), .B1(new_n519), .B2(new_n322), .ZN(new_n520));
  AOI21_X1  g0320(.A(new_n489), .B1(new_n500), .B2(new_n520), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n519), .A2(new_n322), .ZN(new_n522));
  INV_X1    g0322(.A(new_n505), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n499), .A2(new_n312), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n498), .A2(new_n314), .ZN(new_n526));
  NAND3_X1  g0326(.A1(new_n524), .A2(new_n525), .A3(new_n526), .ZN(new_n527));
  INV_X1    g0327(.A(KEYINPUT91), .ZN(new_n528));
  INV_X1    g0328(.A(KEYINPUT21), .ZN(new_n529));
  OAI21_X1  g0329(.A(G169), .B1(new_n460), .B2(new_n469), .ZN(new_n530));
  OAI211_X1 g0330(.A(new_n528), .B(new_n529), .C1(new_n486), .C2(new_n530), .ZN(new_n531));
  OAI21_X1  g0331(.A(new_n528), .B1(new_n486), .B2(new_n530), .ZN(new_n532));
  NOR3_X1   g0332(.A1(new_n460), .A2(new_n469), .A3(new_n314), .ZN(new_n533));
  AOI22_X1  g0333(.A1(new_n532), .A2(KEYINPUT21), .B1(new_n487), .B2(new_n533), .ZN(new_n534));
  NAND4_X1  g0334(.A1(new_n521), .A2(new_n527), .A3(new_n531), .A4(new_n534), .ZN(new_n535));
  AOI21_X1  g0335(.A(G33), .B1(new_n402), .B2(new_n404), .ZN(new_n536));
  AOI21_X1  g0336(.A(KEYINPUT3), .B1(new_n398), .B2(new_n400), .ZN(new_n537));
  OAI211_X1 g0337(.A(KEYINPUT7), .B(new_n208), .C1(new_n536), .C2(new_n537), .ZN(new_n538));
  INV_X1    g0338(.A(new_n422), .ZN(new_n539));
  AOI21_X1  g0339(.A(new_n375), .B1(new_n538), .B2(new_n539), .ZN(new_n540));
  INV_X1    g0340(.A(KEYINPUT6), .ZN(new_n541));
  NOR3_X1   g0341(.A1(new_n541), .A2(new_n342), .A3(G107), .ZN(new_n542));
  XNOR2_X1  g0342(.A(G97), .B(G107), .ZN(new_n543));
  AOI21_X1  g0343(.A(new_n542), .B1(new_n543), .B2(new_n541), .ZN(new_n544));
  OAI22_X1  g0344(.A1(new_n544), .A2(new_n208), .B1(new_n220), .B2(new_n364), .ZN(new_n545));
  OAI21_X1  g0345(.A(new_n322), .B1(new_n540), .B2(new_n545), .ZN(new_n546));
  INV_X1    g0346(.A(KEYINPUT85), .ZN(new_n547));
  NOR2_X1   g0347(.A1(new_n293), .A2(G97), .ZN(new_n548));
  INV_X1    g0348(.A(new_n504), .ZN(new_n549));
  AOI21_X1  g0349(.A(new_n548), .B1(new_n549), .B2(G97), .ZN(new_n550));
  NAND3_X1  g0350(.A1(new_n546), .A2(new_n547), .A3(new_n550), .ZN(new_n551));
  INV_X1    g0351(.A(new_n551), .ZN(new_n552));
  AOI21_X1  g0352(.A(new_n547), .B1(new_n546), .B2(new_n550), .ZN(new_n553));
  NOR2_X1   g0353(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  INV_X1    g0354(.A(KEYINPUT4), .ZN(new_n555));
  NOR3_X1   g0355(.A1(new_n555), .A2(new_n221), .A3(G1698), .ZN(new_n556));
  AOI22_X1  g0356(.A1(new_n258), .A2(new_n556), .B1(G33), .B2(G283), .ZN(new_n557));
  AOI21_X1  g0357(.A(new_n555), .B1(new_n258), .B2(G250), .ZN(new_n558));
  OAI21_X1  g0358(.A(new_n557), .B1(new_n558), .B2(new_n259), .ZN(new_n559));
  AOI21_X1  g0359(.A(KEYINPUT4), .B1(new_n456), .B2(G244), .ZN(new_n560));
  OAI21_X1  g0360(.A(new_n344), .B1(new_n559), .B2(new_n560), .ZN(new_n561));
  AOI21_X1  g0361(.A(new_n465), .B1(new_n494), .B2(G257), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n563), .A2(G200), .ZN(new_n564));
  AND2_X1   g0364(.A1(new_n561), .A2(new_n562), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n565), .A2(G190), .ZN(new_n566));
  NAND3_X1  g0366(.A1(new_n554), .A2(new_n564), .A3(new_n566), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n221), .A2(G1698), .ZN(new_n568));
  OAI211_X1 g0368(.A(new_n456), .B(new_n568), .C1(G238), .C2(G1698), .ZN(new_n569));
  AOI21_X1  g0369(.A(new_n253), .B1(new_n569), .B2(new_n515), .ZN(new_n570));
  INV_X1    g0370(.A(G45), .ZN(new_n571));
  OAI21_X1  g0371(.A(new_n223), .B1(new_n571), .B2(G1), .ZN(new_n572));
  NAND3_X1  g0372(.A1(new_n207), .A2(new_n464), .A3(G45), .ZN(new_n573));
  AND3_X1   g0373(.A1(new_n253), .A2(new_n572), .A3(new_n573), .ZN(new_n574));
  OAI21_X1  g0374(.A(new_n277), .B1(new_n570), .B2(new_n574), .ZN(new_n575));
  NAND3_X1  g0375(.A1(new_n456), .A2(new_n208), .A3(G68), .ZN(new_n576));
  NOR3_X1   g0376(.A1(G87), .A2(G97), .A3(G107), .ZN(new_n577));
  XNOR2_X1  g0377(.A(new_n577), .B(KEYINPUT87), .ZN(new_n578));
  OAI21_X1  g0378(.A(new_n208), .B1(new_n251), .B2(new_n342), .ZN(new_n579));
  NAND3_X1  g0379(.A1(new_n578), .A2(KEYINPUT19), .A3(new_n579), .ZN(new_n580));
  NOR2_X1   g0380(.A1(new_n287), .A2(new_n342), .ZN(new_n581));
  OAI211_X1 g0381(.A(new_n576), .B(new_n580), .C1(KEYINPUT19), .C2(new_n581), .ZN(new_n582));
  AOI22_X1  g0382(.A1(new_n582), .A2(new_n322), .B1(new_n321), .B2(new_n365), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n549), .A2(G87), .ZN(new_n584));
  NAND3_X1  g0384(.A1(new_n575), .A2(new_n583), .A3(new_n584), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n585), .A2(KEYINPUT88), .ZN(new_n586));
  INV_X1    g0386(.A(KEYINPUT88), .ZN(new_n587));
  NAND4_X1  g0387(.A1(new_n575), .A2(new_n583), .A3(new_n587), .A4(new_n584), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n569), .A2(new_n515), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n589), .A2(new_n344), .ZN(new_n590));
  INV_X1    g0390(.A(new_n574), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  NOR2_X1   g0392(.A1(new_n592), .A2(new_n358), .ZN(new_n593));
  INV_X1    g0393(.A(new_n593), .ZN(new_n594));
  NAND3_X1  g0394(.A1(new_n586), .A2(new_n588), .A3(new_n594), .ZN(new_n595));
  NOR2_X1   g0395(.A1(new_n570), .A2(new_n574), .ZN(new_n596));
  AOI21_X1  g0396(.A(KEYINPUT86), .B1(new_n596), .B2(new_n314), .ZN(new_n597));
  INV_X1    g0397(.A(KEYINPUT86), .ZN(new_n598));
  NOR4_X1   g0398(.A1(new_n570), .A2(new_n598), .A3(G179), .A4(new_n574), .ZN(new_n599));
  NOR2_X1   g0399(.A1(new_n597), .A2(new_n599), .ZN(new_n600));
  INV_X1    g0400(.A(new_n365), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n549), .A2(new_n601), .ZN(new_n602));
  AOI22_X1  g0402(.A1(new_n592), .A2(new_n312), .B1(new_n583), .B2(new_n602), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n600), .A2(new_n603), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n563), .A2(G169), .ZN(new_n605));
  OAI21_X1  g0405(.A(new_n605), .B1(new_n314), .B2(new_n563), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n546), .A2(new_n550), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  NAND4_X1  g0408(.A1(new_n567), .A2(new_n595), .A3(new_n604), .A4(new_n608), .ZN(new_n609));
  INV_X1    g0409(.A(KEYINPUT89), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  AOI21_X1  g0411(.A(new_n593), .B1(new_n585), .B2(KEYINPUT88), .ZN(new_n612));
  AOI22_X1  g0412(.A1(new_n612), .A2(new_n588), .B1(new_n600), .B2(new_n603), .ZN(new_n613));
  NAND4_X1  g0413(.A1(new_n613), .A2(KEYINPUT89), .A3(new_n608), .A4(new_n567), .ZN(new_n614));
  AOI21_X1  g0414(.A(new_n535), .B1(new_n611), .B2(new_n614), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n455), .A2(new_n615), .ZN(new_n616));
  XOR2_X1   g0416(.A(new_n616), .B(KEYINPUT93), .Z(G372));
  NAND2_X1  g0417(.A1(new_n534), .A2(new_n531), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n525), .A2(new_n526), .ZN(new_n619));
  NOR2_X1   g0419(.A1(new_n619), .A2(new_n520), .ZN(new_n620));
  NOR2_X1   g0420(.A1(new_n618), .A2(new_n620), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n520), .A2(new_n500), .ZN(new_n622));
  OR2_X1    g0422(.A1(new_n585), .A2(new_n593), .ZN(new_n623));
  NAND4_X1  g0423(.A1(new_n567), .A2(new_n622), .A3(new_n608), .A4(new_n623), .ZN(new_n624));
  NOR2_X1   g0424(.A1(new_n621), .A2(new_n624), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n596), .A2(new_n314), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n603), .A2(new_n626), .ZN(new_n627));
  OR2_X1    g0427(.A1(new_n552), .A2(new_n553), .ZN(new_n628));
  NAND3_X1  g0428(.A1(new_n623), .A2(new_n606), .A3(new_n628), .ZN(new_n629));
  OAI21_X1  g0429(.A(new_n627), .B1(new_n629), .B2(KEYINPUT26), .ZN(new_n630));
  INV_X1    g0430(.A(new_n630), .ZN(new_n631));
  INV_X1    g0431(.A(new_n608), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n613), .A2(new_n632), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n633), .A2(KEYINPUT26), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n631), .A2(new_n634), .ZN(new_n635));
  OAI21_X1  g0435(.A(new_n455), .B1(new_n625), .B2(new_n635), .ZN(new_n636));
  INV_X1    g0436(.A(new_n316), .ZN(new_n637));
  INV_X1    g0437(.A(new_n355), .ZN(new_n638));
  INV_X1    g0438(.A(new_n386), .ZN(new_n639));
  AOI21_X1  g0439(.A(new_n638), .B1(new_n359), .B2(new_n639), .ZN(new_n640));
  INV_X1    g0440(.A(new_n453), .ZN(new_n641));
  OAI21_X1  g0441(.A(new_n442), .B1(new_n640), .B2(new_n641), .ZN(new_n642));
  AOI21_X1  g0442(.A(new_n637), .B1(new_n642), .B2(new_n311), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n636), .A2(new_n643), .ZN(G369));
  INV_X1    g0444(.A(G13), .ZN(new_n645));
  NOR3_X1   g0445(.A1(new_n645), .A2(G1), .A3(G20), .ZN(new_n646));
  INV_X1    g0446(.A(new_n646), .ZN(new_n647));
  INV_X1    g0447(.A(KEYINPUT94), .ZN(new_n648));
  AND3_X1   g0448(.A1(new_n647), .A2(new_n648), .A3(KEYINPUT27), .ZN(new_n649));
  AOI21_X1  g0449(.A(new_n648), .B1(new_n647), .B2(KEYINPUT27), .ZN(new_n650));
  OAI221_X1 g0450(.A(G213), .B1(KEYINPUT27), .B2(new_n647), .C1(new_n649), .C2(new_n650), .ZN(new_n651));
  INV_X1    g0451(.A(G343), .ZN(new_n652));
  NOR2_X1   g0452(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  INV_X1    g0453(.A(new_n653), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n620), .A2(new_n654), .ZN(new_n655));
  INV_X1    g0455(.A(new_n655), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n524), .A2(new_n653), .ZN(new_n657));
  INV_X1    g0457(.A(new_n619), .ZN(new_n658));
  AOI22_X1  g0458(.A1(new_n657), .A2(new_n622), .B1(new_n658), .B2(new_n524), .ZN(new_n659));
  NOR2_X1   g0459(.A1(new_n656), .A2(new_n659), .ZN(new_n660));
  NOR2_X1   g0460(.A1(new_n486), .A2(new_n654), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n618), .A2(new_n661), .ZN(new_n662));
  OAI211_X1 g0462(.A(new_n534), .B(new_n531), .C1(new_n486), .C2(new_n654), .ZN(new_n663));
  AOI21_X1  g0463(.A(new_n489), .B1(new_n662), .B2(new_n663), .ZN(new_n664));
  NAND3_X1  g0464(.A1(new_n664), .A2(KEYINPUT95), .A3(G330), .ZN(new_n665));
  INV_X1    g0465(.A(new_n665), .ZN(new_n666));
  AOI21_X1  g0466(.A(KEYINPUT95), .B1(new_n664), .B2(G330), .ZN(new_n667));
  OAI21_X1  g0467(.A(new_n660), .B1(new_n666), .B2(new_n667), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n618), .A2(new_n654), .ZN(new_n669));
  OAI21_X1  g0469(.A(new_n655), .B1(new_n659), .B2(new_n669), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n670), .A2(KEYINPUT96), .ZN(new_n671));
  INV_X1    g0471(.A(KEYINPUT96), .ZN(new_n672));
  OAI211_X1 g0472(.A(new_n672), .B(new_n655), .C1(new_n659), .C2(new_n669), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n671), .A2(new_n673), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n668), .A2(new_n674), .ZN(G399));
  INV_X1    g0475(.A(new_n211), .ZN(new_n676));
  NOR2_X1   g0476(.A1(new_n676), .A2(new_n268), .ZN(new_n677));
  INV_X1    g0477(.A(new_n677), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n678), .A2(G1), .ZN(new_n679));
  OR2_X1    g0479(.A1(new_n578), .A2(G116), .ZN(new_n680));
  OAI22_X1  g0480(.A1(new_n679), .A2(new_n680), .B1(new_n218), .B2(new_n678), .ZN(new_n681));
  XNOR2_X1  g0481(.A(new_n681), .B(KEYINPUT28), .ZN(new_n682));
  NOR3_X1   g0482(.A1(new_n470), .A2(new_n596), .A3(G179), .ZN(new_n683));
  NAND3_X1  g0483(.A1(new_n683), .A2(new_n563), .A3(new_n499), .ZN(new_n684));
  INV_X1    g0484(.A(KEYINPUT30), .ZN(new_n685));
  NOR2_X1   g0485(.A1(new_n493), .A2(new_n496), .ZN(new_n686));
  NAND3_X1  g0486(.A1(new_n533), .A2(new_n596), .A3(new_n686), .ZN(new_n687));
  OAI21_X1  g0487(.A(new_n685), .B1(new_n687), .B2(new_n563), .ZN(new_n688));
  AND2_X1   g0488(.A1(new_n686), .A2(new_n596), .ZN(new_n689));
  NAND4_X1  g0489(.A1(new_n689), .A2(KEYINPUT30), .A3(new_n565), .A4(new_n533), .ZN(new_n690));
  NAND3_X1  g0490(.A1(new_n684), .A2(new_n688), .A3(new_n690), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n691), .A2(new_n653), .ZN(new_n692));
  INV_X1    g0492(.A(KEYINPUT31), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  NAND3_X1  g0494(.A1(new_n691), .A2(KEYINPUT31), .A3(new_n653), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  AOI21_X1  g0496(.A(new_n696), .B1(new_n615), .B2(new_n654), .ZN(new_n697));
  INV_X1    g0497(.A(G330), .ZN(new_n698));
  NOR2_X1   g0498(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  OAI21_X1  g0499(.A(new_n654), .B1(new_n635), .B2(new_n625), .ZN(new_n700));
  INV_X1    g0500(.A(KEYINPUT29), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  INV_X1    g0502(.A(KEYINPUT97), .ZN(new_n703));
  INV_X1    g0503(.A(new_n627), .ZN(new_n704));
  AOI21_X1  g0504(.A(new_n704), .B1(new_n629), .B2(KEYINPUT26), .ZN(new_n705));
  INV_X1    g0505(.A(KEYINPUT26), .ZN(new_n706));
  NAND3_X1  g0506(.A1(new_n613), .A2(new_n706), .A3(new_n632), .ZN(new_n707));
  OAI211_X1 g0507(.A(new_n705), .B(new_n707), .C1(new_n621), .C2(new_n624), .ZN(new_n708));
  AND2_X1   g0508(.A1(new_n708), .A2(new_n654), .ZN(new_n709));
  AOI22_X1  g0509(.A1(new_n702), .A2(new_n703), .B1(KEYINPUT29), .B2(new_n709), .ZN(new_n710));
  NAND3_X1  g0510(.A1(new_n700), .A2(KEYINPUT97), .A3(new_n701), .ZN(new_n711));
  AOI21_X1  g0511(.A(new_n699), .B1(new_n710), .B2(new_n711), .ZN(new_n712));
  OAI21_X1  g0512(.A(new_n682), .B1(new_n712), .B2(G1), .ZN(G364));
  NOR2_X1   g0513(.A1(new_n666), .A2(new_n667), .ZN(new_n714));
  NOR2_X1   g0514(.A1(new_n645), .A2(G20), .ZN(new_n715));
  AOI21_X1  g0515(.A(new_n207), .B1(new_n715), .B2(G45), .ZN(new_n716));
  INV_X1    g0516(.A(new_n716), .ZN(new_n717));
  NOR2_X1   g0517(.A1(new_n677), .A2(new_n717), .ZN(new_n718));
  INV_X1    g0518(.A(new_n718), .ZN(new_n719));
  OAI211_X1 g0519(.A(new_n714), .B(new_n719), .C1(G330), .C2(new_n664), .ZN(new_n720));
  AOI21_X1  g0520(.A(new_n214), .B1(G20), .B2(new_n312), .ZN(new_n721));
  NOR2_X1   g0521(.A1(G179), .A2(G200), .ZN(new_n722));
  AOI21_X1  g0522(.A(new_n208), .B1(new_n722), .B2(G190), .ZN(new_n723));
  INV_X1    g0523(.A(new_n723), .ZN(new_n724));
  NAND3_X1  g0524(.A1(G20), .A2(G179), .A3(G200), .ZN(new_n725));
  NOR2_X1   g0525(.A1(new_n725), .A2(new_n358), .ZN(new_n726));
  AOI22_X1  g0526(.A1(new_n724), .A2(G294), .B1(G326), .B2(new_n726), .ZN(new_n727));
  NOR2_X1   g0527(.A1(new_n725), .A2(G190), .ZN(new_n728));
  INV_X1    g0528(.A(new_n728), .ZN(new_n729));
  XOR2_X1   g0529(.A(KEYINPUT33), .B(G317), .Z(new_n730));
  OAI21_X1  g0530(.A(new_n727), .B1(new_n729), .B2(new_n730), .ZN(new_n731));
  NOR2_X1   g0531(.A1(new_n314), .A2(G200), .ZN(new_n732));
  NAND3_X1  g0532(.A1(new_n732), .A2(G20), .A3(G190), .ZN(new_n733));
  INV_X1    g0533(.A(G322), .ZN(new_n734));
  NOR2_X1   g0534(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  NOR2_X1   g0535(.A1(new_n208), .A2(G190), .ZN(new_n736));
  NAND2_X1  g0536(.A1(new_n736), .A2(new_n722), .ZN(new_n737));
  INV_X1    g0537(.A(new_n737), .ZN(new_n738));
  AOI21_X1  g0538(.A(new_n735), .B1(G329), .B2(new_n738), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n736), .A2(new_n732), .ZN(new_n740));
  INV_X1    g0540(.A(new_n740), .ZN(new_n741));
  AOI21_X1  g0541(.A(new_n258), .B1(new_n741), .B2(G311), .ZN(new_n742));
  INV_X1    g0542(.A(G303), .ZN(new_n743));
  NOR2_X1   g0543(.A1(new_n208), .A2(G179), .ZN(new_n744));
  NAND3_X1  g0544(.A1(new_n277), .A2(G190), .A3(new_n744), .ZN(new_n745));
  OAI211_X1 g0545(.A(new_n739), .B(new_n742), .C1(new_n743), .C2(new_n745), .ZN(new_n746));
  NAND3_X1  g0546(.A1(new_n277), .A2(new_n358), .A3(new_n744), .ZN(new_n747));
  INV_X1    g0547(.A(new_n747), .ZN(new_n748));
  AOI211_X1 g0548(.A(new_n731), .B(new_n746), .C1(G283), .C2(new_n748), .ZN(new_n749));
  INV_X1    g0549(.A(new_n745), .ZN(new_n750));
  NAND2_X1  g0550(.A1(new_n750), .A2(G87), .ZN(new_n751));
  NAND2_X1  g0551(.A1(new_n748), .A2(G107), .ZN(new_n752));
  NAND2_X1  g0552(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  INV_X1    g0553(.A(G159), .ZN(new_n754));
  OR3_X1    g0554(.A1(new_n737), .A2(KEYINPUT32), .A3(new_n754), .ZN(new_n755));
  OAI21_X1  g0555(.A(KEYINPUT32), .B1(new_n737), .B2(new_n754), .ZN(new_n756));
  OAI211_X1 g0556(.A(new_n755), .B(new_n756), .C1(new_n342), .C2(new_n723), .ZN(new_n757));
  OAI221_X1 g0557(.A(new_n258), .B1(new_n740), .B2(new_n220), .C1(new_n202), .C2(new_n733), .ZN(new_n758));
  INV_X1    g0558(.A(new_n726), .ZN(new_n759));
  OAI22_X1  g0559(.A1(new_n729), .A2(new_n203), .B1(new_n759), .B2(new_n201), .ZN(new_n760));
  NOR4_X1   g0560(.A1(new_n753), .A2(new_n757), .A3(new_n758), .A4(new_n760), .ZN(new_n761));
  OAI21_X1  g0561(.A(new_n721), .B1(new_n749), .B2(new_n761), .ZN(new_n762));
  NAND2_X1  g0562(.A1(new_n211), .A2(new_n258), .ZN(new_n763));
  XNOR2_X1  g0563(.A(new_n763), .B(KEYINPUT98), .ZN(new_n764));
  AOI22_X1  g0564(.A1(new_n764), .A2(G355), .B1(new_n472), .B2(new_n676), .ZN(new_n765));
  NOR2_X1   g0565(.A1(new_n246), .A2(new_n571), .ZN(new_n766));
  NOR2_X1   g0566(.A1(new_n676), .A2(new_n456), .ZN(new_n767));
  OAI21_X1  g0567(.A(new_n767), .B1(G45), .B2(new_n218), .ZN(new_n768));
  OAI21_X1  g0568(.A(new_n765), .B1(new_n766), .B2(new_n768), .ZN(new_n769));
  NOR2_X1   g0569(.A1(G13), .A2(G33), .ZN(new_n770));
  INV_X1    g0570(.A(new_n770), .ZN(new_n771));
  NOR2_X1   g0571(.A1(new_n771), .A2(G20), .ZN(new_n772));
  NOR2_X1   g0572(.A1(new_n772), .A2(new_n721), .ZN(new_n773));
  AOI21_X1  g0573(.A(new_n719), .B1(new_n769), .B2(new_n773), .ZN(new_n774));
  INV_X1    g0574(.A(new_n772), .ZN(new_n775));
  OAI211_X1 g0575(.A(new_n762), .B(new_n774), .C1(new_n664), .C2(new_n775), .ZN(new_n776));
  AND2_X1   g0576(.A1(new_n720), .A2(new_n776), .ZN(new_n777));
  INV_X1    g0577(.A(new_n777), .ZN(G396));
  NOR2_X1   g0578(.A1(new_n386), .A2(new_n653), .ZN(new_n779));
  NAND2_X1  g0579(.A1(new_n385), .A2(new_n653), .ZN(new_n780));
  NAND2_X1  g0580(.A1(new_n382), .A2(new_n780), .ZN(new_n781));
  AOI21_X1  g0581(.A(new_n779), .B1(new_n781), .B2(new_n386), .ZN(new_n782));
  INV_X1    g0582(.A(new_n782), .ZN(new_n783));
  NOR2_X1   g0583(.A1(new_n700), .A2(new_n783), .ZN(new_n784));
  INV_X1    g0584(.A(new_n784), .ZN(new_n785));
  NAND2_X1  g0585(.A1(new_n700), .A2(new_n783), .ZN(new_n786));
  NAND2_X1  g0586(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  INV_X1    g0587(.A(new_n697), .ZN(new_n788));
  NAND2_X1  g0588(.A1(new_n788), .A2(G330), .ZN(new_n789));
  AOI21_X1  g0589(.A(new_n718), .B1(new_n787), .B2(new_n789), .ZN(new_n790));
  OAI21_X1  g0590(.A(new_n790), .B1(new_n789), .B2(new_n787), .ZN(new_n791));
  NOR2_X1   g0591(.A1(new_n721), .A2(new_n770), .ZN(new_n792));
  AOI21_X1  g0592(.A(new_n719), .B1(new_n220), .B2(new_n792), .ZN(new_n793));
  INV_X1    g0593(.A(new_n721), .ZN(new_n794));
  INV_X1    g0594(.A(new_n733), .ZN(new_n795));
  AOI22_X1  g0595(.A1(new_n795), .A2(G143), .B1(new_n741), .B2(G159), .ZN(new_n796));
  INV_X1    g0596(.A(G150), .ZN(new_n797));
  INV_X1    g0597(.A(G137), .ZN(new_n798));
  OAI221_X1 g0598(.A(new_n796), .B1(new_n729), .B2(new_n797), .C1(new_n798), .C2(new_n759), .ZN(new_n799));
  XNOR2_X1  g0599(.A(new_n799), .B(KEYINPUT34), .ZN(new_n800));
  NOR2_X1   g0600(.A1(new_n747), .A2(new_n203), .ZN(new_n801));
  NAND2_X1  g0601(.A1(new_n401), .A2(new_n405), .ZN(new_n802));
  AOI21_X1  g0602(.A(new_n802), .B1(G132), .B2(new_n738), .ZN(new_n803));
  OAI21_X1  g0603(.A(new_n803), .B1(new_n202), .B2(new_n723), .ZN(new_n804));
  AOI211_X1 g0604(.A(new_n801), .B(new_n804), .C1(G50), .C2(new_n750), .ZN(new_n805));
  NOR2_X1   g0605(.A1(new_n747), .A2(new_n222), .ZN(new_n806));
  AOI22_X1  g0606(.A1(new_n741), .A2(G116), .B1(new_n738), .B2(G311), .ZN(new_n807));
  INV_X1    g0607(.A(G294), .ZN(new_n808));
  OAI211_X1 g0608(.A(new_n807), .B(new_n257), .C1(new_n808), .C2(new_n733), .ZN(new_n809));
  AOI211_X1 g0609(.A(new_n806), .B(new_n809), .C1(G107), .C2(new_n750), .ZN(new_n810));
  OAI22_X1  g0610(.A1(new_n729), .A2(new_n480), .B1(new_n723), .B2(new_n342), .ZN(new_n811));
  AOI21_X1  g0611(.A(new_n811), .B1(G303), .B2(new_n726), .ZN(new_n812));
  AOI22_X1  g0612(.A1(new_n800), .A2(new_n805), .B1(new_n810), .B2(new_n812), .ZN(new_n813));
  OAI221_X1 g0613(.A(new_n793), .B1(new_n794), .B2(new_n813), .C1(new_n782), .C2(new_n771), .ZN(new_n814));
  AND2_X1   g0614(.A1(new_n791), .A2(new_n814), .ZN(new_n815));
  INV_X1    g0615(.A(new_n815), .ZN(G384));
  NOR2_X1   g0616(.A1(new_n715), .A2(new_n207), .ZN(new_n817));
  INV_X1    g0617(.A(new_n412), .ZN(new_n818));
  NAND3_X1  g0618(.A1(new_n802), .A2(new_n208), .A3(new_n818), .ZN(new_n819));
  OAI211_X1 g0619(.A(new_n819), .B(G68), .C1(new_n407), .C2(new_n406), .ZN(new_n820));
  AOI21_X1  g0620(.A(KEYINPUT16), .B1(new_n820), .B2(new_n424), .ZN(new_n821));
  OAI21_X1  g0621(.A(new_n390), .B1(new_n415), .B2(new_n821), .ZN(new_n822));
  INV_X1    g0622(.A(new_n651), .ZN(new_n823));
  NAND2_X1  g0623(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  AOI21_X1  g0624(.A(new_n824), .B1(new_n442), .B2(new_n453), .ZN(new_n825));
  INV_X1    g0625(.A(new_n825), .ZN(new_n826));
  AOI21_X1  g0626(.A(new_n280), .B1(new_n820), .B2(new_n397), .ZN(new_n827));
  AOI21_X1  g0627(.A(new_n203), .B1(new_n538), .B2(new_n539), .ZN(new_n828));
  OAI21_X1  g0628(.A(new_n396), .B1(new_n828), .B2(new_n395), .ZN(new_n829));
  AOI21_X1  g0629(.A(new_n389), .B1(new_n827), .B2(new_n829), .ZN(new_n830));
  INV_X1    g0630(.A(new_n439), .ZN(new_n831));
  OAI21_X1  g0631(.A(new_n447), .B1(new_n830), .B2(new_n831), .ZN(new_n832));
  NOR2_X1   g0632(.A1(new_n830), .A2(new_n651), .ZN(new_n833));
  NOR3_X1   g0633(.A1(new_n832), .A2(new_n833), .A3(KEYINPUT37), .ZN(new_n834));
  INV_X1    g0634(.A(KEYINPUT101), .ZN(new_n835));
  OAI21_X1  g0635(.A(new_n424), .B1(new_n408), .B2(new_n413), .ZN(new_n836));
  NAND2_X1  g0636(.A1(new_n836), .A2(new_n396), .ZN(new_n837));
  AOI21_X1  g0637(.A(new_n389), .B1(new_n837), .B2(new_n827), .ZN(new_n838));
  NAND3_X1  g0638(.A1(new_n436), .A2(new_n438), .A3(new_n651), .ZN(new_n839));
  INV_X1    g0639(.A(new_n839), .ZN(new_n840));
  OAI21_X1  g0640(.A(new_n447), .B1(new_n838), .B2(new_n840), .ZN(new_n841));
  AOI21_X1  g0641(.A(new_n835), .B1(new_n841), .B2(KEYINPUT37), .ZN(new_n842));
  NOR2_X1   g0642(.A1(new_n834), .A2(new_n842), .ZN(new_n843));
  NAND3_X1  g0643(.A1(new_n841), .A2(new_n835), .A3(KEYINPUT37), .ZN(new_n844));
  AOI21_X1  g0644(.A(KEYINPUT102), .B1(new_n843), .B2(new_n844), .ZN(new_n845));
  AOI22_X1  g0645(.A1(new_n822), .A2(new_n839), .B1(new_n830), .B2(new_n446), .ZN(new_n846));
  INV_X1    g0646(.A(KEYINPUT37), .ZN(new_n847));
  OAI21_X1  g0647(.A(KEYINPUT101), .B1(new_n846), .B2(new_n847), .ZN(new_n848));
  NAND2_X1  g0648(.A1(new_n426), .A2(new_n823), .ZN(new_n849));
  NAND4_X1  g0649(.A1(new_n440), .A2(new_n849), .A3(new_n847), .A4(new_n447), .ZN(new_n850));
  NAND4_X1  g0650(.A1(new_n848), .A2(KEYINPUT102), .A3(new_n844), .A4(new_n850), .ZN(new_n851));
  INV_X1    g0651(.A(new_n851), .ZN(new_n852));
  OAI211_X1 g0652(.A(KEYINPUT38), .B(new_n826), .C1(new_n845), .C2(new_n852), .ZN(new_n853));
  NAND2_X1  g0653(.A1(new_n853), .A2(KEYINPUT105), .ZN(new_n854));
  INV_X1    g0654(.A(KEYINPUT39), .ZN(new_n855));
  INV_X1    g0655(.A(KEYINPUT102), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n822), .A2(new_n839), .ZN(new_n857));
  AOI21_X1  g0657(.A(new_n847), .B1(new_n857), .B2(new_n447), .ZN(new_n858));
  OAI21_X1  g0658(.A(new_n850), .B1(new_n858), .B2(new_n835), .ZN(new_n859));
  INV_X1    g0659(.A(new_n844), .ZN(new_n860));
  OAI21_X1  g0660(.A(new_n856), .B1(new_n859), .B2(new_n860), .ZN(new_n861));
  AOI21_X1  g0661(.A(new_n825), .B1(new_n861), .B2(new_n851), .ZN(new_n862));
  INV_X1    g0662(.A(KEYINPUT105), .ZN(new_n863));
  NAND3_X1  g0663(.A1(new_n862), .A2(new_n863), .A3(KEYINPUT38), .ZN(new_n864));
  INV_X1    g0664(.A(KEYINPUT38), .ZN(new_n865));
  AOI21_X1  g0665(.A(new_n849), .B1(new_n442), .B2(new_n453), .ZN(new_n866));
  OAI21_X1  g0666(.A(KEYINPUT37), .B1(new_n832), .B2(new_n833), .ZN(new_n867));
  AND2_X1   g0667(.A1(new_n867), .A2(new_n850), .ZN(new_n868));
  OAI21_X1  g0668(.A(new_n865), .B1(new_n866), .B2(new_n868), .ZN(new_n869));
  NAND4_X1  g0669(.A1(new_n854), .A2(new_n855), .A3(new_n864), .A4(new_n869), .ZN(new_n870));
  INV_X1    g0670(.A(KEYINPUT103), .ZN(new_n871));
  AOI21_X1  g0671(.A(new_n871), .B1(new_n862), .B2(KEYINPUT38), .ZN(new_n872));
  OAI21_X1  g0672(.A(new_n826), .B1(new_n845), .B2(new_n852), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n873), .A2(new_n865), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n872), .A2(new_n874), .ZN(new_n875));
  NOR3_X1   g0675(.A1(new_n862), .A2(KEYINPUT103), .A3(KEYINPUT38), .ZN(new_n876));
  INV_X1    g0676(.A(new_n876), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n875), .A2(new_n877), .ZN(new_n878));
  OAI21_X1  g0678(.A(new_n870), .B1(new_n878), .B2(new_n855), .ZN(new_n879));
  NAND3_X1  g0679(.A1(new_n879), .A2(new_n638), .A3(new_n654), .ZN(new_n880));
  INV_X1    g0680(.A(KEYINPUT104), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n853), .A2(KEYINPUT103), .ZN(new_n882));
  NOR2_X1   g0682(.A1(new_n862), .A2(KEYINPUT38), .ZN(new_n883));
  NOR2_X1   g0683(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  OAI21_X1  g0684(.A(new_n881), .B1(new_n884), .B2(new_n876), .ZN(new_n885));
  XNOR2_X1  g0685(.A(new_n779), .B(KEYINPUT99), .ZN(new_n886));
  AOI21_X1  g0686(.A(new_n630), .B1(KEYINPUT26), .B2(new_n633), .ZN(new_n887));
  INV_X1    g0687(.A(new_n625), .ZN(new_n888));
  AOI21_X1  g0688(.A(new_n653), .B1(new_n887), .B2(new_n888), .ZN(new_n889));
  AOI21_X1  g0689(.A(new_n886), .B1(new_n889), .B2(new_n782), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n334), .A2(new_n653), .ZN(new_n891));
  NAND3_X1  g0691(.A1(new_n355), .A2(new_n359), .A3(new_n891), .ZN(new_n892));
  INV_X1    g0692(.A(new_n891), .ZN(new_n893));
  OAI21_X1  g0693(.A(new_n893), .B1(new_n352), .B2(new_n354), .ZN(new_n894));
  INV_X1    g0694(.A(KEYINPUT100), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  OAI211_X1 g0696(.A(new_n893), .B(KEYINPUT100), .C1(new_n352), .C2(new_n354), .ZN(new_n897));
  NAND3_X1  g0697(.A1(new_n892), .A2(new_n896), .A3(new_n897), .ZN(new_n898));
  INV_X1    g0698(.A(new_n898), .ZN(new_n899));
  NOR2_X1   g0699(.A1(new_n890), .A2(new_n899), .ZN(new_n900));
  NAND3_X1  g0700(.A1(new_n875), .A2(new_n877), .A3(KEYINPUT104), .ZN(new_n901));
  NAND3_X1  g0701(.A1(new_n885), .A2(new_n900), .A3(new_n901), .ZN(new_n902));
  OR2_X1    g0702(.A1(new_n442), .A2(new_n823), .ZN(new_n903));
  NAND3_X1  g0703(.A1(new_n880), .A2(new_n902), .A3(new_n903), .ZN(new_n904));
  OAI21_X1  g0704(.A(new_n703), .B1(new_n889), .B2(KEYINPUT29), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n709), .A2(KEYINPUT29), .ZN(new_n906));
  NAND4_X1  g0706(.A1(new_n905), .A2(new_n711), .A3(new_n455), .A4(new_n906), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n907), .A2(new_n643), .ZN(new_n908));
  XNOR2_X1  g0708(.A(new_n904), .B(new_n908), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n898), .A2(new_n782), .ZN(new_n910));
  NOR2_X1   g0710(.A1(new_n697), .A2(new_n910), .ZN(new_n911));
  NAND3_X1  g0711(.A1(new_n885), .A2(new_n901), .A3(new_n911), .ZN(new_n912));
  INV_X1    g0712(.A(KEYINPUT40), .ZN(new_n913));
  NAND3_X1  g0713(.A1(new_n854), .A2(new_n864), .A3(new_n869), .ZN(new_n914));
  NOR3_X1   g0714(.A1(new_n697), .A2(new_n910), .A3(new_n913), .ZN(new_n915));
  AOI22_X1  g0715(.A1(new_n912), .A2(new_n913), .B1(new_n914), .B2(new_n915), .ZN(new_n916));
  AND2_X1   g0716(.A1(new_n455), .A2(new_n788), .ZN(new_n917));
  AOI21_X1  g0717(.A(new_n698), .B1(new_n916), .B2(new_n917), .ZN(new_n918));
  OAI21_X1  g0718(.A(new_n918), .B1(new_n916), .B2(new_n917), .ZN(new_n919));
  AOI21_X1  g0719(.A(new_n817), .B1(new_n909), .B2(new_n919), .ZN(new_n920));
  OAI21_X1  g0720(.A(new_n920), .B1(new_n909), .B2(new_n919), .ZN(new_n921));
  INV_X1    g0721(.A(new_n544), .ZN(new_n922));
  AOI211_X1 g0722(.A(new_n472), .B(new_n217), .C1(new_n922), .C2(KEYINPUT35), .ZN(new_n923));
  OAI21_X1  g0723(.A(new_n923), .B1(KEYINPUT35), .B2(new_n922), .ZN(new_n924));
  XNOR2_X1  g0724(.A(new_n924), .B(KEYINPUT36), .ZN(new_n925));
  NOR3_X1   g0725(.A1(new_n391), .A2(new_n218), .A3(new_n220), .ZN(new_n926));
  NOR2_X1   g0726(.A1(new_n203), .A2(G50), .ZN(new_n927));
  OAI211_X1 g0727(.A(G1), .B(new_n645), .C1(new_n926), .C2(new_n927), .ZN(new_n928));
  NAND3_X1  g0728(.A1(new_n921), .A2(new_n925), .A3(new_n928), .ZN(G367));
  NAND2_X1  g0729(.A1(new_n583), .A2(new_n584), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n930), .A2(new_n653), .ZN(new_n931));
  NAND3_X1  g0731(.A1(new_n623), .A2(new_n627), .A3(new_n931), .ZN(new_n932));
  OAI21_X1  g0732(.A(new_n932), .B1(new_n627), .B2(new_n931), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n933), .A2(KEYINPUT43), .ZN(new_n934));
  NOR2_X1   g0734(.A1(new_n554), .A2(new_n654), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n935), .A2(new_n606), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n936), .A2(KEYINPUT106), .ZN(new_n937));
  INV_X1    g0737(.A(KEYINPUT106), .ZN(new_n938));
  NAND3_X1  g0738(.A1(new_n935), .A2(new_n938), .A3(new_n606), .ZN(new_n939));
  OAI211_X1 g0739(.A(new_n567), .B(new_n608), .C1(new_n554), .C2(new_n654), .ZN(new_n940));
  NAND3_X1  g0740(.A1(new_n937), .A2(new_n939), .A3(new_n940), .ZN(new_n941));
  INV_X1    g0741(.A(new_n669), .ZN(new_n942));
  NAND3_X1  g0742(.A1(new_n660), .A2(new_n941), .A3(new_n942), .ZN(new_n943));
  XNOR2_X1  g0743(.A(new_n943), .B(KEYINPUT42), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n941), .A2(new_n620), .ZN(new_n945));
  AOI21_X1  g0745(.A(new_n653), .B1(new_n945), .B2(new_n608), .ZN(new_n946));
  OAI21_X1  g0746(.A(new_n934), .B1(new_n944), .B2(new_n946), .ZN(new_n947));
  NOR2_X1   g0747(.A1(new_n933), .A2(KEYINPUT43), .ZN(new_n948));
  XNOR2_X1  g0748(.A(new_n947), .B(new_n948), .ZN(new_n949));
  INV_X1    g0749(.A(new_n941), .ZN(new_n950));
  NOR2_X1   g0750(.A1(new_n668), .A2(new_n950), .ZN(new_n951));
  XNOR2_X1  g0751(.A(new_n949), .B(new_n951), .ZN(new_n952));
  XOR2_X1   g0752(.A(new_n677), .B(KEYINPUT41), .Z(new_n953));
  INV_X1    g0753(.A(new_n660), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n664), .A2(G330), .ZN(new_n955));
  INV_X1    g0755(.A(KEYINPUT95), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n955), .A2(new_n956), .ZN(new_n957));
  AOI21_X1  g0757(.A(new_n954), .B1(new_n957), .B2(new_n665), .ZN(new_n958));
  AOI21_X1  g0758(.A(new_n950), .B1(new_n671), .B2(new_n673), .ZN(new_n959));
  NOR2_X1   g0759(.A1(new_n959), .A2(KEYINPUT45), .ZN(new_n960));
  INV_X1    g0760(.A(KEYINPUT45), .ZN(new_n961));
  AOI211_X1 g0761(.A(new_n961), .B(new_n950), .C1(new_n671), .C2(new_n673), .ZN(new_n962));
  NOR2_X1   g0762(.A1(new_n960), .A2(new_n962), .ZN(new_n963));
  NAND3_X1  g0763(.A1(new_n671), .A2(new_n673), .A3(new_n950), .ZN(new_n964));
  XOR2_X1   g0764(.A(KEYINPUT107), .B(KEYINPUT44), .Z(new_n965));
  INV_X1    g0765(.A(new_n965), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n964), .A2(new_n966), .ZN(new_n967));
  NAND4_X1  g0767(.A1(new_n671), .A2(new_n673), .A3(new_n950), .A4(new_n965), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n967), .A2(new_n968), .ZN(new_n969));
  OAI21_X1  g0769(.A(new_n958), .B1(new_n963), .B2(new_n969), .ZN(new_n970));
  XNOR2_X1  g0770(.A(new_n959), .B(KEYINPUT45), .ZN(new_n971));
  AND2_X1   g0771(.A1(new_n967), .A2(new_n968), .ZN(new_n972));
  NAND3_X1  g0772(.A1(new_n971), .A2(new_n972), .A3(new_n668), .ZN(new_n973));
  AND2_X1   g0773(.A1(new_n970), .A2(new_n973), .ZN(new_n974));
  NOR3_X1   g0774(.A1(new_n666), .A2(new_n667), .A3(new_n660), .ZN(new_n975));
  OAI21_X1  g0775(.A(new_n942), .B1(new_n975), .B2(new_n958), .ZN(new_n976));
  NAND3_X1  g0776(.A1(new_n957), .A2(new_n665), .A3(new_n954), .ZN(new_n977));
  NAND3_X1  g0777(.A1(new_n668), .A2(new_n669), .A3(new_n977), .ZN(new_n978));
  AND2_X1   g0778(.A1(new_n976), .A2(new_n978), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n905), .A2(new_n906), .ZN(new_n980));
  INV_X1    g0780(.A(new_n711), .ZN(new_n981));
  OAI21_X1  g0781(.A(new_n789), .B1(new_n980), .B2(new_n981), .ZN(new_n982));
  OAI21_X1  g0782(.A(KEYINPUT108), .B1(new_n979), .B2(new_n982), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n976), .A2(new_n978), .ZN(new_n984));
  INV_X1    g0784(.A(KEYINPUT108), .ZN(new_n985));
  NAND3_X1  g0785(.A1(new_n712), .A2(new_n984), .A3(new_n985), .ZN(new_n986));
  NAND3_X1  g0786(.A1(new_n974), .A2(new_n983), .A3(new_n986), .ZN(new_n987));
  AOI21_X1  g0787(.A(new_n953), .B1(new_n987), .B2(new_n712), .ZN(new_n988));
  OAI21_X1  g0788(.A(new_n952), .B1(new_n988), .B2(new_n717), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n242), .A2(new_n767), .ZN(new_n990));
  AOI211_X1 g0790(.A(new_n772), .B(new_n721), .C1(new_n676), .C2(new_n601), .ZN(new_n991));
  AOI21_X1  g0791(.A(new_n719), .B1(new_n990), .B2(new_n991), .ZN(new_n992));
  OAI22_X1  g0792(.A1(new_n733), .A2(new_n797), .B1(new_n740), .B2(new_n201), .ZN(new_n993));
  AOI211_X1 g0793(.A(new_n257), .B(new_n993), .C1(G137), .C2(new_n738), .ZN(new_n994));
  INV_X1    g0794(.A(G143), .ZN(new_n995));
  OAI22_X1  g0795(.A1(new_n729), .A2(new_n754), .B1(new_n759), .B2(new_n995), .ZN(new_n996));
  NOR2_X1   g0796(.A1(new_n723), .A2(new_n203), .ZN(new_n997));
  NOR2_X1   g0797(.A1(new_n996), .A2(new_n997), .ZN(new_n998));
  NAND2_X1  g0798(.A1(new_n748), .A2(G77), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n750), .A2(G58), .ZN(new_n1000));
  NAND4_X1  g0800(.A1(new_n994), .A2(new_n998), .A3(new_n999), .A4(new_n1000), .ZN(new_n1001));
  NAND2_X1  g0801(.A1(new_n748), .A2(G97), .ZN(new_n1002));
  AOI21_X1  g0802(.A(new_n456), .B1(G317), .B2(new_n738), .ZN(new_n1003));
  NAND2_X1  g0803(.A1(new_n1002), .A2(new_n1003), .ZN(new_n1004));
  XNOR2_X1  g0804(.A(new_n1004), .B(KEYINPUT109), .ZN(new_n1005));
  NAND3_X1  g0805(.A1(new_n750), .A2(KEYINPUT46), .A3(G116), .ZN(new_n1006));
  INV_X1    g0806(.A(KEYINPUT46), .ZN(new_n1007));
  OAI21_X1  g0807(.A(new_n1007), .B1(new_n745), .B2(new_n472), .ZN(new_n1008));
  OAI22_X1  g0808(.A1(new_n733), .A2(new_n743), .B1(new_n740), .B2(new_n480), .ZN(new_n1009));
  AOI21_X1  g0809(.A(new_n1009), .B1(G107), .B2(new_n724), .ZN(new_n1010));
  AOI22_X1  g0810(.A1(new_n728), .A2(G294), .B1(new_n726), .B2(G311), .ZN(new_n1011));
  NAND4_X1  g0811(.A1(new_n1006), .A2(new_n1008), .A3(new_n1010), .A4(new_n1011), .ZN(new_n1012));
  OAI21_X1  g0812(.A(new_n1001), .B1(new_n1005), .B2(new_n1012), .ZN(new_n1013));
  XOR2_X1   g0813(.A(new_n1013), .B(KEYINPUT110), .Z(new_n1014));
  XNOR2_X1  g0814(.A(new_n1014), .B(KEYINPUT47), .ZN(new_n1015));
  OAI221_X1 g0815(.A(new_n992), .B1(new_n933), .B2(new_n775), .C1(new_n1015), .C2(new_n794), .ZN(new_n1016));
  NAND2_X1  g0816(.A1(new_n989), .A2(new_n1016), .ZN(G387));
  NAND2_X1  g0817(.A1(new_n979), .A2(new_n982), .ZN(new_n1018));
  NAND2_X1  g0818(.A1(new_n712), .A2(new_n984), .ZN(new_n1019));
  NAND3_X1  g0819(.A1(new_n1018), .A2(new_n677), .A3(new_n1019), .ZN(new_n1020));
  NOR2_X1   g0820(.A1(new_n281), .A2(G50), .ZN(new_n1021));
  XOR2_X1   g0821(.A(new_n1021), .B(KEYINPUT50), .Z(new_n1022));
  OAI21_X1  g0822(.A(new_n571), .B1(new_n203), .B2(new_n220), .ZN(new_n1023));
  NOR3_X1   g0823(.A1(new_n1022), .A2(new_n680), .A3(new_n1023), .ZN(new_n1024));
  INV_X1    g0824(.A(new_n237), .ZN(new_n1025));
  OAI21_X1  g0825(.A(new_n767), .B1(new_n1025), .B2(new_n571), .ZN(new_n1026));
  NAND2_X1  g0826(.A1(new_n764), .A2(new_n680), .ZN(new_n1027));
  AOI21_X1  g0827(.A(new_n1024), .B1(new_n1026), .B2(new_n1027), .ZN(new_n1028));
  NOR2_X1   g0828(.A1(new_n211), .A2(G107), .ZN(new_n1029));
  OAI21_X1  g0829(.A(new_n773), .B1(new_n1028), .B2(new_n1029), .ZN(new_n1030));
  NOR2_X1   g0830(.A1(new_n723), .A2(new_n365), .ZN(new_n1031));
  OAI221_X1 g0831(.A(new_n456), .B1(new_n201), .B2(new_n733), .C1(new_n797), .C2(new_n737), .ZN(new_n1032));
  AOI211_X1 g0832(.A(new_n1031), .B(new_n1032), .C1(G159), .C2(new_n726), .ZN(new_n1033));
  OAI22_X1  g0833(.A1(new_n285), .A2(new_n729), .B1(new_n203), .B2(new_n740), .ZN(new_n1034));
  XNOR2_X1  g0834(.A(new_n1034), .B(KEYINPUT111), .ZN(new_n1035));
  NAND2_X1  g0835(.A1(new_n750), .A2(G77), .ZN(new_n1036));
  NAND4_X1  g0836(.A1(new_n1033), .A2(new_n1002), .A3(new_n1035), .A4(new_n1036), .ZN(new_n1037));
  AOI21_X1  g0837(.A(new_n456), .B1(G326), .B2(new_n738), .ZN(new_n1038));
  OAI22_X1  g0838(.A1(new_n745), .A2(new_n808), .B1(new_n480), .B2(new_n723), .ZN(new_n1039));
  AOI22_X1  g0839(.A1(new_n795), .A2(G317), .B1(new_n741), .B2(G303), .ZN(new_n1040));
  NAND2_X1  g0840(.A1(new_n728), .A2(G311), .ZN(new_n1041));
  OAI211_X1 g0841(.A(new_n1040), .B(new_n1041), .C1(new_n734), .C2(new_n759), .ZN(new_n1042));
  INV_X1    g0842(.A(KEYINPUT48), .ZN(new_n1043));
  AOI21_X1  g0843(.A(new_n1039), .B1(new_n1042), .B2(new_n1043), .ZN(new_n1044));
  OAI21_X1  g0844(.A(new_n1044), .B1(new_n1043), .B2(new_n1042), .ZN(new_n1045));
  INV_X1    g0845(.A(KEYINPUT49), .ZN(new_n1046));
  OAI221_X1 g0846(.A(new_n1038), .B1(new_n472), .B2(new_n747), .C1(new_n1045), .C2(new_n1046), .ZN(new_n1047));
  AND2_X1   g0847(.A1(new_n1045), .A2(new_n1046), .ZN(new_n1048));
  OAI21_X1  g0848(.A(new_n1037), .B1(new_n1047), .B2(new_n1048), .ZN(new_n1049));
  AOI21_X1  g0849(.A(new_n719), .B1(new_n1049), .B2(new_n721), .ZN(new_n1050));
  OAI211_X1 g0850(.A(new_n1030), .B(new_n1050), .C1(new_n660), .C2(new_n775), .ZN(new_n1051));
  OAI211_X1 g0851(.A(new_n1020), .B(new_n1051), .C1(new_n716), .C2(new_n979), .ZN(G393));
  NAND2_X1  g0852(.A1(new_n970), .A2(new_n973), .ZN(new_n1053));
  AOI21_X1  g0853(.A(new_n678), .B1(new_n1053), .B2(new_n1019), .ZN(new_n1054));
  NAND2_X1  g0854(.A1(new_n987), .A2(new_n1054), .ZN(new_n1055));
  NAND2_X1  g0855(.A1(new_n974), .A2(new_n717), .ZN(new_n1056));
  INV_X1    g0856(.A(new_n767), .ZN(new_n1057));
  OAI221_X1 g0857(.A(new_n773), .B1(new_n342), .B2(new_n211), .C1(new_n1057), .C2(new_n249), .ZN(new_n1058));
  NAND2_X1  g0858(.A1(new_n1058), .A2(new_n718), .ZN(new_n1059));
  AOI21_X1  g0859(.A(new_n806), .B1(G68), .B2(new_n750), .ZN(new_n1060));
  OAI22_X1  g0860(.A1(new_n759), .A2(new_n797), .B1(new_n733), .B2(new_n754), .ZN(new_n1061));
  XNOR2_X1  g0861(.A(new_n1061), .B(KEYINPUT51), .ZN(new_n1062));
  OAI22_X1  g0862(.A1(new_n740), .A2(new_n281), .B1(new_n737), .B2(new_n995), .ZN(new_n1063));
  NOR2_X1   g0863(.A1(new_n1063), .A2(new_n802), .ZN(new_n1064));
  NOR2_X1   g0864(.A1(new_n723), .A2(new_n220), .ZN(new_n1065));
  AOI21_X1  g0865(.A(new_n1065), .B1(new_n728), .B2(G50), .ZN(new_n1066));
  NAND4_X1  g0866(.A1(new_n1060), .A2(new_n1062), .A3(new_n1064), .A4(new_n1066), .ZN(new_n1067));
  AOI22_X1  g0867(.A1(new_n795), .A2(G311), .B1(G317), .B2(new_n726), .ZN(new_n1068));
  XNOR2_X1  g0868(.A(new_n1068), .B(KEYINPUT112), .ZN(new_n1069));
  XOR2_X1   g0869(.A(new_n1069), .B(KEYINPUT52), .Z(new_n1070));
  NAND2_X1  g0870(.A1(new_n750), .A2(G283), .ZN(new_n1071));
  OAI21_X1  g0871(.A(new_n257), .B1(new_n737), .B2(new_n734), .ZN(new_n1072));
  AOI21_X1  g0872(.A(new_n1072), .B1(G294), .B2(new_n741), .ZN(new_n1073));
  AOI22_X1  g0873(.A1(new_n724), .A2(G116), .B1(G303), .B2(new_n728), .ZN(new_n1074));
  NAND4_X1  g0874(.A1(new_n752), .A2(new_n1071), .A3(new_n1073), .A4(new_n1074), .ZN(new_n1075));
  OAI21_X1  g0875(.A(new_n1067), .B1(new_n1070), .B2(new_n1075), .ZN(new_n1076));
  AOI21_X1  g0876(.A(new_n1059), .B1(new_n1076), .B2(new_n721), .ZN(new_n1077));
  OAI21_X1  g0877(.A(new_n1077), .B1(new_n941), .B2(new_n775), .ZN(new_n1078));
  NAND3_X1  g0878(.A1(new_n1055), .A2(new_n1056), .A3(new_n1078), .ZN(G390));
  INV_X1    g0879(.A(new_n792), .ZN(new_n1080));
  OAI21_X1  g0880(.A(new_n718), .B1(new_n286), .B2(new_n1080), .ZN(new_n1081));
  AND2_X1   g0881(.A1(new_n795), .A2(G132), .ZN(new_n1082));
  AOI211_X1 g0882(.A(new_n257), .B(new_n1082), .C1(G125), .C2(new_n738), .ZN(new_n1083));
  INV_X1    g0883(.A(G128), .ZN(new_n1084));
  OAI22_X1  g0884(.A1(new_n729), .A2(new_n798), .B1(new_n759), .B2(new_n1084), .ZN(new_n1085));
  AOI21_X1  g0885(.A(new_n1085), .B1(G159), .B2(new_n724), .ZN(new_n1086));
  XNOR2_X1  g0886(.A(KEYINPUT54), .B(G143), .ZN(new_n1087));
  XNOR2_X1  g0887(.A(new_n1087), .B(KEYINPUT116), .ZN(new_n1088));
  NAND2_X1  g0888(.A1(new_n1088), .A2(new_n741), .ZN(new_n1089));
  NAND2_X1  g0889(.A1(new_n748), .A2(G50), .ZN(new_n1090));
  NAND4_X1  g0890(.A1(new_n1083), .A2(new_n1086), .A3(new_n1089), .A4(new_n1090), .ZN(new_n1091));
  NAND2_X1  g0891(.A1(new_n750), .A2(G150), .ZN(new_n1092));
  XNOR2_X1  g0892(.A(new_n1092), .B(KEYINPUT53), .ZN(new_n1093));
  OAI22_X1  g0893(.A1(new_n740), .A2(new_n342), .B1(new_n737), .B2(new_n808), .ZN(new_n1094));
  AOI211_X1 g0894(.A(new_n258), .B(new_n1094), .C1(G116), .C2(new_n795), .ZN(new_n1095));
  OAI211_X1 g0895(.A(new_n1095), .B(new_n751), .C1(new_n203), .C2(new_n747), .ZN(new_n1096));
  AOI21_X1  g0896(.A(new_n1065), .B1(new_n728), .B2(G107), .ZN(new_n1097));
  OAI21_X1  g0897(.A(new_n1097), .B1(new_n480), .B2(new_n759), .ZN(new_n1098));
  OAI22_X1  g0898(.A1(new_n1091), .A2(new_n1093), .B1(new_n1096), .B2(new_n1098), .ZN(new_n1099));
  AOI21_X1  g0899(.A(new_n1081), .B1(new_n1099), .B2(new_n721), .ZN(new_n1100));
  OAI21_X1  g0900(.A(new_n1100), .B1(new_n879), .B2(new_n771), .ZN(new_n1101));
  NAND2_X1  g0901(.A1(new_n638), .A2(new_n654), .ZN(new_n1102));
  OAI21_X1  g0902(.A(new_n1102), .B1(new_n890), .B2(new_n899), .ZN(new_n1103));
  OAI211_X1 g0903(.A(new_n1103), .B(new_n870), .C1(new_n855), .C2(new_n878), .ZN(new_n1104));
  XOR2_X1   g0904(.A(new_n898), .B(KEYINPUT113), .Z(new_n1105));
  NAND2_X1  g0905(.A1(new_n781), .A2(new_n386), .ZN(new_n1106));
  AOI21_X1  g0906(.A(new_n779), .B1(new_n709), .B2(new_n1106), .ZN(new_n1107));
  OAI211_X1 g0907(.A(new_n914), .B(new_n1102), .C1(new_n1105), .C2(new_n1107), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n1104), .A2(new_n1108), .ZN(new_n1109));
  NAND3_X1  g0909(.A1(new_n699), .A2(new_n782), .A3(new_n898), .ZN(new_n1110));
  INV_X1    g0910(.A(new_n1110), .ZN(new_n1111));
  NAND2_X1  g0911(.A1(new_n1109), .A2(new_n1111), .ZN(new_n1112));
  NAND3_X1  g0912(.A1(new_n1104), .A2(new_n1110), .A3(new_n1108), .ZN(new_n1113));
  NAND2_X1  g0913(.A1(new_n1112), .A2(new_n1113), .ZN(new_n1114));
  OAI21_X1  g0914(.A(new_n1101), .B1(new_n1114), .B2(new_n716), .ZN(new_n1115));
  INV_X1    g0915(.A(KEYINPUT114), .ZN(new_n1116));
  AND3_X1   g0916(.A1(new_n699), .A2(new_n1116), .A3(new_n455), .ZN(new_n1117));
  AOI21_X1  g0917(.A(new_n1116), .B1(new_n699), .B2(new_n455), .ZN(new_n1118));
  OAI211_X1 g0918(.A(new_n907), .B(new_n643), .C1(new_n1117), .C2(new_n1118), .ZN(new_n1119));
  AOI21_X1  g0919(.A(new_n898), .B1(new_n699), .B2(new_n782), .ZN(new_n1120));
  OAI22_X1  g0920(.A1(new_n1111), .A2(new_n1120), .B1(new_n784), .B2(new_n886), .ZN(new_n1121));
  OAI21_X1  g0921(.A(new_n1105), .B1(new_n789), .B2(new_n783), .ZN(new_n1122));
  NAND3_X1  g0922(.A1(new_n1122), .A2(new_n1110), .A3(new_n1107), .ZN(new_n1123));
  AOI21_X1  g0923(.A(new_n1119), .B1(new_n1121), .B2(new_n1123), .ZN(new_n1124));
  NAND3_X1  g0924(.A1(new_n1124), .A2(new_n1112), .A3(new_n1113), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n1125), .A2(new_n677), .ZN(new_n1126));
  INV_X1    g0926(.A(KEYINPUT115), .ZN(new_n1127));
  INV_X1    g0927(.A(new_n1124), .ZN(new_n1128));
  AOI22_X1  g0928(.A1(new_n1126), .A2(new_n1127), .B1(new_n1114), .B2(new_n1128), .ZN(new_n1129));
  NAND3_X1  g0929(.A1(new_n1125), .A2(KEYINPUT115), .A3(new_n677), .ZN(new_n1130));
  AOI21_X1  g0930(.A(new_n1115), .B1(new_n1129), .B2(new_n1130), .ZN(new_n1131));
  INV_X1    g0931(.A(new_n1131), .ZN(G378));
  NAND2_X1  g0932(.A1(new_n299), .A2(new_n823), .ZN(new_n1133));
  XOR2_X1   g0933(.A(new_n1133), .B(KEYINPUT55), .Z(new_n1134));
  XNOR2_X1  g0934(.A(new_n317), .B(new_n1134), .ZN(new_n1135));
  XNOR2_X1  g0935(.A(KEYINPUT119), .B(KEYINPUT56), .ZN(new_n1136));
  XNOR2_X1  g0936(.A(new_n1135), .B(new_n1136), .ZN(new_n1137));
  AOI21_X1  g0937(.A(new_n698), .B1(new_n915), .B2(new_n914), .ZN(new_n1138));
  INV_X1    g0938(.A(new_n1138), .ZN(new_n1139));
  AOI21_X1  g0939(.A(new_n1139), .B1(new_n912), .B2(new_n913), .ZN(new_n1140));
  OAI21_X1  g0940(.A(new_n1137), .B1(new_n1140), .B2(KEYINPUT120), .ZN(new_n1141));
  INV_X1    g0941(.A(KEYINPUT120), .ZN(new_n1142));
  AOI211_X1 g0942(.A(new_n1142), .B(new_n1139), .C1(new_n913), .C2(new_n912), .ZN(new_n1143));
  NOR2_X1   g0943(.A1(new_n1141), .A2(new_n1143), .ZN(new_n1144));
  AND3_X1   g0944(.A1(new_n875), .A2(new_n877), .A3(KEYINPUT104), .ZN(new_n1145));
  AOI21_X1  g0945(.A(KEYINPUT104), .B1(new_n875), .B2(new_n877), .ZN(new_n1146));
  INV_X1    g0946(.A(new_n911), .ZN(new_n1147));
  NOR3_X1   g0947(.A1(new_n1145), .A2(new_n1146), .A3(new_n1147), .ZN(new_n1148));
  OAI21_X1  g0948(.A(new_n1138), .B1(new_n1148), .B2(KEYINPUT40), .ZN(new_n1149));
  NOR3_X1   g0949(.A1(new_n1149), .A2(new_n1142), .A3(new_n1137), .ZN(new_n1150));
  OAI21_X1  g0950(.A(new_n904), .B1(new_n1144), .B2(new_n1150), .ZN(new_n1151));
  NAND2_X1  g0951(.A1(new_n1149), .A2(new_n1142), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n1140), .A2(KEYINPUT120), .ZN(new_n1153));
  NAND3_X1  g0953(.A1(new_n1152), .A2(new_n1153), .A3(new_n1137), .ZN(new_n1154));
  NAND2_X1  g0954(.A1(new_n1141), .A2(new_n1143), .ZN(new_n1155));
  INV_X1    g0955(.A(new_n904), .ZN(new_n1156));
  NAND3_X1  g0956(.A1(new_n1154), .A2(new_n1155), .A3(new_n1156), .ZN(new_n1157));
  INV_X1    g0957(.A(new_n1119), .ZN(new_n1158));
  NAND2_X1  g0958(.A1(new_n1125), .A2(new_n1158), .ZN(new_n1159));
  NAND3_X1  g0959(.A1(new_n1151), .A2(new_n1157), .A3(new_n1159), .ZN(new_n1160));
  INV_X1    g0960(.A(KEYINPUT57), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n1160), .A2(new_n1161), .ZN(new_n1162));
  NAND4_X1  g0962(.A1(new_n1151), .A2(new_n1157), .A3(KEYINPUT57), .A4(new_n1159), .ZN(new_n1163));
  NAND3_X1  g0963(.A1(new_n1162), .A2(new_n677), .A3(new_n1163), .ZN(new_n1164));
  NAND3_X1  g0964(.A1(new_n1151), .A2(new_n717), .A3(new_n1157), .ZN(new_n1165));
  OAI21_X1  g0965(.A(new_n718), .B1(G50), .B2(new_n1080), .ZN(new_n1166));
  NOR2_X1   g0966(.A1(new_n456), .A2(new_n268), .ZN(new_n1167));
  AOI211_X1 g0967(.A(G50), .B(new_n1167), .C1(new_n251), .C2(new_n252), .ZN(new_n1168));
  NAND2_X1  g0968(.A1(new_n748), .A2(G58), .ZN(new_n1169));
  AND2_X1   g0969(.A1(new_n1169), .A2(new_n1167), .ZN(new_n1170));
  NOR2_X1   g0970(.A1(new_n759), .A2(new_n472), .ZN(new_n1171));
  AOI211_X1 g0971(.A(new_n997), .B(new_n1171), .C1(G97), .C2(new_n728), .ZN(new_n1172));
  OAI22_X1  g0972(.A1(new_n740), .A2(new_n365), .B1(new_n737), .B2(new_n480), .ZN(new_n1173));
  AOI21_X1  g0973(.A(new_n1173), .B1(G107), .B2(new_n795), .ZN(new_n1174));
  NAND4_X1  g0974(.A1(new_n1170), .A2(new_n1036), .A3(new_n1172), .A4(new_n1174), .ZN(new_n1175));
  INV_X1    g0975(.A(KEYINPUT58), .ZN(new_n1176));
  AOI21_X1  g0976(.A(new_n1168), .B1(new_n1175), .B2(new_n1176), .ZN(new_n1177));
  AOI22_X1  g0977(.A1(new_n724), .A2(G150), .B1(G125), .B2(new_n726), .ZN(new_n1178));
  XNOR2_X1  g0978(.A(new_n1178), .B(KEYINPUT117), .ZN(new_n1179));
  NAND2_X1  g0979(.A1(new_n750), .A2(new_n1088), .ZN(new_n1180));
  OAI22_X1  g0980(.A1(new_n733), .A2(new_n1084), .B1(new_n740), .B2(new_n798), .ZN(new_n1181));
  AOI21_X1  g0981(.A(new_n1181), .B1(G132), .B2(new_n728), .ZN(new_n1182));
  NAND3_X1  g0982(.A1(new_n1179), .A2(new_n1180), .A3(new_n1182), .ZN(new_n1183));
  NOR2_X1   g0983(.A1(new_n1183), .A2(KEYINPUT59), .ZN(new_n1184));
  NAND2_X1  g0984(.A1(new_n1183), .A2(KEYINPUT59), .ZN(new_n1185));
  AOI211_X1 g0985(.A(G33), .B(G41), .C1(new_n738), .C2(G124), .ZN(new_n1186));
  OAI21_X1  g0986(.A(new_n1186), .B1(new_n754), .B2(new_n747), .ZN(new_n1187));
  XNOR2_X1  g0987(.A(new_n1187), .B(KEYINPUT118), .ZN(new_n1188));
  NAND2_X1  g0988(.A1(new_n1185), .A2(new_n1188), .ZN(new_n1189));
  OAI221_X1 g0989(.A(new_n1177), .B1(new_n1176), .B2(new_n1175), .C1(new_n1184), .C2(new_n1189), .ZN(new_n1190));
  AOI21_X1  g0990(.A(new_n1166), .B1(new_n1190), .B2(new_n721), .ZN(new_n1191));
  OAI21_X1  g0991(.A(new_n1191), .B1(new_n1137), .B2(new_n771), .ZN(new_n1192));
  NAND2_X1  g0992(.A1(new_n1165), .A2(new_n1192), .ZN(new_n1193));
  INV_X1    g0993(.A(new_n1193), .ZN(new_n1194));
  NAND2_X1  g0994(.A1(new_n1164), .A2(new_n1194), .ZN(G375));
  NAND2_X1  g0995(.A1(new_n1121), .A2(new_n1123), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(new_n1105), .A2(new_n770), .ZN(new_n1197));
  OAI21_X1  g0997(.A(new_n718), .B1(G68), .B2(new_n1080), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(new_n1169), .A2(new_n456), .ZN(new_n1199));
  XOR2_X1   g0999(.A(new_n1199), .B(KEYINPUT121), .Z(new_n1200));
  NAND2_X1  g1000(.A1(new_n750), .A2(G159), .ZN(new_n1201));
  OAI22_X1  g1001(.A1(new_n733), .A2(new_n798), .B1(new_n737), .B2(new_n1084), .ZN(new_n1202));
  AOI21_X1  g1002(.A(new_n1202), .B1(G150), .B2(new_n741), .ZN(new_n1203));
  AOI22_X1  g1003(.A1(new_n724), .A2(G50), .B1(G132), .B2(new_n726), .ZN(new_n1204));
  NAND2_X1  g1004(.A1(new_n1088), .A2(new_n728), .ZN(new_n1205));
  NAND4_X1  g1005(.A1(new_n1201), .A2(new_n1203), .A3(new_n1204), .A4(new_n1205), .ZN(new_n1206));
  AOI21_X1  g1006(.A(new_n1031), .B1(new_n728), .B2(G116), .ZN(new_n1207));
  OAI21_X1  g1007(.A(new_n1207), .B1(new_n808), .B2(new_n759), .ZN(new_n1208));
  OAI22_X1  g1008(.A1(new_n740), .A2(new_n375), .B1(new_n737), .B2(new_n743), .ZN(new_n1209));
  AOI211_X1 g1009(.A(new_n258), .B(new_n1209), .C1(G283), .C2(new_n795), .ZN(new_n1210));
  OAI211_X1 g1010(.A(new_n1210), .B(new_n999), .C1(new_n342), .C2(new_n745), .ZN(new_n1211));
  OAI22_X1  g1011(.A1(new_n1200), .A2(new_n1206), .B1(new_n1208), .B2(new_n1211), .ZN(new_n1212));
  AOI21_X1  g1012(.A(new_n1198), .B1(new_n1212), .B2(new_n721), .ZN(new_n1213));
  AOI22_X1  g1013(.A1(new_n1196), .A2(new_n717), .B1(new_n1197), .B2(new_n1213), .ZN(new_n1214));
  INV_X1    g1014(.A(new_n953), .ZN(new_n1215));
  NAND2_X1  g1015(.A1(new_n1128), .A2(new_n1215), .ZN(new_n1216));
  NOR2_X1   g1016(.A1(new_n1196), .A2(new_n1158), .ZN(new_n1217));
  OAI21_X1  g1017(.A(new_n1214), .B1(new_n1216), .B2(new_n1217), .ZN(G381));
  NOR2_X1   g1018(.A1(G375), .A2(G378), .ZN(new_n1219));
  AND3_X1   g1019(.A1(new_n1055), .A2(new_n1056), .A3(new_n1078), .ZN(new_n1220));
  NAND3_X1  g1020(.A1(new_n989), .A2(new_n1220), .A3(new_n1016), .ZN(new_n1221));
  OR3_X1    g1021(.A1(G393), .A2(G396), .A3(G384), .ZN(new_n1222));
  NOR3_X1   g1022(.A1(new_n1221), .A2(G381), .A3(new_n1222), .ZN(new_n1223));
  NAND2_X1  g1023(.A1(new_n1219), .A2(new_n1223), .ZN(G407));
  OAI21_X1  g1024(.A(new_n1219), .B1(new_n652), .B2(new_n1223), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(new_n1225), .A2(G213), .ZN(G409));
  XNOR2_X1  g1026(.A(G393), .B(new_n777), .ZN(new_n1227));
  INV_X1    g1027(.A(new_n1227), .ZN(new_n1228));
  AND3_X1   g1028(.A1(new_n989), .A2(new_n1016), .A3(new_n1220), .ZN(new_n1229));
  AOI21_X1  g1029(.A(new_n1220), .B1(new_n989), .B2(new_n1016), .ZN(new_n1230));
  NOR3_X1   g1030(.A1(new_n1229), .A2(new_n1230), .A3(KEYINPUT123), .ZN(new_n1231));
  INV_X1    g1031(.A(KEYINPUT123), .ZN(new_n1232));
  INV_X1    g1032(.A(new_n951), .ZN(new_n1233));
  XNOR2_X1  g1033(.A(new_n949), .B(new_n1233), .ZN(new_n1234));
  AND3_X1   g1034(.A1(new_n712), .A2(new_n984), .A3(new_n985), .ZN(new_n1235));
  AOI21_X1  g1035(.A(new_n985), .B1(new_n712), .B2(new_n984), .ZN(new_n1236));
  NOR3_X1   g1036(.A1(new_n1235), .A2(new_n1236), .A3(new_n1053), .ZN(new_n1237));
  OAI21_X1  g1037(.A(new_n1215), .B1(new_n1237), .B2(new_n982), .ZN(new_n1238));
  AOI21_X1  g1038(.A(new_n1234), .B1(new_n1238), .B2(new_n716), .ZN(new_n1239));
  INV_X1    g1039(.A(new_n1016), .ZN(new_n1240));
  OAI21_X1  g1040(.A(G390), .B1(new_n1239), .B2(new_n1240), .ZN(new_n1241));
  AOI21_X1  g1041(.A(new_n1232), .B1(new_n1241), .B2(new_n1221), .ZN(new_n1242));
  OAI21_X1  g1042(.A(new_n1228), .B1(new_n1231), .B2(new_n1242), .ZN(new_n1243));
  OAI21_X1  g1043(.A(KEYINPUT123), .B1(new_n1229), .B2(new_n1230), .ZN(new_n1244));
  NAND3_X1  g1044(.A1(new_n1241), .A2(new_n1232), .A3(new_n1221), .ZN(new_n1245));
  NAND3_X1  g1045(.A1(new_n1244), .A2(new_n1227), .A3(new_n1245), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(new_n1243), .A2(new_n1246), .ZN(new_n1247));
  XNOR2_X1  g1047(.A(new_n1247), .B(KEYINPUT125), .ZN(new_n1248));
  INV_X1    g1048(.A(G213), .ZN(new_n1249));
  NOR2_X1   g1049(.A1(new_n1249), .A2(G343), .ZN(new_n1250));
  INV_X1    g1050(.A(new_n1250), .ZN(new_n1251));
  AOI21_X1  g1051(.A(new_n678), .B1(new_n1160), .B2(new_n1161), .ZN(new_n1252));
  AOI211_X1 g1052(.A(new_n1131), .B(new_n1193), .C1(new_n1252), .C2(new_n1163), .ZN(new_n1253));
  OAI211_X1 g1053(.A(new_n1165), .B(new_n1192), .C1(new_n1160), .C2(new_n953), .ZN(new_n1254));
  NAND2_X1  g1054(.A1(new_n1254), .A2(new_n1131), .ZN(new_n1255));
  INV_X1    g1055(.A(new_n1255), .ZN(new_n1256));
  OAI21_X1  g1056(.A(new_n1251), .B1(new_n1253), .B2(new_n1256), .ZN(new_n1257));
  OAI21_X1  g1057(.A(new_n1128), .B1(new_n1217), .B2(KEYINPUT60), .ZN(new_n1258));
  INV_X1    g1058(.A(KEYINPUT122), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(new_n1258), .A2(new_n1259), .ZN(new_n1260));
  OAI211_X1 g1060(.A(new_n1128), .B(KEYINPUT122), .C1(new_n1217), .C2(KEYINPUT60), .ZN(new_n1261));
  AOI21_X1  g1061(.A(new_n678), .B1(new_n1217), .B2(KEYINPUT60), .ZN(new_n1262));
  NAND3_X1  g1062(.A1(new_n1260), .A2(new_n1261), .A3(new_n1262), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n1263), .A2(new_n1214), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(new_n1264), .A2(new_n815), .ZN(new_n1265));
  NAND3_X1  g1065(.A1(new_n1263), .A2(G384), .A3(new_n1214), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(new_n1265), .A2(new_n1266), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(new_n1250), .A2(G2897), .ZN(new_n1268));
  XNOR2_X1  g1068(.A(new_n1267), .B(new_n1268), .ZN(new_n1269));
  AOI21_X1  g1069(.A(KEYINPUT61), .B1(new_n1257), .B2(new_n1269), .ZN(new_n1270));
  INV_X1    g1070(.A(new_n1267), .ZN(new_n1271));
  OAI211_X1 g1071(.A(new_n1251), .B(new_n1271), .C1(new_n1253), .C2(new_n1256), .ZN(new_n1272));
  NAND2_X1  g1072(.A1(new_n1272), .A2(KEYINPUT62), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(new_n1270), .A2(new_n1273), .ZN(new_n1274));
  NOR2_X1   g1074(.A1(new_n1272), .A2(KEYINPUT62), .ZN(new_n1275));
  OAI21_X1  g1075(.A(new_n1248), .B1(new_n1274), .B2(new_n1275), .ZN(new_n1276));
  INV_X1    g1076(.A(KEYINPUT124), .ZN(new_n1277));
  INV_X1    g1077(.A(KEYINPUT63), .ZN(new_n1278));
  NOR2_X1   g1078(.A1(new_n1267), .A2(new_n1278), .ZN(new_n1279));
  OAI211_X1 g1079(.A(new_n1251), .B(new_n1279), .C1(new_n1253), .C2(new_n1256), .ZN(new_n1280));
  INV_X1    g1080(.A(new_n1246), .ZN(new_n1281));
  AOI21_X1  g1081(.A(new_n1227), .B1(new_n1244), .B2(new_n1245), .ZN(new_n1282));
  NOR2_X1   g1082(.A1(new_n1281), .A2(new_n1282), .ZN(new_n1283));
  NAND2_X1  g1083(.A1(new_n1280), .A2(new_n1283), .ZN(new_n1284));
  NAND3_X1  g1084(.A1(new_n1164), .A2(G378), .A3(new_n1194), .ZN(new_n1285));
  AOI21_X1  g1085(.A(new_n1250), .B1(new_n1285), .B2(new_n1255), .ZN(new_n1286));
  AOI21_X1  g1086(.A(KEYINPUT63), .B1(new_n1286), .B2(new_n1271), .ZN(new_n1287));
  NOR2_X1   g1087(.A1(new_n1284), .A2(new_n1287), .ZN(new_n1288));
  AOI21_X1  g1088(.A(new_n1277), .B1(new_n1288), .B2(new_n1270), .ZN(new_n1289));
  AOI21_X1  g1089(.A(new_n1247), .B1(new_n1286), .B2(new_n1279), .ZN(new_n1290));
  NAND2_X1  g1090(.A1(new_n1272), .A2(new_n1278), .ZN(new_n1291));
  AND4_X1   g1091(.A1(new_n1277), .A2(new_n1270), .A3(new_n1290), .A4(new_n1291), .ZN(new_n1292));
  OAI21_X1  g1092(.A(new_n1276), .B1(new_n1289), .B2(new_n1292), .ZN(G405));
  NAND2_X1  g1093(.A1(G375), .A2(new_n1131), .ZN(new_n1294));
  XNOR2_X1  g1094(.A(new_n1294), .B(new_n1271), .ZN(new_n1295));
  INV_X1    g1095(.A(KEYINPUT126), .ZN(new_n1296));
  NAND2_X1  g1096(.A1(new_n1285), .A2(new_n1296), .ZN(new_n1297));
  AND2_X1   g1097(.A1(new_n1295), .A2(new_n1297), .ZN(new_n1298));
  NOR2_X1   g1098(.A1(new_n1295), .A2(new_n1297), .ZN(new_n1299));
  OAI21_X1  g1099(.A(new_n1247), .B1(new_n1298), .B2(new_n1299), .ZN(new_n1300));
  XNOR2_X1  g1100(.A(new_n1294), .B(new_n1267), .ZN(new_n1301));
  NAND3_X1  g1101(.A1(new_n1301), .A2(new_n1296), .A3(new_n1285), .ZN(new_n1302));
  NAND2_X1  g1102(.A1(new_n1295), .A2(new_n1297), .ZN(new_n1303));
  NAND3_X1  g1103(.A1(new_n1302), .A2(new_n1283), .A3(new_n1303), .ZN(new_n1304));
  NAND2_X1  g1104(.A1(new_n1300), .A2(new_n1304), .ZN(G402));
endmodule


