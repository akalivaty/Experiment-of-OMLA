

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
         n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
         n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
         n1043, n1044;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NOR2_X1 U560 ( .A1(n666), .A2(n555), .ZN(n653) );
  XOR2_X1 U561 ( .A(n725), .B(KEYINPUT28), .Z(n526) );
  NOR2_X2 U562 ( .A1(G651), .A2(n666), .ZN(n550) );
  XOR2_X2 U563 ( .A(G543), .B(KEYINPUT0), .Z(n666) );
  XNOR2_X2 U564 ( .A(n704), .B(n796), .ZN(n705) );
  OR2_X2 U565 ( .A1(n703), .A2(n702), .ZN(n796) );
  OR2_X1 U566 ( .A1(n597), .A2(n596), .ZN(n599) );
  INV_X1 U567 ( .A(KEYINPUT17), .ZN(n531) );
  NOR2_X1 U568 ( .A1(G2105), .A2(G2104), .ZN(n532) );
  INV_X1 U569 ( .A(n1002), .ZN(n781) );
  NAND2_X1 U570 ( .A1(n879), .A2(G137), .ZN(n573) );
  INV_X1 U571 ( .A(KEYINPUT23), .ZN(n570) );
  NOR2_X1 U572 ( .A1(n781), .A2(n780), .ZN(n527) );
  XNOR2_X1 U573 ( .A(n610), .B(KEYINPUT5), .ZN(n528) );
  AND2_X1 U574 ( .A1(n992), .A2(n840), .ZN(n529) );
  XOR2_X1 U575 ( .A(KEYINPUT6), .B(n606), .Z(n530) );
  INV_X1 U576 ( .A(KEYINPUT26), .ZN(n709) );
  OR2_X1 U577 ( .A1(n995), .A2(n716), .ZN(n715) );
  INV_X1 U578 ( .A(KEYINPUT96), .ZN(n748) );
  NAND2_X1 U579 ( .A1(G8), .A2(n755), .ZN(n753) );
  BUF_X1 U580 ( .A(n753), .Z(n791) );
  XNOR2_X1 U581 ( .A(KEYINPUT15), .B(KEYINPUT73), .ZN(n598) );
  INV_X1 U582 ( .A(G2105), .ZN(n535) );
  NOR2_X1 U583 ( .A1(n827), .A2(n529), .ZN(n828) );
  XNOR2_X1 U584 ( .A(n599), .B(n598), .ZN(n995) );
  XOR2_X1 U585 ( .A(KEYINPUT1), .B(n549), .Z(n670) );
  NAND2_X1 U586 ( .A1(n530), .A2(n528), .ZN(n611) );
  XNOR2_X1 U587 ( .A(n571), .B(n570), .ZN(n572) );
  XNOR2_X1 U588 ( .A(n611), .B(KEYINPUT7), .ZN(n612) );
  XNOR2_X2 U589 ( .A(n532), .B(n531), .ZN(n879) );
  NAND2_X1 U590 ( .A1(G138), .A2(n879), .ZN(n534) );
  AND2_X4 U591 ( .A1(n535), .A2(G2104), .ZN(n881) );
  NAND2_X1 U592 ( .A1(G102), .A2(n881), .ZN(n533) );
  NAND2_X1 U593 ( .A1(n534), .A2(n533), .ZN(n539) );
  NOR2_X2 U594 ( .A1(G2104), .A2(n535), .ZN(n885) );
  NAND2_X1 U595 ( .A1(G126), .A2(n885), .ZN(n537) );
  AND2_X1 U596 ( .A1(G2105), .A2(G2104), .ZN(n888) );
  NAND2_X1 U597 ( .A1(G114), .A2(n888), .ZN(n536) );
  NAND2_X1 U598 ( .A1(n537), .A2(n536), .ZN(n538) );
  NOR2_X1 U599 ( .A1(n539), .A2(n538), .ZN(G164) );
  XOR2_X1 U600 ( .A(G2443), .B(G2446), .Z(n541) );
  XNOR2_X1 U601 ( .A(G2427), .B(G2451), .ZN(n540) );
  XNOR2_X1 U602 ( .A(n541), .B(n540), .ZN(n547) );
  XOR2_X1 U603 ( .A(G2430), .B(G2454), .Z(n543) );
  XNOR2_X1 U604 ( .A(G1341), .B(G1348), .ZN(n542) );
  XNOR2_X1 U605 ( .A(n543), .B(n542), .ZN(n545) );
  XOR2_X1 U606 ( .A(G2435), .B(G2438), .Z(n544) );
  XNOR2_X1 U607 ( .A(n545), .B(n544), .ZN(n546) );
  XOR2_X1 U608 ( .A(n547), .B(n546), .Z(n548) );
  AND2_X1 U609 ( .A1(G14), .A2(n548), .ZN(G401) );
  INV_X1 U610 ( .A(G651), .ZN(n555) );
  NOR2_X1 U611 ( .A1(G543), .A2(n555), .ZN(n549) );
  NAND2_X1 U612 ( .A1(G64), .A2(n670), .ZN(n553) );
  XNOR2_X1 U613 ( .A(n550), .B(KEYINPUT64), .ZN(n588) );
  INV_X1 U614 ( .A(n588), .ZN(n551) );
  INV_X1 U615 ( .A(n551), .ZN(n664) );
  NAND2_X1 U616 ( .A1(G52), .A2(n664), .ZN(n552) );
  NAND2_X1 U617 ( .A1(n553), .A2(n552), .ZN(n554) );
  XNOR2_X1 U618 ( .A(KEYINPUT66), .B(n554), .ZN(n562) );
  XNOR2_X1 U619 ( .A(KEYINPUT68), .B(KEYINPUT9), .ZN(n560) );
  NAND2_X1 U620 ( .A1(n653), .A2(G77), .ZN(n558) );
  NOR2_X1 U621 ( .A1(G651), .A2(G543), .ZN(n656) );
  NAND2_X1 U622 ( .A1(n656), .A2(G90), .ZN(n556) );
  XOR2_X1 U623 ( .A(KEYINPUT67), .B(n556), .Z(n557) );
  NAND2_X1 U624 ( .A1(n558), .A2(n557), .ZN(n559) );
  XOR2_X1 U625 ( .A(n560), .B(n559), .Z(n561) );
  NOR2_X1 U626 ( .A1(n562), .A2(n561), .ZN(G171) );
  AND2_X1 U627 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U628 ( .A(G57), .ZN(G237) );
  INV_X1 U629 ( .A(G108), .ZN(G238) );
  INV_X1 U630 ( .A(G120), .ZN(G236) );
  NAND2_X1 U631 ( .A1(G62), .A2(n670), .ZN(n564) );
  NAND2_X1 U632 ( .A1(G50), .A2(n664), .ZN(n563) );
  NAND2_X1 U633 ( .A1(n564), .A2(n563), .ZN(n569) );
  NAND2_X1 U634 ( .A1(G88), .A2(n656), .ZN(n566) );
  NAND2_X1 U635 ( .A1(G75), .A2(n653), .ZN(n565) );
  NAND2_X1 U636 ( .A1(n566), .A2(n565), .ZN(n567) );
  XOR2_X1 U637 ( .A(KEYINPUT81), .B(n567), .Z(n568) );
  NOR2_X1 U638 ( .A1(n569), .A2(n568), .ZN(G166) );
  NAND2_X1 U639 ( .A1(G101), .A2(n881), .ZN(n571) );
  NAND2_X1 U640 ( .A1(n573), .A2(n572), .ZN(n703) );
  NAND2_X1 U641 ( .A1(G125), .A2(n885), .ZN(n575) );
  NAND2_X1 U642 ( .A1(G113), .A2(n888), .ZN(n574) );
  NAND2_X1 U643 ( .A1(n575), .A2(n574), .ZN(n701) );
  NOR2_X1 U644 ( .A1(n703), .A2(n701), .ZN(G160) );
  NAND2_X1 U645 ( .A1(G7), .A2(G661), .ZN(n576) );
  XNOR2_X1 U646 ( .A(n576), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U647 ( .A(G223), .ZN(n846) );
  NAND2_X1 U648 ( .A1(n846), .A2(G567), .ZN(n577) );
  XOR2_X1 U649 ( .A(KEYINPUT11), .B(n577), .Z(G234) );
  NAND2_X1 U650 ( .A1(n656), .A2(G81), .ZN(n578) );
  XNOR2_X1 U651 ( .A(n578), .B(KEYINPUT12), .ZN(n580) );
  NAND2_X1 U652 ( .A1(G68), .A2(n653), .ZN(n579) );
  NAND2_X1 U653 ( .A1(n580), .A2(n579), .ZN(n581) );
  XNOR2_X1 U654 ( .A(KEYINPUT13), .B(n581), .ZN(n587) );
  NAND2_X1 U655 ( .A1(G56), .A2(n670), .ZN(n582) );
  XOR2_X1 U656 ( .A(KEYINPUT14), .B(n582), .Z(n585) );
  NAND2_X1 U657 ( .A1(G43), .A2(n664), .ZN(n583) );
  XNOR2_X1 U658 ( .A(KEYINPUT69), .B(n583), .ZN(n584) );
  NOR2_X1 U659 ( .A1(n585), .A2(n584), .ZN(n586) );
  NAND2_X1 U660 ( .A1(n587), .A2(n586), .ZN(n1001) );
  INV_X1 U661 ( .A(G860), .ZN(n637) );
  OR2_X1 U662 ( .A1(n1001), .A2(n637), .ZN(G153) );
  NAND2_X1 U663 ( .A1(n588), .A2(G54), .ZN(n589) );
  XOR2_X1 U664 ( .A(n589), .B(KEYINPUT71), .Z(n591) );
  NAND2_X1 U665 ( .A1(n653), .A2(G79), .ZN(n590) );
  NAND2_X1 U666 ( .A1(n591), .A2(n590), .ZN(n592) );
  XNOR2_X1 U667 ( .A(n592), .B(KEYINPUT72), .ZN(n597) );
  NAND2_X1 U668 ( .A1(G66), .A2(n670), .ZN(n595) );
  NAND2_X1 U669 ( .A1(n656), .A2(G92), .ZN(n593) );
  XNOR2_X1 U670 ( .A(KEYINPUT70), .B(n593), .ZN(n594) );
  NAND2_X1 U671 ( .A1(n595), .A2(n594), .ZN(n596) );
  INV_X1 U672 ( .A(n995), .ZN(n635) );
  NOR2_X1 U673 ( .A1(n635), .A2(G868), .ZN(n600) );
  XNOR2_X1 U674 ( .A(n600), .B(KEYINPUT74), .ZN(n602) );
  INV_X1 U675 ( .A(G868), .ZN(n682) );
  NOR2_X1 U676 ( .A1(n682), .A2(G171), .ZN(n601) );
  NOR2_X1 U677 ( .A1(n602), .A2(n601), .ZN(n603) );
  XNOR2_X1 U678 ( .A(KEYINPUT75), .B(n603), .ZN(G284) );
  INV_X1 U679 ( .A(G171), .ZN(G301) );
  NAND2_X1 U680 ( .A1(G63), .A2(n670), .ZN(n605) );
  NAND2_X1 U681 ( .A1(G51), .A2(n664), .ZN(n604) );
  NAND2_X1 U682 ( .A1(n605), .A2(n604), .ZN(n606) );
  NAND2_X1 U683 ( .A1(n656), .A2(G89), .ZN(n607) );
  XNOR2_X1 U684 ( .A(n607), .B(KEYINPUT4), .ZN(n609) );
  NAND2_X1 U685 ( .A1(G76), .A2(n653), .ZN(n608) );
  NAND2_X1 U686 ( .A1(n609), .A2(n608), .ZN(n610) );
  XNOR2_X1 U687 ( .A(KEYINPUT76), .B(n612), .ZN(G168) );
  XOR2_X1 U688 ( .A(KEYINPUT8), .B(G168), .Z(G286) );
  NAND2_X1 U689 ( .A1(G65), .A2(n670), .ZN(n614) );
  NAND2_X1 U690 ( .A1(G53), .A2(n664), .ZN(n613) );
  NAND2_X1 U691 ( .A1(n614), .A2(n613), .ZN(n618) );
  NAND2_X1 U692 ( .A1(G91), .A2(n656), .ZN(n616) );
  NAND2_X1 U693 ( .A1(G78), .A2(n653), .ZN(n615) );
  NAND2_X1 U694 ( .A1(n616), .A2(n615), .ZN(n617) );
  NOR2_X1 U695 ( .A1(n618), .A2(n617), .ZN(n988) );
  INV_X1 U696 ( .A(n988), .ZN(G299) );
  NAND2_X1 U697 ( .A1(G868), .A2(G286), .ZN(n620) );
  NAND2_X1 U698 ( .A1(G299), .A2(n682), .ZN(n619) );
  NAND2_X1 U699 ( .A1(n620), .A2(n619), .ZN(G297) );
  NAND2_X1 U700 ( .A1(n637), .A2(G559), .ZN(n621) );
  NAND2_X1 U701 ( .A1(n621), .A2(n635), .ZN(n622) );
  XNOR2_X1 U702 ( .A(n622), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U703 ( .A1(G868), .A2(n1001), .ZN(n625) );
  NAND2_X1 U704 ( .A1(G868), .A2(n635), .ZN(n623) );
  NOR2_X1 U705 ( .A1(G559), .A2(n623), .ZN(n624) );
  NOR2_X1 U706 ( .A1(n625), .A2(n624), .ZN(G282) );
  NAND2_X1 U707 ( .A1(n885), .A2(G123), .ZN(n626) );
  XNOR2_X1 U708 ( .A(n626), .B(KEYINPUT18), .ZN(n628) );
  NAND2_X1 U709 ( .A1(G111), .A2(n888), .ZN(n627) );
  NAND2_X1 U710 ( .A1(n628), .A2(n627), .ZN(n632) );
  NAND2_X1 U711 ( .A1(G135), .A2(n879), .ZN(n630) );
  NAND2_X1 U712 ( .A1(G99), .A2(n881), .ZN(n629) );
  NAND2_X1 U713 ( .A1(n630), .A2(n629), .ZN(n631) );
  NOR2_X1 U714 ( .A1(n632), .A2(n631), .ZN(n946) );
  XNOR2_X1 U715 ( .A(G2096), .B(n946), .ZN(n634) );
  INV_X1 U716 ( .A(G2100), .ZN(n633) );
  NAND2_X1 U717 ( .A1(n634), .A2(n633), .ZN(G156) );
  NAND2_X1 U718 ( .A1(G559), .A2(n635), .ZN(n636) );
  XOR2_X1 U719 ( .A(n1001), .B(n636), .Z(n679) );
  NAND2_X1 U720 ( .A1(n637), .A2(n679), .ZN(n645) );
  NAND2_X1 U721 ( .A1(G67), .A2(n670), .ZN(n639) );
  NAND2_X1 U722 ( .A1(G55), .A2(n664), .ZN(n638) );
  NAND2_X1 U723 ( .A1(n639), .A2(n638), .ZN(n644) );
  NAND2_X1 U724 ( .A1(G93), .A2(n656), .ZN(n641) );
  NAND2_X1 U725 ( .A1(G80), .A2(n653), .ZN(n640) );
  NAND2_X1 U726 ( .A1(n641), .A2(n640), .ZN(n642) );
  XOR2_X1 U727 ( .A(KEYINPUT77), .B(n642), .Z(n643) );
  NOR2_X1 U728 ( .A1(n644), .A2(n643), .ZN(n681) );
  XOR2_X1 U729 ( .A(n645), .B(n681), .Z(G145) );
  NAND2_X1 U730 ( .A1(G85), .A2(n656), .ZN(n647) );
  NAND2_X1 U731 ( .A1(G72), .A2(n653), .ZN(n646) );
  NAND2_X1 U732 ( .A1(n647), .A2(n646), .ZN(n648) );
  XNOR2_X1 U733 ( .A(KEYINPUT65), .B(n648), .ZN(n652) );
  NAND2_X1 U734 ( .A1(n664), .A2(G47), .ZN(n650) );
  NAND2_X1 U735 ( .A1(G60), .A2(n670), .ZN(n649) );
  AND2_X1 U736 ( .A1(n650), .A2(n649), .ZN(n651) );
  NAND2_X1 U737 ( .A1(n652), .A2(n651), .ZN(G290) );
  XOR2_X1 U738 ( .A(KEYINPUT79), .B(KEYINPUT2), .Z(n655) );
  NAND2_X1 U739 ( .A1(G73), .A2(n653), .ZN(n654) );
  XNOR2_X1 U740 ( .A(n655), .B(n654), .ZN(n663) );
  NAND2_X1 U741 ( .A1(G86), .A2(n656), .ZN(n658) );
  NAND2_X1 U742 ( .A1(G61), .A2(n670), .ZN(n657) );
  NAND2_X1 U743 ( .A1(n658), .A2(n657), .ZN(n661) );
  NAND2_X1 U744 ( .A1(n664), .A2(G48), .ZN(n659) );
  XOR2_X1 U745 ( .A(KEYINPUT80), .B(n659), .Z(n660) );
  NOR2_X1 U746 ( .A1(n661), .A2(n660), .ZN(n662) );
  NAND2_X1 U747 ( .A1(n663), .A2(n662), .ZN(G305) );
  NAND2_X1 U748 ( .A1(n664), .A2(G49), .ZN(n665) );
  XNOR2_X1 U749 ( .A(n665), .B(KEYINPUT78), .ZN(n672) );
  NAND2_X1 U750 ( .A1(G87), .A2(n666), .ZN(n668) );
  NAND2_X1 U751 ( .A1(G74), .A2(G651), .ZN(n667) );
  NAND2_X1 U752 ( .A1(n668), .A2(n667), .ZN(n669) );
  NOR2_X1 U753 ( .A1(n670), .A2(n669), .ZN(n671) );
  NAND2_X1 U754 ( .A1(n672), .A2(n671), .ZN(G288) );
  XNOR2_X1 U755 ( .A(G166), .B(G290), .ZN(n678) );
  XNOR2_X1 U756 ( .A(KEYINPUT82), .B(KEYINPUT19), .ZN(n674) );
  XNOR2_X1 U757 ( .A(G305), .B(n988), .ZN(n673) );
  XNOR2_X1 U758 ( .A(n674), .B(n673), .ZN(n675) );
  XNOR2_X1 U759 ( .A(n681), .B(n675), .ZN(n676) );
  XNOR2_X1 U760 ( .A(n676), .B(G288), .ZN(n677) );
  XNOR2_X1 U761 ( .A(n678), .B(n677), .ZN(n898) );
  XOR2_X1 U762 ( .A(n898), .B(n679), .Z(n680) );
  NOR2_X1 U763 ( .A1(n682), .A2(n680), .ZN(n684) );
  AND2_X1 U764 ( .A1(n682), .A2(n681), .ZN(n683) );
  NOR2_X1 U765 ( .A1(n684), .A2(n683), .ZN(G295) );
  NAND2_X1 U766 ( .A1(G2078), .A2(G2084), .ZN(n685) );
  XOR2_X1 U767 ( .A(KEYINPUT20), .B(n685), .Z(n686) );
  NAND2_X1 U768 ( .A1(G2090), .A2(n686), .ZN(n687) );
  XNOR2_X1 U769 ( .A(KEYINPUT21), .B(n687), .ZN(n688) );
  NAND2_X1 U770 ( .A1(n688), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U771 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U772 ( .A1(G236), .A2(G238), .ZN(n689) );
  NAND2_X1 U773 ( .A1(G69), .A2(n689), .ZN(n690) );
  NOR2_X1 U774 ( .A1(n690), .A2(G237), .ZN(n691) );
  XNOR2_X1 U775 ( .A(n691), .B(KEYINPUT85), .ZN(n850) );
  NAND2_X1 U776 ( .A1(n850), .A2(G567), .ZN(n698) );
  XOR2_X1 U777 ( .A(KEYINPUT83), .B(KEYINPUT22), .Z(n693) );
  NAND2_X1 U778 ( .A1(G132), .A2(G82), .ZN(n692) );
  XNOR2_X1 U779 ( .A(n693), .B(n692), .ZN(n694) );
  NOR2_X1 U780 ( .A1(G218), .A2(n694), .ZN(n695) );
  NAND2_X1 U781 ( .A1(G96), .A2(n695), .ZN(n696) );
  XNOR2_X1 U782 ( .A(KEYINPUT84), .B(n696), .ZN(n851) );
  NAND2_X1 U783 ( .A1(n851), .A2(G2106), .ZN(n697) );
  NAND2_X1 U784 ( .A1(n698), .A2(n697), .ZN(n930) );
  NAND2_X1 U785 ( .A1(G483), .A2(G661), .ZN(n699) );
  NOR2_X1 U786 ( .A1(n930), .A2(n699), .ZN(n849) );
  NAND2_X1 U787 ( .A1(n849), .A2(G36), .ZN(G176) );
  INV_X1 U788 ( .A(G166), .ZN(G303) );
  XNOR2_X1 U789 ( .A(KEYINPUT40), .B(KEYINPUT102), .ZN(n845) );
  INV_X1 U790 ( .A(KEYINPUT90), .ZN(n704) );
  INV_X1 U791 ( .A(G40), .ZN(n700) );
  OR2_X1 U792 ( .A1(n701), .A2(n700), .ZN(n702) );
  NOR2_X1 U793 ( .A1(G164), .A2(G1384), .ZN(n797) );
  NAND2_X2 U794 ( .A1(n705), .A2(n797), .ZN(n755) );
  NOR2_X1 U795 ( .A1(G2084), .A2(n755), .ZN(n735) );
  NAND2_X1 U796 ( .A1(G8), .A2(n735), .ZN(n706) );
  XOR2_X1 U797 ( .A(KEYINPUT92), .B(n706), .Z(n751) );
  NAND2_X1 U798 ( .A1(G1348), .A2(n755), .ZN(n708) );
  INV_X2 U799 ( .A(n755), .ZN(n729) );
  NAND2_X1 U800 ( .A1(G2067), .A2(n729), .ZN(n707) );
  NAND2_X1 U801 ( .A1(n708), .A2(n707), .ZN(n716) );
  INV_X1 U802 ( .A(G1996), .ZN(n959) );
  NOR2_X1 U803 ( .A1(n755), .A2(n959), .ZN(n710) );
  XNOR2_X1 U804 ( .A(n710), .B(n709), .ZN(n712) );
  NAND2_X1 U805 ( .A1(n755), .A2(G1341), .ZN(n711) );
  NAND2_X1 U806 ( .A1(n712), .A2(n711), .ZN(n713) );
  OR2_X1 U807 ( .A1(n1001), .A2(n713), .ZN(n714) );
  NAND2_X1 U808 ( .A1(n715), .A2(n714), .ZN(n718) );
  NAND2_X1 U809 ( .A1(n995), .A2(n716), .ZN(n717) );
  NAND2_X1 U810 ( .A1(n718), .A2(n717), .ZN(n723) );
  NAND2_X1 U811 ( .A1(n729), .A2(G2072), .ZN(n719) );
  XNOR2_X1 U812 ( .A(n719), .B(KEYINPUT27), .ZN(n721) );
  INV_X1 U813 ( .A(G1956), .ZN(n1013) );
  NOR2_X1 U814 ( .A1(n1013), .A2(n729), .ZN(n720) );
  NOR2_X1 U815 ( .A1(n721), .A2(n720), .ZN(n724) );
  NAND2_X1 U816 ( .A1(n988), .A2(n724), .ZN(n722) );
  NAND2_X1 U817 ( .A1(n723), .A2(n722), .ZN(n726) );
  NOR2_X1 U818 ( .A1(n988), .A2(n724), .ZN(n725) );
  NAND2_X1 U819 ( .A1(n726), .A2(n526), .ZN(n728) );
  XOR2_X1 U820 ( .A(KEYINPUT29), .B(KEYINPUT93), .Z(n727) );
  XNOR2_X1 U821 ( .A(n728), .B(n727), .ZN(n733) );
  NAND2_X1 U822 ( .A1(G1961), .A2(n755), .ZN(n731) );
  XOR2_X1 U823 ( .A(G2078), .B(KEYINPUT25), .Z(n961) );
  NAND2_X1 U824 ( .A1(n729), .A2(n961), .ZN(n730) );
  NAND2_X1 U825 ( .A1(n731), .A2(n730), .ZN(n734) );
  NOR2_X1 U826 ( .A1(G301), .A2(n734), .ZN(n732) );
  NOR2_X1 U827 ( .A1(n733), .A2(n732), .ZN(n744) );
  AND2_X1 U828 ( .A1(G301), .A2(n734), .ZN(n741) );
  NOR2_X1 U829 ( .A1(G1966), .A2(n753), .ZN(n746) );
  NOR2_X1 U830 ( .A1(n746), .A2(n735), .ZN(n736) );
  XNOR2_X1 U831 ( .A(n736), .B(KEYINPUT94), .ZN(n737) );
  NAND2_X1 U832 ( .A1(n737), .A2(G8), .ZN(n738) );
  XNOR2_X1 U833 ( .A(n738), .B(KEYINPUT30), .ZN(n739) );
  NOR2_X1 U834 ( .A1(n739), .A2(G168), .ZN(n740) );
  NOR2_X1 U835 ( .A1(n741), .A2(n740), .ZN(n742) );
  XNOR2_X1 U836 ( .A(n742), .B(KEYINPUT31), .ZN(n743) );
  NOR2_X1 U837 ( .A1(n744), .A2(n743), .ZN(n745) );
  XNOR2_X1 U838 ( .A(n745), .B(KEYINPUT95), .ZN(n759) );
  INV_X1 U839 ( .A(n759), .ZN(n747) );
  NOR2_X1 U840 ( .A1(n747), .A2(n746), .ZN(n749) );
  XNOR2_X1 U841 ( .A(n749), .B(n748), .ZN(n750) );
  NOR2_X1 U842 ( .A1(n751), .A2(n750), .ZN(n752) );
  XNOR2_X1 U843 ( .A(n752), .B(KEYINPUT97), .ZN(n765) );
  NOR2_X1 U844 ( .A1(G1971), .A2(n791), .ZN(n754) );
  XNOR2_X1 U845 ( .A(n754), .B(KEYINPUT98), .ZN(n757) );
  NOR2_X1 U846 ( .A1(n755), .A2(G2090), .ZN(n756) );
  NOR2_X1 U847 ( .A1(n757), .A2(n756), .ZN(n758) );
  NAND2_X1 U848 ( .A1(G303), .A2(n758), .ZN(n761) );
  NAND2_X1 U849 ( .A1(n759), .A2(G286), .ZN(n760) );
  NAND2_X1 U850 ( .A1(n761), .A2(n760), .ZN(n762) );
  NAND2_X1 U851 ( .A1(n762), .A2(G8), .ZN(n763) );
  XNOR2_X1 U852 ( .A(KEYINPUT32), .B(n763), .ZN(n764) );
  NAND2_X1 U853 ( .A1(n765), .A2(n764), .ZN(n783) );
  NOR2_X1 U854 ( .A1(G1976), .A2(G288), .ZN(n984) );
  NOR2_X1 U855 ( .A1(G1971), .A2(G303), .ZN(n766) );
  NOR2_X1 U856 ( .A1(n984), .A2(n766), .ZN(n767) );
  NAND2_X1 U857 ( .A1(n783), .A2(n767), .ZN(n769) );
  NAND2_X1 U858 ( .A1(G288), .A2(G1976), .ZN(n768) );
  XOR2_X1 U859 ( .A(KEYINPUT99), .B(n768), .Z(n985) );
  NAND2_X1 U860 ( .A1(n769), .A2(n985), .ZN(n770) );
  XNOR2_X1 U861 ( .A(KEYINPUT100), .B(n770), .ZN(n772) );
  OR2_X1 U862 ( .A1(n791), .A2(KEYINPUT101), .ZN(n771) );
  NOR2_X1 U863 ( .A1(n772), .A2(n771), .ZN(n773) );
  NOR2_X1 U864 ( .A1(n773), .A2(KEYINPUT33), .ZN(n774) );
  INV_X1 U865 ( .A(n774), .ZN(n782) );
  XOR2_X1 U866 ( .A(G1981), .B(G305), .Z(n1002) );
  INV_X1 U867 ( .A(KEYINPUT101), .ZN(n776) );
  NAND2_X1 U868 ( .A1(n984), .A2(KEYINPUT33), .ZN(n775) );
  NAND2_X1 U869 ( .A1(n776), .A2(n775), .ZN(n778) );
  NAND2_X1 U870 ( .A1(n984), .A2(KEYINPUT101), .ZN(n777) );
  NAND2_X1 U871 ( .A1(n778), .A2(n777), .ZN(n779) );
  NOR2_X1 U872 ( .A1(n791), .A2(n779), .ZN(n780) );
  NAND2_X1 U873 ( .A1(n782), .A2(n527), .ZN(n788) );
  NOR2_X1 U874 ( .A1(G2090), .A2(G303), .ZN(n784) );
  NAND2_X1 U875 ( .A1(G8), .A2(n784), .ZN(n785) );
  NAND2_X1 U876 ( .A1(n783), .A2(n785), .ZN(n786) );
  NAND2_X1 U877 ( .A1(n786), .A2(n791), .ZN(n787) );
  NAND2_X1 U878 ( .A1(n788), .A2(n787), .ZN(n794) );
  NOR2_X1 U879 ( .A1(G1981), .A2(G305), .ZN(n789) );
  XOR2_X1 U880 ( .A(n789), .B(KEYINPUT24), .Z(n790) );
  NOR2_X1 U881 ( .A1(n791), .A2(n790), .ZN(n792) );
  XOR2_X1 U882 ( .A(KEYINPUT91), .B(n792), .Z(n793) );
  NOR2_X1 U883 ( .A1(n794), .A2(n793), .ZN(n795) );
  INV_X1 U884 ( .A(n795), .ZN(n829) );
  NOR2_X1 U885 ( .A1(n797), .A2(n796), .ZN(n840) );
  NAND2_X1 U886 ( .A1(G140), .A2(n879), .ZN(n799) );
  NAND2_X1 U887 ( .A1(G104), .A2(n881), .ZN(n798) );
  NAND2_X1 U888 ( .A1(n799), .A2(n798), .ZN(n800) );
  XNOR2_X1 U889 ( .A(KEYINPUT34), .B(n800), .ZN(n805) );
  NAND2_X1 U890 ( .A1(G128), .A2(n885), .ZN(n802) );
  NAND2_X1 U891 ( .A1(G116), .A2(n888), .ZN(n801) );
  NAND2_X1 U892 ( .A1(n802), .A2(n801), .ZN(n803) );
  XOR2_X1 U893 ( .A(KEYINPUT35), .B(n803), .Z(n804) );
  NOR2_X1 U894 ( .A1(n805), .A2(n804), .ZN(n806) );
  XNOR2_X1 U895 ( .A(KEYINPUT36), .B(n806), .ZN(n893) );
  XNOR2_X1 U896 ( .A(G2067), .B(KEYINPUT37), .ZN(n838) );
  NOR2_X1 U897 ( .A1(n893), .A2(n838), .ZN(n937) );
  NAND2_X1 U898 ( .A1(n840), .A2(n937), .ZN(n836) );
  XOR2_X1 U899 ( .A(KEYINPUT88), .B(KEYINPUT38), .Z(n808) );
  NAND2_X1 U900 ( .A1(G105), .A2(n881), .ZN(n807) );
  XNOR2_X1 U901 ( .A(n808), .B(n807), .ZN(n812) );
  NAND2_X1 U902 ( .A1(G141), .A2(n879), .ZN(n810) );
  NAND2_X1 U903 ( .A1(G129), .A2(n885), .ZN(n809) );
  NAND2_X1 U904 ( .A1(n810), .A2(n809), .ZN(n811) );
  NOR2_X1 U905 ( .A1(n812), .A2(n811), .ZN(n814) );
  NAND2_X1 U906 ( .A1(n888), .A2(G117), .ZN(n813) );
  NAND2_X1 U907 ( .A1(n814), .A2(n813), .ZN(n875) );
  NAND2_X1 U908 ( .A1(G1996), .A2(n875), .ZN(n824) );
  NAND2_X1 U909 ( .A1(G131), .A2(n879), .ZN(n816) );
  NAND2_X1 U910 ( .A1(G95), .A2(n881), .ZN(n815) );
  NAND2_X1 U911 ( .A1(n816), .A2(n815), .ZN(n821) );
  NAND2_X1 U912 ( .A1(G119), .A2(n885), .ZN(n818) );
  NAND2_X1 U913 ( .A1(G107), .A2(n888), .ZN(n817) );
  NAND2_X1 U914 ( .A1(n818), .A2(n817), .ZN(n819) );
  XNOR2_X1 U915 ( .A(KEYINPUT86), .B(n819), .ZN(n820) );
  NOR2_X1 U916 ( .A1(n821), .A2(n820), .ZN(n822) );
  XNOR2_X1 U917 ( .A(n822), .B(KEYINPUT87), .ZN(n869) );
  NAND2_X1 U918 ( .A1(G1991), .A2(n869), .ZN(n823) );
  NAND2_X1 U919 ( .A1(n824), .A2(n823), .ZN(n825) );
  XNOR2_X1 U920 ( .A(KEYINPUT89), .B(n825), .ZN(n943) );
  INV_X1 U921 ( .A(n943), .ZN(n826) );
  NAND2_X1 U922 ( .A1(n826), .A2(n840), .ZN(n830) );
  NAND2_X1 U923 ( .A1(n836), .A2(n830), .ZN(n827) );
  XNOR2_X1 U924 ( .A(G1986), .B(G290), .ZN(n992) );
  NAND2_X1 U925 ( .A1(n829), .A2(n828), .ZN(n843) );
  NOR2_X1 U926 ( .A1(G1996), .A2(n875), .ZN(n932) );
  INV_X1 U927 ( .A(n830), .ZN(n833) );
  NOR2_X1 U928 ( .A1(G1991), .A2(n869), .ZN(n945) );
  NOR2_X1 U929 ( .A1(G1986), .A2(G290), .ZN(n831) );
  NOR2_X1 U930 ( .A1(n945), .A2(n831), .ZN(n832) );
  NOR2_X1 U931 ( .A1(n833), .A2(n832), .ZN(n834) );
  NOR2_X1 U932 ( .A1(n932), .A2(n834), .ZN(n835) );
  XNOR2_X1 U933 ( .A(n835), .B(KEYINPUT39), .ZN(n837) );
  NAND2_X1 U934 ( .A1(n837), .A2(n836), .ZN(n839) );
  NAND2_X1 U935 ( .A1(n893), .A2(n838), .ZN(n936) );
  NAND2_X1 U936 ( .A1(n839), .A2(n936), .ZN(n841) );
  NAND2_X1 U937 ( .A1(n841), .A2(n840), .ZN(n842) );
  NAND2_X1 U938 ( .A1(n843), .A2(n842), .ZN(n844) );
  XNOR2_X1 U939 ( .A(n845), .B(n844), .ZN(G329) );
  NAND2_X1 U940 ( .A1(G2106), .A2(n846), .ZN(G217) );
  AND2_X1 U941 ( .A1(G15), .A2(G2), .ZN(n847) );
  NAND2_X1 U942 ( .A1(G661), .A2(n847), .ZN(G259) );
  NAND2_X1 U943 ( .A1(G3), .A2(G1), .ZN(n848) );
  NAND2_X1 U944 ( .A1(n849), .A2(n848), .ZN(G188) );
  INV_X1 U946 ( .A(G132), .ZN(G219) );
  INV_X1 U947 ( .A(G96), .ZN(G221) );
  INV_X1 U948 ( .A(G82), .ZN(G220) );
  NOR2_X1 U949 ( .A1(n851), .A2(n850), .ZN(G325) );
  INV_X1 U950 ( .A(G325), .ZN(G261) );
  NAND2_X1 U951 ( .A1(n885), .A2(G124), .ZN(n852) );
  XNOR2_X1 U952 ( .A(n852), .B(KEYINPUT44), .ZN(n854) );
  NAND2_X1 U953 ( .A1(G112), .A2(n888), .ZN(n853) );
  NAND2_X1 U954 ( .A1(n854), .A2(n853), .ZN(n858) );
  NAND2_X1 U955 ( .A1(G136), .A2(n879), .ZN(n856) );
  NAND2_X1 U956 ( .A1(G100), .A2(n881), .ZN(n855) );
  NAND2_X1 U957 ( .A1(n856), .A2(n855), .ZN(n857) );
  NOR2_X1 U958 ( .A1(n858), .A2(n857), .ZN(G162) );
  NAND2_X1 U959 ( .A1(n881), .A2(G103), .ZN(n859) );
  XNOR2_X1 U960 ( .A(KEYINPUT109), .B(n859), .ZN(n867) );
  NAND2_X1 U961 ( .A1(G127), .A2(n885), .ZN(n861) );
  NAND2_X1 U962 ( .A1(G115), .A2(n888), .ZN(n860) );
  NAND2_X1 U963 ( .A1(n861), .A2(n860), .ZN(n862) );
  XNOR2_X1 U964 ( .A(n862), .B(KEYINPUT47), .ZN(n863) );
  XNOR2_X1 U965 ( .A(n863), .B(KEYINPUT110), .ZN(n865) );
  NAND2_X1 U966 ( .A1(n879), .A2(G139), .ZN(n864) );
  NAND2_X1 U967 ( .A1(n865), .A2(n864), .ZN(n866) );
  NOR2_X1 U968 ( .A1(n867), .A2(n866), .ZN(n939) );
  XOR2_X1 U969 ( .A(G164), .B(n939), .Z(n868) );
  XNOR2_X1 U970 ( .A(n869), .B(n868), .ZN(n873) );
  XOR2_X1 U971 ( .A(KEYINPUT46), .B(KEYINPUT111), .Z(n871) );
  XNOR2_X1 U972 ( .A(KEYINPUT112), .B(KEYINPUT48), .ZN(n870) );
  XNOR2_X1 U973 ( .A(n871), .B(n870), .ZN(n872) );
  XOR2_X1 U974 ( .A(n873), .B(n872), .Z(n878) );
  XOR2_X1 U975 ( .A(n946), .B(G162), .Z(n874) );
  XNOR2_X1 U976 ( .A(n875), .B(n874), .ZN(n876) );
  XNOR2_X1 U977 ( .A(G160), .B(n876), .ZN(n877) );
  XNOR2_X1 U978 ( .A(n878), .B(n877), .ZN(n895) );
  NAND2_X1 U979 ( .A1(n879), .A2(G142), .ZN(n880) );
  XNOR2_X1 U980 ( .A(n880), .B(KEYINPUT108), .ZN(n883) );
  NAND2_X1 U981 ( .A1(G106), .A2(n881), .ZN(n882) );
  NAND2_X1 U982 ( .A1(n883), .A2(n882), .ZN(n884) );
  XNOR2_X1 U983 ( .A(n884), .B(KEYINPUT45), .ZN(n887) );
  NAND2_X1 U984 ( .A1(G130), .A2(n885), .ZN(n886) );
  NAND2_X1 U985 ( .A1(n887), .A2(n886), .ZN(n891) );
  NAND2_X1 U986 ( .A1(G118), .A2(n888), .ZN(n889) );
  XNOR2_X1 U987 ( .A(KEYINPUT107), .B(n889), .ZN(n890) );
  NOR2_X1 U988 ( .A1(n891), .A2(n890), .ZN(n892) );
  XOR2_X1 U989 ( .A(n893), .B(n892), .Z(n894) );
  XNOR2_X1 U990 ( .A(n895), .B(n894), .ZN(n896) );
  NOR2_X1 U991 ( .A1(G37), .A2(n896), .ZN(G395) );
  XNOR2_X1 U992 ( .A(G171), .B(n1001), .ZN(n897) );
  XNOR2_X1 U993 ( .A(n897), .B(G286), .ZN(n900) );
  XNOR2_X1 U994 ( .A(n995), .B(n898), .ZN(n899) );
  XNOR2_X1 U995 ( .A(n900), .B(n899), .ZN(n901) );
  NOR2_X1 U996 ( .A1(G37), .A2(n901), .ZN(G397) );
  XNOR2_X1 U997 ( .A(G1966), .B(G2474), .ZN(n911) );
  XOR2_X1 U998 ( .A(G1961), .B(G1976), .Z(n903) );
  XNOR2_X1 U999 ( .A(G1986), .B(G1981), .ZN(n902) );
  XNOR2_X1 U1000 ( .A(n903), .B(n902), .ZN(n907) );
  XOR2_X1 U1001 ( .A(G1956), .B(G1971), .Z(n905) );
  XNOR2_X1 U1002 ( .A(G1996), .B(G1991), .ZN(n904) );
  XNOR2_X1 U1003 ( .A(n905), .B(n904), .ZN(n906) );
  XOR2_X1 U1004 ( .A(n907), .B(n906), .Z(n909) );
  XNOR2_X1 U1005 ( .A(KEYINPUT106), .B(KEYINPUT41), .ZN(n908) );
  XNOR2_X1 U1006 ( .A(n909), .B(n908), .ZN(n910) );
  XNOR2_X1 U1007 ( .A(n911), .B(n910), .ZN(G229) );
  XNOR2_X1 U1008 ( .A(G2067), .B(G2090), .ZN(n912) );
  XNOR2_X1 U1009 ( .A(n912), .B(KEYINPUT103), .ZN(n922) );
  XOR2_X1 U1010 ( .A(KEYINPUT104), .B(KEYINPUT105), .Z(n914) );
  XNOR2_X1 U1011 ( .A(KEYINPUT42), .B(G2096), .ZN(n913) );
  XNOR2_X1 U1012 ( .A(n914), .B(n913), .ZN(n918) );
  XOR2_X1 U1013 ( .A(G2100), .B(G2084), .Z(n916) );
  XNOR2_X1 U1014 ( .A(G2072), .B(G2078), .ZN(n915) );
  XNOR2_X1 U1015 ( .A(n916), .B(n915), .ZN(n917) );
  XOR2_X1 U1016 ( .A(n918), .B(n917), .Z(n920) );
  XNOR2_X1 U1017 ( .A(G2678), .B(KEYINPUT43), .ZN(n919) );
  XNOR2_X1 U1018 ( .A(n920), .B(n919), .ZN(n921) );
  XNOR2_X1 U1019 ( .A(n922), .B(n921), .ZN(G227) );
  NOR2_X1 U1020 ( .A1(G395), .A2(G397), .ZN(n923) );
  XNOR2_X1 U1021 ( .A(KEYINPUT114), .B(n923), .ZN(n929) );
  NOR2_X1 U1022 ( .A1(n930), .A2(G401), .ZN(n924) );
  XNOR2_X1 U1023 ( .A(n924), .B(KEYINPUT113), .ZN(n927) );
  NOR2_X1 U1024 ( .A1(G229), .A2(G227), .ZN(n925) );
  XNOR2_X1 U1025 ( .A(KEYINPUT49), .B(n925), .ZN(n926) );
  NOR2_X1 U1026 ( .A1(n927), .A2(n926), .ZN(n928) );
  NAND2_X1 U1027 ( .A1(n929), .A2(n928), .ZN(G225) );
  INV_X1 U1028 ( .A(G225), .ZN(G308) );
  INV_X1 U1029 ( .A(n930), .ZN(G319) );
  INV_X1 U1030 ( .A(G69), .ZN(G235) );
  XNOR2_X1 U1031 ( .A(G160), .B(G2084), .ZN(n935) );
  XOR2_X1 U1032 ( .A(G2090), .B(G162), .Z(n931) );
  NOR2_X1 U1033 ( .A1(n932), .A2(n931), .ZN(n933) );
  XOR2_X1 U1034 ( .A(KEYINPUT51), .B(n933), .Z(n934) );
  NAND2_X1 U1035 ( .A1(n935), .A2(n934), .ZN(n953) );
  INV_X1 U1036 ( .A(n936), .ZN(n938) );
  NOR2_X1 U1037 ( .A1(n938), .A2(n937), .ZN(n951) );
  XOR2_X1 U1038 ( .A(G2072), .B(n939), .Z(n941) );
  XOR2_X1 U1039 ( .A(G164), .B(G2078), .Z(n940) );
  NOR2_X1 U1040 ( .A1(n941), .A2(n940), .ZN(n942) );
  XNOR2_X1 U1041 ( .A(KEYINPUT50), .B(n942), .ZN(n944) );
  NAND2_X1 U1042 ( .A1(n944), .A2(n943), .ZN(n949) );
  NOR2_X1 U1043 ( .A1(n946), .A2(n945), .ZN(n947) );
  XNOR2_X1 U1044 ( .A(KEYINPUT115), .B(n947), .ZN(n948) );
  NOR2_X1 U1045 ( .A1(n949), .A2(n948), .ZN(n950) );
  NAND2_X1 U1046 ( .A1(n951), .A2(n950), .ZN(n952) );
  NOR2_X1 U1047 ( .A1(n953), .A2(n952), .ZN(n954) );
  XNOR2_X1 U1048 ( .A(KEYINPUT52), .B(n954), .ZN(n955) );
  XOR2_X1 U1049 ( .A(KEYINPUT55), .B(KEYINPUT116), .Z(n980) );
  NAND2_X1 U1050 ( .A1(n955), .A2(n980), .ZN(n956) );
  NAND2_X1 U1051 ( .A1(n956), .A2(G29), .ZN(n1043) );
  XNOR2_X1 U1052 ( .A(KEYINPUT54), .B(KEYINPUT121), .ZN(n957) );
  XNOR2_X1 U1053 ( .A(n957), .B(G34), .ZN(n958) );
  XNOR2_X1 U1054 ( .A(G2084), .B(n958), .ZN(n978) );
  XNOR2_X1 U1055 ( .A(G2090), .B(G35), .ZN(n976) );
  XNOR2_X1 U1056 ( .A(KEYINPUT119), .B(G32), .ZN(n960) );
  XNOR2_X1 U1057 ( .A(n960), .B(n959), .ZN(n963) );
  XNOR2_X1 U1058 ( .A(G27), .B(n961), .ZN(n962) );
  NOR2_X1 U1059 ( .A1(n963), .A2(n962), .ZN(n964) );
  XNOR2_X1 U1060 ( .A(KEYINPUT120), .B(n964), .ZN(n968) );
  XNOR2_X1 U1061 ( .A(G2067), .B(G26), .ZN(n966) );
  XNOR2_X1 U1062 ( .A(G33), .B(G2072), .ZN(n965) );
  NOR2_X1 U1063 ( .A1(n966), .A2(n965), .ZN(n967) );
  NAND2_X1 U1064 ( .A1(n968), .A2(n967), .ZN(n973) );
  XNOR2_X1 U1065 ( .A(G1991), .B(G25), .ZN(n969) );
  XNOR2_X1 U1066 ( .A(n969), .B(KEYINPUT117), .ZN(n970) );
  NAND2_X1 U1067 ( .A1(G28), .A2(n970), .ZN(n971) );
  XNOR2_X1 U1068 ( .A(KEYINPUT118), .B(n971), .ZN(n972) );
  NOR2_X1 U1069 ( .A1(n973), .A2(n972), .ZN(n974) );
  XNOR2_X1 U1070 ( .A(KEYINPUT53), .B(n974), .ZN(n975) );
  NOR2_X1 U1071 ( .A1(n976), .A2(n975), .ZN(n977) );
  NAND2_X1 U1072 ( .A1(n978), .A2(n977), .ZN(n979) );
  XNOR2_X1 U1073 ( .A(n980), .B(n979), .ZN(n982) );
  INV_X1 U1074 ( .A(G29), .ZN(n981) );
  NAND2_X1 U1075 ( .A1(n982), .A2(n981), .ZN(n983) );
  NAND2_X1 U1076 ( .A1(G11), .A2(n983), .ZN(n1041) );
  XNOR2_X1 U1077 ( .A(G16), .B(KEYINPUT56), .ZN(n1011) );
  INV_X1 U1078 ( .A(n984), .ZN(n986) );
  NAND2_X1 U1079 ( .A1(n986), .A2(n985), .ZN(n987) );
  XNOR2_X1 U1080 ( .A(n987), .B(KEYINPUT123), .ZN(n994) );
  XNOR2_X1 U1081 ( .A(n988), .B(G1956), .ZN(n990) );
  XNOR2_X1 U1082 ( .A(G1971), .B(G166), .ZN(n989) );
  NAND2_X1 U1083 ( .A1(n990), .A2(n989), .ZN(n991) );
  NOR2_X1 U1084 ( .A1(n992), .A2(n991), .ZN(n993) );
  NAND2_X1 U1085 ( .A1(n994), .A2(n993), .ZN(n999) );
  XOR2_X1 U1086 ( .A(n995), .B(G1348), .Z(n997) );
  XNOR2_X1 U1087 ( .A(G171), .B(G1961), .ZN(n996) );
  NAND2_X1 U1088 ( .A1(n997), .A2(n996), .ZN(n998) );
  NOR2_X1 U1089 ( .A1(n999), .A2(n998), .ZN(n1000) );
  XNOR2_X1 U1090 ( .A(KEYINPUT124), .B(n1000), .ZN(n1009) );
  XNOR2_X1 U1091 ( .A(n1001), .B(G1341), .ZN(n1007) );
  XNOR2_X1 U1092 ( .A(G1966), .B(G168), .ZN(n1003) );
  NAND2_X1 U1093 ( .A1(n1003), .A2(n1002), .ZN(n1005) );
  XOR2_X1 U1094 ( .A(KEYINPUT57), .B(KEYINPUT122), .Z(n1004) );
  XNOR2_X1 U1095 ( .A(n1005), .B(n1004), .ZN(n1006) );
  NOR2_X1 U1096 ( .A1(n1007), .A2(n1006), .ZN(n1008) );
  NAND2_X1 U1097 ( .A1(n1009), .A2(n1008), .ZN(n1010) );
  NAND2_X1 U1098 ( .A1(n1011), .A2(n1010), .ZN(n1039) );
  INV_X1 U1099 ( .A(G16), .ZN(n1037) );
  XNOR2_X1 U1100 ( .A(KEYINPUT61), .B(KEYINPUT127), .ZN(n1035) );
  XNOR2_X1 U1101 ( .A(KEYINPUT125), .B(G1966), .ZN(n1012) );
  XNOR2_X1 U1102 ( .A(n1012), .B(G21), .ZN(n1033) );
  XOR2_X1 U1103 ( .A(G1961), .B(G5), .Z(n1023) );
  XNOR2_X1 U1104 ( .A(G20), .B(n1013), .ZN(n1017) );
  XNOR2_X1 U1105 ( .A(G1981), .B(G6), .ZN(n1015) );
  XNOR2_X1 U1106 ( .A(G1341), .B(G19), .ZN(n1014) );
  NOR2_X1 U1107 ( .A1(n1015), .A2(n1014), .ZN(n1016) );
  NAND2_X1 U1108 ( .A1(n1017), .A2(n1016), .ZN(n1020) );
  XOR2_X1 U1109 ( .A(KEYINPUT59), .B(G1348), .Z(n1018) );
  XNOR2_X1 U1110 ( .A(G4), .B(n1018), .ZN(n1019) );
  NOR2_X1 U1111 ( .A1(n1020), .A2(n1019), .ZN(n1021) );
  XNOR2_X1 U1112 ( .A(KEYINPUT60), .B(n1021), .ZN(n1022) );
  NAND2_X1 U1113 ( .A1(n1023), .A2(n1022), .ZN(n1031) );
  XNOR2_X1 U1114 ( .A(G1986), .B(G24), .ZN(n1025) );
  XNOR2_X1 U1115 ( .A(G1971), .B(G22), .ZN(n1024) );
  NOR2_X1 U1116 ( .A1(n1025), .A2(n1024), .ZN(n1028) );
  XOR2_X1 U1117 ( .A(G1976), .B(KEYINPUT126), .Z(n1026) );
  XNOR2_X1 U1118 ( .A(G23), .B(n1026), .ZN(n1027) );
  NAND2_X1 U1119 ( .A1(n1028), .A2(n1027), .ZN(n1029) );
  XNOR2_X1 U1120 ( .A(KEYINPUT58), .B(n1029), .ZN(n1030) );
  NOR2_X1 U1121 ( .A1(n1031), .A2(n1030), .ZN(n1032) );
  NAND2_X1 U1122 ( .A1(n1033), .A2(n1032), .ZN(n1034) );
  XNOR2_X1 U1123 ( .A(n1035), .B(n1034), .ZN(n1036) );
  NAND2_X1 U1124 ( .A1(n1037), .A2(n1036), .ZN(n1038) );
  NAND2_X1 U1125 ( .A1(n1039), .A2(n1038), .ZN(n1040) );
  NOR2_X1 U1126 ( .A1(n1041), .A2(n1040), .ZN(n1042) );
  NAND2_X1 U1127 ( .A1(n1043), .A2(n1042), .ZN(n1044) );
  XOR2_X1 U1128 ( .A(KEYINPUT62), .B(n1044), .Z(G311) );
  INV_X1 U1129 ( .A(G311), .ZN(G150) );
endmodule

