//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 0 1 0 0 0 1 0 1 1 1 0 1 1 0 0 0 1 0 1 1 0 0 1 0 1 0 0 1 1 1 0 1 0 0 1 1 0 1 0 1 0 0 0 1 0 1 0 1 0 1 0 0 0 0 1 0 0 0 1 0 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:26:22 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n742, new_n743, new_n744, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n757, new_n758, new_n759, new_n761, new_n762,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n777, new_n778,
    new_n779, new_n780, new_n781, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n795, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n819, new_n820, new_n821, new_n822, new_n823, new_n824,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n946, new_n947, new_n948, new_n949, new_n950, new_n951, new_n952,
    new_n953, new_n954, new_n955, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n967, new_n968,
    new_n969, new_n971, new_n972, new_n973, new_n974, new_n975, new_n976,
    new_n977, new_n978, new_n979, new_n980, new_n982, new_n983, new_n984,
    new_n985, new_n986, new_n987, new_n988, new_n989, new_n990, new_n991,
    new_n992, new_n993, new_n995, new_n996, new_n997, new_n998, new_n999,
    new_n1000, new_n1001, new_n1002, new_n1003, new_n1004, new_n1005,
    new_n1006, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1022, new_n1023, new_n1024,
    new_n1025, new_n1026, new_n1027, new_n1028, new_n1029, new_n1030,
    new_n1031, new_n1033, new_n1034, new_n1035, new_n1036, new_n1037,
    new_n1038, new_n1039, new_n1040, new_n1041;
  XNOR2_X1  g000(.A(KEYINPUT9), .B(G234), .ZN(new_n187));
  INV_X1    g001(.A(G217), .ZN(new_n188));
  NOR3_X1   g002(.A1(new_n187), .A2(new_n188), .A3(G953), .ZN(new_n189));
  INV_X1    g003(.A(new_n189), .ZN(new_n190));
  OR2_X1    g004(.A1(KEYINPUT90), .A2(KEYINPUT13), .ZN(new_n191));
  INV_X1    g005(.A(G143), .ZN(new_n192));
  NAND2_X1  g006(.A1(KEYINPUT90), .A2(KEYINPUT13), .ZN(new_n193));
  NAND4_X1  g007(.A1(new_n191), .A2(G128), .A3(new_n192), .A4(new_n193), .ZN(new_n194));
  AND2_X1   g008(.A1(new_n191), .A2(new_n193), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n192), .A2(G128), .ZN(new_n196));
  INV_X1    g010(.A(G128), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n197), .A2(G143), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n196), .A2(new_n198), .ZN(new_n199));
  OAI211_X1 g013(.A(new_n194), .B(G134), .C1(new_n195), .C2(new_n199), .ZN(new_n200));
  INV_X1    g014(.A(G134), .ZN(new_n201));
  NAND3_X1  g015(.A1(new_n196), .A2(new_n198), .A3(new_n201), .ZN(new_n202));
  INV_X1    g016(.A(G107), .ZN(new_n203));
  INV_X1    g017(.A(G122), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n204), .A2(G116), .ZN(new_n205));
  INV_X1    g019(.A(G116), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n206), .A2(G122), .ZN(new_n207));
  AOI21_X1  g021(.A(new_n203), .B1(new_n205), .B2(new_n207), .ZN(new_n208));
  AND3_X1   g022(.A1(new_n205), .A2(new_n207), .A3(new_n203), .ZN(new_n209));
  OAI211_X1 g023(.A(new_n200), .B(new_n202), .C1(new_n208), .C2(new_n209), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n199), .A2(G134), .ZN(new_n211));
  AOI21_X1  g025(.A(new_n209), .B1(new_n211), .B2(new_n202), .ZN(new_n212));
  OAI21_X1  g026(.A(new_n205), .B1(new_n207), .B2(KEYINPUT14), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n207), .A2(KEYINPUT14), .ZN(new_n214));
  INV_X1    g028(.A(KEYINPUT91), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n214), .A2(new_n215), .ZN(new_n216));
  NAND3_X1  g030(.A1(new_n207), .A2(KEYINPUT91), .A3(KEYINPUT14), .ZN(new_n217));
  AOI21_X1  g031(.A(new_n213), .B1(new_n216), .B2(new_n217), .ZN(new_n218));
  OAI21_X1  g032(.A(new_n212), .B1(new_n218), .B2(new_n203), .ZN(new_n219));
  INV_X1    g033(.A(KEYINPUT92), .ZN(new_n220));
  NAND3_X1  g034(.A1(new_n210), .A2(new_n219), .A3(new_n220), .ZN(new_n221));
  INV_X1    g035(.A(new_n221), .ZN(new_n222));
  AOI21_X1  g036(.A(new_n220), .B1(new_n210), .B2(new_n219), .ZN(new_n223));
  OAI21_X1  g037(.A(new_n190), .B1(new_n222), .B2(new_n223), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n210), .A2(new_n219), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n225), .A2(KEYINPUT92), .ZN(new_n226));
  NAND3_X1  g040(.A1(new_n226), .A2(new_n189), .A3(new_n221), .ZN(new_n227));
  XNOR2_X1  g041(.A(KEYINPUT72), .B(G902), .ZN(new_n228));
  NAND3_X1  g042(.A1(new_n224), .A2(new_n227), .A3(new_n228), .ZN(new_n229));
  INV_X1    g043(.A(KEYINPUT93), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n229), .A2(new_n230), .ZN(new_n231));
  INV_X1    g045(.A(G478), .ZN(new_n232));
  NOR2_X1   g046(.A1(new_n232), .A2(KEYINPUT15), .ZN(new_n233));
  NAND4_X1  g047(.A1(new_n224), .A2(new_n227), .A3(KEYINPUT93), .A4(new_n228), .ZN(new_n234));
  NAND3_X1  g048(.A1(new_n231), .A2(new_n233), .A3(new_n234), .ZN(new_n235));
  INV_X1    g049(.A(G952), .ZN(new_n236));
  AOI211_X1 g050(.A(G953), .B(new_n236), .C1(G234), .C2(G237), .ZN(new_n237));
  XOR2_X1   g051(.A(KEYINPUT21), .B(G898), .Z(new_n238));
  XNOR2_X1  g052(.A(new_n238), .B(KEYINPUT94), .ZN(new_n239));
  INV_X1    g053(.A(new_n239), .ZN(new_n240));
  INV_X1    g054(.A(G953), .ZN(new_n241));
  AOI211_X1 g055(.A(new_n241), .B(new_n228), .C1(G234), .C2(G237), .ZN(new_n242));
  AOI21_X1  g056(.A(new_n237), .B1(new_n240), .B2(new_n242), .ZN(new_n243));
  INV_X1    g057(.A(new_n243), .ZN(new_n244));
  OR2_X1    g058(.A1(new_n229), .A2(new_n233), .ZN(new_n245));
  AND3_X1   g059(.A1(new_n235), .A2(new_n244), .A3(new_n245), .ZN(new_n246));
  INV_X1    g060(.A(KEYINPUT20), .ZN(new_n247));
  XNOR2_X1  g061(.A(G113), .B(G122), .ZN(new_n248));
  INV_X1    g062(.A(G104), .ZN(new_n249));
  XNOR2_X1  g063(.A(new_n248), .B(new_n249), .ZN(new_n250));
  INV_X1    g064(.A(G140), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n251), .A2(G125), .ZN(new_n252));
  INV_X1    g066(.A(G125), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n253), .A2(G140), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n252), .A2(new_n254), .ZN(new_n255));
  INV_X1    g069(.A(KEYINPUT76), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  NAND3_X1  g071(.A1(new_n252), .A2(new_n254), .A3(KEYINPUT76), .ZN(new_n258));
  AND2_X1   g072(.A1(KEYINPUT65), .A2(G146), .ZN(new_n259));
  NOR2_X1   g073(.A1(KEYINPUT65), .A2(G146), .ZN(new_n260));
  NOR2_X1   g074(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  NAND3_X1  g075(.A1(new_n257), .A2(new_n258), .A3(new_n261), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n255), .A2(G146), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n262), .A2(new_n263), .ZN(new_n264));
  NOR2_X1   g078(.A1(G237), .A2(G953), .ZN(new_n265));
  AND2_X1   g079(.A1(new_n192), .A2(KEYINPUT87), .ZN(new_n266));
  NOR2_X1   g080(.A1(new_n192), .A2(KEYINPUT87), .ZN(new_n267));
  OAI211_X1 g081(.A(G214), .B(new_n265), .C1(new_n266), .C2(new_n267), .ZN(new_n268));
  INV_X1    g082(.A(KEYINPUT18), .ZN(new_n269));
  INV_X1    g083(.A(G131), .ZN(new_n270));
  NOR2_X1   g084(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n265), .A2(G214), .ZN(new_n272));
  OAI21_X1  g086(.A(new_n272), .B1(KEYINPUT87), .B2(new_n192), .ZN(new_n273));
  NAND3_X1  g087(.A1(new_n268), .A2(new_n271), .A3(new_n273), .ZN(new_n274));
  INV_X1    g088(.A(new_n274), .ZN(new_n275));
  AOI21_X1  g089(.A(new_n271), .B1(new_n268), .B2(new_n273), .ZN(new_n276));
  OAI21_X1  g090(.A(new_n264), .B1(new_n275), .B2(new_n276), .ZN(new_n277));
  NAND3_X1  g091(.A1(new_n252), .A2(new_n254), .A3(KEYINPUT16), .ZN(new_n278));
  INV_X1    g092(.A(KEYINPUT16), .ZN(new_n279));
  NAND3_X1  g093(.A1(new_n279), .A2(new_n251), .A3(G125), .ZN(new_n280));
  INV_X1    g094(.A(KEYINPUT74), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  NAND4_X1  g096(.A1(new_n279), .A2(new_n251), .A3(KEYINPUT74), .A4(G125), .ZN(new_n283));
  NAND3_X1  g097(.A1(new_n278), .A2(new_n282), .A3(new_n283), .ZN(new_n284));
  INV_X1    g098(.A(G146), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  NAND4_X1  g100(.A1(new_n278), .A2(new_n282), .A3(G146), .A4(new_n283), .ZN(new_n287));
  NAND3_X1  g101(.A1(new_n286), .A2(KEYINPUT75), .A3(new_n287), .ZN(new_n288));
  INV_X1    g102(.A(KEYINPUT75), .ZN(new_n289));
  NAND3_X1  g103(.A1(new_n284), .A2(new_n289), .A3(new_n285), .ZN(new_n290));
  AND2_X1   g104(.A1(new_n288), .A2(new_n290), .ZN(new_n291));
  XNOR2_X1  g105(.A(KEYINPUT87), .B(G143), .ZN(new_n292));
  NOR2_X1   g106(.A1(new_n292), .A2(new_n272), .ZN(new_n293));
  AOI21_X1  g107(.A(new_n267), .B1(G214), .B2(new_n265), .ZN(new_n294));
  OAI21_X1  g108(.A(G131), .B1(new_n293), .B2(new_n294), .ZN(new_n295));
  NAND3_X1  g109(.A1(new_n268), .A2(new_n270), .A3(new_n273), .ZN(new_n296));
  INV_X1    g110(.A(KEYINPUT17), .ZN(new_n297));
  NAND3_X1  g111(.A1(new_n295), .A2(new_n296), .A3(new_n297), .ZN(new_n298));
  OAI211_X1 g112(.A(KEYINPUT17), .B(G131), .C1(new_n293), .C2(new_n294), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n298), .A2(new_n299), .ZN(new_n300));
  OAI211_X1 g114(.A(new_n250), .B(new_n277), .C1(new_n291), .C2(new_n300), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n295), .A2(new_n296), .ZN(new_n302));
  INV_X1    g116(.A(KEYINPUT19), .ZN(new_n303));
  NAND3_X1  g117(.A1(new_n257), .A2(new_n258), .A3(new_n303), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n255), .A2(KEYINPUT19), .ZN(new_n305));
  NAND3_X1  g119(.A1(new_n304), .A2(new_n261), .A3(new_n305), .ZN(new_n306));
  NAND3_X1  g120(.A1(new_n302), .A2(new_n306), .A3(new_n287), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n307), .A2(new_n277), .ZN(new_n308));
  INV_X1    g122(.A(new_n250), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n308), .A2(new_n309), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n301), .A2(new_n310), .ZN(new_n311));
  NOR2_X1   g125(.A1(G475), .A2(G902), .ZN(new_n312));
  AOI21_X1  g126(.A(new_n247), .B1(new_n311), .B2(new_n312), .ZN(new_n313));
  INV_X1    g127(.A(new_n312), .ZN(new_n314));
  AOI211_X1 g128(.A(KEYINPUT20), .B(new_n314), .C1(new_n301), .C2(new_n310), .ZN(new_n315));
  OAI21_X1  g129(.A(new_n277), .B1(new_n291), .B2(new_n300), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n316), .A2(new_n309), .ZN(new_n317));
  AOI21_X1  g131(.A(G902), .B1(new_n317), .B2(new_n301), .ZN(new_n318));
  XOR2_X1   g132(.A(KEYINPUT88), .B(G475), .Z(new_n319));
  OAI22_X1  g133(.A1(new_n313), .A2(new_n315), .B1(new_n318), .B2(new_n319), .ZN(new_n320));
  INV_X1    g134(.A(KEYINPUT89), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n320), .A2(new_n321), .ZN(new_n322));
  AOI21_X1  g136(.A(new_n250), .B1(new_n307), .B2(new_n277), .ZN(new_n323));
  INV_X1    g137(.A(new_n276), .ZN(new_n324));
  AOI22_X1  g138(.A1(new_n324), .A2(new_n274), .B1(new_n262), .B2(new_n263), .ZN(new_n325));
  AND2_X1   g139(.A1(new_n298), .A2(new_n299), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n288), .A2(new_n290), .ZN(new_n327));
  AOI21_X1  g141(.A(new_n325), .B1(new_n326), .B2(new_n327), .ZN(new_n328));
  AOI21_X1  g142(.A(new_n323), .B1(new_n328), .B2(new_n250), .ZN(new_n329));
  OAI21_X1  g143(.A(KEYINPUT20), .B1(new_n329), .B2(new_n314), .ZN(new_n330));
  NAND3_X1  g144(.A1(new_n311), .A2(new_n247), .A3(new_n312), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n330), .A2(new_n331), .ZN(new_n332));
  INV_X1    g146(.A(G902), .ZN(new_n333));
  NOR2_X1   g147(.A1(new_n328), .A2(new_n250), .ZN(new_n334));
  INV_X1    g148(.A(new_n301), .ZN(new_n335));
  OAI21_X1  g149(.A(new_n333), .B1(new_n334), .B2(new_n335), .ZN(new_n336));
  INV_X1    g150(.A(new_n319), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n336), .A2(new_n337), .ZN(new_n338));
  NAND3_X1  g152(.A1(new_n332), .A2(new_n338), .A3(KEYINPUT89), .ZN(new_n339));
  NAND3_X1  g153(.A1(new_n246), .A2(new_n322), .A3(new_n339), .ZN(new_n340));
  OAI21_X1  g154(.A(G210), .B1(G237), .B2(G902), .ZN(new_n341));
  INV_X1    g155(.A(new_n341), .ZN(new_n342));
  INV_X1    g156(.A(KEYINPUT1), .ZN(new_n343));
  INV_X1    g157(.A(KEYINPUT66), .ZN(new_n344));
  OAI21_X1  g158(.A(new_n344), .B1(new_n285), .B2(G143), .ZN(new_n345));
  AOI21_X1  g159(.A(new_n345), .B1(new_n261), .B2(G143), .ZN(new_n346));
  INV_X1    g160(.A(KEYINPUT65), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n347), .A2(new_n285), .ZN(new_n348));
  NAND2_X1  g162(.A1(KEYINPUT65), .A2(G146), .ZN(new_n349));
  NAND4_X1  g163(.A1(new_n348), .A2(KEYINPUT66), .A3(G143), .A4(new_n349), .ZN(new_n350));
  INV_X1    g164(.A(new_n350), .ZN(new_n351));
  OAI211_X1 g165(.A(new_n343), .B(G128), .C1(new_n346), .C2(new_n351), .ZN(new_n352));
  OAI21_X1  g166(.A(new_n192), .B1(new_n259), .B2(new_n260), .ZN(new_n353));
  INV_X1    g167(.A(KEYINPUT64), .ZN(new_n354));
  OAI21_X1  g168(.A(new_n354), .B1(new_n192), .B2(G146), .ZN(new_n355));
  NAND3_X1  g169(.A1(new_n285), .A2(KEYINPUT64), .A3(G143), .ZN(new_n356));
  NAND3_X1  g170(.A1(new_n353), .A2(new_n355), .A3(new_n356), .ZN(new_n357));
  AOI21_X1  g171(.A(new_n343), .B1(new_n261), .B2(G143), .ZN(new_n358));
  OAI21_X1  g172(.A(new_n357), .B1(new_n358), .B2(new_n197), .ZN(new_n359));
  NAND3_X1  g173(.A1(new_n352), .A2(new_n359), .A3(new_n253), .ZN(new_n360));
  NAND2_X1  g174(.A1(KEYINPUT0), .A2(G128), .ZN(new_n361));
  NAND3_X1  g175(.A1(new_n348), .A2(G143), .A3(new_n349), .ZN(new_n362));
  INV_X1    g176(.A(new_n345), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n362), .A2(new_n363), .ZN(new_n364));
  AOI21_X1  g178(.A(new_n361), .B1(new_n364), .B2(new_n350), .ZN(new_n365));
  INV_X1    g179(.A(new_n361), .ZN(new_n366));
  NOR2_X1   g180(.A1(KEYINPUT0), .A2(G128), .ZN(new_n367));
  OR2_X1    g181(.A1(new_n366), .A2(new_n367), .ZN(new_n368));
  AND2_X1   g182(.A1(new_n355), .A2(new_n356), .ZN(new_n369));
  AOI21_X1  g183(.A(new_n368), .B1(new_n369), .B2(new_n353), .ZN(new_n370));
  OAI21_X1  g184(.A(G125), .B1(new_n365), .B2(new_n370), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n360), .A2(new_n371), .ZN(new_n372));
  INV_X1    g186(.A(G224), .ZN(new_n373));
  NOR2_X1   g187(.A1(new_n373), .A2(G953), .ZN(new_n374));
  XOR2_X1   g188(.A(new_n372), .B(new_n374), .Z(new_n375));
  XNOR2_X1  g189(.A(KEYINPUT2), .B(G113), .ZN(new_n376));
  INV_X1    g190(.A(new_n376), .ZN(new_n377));
  INV_X1    g191(.A(KEYINPUT69), .ZN(new_n378));
  INV_X1    g192(.A(G119), .ZN(new_n379));
  OAI21_X1  g193(.A(new_n378), .B1(new_n379), .B2(G116), .ZN(new_n380));
  XNOR2_X1  g194(.A(KEYINPUT68), .B(G119), .ZN(new_n381));
  AOI21_X1  g195(.A(new_n380), .B1(new_n381), .B2(G116), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n379), .A2(KEYINPUT68), .ZN(new_n383));
  INV_X1    g197(.A(KEYINPUT68), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n384), .A2(G119), .ZN(new_n385));
  AND4_X1   g199(.A1(KEYINPUT69), .A2(new_n383), .A3(new_n385), .A4(G116), .ZN(new_n386));
  OAI21_X1  g200(.A(new_n377), .B1(new_n382), .B2(new_n386), .ZN(new_n387));
  NAND3_X1  g201(.A1(new_n383), .A2(new_n385), .A3(G116), .ZN(new_n388));
  INV_X1    g202(.A(new_n380), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n388), .A2(new_n389), .ZN(new_n390));
  NAND3_X1  g204(.A1(new_n381), .A2(KEYINPUT69), .A3(G116), .ZN(new_n391));
  NAND3_X1  g205(.A1(new_n390), .A2(new_n391), .A3(new_n376), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n387), .A2(new_n392), .ZN(new_n393));
  INV_X1    g207(.A(G101), .ZN(new_n394));
  OAI21_X1  g208(.A(KEYINPUT3), .B1(new_n249), .B2(G107), .ZN(new_n395));
  INV_X1    g209(.A(KEYINPUT3), .ZN(new_n396));
  NAND3_X1  g210(.A1(new_n396), .A2(new_n203), .A3(G104), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n249), .A2(G107), .ZN(new_n398));
  NAND3_X1  g212(.A1(new_n395), .A2(new_n397), .A3(new_n398), .ZN(new_n399));
  AOI21_X1  g213(.A(new_n394), .B1(new_n399), .B2(KEYINPUT79), .ZN(new_n400));
  INV_X1    g214(.A(KEYINPUT4), .ZN(new_n401));
  INV_X1    g215(.A(KEYINPUT79), .ZN(new_n402));
  NAND4_X1  g216(.A1(new_n395), .A2(new_n397), .A3(new_n402), .A4(new_n398), .ZN(new_n403));
  NAND3_X1  g217(.A1(new_n400), .A2(new_n401), .A3(new_n403), .ZN(new_n404));
  AND2_X1   g218(.A1(new_n400), .A2(new_n403), .ZN(new_n405));
  NAND4_X1  g219(.A1(new_n395), .A2(new_n397), .A3(new_n394), .A4(new_n398), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n406), .A2(KEYINPUT4), .ZN(new_n407));
  OAI211_X1 g221(.A(new_n393), .B(new_n404), .C1(new_n405), .C2(new_n407), .ZN(new_n408));
  AOI21_X1  g222(.A(new_n376), .B1(new_n390), .B2(new_n391), .ZN(new_n409));
  NOR2_X1   g223(.A1(new_n249), .A2(G107), .ZN(new_n410));
  NOR2_X1   g224(.A1(new_n203), .A2(G104), .ZN(new_n411));
  OAI21_X1  g225(.A(G101), .B1(new_n410), .B2(new_n411), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n406), .A2(new_n412), .ZN(new_n413));
  NOR2_X1   g227(.A1(new_n409), .A2(new_n413), .ZN(new_n414));
  INV_X1    g228(.A(KEYINPUT5), .ZN(new_n415));
  AOI21_X1  g229(.A(new_n415), .B1(new_n390), .B2(new_n391), .ZN(new_n416));
  NAND4_X1  g230(.A1(new_n383), .A2(new_n385), .A3(new_n415), .A4(G116), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n417), .A2(G113), .ZN(new_n418));
  OAI21_X1  g232(.A(new_n414), .B1(new_n416), .B2(new_n418), .ZN(new_n419));
  XNOR2_X1  g233(.A(G110), .B(G122), .ZN(new_n420));
  NAND3_X1  g234(.A1(new_n408), .A2(new_n419), .A3(new_n420), .ZN(new_n421));
  INV_X1    g235(.A(KEYINPUT6), .ZN(new_n422));
  NOR2_X1   g236(.A1(new_n422), .A2(KEYINPUT83), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n421), .A2(new_n423), .ZN(new_n424));
  AOI21_X1  g238(.A(new_n420), .B1(new_n408), .B2(new_n419), .ZN(new_n425));
  INV_X1    g239(.A(new_n425), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n424), .A2(new_n426), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n425), .A2(new_n423), .ZN(new_n428));
  AOI21_X1  g242(.A(new_n375), .B1(new_n427), .B2(new_n428), .ZN(new_n429));
  OAI21_X1  g243(.A(KEYINPUT7), .B1(new_n373), .B2(G953), .ZN(new_n430));
  INV_X1    g244(.A(new_n430), .ZN(new_n431));
  NAND3_X1  g245(.A1(new_n360), .A2(new_n371), .A3(new_n431), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n432), .A2(KEYINPUT86), .ZN(new_n433));
  INV_X1    g247(.A(KEYINPUT86), .ZN(new_n434));
  NAND4_X1  g248(.A1(new_n360), .A2(new_n371), .A3(new_n434), .A4(new_n431), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n372), .A2(new_n430), .ZN(new_n436));
  NAND4_X1  g250(.A1(new_n421), .A2(new_n433), .A3(new_n435), .A4(new_n436), .ZN(new_n437));
  XNOR2_X1  g251(.A(new_n420), .B(KEYINPUT8), .ZN(new_n438));
  INV_X1    g252(.A(new_n438), .ZN(new_n439));
  OAI21_X1  g253(.A(KEYINPUT5), .B1(new_n382), .B2(new_n386), .ZN(new_n440));
  INV_X1    g254(.A(KEYINPUT84), .ZN(new_n441));
  NAND3_X1  g255(.A1(new_n417), .A2(new_n441), .A3(G113), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n418), .A2(KEYINPUT84), .ZN(new_n443));
  NAND3_X1  g257(.A1(new_n440), .A2(new_n442), .A3(new_n443), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n444), .A2(new_n414), .ZN(new_n445));
  INV_X1    g259(.A(KEYINPUT85), .ZN(new_n446));
  OAI21_X1  g260(.A(new_n387), .B1(new_n416), .B2(new_n418), .ZN(new_n447));
  AOI22_X1  g261(.A1(new_n445), .A2(new_n446), .B1(new_n413), .B2(new_n447), .ZN(new_n448));
  NAND3_X1  g262(.A1(new_n444), .A2(new_n414), .A3(KEYINPUT85), .ZN(new_n449));
  AOI21_X1  g263(.A(new_n439), .B1(new_n448), .B2(new_n449), .ZN(new_n450));
  OAI21_X1  g264(.A(new_n333), .B1(new_n437), .B2(new_n450), .ZN(new_n451));
  OAI21_X1  g265(.A(new_n342), .B1(new_n429), .B2(new_n451), .ZN(new_n452));
  AND4_X1   g266(.A1(new_n421), .A2(new_n433), .A3(new_n435), .A4(new_n436), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n448), .A2(new_n449), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n454), .A2(new_n438), .ZN(new_n455));
  AOI21_X1  g269(.A(G902), .B1(new_n453), .B2(new_n455), .ZN(new_n456));
  XNOR2_X1  g270(.A(new_n372), .B(new_n374), .ZN(new_n457));
  AOI21_X1  g271(.A(new_n425), .B1(new_n423), .B2(new_n421), .ZN(new_n458));
  AND2_X1   g272(.A1(new_n425), .A2(new_n423), .ZN(new_n459));
  OAI21_X1  g273(.A(new_n457), .B1(new_n458), .B2(new_n459), .ZN(new_n460));
  NAND3_X1  g274(.A1(new_n456), .A2(new_n460), .A3(new_n341), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n452), .A2(new_n461), .ZN(new_n462));
  OAI21_X1  g276(.A(G214), .B1(G237), .B2(G902), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  NOR2_X1   g278(.A1(new_n340), .A2(new_n464), .ZN(new_n465));
  OAI21_X1  g279(.A(G221), .B1(new_n187), .B2(G902), .ZN(new_n466));
  INV_X1    g280(.A(new_n466), .ZN(new_n467));
  INV_X1    g281(.A(G469), .ZN(new_n468));
  NOR2_X1   g282(.A1(new_n468), .A2(new_n333), .ZN(new_n469));
  INV_X1    g283(.A(KEYINPUT10), .ZN(new_n470));
  INV_X1    g284(.A(new_n413), .ZN(new_n471));
  OAI21_X1  g285(.A(KEYINPUT1), .B1(new_n192), .B2(G146), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n472), .A2(G128), .ZN(new_n473));
  AND3_X1   g287(.A1(new_n364), .A2(new_n350), .A3(new_n473), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n343), .A2(G128), .ZN(new_n475));
  AOI21_X1  g289(.A(new_n475), .B1(new_n364), .B2(new_n350), .ZN(new_n476));
  OAI211_X1 g290(.A(new_n470), .B(new_n471), .C1(new_n474), .C2(new_n476), .ZN(new_n477));
  AOI21_X1  g291(.A(new_n413), .B1(new_n352), .B2(new_n359), .ZN(new_n478));
  OAI21_X1  g292(.A(new_n477), .B1(new_n478), .B2(new_n470), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n399), .A2(KEYINPUT79), .ZN(new_n480));
  AND4_X1   g294(.A1(new_n401), .A2(new_n480), .A3(G101), .A4(new_n403), .ZN(new_n481));
  AOI21_X1  g295(.A(new_n407), .B1(new_n400), .B2(new_n403), .ZN(new_n482));
  NOR2_X1   g296(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  NOR2_X1   g297(.A1(new_n365), .A2(new_n370), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  INV_X1    g299(.A(KEYINPUT11), .ZN(new_n486));
  OAI21_X1  g300(.A(new_n486), .B1(new_n201), .B2(G137), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n201), .A2(G137), .ZN(new_n488));
  INV_X1    g302(.A(G137), .ZN(new_n489));
  NAND3_X1  g303(.A1(new_n489), .A2(KEYINPUT11), .A3(G134), .ZN(new_n490));
  NAND3_X1  g304(.A1(new_n487), .A2(new_n488), .A3(new_n490), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n491), .A2(G131), .ZN(new_n492));
  NAND4_X1  g306(.A1(new_n487), .A2(new_n490), .A3(new_n270), .A4(new_n488), .ZN(new_n493));
  NAND3_X1  g307(.A1(new_n492), .A2(KEYINPUT67), .A3(new_n493), .ZN(new_n494));
  INV_X1    g308(.A(KEYINPUT80), .ZN(new_n495));
  INV_X1    g309(.A(KEYINPUT67), .ZN(new_n496));
  NAND3_X1  g310(.A1(new_n491), .A2(new_n496), .A3(G131), .ZN(new_n497));
  AND3_X1   g311(.A1(new_n494), .A2(new_n495), .A3(new_n497), .ZN(new_n498));
  AOI21_X1  g312(.A(new_n495), .B1(new_n494), .B2(new_n497), .ZN(new_n499));
  NOR2_X1   g313(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  NAND3_X1  g314(.A1(new_n479), .A2(new_n485), .A3(new_n500), .ZN(new_n501));
  INV_X1    g315(.A(KEYINPUT81), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n362), .A2(KEYINPUT1), .ZN(new_n504));
  AOI22_X1  g318(.A1(new_n504), .A2(G128), .B1(new_n369), .B2(new_n353), .ZN(new_n505));
  OAI21_X1  g319(.A(new_n471), .B1(new_n505), .B2(new_n476), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n506), .A2(KEYINPUT10), .ZN(new_n507));
  AOI22_X1  g321(.A1(new_n507), .A2(new_n477), .B1(new_n483), .B2(new_n484), .ZN(new_n508));
  NAND3_X1  g322(.A1(new_n508), .A2(KEYINPUT81), .A3(new_n500), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n503), .A2(new_n509), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n494), .A2(new_n497), .ZN(new_n511));
  INV_X1    g325(.A(new_n511), .ZN(new_n512));
  NOR3_X1   g326(.A1(new_n505), .A2(new_n476), .A3(new_n471), .ZN(new_n513));
  NAND3_X1  g327(.A1(new_n364), .A2(new_n350), .A3(new_n473), .ZN(new_n514));
  AOI21_X1  g328(.A(new_n413), .B1(new_n352), .B2(new_n514), .ZN(new_n515));
  OAI21_X1  g329(.A(new_n512), .B1(new_n513), .B2(new_n515), .ZN(new_n516));
  INV_X1    g330(.A(KEYINPUT12), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  OAI21_X1  g332(.A(new_n471), .B1(new_n474), .B2(new_n476), .ZN(new_n519));
  NAND3_X1  g333(.A1(new_n352), .A2(new_n359), .A3(new_n413), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  NAND3_X1  g335(.A1(new_n521), .A2(KEYINPUT12), .A3(new_n512), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n518), .A2(new_n522), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n510), .A2(new_n523), .ZN(new_n524));
  XNOR2_X1  g338(.A(G110), .B(G140), .ZN(new_n525));
  INV_X1    g339(.A(G227), .ZN(new_n526));
  NOR2_X1   g340(.A1(new_n526), .A2(G953), .ZN(new_n527));
  XNOR2_X1  g341(.A(new_n525), .B(new_n527), .ZN(new_n528));
  AOI21_X1  g342(.A(new_n528), .B1(new_n503), .B2(new_n509), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n479), .A2(new_n485), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n530), .A2(new_n512), .ZN(new_n531));
  AOI22_X1  g345(.A1(new_n524), .A2(new_n528), .B1(new_n529), .B2(new_n531), .ZN(new_n532));
  AOI21_X1  g346(.A(new_n469), .B1(new_n532), .B2(G469), .ZN(new_n533));
  AOI21_X1  g347(.A(KEYINPUT81), .B1(new_n508), .B2(new_n500), .ZN(new_n534));
  AND4_X1   g348(.A1(KEYINPUT81), .A2(new_n479), .A3(new_n485), .A4(new_n500), .ZN(new_n535));
  OAI21_X1  g349(.A(new_n531), .B1(new_n534), .B2(new_n535), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n536), .A2(new_n528), .ZN(new_n537));
  INV_X1    g351(.A(new_n528), .ZN(new_n538));
  INV_X1    g352(.A(KEYINPUT82), .ZN(new_n539));
  AOI21_X1  g353(.A(KEYINPUT12), .B1(new_n521), .B2(new_n512), .ZN(new_n540));
  AOI211_X1 g354(.A(new_n517), .B(new_n511), .C1(new_n519), .C2(new_n520), .ZN(new_n541));
  OAI21_X1  g355(.A(new_n539), .B1(new_n540), .B2(new_n541), .ZN(new_n542));
  NAND3_X1  g356(.A1(new_n518), .A2(KEYINPUT82), .A3(new_n522), .ZN(new_n543));
  NAND4_X1  g357(.A1(new_n510), .A2(new_n538), .A3(new_n542), .A4(new_n543), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n537), .A2(new_n544), .ZN(new_n545));
  NAND3_X1  g359(.A1(new_n545), .A2(new_n468), .A3(new_n228), .ZN(new_n546));
  AOI21_X1  g360(.A(new_n467), .B1(new_n533), .B2(new_n546), .ZN(new_n547));
  OAI21_X1  g361(.A(new_n366), .B1(new_n346), .B2(new_n351), .ZN(new_n548));
  INV_X1    g362(.A(new_n368), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n357), .A2(new_n549), .ZN(new_n550));
  NAND4_X1  g364(.A1(new_n548), .A2(new_n494), .A3(new_n550), .A4(new_n497), .ZN(new_n551));
  INV_X1    g365(.A(new_n488), .ZN(new_n552));
  NOR2_X1   g366(.A1(new_n201), .A2(G137), .ZN(new_n553));
  OAI21_X1  g367(.A(G131), .B1(new_n552), .B2(new_n553), .ZN(new_n554));
  AND2_X1   g368(.A1(new_n554), .A2(new_n493), .ZN(new_n555));
  OAI21_X1  g369(.A(new_n555), .B1(new_n505), .B2(new_n476), .ZN(new_n556));
  NOR3_X1   g370(.A1(new_n382), .A2(new_n386), .A3(new_n377), .ZN(new_n557));
  NOR2_X1   g371(.A1(new_n557), .A2(new_n409), .ZN(new_n558));
  AND3_X1   g372(.A1(new_n551), .A2(new_n556), .A3(new_n558), .ZN(new_n559));
  AOI21_X1  g373(.A(new_n558), .B1(new_n551), .B2(new_n556), .ZN(new_n560));
  OAI21_X1  g374(.A(KEYINPUT28), .B1(new_n559), .B2(new_n560), .ZN(new_n561));
  INV_X1    g375(.A(KEYINPUT71), .ZN(new_n562));
  OAI21_X1  g376(.A(new_n562), .B1(new_n559), .B2(KEYINPUT28), .ZN(new_n563));
  NAND3_X1  g377(.A1(new_n551), .A2(new_n556), .A3(new_n558), .ZN(new_n564));
  INV_X1    g378(.A(KEYINPUT28), .ZN(new_n565));
  NAND3_X1  g379(.A1(new_n564), .A2(KEYINPUT71), .A3(new_n565), .ZN(new_n566));
  NAND3_X1  g380(.A1(new_n561), .A2(new_n563), .A3(new_n566), .ZN(new_n567));
  XNOR2_X1  g381(.A(KEYINPUT26), .B(G101), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n265), .A2(G210), .ZN(new_n569));
  XNOR2_X1  g383(.A(new_n568), .B(new_n569), .ZN(new_n570));
  XNOR2_X1  g384(.A(KEYINPUT70), .B(KEYINPUT27), .ZN(new_n571));
  XNOR2_X1  g385(.A(new_n570), .B(new_n571), .ZN(new_n572));
  INV_X1    g386(.A(new_n572), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n567), .A2(new_n573), .ZN(new_n574));
  INV_X1    g388(.A(KEYINPUT30), .ZN(new_n575));
  AND3_X1   g389(.A1(new_n551), .A2(new_n556), .A3(new_n575), .ZN(new_n576));
  AOI21_X1  g390(.A(new_n575), .B1(new_n551), .B2(new_n556), .ZN(new_n577));
  OAI21_X1  g391(.A(new_n393), .B1(new_n576), .B2(new_n577), .ZN(new_n578));
  NAND3_X1  g392(.A1(new_n578), .A2(new_n564), .A3(new_n572), .ZN(new_n579));
  AOI21_X1  g393(.A(KEYINPUT29), .B1(new_n574), .B2(new_n579), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n573), .A2(KEYINPUT29), .ZN(new_n581));
  OAI21_X1  g395(.A(new_n228), .B1(new_n567), .B2(new_n581), .ZN(new_n582));
  OAI21_X1  g396(.A(G472), .B1(new_n580), .B2(new_n582), .ZN(new_n583));
  NOR2_X1   g397(.A1(G472), .A2(G902), .ZN(new_n584));
  INV_X1    g398(.A(new_n584), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n551), .A2(new_n556), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n586), .A2(KEYINPUT30), .ZN(new_n587));
  NAND3_X1  g401(.A1(new_n551), .A2(new_n556), .A3(new_n575), .ZN(new_n588));
  AOI21_X1  g402(.A(new_n558), .B1(new_n587), .B2(new_n588), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n564), .A2(new_n573), .ZN(new_n590));
  NOR3_X1   g404(.A1(new_n589), .A2(KEYINPUT31), .A3(new_n590), .ZN(new_n591));
  INV_X1    g405(.A(KEYINPUT31), .ZN(new_n592));
  INV_X1    g406(.A(new_n590), .ZN(new_n593));
  AOI21_X1  g407(.A(new_n592), .B1(new_n578), .B2(new_n593), .ZN(new_n594));
  NOR2_X1   g408(.A1(new_n591), .A2(new_n594), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n567), .A2(new_n572), .ZN(new_n596));
  AOI211_X1 g410(.A(KEYINPUT32), .B(new_n585), .C1(new_n595), .C2(new_n596), .ZN(new_n597));
  INV_X1    g411(.A(KEYINPUT32), .ZN(new_n598));
  OAI21_X1  g412(.A(KEYINPUT31), .B1(new_n589), .B2(new_n590), .ZN(new_n599));
  NAND3_X1  g413(.A1(new_n578), .A2(new_n593), .A3(new_n592), .ZN(new_n600));
  NAND3_X1  g414(.A1(new_n596), .A2(new_n599), .A3(new_n600), .ZN(new_n601));
  AOI21_X1  g415(.A(new_n598), .B1(new_n601), .B2(new_n584), .ZN(new_n602));
  OAI21_X1  g416(.A(new_n583), .B1(new_n597), .B2(new_n602), .ZN(new_n603));
  AOI21_X1  g417(.A(new_n188), .B1(new_n228), .B2(G234), .ZN(new_n604));
  NAND3_X1  g418(.A1(new_n383), .A2(new_n385), .A3(G128), .ZN(new_n605));
  NAND3_X1  g419(.A1(new_n197), .A2(KEYINPUT23), .A3(G119), .ZN(new_n606));
  AOI21_X1  g420(.A(G128), .B1(new_n383), .B2(new_n385), .ZN(new_n607));
  OAI211_X1 g421(.A(new_n605), .B(new_n606), .C1(new_n607), .C2(KEYINPUT23), .ZN(new_n608));
  INV_X1    g422(.A(KEYINPUT73), .ZN(new_n609));
  OAI21_X1  g423(.A(new_n609), .B1(new_n379), .B2(G128), .ZN(new_n610));
  NAND3_X1  g424(.A1(new_n197), .A2(KEYINPUT73), .A3(G119), .ZN(new_n611));
  AND3_X1   g425(.A1(new_n605), .A2(new_n610), .A3(new_n611), .ZN(new_n612));
  XOR2_X1   g426(.A(KEYINPUT24), .B(G110), .Z(new_n613));
  AOI22_X1  g427(.A1(G110), .A2(new_n608), .B1(new_n612), .B2(new_n613), .ZN(new_n614));
  NAND3_X1  g428(.A1(new_n614), .A2(new_n288), .A3(new_n290), .ZN(new_n615));
  OAI22_X1  g429(.A1(new_n608), .A2(G110), .B1(new_n612), .B2(new_n613), .ZN(new_n616));
  NAND3_X1  g430(.A1(new_n616), .A2(new_n287), .A3(new_n262), .ZN(new_n617));
  NAND3_X1  g431(.A1(new_n241), .A2(G221), .A3(G234), .ZN(new_n618));
  XNOR2_X1  g432(.A(new_n618), .B(KEYINPUT77), .ZN(new_n619));
  XNOR2_X1  g433(.A(KEYINPUT22), .B(G137), .ZN(new_n620));
  XNOR2_X1  g434(.A(new_n619), .B(new_n620), .ZN(new_n621));
  AND3_X1   g435(.A1(new_n615), .A2(new_n617), .A3(new_n621), .ZN(new_n622));
  AOI21_X1  g436(.A(new_n621), .B1(new_n615), .B2(new_n617), .ZN(new_n623));
  NOR2_X1   g437(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  AOI21_X1  g438(.A(KEYINPUT25), .B1(new_n624), .B2(new_n228), .ZN(new_n625));
  INV_X1    g439(.A(KEYINPUT25), .ZN(new_n626));
  INV_X1    g440(.A(new_n228), .ZN(new_n627));
  NOR4_X1   g441(.A1(new_n622), .A2(new_n623), .A3(new_n626), .A4(new_n627), .ZN(new_n628));
  OAI21_X1  g442(.A(new_n604), .B1(new_n625), .B2(new_n628), .ZN(new_n629));
  INV_X1    g443(.A(KEYINPUT78), .ZN(new_n630));
  NAND2_X1  g444(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  OAI211_X1 g445(.A(KEYINPUT78), .B(new_n604), .C1(new_n625), .C2(new_n628), .ZN(new_n632));
  NOR2_X1   g446(.A1(new_n604), .A2(G902), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n624), .A2(new_n633), .ZN(new_n634));
  NAND3_X1  g448(.A1(new_n631), .A2(new_n632), .A3(new_n634), .ZN(new_n635));
  INV_X1    g449(.A(new_n635), .ZN(new_n636));
  NAND4_X1  g450(.A1(new_n465), .A2(new_n547), .A3(new_n603), .A4(new_n636), .ZN(new_n637));
  XNOR2_X1  g451(.A(new_n637), .B(G101), .ZN(G3));
  INV_X1    g452(.A(new_n463), .ZN(new_n639));
  AOI21_X1  g453(.A(new_n639), .B1(new_n452), .B2(new_n461), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n640), .A2(new_n244), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n322), .A2(new_n339), .ZN(new_n642));
  AND3_X1   g456(.A1(new_n224), .A2(new_n227), .A3(KEYINPUT33), .ZN(new_n643));
  AOI21_X1  g457(.A(KEYINPUT33), .B1(new_n224), .B2(new_n227), .ZN(new_n644));
  OAI211_X1 g458(.A(G478), .B(new_n228), .C1(new_n643), .C2(new_n644), .ZN(new_n645));
  NAND3_X1  g459(.A1(new_n231), .A2(new_n232), .A3(new_n234), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  AOI21_X1  g461(.A(KEYINPUT95), .B1(new_n642), .B2(new_n647), .ZN(new_n648));
  INV_X1    g462(.A(new_n648), .ZN(new_n649));
  NAND3_X1  g463(.A1(new_n642), .A2(KEYINPUT95), .A3(new_n647), .ZN(new_n650));
  AOI21_X1  g464(.A(new_n641), .B1(new_n649), .B2(new_n650), .ZN(new_n651));
  NAND2_X1  g465(.A1(new_n586), .A2(new_n393), .ZN(new_n652));
  AOI21_X1  g466(.A(new_n565), .B1(new_n652), .B2(new_n564), .ZN(new_n653));
  AND3_X1   g467(.A1(new_n564), .A2(KEYINPUT71), .A3(new_n565), .ZN(new_n654));
  NOR2_X1   g468(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  AOI21_X1  g469(.A(new_n573), .B1(new_n655), .B2(new_n563), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n599), .A2(new_n600), .ZN(new_n657));
  OAI21_X1  g471(.A(new_n584), .B1(new_n656), .B2(new_n657), .ZN(new_n658));
  AOI21_X1  g472(.A(new_n627), .B1(new_n595), .B2(new_n596), .ZN(new_n659));
  INV_X1    g473(.A(G472), .ZN(new_n660));
  OAI21_X1  g474(.A(new_n658), .B1(new_n659), .B2(new_n660), .ZN(new_n661));
  NOR2_X1   g475(.A1(new_n661), .A2(new_n635), .ZN(new_n662));
  NAND3_X1  g476(.A1(new_n651), .A2(new_n547), .A3(new_n662), .ZN(new_n663));
  XOR2_X1   g477(.A(KEYINPUT34), .B(G104), .Z(new_n664));
  XNOR2_X1  g478(.A(new_n663), .B(new_n664), .ZN(G6));
  NAND2_X1  g479(.A1(new_n235), .A2(new_n245), .ZN(new_n666));
  NAND2_X1  g480(.A1(new_n313), .A2(KEYINPUT96), .ZN(new_n667));
  INV_X1    g481(.A(KEYINPUT96), .ZN(new_n668));
  NAND3_X1  g482(.A1(new_n330), .A2(new_n331), .A3(new_n668), .ZN(new_n669));
  NAND4_X1  g483(.A1(new_n666), .A2(new_n338), .A3(new_n667), .A4(new_n669), .ZN(new_n670));
  NOR2_X1   g484(.A1(new_n641), .A2(new_n670), .ZN(new_n671));
  NAND3_X1  g485(.A1(new_n671), .A2(new_n547), .A3(new_n662), .ZN(new_n672));
  XOR2_X1   g486(.A(KEYINPUT35), .B(G107), .Z(new_n673));
  XNOR2_X1  g487(.A(new_n672), .B(new_n673), .ZN(G9));
  INV_X1    g488(.A(new_n621), .ZN(new_n675));
  NOR2_X1   g489(.A1(new_n675), .A2(KEYINPUT36), .ZN(new_n676));
  XNOR2_X1  g490(.A(new_n676), .B(KEYINPUT97), .ZN(new_n677));
  NAND2_X1  g491(.A1(new_n615), .A2(new_n617), .ZN(new_n678));
  XNOR2_X1  g492(.A(new_n677), .B(new_n678), .ZN(new_n679));
  NAND2_X1  g493(.A1(new_n679), .A2(new_n633), .ZN(new_n680));
  AND3_X1   g494(.A1(new_n680), .A2(new_n631), .A3(new_n632), .ZN(new_n681));
  NOR2_X1   g495(.A1(new_n681), .A2(new_n661), .ZN(new_n682));
  NAND3_X1  g496(.A1(new_n682), .A2(new_n547), .A3(new_n465), .ZN(new_n683));
  XOR2_X1   g497(.A(KEYINPUT37), .B(G110), .Z(new_n684));
  XNOR2_X1  g498(.A(new_n683), .B(new_n684), .ZN(G12));
  AOI211_X1 g499(.A(G469), .B(new_n627), .C1(new_n537), .C2(new_n544), .ZN(new_n686));
  NAND3_X1  g500(.A1(new_n510), .A2(new_n531), .A3(new_n538), .ZN(new_n687));
  AOI22_X1  g501(.A1(new_n503), .A2(new_n509), .B1(new_n522), .B2(new_n518), .ZN(new_n688));
  OAI211_X1 g502(.A(new_n687), .B(G469), .C1(new_n538), .C2(new_n688), .ZN(new_n689));
  INV_X1    g503(.A(new_n469), .ZN(new_n690));
  NAND2_X1  g504(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  OAI211_X1 g505(.A(new_n466), .B(new_n640), .C1(new_n686), .C2(new_n691), .ZN(new_n692));
  INV_X1    g506(.A(new_n692), .ZN(new_n693));
  NAND2_X1  g507(.A1(new_n658), .A2(KEYINPUT32), .ZN(new_n694));
  NAND3_X1  g508(.A1(new_n601), .A2(new_n598), .A3(new_n584), .ZN(new_n695));
  NAND2_X1  g509(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  AOI21_X1  g510(.A(new_n681), .B1(new_n583), .B2(new_n696), .ZN(new_n697));
  INV_X1    g511(.A(new_n666), .ZN(new_n698));
  NAND2_X1  g512(.A1(new_n669), .A2(new_n667), .ZN(new_n699));
  INV_X1    g513(.A(G900), .ZN(new_n700));
  NAND2_X1  g514(.A1(new_n242), .A2(new_n700), .ZN(new_n701));
  INV_X1    g515(.A(new_n237), .ZN(new_n702));
  NAND2_X1  g516(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  NAND2_X1  g517(.A1(new_n338), .A2(new_n703), .ZN(new_n704));
  NOR3_X1   g518(.A1(new_n698), .A2(new_n699), .A3(new_n704), .ZN(new_n705));
  NAND3_X1  g519(.A1(new_n693), .A2(new_n697), .A3(new_n705), .ZN(new_n706));
  XOR2_X1   g520(.A(KEYINPUT98), .B(G128), .Z(new_n707));
  XNOR2_X1  g521(.A(new_n706), .B(new_n707), .ZN(G30));
  XNOR2_X1  g522(.A(new_n703), .B(KEYINPUT39), .ZN(new_n709));
  NAND2_X1  g523(.A1(new_n547), .A2(new_n709), .ZN(new_n710));
  INV_X1    g524(.A(KEYINPUT104), .ZN(new_n711));
  XNOR2_X1  g525(.A(new_n710), .B(new_n711), .ZN(new_n712));
  NAND2_X1  g526(.A1(new_n712), .A2(KEYINPUT40), .ZN(new_n713));
  XNOR2_X1  g527(.A(new_n710), .B(KEYINPUT104), .ZN(new_n714));
  INV_X1    g528(.A(KEYINPUT40), .ZN(new_n715));
  NAND2_X1  g529(.A1(new_n714), .A2(new_n715), .ZN(new_n716));
  XOR2_X1   g530(.A(KEYINPUT99), .B(KEYINPUT38), .Z(new_n717));
  XNOR2_X1  g531(.A(new_n462), .B(new_n717), .ZN(new_n718));
  NAND3_X1  g532(.A1(new_n680), .A2(new_n631), .A3(new_n632), .ZN(new_n719));
  NOR2_X1   g533(.A1(new_n719), .A2(new_n639), .ZN(new_n720));
  AND4_X1   g534(.A1(new_n642), .A2(new_n718), .A3(new_n666), .A4(new_n720), .ZN(new_n721));
  NAND3_X1  g535(.A1(new_n713), .A2(new_n716), .A3(new_n721), .ZN(new_n722));
  OAI21_X1  g536(.A(new_n572), .B1(new_n559), .B2(new_n560), .ZN(new_n723));
  OAI211_X1 g537(.A(KEYINPUT100), .B(new_n723), .C1(new_n589), .C2(new_n590), .ZN(new_n724));
  NAND2_X1  g538(.A1(new_n724), .A2(new_n333), .ZN(new_n725));
  NAND2_X1  g539(.A1(new_n578), .A2(new_n593), .ZN(new_n726));
  AOI21_X1  g540(.A(KEYINPUT100), .B1(new_n726), .B2(new_n723), .ZN(new_n727));
  OAI211_X1 g541(.A(KEYINPUT101), .B(G472), .C1(new_n725), .C2(new_n727), .ZN(new_n728));
  OAI21_X1  g542(.A(G472), .B1(new_n725), .B2(new_n727), .ZN(new_n729));
  INV_X1    g543(.A(KEYINPUT101), .ZN(new_n730));
  NAND2_X1  g544(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  OAI211_X1 g545(.A(new_n728), .B(new_n731), .C1(new_n597), .C2(new_n602), .ZN(new_n732));
  INV_X1    g546(.A(KEYINPUT102), .ZN(new_n733));
  NAND2_X1  g547(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  NAND4_X1  g548(.A1(new_n696), .A2(KEYINPUT102), .A3(new_n728), .A4(new_n731), .ZN(new_n735));
  NAND2_X1  g549(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  XNOR2_X1  g550(.A(new_n736), .B(KEYINPUT103), .ZN(new_n737));
  INV_X1    g551(.A(new_n737), .ZN(new_n738));
  OR2_X1    g552(.A1(new_n722), .A2(new_n738), .ZN(new_n739));
  XNOR2_X1  g553(.A(KEYINPUT105), .B(G143), .ZN(new_n740));
  XNOR2_X1  g554(.A(new_n739), .B(new_n740), .ZN(G45));
  INV_X1    g555(.A(new_n703), .ZN(new_n742));
  AOI221_X4 g556(.A(new_n742), .B1(new_n646), .B2(new_n645), .C1(new_n322), .C2(new_n339), .ZN(new_n743));
  NAND3_X1  g557(.A1(new_n693), .A2(new_n697), .A3(new_n743), .ZN(new_n744));
  XNOR2_X1  g558(.A(new_n744), .B(G146), .ZN(G48));
  AOI21_X1  g559(.A(new_n635), .B1(new_n696), .B2(new_n583), .ZN(new_n746));
  AND2_X1   g560(.A1(new_n542), .A2(new_n543), .ZN(new_n747));
  AOI22_X1  g561(.A1(new_n529), .A2(new_n747), .B1(new_n536), .B2(new_n528), .ZN(new_n748));
  OAI21_X1  g562(.A(G469), .B1(new_n748), .B2(new_n627), .ZN(new_n749));
  NAND3_X1  g563(.A1(new_n749), .A2(new_n466), .A3(new_n546), .ZN(new_n750));
  INV_X1    g564(.A(KEYINPUT106), .ZN(new_n751));
  NAND2_X1  g565(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  NAND4_X1  g566(.A1(new_n749), .A2(new_n546), .A3(KEYINPUT106), .A4(new_n466), .ZN(new_n753));
  NAND4_X1  g567(.A1(new_n651), .A2(new_n746), .A3(new_n752), .A4(new_n753), .ZN(new_n754));
  XNOR2_X1  g568(.A(KEYINPUT41), .B(G113), .ZN(new_n755));
  XNOR2_X1  g569(.A(new_n754), .B(new_n755), .ZN(G15));
  NAND4_X1  g570(.A1(new_n752), .A2(new_n746), .A3(new_n671), .A4(new_n753), .ZN(new_n757));
  XNOR2_X1  g571(.A(new_n757), .B(KEYINPUT107), .ZN(new_n758));
  XNOR2_X1  g572(.A(KEYINPUT108), .B(G116), .ZN(new_n759));
  XNOR2_X1  g573(.A(new_n758), .B(new_n759), .ZN(G18));
  NAND4_X1  g574(.A1(new_n697), .A2(new_n752), .A3(new_n465), .A4(new_n753), .ZN(new_n761));
  XNOR2_X1  g575(.A(KEYINPUT109), .B(G119), .ZN(new_n762));
  XNOR2_X1  g576(.A(new_n761), .B(new_n762), .ZN(G21));
  OAI21_X1  g577(.A(KEYINPUT110), .B1(new_n659), .B2(new_n660), .ZN(new_n764));
  OAI21_X1  g578(.A(new_n228), .B1(new_n656), .B2(new_n657), .ZN(new_n765));
  INV_X1    g579(.A(KEYINPUT110), .ZN(new_n766));
  NAND3_X1  g580(.A1(new_n765), .A2(new_n766), .A3(G472), .ZN(new_n767));
  NAND3_X1  g581(.A1(new_n764), .A2(new_n658), .A3(new_n767), .ZN(new_n768));
  INV_X1    g582(.A(KEYINPUT111), .ZN(new_n769));
  NAND2_X1  g583(.A1(new_n635), .A2(new_n769), .ZN(new_n770));
  NAND4_X1  g584(.A1(new_n631), .A2(KEYINPUT111), .A3(new_n632), .A4(new_n634), .ZN(new_n771));
  AOI21_X1  g585(.A(new_n768), .B1(new_n770), .B2(new_n771), .ZN(new_n772));
  NAND3_X1  g586(.A1(new_n642), .A2(new_n640), .A3(new_n666), .ZN(new_n773));
  NOR2_X1   g587(.A1(new_n773), .A2(new_n243), .ZN(new_n774));
  NAND4_X1  g588(.A1(new_n772), .A2(new_n752), .A3(new_n753), .A4(new_n774), .ZN(new_n775));
  XNOR2_X1  g589(.A(new_n775), .B(G122), .ZN(G24));
  NAND4_X1  g590(.A1(new_n764), .A2(new_n719), .A3(new_n658), .A4(new_n767), .ZN(new_n777));
  NAND3_X1  g591(.A1(new_n642), .A2(new_n647), .A3(new_n703), .ZN(new_n778));
  NOR2_X1   g592(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  NAND4_X1  g593(.A1(new_n779), .A2(new_n640), .A3(new_n752), .A4(new_n753), .ZN(new_n780));
  XOR2_X1   g594(.A(KEYINPUT112), .B(G125), .Z(new_n781));
  XNOR2_X1  g595(.A(new_n780), .B(new_n781), .ZN(G27));
  NAND2_X1  g596(.A1(new_n770), .A2(new_n771), .ZN(new_n783));
  NAND2_X1  g597(.A1(new_n783), .A2(new_n603), .ZN(new_n784));
  NOR2_X1   g598(.A1(new_n462), .A2(new_n639), .ZN(new_n785));
  NAND3_X1  g599(.A1(new_n547), .A2(new_n743), .A3(new_n785), .ZN(new_n786));
  OAI21_X1  g600(.A(KEYINPUT42), .B1(new_n784), .B2(new_n786), .ZN(new_n787));
  OAI21_X1  g601(.A(new_n466), .B1(new_n686), .B2(new_n691), .ZN(new_n788));
  INV_X1    g602(.A(new_n785), .ZN(new_n789));
  NOR2_X1   g603(.A1(new_n788), .A2(new_n789), .ZN(new_n790));
  NOR2_X1   g604(.A1(new_n778), .A2(KEYINPUT42), .ZN(new_n791));
  NAND3_X1  g605(.A1(new_n790), .A2(new_n746), .A3(new_n791), .ZN(new_n792));
  NAND2_X1  g606(.A1(new_n787), .A2(new_n792), .ZN(new_n793));
  XNOR2_X1  g607(.A(new_n793), .B(new_n270), .ZN(G33));
  NAND3_X1  g608(.A1(new_n790), .A2(new_n746), .A3(new_n705), .ZN(new_n795));
  XNOR2_X1  g609(.A(new_n795), .B(G134), .ZN(G36));
  NAND3_X1  g610(.A1(new_n322), .A2(new_n339), .A3(new_n647), .ZN(new_n797));
  OR2_X1    g611(.A1(new_n797), .A2(KEYINPUT43), .ZN(new_n798));
  NAND2_X1  g612(.A1(new_n797), .A2(KEYINPUT43), .ZN(new_n799));
  NAND4_X1  g613(.A1(new_n798), .A2(new_n661), .A3(new_n719), .A4(new_n799), .ZN(new_n800));
  INV_X1    g614(.A(KEYINPUT44), .ZN(new_n801));
  AOI21_X1  g615(.A(new_n789), .B1(new_n800), .B2(new_n801), .ZN(new_n802));
  OAI21_X1  g616(.A(new_n802), .B1(new_n801), .B2(new_n800), .ZN(new_n803));
  NAND2_X1  g617(.A1(new_n532), .A2(KEYINPUT45), .ZN(new_n804));
  INV_X1    g618(.A(KEYINPUT45), .ZN(new_n805));
  AND3_X1   g619(.A1(new_n510), .A2(new_n531), .A3(new_n538), .ZN(new_n806));
  AOI21_X1  g620(.A(new_n538), .B1(new_n510), .B2(new_n523), .ZN(new_n807));
  OAI21_X1  g621(.A(new_n805), .B1(new_n806), .B2(new_n807), .ZN(new_n808));
  NAND3_X1  g622(.A1(new_n804), .A2(G469), .A3(new_n808), .ZN(new_n809));
  NAND2_X1  g623(.A1(new_n809), .A2(new_n690), .ZN(new_n810));
  INV_X1    g624(.A(KEYINPUT46), .ZN(new_n811));
  AOI21_X1  g625(.A(new_n686), .B1(new_n810), .B2(new_n811), .ZN(new_n812));
  NAND3_X1  g626(.A1(new_n809), .A2(KEYINPUT46), .A3(new_n690), .ZN(new_n813));
  NAND2_X1  g627(.A1(new_n812), .A2(new_n813), .ZN(new_n814));
  NAND3_X1  g628(.A1(new_n814), .A2(new_n466), .A3(new_n709), .ZN(new_n815));
  OR2_X1    g629(.A1(new_n803), .A2(new_n815), .ZN(new_n816));
  XNOR2_X1  g630(.A(KEYINPUT113), .B(G137), .ZN(new_n817));
  XNOR2_X1  g631(.A(new_n816), .B(new_n817), .ZN(G39));
  AOI21_X1  g632(.A(KEYINPUT47), .B1(new_n814), .B2(new_n466), .ZN(new_n819));
  INV_X1    g633(.A(KEYINPUT47), .ZN(new_n820));
  AOI211_X1 g634(.A(new_n820), .B(new_n467), .C1(new_n812), .C2(new_n813), .ZN(new_n821));
  OR2_X1    g635(.A1(new_n819), .A2(new_n821), .ZN(new_n822));
  NOR4_X1   g636(.A1(new_n603), .A2(new_n789), .A3(new_n778), .A4(new_n636), .ZN(new_n823));
  NAND2_X1  g637(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  XNOR2_X1  g638(.A(new_n824), .B(G140), .ZN(G42));
  INV_X1    g639(.A(KEYINPUT115), .ZN(new_n826));
  INV_X1    g640(.A(KEYINPUT53), .ZN(new_n827));
  XOR2_X1   g641(.A(new_n703), .B(KEYINPUT114), .Z(new_n828));
  NAND4_X1  g642(.A1(new_n680), .A2(new_n631), .A3(new_n632), .A4(new_n828), .ZN(new_n829));
  NOR3_X1   g643(.A1(new_n788), .A2(new_n773), .A3(new_n829), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n736), .A2(new_n830), .ZN(new_n831));
  OAI211_X1 g645(.A(new_n693), .B(new_n697), .C1(new_n705), .C2(new_n743), .ZN(new_n832));
  NAND3_X1  g646(.A1(new_n780), .A2(new_n831), .A3(new_n832), .ZN(new_n833));
  INV_X1    g647(.A(KEYINPUT52), .ZN(new_n834));
  NAND2_X1  g648(.A1(new_n833), .A2(new_n834), .ZN(new_n835));
  NAND4_X1  g649(.A1(new_n780), .A2(new_n831), .A3(KEYINPUT52), .A4(new_n832), .ZN(new_n836));
  NAND2_X1  g650(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  INV_X1    g651(.A(new_n837), .ZN(new_n838));
  NOR3_X1   g652(.A1(new_n699), .A2(new_n666), .A3(new_n704), .ZN(new_n839));
  AND3_X1   g653(.A1(new_n603), .A2(new_n719), .A3(new_n839), .ZN(new_n840));
  OAI21_X1  g654(.A(new_n790), .B1(new_n779), .B2(new_n840), .ZN(new_n841));
  NAND4_X1  g655(.A1(new_n841), .A2(new_n787), .A3(new_n792), .A4(new_n795), .ZN(new_n842));
  INV_X1    g656(.A(new_n842), .ZN(new_n843));
  INV_X1    g657(.A(new_n768), .ZN(new_n844));
  NAND4_X1  g658(.A1(new_n844), .A2(new_n752), .A3(new_n753), .A4(new_n783), .ZN(new_n845));
  INV_X1    g659(.A(new_n774), .ZN(new_n846));
  NAND3_X1  g660(.A1(new_n752), .A2(new_n746), .A3(new_n753), .ZN(new_n847));
  INV_X1    g661(.A(new_n641), .ZN(new_n848));
  INV_X1    g662(.A(new_n650), .ZN(new_n849));
  OAI21_X1  g663(.A(new_n848), .B1(new_n849), .B2(new_n648), .ZN(new_n850));
  OAI22_X1  g664(.A1(new_n845), .A2(new_n846), .B1(new_n847), .B2(new_n850), .ZN(new_n851));
  NAND2_X1  g665(.A1(new_n642), .A2(new_n647), .ZN(new_n852));
  NAND3_X1  g666(.A1(new_n322), .A2(new_n339), .A3(new_n666), .ZN(new_n853));
  NAND2_X1  g667(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  NAND4_X1  g668(.A1(new_n854), .A2(new_n848), .A3(new_n662), .A4(new_n547), .ZN(new_n855));
  NAND4_X1  g669(.A1(new_n761), .A2(new_n637), .A3(new_n683), .A4(new_n855), .ZN(new_n856));
  NOR2_X1   g670(.A1(new_n851), .A2(new_n856), .ZN(new_n857));
  INV_X1    g671(.A(KEYINPUT107), .ZN(new_n858));
  XNOR2_X1  g672(.A(new_n757), .B(new_n858), .ZN(new_n859));
  NAND3_X1  g673(.A1(new_n843), .A2(new_n857), .A3(new_n859), .ZN(new_n860));
  OAI21_X1  g674(.A(new_n827), .B1(new_n838), .B2(new_n860), .ZN(new_n861));
  AND3_X1   g675(.A1(new_n855), .A2(new_n637), .A3(new_n683), .ZN(new_n862));
  NAND4_X1  g676(.A1(new_n862), .A2(new_n754), .A3(new_n775), .A4(new_n761), .ZN(new_n863));
  NOR3_X1   g677(.A1(new_n863), .A2(new_n758), .A3(new_n842), .ZN(new_n864));
  NAND3_X1  g678(.A1(new_n864), .A2(KEYINPUT53), .A3(new_n837), .ZN(new_n865));
  AND3_X1   g679(.A1(new_n861), .A2(KEYINPUT54), .A3(new_n865), .ZN(new_n866));
  AOI21_X1  g680(.A(KEYINPUT54), .B1(new_n861), .B2(new_n865), .ZN(new_n867));
  OAI21_X1  g681(.A(new_n826), .B1(new_n866), .B2(new_n867), .ZN(new_n868));
  INV_X1    g682(.A(KEYINPUT54), .ZN(new_n869));
  NOR2_X1   g683(.A1(new_n863), .A2(new_n758), .ZN(new_n870));
  AND4_X1   g684(.A1(KEYINPUT53), .A2(new_n870), .A3(new_n837), .A4(new_n843), .ZN(new_n871));
  AOI21_X1  g685(.A(KEYINPUT53), .B1(new_n864), .B2(new_n837), .ZN(new_n872));
  OAI21_X1  g686(.A(new_n869), .B1(new_n871), .B2(new_n872), .ZN(new_n873));
  NAND3_X1  g687(.A1(new_n861), .A2(KEYINPUT54), .A3(new_n865), .ZN(new_n874));
  NAND3_X1  g688(.A1(new_n873), .A2(KEYINPUT115), .A3(new_n874), .ZN(new_n875));
  AND2_X1   g689(.A1(new_n752), .A2(new_n753), .ZN(new_n876));
  NAND2_X1  g690(.A1(new_n876), .A2(new_n785), .ZN(new_n877));
  INV_X1    g691(.A(new_n877), .ZN(new_n878));
  INV_X1    g692(.A(new_n777), .ZN(new_n879));
  NAND3_X1  g693(.A1(new_n798), .A2(new_n237), .A3(new_n799), .ZN(new_n880));
  INV_X1    g694(.A(new_n880), .ZN(new_n881));
  NAND4_X1  g695(.A1(new_n878), .A2(KEYINPUT118), .A3(new_n879), .A4(new_n881), .ZN(new_n882));
  INV_X1    g696(.A(KEYINPUT118), .ZN(new_n883));
  NAND3_X1  g697(.A1(new_n876), .A2(new_n881), .A3(new_n785), .ZN(new_n884));
  OAI21_X1  g698(.A(new_n883), .B1(new_n884), .B2(new_n777), .ZN(new_n885));
  NAND2_X1  g699(.A1(new_n882), .A2(new_n885), .ZN(new_n886));
  NOR2_X1   g700(.A1(new_n635), .A2(new_n702), .ZN(new_n887));
  INV_X1    g701(.A(new_n887), .ZN(new_n888));
  NOR2_X1   g702(.A1(new_n877), .A2(new_n888), .ZN(new_n889));
  NOR2_X1   g703(.A1(new_n642), .A2(new_n647), .ZN(new_n890));
  NAND3_X1  g704(.A1(new_n738), .A2(new_n889), .A3(new_n890), .ZN(new_n891));
  NAND2_X1  g705(.A1(new_n886), .A2(new_n891), .ZN(new_n892));
  INV_X1    g706(.A(KEYINPUT116), .ZN(new_n893));
  NAND2_X1  g707(.A1(new_n772), .A2(new_n785), .ZN(new_n894));
  OAI21_X1  g708(.A(new_n893), .B1(new_n894), .B2(new_n880), .ZN(new_n895));
  NAND4_X1  g709(.A1(new_n881), .A2(new_n772), .A3(KEYINPUT116), .A4(new_n785), .ZN(new_n896));
  NAND2_X1  g710(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  NOR2_X1   g711(.A1(new_n819), .A2(new_n821), .ZN(new_n898));
  NAND2_X1  g712(.A1(new_n749), .A2(new_n546), .ZN(new_n899));
  NOR2_X1   g713(.A1(new_n899), .A2(new_n466), .ZN(new_n900));
  INV_X1    g714(.A(new_n900), .ZN(new_n901));
  AOI21_X1  g715(.A(new_n897), .B1(new_n898), .B2(new_n901), .ZN(new_n902));
  NOR2_X1   g716(.A1(new_n892), .A2(new_n902), .ZN(new_n903));
  NOR2_X1   g717(.A1(new_n845), .A2(new_n880), .ZN(new_n904));
  NOR2_X1   g718(.A1(new_n718), .A2(new_n463), .ZN(new_n905));
  NAND2_X1  g719(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  INV_X1    g720(.A(KEYINPUT50), .ZN(new_n907));
  NAND2_X1  g721(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  NAND3_X1  g722(.A1(new_n904), .A2(KEYINPUT50), .A3(new_n905), .ZN(new_n909));
  NAND2_X1  g723(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  INV_X1    g724(.A(KEYINPUT117), .ZN(new_n911));
  NAND2_X1  g725(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  NAND3_X1  g726(.A1(new_n908), .A2(KEYINPUT117), .A3(new_n909), .ZN(new_n913));
  NAND2_X1  g727(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  AOI21_X1  g728(.A(KEYINPUT51), .B1(new_n903), .B2(new_n914), .ZN(new_n915));
  NOR3_X1   g729(.A1(new_n737), .A2(new_n877), .A3(new_n888), .ZN(new_n916));
  AOI22_X1  g730(.A1(new_n916), .A2(new_n890), .B1(new_n882), .B2(new_n885), .ZN(new_n917));
  OAI211_X1 g731(.A(new_n895), .B(new_n896), .C1(new_n822), .C2(new_n900), .ZN(new_n918));
  INV_X1    g732(.A(KEYINPUT51), .ZN(new_n919));
  AOI21_X1  g733(.A(new_n919), .B1(new_n908), .B2(new_n909), .ZN(new_n920));
  NAND3_X1  g734(.A1(new_n917), .A2(new_n918), .A3(new_n920), .ZN(new_n921));
  NOR2_X1   g735(.A1(new_n849), .A2(new_n648), .ZN(new_n922));
  INV_X1    g736(.A(new_n922), .ZN(new_n923));
  NAND3_X1  g737(.A1(new_n738), .A2(new_n923), .A3(new_n889), .ZN(new_n924));
  NOR2_X1   g738(.A1(new_n884), .A2(new_n784), .ZN(new_n925));
  INV_X1    g739(.A(KEYINPUT48), .ZN(new_n926));
  NOR2_X1   g740(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  NOR3_X1   g741(.A1(new_n884), .A2(KEYINPUT48), .A3(new_n784), .ZN(new_n928));
  OAI21_X1  g742(.A(new_n924), .B1(new_n927), .B2(new_n928), .ZN(new_n929));
  NAND2_X1  g743(.A1(new_n904), .A2(new_n640), .ZN(new_n930));
  NAND2_X1  g744(.A1(new_n930), .A2(KEYINPUT119), .ZN(new_n931));
  INV_X1    g745(.A(KEYINPUT119), .ZN(new_n932));
  NAND3_X1  g746(.A1(new_n904), .A2(new_n932), .A3(new_n640), .ZN(new_n933));
  NAND4_X1  g747(.A1(new_n931), .A2(G952), .A3(new_n241), .A4(new_n933), .ZN(new_n934));
  NOR2_X1   g748(.A1(new_n929), .A2(new_n934), .ZN(new_n935));
  NAND2_X1  g749(.A1(new_n921), .A2(new_n935), .ZN(new_n936));
  NOR2_X1   g750(.A1(new_n915), .A2(new_n936), .ZN(new_n937));
  NAND3_X1  g751(.A1(new_n868), .A2(new_n875), .A3(new_n937), .ZN(new_n938));
  NAND2_X1  g752(.A1(new_n236), .A2(new_n241), .ZN(new_n939));
  XNOR2_X1  g753(.A(new_n939), .B(KEYINPUT120), .ZN(new_n940));
  NAND2_X1  g754(.A1(new_n938), .A2(new_n940), .ZN(new_n941));
  XOR2_X1   g755(.A(new_n899), .B(KEYINPUT49), .Z(new_n942));
  NOR4_X1   g756(.A1(new_n718), .A2(new_n467), .A3(new_n639), .A4(new_n797), .ZN(new_n943));
  NAND4_X1  g757(.A1(new_n738), .A2(new_n783), .A3(new_n942), .A4(new_n943), .ZN(new_n944));
  NAND2_X1  g758(.A1(new_n941), .A2(new_n944), .ZN(G75));
  AOI21_X1  g759(.A(new_n228), .B1(new_n861), .B2(new_n865), .ZN(new_n946));
  NAND2_X1  g760(.A1(new_n946), .A2(new_n342), .ZN(new_n947));
  INV_X1    g761(.A(KEYINPUT56), .ZN(new_n948));
  NAND2_X1  g762(.A1(new_n427), .A2(new_n428), .ZN(new_n949));
  XNOR2_X1  g763(.A(new_n949), .B(KEYINPUT121), .ZN(new_n950));
  XNOR2_X1  g764(.A(new_n950), .B(KEYINPUT55), .ZN(new_n951));
  XNOR2_X1  g765(.A(new_n951), .B(new_n457), .ZN(new_n952));
  AND3_X1   g766(.A1(new_n947), .A2(new_n948), .A3(new_n952), .ZN(new_n953));
  AOI21_X1  g767(.A(new_n952), .B1(new_n947), .B2(new_n948), .ZN(new_n954));
  NOR2_X1   g768(.A1(new_n241), .A2(G952), .ZN(new_n955));
  NOR3_X1   g769(.A1(new_n953), .A2(new_n954), .A3(new_n955), .ZN(G51));
  XNOR2_X1  g770(.A(new_n469), .B(KEYINPUT57), .ZN(new_n957));
  NAND3_X1  g771(.A1(new_n873), .A2(new_n874), .A3(new_n957), .ZN(new_n958));
  NAND2_X1  g772(.A1(new_n958), .A2(KEYINPUT122), .ZN(new_n959));
  INV_X1    g773(.A(KEYINPUT122), .ZN(new_n960));
  NAND4_X1  g774(.A1(new_n873), .A2(new_n960), .A3(new_n874), .A4(new_n957), .ZN(new_n961));
  XNOR2_X1  g775(.A(new_n748), .B(KEYINPUT123), .ZN(new_n962));
  NAND3_X1  g776(.A1(new_n959), .A2(new_n961), .A3(new_n962), .ZN(new_n963));
  INV_X1    g777(.A(new_n809), .ZN(new_n964));
  NAND2_X1  g778(.A1(new_n946), .A2(new_n964), .ZN(new_n965));
  AOI21_X1  g779(.A(new_n955), .B1(new_n963), .B2(new_n965), .ZN(G54));
  NAND3_X1  g780(.A1(new_n946), .A2(KEYINPUT58), .A3(G475), .ZN(new_n967));
  AND2_X1   g781(.A1(new_n967), .A2(new_n329), .ZN(new_n968));
  NOR2_X1   g782(.A1(new_n967), .A2(new_n329), .ZN(new_n969));
  NOR3_X1   g783(.A1(new_n968), .A2(new_n969), .A3(new_n955), .ZN(G60));
  NOR2_X1   g784(.A1(new_n643), .A2(new_n644), .ZN(new_n971));
  INV_X1    g785(.A(new_n971), .ZN(new_n972));
  NAND2_X1  g786(.A1(G478), .A2(G902), .ZN(new_n973));
  XNOR2_X1  g787(.A(new_n973), .B(KEYINPUT59), .ZN(new_n974));
  NAND4_X1  g788(.A1(new_n873), .A2(new_n972), .A3(new_n874), .A4(new_n974), .ZN(new_n975));
  INV_X1    g789(.A(new_n955), .ZN(new_n976));
  NAND2_X1  g790(.A1(new_n975), .A2(new_n976), .ZN(new_n977));
  INV_X1    g791(.A(new_n875), .ZN(new_n978));
  AOI21_X1  g792(.A(KEYINPUT115), .B1(new_n873), .B2(new_n874), .ZN(new_n979));
  OAI21_X1  g793(.A(new_n974), .B1(new_n978), .B2(new_n979), .ZN(new_n980));
  AOI21_X1  g794(.A(new_n977), .B1(new_n980), .B2(new_n971), .ZN(G63));
  NOR2_X1   g795(.A1(new_n871), .A2(new_n872), .ZN(new_n982));
  NAND2_X1  g796(.A1(G217), .A2(G902), .ZN(new_n983));
  XNOR2_X1  g797(.A(new_n983), .B(KEYINPUT60), .ZN(new_n984));
  OAI22_X1  g798(.A1(new_n982), .A2(new_n984), .B1(new_n622), .B2(new_n623), .ZN(new_n985));
  NAND2_X1  g799(.A1(new_n861), .A2(new_n865), .ZN(new_n986));
  INV_X1    g800(.A(new_n984), .ZN(new_n987));
  XNOR2_X1  g801(.A(new_n679), .B(KEYINPUT124), .ZN(new_n988));
  NAND3_X1  g802(.A1(new_n986), .A2(new_n987), .A3(new_n988), .ZN(new_n989));
  NAND3_X1  g803(.A1(new_n985), .A2(new_n976), .A3(new_n989), .ZN(new_n990));
  INV_X1    g804(.A(KEYINPUT61), .ZN(new_n991));
  NAND2_X1  g805(.A1(new_n990), .A2(new_n991), .ZN(new_n992));
  NAND4_X1  g806(.A1(new_n985), .A2(KEYINPUT61), .A3(new_n976), .A4(new_n989), .ZN(new_n993));
  NAND2_X1  g807(.A1(new_n992), .A2(new_n993), .ZN(G66));
  OAI21_X1  g808(.A(new_n241), .B1(new_n863), .B2(new_n758), .ZN(new_n995));
  INV_X1    g809(.A(KEYINPUT125), .ZN(new_n996));
  XNOR2_X1  g810(.A(new_n995), .B(new_n996), .ZN(new_n997));
  OAI21_X1  g811(.A(G953), .B1(new_n240), .B2(new_n373), .ZN(new_n998));
  NAND2_X1  g812(.A1(new_n997), .A2(new_n998), .ZN(new_n999));
  NAND2_X1  g813(.A1(new_n999), .A2(KEYINPUT126), .ZN(new_n1000));
  INV_X1    g814(.A(KEYINPUT126), .ZN(new_n1001));
  NAND3_X1  g815(.A1(new_n997), .A2(new_n1001), .A3(new_n998), .ZN(new_n1002));
  NAND2_X1  g816(.A1(new_n1000), .A2(new_n1002), .ZN(new_n1003));
  INV_X1    g817(.A(new_n950), .ZN(new_n1004));
  INV_X1    g818(.A(G898), .ZN(new_n1005));
  AOI21_X1  g819(.A(new_n1004), .B1(new_n1005), .B2(G953), .ZN(new_n1006));
  XNOR2_X1  g820(.A(new_n1003), .B(new_n1006), .ZN(G69));
  NOR2_X1   g821(.A1(new_n576), .A2(new_n577), .ZN(new_n1008));
  NAND2_X1  g822(.A1(new_n304), .A2(new_n305), .ZN(new_n1009));
  XOR2_X1   g823(.A(new_n1008), .B(new_n1009), .Z(new_n1010));
  NAND4_X1  g824(.A1(new_n714), .A2(new_n746), .A3(new_n785), .A4(new_n854), .ZN(new_n1011));
  NAND3_X1  g825(.A1(new_n824), .A2(new_n816), .A3(new_n1011), .ZN(new_n1012));
  AND2_X1   g826(.A1(new_n780), .A2(new_n832), .ZN(new_n1013));
  NAND3_X1  g827(.A1(new_n739), .A2(KEYINPUT62), .A3(new_n1013), .ZN(new_n1014));
  OAI21_X1  g828(.A(new_n1013), .B1(new_n722), .B2(new_n738), .ZN(new_n1015));
  INV_X1    g829(.A(KEYINPUT62), .ZN(new_n1016));
  NAND2_X1  g830(.A1(new_n1015), .A2(new_n1016), .ZN(new_n1017));
  AOI21_X1  g831(.A(new_n1012), .B1(new_n1014), .B2(new_n1017), .ZN(new_n1018));
  OAI21_X1  g832(.A(new_n1010), .B1(new_n1018), .B2(G953), .ZN(new_n1019));
  INV_X1    g833(.A(new_n824), .ZN(new_n1020));
  OR3_X1    g834(.A1(new_n815), .A2(new_n773), .A3(new_n784), .ZN(new_n1021));
  NAND4_X1  g835(.A1(new_n1021), .A2(new_n787), .A3(new_n792), .A4(new_n795), .ZN(new_n1022));
  NAND2_X1  g836(.A1(new_n816), .A2(new_n1013), .ZN(new_n1023));
  NOR3_X1   g837(.A1(new_n1020), .A2(new_n1022), .A3(new_n1023), .ZN(new_n1024));
  NAND2_X1  g838(.A1(new_n1024), .A2(new_n241), .ZN(new_n1025));
  AOI21_X1  g839(.A(new_n1010), .B1(G900), .B2(G953), .ZN(new_n1026));
  NAND2_X1  g840(.A1(new_n1025), .A2(new_n1026), .ZN(new_n1027));
  OAI21_X1  g841(.A(G953), .B1(new_n526), .B2(new_n700), .ZN(new_n1028));
  XNOR2_X1  g842(.A(new_n1028), .B(KEYINPUT127), .ZN(new_n1029));
  AND3_X1   g843(.A1(new_n1019), .A2(new_n1027), .A3(new_n1029), .ZN(new_n1030));
  AOI21_X1  g844(.A(new_n1029), .B1(new_n1019), .B2(new_n1027), .ZN(new_n1031));
  NOR2_X1   g845(.A1(new_n1030), .A2(new_n1031), .ZN(G72));
  OAI21_X1  g846(.A(new_n573), .B1(new_n589), .B2(new_n559), .ZN(new_n1033));
  NAND2_X1  g847(.A1(new_n1018), .A2(new_n870), .ZN(new_n1034));
  NAND2_X1  g848(.A1(G472), .A2(G902), .ZN(new_n1035));
  XOR2_X1   g849(.A(new_n1035), .B(KEYINPUT63), .Z(new_n1036));
  AOI21_X1  g850(.A(new_n1033), .B1(new_n1034), .B2(new_n1036), .ZN(new_n1037));
  INV_X1    g851(.A(new_n1036), .ZN(new_n1038));
  AOI21_X1  g852(.A(new_n1038), .B1(new_n1024), .B2(new_n870), .ZN(new_n1039));
  OAI21_X1  g853(.A(new_n976), .B1(new_n1039), .B2(new_n579), .ZN(new_n1040));
  AND4_X1   g854(.A1(new_n579), .A2(new_n986), .A3(new_n1033), .A4(new_n1036), .ZN(new_n1041));
  NOR3_X1   g855(.A1(new_n1037), .A2(new_n1040), .A3(new_n1041), .ZN(G57));
endmodule


