//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 1 1 1 0 0 1 1 1 1 0 1 0 1 1 1 0 0 0 0 0 0 1 1 1 0 1 1 0 0 1 1 0 0 1 0 1 0 0 0 1 1 0 1 1 0 0 1 1 1 0 0 0 1 1 1 1 1 1 0 1 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:38:58 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n205, new_n206, new_n207, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n244, new_n245,
    new_n246, new_n248, new_n249, new_n250, new_n251, new_n252, new_n253,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1249, new_n1250, new_n1251, new_n1252, new_n1253, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1313, new_n1314;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  INV_X1    g0004(.A(G97), .ZN(new_n205));
  INV_X1    g0005(.A(G107), .ZN(new_n206));
  NAND2_X1  g0006(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  NAND2_X1  g0007(.A1(new_n207), .A2(G87), .ZN(G355));
  INV_X1    g0008(.A(G1), .ZN(new_n209));
  INV_X1    g0009(.A(G20), .ZN(new_n210));
  NOR2_X1   g0010(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  INV_X1    g0011(.A(new_n211), .ZN(new_n212));
  NOR2_X1   g0012(.A1(new_n212), .A2(G13), .ZN(new_n213));
  OAI211_X1 g0013(.A(new_n213), .B(G250), .C1(G257), .C2(G264), .ZN(new_n214));
  XOR2_X1   g0014(.A(new_n214), .B(KEYINPUT64), .Z(new_n215));
  XNOR2_X1  g0015(.A(new_n215), .B(KEYINPUT0), .ZN(new_n216));
  NAND2_X1  g0016(.A1(G1), .A2(G13), .ZN(new_n217));
  NOR2_X1   g0017(.A1(new_n217), .A2(new_n210), .ZN(new_n218));
  NOR3_X1   g0018(.A1(KEYINPUT65), .A2(G58), .A3(G68), .ZN(new_n219));
  INV_X1    g0019(.A(new_n219), .ZN(new_n220));
  OAI21_X1  g0020(.A(KEYINPUT65), .B1(G58), .B2(G68), .ZN(new_n221));
  AOI21_X1  g0021(.A(new_n202), .B1(new_n220), .B2(new_n221), .ZN(new_n222));
  AOI21_X1  g0022(.A(new_n216), .B1(new_n218), .B2(new_n222), .ZN(new_n223));
  AOI22_X1  g0023(.A1(G68), .A2(G238), .B1(G116), .B2(G270), .ZN(new_n224));
  INV_X1    g0024(.A(G226), .ZN(new_n225));
  INV_X1    g0025(.A(G77), .ZN(new_n226));
  INV_X1    g0026(.A(G244), .ZN(new_n227));
  OAI221_X1 g0027(.A(new_n224), .B1(new_n202), .B2(new_n225), .C1(new_n226), .C2(new_n227), .ZN(new_n228));
  NAND2_X1  g0028(.A1(new_n228), .A2(KEYINPUT66), .ZN(new_n229));
  AOI22_X1  g0029(.A1(G87), .A2(G250), .B1(G107), .B2(G264), .ZN(new_n230));
  AOI22_X1  g0030(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n231));
  NAND3_X1  g0031(.A1(new_n229), .A2(new_n230), .A3(new_n231), .ZN(new_n232));
  NOR2_X1   g0032(.A1(new_n228), .A2(KEYINPUT66), .ZN(new_n233));
  OAI21_X1  g0033(.A(new_n212), .B1(new_n232), .B2(new_n233), .ZN(new_n234));
  OAI21_X1  g0034(.A(new_n223), .B1(KEYINPUT1), .B2(new_n234), .ZN(new_n235));
  AOI21_X1  g0035(.A(new_n235), .B1(KEYINPUT1), .B2(new_n234), .ZN(G361));
  XNOR2_X1  g0036(.A(G238), .B(G244), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n237), .B(KEYINPUT2), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n238), .B(G226), .ZN(new_n239));
  INV_X1    g0039(.A(G232), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n241), .B(KEYINPUT67), .ZN(new_n242));
  XOR2_X1   g0042(.A(G250), .B(G257), .Z(new_n243));
  XNOR2_X1  g0043(.A(G264), .B(G270), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  INV_X1    g0045(.A(new_n245), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n242), .B(new_n246), .ZN(G358));
  XOR2_X1   g0047(.A(G68), .B(G77), .Z(new_n248));
  XNOR2_X1  g0048(.A(G50), .B(G58), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n248), .B(new_n249), .ZN(new_n250));
  XOR2_X1   g0050(.A(G87), .B(G97), .Z(new_n251));
  XNOR2_X1  g0051(.A(G107), .B(G116), .ZN(new_n252));
  XNOR2_X1  g0052(.A(new_n251), .B(new_n252), .ZN(new_n253));
  XNOR2_X1  g0053(.A(new_n250), .B(new_n253), .ZN(G351));
  AND2_X1   g0054(.A1(KEYINPUT3), .A2(G33), .ZN(new_n255));
  NOR2_X1   g0055(.A1(KEYINPUT3), .A2(G33), .ZN(new_n256));
  NOR2_X1   g0056(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n257), .A2(G77), .ZN(new_n258));
  INV_X1    g0058(.A(KEYINPUT68), .ZN(new_n259));
  INV_X1    g0059(.A(G1698), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  NAND2_X1  g0061(.A1(KEYINPUT68), .A2(G1698), .ZN(new_n262));
  OAI211_X1 g0062(.A(new_n261), .B(new_n262), .C1(new_n255), .C2(new_n256), .ZN(new_n263));
  INV_X1    g0063(.A(G222), .ZN(new_n264));
  OR2_X1    g0064(.A1(KEYINPUT3), .A2(G33), .ZN(new_n265));
  NAND2_X1  g0065(.A1(KEYINPUT3), .A2(G33), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n265), .A2(new_n266), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n267), .A2(G1698), .ZN(new_n268));
  INV_X1    g0068(.A(G223), .ZN(new_n269));
  OAI221_X1 g0069(.A(new_n258), .B1(new_n263), .B2(new_n264), .C1(new_n268), .C2(new_n269), .ZN(new_n270));
  AOI21_X1  g0070(.A(new_n217), .B1(G33), .B2(G41), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  OAI211_X1 g0072(.A(new_n209), .B(G274), .C1(G41), .C2(G45), .ZN(new_n273));
  INV_X1    g0073(.A(new_n273), .ZN(new_n274));
  OR2_X1    g0074(.A1(G41), .A2(G45), .ZN(new_n275));
  AND2_X1   g0075(.A1(G1), .A2(G13), .ZN(new_n276));
  NAND2_X1  g0076(.A1(G33), .A2(G41), .ZN(new_n277));
  AOI22_X1  g0077(.A1(new_n275), .A2(new_n209), .B1(new_n276), .B2(new_n277), .ZN(new_n278));
  AOI21_X1  g0078(.A(new_n274), .B1(new_n278), .B2(G226), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n272), .A2(new_n279), .ZN(new_n280));
  INV_X1    g0080(.A(G200), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  OAI21_X1  g0082(.A(new_n282), .B1(G190), .B2(new_n280), .ZN(new_n283));
  AOI21_X1  g0083(.A(KEYINPUT10), .B1(new_n283), .B2(KEYINPUT69), .ZN(new_n284));
  NOR2_X1   g0084(.A1(G20), .A2(G33), .ZN(new_n285));
  AOI22_X1  g0085(.A1(new_n203), .A2(G20), .B1(G150), .B2(new_n285), .ZN(new_n286));
  XNOR2_X1  g0086(.A(KEYINPUT8), .B(G58), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n210), .A2(G33), .ZN(new_n288));
  OAI21_X1  g0088(.A(new_n286), .B1(new_n287), .B2(new_n288), .ZN(new_n289));
  NAND3_X1  g0089(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n290), .A2(new_n217), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n289), .A2(new_n291), .ZN(new_n292));
  INV_X1    g0092(.A(G13), .ZN(new_n293));
  NOR3_X1   g0093(.A1(new_n293), .A2(new_n210), .A3(G1), .ZN(new_n294));
  INV_X1    g0094(.A(new_n294), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n295), .A2(new_n202), .ZN(new_n296));
  AOI21_X1  g0096(.A(new_n291), .B1(new_n209), .B2(G20), .ZN(new_n297));
  OAI21_X1  g0097(.A(new_n296), .B1(new_n297), .B2(new_n202), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n292), .A2(new_n298), .ZN(new_n299));
  XNOR2_X1  g0099(.A(new_n299), .B(KEYINPUT9), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n283), .A2(new_n300), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n284), .A2(new_n301), .ZN(new_n302));
  OAI211_X1 g0102(.A(new_n283), .B(new_n300), .C1(KEYINPUT69), .C2(KEYINPUT10), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n280), .A2(G169), .ZN(new_n304));
  INV_X1    g0104(.A(G179), .ZN(new_n305));
  OAI21_X1  g0105(.A(new_n304), .B1(new_n305), .B2(new_n280), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n306), .A2(new_n299), .ZN(new_n307));
  NAND2_X1  g0107(.A1(G20), .A2(G77), .ZN(new_n308));
  INV_X1    g0108(.A(new_n285), .ZN(new_n309));
  XNOR2_X1  g0109(.A(KEYINPUT15), .B(G87), .ZN(new_n310));
  OAI221_X1 g0110(.A(new_n308), .B1(new_n287), .B2(new_n309), .C1(new_n288), .C2(new_n310), .ZN(new_n311));
  AND2_X1   g0111(.A1(new_n311), .A2(new_n291), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n297), .A2(G77), .ZN(new_n313));
  OAI21_X1  g0113(.A(new_n313), .B1(G77), .B2(new_n295), .ZN(new_n314));
  NOR2_X1   g0114(.A1(new_n312), .A2(new_n314), .ZN(new_n315));
  INV_X1    g0115(.A(new_n278), .ZN(new_n316));
  OAI21_X1  g0116(.A(new_n273), .B1(new_n316), .B2(new_n227), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n257), .A2(G107), .ZN(new_n318));
  INV_X1    g0118(.A(G238), .ZN(new_n319));
  OAI221_X1 g0119(.A(new_n318), .B1(new_n263), .B2(new_n240), .C1(new_n268), .C2(new_n319), .ZN(new_n320));
  AOI21_X1  g0120(.A(new_n317), .B1(new_n320), .B2(new_n271), .ZN(new_n321));
  INV_X1    g0121(.A(G190), .ZN(new_n322));
  AND2_X1   g0122(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  NOR2_X1   g0123(.A1(new_n321), .A2(G200), .ZN(new_n324));
  OAI21_X1  g0124(.A(new_n315), .B1(new_n323), .B2(new_n324), .ZN(new_n325));
  INV_X1    g0125(.A(new_n315), .ZN(new_n326));
  AND2_X1   g0126(.A1(new_n321), .A2(G179), .ZN(new_n327));
  INV_X1    g0127(.A(G169), .ZN(new_n328));
  NOR2_X1   g0128(.A1(new_n321), .A2(new_n328), .ZN(new_n329));
  OAI21_X1  g0129(.A(new_n326), .B1(new_n327), .B2(new_n329), .ZN(new_n330));
  AND2_X1   g0130(.A1(new_n325), .A2(new_n330), .ZN(new_n331));
  NAND4_X1  g0131(.A1(new_n302), .A2(new_n303), .A3(new_n307), .A4(new_n331), .ZN(new_n332));
  OAI22_X1  g0132(.A1(new_n288), .A2(new_n226), .B1(new_n210), .B2(G68), .ZN(new_n333));
  OAI22_X1  g0133(.A1(new_n333), .A2(KEYINPUT71), .B1(new_n202), .B2(new_n309), .ZN(new_n334));
  AND2_X1   g0134(.A1(new_n333), .A2(KEYINPUT71), .ZN(new_n335));
  OAI21_X1  g0135(.A(new_n291), .B1(new_n334), .B2(new_n335), .ZN(new_n336));
  XOR2_X1   g0136(.A(KEYINPUT72), .B(KEYINPUT11), .Z(new_n337));
  OR2_X1    g0137(.A1(new_n336), .A2(new_n337), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n336), .A2(new_n337), .ZN(new_n339));
  NOR2_X1   g0139(.A1(new_n293), .A2(G1), .ZN(new_n340));
  INV_X1    g0140(.A(G68), .ZN(new_n341));
  NAND3_X1  g0141(.A1(new_n340), .A2(G20), .A3(new_n341), .ZN(new_n342));
  XOR2_X1   g0142(.A(new_n342), .B(KEYINPUT12), .Z(new_n343));
  AOI21_X1  g0143(.A(new_n343), .B1(G68), .B2(new_n297), .ZN(new_n344));
  NAND3_X1  g0144(.A1(new_n338), .A2(new_n339), .A3(new_n344), .ZN(new_n345));
  INV_X1    g0145(.A(new_n345), .ZN(new_n346));
  NAND3_X1  g0146(.A1(new_n277), .A2(G1), .A3(G13), .ZN(new_n347));
  OAI21_X1  g0147(.A(new_n209), .B1(G41), .B2(G45), .ZN(new_n348));
  NAND3_X1  g0148(.A1(new_n347), .A2(G238), .A3(new_n348), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n273), .A2(KEYINPUT70), .ZN(new_n350));
  INV_X1    g0150(.A(KEYINPUT70), .ZN(new_n351));
  NAND4_X1  g0151(.A1(new_n275), .A2(new_n351), .A3(new_n209), .A4(G274), .ZN(new_n352));
  NAND3_X1  g0152(.A1(new_n349), .A2(new_n350), .A3(new_n352), .ZN(new_n353));
  OAI211_X1 g0153(.A(G232), .B(G1698), .C1(new_n255), .C2(new_n256), .ZN(new_n354));
  NAND2_X1  g0154(.A1(G33), .A2(G97), .ZN(new_n355));
  OAI21_X1  g0155(.A(G226), .B1(new_n255), .B2(new_n256), .ZN(new_n356));
  XNOR2_X1  g0156(.A(KEYINPUT68), .B(G1698), .ZN(new_n357));
  OAI211_X1 g0157(.A(new_n354), .B(new_n355), .C1(new_n356), .C2(new_n357), .ZN(new_n358));
  AOI211_X1 g0158(.A(KEYINPUT13), .B(new_n353), .C1(new_n271), .C2(new_n358), .ZN(new_n359));
  INV_X1    g0159(.A(KEYINPUT13), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n358), .A2(new_n271), .ZN(new_n361));
  INV_X1    g0161(.A(new_n353), .ZN(new_n362));
  AOI21_X1  g0162(.A(new_n360), .B1(new_n361), .B2(new_n362), .ZN(new_n363));
  OAI21_X1  g0163(.A(G169), .B1(new_n359), .B2(new_n363), .ZN(new_n364));
  INV_X1    g0164(.A(KEYINPUT14), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  OAI211_X1 g0166(.A(KEYINPUT14), .B(G169), .C1(new_n359), .C2(new_n363), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n366), .A2(new_n367), .ZN(new_n368));
  INV_X1    g0168(.A(new_n355), .ZN(new_n369));
  AOI21_X1  g0169(.A(new_n225), .B1(new_n265), .B2(new_n266), .ZN(new_n370));
  AND2_X1   g0170(.A1(KEYINPUT68), .A2(G1698), .ZN(new_n371));
  NOR2_X1   g0171(.A1(KEYINPUT68), .A2(G1698), .ZN(new_n372));
  NOR2_X1   g0172(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  AOI21_X1  g0173(.A(new_n369), .B1(new_n370), .B2(new_n373), .ZN(new_n374));
  AOI21_X1  g0174(.A(new_n347), .B1(new_n374), .B2(new_n354), .ZN(new_n375));
  OAI21_X1  g0175(.A(KEYINPUT13), .B1(new_n375), .B2(new_n353), .ZN(new_n376));
  NAND3_X1  g0176(.A1(new_n361), .A2(new_n360), .A3(new_n362), .ZN(new_n377));
  NAND3_X1  g0177(.A1(new_n376), .A2(new_n377), .A3(G179), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n378), .A2(KEYINPUT73), .ZN(new_n379));
  INV_X1    g0179(.A(KEYINPUT73), .ZN(new_n380));
  NAND4_X1  g0180(.A1(new_n376), .A2(new_n377), .A3(new_n380), .A4(G179), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n379), .A2(new_n381), .ZN(new_n382));
  AOI21_X1  g0182(.A(new_n346), .B1(new_n368), .B2(new_n382), .ZN(new_n383));
  AOI21_X1  g0183(.A(G200), .B1(new_n376), .B2(new_n377), .ZN(new_n384));
  NOR3_X1   g0184(.A1(new_n359), .A2(new_n363), .A3(G190), .ZN(new_n385));
  OAI21_X1  g0185(.A(new_n346), .B1(new_n384), .B2(new_n385), .ZN(new_n386));
  INV_X1    g0186(.A(new_n386), .ZN(new_n387));
  NOR3_X1   g0187(.A1(new_n332), .A2(new_n383), .A3(new_n387), .ZN(new_n388));
  NAND4_X1  g0188(.A1(new_n265), .A2(KEYINPUT7), .A3(new_n210), .A4(new_n266), .ZN(new_n389));
  INV_X1    g0189(.A(KEYINPUT74), .ZN(new_n390));
  NOR2_X1   g0190(.A1(new_n389), .A2(new_n390), .ZN(new_n391));
  NOR3_X1   g0191(.A1(new_n255), .A2(new_n256), .A3(G20), .ZN(new_n392));
  OAI21_X1  g0192(.A(KEYINPUT74), .B1(new_n392), .B2(KEYINPUT7), .ZN(new_n393));
  AOI21_X1  g0193(.A(new_n391), .B1(new_n393), .B2(new_n389), .ZN(new_n394));
  OAI21_X1  g0194(.A(KEYINPUT75), .B1(new_n394), .B2(new_n341), .ZN(new_n395));
  XNOR2_X1  g0195(.A(G58), .B(G68), .ZN(new_n396));
  AOI22_X1  g0196(.A1(new_n396), .A2(G20), .B1(G159), .B2(new_n285), .ZN(new_n397));
  NAND3_X1  g0197(.A1(new_n392), .A2(KEYINPUT74), .A3(KEYINPUT7), .ZN(new_n398));
  NAND3_X1  g0198(.A1(new_n265), .A2(new_n210), .A3(new_n266), .ZN(new_n399));
  INV_X1    g0199(.A(KEYINPUT7), .ZN(new_n400));
  AOI21_X1  g0200(.A(new_n390), .B1(new_n399), .B2(new_n400), .ZN(new_n401));
  INV_X1    g0201(.A(new_n389), .ZN(new_n402));
  OAI21_X1  g0202(.A(new_n398), .B1(new_n401), .B2(new_n402), .ZN(new_n403));
  INV_X1    g0203(.A(KEYINPUT75), .ZN(new_n404));
  NAND3_X1  g0204(.A1(new_n403), .A2(new_n404), .A3(G68), .ZN(new_n405));
  NAND4_X1  g0205(.A1(new_n395), .A2(KEYINPUT16), .A3(new_n397), .A4(new_n405), .ZN(new_n406));
  INV_X1    g0206(.A(KEYINPUT16), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n399), .A2(new_n400), .ZN(new_n408));
  AOI21_X1  g0208(.A(new_n341), .B1(new_n408), .B2(new_n389), .ZN(new_n409));
  INV_X1    g0209(.A(new_n397), .ZN(new_n410));
  OAI21_X1  g0210(.A(new_n407), .B1(new_n409), .B2(new_n410), .ZN(new_n411));
  NAND3_X1  g0211(.A1(new_n406), .A2(new_n411), .A3(new_n291), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n295), .A2(new_n287), .ZN(new_n413));
  OAI21_X1  g0213(.A(new_n413), .B1(new_n297), .B2(new_n287), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n412), .A2(new_n414), .ZN(new_n415));
  INV_X1    g0215(.A(KEYINPUT77), .ZN(new_n416));
  AOI21_X1  g0216(.A(new_n416), .B1(new_n278), .B2(G232), .ZN(new_n417));
  NAND4_X1  g0217(.A1(new_n347), .A2(new_n348), .A3(new_n416), .A4(G232), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n418), .A2(new_n273), .ZN(new_n419));
  NOR2_X1   g0219(.A1(new_n417), .A2(new_n419), .ZN(new_n420));
  OAI211_X1 g0220(.A(G226), .B(G1698), .C1(new_n255), .C2(new_n256), .ZN(new_n421));
  NAND2_X1  g0221(.A1(G33), .A2(G87), .ZN(new_n422));
  OAI211_X1 g0222(.A(new_n421), .B(new_n422), .C1(new_n263), .C2(new_n269), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n423), .A2(new_n271), .ZN(new_n424));
  AND3_X1   g0224(.A1(new_n420), .A2(new_n424), .A3(KEYINPUT78), .ZN(new_n425));
  AOI21_X1  g0225(.A(KEYINPUT78), .B1(new_n420), .B2(new_n424), .ZN(new_n426));
  NOR3_X1   g0226(.A1(new_n425), .A2(new_n426), .A3(G169), .ZN(new_n427));
  INV_X1    g0227(.A(KEYINPUT76), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n424), .A2(new_n428), .ZN(new_n429));
  NAND3_X1  g0229(.A1(new_n423), .A2(KEYINPUT76), .A3(new_n271), .ZN(new_n430));
  NAND4_X1  g0230(.A1(new_n429), .A2(new_n305), .A3(new_n420), .A4(new_n430), .ZN(new_n431));
  INV_X1    g0231(.A(new_n431), .ZN(new_n432));
  OAI21_X1  g0232(.A(KEYINPUT79), .B1(new_n427), .B2(new_n432), .ZN(new_n433));
  INV_X1    g0233(.A(new_n426), .ZN(new_n434));
  NAND3_X1  g0234(.A1(new_n420), .A2(new_n424), .A3(KEYINPUT78), .ZN(new_n435));
  NAND3_X1  g0235(.A1(new_n434), .A2(new_n328), .A3(new_n435), .ZN(new_n436));
  INV_X1    g0236(.A(KEYINPUT79), .ZN(new_n437));
  NAND3_X1  g0237(.A1(new_n436), .A2(new_n431), .A3(new_n437), .ZN(new_n438));
  NAND3_X1  g0238(.A1(new_n415), .A2(new_n433), .A3(new_n438), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n439), .A2(KEYINPUT18), .ZN(new_n440));
  INV_X1    g0240(.A(KEYINPUT18), .ZN(new_n441));
  NAND4_X1  g0241(.A1(new_n415), .A2(new_n433), .A3(new_n441), .A4(new_n438), .ZN(new_n442));
  AND2_X1   g0242(.A1(new_n440), .A2(new_n442), .ZN(new_n443));
  INV_X1    g0243(.A(KEYINPUT80), .ZN(new_n444));
  NOR3_X1   g0244(.A1(new_n425), .A2(new_n426), .A3(G200), .ZN(new_n445));
  NOR3_X1   g0245(.A1(new_n417), .A2(new_n419), .A3(G190), .ZN(new_n446));
  NAND3_X1  g0246(.A1(new_n429), .A2(new_n430), .A3(new_n446), .ZN(new_n447));
  INV_X1    g0247(.A(new_n447), .ZN(new_n448));
  OAI21_X1  g0248(.A(new_n444), .B1(new_n445), .B2(new_n448), .ZN(new_n449));
  NAND3_X1  g0249(.A1(new_n434), .A2(new_n281), .A3(new_n435), .ZN(new_n450));
  NAND3_X1  g0250(.A1(new_n450), .A2(new_n447), .A3(KEYINPUT80), .ZN(new_n451));
  NAND4_X1  g0251(.A1(new_n449), .A2(new_n451), .A3(new_n412), .A4(new_n414), .ZN(new_n452));
  INV_X1    g0252(.A(KEYINPUT17), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  AND2_X1   g0254(.A1(new_n412), .A2(new_n414), .ZN(new_n455));
  NAND4_X1  g0255(.A1(new_n455), .A2(KEYINPUT17), .A3(new_n449), .A4(new_n451), .ZN(new_n456));
  AND2_X1   g0256(.A1(new_n454), .A2(new_n456), .ZN(new_n457));
  NAND3_X1  g0257(.A1(new_n388), .A2(new_n443), .A3(new_n457), .ZN(new_n458));
  INV_X1    g0258(.A(new_n458), .ZN(new_n459));
  INV_X1    g0259(.A(G33), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n460), .A2(G97), .ZN(new_n461));
  NAND2_X1  g0261(.A1(G33), .A2(G283), .ZN(new_n462));
  AOI21_X1  g0262(.A(G20), .B1(new_n461), .B2(new_n462), .ZN(new_n463));
  INV_X1    g0263(.A(G116), .ZN(new_n464));
  NOR2_X1   g0264(.A1(new_n210), .A2(new_n464), .ZN(new_n465));
  OAI21_X1  g0265(.A(new_n291), .B1(new_n463), .B2(new_n465), .ZN(new_n466));
  INV_X1    g0266(.A(KEYINPUT20), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  OAI211_X1 g0268(.A(KEYINPUT20), .B(new_n291), .C1(new_n463), .C2(new_n465), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  NOR2_X1   g0270(.A1(new_n295), .A2(G116), .ZN(new_n471));
  NOR2_X1   g0271(.A1(new_n460), .A2(G1), .ZN(new_n472));
  NOR3_X1   g0272(.A1(new_n294), .A2(new_n291), .A3(new_n472), .ZN(new_n473));
  AOI21_X1  g0273(.A(new_n471), .B1(new_n473), .B2(G116), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n470), .A2(new_n474), .ZN(new_n475));
  OAI211_X1 g0275(.A(G264), .B(G1698), .C1(new_n255), .C2(new_n256), .ZN(new_n476));
  NAND3_X1  g0276(.A1(new_n265), .A2(G303), .A3(new_n266), .ZN(new_n477));
  INV_X1    g0277(.A(G257), .ZN(new_n478));
  OAI211_X1 g0278(.A(new_n476), .B(new_n477), .C1(new_n263), .C2(new_n478), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n479), .A2(new_n271), .ZN(new_n480));
  XNOR2_X1  g0280(.A(KEYINPUT5), .B(G41), .ZN(new_n481));
  INV_X1    g0281(.A(G45), .ZN(new_n482));
  NOR2_X1   g0282(.A1(new_n482), .A2(G1), .ZN(new_n483));
  AOI22_X1  g0283(.A1(new_n481), .A2(new_n483), .B1(new_n276), .B2(new_n277), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n209), .A2(G45), .ZN(new_n485));
  OR2_X1    g0285(.A1(KEYINPUT5), .A2(G41), .ZN(new_n486));
  NAND2_X1  g0286(.A1(KEYINPUT5), .A2(G41), .ZN(new_n487));
  AOI21_X1  g0287(.A(new_n485), .B1(new_n486), .B2(new_n487), .ZN(new_n488));
  AOI22_X1  g0288(.A1(new_n484), .A2(G270), .B1(G274), .B2(new_n488), .ZN(new_n489));
  NAND4_X1  g0289(.A1(new_n475), .A2(G179), .A3(new_n480), .A4(new_n489), .ZN(new_n490));
  AOI21_X1  g0290(.A(new_n328), .B1(new_n470), .B2(new_n474), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n480), .A2(new_n489), .ZN(new_n492));
  AOI21_X1  g0292(.A(KEYINPUT86), .B1(new_n491), .B2(new_n492), .ZN(new_n493));
  INV_X1    g0293(.A(KEYINPUT21), .ZN(new_n494));
  OAI21_X1  g0294(.A(new_n490), .B1(new_n493), .B2(new_n494), .ZN(new_n495));
  AOI211_X1 g0295(.A(KEYINPUT86), .B(KEYINPUT21), .C1(new_n491), .C2(new_n492), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n492), .A2(new_n281), .ZN(new_n497));
  NAND3_X1  g0297(.A1(new_n480), .A2(new_n322), .A3(new_n489), .ZN(new_n498));
  AOI21_X1  g0298(.A(new_n475), .B1(new_n497), .B2(new_n498), .ZN(new_n499));
  NOR3_X1   g0299(.A1(new_n495), .A2(new_n496), .A3(new_n499), .ZN(new_n500));
  INV_X1    g0300(.A(G294), .ZN(new_n501));
  NOR2_X1   g0301(.A1(new_n460), .A2(new_n501), .ZN(new_n502));
  NOR2_X1   g0302(.A1(new_n257), .A2(new_n357), .ZN(new_n503));
  AOI21_X1  g0303(.A(new_n502), .B1(new_n503), .B2(G250), .ZN(new_n504));
  OAI211_X1 g0304(.A(G257), .B(G1698), .C1(new_n255), .C2(new_n256), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n505), .A2(KEYINPUT89), .ZN(new_n506));
  INV_X1    g0306(.A(KEYINPUT89), .ZN(new_n507));
  NAND4_X1  g0307(.A1(new_n267), .A2(new_n507), .A3(G257), .A4(G1698), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n506), .A2(new_n508), .ZN(new_n509));
  AOI21_X1  g0309(.A(new_n347), .B1(new_n504), .B2(new_n509), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n484), .A2(G264), .ZN(new_n511));
  INV_X1    g0311(.A(new_n511), .ZN(new_n512));
  NOR2_X1   g0312(.A1(new_n510), .A2(new_n512), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n488), .A2(G274), .ZN(new_n514));
  NAND3_X1  g0314(.A1(new_n513), .A2(G179), .A3(new_n514), .ZN(new_n515));
  INV_X1    g0315(.A(G250), .ZN(new_n516));
  OAI22_X1  g0316(.A1(new_n263), .A2(new_n516), .B1(new_n460), .B2(new_n501), .ZN(new_n517));
  AOI21_X1  g0317(.A(new_n517), .B1(new_n508), .B2(new_n506), .ZN(new_n518));
  OAI211_X1 g0318(.A(new_n514), .B(new_n511), .C1(new_n518), .C2(new_n347), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n519), .A2(G169), .ZN(new_n520));
  OAI211_X1 g0320(.A(new_n210), .B(G87), .C1(new_n255), .C2(new_n256), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n521), .A2(KEYINPUT87), .ZN(new_n522));
  INV_X1    g0322(.A(KEYINPUT87), .ZN(new_n523));
  NAND4_X1  g0323(.A1(new_n267), .A2(new_n523), .A3(new_n210), .A4(G87), .ZN(new_n524));
  NAND3_X1  g0324(.A1(new_n522), .A2(new_n524), .A3(KEYINPUT22), .ZN(new_n525));
  INV_X1    g0325(.A(KEYINPUT22), .ZN(new_n526));
  NAND3_X1  g0326(.A1(new_n521), .A2(KEYINPUT87), .A3(new_n526), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n206), .A2(G20), .ZN(new_n528));
  NAND3_X1  g0328(.A1(new_n528), .A2(KEYINPUT88), .A3(KEYINPUT23), .ZN(new_n529));
  INV_X1    g0329(.A(new_n529), .ZN(new_n530));
  NAND2_X1  g0330(.A1(G33), .A2(G116), .ZN(new_n531));
  OAI22_X1  g0331(.A1(new_n528), .A2(KEYINPUT23), .B1(G20), .B2(new_n531), .ZN(new_n532));
  AOI21_X1  g0332(.A(KEYINPUT88), .B1(new_n528), .B2(KEYINPUT23), .ZN(new_n533));
  NOR3_X1   g0333(.A1(new_n530), .A2(new_n532), .A3(new_n533), .ZN(new_n534));
  NAND3_X1  g0334(.A1(new_n525), .A2(new_n527), .A3(new_n534), .ZN(new_n535));
  INV_X1    g0335(.A(KEYINPUT24), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  NAND4_X1  g0337(.A1(new_n525), .A2(KEYINPUT24), .A3(new_n534), .A4(new_n527), .ZN(new_n538));
  NAND3_X1  g0338(.A1(new_n537), .A2(new_n291), .A3(new_n538), .ZN(new_n539));
  INV_X1    g0339(.A(new_n340), .ZN(new_n540));
  NOR2_X1   g0340(.A1(new_n540), .A2(new_n528), .ZN(new_n541));
  XOR2_X1   g0341(.A(new_n541), .B(KEYINPUT25), .Z(new_n542));
  AOI21_X1  g0342(.A(new_n542), .B1(G107), .B2(new_n473), .ZN(new_n543));
  AOI22_X1  g0343(.A1(new_n515), .A2(new_n520), .B1(new_n539), .B2(new_n543), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n539), .A2(new_n543), .ZN(new_n545));
  INV_X1    g0345(.A(new_n545), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n519), .A2(new_n281), .ZN(new_n547));
  OAI21_X1  g0347(.A(new_n547), .B1(G190), .B2(new_n519), .ZN(new_n548));
  AOI21_X1  g0348(.A(new_n544), .B1(new_n546), .B2(new_n548), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n310), .A2(new_n294), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n473), .A2(G87), .ZN(new_n551));
  OAI211_X1 g0351(.A(new_n210), .B(G68), .C1(new_n255), .C2(new_n256), .ZN(new_n552));
  INV_X1    g0352(.A(KEYINPUT19), .ZN(new_n553));
  OAI21_X1  g0353(.A(new_n553), .B1(new_n355), .B2(G20), .ZN(new_n554));
  NAND3_X1  g0354(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n555));
  INV_X1    g0355(.A(KEYINPUT84), .ZN(new_n556));
  NAND3_X1  g0356(.A1(new_n555), .A2(new_n556), .A3(new_n210), .ZN(new_n557));
  NOR2_X1   g0357(.A1(G87), .A2(G97), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n558), .A2(new_n206), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n557), .A2(new_n559), .ZN(new_n560));
  AOI21_X1  g0360(.A(new_n556), .B1(new_n555), .B2(new_n210), .ZN(new_n561));
  OAI211_X1 g0361(.A(new_n552), .B(new_n554), .C1(new_n560), .C2(new_n561), .ZN(new_n562));
  OAI21_X1  g0362(.A(new_n291), .B1(new_n562), .B2(KEYINPUT85), .ZN(new_n563));
  INV_X1    g0363(.A(KEYINPUT85), .ZN(new_n564));
  AND2_X1   g0364(.A1(new_n552), .A2(new_n554), .ZN(new_n565));
  INV_X1    g0365(.A(new_n561), .ZN(new_n566));
  NAND3_X1  g0366(.A1(new_n566), .A2(new_n557), .A3(new_n559), .ZN(new_n567));
  AOI21_X1  g0367(.A(new_n564), .B1(new_n565), .B2(new_n567), .ZN(new_n568));
  OAI211_X1 g0368(.A(new_n550), .B(new_n551), .C1(new_n563), .C2(new_n568), .ZN(new_n569));
  INV_X1    g0369(.A(new_n569), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n485), .A2(G250), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n483), .A2(G274), .ZN(new_n572));
  AOI21_X1  g0372(.A(new_n271), .B1(new_n571), .B2(new_n572), .ZN(new_n573));
  OAI211_X1 g0373(.A(G244), .B(G1698), .C1(new_n255), .C2(new_n256), .ZN(new_n574));
  OAI211_X1 g0374(.A(new_n531), .B(new_n574), .C1(new_n263), .C2(new_n319), .ZN(new_n575));
  AOI21_X1  g0375(.A(new_n573), .B1(new_n575), .B2(new_n271), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n576), .A2(new_n322), .ZN(new_n577));
  OAI21_X1  g0377(.A(new_n577), .B1(G200), .B2(new_n576), .ZN(new_n578));
  NOR2_X1   g0378(.A1(new_n576), .A2(G169), .ZN(new_n579));
  AOI211_X1 g0379(.A(G179), .B(new_n573), .C1(new_n575), .C2(new_n271), .ZN(new_n580));
  NOR2_X1   g0380(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  INV_X1    g0381(.A(new_n310), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n473), .A2(new_n582), .ZN(new_n583));
  OAI211_X1 g0383(.A(new_n550), .B(new_n583), .C1(new_n563), .C2(new_n568), .ZN(new_n584));
  AOI22_X1  g0384(.A1(new_n570), .A2(new_n578), .B1(new_n581), .B2(new_n584), .ZN(new_n585));
  NOR2_X1   g0385(.A1(new_n295), .A2(G97), .ZN(new_n586));
  AOI21_X1  g0386(.A(new_n586), .B1(new_n473), .B2(G97), .ZN(new_n587));
  INV_X1    g0387(.A(new_n587), .ZN(new_n588));
  XNOR2_X1  g0388(.A(G97), .B(G107), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n589), .A2(KEYINPUT82), .ZN(new_n590));
  INV_X1    g0390(.A(KEYINPUT6), .ZN(new_n591));
  INV_X1    g0391(.A(KEYINPUT82), .ZN(new_n592));
  NAND2_X1  g0392(.A1(G97), .A2(G107), .ZN(new_n593));
  NAND3_X1  g0393(.A1(new_n207), .A2(new_n592), .A3(new_n593), .ZN(new_n594));
  NAND3_X1  g0394(.A1(new_n590), .A2(new_n591), .A3(new_n594), .ZN(new_n595));
  NAND3_X1  g0395(.A1(new_n206), .A2(KEYINPUT6), .A3(G97), .ZN(new_n596));
  INV_X1    g0396(.A(KEYINPUT81), .ZN(new_n597));
  XNOR2_X1  g0397(.A(new_n596), .B(new_n597), .ZN(new_n598));
  AOI21_X1  g0398(.A(new_n210), .B1(new_n595), .B2(new_n598), .ZN(new_n599));
  INV_X1    g0399(.A(new_n599), .ZN(new_n600));
  AOI21_X1  g0400(.A(new_n206), .B1(new_n408), .B2(new_n389), .ZN(new_n601));
  NOR2_X1   g0401(.A1(new_n309), .A2(new_n226), .ZN(new_n602));
  NOR2_X1   g0402(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n600), .A2(new_n603), .ZN(new_n604));
  AOI21_X1  g0404(.A(new_n588), .B1(new_n604), .B2(new_n291), .ZN(new_n605));
  AOI21_X1  g0405(.A(new_n260), .B1(new_n265), .B2(new_n266), .ZN(new_n606));
  AOI22_X1  g0406(.A1(new_n606), .A2(G250), .B1(G33), .B2(G283), .ZN(new_n607));
  NAND2_X1  g0407(.A1(KEYINPUT83), .A2(KEYINPUT4), .ZN(new_n608));
  NOR2_X1   g0408(.A1(KEYINPUT83), .A2(KEYINPUT4), .ZN(new_n609));
  OAI21_X1  g0409(.A(G244), .B1(new_n255), .B2(new_n256), .ZN(new_n610));
  OAI211_X1 g0410(.A(new_n608), .B(new_n609), .C1(new_n610), .C2(new_n357), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n607), .A2(new_n611), .ZN(new_n612));
  NAND3_X1  g0412(.A1(new_n267), .A2(new_n373), .A3(G244), .ZN(new_n613));
  AOI21_X1  g0413(.A(new_n609), .B1(new_n613), .B2(new_n608), .ZN(new_n614));
  OAI21_X1  g0414(.A(new_n271), .B1(new_n612), .B2(new_n614), .ZN(new_n615));
  AOI22_X1  g0415(.A1(new_n484), .A2(G257), .B1(G274), .B2(new_n488), .ZN(new_n616));
  AND3_X1   g0416(.A1(new_n615), .A2(new_n322), .A3(new_n616), .ZN(new_n617));
  AOI21_X1  g0417(.A(G200), .B1(new_n615), .B2(new_n616), .ZN(new_n618));
  OAI21_X1  g0418(.A(new_n605), .B1(new_n617), .B2(new_n618), .ZN(new_n619));
  NOR3_X1   g0419(.A1(new_n599), .A2(new_n602), .A3(new_n601), .ZN(new_n620));
  INV_X1    g0420(.A(new_n291), .ZN(new_n621));
  OAI21_X1  g0421(.A(new_n587), .B1(new_n620), .B2(new_n621), .ZN(new_n622));
  AND3_X1   g0422(.A1(new_n615), .A2(G179), .A3(new_n616), .ZN(new_n623));
  AOI21_X1  g0423(.A(new_n328), .B1(new_n615), .B2(new_n616), .ZN(new_n624));
  OAI21_X1  g0424(.A(new_n622), .B1(new_n623), .B2(new_n624), .ZN(new_n625));
  AND3_X1   g0425(.A1(new_n585), .A2(new_n619), .A3(new_n625), .ZN(new_n626));
  AND4_X1   g0426(.A1(new_n459), .A2(new_n500), .A3(new_n549), .A4(new_n626), .ZN(G372));
  AND2_X1   g0427(.A1(new_n302), .A2(new_n303), .ZN(new_n628));
  INV_X1    g0428(.A(new_n383), .ZN(new_n629));
  AOI21_X1  g0429(.A(new_n387), .B1(new_n629), .B2(new_n330), .ZN(new_n630));
  AND2_X1   g0430(.A1(new_n457), .A2(new_n630), .ZN(new_n631));
  INV_X1    g0431(.A(new_n443), .ZN(new_n632));
  OAI21_X1  g0432(.A(new_n628), .B1(new_n631), .B2(new_n632), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n633), .A2(new_n307), .ZN(new_n634));
  AND2_X1   g0434(.A1(new_n570), .A2(new_n578), .ZN(new_n635));
  NOR2_X1   g0435(.A1(new_n635), .A2(KEYINPUT26), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n546), .A2(new_n548), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n637), .A2(new_n619), .ZN(new_n638));
  AOI21_X1  g0438(.A(new_n328), .B1(new_n513), .B2(new_n514), .ZN(new_n639));
  NOR2_X1   g0439(.A1(new_n519), .A2(new_n305), .ZN(new_n640));
  OAI21_X1  g0440(.A(new_n545), .B1(new_n639), .B2(new_n640), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n641), .A2(KEYINPUT91), .ZN(new_n642));
  INV_X1    g0442(.A(KEYINPUT91), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n544), .A2(new_n643), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n642), .A2(new_n644), .ZN(new_n645));
  NOR2_X1   g0445(.A1(new_n495), .A2(new_n496), .ZN(new_n646));
  AOI21_X1  g0446(.A(new_n638), .B1(new_n645), .B2(new_n646), .ZN(new_n647));
  INV_X1    g0447(.A(new_n625), .ZN(new_n648));
  OAI21_X1  g0448(.A(new_n636), .B1(new_n647), .B2(new_n648), .ZN(new_n649));
  INV_X1    g0449(.A(KEYINPUT26), .ZN(new_n650));
  AOI21_X1  g0450(.A(new_n650), .B1(new_n648), .B2(new_n585), .ZN(new_n651));
  NOR3_X1   g0451(.A1(new_n576), .A2(KEYINPUT90), .A3(G169), .ZN(new_n652));
  OR2_X1    g0452(.A1(new_n580), .A2(KEYINPUT90), .ZN(new_n653));
  INV_X1    g0453(.A(new_n579), .ZN(new_n654));
  AOI21_X1  g0454(.A(new_n652), .B1(new_n653), .B2(new_n654), .ZN(new_n655));
  AOI21_X1  g0455(.A(new_n651), .B1(new_n584), .B2(new_n655), .ZN(new_n656));
  AOI21_X1  g0456(.A(new_n458), .B1(new_n649), .B2(new_n656), .ZN(new_n657));
  OR2_X1    g0457(.A1(new_n634), .A2(new_n657), .ZN(G369));
  OR3_X1    g0458(.A1(new_n540), .A2(KEYINPUT27), .A3(G20), .ZN(new_n659));
  OAI21_X1  g0459(.A(KEYINPUT27), .B1(new_n540), .B2(G20), .ZN(new_n660));
  NAND3_X1  g0460(.A1(new_n659), .A2(G213), .A3(new_n660), .ZN(new_n661));
  INV_X1    g0461(.A(G343), .ZN(new_n662));
  NOR2_X1   g0462(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n545), .A2(new_n663), .ZN(new_n664));
  NAND3_X1  g0464(.A1(new_n637), .A2(new_n641), .A3(new_n664), .ZN(new_n665));
  XNOR2_X1  g0465(.A(new_n665), .B(KEYINPUT92), .ZN(new_n666));
  OAI211_X1 g0466(.A(new_n545), .B(new_n663), .C1(new_n639), .C2(new_n640), .ZN(new_n667));
  XNOR2_X1  g0467(.A(new_n667), .B(KEYINPUT93), .ZN(new_n668));
  INV_X1    g0468(.A(new_n668), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n666), .A2(new_n669), .ZN(new_n670));
  NOR2_X1   g0470(.A1(new_n646), .A2(new_n663), .ZN(new_n671));
  INV_X1    g0471(.A(new_n645), .ZN(new_n672));
  INV_X1    g0472(.A(new_n663), .ZN(new_n673));
  AOI22_X1  g0473(.A1(new_n670), .A2(new_n671), .B1(new_n672), .B2(new_n673), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n475), .A2(new_n663), .ZN(new_n675));
  INV_X1    g0475(.A(new_n675), .ZN(new_n676));
  OR2_X1    g0476(.A1(new_n500), .A2(new_n676), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n646), .A2(new_n676), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  INV_X1    g0479(.A(G330), .ZN(new_n680));
  NOR2_X1   g0480(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n670), .A2(new_n681), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n674), .A2(new_n682), .ZN(G399));
  INV_X1    g0483(.A(new_n213), .ZN(new_n684));
  NOR2_X1   g0484(.A1(new_n684), .A2(G41), .ZN(new_n685));
  INV_X1    g0485(.A(new_n685), .ZN(new_n686));
  NAND3_X1  g0486(.A1(new_n558), .A2(new_n206), .A3(new_n464), .ZN(new_n687));
  INV_X1    g0487(.A(new_n687), .ZN(new_n688));
  NAND3_X1  g0488(.A1(new_n686), .A2(G1), .A3(new_n688), .ZN(new_n689));
  INV_X1    g0489(.A(new_n222), .ZN(new_n690));
  OAI21_X1  g0490(.A(new_n689), .B1(new_n690), .B2(new_n686), .ZN(new_n691));
  XNOR2_X1  g0491(.A(new_n691), .B(KEYINPUT28), .ZN(new_n692));
  AOI21_X1  g0492(.A(new_n663), .B1(new_n649), .B2(new_n656), .ZN(new_n693));
  INV_X1    g0493(.A(KEYINPUT29), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  AOI21_X1  g0495(.A(new_n635), .B1(new_n584), .B2(new_n655), .ZN(new_n696));
  AND2_X1   g0496(.A1(new_n619), .A2(new_n625), .ZN(new_n697));
  NAND3_X1  g0497(.A1(new_n696), .A2(new_n697), .A3(new_n637), .ZN(new_n698));
  NOR3_X1   g0498(.A1(new_n544), .A2(new_n495), .A3(new_n496), .ZN(new_n699));
  NOR2_X1   g0499(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  NAND3_X1  g0500(.A1(new_n648), .A2(new_n650), .A3(new_n585), .ZN(new_n701));
  OAI21_X1  g0501(.A(KEYINPUT26), .B1(new_n625), .B2(new_n635), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n655), .A2(new_n584), .ZN(new_n703));
  NAND3_X1  g0503(.A1(new_n701), .A2(new_n702), .A3(new_n703), .ZN(new_n704));
  OAI21_X1  g0504(.A(new_n673), .B1(new_n700), .B2(new_n704), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n705), .A2(KEYINPUT29), .ZN(new_n706));
  INV_X1    g0506(.A(KEYINPUT31), .ZN(new_n707));
  NAND3_X1  g0507(.A1(new_n480), .A2(G179), .A3(new_n489), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n708), .A2(KEYINPUT94), .ZN(new_n709));
  INV_X1    g0509(.A(KEYINPUT94), .ZN(new_n710));
  NAND4_X1  g0510(.A1(new_n480), .A2(new_n489), .A3(new_n710), .A4(G179), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n709), .A2(new_n711), .ZN(new_n712));
  INV_X1    g0512(.A(new_n576), .ZN(new_n713));
  NOR3_X1   g0513(.A1(new_n713), .A2(new_n510), .A3(new_n512), .ZN(new_n714));
  AND2_X1   g0514(.A1(new_n615), .A2(new_n616), .ZN(new_n715));
  NAND4_X1  g0515(.A1(new_n712), .A2(KEYINPUT30), .A3(new_n714), .A4(new_n715), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n615), .A2(new_n616), .ZN(new_n717));
  AOI21_X1  g0517(.A(G179), .B1(new_n480), .B2(new_n489), .ZN(new_n718));
  NAND4_X1  g0518(.A1(new_n519), .A2(new_n717), .A3(new_n713), .A4(new_n718), .ZN(new_n719));
  NAND2_X1  g0519(.A1(new_n716), .A2(new_n719), .ZN(new_n720));
  OAI211_X1 g0520(.A(new_n511), .B(new_n576), .C1(new_n518), .C2(new_n347), .ZN(new_n721));
  NOR2_X1   g0521(.A1(new_n721), .A2(new_n717), .ZN(new_n722));
  AOI21_X1  g0522(.A(KEYINPUT30), .B1(new_n722), .B2(new_n712), .ZN(new_n723));
  OAI211_X1 g0523(.A(new_n707), .B(new_n663), .C1(new_n720), .C2(new_n723), .ZN(new_n724));
  INV_X1    g0524(.A(new_n724), .ZN(new_n725));
  NAND4_X1  g0525(.A1(new_n549), .A2(new_n626), .A3(new_n500), .A4(new_n673), .ZN(new_n726));
  INV_X1    g0526(.A(KEYINPUT30), .ZN(new_n727));
  INV_X1    g0527(.A(new_n712), .ZN(new_n728));
  NAND4_X1  g0528(.A1(new_n513), .A2(new_n576), .A3(new_n615), .A4(new_n616), .ZN(new_n729));
  OAI21_X1  g0529(.A(new_n727), .B1(new_n728), .B2(new_n729), .ZN(new_n730));
  NAND3_X1  g0530(.A1(new_n730), .A2(new_n716), .A3(new_n719), .ZN(new_n731));
  AOI21_X1  g0531(.A(new_n707), .B1(new_n731), .B2(new_n663), .ZN(new_n732));
  AOI21_X1  g0532(.A(new_n725), .B1(new_n726), .B2(new_n732), .ZN(new_n733));
  NAND2_X1  g0533(.A1(new_n733), .A2(G330), .ZN(new_n734));
  NAND3_X1  g0534(.A1(new_n695), .A2(new_n706), .A3(new_n734), .ZN(new_n735));
  INV_X1    g0535(.A(new_n735), .ZN(new_n736));
  OAI21_X1  g0536(.A(new_n692), .B1(new_n736), .B2(G1), .ZN(G364));
  XNOR2_X1  g0537(.A(new_n681), .B(KEYINPUT95), .ZN(new_n738));
  INV_X1    g0538(.A(new_n738), .ZN(new_n739));
  NOR2_X1   g0539(.A1(new_n293), .A2(G20), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n740), .A2(G45), .ZN(new_n741));
  NAND3_X1  g0541(.A1(new_n686), .A2(G1), .A3(new_n741), .ZN(new_n742));
  INV_X1    g0542(.A(new_n679), .ZN(new_n743));
  OAI211_X1 g0543(.A(new_n739), .B(new_n742), .C1(G330), .C2(new_n743), .ZN(new_n744));
  INV_X1    g0544(.A(new_n742), .ZN(new_n745));
  NOR2_X1   g0545(.A1(G13), .A2(G33), .ZN(new_n746));
  INV_X1    g0546(.A(new_n746), .ZN(new_n747));
  NOR2_X1   g0547(.A1(new_n747), .A2(G20), .ZN(new_n748));
  AOI21_X1  g0548(.A(new_n217), .B1(G20), .B2(new_n328), .ZN(new_n749));
  NOR2_X1   g0549(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  INV_X1    g0550(.A(new_n750), .ZN(new_n751));
  NAND2_X1  g0551(.A1(new_n213), .A2(new_n267), .ZN(new_n752));
  INV_X1    g0552(.A(G355), .ZN(new_n753));
  OAI22_X1  g0553(.A1(new_n752), .A2(new_n753), .B1(G116), .B2(new_n213), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n250), .A2(G45), .ZN(new_n755));
  OAI21_X1  g0555(.A(new_n755), .B1(G45), .B2(new_n222), .ZN(new_n756));
  NOR2_X1   g0556(.A1(new_n684), .A2(new_n267), .ZN(new_n757));
  AOI21_X1  g0557(.A(new_n754), .B1(new_n756), .B2(new_n757), .ZN(new_n758));
  NOR2_X1   g0558(.A1(new_n210), .A2(G190), .ZN(new_n759));
  NOR2_X1   g0559(.A1(G179), .A2(G200), .ZN(new_n760));
  NAND2_X1  g0560(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  INV_X1    g0561(.A(G159), .ZN(new_n762));
  NOR2_X1   g0562(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  XNOR2_X1  g0563(.A(new_n763), .B(KEYINPUT32), .ZN(new_n764));
  NOR2_X1   g0564(.A1(new_n305), .A2(G200), .ZN(new_n765));
  NAND2_X1  g0565(.A1(new_n759), .A2(new_n765), .ZN(new_n766));
  INV_X1    g0566(.A(new_n766), .ZN(new_n767));
  NOR2_X1   g0567(.A1(new_n281), .A2(G179), .ZN(new_n768));
  NAND2_X1  g0568(.A1(new_n768), .A2(new_n759), .ZN(new_n769));
  INV_X1    g0569(.A(new_n769), .ZN(new_n770));
  AOI22_X1  g0570(.A1(G77), .A2(new_n767), .B1(new_n770), .B2(G107), .ZN(new_n771));
  NOR2_X1   g0571(.A1(new_n305), .A2(new_n281), .ZN(new_n772));
  NAND2_X1  g0572(.A1(G20), .A2(G190), .ZN(new_n773));
  INV_X1    g0573(.A(new_n773), .ZN(new_n774));
  NAND2_X1  g0574(.A1(new_n772), .A2(new_n774), .ZN(new_n775));
  OAI211_X1 g0575(.A(new_n764), .B(new_n771), .C1(new_n202), .C2(new_n775), .ZN(new_n776));
  AOI21_X1  g0576(.A(new_n210), .B1(new_n760), .B2(G190), .ZN(new_n777));
  NOR2_X1   g0577(.A1(new_n777), .A2(new_n205), .ZN(new_n778));
  NAND2_X1  g0578(.A1(new_n772), .A2(new_n759), .ZN(new_n779));
  OAI21_X1  g0579(.A(new_n267), .B1(new_n779), .B2(new_n341), .ZN(new_n780));
  INV_X1    g0580(.A(G58), .ZN(new_n781));
  NAND2_X1  g0581(.A1(new_n765), .A2(new_n774), .ZN(new_n782));
  NAND2_X1  g0582(.A1(new_n768), .A2(new_n774), .ZN(new_n783));
  INV_X1    g0583(.A(G87), .ZN(new_n784));
  OAI22_X1  g0584(.A1(new_n781), .A2(new_n782), .B1(new_n783), .B2(new_n784), .ZN(new_n785));
  NOR4_X1   g0585(.A1(new_n776), .A2(new_n778), .A3(new_n780), .A4(new_n785), .ZN(new_n786));
  INV_X1    g0586(.A(new_n761), .ZN(new_n787));
  OR2_X1    g0587(.A1(new_n787), .A2(KEYINPUT97), .ZN(new_n788));
  NAND2_X1  g0588(.A1(new_n787), .A2(KEYINPUT97), .ZN(new_n789));
  NAND2_X1  g0589(.A1(new_n788), .A2(new_n789), .ZN(new_n790));
  INV_X1    g0590(.A(new_n790), .ZN(new_n791));
  AOI22_X1  g0591(.A1(new_n791), .A2(G329), .B1(G283), .B2(new_n770), .ZN(new_n792));
  XOR2_X1   g0592(.A(new_n792), .B(KEYINPUT98), .Z(new_n793));
  INV_X1    g0593(.A(G303), .ZN(new_n794));
  OAI21_X1  g0594(.A(new_n257), .B1(new_n783), .B2(new_n794), .ZN(new_n795));
  XNOR2_X1  g0595(.A(new_n795), .B(KEYINPUT96), .ZN(new_n796));
  NOR2_X1   g0596(.A1(new_n777), .A2(new_n501), .ZN(new_n797));
  INV_X1    g0597(.A(G326), .ZN(new_n798));
  INV_X1    g0598(.A(G322), .ZN(new_n799));
  OAI22_X1  g0599(.A1(new_n775), .A2(new_n798), .B1(new_n782), .B2(new_n799), .ZN(new_n800));
  XOR2_X1   g0600(.A(KEYINPUT33), .B(G317), .Z(new_n801));
  INV_X1    g0601(.A(G311), .ZN(new_n802));
  OAI22_X1  g0602(.A1(new_n801), .A2(new_n779), .B1(new_n766), .B2(new_n802), .ZN(new_n803));
  NOR4_X1   g0603(.A1(new_n796), .A2(new_n797), .A3(new_n800), .A4(new_n803), .ZN(new_n804));
  AOI21_X1  g0604(.A(new_n786), .B1(new_n793), .B2(new_n804), .ZN(new_n805));
  INV_X1    g0605(.A(new_n749), .ZN(new_n806));
  OAI221_X1 g0606(.A(new_n745), .B1(new_n751), .B2(new_n758), .C1(new_n805), .C2(new_n806), .ZN(new_n807));
  XOR2_X1   g0607(.A(new_n807), .B(KEYINPUT99), .Z(new_n808));
  INV_X1    g0608(.A(new_n748), .ZN(new_n809));
  OAI21_X1  g0609(.A(new_n808), .B1(new_n743), .B2(new_n809), .ZN(new_n810));
  NAND2_X1  g0610(.A1(new_n744), .A2(new_n810), .ZN(G396));
  OAI22_X1  g0611(.A1(new_n775), .A2(new_n794), .B1(new_n766), .B2(new_n464), .ZN(new_n812));
  OAI22_X1  g0612(.A1(new_n769), .A2(new_n784), .B1(new_n783), .B2(new_n206), .ZN(new_n813));
  OAI21_X1  g0613(.A(new_n257), .B1(new_n782), .B2(new_n501), .ZN(new_n814));
  NOR4_X1   g0614(.A1(new_n812), .A2(new_n813), .A3(new_n814), .A4(new_n778), .ZN(new_n815));
  INV_X1    g0615(.A(G283), .ZN(new_n816));
  AND2_X1   g0616(.A1(new_n779), .A2(KEYINPUT100), .ZN(new_n817));
  NOR2_X1   g0617(.A1(new_n779), .A2(KEYINPUT100), .ZN(new_n818));
  NOR2_X1   g0618(.A1(new_n817), .A2(new_n818), .ZN(new_n819));
  OAI221_X1 g0619(.A(new_n815), .B1(new_n816), .B2(new_n819), .C1(new_n802), .C2(new_n790), .ZN(new_n820));
  INV_X1    g0620(.A(new_n779), .ZN(new_n821));
  INV_X1    g0621(.A(new_n782), .ZN(new_n822));
  AOI22_X1  g0622(.A1(G150), .A2(new_n821), .B1(new_n822), .B2(G143), .ZN(new_n823));
  INV_X1    g0623(.A(G137), .ZN(new_n824));
  OAI221_X1 g0624(.A(new_n823), .B1(new_n824), .B2(new_n775), .C1(new_n762), .C2(new_n766), .ZN(new_n825));
  XOR2_X1   g0625(.A(new_n825), .B(KEYINPUT34), .Z(new_n826));
  NOR2_X1   g0626(.A1(new_n769), .A2(new_n341), .ZN(new_n827));
  OAI21_X1  g0627(.A(new_n267), .B1(new_n783), .B2(new_n202), .ZN(new_n828));
  INV_X1    g0628(.A(new_n777), .ZN(new_n829));
  AOI211_X1 g0629(.A(new_n827), .B(new_n828), .C1(G58), .C2(new_n829), .ZN(new_n830));
  INV_X1    g0630(.A(G132), .ZN(new_n831));
  OAI21_X1  g0631(.A(new_n830), .B1(new_n831), .B2(new_n790), .ZN(new_n832));
  OAI21_X1  g0632(.A(new_n820), .B1(new_n826), .B2(new_n832), .ZN(new_n833));
  NAND2_X1  g0633(.A1(new_n833), .A2(new_n749), .ZN(new_n834));
  NOR2_X1   g0634(.A1(new_n749), .A2(new_n746), .ZN(new_n835));
  AOI21_X1  g0635(.A(new_n742), .B1(new_n226), .B2(new_n835), .ZN(new_n836));
  OAI211_X1 g0636(.A(new_n325), .B(new_n330), .C1(new_n315), .C2(new_n673), .ZN(new_n837));
  XNOR2_X1  g0637(.A(new_n837), .B(KEYINPUT101), .ZN(new_n838));
  OR2_X1    g0638(.A1(new_n330), .A2(new_n673), .ZN(new_n839));
  NAND2_X1  g0639(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  OAI211_X1 g0640(.A(new_n834), .B(new_n836), .C1(new_n840), .C2(new_n747), .ZN(new_n841));
  INV_X1    g0641(.A(new_n841), .ZN(new_n842));
  INV_X1    g0642(.A(new_n840), .ZN(new_n843));
  XNOR2_X1  g0643(.A(new_n693), .B(new_n843), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n726), .A2(new_n732), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n845), .A2(new_n724), .ZN(new_n846));
  NOR2_X1   g0646(.A1(new_n846), .A2(new_n680), .ZN(new_n847));
  NOR2_X1   g0647(.A1(new_n844), .A2(new_n847), .ZN(new_n848));
  INV_X1    g0648(.A(new_n848), .ZN(new_n849));
  AOI21_X1  g0649(.A(new_n745), .B1(new_n844), .B2(new_n847), .ZN(new_n850));
  AOI21_X1  g0650(.A(new_n842), .B1(new_n849), .B2(new_n850), .ZN(new_n851));
  INV_X1    g0651(.A(new_n851), .ZN(G384));
  NOR2_X1   g0652(.A1(new_n740), .A2(new_n209), .ZN(new_n853));
  NAND4_X1  g0653(.A1(new_n454), .A2(new_n440), .A3(new_n442), .A4(new_n456), .ZN(new_n854));
  AND2_X1   g0654(.A1(new_n405), .A2(new_n397), .ZN(new_n855));
  AOI21_X1  g0655(.A(KEYINPUT16), .B1(new_n855), .B2(new_n395), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n406), .A2(new_n291), .ZN(new_n857));
  OAI21_X1  g0657(.A(new_n414), .B1(new_n856), .B2(new_n857), .ZN(new_n858));
  INV_X1    g0658(.A(new_n661), .ZN(new_n859));
  AND2_X1   g0659(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n854), .A2(new_n860), .ZN(new_n861));
  INV_X1    g0661(.A(KEYINPUT37), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n415), .A2(new_n859), .ZN(new_n863));
  NAND4_X1  g0663(.A1(new_n452), .A2(new_n439), .A3(new_n862), .A4(new_n863), .ZN(new_n864));
  NOR3_X1   g0664(.A1(new_n427), .A2(new_n432), .A3(KEYINPUT79), .ZN(new_n865));
  AOI21_X1  g0665(.A(new_n437), .B1(new_n436), .B2(new_n431), .ZN(new_n866));
  OAI21_X1  g0666(.A(new_n661), .B1(new_n865), .B2(new_n866), .ZN(new_n867));
  NOR3_X1   g0667(.A1(new_n445), .A2(new_n444), .A3(new_n448), .ZN(new_n868));
  AOI21_X1  g0668(.A(KEYINPUT80), .B1(new_n450), .B2(new_n447), .ZN(new_n869));
  NOR2_X1   g0669(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  AOI22_X1  g0670(.A1(new_n867), .A2(new_n858), .B1(new_n870), .B2(new_n455), .ZN(new_n871));
  OAI21_X1  g0671(.A(new_n864), .B1(new_n871), .B2(new_n862), .ZN(new_n872));
  AND3_X1   g0672(.A1(new_n861), .A2(KEYINPUT38), .A3(new_n872), .ZN(new_n873));
  INV_X1    g0673(.A(new_n863), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n854), .A2(new_n874), .ZN(new_n875));
  NAND3_X1  g0675(.A1(new_n452), .A2(new_n439), .A3(new_n863), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n876), .A2(KEYINPUT37), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n877), .A2(new_n864), .ZN(new_n878));
  AOI21_X1  g0678(.A(KEYINPUT38), .B1(new_n875), .B2(new_n878), .ZN(new_n879));
  OAI21_X1  g0679(.A(KEYINPUT104), .B1(new_n873), .B2(new_n879), .ZN(new_n880));
  NAND3_X1  g0680(.A1(new_n861), .A2(new_n872), .A3(KEYINPUT38), .ZN(new_n881));
  INV_X1    g0681(.A(KEYINPUT104), .ZN(new_n882));
  AOI22_X1  g0682(.A1(new_n854), .A2(new_n874), .B1(new_n877), .B2(new_n864), .ZN(new_n883));
  OAI211_X1 g0683(.A(new_n881), .B(new_n882), .C1(KEYINPUT38), .C2(new_n883), .ZN(new_n884));
  INV_X1    g0684(.A(KEYINPUT102), .ZN(new_n885));
  OAI21_X1  g0685(.A(new_n885), .B1(new_n383), .B2(new_n387), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n345), .A2(new_n663), .ZN(new_n887));
  AOI22_X1  g0687(.A1(new_n366), .A2(new_n367), .B1(new_n379), .B2(new_n381), .ZN(new_n888));
  OAI211_X1 g0688(.A(KEYINPUT102), .B(new_n386), .C1(new_n888), .C2(new_n346), .ZN(new_n889));
  AND3_X1   g0689(.A1(new_n886), .A2(new_n887), .A3(new_n889), .ZN(new_n890));
  AOI21_X1  g0690(.A(new_n887), .B1(new_n886), .B2(new_n889), .ZN(new_n891));
  OAI211_X1 g0691(.A(new_n733), .B(new_n840), .C1(new_n890), .C2(new_n891), .ZN(new_n892));
  INV_X1    g0692(.A(KEYINPUT40), .ZN(new_n893));
  NOR2_X1   g0693(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  NAND3_X1  g0694(.A1(new_n880), .A2(new_n884), .A3(new_n894), .ZN(new_n895));
  INV_X1    g0695(.A(new_n892), .ZN(new_n896));
  AOI21_X1  g0696(.A(KEYINPUT38), .B1(new_n861), .B2(new_n872), .ZN(new_n897));
  OAI21_X1  g0697(.A(new_n896), .B1(new_n873), .B2(new_n897), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n898), .A2(new_n893), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n895), .A2(new_n899), .ZN(new_n900));
  NOR2_X1   g0700(.A1(new_n458), .A2(new_n846), .ZN(new_n901));
  XNOR2_X1  g0701(.A(new_n900), .B(new_n901), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n902), .A2(G330), .ZN(new_n903));
  XOR2_X1   g0703(.A(new_n903), .B(KEYINPUT105), .Z(new_n904));
  INV_X1    g0704(.A(new_n904), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n861), .A2(new_n872), .ZN(new_n906));
  INV_X1    g0706(.A(KEYINPUT38), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  INV_X1    g0708(.A(KEYINPUT103), .ZN(new_n909));
  OAI211_X1 g0709(.A(new_n908), .B(new_n881), .C1(new_n909), .C2(new_n879), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n910), .A2(KEYINPUT39), .ZN(new_n911));
  NOR2_X1   g0711(.A1(new_n873), .A2(new_n879), .ZN(new_n912));
  NOR2_X1   g0712(.A1(KEYINPUT103), .A2(KEYINPUT39), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n911), .A2(new_n914), .ZN(new_n915));
  NOR2_X1   g0715(.A1(new_n629), .A2(new_n663), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  OR2_X1    g0717(.A1(new_n330), .A2(new_n663), .ZN(new_n918));
  INV_X1    g0718(.A(new_n918), .ZN(new_n919));
  AOI21_X1  g0719(.A(new_n919), .B1(new_n693), .B2(new_n840), .ZN(new_n920));
  NOR2_X1   g0720(.A1(new_n890), .A2(new_n891), .ZN(new_n921));
  NOR2_X1   g0721(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n908), .A2(new_n881), .ZN(new_n923));
  AOI22_X1  g0723(.A1(new_n922), .A2(new_n923), .B1(new_n632), .B2(new_n661), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n917), .A2(new_n924), .ZN(new_n925));
  AOI21_X1  g0725(.A(new_n458), .B1(new_n695), .B2(new_n706), .ZN(new_n926));
  NOR2_X1   g0726(.A1(new_n926), .A2(new_n634), .ZN(new_n927));
  XOR2_X1   g0727(.A(new_n925), .B(new_n927), .Z(new_n928));
  AOI21_X1  g0728(.A(new_n853), .B1(new_n905), .B2(new_n928), .ZN(new_n929));
  OAI21_X1  g0729(.A(new_n929), .B1(new_n905), .B2(new_n928), .ZN(new_n930));
  OAI21_X1  g0730(.A(G77), .B1(new_n781), .B2(new_n341), .ZN(new_n931));
  OAI22_X1  g0731(.A1(new_n690), .A2(new_n931), .B1(G50), .B2(new_n341), .ZN(new_n932));
  NAND3_X1  g0732(.A1(new_n932), .A2(G1), .A3(new_n293), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n595), .A2(new_n598), .ZN(new_n934));
  OAI211_X1 g0734(.A(G116), .B(new_n218), .C1(new_n934), .C2(KEYINPUT35), .ZN(new_n935));
  AOI21_X1  g0735(.A(new_n935), .B1(KEYINPUT35), .B2(new_n934), .ZN(new_n936));
  XOR2_X1   g0736(.A(new_n936), .B(KEYINPUT36), .Z(new_n937));
  NAND3_X1  g0737(.A1(new_n930), .A2(new_n933), .A3(new_n937), .ZN(G367));
  OAI21_X1  g0738(.A(new_n697), .B1(new_n605), .B2(new_n673), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n648), .A2(new_n663), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n939), .A2(new_n940), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n941), .A2(KEYINPUT106), .ZN(new_n942));
  INV_X1    g0742(.A(KEYINPUT106), .ZN(new_n943));
  NAND3_X1  g0743(.A1(new_n939), .A2(new_n943), .A3(new_n940), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n942), .A2(new_n944), .ZN(new_n945));
  INV_X1    g0745(.A(new_n945), .ZN(new_n946));
  NOR2_X1   g0746(.A1(new_n682), .A2(new_n946), .ZN(new_n947));
  XNOR2_X1  g0747(.A(new_n947), .B(KEYINPUT107), .ZN(new_n948));
  NOR2_X1   g0748(.A1(new_n570), .A2(new_n673), .ZN(new_n949));
  NOR2_X1   g0749(.A1(new_n696), .A2(new_n949), .ZN(new_n950));
  AND2_X1   g0750(.A1(new_n703), .A2(new_n949), .ZN(new_n951));
  NOR2_X1   g0751(.A1(new_n950), .A2(new_n951), .ZN(new_n952));
  INV_X1    g0752(.A(new_n952), .ZN(new_n953));
  INV_X1    g0753(.A(KEYINPUT43), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n953), .A2(new_n954), .ZN(new_n955));
  XNOR2_X1  g0755(.A(new_n948), .B(new_n955), .ZN(new_n956));
  AOI21_X1  g0756(.A(new_n648), .B1(new_n945), .B2(new_n544), .ZN(new_n957));
  NAND3_X1  g0757(.A1(new_n945), .A2(new_n670), .A3(new_n671), .ZN(new_n958));
  OAI22_X1  g0758(.A1(new_n957), .A2(new_n663), .B1(new_n958), .B2(KEYINPUT42), .ZN(new_n959));
  AND2_X1   g0759(.A1(new_n958), .A2(KEYINPUT42), .ZN(new_n960));
  OAI22_X1  g0760(.A1(new_n959), .A2(new_n960), .B1(new_n954), .B2(new_n953), .ZN(new_n961));
  XNOR2_X1  g0761(.A(new_n956), .B(new_n961), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n741), .A2(G1), .ZN(new_n963));
  INV_X1    g0763(.A(new_n963), .ZN(new_n964));
  XNOR2_X1  g0764(.A(KEYINPUT108), .B(KEYINPUT41), .ZN(new_n965));
  XOR2_X1   g0765(.A(new_n685), .B(new_n965), .Z(new_n966));
  NAND2_X1  g0766(.A1(new_n670), .A2(new_n671), .ZN(new_n967));
  OR2_X1    g0767(.A1(new_n665), .A2(KEYINPUT92), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n665), .A2(KEYINPUT92), .ZN(new_n969));
  AOI21_X1  g0769(.A(new_n668), .B1(new_n968), .B2(new_n969), .ZN(new_n970));
  INV_X1    g0770(.A(new_n671), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n970), .A2(new_n971), .ZN(new_n972));
  NAND4_X1  g0772(.A1(new_n967), .A2(KEYINPUT109), .A3(new_n972), .A4(new_n681), .ZN(new_n973));
  AND2_X1   g0773(.A1(new_n967), .A2(new_n972), .ZN(new_n974));
  OAI21_X1  g0774(.A(new_n973), .B1(new_n974), .B2(new_n738), .ZN(new_n975));
  AOI21_X1  g0775(.A(KEYINPUT109), .B1(new_n974), .B2(new_n681), .ZN(new_n976));
  NOR3_X1   g0776(.A1(new_n975), .A2(new_n976), .A3(new_n735), .ZN(new_n977));
  INV_X1    g0777(.A(new_n682), .ZN(new_n978));
  NAND2_X1  g0778(.A1(new_n672), .A2(new_n673), .ZN(new_n979));
  OAI211_X1 g0779(.A(new_n945), .B(new_n979), .C1(new_n970), .C2(new_n971), .ZN(new_n980));
  XNOR2_X1  g0780(.A(new_n980), .B(KEYINPUT45), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n967), .A2(new_n979), .ZN(new_n982));
  INV_X1    g0782(.A(KEYINPUT44), .ZN(new_n983));
  NAND3_X1  g0783(.A1(new_n982), .A2(new_n983), .A3(new_n946), .ZN(new_n984));
  OAI21_X1  g0784(.A(KEYINPUT44), .B1(new_n674), .B2(new_n945), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n984), .A2(new_n985), .ZN(new_n986));
  OAI21_X1  g0786(.A(new_n978), .B1(new_n981), .B2(new_n986), .ZN(new_n987));
  INV_X1    g0787(.A(KEYINPUT45), .ZN(new_n988));
  XNOR2_X1  g0788(.A(new_n980), .B(new_n988), .ZN(new_n989));
  NAND4_X1  g0789(.A1(new_n989), .A2(new_n682), .A3(new_n985), .A4(new_n984), .ZN(new_n990));
  NAND3_X1  g0790(.A1(new_n977), .A2(new_n987), .A3(new_n990), .ZN(new_n991));
  AOI21_X1  g0791(.A(new_n966), .B1(new_n991), .B2(new_n736), .ZN(new_n992));
  INV_X1    g0792(.A(KEYINPUT110), .ZN(new_n993));
  OAI21_X1  g0793(.A(new_n964), .B1(new_n992), .B2(new_n993), .ZN(new_n994));
  AOI211_X1 g0794(.A(KEYINPUT110), .B(new_n966), .C1(new_n991), .C2(new_n736), .ZN(new_n995));
  OAI21_X1  g0795(.A(new_n962), .B1(new_n994), .B2(new_n995), .ZN(new_n996));
  NAND2_X1  g0796(.A1(new_n246), .A2(new_n757), .ZN(new_n997));
  AOI21_X1  g0797(.A(new_n751), .B1(new_n684), .B2(new_n582), .ZN(new_n998));
  AOI21_X1  g0798(.A(new_n742), .B1(new_n997), .B2(new_n998), .ZN(new_n999));
  INV_X1    g0799(.A(new_n783), .ZN(new_n1000));
  AOI22_X1  g0800(.A1(new_n767), .A2(G50), .B1(new_n1000), .B2(G58), .ZN(new_n1001));
  INV_X1    g0801(.A(G143), .ZN(new_n1002));
  OAI21_X1  g0802(.A(new_n1001), .B1(new_n1002), .B2(new_n775), .ZN(new_n1003));
  INV_X1    g0803(.A(new_n819), .ZN(new_n1004));
  AOI21_X1  g0804(.A(new_n1003), .B1(G159), .B2(new_n1004), .ZN(new_n1005));
  NAND2_X1  g0805(.A1(new_n829), .A2(G68), .ZN(new_n1006));
  INV_X1    g0806(.A(G150), .ZN(new_n1007));
  OAI22_X1  g0807(.A1(new_n769), .A2(new_n226), .B1(new_n782), .B2(new_n1007), .ZN(new_n1008));
  AOI211_X1 g0808(.A(new_n257), .B(new_n1008), .C1(G137), .C2(new_n787), .ZN(new_n1009));
  NAND3_X1  g0809(.A1(new_n1005), .A2(new_n1006), .A3(new_n1009), .ZN(new_n1010));
  INV_X1    g0810(.A(G317), .ZN(new_n1011));
  OAI22_X1  g0811(.A1(new_n769), .A2(new_n205), .B1(new_n761), .B2(new_n1011), .ZN(new_n1012));
  OAI22_X1  g0812(.A1(new_n766), .A2(new_n816), .B1(new_n782), .B2(new_n794), .ZN(new_n1013));
  AOI211_X1 g0813(.A(new_n1012), .B(new_n1013), .C1(new_n1004), .C2(G294), .ZN(new_n1014));
  OAI21_X1  g0814(.A(new_n257), .B1(new_n775), .B2(new_n802), .ZN(new_n1015));
  NOR2_X1   g0815(.A1(new_n783), .A2(new_n464), .ZN(new_n1016));
  OAI22_X1  g0816(.A1(new_n1016), .A2(KEYINPUT46), .B1(new_n206), .B2(new_n777), .ZN(new_n1017));
  AOI211_X1 g0817(.A(new_n1015), .B(new_n1017), .C1(KEYINPUT46), .C2(new_n1016), .ZN(new_n1018));
  NAND2_X1  g0818(.A1(new_n1014), .A2(new_n1018), .ZN(new_n1019));
  AOI21_X1  g0819(.A(KEYINPUT47), .B1(new_n1010), .B2(new_n1019), .ZN(new_n1020));
  NAND3_X1  g0820(.A1(new_n1010), .A2(new_n1019), .A3(KEYINPUT47), .ZN(new_n1021));
  NAND2_X1  g0821(.A1(new_n1021), .A2(new_n749), .ZN(new_n1022));
  OAI221_X1 g0822(.A(new_n999), .B1(new_n1020), .B2(new_n1022), .C1(new_n952), .C2(new_n809), .ZN(new_n1023));
  NAND2_X1  g0823(.A1(new_n996), .A2(new_n1023), .ZN(G387));
  NOR2_X1   g0824(.A1(new_n977), .A2(new_n686), .ZN(new_n1025));
  NOR2_X1   g0825(.A1(new_n975), .A2(new_n976), .ZN(new_n1026));
  OAI21_X1  g0826(.A(new_n1025), .B1(new_n736), .B2(new_n1026), .ZN(new_n1027));
  NAND2_X1  g0827(.A1(new_n970), .A2(new_n748), .ZN(new_n1028));
  OAI22_X1  g0828(.A1(new_n752), .A2(new_n688), .B1(G107), .B2(new_n213), .ZN(new_n1029));
  NAND2_X1  g0829(.A1(new_n241), .A2(G45), .ZN(new_n1030));
  INV_X1    g0830(.A(new_n757), .ZN(new_n1031));
  NOR2_X1   g0831(.A1(new_n287), .A2(G50), .ZN(new_n1032));
  XNOR2_X1  g0832(.A(new_n1032), .B(KEYINPUT50), .ZN(new_n1033));
  AOI211_X1 g0833(.A(G45), .B(new_n687), .C1(G68), .C2(G77), .ZN(new_n1034));
  AOI21_X1  g0834(.A(new_n1031), .B1(new_n1033), .B2(new_n1034), .ZN(new_n1035));
  AOI21_X1  g0835(.A(new_n1029), .B1(new_n1030), .B2(new_n1035), .ZN(new_n1036));
  OAI21_X1  g0836(.A(new_n745), .B1(new_n1036), .B2(new_n751), .ZN(new_n1037));
  OAI22_X1  g0837(.A1(new_n775), .A2(new_n762), .B1(new_n766), .B2(new_n341), .ZN(new_n1038));
  OAI22_X1  g0838(.A1(new_n779), .A2(new_n287), .B1(new_n782), .B2(new_n202), .ZN(new_n1039));
  NOR2_X1   g0839(.A1(new_n777), .A2(new_n310), .ZN(new_n1040));
  NOR3_X1   g0840(.A1(new_n1038), .A2(new_n1039), .A3(new_n1040), .ZN(new_n1041));
  NAND2_X1  g0841(.A1(new_n1000), .A2(G77), .ZN(new_n1042));
  OAI21_X1  g0842(.A(new_n1042), .B1(new_n1007), .B2(new_n761), .ZN(new_n1043));
  OAI21_X1  g0843(.A(new_n267), .B1(new_n769), .B2(new_n205), .ZN(new_n1044));
  NOR2_X1   g0844(.A1(new_n1043), .A2(new_n1044), .ZN(new_n1045));
  INV_X1    g0845(.A(KEYINPUT111), .ZN(new_n1046));
  NOR2_X1   g0846(.A1(new_n1045), .A2(new_n1046), .ZN(new_n1047));
  NOR3_X1   g0847(.A1(new_n1043), .A2(KEYINPUT111), .A3(new_n1044), .ZN(new_n1048));
  OAI21_X1  g0848(.A(new_n1041), .B1(new_n1047), .B2(new_n1048), .ZN(new_n1049));
  XNOR2_X1  g0849(.A(new_n1049), .B(KEYINPUT112), .ZN(new_n1050));
  AOI21_X1  g0850(.A(new_n267), .B1(new_n770), .B2(G116), .ZN(new_n1051));
  OAI22_X1  g0851(.A1(new_n783), .A2(new_n501), .B1(new_n777), .B2(new_n816), .ZN(new_n1052));
  INV_X1    g0852(.A(new_n775), .ZN(new_n1053));
  AOI22_X1  g0853(.A1(new_n1053), .A2(G322), .B1(new_n767), .B2(G303), .ZN(new_n1054));
  OAI21_X1  g0854(.A(new_n1054), .B1(new_n1011), .B2(new_n782), .ZN(new_n1055));
  AOI21_X1  g0855(.A(new_n1055), .B1(G311), .B2(new_n1004), .ZN(new_n1056));
  AOI21_X1  g0856(.A(new_n1052), .B1(new_n1056), .B2(KEYINPUT48), .ZN(new_n1057));
  OAI21_X1  g0857(.A(new_n1057), .B1(KEYINPUT48), .B2(new_n1056), .ZN(new_n1058));
  INV_X1    g0858(.A(KEYINPUT49), .ZN(new_n1059));
  OAI221_X1 g0859(.A(new_n1051), .B1(new_n798), .B2(new_n761), .C1(new_n1058), .C2(new_n1059), .ZN(new_n1060));
  AND2_X1   g0860(.A1(new_n1058), .A2(new_n1059), .ZN(new_n1061));
  OAI21_X1  g0861(.A(new_n1050), .B1(new_n1060), .B2(new_n1061), .ZN(new_n1062));
  AOI21_X1  g0862(.A(new_n1037), .B1(new_n1062), .B2(new_n749), .ZN(new_n1063));
  AOI22_X1  g0863(.A1(new_n1026), .A2(new_n963), .B1(new_n1028), .B2(new_n1063), .ZN(new_n1064));
  NAND2_X1  g0864(.A1(new_n1027), .A2(new_n1064), .ZN(G393));
  OAI221_X1 g0865(.A(new_n750), .B1(new_n205), .B2(new_n213), .C1(new_n1031), .C2(new_n253), .ZN(new_n1066));
  NAND2_X1  g0866(.A1(new_n1066), .A2(new_n745), .ZN(new_n1067));
  NAND2_X1  g0867(.A1(new_n1004), .A2(G50), .ZN(new_n1068));
  OAI22_X1  g0868(.A1(new_n775), .A2(new_n1007), .B1(new_n782), .B2(new_n762), .ZN(new_n1069));
  XNOR2_X1  g0869(.A(new_n1069), .B(KEYINPUT51), .ZN(new_n1070));
  OAI22_X1  g0870(.A1(new_n783), .A2(new_n341), .B1(new_n761), .B2(new_n1002), .ZN(new_n1071));
  INV_X1    g0871(.A(new_n287), .ZN(new_n1072));
  AOI21_X1  g0872(.A(new_n1071), .B1(new_n1072), .B2(new_n767), .ZN(new_n1073));
  OAI21_X1  g0873(.A(new_n267), .B1(new_n769), .B2(new_n784), .ZN(new_n1074));
  AOI21_X1  g0874(.A(new_n1074), .B1(G77), .B2(new_n829), .ZN(new_n1075));
  NAND4_X1  g0875(.A1(new_n1068), .A2(new_n1070), .A3(new_n1073), .A4(new_n1075), .ZN(new_n1076));
  AOI22_X1  g0876(.A1(G283), .A2(new_n1000), .B1(new_n787), .B2(G322), .ZN(new_n1077));
  OAI211_X1 g0877(.A(new_n1077), .B(new_n257), .C1(new_n206), .C2(new_n769), .ZN(new_n1078));
  XNOR2_X1  g0878(.A(new_n1078), .B(KEYINPUT113), .ZN(new_n1079));
  OAI22_X1  g0879(.A1(new_n775), .A2(new_n1011), .B1(new_n782), .B2(new_n802), .ZN(new_n1080));
  XNOR2_X1  g0880(.A(new_n1080), .B(KEYINPUT52), .ZN(new_n1081));
  AOI22_X1  g0881(.A1(G294), .A2(new_n767), .B1(new_n829), .B2(G116), .ZN(new_n1082));
  OAI211_X1 g0882(.A(new_n1081), .B(new_n1082), .C1(new_n794), .C2(new_n819), .ZN(new_n1083));
  OAI21_X1  g0883(.A(new_n1076), .B1(new_n1079), .B2(new_n1083), .ZN(new_n1084));
  AOI21_X1  g0884(.A(new_n1067), .B1(new_n1084), .B2(new_n749), .ZN(new_n1085));
  OAI21_X1  g0885(.A(new_n1085), .B1(new_n945), .B2(new_n809), .ZN(new_n1086));
  NAND2_X1  g0886(.A1(new_n987), .A2(new_n990), .ZN(new_n1087));
  OAI21_X1  g0887(.A(new_n1086), .B1(new_n1087), .B2(new_n964), .ZN(new_n1088));
  INV_X1    g0888(.A(new_n1087), .ZN(new_n1089));
  OR2_X1    g0889(.A1(new_n1089), .A2(new_n977), .ZN(new_n1090));
  AND2_X1   g0890(.A1(new_n991), .A2(new_n685), .ZN(new_n1091));
  AOI21_X1  g0891(.A(new_n1088), .B1(new_n1090), .B2(new_n1091), .ZN(new_n1092));
  INV_X1    g0892(.A(new_n1092), .ZN(G390));
  INV_X1    g0893(.A(new_n916), .ZN(new_n1094));
  OAI21_X1  g0894(.A(new_n1094), .B1(new_n920), .B2(new_n921), .ZN(new_n1095));
  NAND3_X1  g0895(.A1(new_n911), .A2(new_n1095), .A3(new_n914), .ZN(new_n1096));
  XOR2_X1   g0896(.A(new_n837), .B(KEYINPUT101), .Z(new_n1097));
  OAI211_X1 g0897(.A(new_n1097), .B(new_n673), .C1(new_n700), .C2(new_n704), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n1098), .A2(new_n918), .ZN(new_n1099));
  OR2_X1    g0899(.A1(new_n890), .A2(new_n891), .ZN(new_n1100));
  AOI21_X1  g0900(.A(new_n916), .B1(new_n1099), .B2(new_n1100), .ZN(new_n1101));
  NAND3_X1  g0901(.A1(new_n1101), .A2(new_n880), .A3(new_n884), .ZN(new_n1102));
  NAND2_X1  g0902(.A1(new_n1096), .A2(new_n1102), .ZN(new_n1103));
  INV_X1    g0903(.A(KEYINPUT114), .ZN(new_n1104));
  NAND4_X1  g0904(.A1(new_n847), .A2(new_n1100), .A3(new_n1104), .A4(new_n840), .ZN(new_n1105));
  OAI21_X1  g0905(.A(new_n840), .B1(new_n890), .B2(new_n891), .ZN(new_n1106));
  OAI21_X1  g0906(.A(KEYINPUT114), .B1(new_n1106), .B2(new_n734), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n1105), .A2(new_n1107), .ZN(new_n1108));
  INV_X1    g0908(.A(new_n1108), .ZN(new_n1109));
  NAND2_X1  g0909(.A1(new_n1103), .A2(new_n1109), .ZN(new_n1110));
  INV_X1    g0910(.A(new_n1106), .ZN(new_n1111));
  NAND2_X1  g0911(.A1(new_n1111), .A2(new_n847), .ZN(new_n1112));
  NAND3_X1  g0912(.A1(new_n1096), .A2(new_n1102), .A3(new_n1112), .ZN(new_n1113));
  NAND2_X1  g0913(.A1(new_n1110), .A2(new_n1113), .ZN(new_n1114));
  OAI21_X1  g0914(.A(new_n921), .B1(new_n734), .B2(new_n843), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n1108), .A2(new_n1115), .ZN(new_n1116));
  INV_X1    g0916(.A(new_n920), .ZN(new_n1117));
  NAND2_X1  g0917(.A1(new_n1116), .A2(new_n1117), .ZN(new_n1118));
  NAND2_X1  g0918(.A1(new_n734), .A2(KEYINPUT115), .ZN(new_n1119));
  INV_X1    g0919(.A(new_n1119), .ZN(new_n1120));
  NOR2_X1   g0920(.A1(new_n734), .A2(KEYINPUT115), .ZN(new_n1121));
  OAI21_X1  g0921(.A(new_n840), .B1(new_n1120), .B2(new_n1121), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n1122), .A2(new_n921), .ZN(new_n1123));
  OAI211_X1 g0923(.A(new_n918), .B(new_n1098), .C1(new_n1106), .C2(new_n734), .ZN(new_n1124));
  INV_X1    g0924(.A(new_n1124), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n1123), .A2(new_n1125), .ZN(new_n1126));
  NAND2_X1  g0926(.A1(new_n1118), .A2(new_n1126), .ZN(new_n1127));
  NOR3_X1   g0927(.A1(new_n458), .A2(new_n680), .A3(new_n846), .ZN(new_n1128));
  NOR3_X1   g0928(.A1(new_n926), .A2(new_n634), .A3(new_n1128), .ZN(new_n1129));
  AOI21_X1  g0929(.A(KEYINPUT116), .B1(new_n1127), .B2(new_n1129), .ZN(new_n1130));
  NAND2_X1  g0930(.A1(new_n1114), .A2(new_n1130), .ZN(new_n1131));
  AOI21_X1  g0931(.A(new_n920), .B1(new_n1108), .B2(new_n1115), .ZN(new_n1132));
  AOI21_X1  g0932(.A(new_n1124), .B1(new_n1122), .B2(new_n921), .ZN(new_n1133));
  OAI21_X1  g0933(.A(new_n1129), .B1(new_n1132), .B2(new_n1133), .ZN(new_n1134));
  INV_X1    g0934(.A(new_n1134), .ZN(new_n1135));
  OAI211_X1 g0935(.A(new_n1110), .B(new_n1113), .C1(new_n1135), .C2(KEYINPUT116), .ZN(new_n1136));
  NAND3_X1  g0936(.A1(new_n1131), .A2(new_n1136), .A3(new_n685), .ZN(new_n1137));
  NAND3_X1  g0937(.A1(new_n1110), .A2(new_n963), .A3(new_n1113), .ZN(new_n1138));
  INV_X1    g0938(.A(new_n835), .ZN(new_n1139));
  INV_X1    g0939(.A(G125), .ZN(new_n1140));
  OAI221_X1 g0940(.A(new_n267), .B1(new_n202), .B2(new_n769), .C1(new_n790), .C2(new_n1140), .ZN(new_n1141));
  XNOR2_X1  g0941(.A(new_n1141), .B(KEYINPUT117), .ZN(new_n1142));
  OR3_X1    g0942(.A1(new_n783), .A2(KEYINPUT53), .A3(new_n1007), .ZN(new_n1143));
  OAI21_X1  g0943(.A(KEYINPUT53), .B1(new_n783), .B2(new_n1007), .ZN(new_n1144));
  OAI211_X1 g0944(.A(new_n1143), .B(new_n1144), .C1(new_n762), .C2(new_n777), .ZN(new_n1145));
  NAND2_X1  g0945(.A1(new_n1053), .A2(G128), .ZN(new_n1146));
  XNOR2_X1  g0946(.A(KEYINPUT54), .B(G143), .ZN(new_n1147));
  OAI221_X1 g0947(.A(new_n1146), .B1(new_n831), .B2(new_n782), .C1(new_n766), .C2(new_n1147), .ZN(new_n1148));
  AOI211_X1 g0948(.A(new_n1145), .B(new_n1148), .C1(G137), .C2(new_n1004), .ZN(new_n1149));
  OAI221_X1 g0949(.A(new_n257), .B1(new_n777), .B2(new_n226), .C1(new_n784), .C2(new_n783), .ZN(new_n1150));
  OAI22_X1  g0950(.A1(new_n775), .A2(new_n816), .B1(new_n782), .B2(new_n464), .ZN(new_n1151));
  NOR2_X1   g0951(.A1(new_n766), .A2(new_n205), .ZN(new_n1152));
  NOR4_X1   g0952(.A1(new_n1150), .A2(new_n827), .A3(new_n1151), .A4(new_n1152), .ZN(new_n1153));
  AOI22_X1  g0953(.A1(new_n791), .A2(G294), .B1(new_n1004), .B2(G107), .ZN(new_n1154));
  AOI22_X1  g0954(.A1(new_n1142), .A2(new_n1149), .B1(new_n1153), .B2(new_n1154), .ZN(new_n1155));
  OAI221_X1 g0955(.A(new_n745), .B1(new_n1072), .B2(new_n1139), .C1(new_n1155), .C2(new_n806), .ZN(new_n1156));
  XOR2_X1   g0956(.A(new_n1156), .B(KEYINPUT118), .Z(new_n1157));
  OAI21_X1  g0957(.A(new_n1157), .B1(new_n915), .B2(new_n747), .ZN(new_n1158));
  AND2_X1   g0958(.A1(new_n1138), .A2(new_n1158), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n1137), .A2(new_n1159), .ZN(G378));
  NAND3_X1  g0960(.A1(new_n895), .A2(new_n899), .A3(G330), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n628), .A2(new_n307), .ZN(new_n1162));
  NAND2_X1  g0962(.A1(new_n299), .A2(new_n859), .ZN(new_n1163));
  XNOR2_X1  g0963(.A(new_n1162), .B(new_n1163), .ZN(new_n1164));
  XOR2_X1   g0964(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1165));
  XNOR2_X1  g0965(.A(new_n1164), .B(new_n1165), .ZN(new_n1166));
  NAND2_X1  g0966(.A1(new_n1161), .A2(new_n1166), .ZN(new_n1167));
  INV_X1    g0967(.A(new_n1166), .ZN(new_n1168));
  NAND4_X1  g0968(.A1(new_n1168), .A2(new_n895), .A3(G330), .A4(new_n899), .ZN(new_n1169));
  NAND2_X1  g0969(.A1(new_n1167), .A2(new_n1169), .ZN(new_n1170));
  NAND2_X1  g0970(.A1(new_n1170), .A2(new_n925), .ZN(new_n1171));
  NAND4_X1  g0971(.A1(new_n1167), .A2(new_n917), .A3(new_n1169), .A4(new_n924), .ZN(new_n1172));
  NAND3_X1  g0972(.A1(new_n1171), .A2(KEYINPUT122), .A3(new_n1172), .ZN(new_n1173));
  INV_X1    g0973(.A(new_n925), .ZN(new_n1174));
  INV_X1    g0974(.A(KEYINPUT122), .ZN(new_n1175));
  NAND4_X1  g0975(.A1(new_n1174), .A2(new_n1175), .A3(new_n1167), .A4(new_n1169), .ZN(new_n1176));
  NAND3_X1  g0976(.A1(new_n1173), .A2(new_n1176), .A3(new_n963), .ZN(new_n1177));
  NOR2_X1   g0977(.A1(new_n267), .A2(G41), .ZN(new_n1178));
  AOI22_X1  g0978(.A1(G97), .A2(new_n821), .B1(new_n822), .B2(G107), .ZN(new_n1179));
  OAI211_X1 g0979(.A(new_n1178), .B(new_n1179), .C1(new_n790), .C2(new_n816), .ZN(new_n1180));
  AOI22_X1  g0980(.A1(new_n1053), .A2(G116), .B1(new_n767), .B2(new_n582), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n770), .A2(G58), .ZN(new_n1182));
  NAND4_X1  g0982(.A1(new_n1181), .A2(new_n1006), .A3(new_n1042), .A4(new_n1182), .ZN(new_n1183));
  NOR2_X1   g0983(.A1(new_n1180), .A2(new_n1183), .ZN(new_n1184));
  XOR2_X1   g0984(.A(new_n1184), .B(KEYINPUT119), .Z(new_n1185));
  INV_X1    g0985(.A(KEYINPUT58), .ZN(new_n1186));
  NAND2_X1  g0986(.A1(new_n1185), .A2(new_n1186), .ZN(new_n1187));
  NOR2_X1   g0987(.A1(G33), .A2(G41), .ZN(new_n1188));
  NOR3_X1   g0988(.A1(new_n1178), .A2(G50), .A3(new_n1188), .ZN(new_n1189));
  OAI22_X1  g0989(.A1(new_n775), .A2(new_n1140), .B1(new_n779), .B2(new_n831), .ZN(new_n1190));
  AOI21_X1  g0990(.A(new_n1190), .B1(G150), .B2(new_n829), .ZN(new_n1191));
  INV_X1    g0991(.A(new_n1147), .ZN(new_n1192));
  AOI22_X1  g0992(.A1(new_n1192), .A2(new_n1000), .B1(new_n822), .B2(G128), .ZN(new_n1193));
  OAI211_X1 g0993(.A(new_n1191), .B(new_n1193), .C1(new_n824), .C2(new_n766), .ZN(new_n1194));
  OR2_X1    g0994(.A1(new_n1194), .A2(KEYINPUT59), .ZN(new_n1195));
  INV_X1    g0995(.A(G124), .ZN(new_n1196));
  OAI221_X1 g0996(.A(new_n1188), .B1(new_n761), .B2(new_n1196), .C1(new_n762), .C2(new_n769), .ZN(new_n1197));
  AOI21_X1  g0997(.A(new_n1197), .B1(new_n1194), .B2(KEYINPUT59), .ZN(new_n1198));
  AOI21_X1  g0998(.A(new_n1189), .B1(new_n1195), .B2(new_n1198), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n1187), .A2(new_n1199), .ZN(new_n1200));
  NOR2_X1   g1000(.A1(new_n1185), .A2(new_n1186), .ZN(new_n1201));
  OAI21_X1  g1001(.A(new_n749), .B1(new_n1200), .B2(new_n1201), .ZN(new_n1202));
  XNOR2_X1  g1002(.A(new_n1202), .B(KEYINPUT120), .ZN(new_n1203));
  AOI21_X1  g1003(.A(new_n742), .B1(new_n202), .B2(new_n835), .ZN(new_n1204));
  OAI211_X1 g1004(.A(new_n1203), .B(new_n1204), .C1(new_n1168), .C2(new_n747), .ZN(new_n1205));
  XOR2_X1   g1005(.A(new_n1205), .B(KEYINPUT121), .Z(new_n1206));
  INV_X1    g1006(.A(new_n1206), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n1177), .A2(new_n1207), .ZN(new_n1208));
  AOI22_X1  g1008(.A1(new_n910), .A2(KEYINPUT39), .B1(new_n912), .B2(new_n913), .ZN(new_n1209));
  AND2_X1   g1009(.A1(new_n880), .A2(new_n884), .ZN(new_n1210));
  AOI22_X1  g1010(.A1(new_n1209), .A2(new_n1095), .B1(new_n1210), .B2(new_n1101), .ZN(new_n1211));
  OAI211_X1 g1011(.A(new_n1113), .B(new_n1127), .C1(new_n1211), .C2(new_n1108), .ZN(new_n1212));
  NAND2_X1  g1012(.A1(new_n1212), .A2(new_n1129), .ZN(new_n1213));
  NAND3_X1  g1013(.A1(new_n1173), .A2(new_n1176), .A3(new_n1213), .ZN(new_n1214));
  INV_X1    g1014(.A(KEYINPUT57), .ZN(new_n1215));
  NAND2_X1  g1015(.A1(new_n1214), .A2(new_n1215), .ZN(new_n1216));
  AOI21_X1  g1016(.A(new_n1215), .B1(new_n1171), .B2(new_n1172), .ZN(new_n1217));
  AOI21_X1  g1017(.A(new_n686), .B1(new_n1217), .B2(new_n1213), .ZN(new_n1218));
  AOI21_X1  g1018(.A(new_n1208), .B1(new_n1216), .B2(new_n1218), .ZN(new_n1219));
  AND2_X1   g1019(.A1(new_n1219), .A2(KEYINPUT123), .ZN(new_n1220));
  NOR2_X1   g1020(.A1(new_n1219), .A2(KEYINPUT123), .ZN(new_n1221));
  NOR2_X1   g1021(.A1(new_n1220), .A2(new_n1221), .ZN(G375));
  NAND2_X1  g1022(.A1(new_n921), .A2(new_n746), .ZN(new_n1223));
  XNOR2_X1  g1023(.A(new_n1223), .B(KEYINPUT124), .ZN(new_n1224));
  INV_X1    g1024(.A(new_n1224), .ZN(new_n1225));
  OAI21_X1  g1025(.A(new_n745), .B1(G68), .B2(new_n1139), .ZN(new_n1226));
  OAI22_X1  g1026(.A1(new_n790), .A2(new_n794), .B1(new_n819), .B2(new_n464), .ZN(new_n1227));
  AOI22_X1  g1027(.A1(G97), .A2(new_n1000), .B1(new_n822), .B2(G283), .ZN(new_n1228));
  OAI221_X1 g1028(.A(new_n1228), .B1(new_n206), .B2(new_n766), .C1(new_n501), .C2(new_n775), .ZN(new_n1229));
  OAI21_X1  g1029(.A(new_n257), .B1(new_n769), .B2(new_n226), .ZN(new_n1230));
  XNOR2_X1  g1030(.A(new_n1230), .B(KEYINPUT125), .ZN(new_n1231));
  OR4_X1    g1031(.A1(new_n1040), .A2(new_n1227), .A3(new_n1229), .A4(new_n1231), .ZN(new_n1232));
  AOI22_X1  g1032(.A1(G132), .A2(new_n1053), .B1(new_n822), .B2(G137), .ZN(new_n1233));
  OAI21_X1  g1033(.A(new_n1233), .B1(new_n819), .B2(new_n1147), .ZN(new_n1234));
  NOR2_X1   g1034(.A1(new_n1234), .A2(KEYINPUT126), .ZN(new_n1235));
  OAI22_X1  g1035(.A1(new_n766), .A2(new_n1007), .B1(new_n783), .B2(new_n762), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n1182), .A2(new_n267), .ZN(new_n1237));
  AOI211_X1 g1037(.A(new_n1236), .B(new_n1237), .C1(G50), .C2(new_n829), .ZN(new_n1238));
  NAND2_X1  g1038(.A1(new_n1234), .A2(KEYINPUT126), .ZN(new_n1239));
  NAND2_X1  g1039(.A1(new_n791), .A2(G128), .ZN(new_n1240));
  NAND3_X1  g1040(.A1(new_n1238), .A2(new_n1239), .A3(new_n1240), .ZN(new_n1241));
  OAI21_X1  g1041(.A(new_n1232), .B1(new_n1235), .B2(new_n1241), .ZN(new_n1242));
  AOI21_X1  g1042(.A(new_n1226), .B1(new_n1242), .B2(new_n749), .ZN(new_n1243));
  AOI22_X1  g1043(.A1(new_n1127), .A2(new_n963), .B1(new_n1225), .B2(new_n1243), .ZN(new_n1244));
  NOR2_X1   g1044(.A1(new_n1127), .A2(new_n1129), .ZN(new_n1245));
  INV_X1    g1045(.A(new_n966), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(new_n1134), .A2(new_n1246), .ZN(new_n1247));
  OAI21_X1  g1047(.A(new_n1244), .B1(new_n1245), .B2(new_n1247), .ZN(G381));
  INV_X1    g1048(.A(G378), .ZN(new_n1249));
  OAI21_X1  g1049(.A(new_n1249), .B1(new_n1220), .B2(new_n1221), .ZN(new_n1250));
  NAND3_X1  g1050(.A1(new_n996), .A2(new_n1023), .A3(new_n1092), .ZN(new_n1251));
  OR2_X1    g1051(.A1(G393), .A2(G396), .ZN(new_n1252));
  OR2_X1    g1052(.A1(new_n1252), .A2(G384), .ZN(new_n1253));
  OR4_X1    g1053(.A1(G381), .A2(new_n1250), .A3(new_n1251), .A4(new_n1253), .ZN(G407));
  OAI211_X1 g1054(.A(G407), .B(G213), .C1(G343), .C2(new_n1250), .ZN(G409));
  NAND2_X1  g1055(.A1(G393), .A2(G396), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(new_n1252), .A2(new_n1256), .ZN(new_n1257));
  INV_X1    g1057(.A(new_n1257), .ZN(new_n1258));
  AND3_X1   g1058(.A1(new_n996), .A2(new_n1023), .A3(new_n1092), .ZN(new_n1259));
  AOI21_X1  g1059(.A(new_n1092), .B1(new_n996), .B2(new_n1023), .ZN(new_n1260));
  OAI21_X1  g1060(.A(new_n1258), .B1(new_n1259), .B2(new_n1260), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(G387), .A2(G390), .ZN(new_n1262));
  NAND3_X1  g1062(.A1(new_n1262), .A2(new_n1251), .A3(new_n1257), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n1261), .A2(new_n1263), .ZN(new_n1264));
  OR4_X1    g1064(.A1(KEYINPUT60), .A2(new_n1129), .A3(new_n1132), .A4(new_n1133), .ZN(new_n1265));
  OAI21_X1  g1065(.A(KEYINPUT60), .B1(new_n1127), .B2(new_n1129), .ZN(new_n1266));
  AND2_X1   g1066(.A1(new_n1265), .A2(new_n1266), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(new_n1134), .A2(new_n685), .ZN(new_n1268));
  OAI211_X1 g1068(.A(G384), .B(new_n1244), .C1(new_n1267), .C2(new_n1268), .ZN(new_n1269));
  AOI21_X1  g1069(.A(new_n1268), .B1(new_n1265), .B2(new_n1266), .ZN(new_n1270));
  INV_X1    g1070(.A(new_n1244), .ZN(new_n1271));
  OAI21_X1  g1071(.A(new_n851), .B1(new_n1270), .B2(new_n1271), .ZN(new_n1272));
  NAND2_X1  g1072(.A1(new_n1269), .A2(new_n1272), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(new_n662), .A2(G213), .ZN(new_n1274));
  INV_X1    g1074(.A(new_n1274), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(new_n1275), .A2(G2897), .ZN(new_n1276));
  XNOR2_X1  g1076(.A(new_n1273), .B(new_n1276), .ZN(new_n1277));
  NAND4_X1  g1077(.A1(new_n1173), .A2(new_n1176), .A3(new_n1213), .A4(new_n1246), .ZN(new_n1278));
  AOI21_X1  g1078(.A(new_n964), .B1(new_n1171), .B2(new_n1172), .ZN(new_n1279));
  NOR2_X1   g1079(.A1(new_n1279), .A2(new_n1206), .ZN(new_n1280));
  AOI21_X1  g1080(.A(G378), .B1(new_n1278), .B2(new_n1280), .ZN(new_n1281));
  AOI21_X1  g1081(.A(new_n1281), .B1(new_n1219), .B2(G378), .ZN(new_n1282));
  OAI21_X1  g1082(.A(new_n1277), .B1(new_n1282), .B2(new_n1275), .ZN(new_n1283));
  NAND2_X1  g1083(.A1(new_n1216), .A2(new_n1218), .ZN(new_n1284));
  INV_X1    g1084(.A(new_n1208), .ZN(new_n1285));
  NAND3_X1  g1085(.A1(new_n1284), .A2(G378), .A3(new_n1285), .ZN(new_n1286));
  NAND2_X1  g1086(.A1(new_n1278), .A2(new_n1280), .ZN(new_n1287));
  NAND2_X1  g1087(.A1(new_n1249), .A2(new_n1287), .ZN(new_n1288));
  NAND2_X1  g1088(.A1(new_n1286), .A2(new_n1288), .ZN(new_n1289));
  INV_X1    g1089(.A(KEYINPUT62), .ZN(new_n1290));
  INV_X1    g1090(.A(new_n1273), .ZN(new_n1291));
  NAND4_X1  g1091(.A1(new_n1289), .A2(new_n1290), .A3(new_n1274), .A4(new_n1291), .ZN(new_n1292));
  INV_X1    g1092(.A(KEYINPUT61), .ZN(new_n1293));
  NAND3_X1  g1093(.A1(new_n1283), .A2(new_n1292), .A3(new_n1293), .ZN(new_n1294));
  AOI211_X1 g1094(.A(new_n1275), .B(new_n1273), .C1(new_n1286), .C2(new_n1288), .ZN(new_n1295));
  NOR2_X1   g1095(.A1(new_n1295), .A2(new_n1290), .ZN(new_n1296));
  OAI21_X1  g1096(.A(new_n1264), .B1(new_n1294), .B2(new_n1296), .ZN(new_n1297));
  AOI21_X1  g1097(.A(new_n1275), .B1(new_n1286), .B2(new_n1288), .ZN(new_n1298));
  NAND2_X1  g1098(.A1(new_n1298), .A2(new_n1291), .ZN(new_n1299));
  INV_X1    g1099(.A(new_n1276), .ZN(new_n1300));
  XNOR2_X1  g1100(.A(new_n1273), .B(new_n1300), .ZN(new_n1301));
  NOR2_X1   g1101(.A1(new_n1298), .A2(new_n1301), .ZN(new_n1302));
  INV_X1    g1102(.A(KEYINPUT63), .ZN(new_n1303));
  OAI21_X1  g1103(.A(new_n1299), .B1(new_n1302), .B2(new_n1303), .ZN(new_n1304));
  NAND3_X1  g1104(.A1(new_n1261), .A2(new_n1263), .A3(new_n1293), .ZN(new_n1305));
  AOI21_X1  g1105(.A(new_n1305), .B1(new_n1295), .B2(KEYINPUT63), .ZN(new_n1306));
  NAND2_X1  g1106(.A1(new_n1304), .A2(new_n1306), .ZN(new_n1307));
  NAND2_X1  g1107(.A1(new_n1297), .A2(new_n1307), .ZN(new_n1308));
  NAND2_X1  g1108(.A1(new_n1308), .A2(KEYINPUT127), .ZN(new_n1309));
  INV_X1    g1109(.A(KEYINPUT127), .ZN(new_n1310));
  NAND3_X1  g1110(.A1(new_n1297), .A2(new_n1307), .A3(new_n1310), .ZN(new_n1311));
  NAND2_X1  g1111(.A1(new_n1309), .A2(new_n1311), .ZN(G405));
  XNOR2_X1  g1112(.A(new_n1264), .B(new_n1273), .ZN(new_n1313));
  OAI21_X1  g1113(.A(new_n1250), .B1(new_n1249), .B2(new_n1219), .ZN(new_n1314));
  XNOR2_X1  g1114(.A(new_n1313), .B(new_n1314), .ZN(G402));
endmodule


