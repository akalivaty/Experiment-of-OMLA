//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 1 0 0 1 0 0 0 1 0 1 1 1 0 1 1 1 1 0 1 1 0 0 0 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 0 0 1 0 1 1 0 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:19:47 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n690, new_n691, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n711, new_n712, new_n713, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n748, new_n749,
    new_n750, new_n751, new_n752, new_n753, new_n755, new_n756, new_n757,
    new_n758, new_n759, new_n760, new_n762, new_n764, new_n765, new_n766,
    new_n767, new_n768, new_n769, new_n770, new_n771, new_n772, new_n773,
    new_n774, new_n775, new_n776, new_n777, new_n778, new_n779, new_n780,
    new_n781, new_n782, new_n783, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n802, new_n803,
    new_n804, new_n805, new_n806, new_n807, new_n808, new_n809, new_n810,
    new_n811, new_n812, new_n813, new_n814, new_n815, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n870, new_n871, new_n873, new_n874, new_n876, new_n877, new_n878,
    new_n879, new_n880, new_n881, new_n882, new_n883, new_n884, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n924, new_n925, new_n926, new_n927, new_n929, new_n930, new_n931,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n940,
    new_n941, new_n942, new_n943, new_n945, new_n946, new_n947, new_n949,
    new_n950, new_n951, new_n952, new_n954, new_n955, new_n956, new_n957,
    new_n958, new_n959, new_n960, new_n961, new_n962, new_n963, new_n964,
    new_n966, new_n967, new_n968, new_n969, new_n971, new_n972, new_n973,
    new_n974, new_n975, new_n976, new_n977, new_n978, new_n979, new_n980,
    new_n981, new_n982, new_n983, new_n984, new_n985, new_n986, new_n988,
    new_n989;
  NAND2_X1  g000(.A1(G183gat), .A2(G190gat), .ZN(new_n202));
  OAI21_X1  g001(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n203));
  INV_X1    g002(.A(KEYINPUT66), .ZN(new_n204));
  AOI21_X1  g003(.A(new_n204), .B1(G169gat), .B2(G176gat), .ZN(new_n205));
  NAND2_X1  g004(.A1(G169gat), .A2(G176gat), .ZN(new_n206));
  NOR2_X1   g005(.A1(new_n206), .A2(KEYINPUT66), .ZN(new_n207));
  OAI21_X1  g006(.A(new_n203), .B1(new_n205), .B2(new_n207), .ZN(new_n208));
  INV_X1    g007(.A(KEYINPUT67), .ZN(new_n209));
  INV_X1    g008(.A(G169gat), .ZN(new_n210));
  INV_X1    g009(.A(G176gat), .ZN(new_n211));
  NAND3_X1  g010(.A1(new_n209), .A2(new_n210), .A3(new_n211), .ZN(new_n212));
  OAI21_X1  g011(.A(KEYINPUT67), .B1(G169gat), .B2(G176gat), .ZN(new_n213));
  AOI21_X1  g012(.A(KEYINPUT26), .B1(new_n212), .B2(new_n213), .ZN(new_n214));
  OAI21_X1  g013(.A(new_n202), .B1(new_n208), .B2(new_n214), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n215), .A2(KEYINPUT69), .ZN(new_n216));
  INV_X1    g015(.A(KEYINPUT28), .ZN(new_n217));
  INV_X1    g016(.A(KEYINPUT27), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n218), .A2(G183gat), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n219), .A2(KEYINPUT68), .ZN(new_n220));
  INV_X1    g019(.A(G190gat), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  INV_X1    g021(.A(G183gat), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n223), .A2(KEYINPUT27), .ZN(new_n224));
  AOI21_X1  g023(.A(KEYINPUT68), .B1(new_n219), .B2(new_n224), .ZN(new_n225));
  OAI21_X1  g024(.A(new_n217), .B1(new_n222), .B2(new_n225), .ZN(new_n226));
  AND2_X1   g025(.A1(new_n219), .A2(new_n224), .ZN(new_n227));
  NAND3_X1  g026(.A1(new_n227), .A2(KEYINPUT28), .A3(new_n221), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n226), .A2(new_n228), .ZN(new_n229));
  INV_X1    g028(.A(KEYINPUT69), .ZN(new_n230));
  OAI211_X1 g029(.A(new_n230), .B(new_n202), .C1(new_n208), .C2(new_n214), .ZN(new_n231));
  NAND3_X1  g030(.A1(new_n216), .A2(new_n229), .A3(new_n231), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n223), .A2(new_n221), .ZN(new_n233));
  NAND3_X1  g032(.A1(new_n233), .A2(KEYINPUT24), .A3(new_n202), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n206), .A2(KEYINPUT66), .ZN(new_n235));
  NAND3_X1  g034(.A1(new_n204), .A2(G169gat), .A3(G176gat), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n235), .A2(new_n236), .ZN(new_n237));
  OR2_X1    g036(.A1(new_n202), .A2(KEYINPUT24), .ZN(new_n238));
  AND3_X1   g037(.A1(new_n234), .A2(new_n237), .A3(new_n238), .ZN(new_n239));
  INV_X1    g038(.A(KEYINPUT23), .ZN(new_n240));
  OAI21_X1  g039(.A(new_n240), .B1(G169gat), .B2(G176gat), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n212), .A2(new_n213), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n242), .A2(KEYINPUT23), .ZN(new_n243));
  NAND4_X1  g042(.A1(new_n239), .A2(KEYINPUT25), .A3(new_n241), .A4(new_n243), .ZN(new_n244));
  INV_X1    g043(.A(KEYINPUT25), .ZN(new_n245));
  NAND4_X1  g044(.A1(new_n234), .A2(new_n237), .A3(new_n241), .A4(new_n238), .ZN(new_n246));
  XNOR2_X1  g045(.A(KEYINPUT64), .B(G169gat), .ZN(new_n247));
  XNOR2_X1  g046(.A(KEYINPUT65), .B(G176gat), .ZN(new_n248));
  AND3_X1   g047(.A1(new_n247), .A2(new_n248), .A3(KEYINPUT23), .ZN(new_n249));
  OAI21_X1  g048(.A(new_n245), .B1(new_n246), .B2(new_n249), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n244), .A2(new_n250), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n232), .A2(new_n251), .ZN(new_n252));
  INV_X1    g051(.A(G113gat), .ZN(new_n253));
  INV_X1    g052(.A(G120gat), .ZN(new_n254));
  AOI21_X1  g053(.A(KEYINPUT1), .B1(new_n253), .B2(new_n254), .ZN(new_n255));
  OAI21_X1  g054(.A(new_n255), .B1(new_n253), .B2(new_n254), .ZN(new_n256));
  INV_X1    g055(.A(G127gat), .ZN(new_n257));
  INV_X1    g056(.A(G134gat), .ZN(new_n258));
  NAND2_X1  g057(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  NAND2_X1  g058(.A1(G127gat), .A2(G134gat), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  AND2_X1   g060(.A1(new_n261), .A2(KEYINPUT70), .ZN(new_n262));
  NOR2_X1   g061(.A1(new_n261), .A2(KEYINPUT70), .ZN(new_n263));
  OAI21_X1  g062(.A(new_n256), .B1(new_n262), .B2(new_n263), .ZN(new_n264));
  XOR2_X1   g063(.A(KEYINPUT71), .B(G120gat), .Z(new_n265));
  NAND2_X1  g064(.A1(new_n265), .A2(G113gat), .ZN(new_n266));
  NAND3_X1  g065(.A1(new_n266), .A2(new_n261), .A3(new_n255), .ZN(new_n267));
  NAND2_X1  g066(.A1(new_n264), .A2(new_n267), .ZN(new_n268));
  INV_X1    g067(.A(new_n268), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n252), .A2(new_n269), .ZN(new_n270));
  NAND3_X1  g069(.A1(new_n232), .A2(new_n268), .A3(new_n251), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  INV_X1    g071(.A(KEYINPUT34), .ZN(new_n273));
  INV_X1    g072(.A(G227gat), .ZN(new_n274));
  INV_X1    g073(.A(G233gat), .ZN(new_n275));
  NOR2_X1   g074(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  INV_X1    g075(.A(new_n276), .ZN(new_n277));
  NAND3_X1  g076(.A1(new_n272), .A2(new_n273), .A3(new_n277), .ZN(new_n278));
  INV_X1    g077(.A(new_n278), .ZN(new_n279));
  AOI21_X1  g078(.A(new_n273), .B1(new_n272), .B2(new_n277), .ZN(new_n280));
  NOR2_X1   g079(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  NAND3_X1  g080(.A1(new_n270), .A2(new_n276), .A3(new_n271), .ZN(new_n282));
  XNOR2_X1  g081(.A(G15gat), .B(G43gat), .ZN(new_n283));
  XNOR2_X1  g082(.A(new_n283), .B(G71gat), .ZN(new_n284));
  INV_X1    g083(.A(G99gat), .ZN(new_n285));
  XNOR2_X1  g084(.A(new_n284), .B(new_n285), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n286), .A2(KEYINPUT33), .ZN(new_n287));
  NAND3_X1  g086(.A1(new_n282), .A2(KEYINPUT32), .A3(new_n287), .ZN(new_n288));
  NAND2_X1  g087(.A1(new_n288), .A2(KEYINPUT73), .ZN(new_n289));
  INV_X1    g088(.A(KEYINPUT73), .ZN(new_n290));
  NAND4_X1  g089(.A1(new_n282), .A2(new_n290), .A3(KEYINPUT32), .A4(new_n287), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n289), .A2(new_n291), .ZN(new_n292));
  AND3_X1   g091(.A1(new_n232), .A2(new_n268), .A3(new_n251), .ZN(new_n293));
  AOI21_X1  g092(.A(new_n268), .B1(new_n232), .B2(new_n251), .ZN(new_n294));
  NOR3_X1   g093(.A1(new_n293), .A2(new_n294), .A3(new_n277), .ZN(new_n295));
  INV_X1    g094(.A(KEYINPUT33), .ZN(new_n296));
  NOR2_X1   g095(.A1(new_n296), .A2(KEYINPUT32), .ZN(new_n297));
  OAI21_X1  g096(.A(new_n286), .B1(new_n295), .B2(new_n297), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n298), .A2(KEYINPUT72), .ZN(new_n299));
  INV_X1    g098(.A(new_n297), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n282), .A2(new_n300), .ZN(new_n301));
  INV_X1    g100(.A(KEYINPUT72), .ZN(new_n302));
  NAND3_X1  g101(.A1(new_n301), .A2(new_n302), .A3(new_n286), .ZN(new_n303));
  AND4_X1   g102(.A1(new_n281), .A2(new_n292), .A3(new_n299), .A4(new_n303), .ZN(new_n304));
  AOI21_X1  g103(.A(new_n302), .B1(new_n301), .B2(new_n286), .ZN(new_n305));
  INV_X1    g104(.A(new_n286), .ZN(new_n306));
  AOI211_X1 g105(.A(KEYINPUT72), .B(new_n306), .C1(new_n282), .C2(new_n300), .ZN(new_n307));
  NOR2_X1   g106(.A1(new_n305), .A2(new_n307), .ZN(new_n308));
  AOI21_X1  g107(.A(new_n281), .B1(new_n308), .B2(new_n292), .ZN(new_n309));
  NOR2_X1   g108(.A1(new_n304), .A2(new_n309), .ZN(new_n310));
  XNOR2_X1  g109(.A(G78gat), .B(G106gat), .ZN(new_n311));
  INV_X1    g110(.A(G50gat), .ZN(new_n312));
  XNOR2_X1  g111(.A(new_n311), .B(new_n312), .ZN(new_n313));
  XNOR2_X1  g112(.A(new_n313), .B(KEYINPUT81), .ZN(new_n314));
  XNOR2_X1  g113(.A(new_n314), .B(KEYINPUT31), .ZN(new_n315));
  INV_X1    g114(.A(KEYINPUT84), .ZN(new_n316));
  NOR2_X1   g115(.A1(new_n315), .A2(new_n316), .ZN(new_n317));
  INV_X1    g116(.A(G228gat), .ZN(new_n318));
  NOR2_X1   g117(.A1(new_n318), .A2(new_n275), .ZN(new_n319));
  INV_X1    g118(.A(new_n319), .ZN(new_n320));
  XOR2_X1   g119(.A(G155gat), .B(G162gat), .Z(new_n321));
  XNOR2_X1  g120(.A(G141gat), .B(G148gat), .ZN(new_n322));
  OAI21_X1  g121(.A(new_n321), .B1(KEYINPUT2), .B2(new_n322), .ZN(new_n323));
  INV_X1    g122(.A(new_n323), .ZN(new_n324));
  INV_X1    g123(.A(KEYINPUT2), .ZN(new_n325));
  XNOR2_X1  g124(.A(KEYINPUT77), .B(G162gat), .ZN(new_n326));
  AOI21_X1  g125(.A(new_n325), .B1(new_n326), .B2(G155gat), .ZN(new_n327));
  INV_X1    g126(.A(KEYINPUT78), .ZN(new_n328));
  AOI21_X1  g127(.A(new_n321), .B1(new_n327), .B2(new_n328), .ZN(new_n329));
  INV_X1    g128(.A(G162gat), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n330), .A2(KEYINPUT77), .ZN(new_n331));
  INV_X1    g130(.A(KEYINPUT77), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n332), .A2(G162gat), .ZN(new_n333));
  NAND3_X1  g132(.A1(new_n331), .A2(new_n333), .A3(G155gat), .ZN(new_n334));
  NAND2_X1  g133(.A1(new_n334), .A2(KEYINPUT2), .ZN(new_n335));
  AOI21_X1  g134(.A(new_n322), .B1(new_n335), .B2(KEYINPUT78), .ZN(new_n336));
  AOI21_X1  g135(.A(new_n324), .B1(new_n329), .B2(new_n336), .ZN(new_n337));
  INV_X1    g136(.A(KEYINPUT29), .ZN(new_n338));
  XNOR2_X1  g137(.A(KEYINPUT76), .B(G211gat), .ZN(new_n339));
  AOI21_X1  g138(.A(KEYINPUT22), .B1(new_n339), .B2(G218gat), .ZN(new_n340));
  INV_X1    g139(.A(G197gat), .ZN(new_n341));
  AND2_X1   g140(.A1(KEYINPUT75), .A2(G204gat), .ZN(new_n342));
  NOR2_X1   g141(.A1(KEYINPUT75), .A2(G204gat), .ZN(new_n343));
  OAI21_X1  g142(.A(new_n341), .B1(new_n342), .B2(new_n343), .ZN(new_n344));
  INV_X1    g143(.A(KEYINPUT75), .ZN(new_n345));
  INV_X1    g144(.A(G204gat), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n345), .A2(new_n346), .ZN(new_n347));
  NAND2_X1  g146(.A1(KEYINPUT75), .A2(G204gat), .ZN(new_n348));
  NAND3_X1  g147(.A1(new_n347), .A2(G197gat), .A3(new_n348), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n344), .A2(new_n349), .ZN(new_n350));
  OAI21_X1  g149(.A(G211gat), .B1(new_n340), .B2(new_n350), .ZN(new_n351));
  INV_X1    g150(.A(G211gat), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n352), .A2(KEYINPUT76), .ZN(new_n353));
  INV_X1    g152(.A(KEYINPUT76), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n354), .A2(G211gat), .ZN(new_n355));
  NAND3_X1  g154(.A1(new_n353), .A2(new_n355), .A3(G218gat), .ZN(new_n356));
  INV_X1    g155(.A(KEYINPUT22), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  NAND4_X1  g157(.A1(new_n358), .A2(new_n352), .A3(new_n349), .A4(new_n344), .ZN(new_n359));
  AND3_X1   g158(.A1(new_n351), .A2(G218gat), .A3(new_n359), .ZN(new_n360));
  AOI21_X1  g159(.A(G218gat), .B1(new_n351), .B2(new_n359), .ZN(new_n361));
  OAI21_X1  g160(.A(new_n338), .B1(new_n360), .B2(new_n361), .ZN(new_n362));
  INV_X1    g161(.A(KEYINPUT3), .ZN(new_n363));
  AOI21_X1  g162(.A(new_n337), .B1(new_n362), .B2(new_n363), .ZN(new_n364));
  INV_X1    g163(.A(new_n361), .ZN(new_n365));
  NAND3_X1  g164(.A1(new_n351), .A2(G218gat), .A3(new_n359), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n365), .A2(new_n366), .ZN(new_n367));
  AOI21_X1  g166(.A(KEYINPUT29), .B1(new_n337), .B2(new_n363), .ZN(new_n368));
  NOR2_X1   g167(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  OAI21_X1  g168(.A(new_n320), .B1(new_n364), .B2(new_n369), .ZN(new_n370));
  INV_X1    g169(.A(KEYINPUT82), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  OAI211_X1 g171(.A(KEYINPUT82), .B(new_n320), .C1(new_n364), .C2(new_n369), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n362), .A2(new_n363), .ZN(new_n374));
  INV_X1    g173(.A(new_n322), .ZN(new_n375));
  OAI21_X1  g174(.A(new_n375), .B1(new_n327), .B2(new_n328), .ZN(new_n376));
  INV_X1    g175(.A(new_n321), .ZN(new_n377));
  OAI21_X1  g176(.A(new_n377), .B1(new_n335), .B2(KEYINPUT78), .ZN(new_n378));
  OAI21_X1  g177(.A(new_n323), .B1(new_n376), .B2(new_n378), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n374), .A2(new_n379), .ZN(new_n380));
  NOR2_X1   g179(.A1(new_n360), .A2(new_n361), .ZN(new_n381));
  OAI211_X1 g180(.A(new_n363), .B(new_n323), .C1(new_n376), .C2(new_n378), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n382), .A2(new_n338), .ZN(new_n383));
  AOI21_X1  g182(.A(KEYINPUT83), .B1(new_n381), .B2(new_n383), .ZN(new_n384));
  AND3_X1   g183(.A1(new_n381), .A2(KEYINPUT83), .A3(new_n383), .ZN(new_n385));
  OAI211_X1 g184(.A(new_n380), .B(new_n319), .C1(new_n384), .C2(new_n385), .ZN(new_n386));
  NAND3_X1  g185(.A1(new_n372), .A2(new_n373), .A3(new_n386), .ZN(new_n387));
  NAND3_X1  g186(.A1(new_n387), .A2(G22gat), .A3(new_n315), .ZN(new_n388));
  INV_X1    g187(.A(G22gat), .ZN(new_n389));
  NAND4_X1  g188(.A1(new_n372), .A2(new_n389), .A3(new_n386), .A4(new_n373), .ZN(new_n390));
  AOI21_X1  g189(.A(new_n317), .B1(new_n388), .B2(new_n390), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n387), .A2(G22gat), .ZN(new_n392));
  AND3_X1   g191(.A1(new_n392), .A2(new_n317), .A3(new_n390), .ZN(new_n393));
  OAI21_X1  g192(.A(new_n310), .B1(new_n391), .B2(new_n393), .ZN(new_n394));
  XNOR2_X1  g193(.A(G1gat), .B(G29gat), .ZN(new_n395));
  XNOR2_X1  g194(.A(new_n395), .B(KEYINPUT0), .ZN(new_n396));
  XNOR2_X1  g195(.A(new_n396), .B(G57gat), .ZN(new_n397));
  INV_X1    g196(.A(G85gat), .ZN(new_n398));
  XNOR2_X1  g197(.A(new_n397), .B(new_n398), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n379), .A2(KEYINPUT3), .ZN(new_n400));
  NAND3_X1  g199(.A1(new_n400), .A2(new_n268), .A3(new_n382), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n401), .A2(KEYINPUT79), .ZN(new_n402));
  INV_X1    g201(.A(KEYINPUT79), .ZN(new_n403));
  NAND4_X1  g202(.A1(new_n400), .A2(new_n403), .A3(new_n268), .A4(new_n382), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n402), .A2(new_n404), .ZN(new_n405));
  NAND2_X1  g204(.A1(G225gat), .A2(G233gat), .ZN(new_n406));
  INV_X1    g205(.A(KEYINPUT4), .ZN(new_n407));
  NAND3_X1  g206(.A1(new_n269), .A2(new_n407), .A3(new_n337), .ZN(new_n408));
  OAI21_X1  g207(.A(KEYINPUT4), .B1(new_n379), .B2(new_n268), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n408), .A2(new_n409), .ZN(new_n410));
  AND4_X1   g209(.A1(KEYINPUT5), .A2(new_n405), .A3(new_n406), .A4(new_n410), .ZN(new_n411));
  INV_X1    g210(.A(KEYINPUT5), .ZN(new_n412));
  XNOR2_X1  g211(.A(new_n379), .B(new_n268), .ZN(new_n413));
  INV_X1    g212(.A(new_n406), .ZN(new_n414));
  AOI21_X1  g213(.A(new_n412), .B1(new_n413), .B2(new_n414), .ZN(new_n415));
  AOI22_X1  g214(.A1(new_n402), .A2(new_n404), .B1(new_n409), .B2(new_n408), .ZN(new_n416));
  AOI21_X1  g215(.A(new_n415), .B1(new_n416), .B2(new_n406), .ZN(new_n417));
  OAI21_X1  g216(.A(new_n399), .B1(new_n411), .B2(new_n417), .ZN(new_n418));
  NAND3_X1  g217(.A1(new_n405), .A2(new_n406), .A3(new_n410), .ZN(new_n419));
  INV_X1    g218(.A(new_n415), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  INV_X1    g220(.A(new_n399), .ZN(new_n422));
  NAND3_X1  g221(.A1(new_n416), .A2(KEYINPUT5), .A3(new_n406), .ZN(new_n423));
  NAND3_X1  g222(.A1(new_n421), .A2(new_n422), .A3(new_n423), .ZN(new_n424));
  INV_X1    g223(.A(KEYINPUT6), .ZN(new_n425));
  NAND4_X1  g224(.A1(new_n418), .A2(KEYINPUT80), .A3(new_n424), .A4(new_n425), .ZN(new_n426));
  NOR2_X1   g225(.A1(new_n411), .A2(new_n417), .ZN(new_n427));
  INV_X1    g226(.A(KEYINPUT80), .ZN(new_n428));
  OAI211_X1 g227(.A(new_n427), .B(new_n422), .C1(new_n428), .C2(KEYINPUT6), .ZN(new_n429));
  NAND2_X1  g228(.A1(new_n426), .A2(new_n429), .ZN(new_n430));
  NAND2_X1  g229(.A1(G226gat), .A2(G233gat), .ZN(new_n431));
  INV_X1    g230(.A(new_n431), .ZN(new_n432));
  AOI211_X1 g231(.A(KEYINPUT29), .B(new_n432), .C1(new_n232), .C2(new_n251), .ZN(new_n433));
  AND3_X1   g232(.A1(new_n232), .A2(new_n432), .A3(new_n251), .ZN(new_n434));
  OAI21_X1  g233(.A(new_n381), .B1(new_n433), .B2(new_n434), .ZN(new_n435));
  NAND3_X1  g234(.A1(new_n252), .A2(new_n338), .A3(new_n431), .ZN(new_n436));
  NAND3_X1  g235(.A1(new_n232), .A2(new_n432), .A3(new_n251), .ZN(new_n437));
  NAND3_X1  g236(.A1(new_n436), .A2(new_n367), .A3(new_n437), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n435), .A2(new_n438), .ZN(new_n439));
  XNOR2_X1  g238(.A(G8gat), .B(G36gat), .ZN(new_n440));
  INV_X1    g239(.A(G64gat), .ZN(new_n441));
  XNOR2_X1  g240(.A(new_n440), .B(new_n441), .ZN(new_n442));
  XOR2_X1   g241(.A(new_n442), .B(G92gat), .Z(new_n443));
  INV_X1    g242(.A(new_n443), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n439), .A2(new_n444), .ZN(new_n445));
  NAND3_X1  g244(.A1(new_n435), .A2(new_n438), .A3(new_n443), .ZN(new_n446));
  NAND3_X1  g245(.A1(new_n445), .A2(KEYINPUT30), .A3(new_n446), .ZN(new_n447));
  INV_X1    g246(.A(KEYINPUT30), .ZN(new_n448));
  NAND3_X1  g247(.A1(new_n439), .A2(new_n448), .A3(new_n444), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n447), .A2(new_n449), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n430), .A2(new_n450), .ZN(new_n451));
  OAI21_X1  g250(.A(KEYINPUT35), .B1(new_n394), .B2(new_n451), .ZN(new_n452));
  INV_X1    g251(.A(new_n281), .ZN(new_n453));
  INV_X1    g252(.A(new_n292), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n299), .A2(new_n303), .ZN(new_n455));
  OAI21_X1  g254(.A(new_n453), .B1(new_n454), .B2(new_n455), .ZN(new_n456));
  INV_X1    g255(.A(KEYINPUT74), .ZN(new_n457));
  NAND3_X1  g256(.A1(new_n308), .A2(new_n281), .A3(new_n292), .ZN(new_n458));
  NAND3_X1  g257(.A1(new_n456), .A2(new_n457), .A3(new_n458), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n309), .A2(KEYINPUT74), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n388), .A2(new_n390), .ZN(new_n462));
  INV_X1    g261(.A(new_n317), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  NAND3_X1  g263(.A1(new_n392), .A2(new_n317), .A3(new_n390), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  NAND3_X1  g265(.A1(new_n418), .A2(new_n425), .A3(new_n424), .ZN(new_n467));
  NAND3_X1  g266(.A1(new_n427), .A2(KEYINPUT6), .A3(new_n422), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  INV_X1    g268(.A(new_n450), .ZN(new_n470));
  NOR2_X1   g269(.A1(new_n470), .A2(KEYINPUT35), .ZN(new_n471));
  NAND4_X1  g270(.A1(new_n461), .A2(new_n466), .A3(new_n469), .A4(new_n471), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n452), .A2(new_n472), .ZN(new_n473));
  INV_X1    g272(.A(KEYINPUT36), .ZN(new_n474));
  AOI21_X1  g273(.A(new_n474), .B1(new_n456), .B2(new_n458), .ZN(new_n475));
  AOI21_X1  g274(.A(new_n475), .B1(new_n461), .B2(new_n474), .ZN(new_n476));
  INV_X1    g275(.A(new_n445), .ZN(new_n477));
  NAND3_X1  g276(.A1(new_n435), .A2(KEYINPUT37), .A3(new_n438), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n478), .A2(new_n443), .ZN(new_n479));
  INV_X1    g278(.A(KEYINPUT37), .ZN(new_n480));
  NOR3_X1   g279(.A1(new_n433), .A2(new_n381), .A3(new_n434), .ZN(new_n481));
  AOI21_X1  g280(.A(new_n367), .B1(new_n436), .B2(new_n437), .ZN(new_n482));
  OAI21_X1  g281(.A(new_n480), .B1(new_n481), .B2(new_n482), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n483), .A2(KEYINPUT85), .ZN(new_n484));
  INV_X1    g283(.A(KEYINPUT85), .ZN(new_n485));
  NAND3_X1  g284(.A1(new_n439), .A2(new_n485), .A3(new_n480), .ZN(new_n486));
  AOI21_X1  g285(.A(new_n479), .B1(new_n484), .B2(new_n486), .ZN(new_n487));
  INV_X1    g286(.A(KEYINPUT38), .ZN(new_n488));
  AOI21_X1  g287(.A(new_n477), .B1(new_n487), .B2(new_n488), .ZN(new_n489));
  INV_X1    g288(.A(new_n479), .ZN(new_n490));
  INV_X1    g289(.A(new_n486), .ZN(new_n491));
  AOI21_X1  g290(.A(new_n485), .B1(new_n439), .B2(new_n480), .ZN(new_n492));
  OAI21_X1  g291(.A(new_n490), .B1(new_n491), .B2(new_n492), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n493), .A2(KEYINPUT38), .ZN(new_n494));
  NAND4_X1  g293(.A1(new_n489), .A2(new_n494), .A3(new_n467), .A4(new_n468), .ZN(new_n495));
  OR3_X1    g294(.A1(new_n416), .A2(KEYINPUT39), .A3(new_n406), .ZN(new_n496));
  OR2_X1    g295(.A1(new_n413), .A2(new_n414), .ZN(new_n497));
  OAI211_X1 g296(.A(KEYINPUT39), .B(new_n497), .C1(new_n416), .C2(new_n406), .ZN(new_n498));
  NAND3_X1  g297(.A1(new_n496), .A2(new_n399), .A3(new_n498), .ZN(new_n499));
  INV_X1    g298(.A(KEYINPUT40), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  NAND4_X1  g300(.A1(new_n496), .A2(KEYINPUT40), .A3(new_n399), .A4(new_n498), .ZN(new_n502));
  NAND4_X1  g301(.A1(new_n501), .A2(new_n470), .A3(new_n424), .A4(new_n502), .ZN(new_n503));
  NAND3_X1  g302(.A1(new_n495), .A2(new_n466), .A3(new_n503), .ZN(new_n504));
  NOR2_X1   g303(.A1(new_n393), .A2(new_n391), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n451), .A2(new_n505), .ZN(new_n506));
  NAND3_X1  g305(.A1(new_n476), .A2(new_n504), .A3(new_n506), .ZN(new_n507));
  INV_X1    g306(.A(KEYINPUT86), .ZN(new_n508));
  AND3_X1   g307(.A1(new_n473), .A2(new_n507), .A3(new_n508), .ZN(new_n509));
  AOI21_X1  g308(.A(new_n508), .B1(new_n473), .B2(new_n507), .ZN(new_n510));
  INV_X1    g309(.A(KEYINPUT92), .ZN(new_n511));
  INV_X1    g310(.A(KEYINPUT14), .ZN(new_n512));
  OAI21_X1  g311(.A(new_n512), .B1(G29gat), .B2(G36gat), .ZN(new_n513));
  INV_X1    g312(.A(G29gat), .ZN(new_n514));
  INV_X1    g313(.A(G36gat), .ZN(new_n515));
  NAND3_X1  g314(.A1(new_n514), .A2(new_n515), .A3(KEYINPUT14), .ZN(new_n516));
  XNOR2_X1  g315(.A(KEYINPUT88), .B(G36gat), .ZN(new_n517));
  OAI211_X1 g316(.A(new_n513), .B(new_n516), .C1(new_n517), .C2(new_n514), .ZN(new_n518));
  INV_X1    g317(.A(KEYINPUT15), .ZN(new_n519));
  XNOR2_X1  g318(.A(new_n518), .B(new_n519), .ZN(new_n520));
  XNOR2_X1  g319(.A(G43gat), .B(G50gat), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  INV_X1    g321(.A(new_n521), .ZN(new_n523));
  OAI21_X1  g322(.A(new_n523), .B1(new_n518), .B2(new_n519), .ZN(new_n524));
  AND2_X1   g323(.A1(new_n522), .A2(new_n524), .ZN(new_n525));
  XNOR2_X1  g324(.A(G15gat), .B(G22gat), .ZN(new_n526));
  OR2_X1    g325(.A1(new_n526), .A2(G1gat), .ZN(new_n527));
  INV_X1    g326(.A(KEYINPUT16), .ZN(new_n528));
  OAI21_X1  g327(.A(new_n526), .B1(new_n528), .B2(G1gat), .ZN(new_n529));
  INV_X1    g328(.A(G8gat), .ZN(new_n530));
  NAND3_X1  g329(.A1(new_n527), .A2(new_n529), .A3(new_n530), .ZN(new_n531));
  INV_X1    g330(.A(KEYINPUT90), .ZN(new_n532));
  XNOR2_X1  g331(.A(new_n531), .B(new_n532), .ZN(new_n533));
  NAND3_X1  g332(.A1(new_n527), .A2(new_n529), .A3(KEYINPUT89), .ZN(new_n534));
  OAI211_X1 g333(.A(new_n534), .B(G8gat), .C1(KEYINPUT89), .C2(new_n527), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n533), .A2(new_n535), .ZN(new_n536));
  NAND3_X1  g335(.A1(new_n525), .A2(KEYINPUT91), .A3(new_n536), .ZN(new_n537));
  INV_X1    g336(.A(new_n537), .ZN(new_n538));
  AOI21_X1  g337(.A(KEYINPUT91), .B1(new_n525), .B2(new_n536), .ZN(new_n539));
  OAI21_X1  g338(.A(new_n511), .B1(new_n538), .B2(new_n539), .ZN(new_n540));
  INV_X1    g339(.A(new_n539), .ZN(new_n541));
  NAND3_X1  g340(.A1(new_n541), .A2(KEYINPUT92), .A3(new_n537), .ZN(new_n542));
  INV_X1    g341(.A(new_n536), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n522), .A2(new_n524), .ZN(new_n544));
  NAND2_X1  g343(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  NAND3_X1  g344(.A1(new_n540), .A2(new_n542), .A3(new_n545), .ZN(new_n546));
  NAND2_X1  g345(.A1(G229gat), .A2(G233gat), .ZN(new_n547));
  XOR2_X1   g346(.A(new_n547), .B(KEYINPUT13), .Z(new_n548));
  NAND2_X1  g347(.A1(new_n546), .A2(new_n548), .ZN(new_n549));
  INV_X1    g348(.A(KEYINPUT17), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n525), .A2(new_n550), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n544), .A2(KEYINPUT17), .ZN(new_n552));
  NAND3_X1  g351(.A1(new_n551), .A2(new_n552), .A3(new_n543), .ZN(new_n553));
  OAI211_X1 g352(.A(new_n553), .B(new_n547), .C1(new_n538), .C2(new_n539), .ZN(new_n554));
  INV_X1    g353(.A(new_n554), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n555), .A2(KEYINPUT18), .ZN(new_n556));
  XNOR2_X1  g355(.A(G113gat), .B(G141gat), .ZN(new_n557));
  XNOR2_X1  g356(.A(new_n557), .B(G197gat), .ZN(new_n558));
  XNOR2_X1  g357(.A(new_n558), .B(KEYINPUT11), .ZN(new_n559));
  XNOR2_X1  g358(.A(new_n559), .B(G169gat), .ZN(new_n560));
  XNOR2_X1  g359(.A(KEYINPUT87), .B(KEYINPUT12), .ZN(new_n561));
  XNOR2_X1  g360(.A(new_n560), .B(new_n561), .ZN(new_n562));
  AND3_X1   g361(.A1(new_n549), .A2(new_n556), .A3(new_n562), .ZN(new_n563));
  INV_X1    g362(.A(KEYINPUT18), .ZN(new_n564));
  NAND2_X1  g363(.A1(new_n554), .A2(new_n564), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n565), .A2(KEYINPUT93), .ZN(new_n566));
  INV_X1    g365(.A(KEYINPUT93), .ZN(new_n567));
  NAND3_X1  g366(.A1(new_n554), .A2(new_n567), .A3(new_n564), .ZN(new_n568));
  NAND2_X1  g367(.A1(new_n566), .A2(new_n568), .ZN(new_n569));
  NAND3_X1  g368(.A1(new_n549), .A2(new_n565), .A3(new_n556), .ZN(new_n570));
  INV_X1    g369(.A(new_n562), .ZN(new_n571));
  AOI22_X1  g370(.A1(new_n563), .A2(new_n569), .B1(new_n570), .B2(new_n571), .ZN(new_n572));
  AOI21_X1  g371(.A(KEYINPUT7), .B1(G85gat), .B2(G92gat), .ZN(new_n573));
  XOR2_X1   g372(.A(KEYINPUT97), .B(G92gat), .Z(new_n574));
  AOI21_X1  g373(.A(new_n573), .B1(new_n574), .B2(new_n398), .ZN(new_n575));
  NAND3_X1  g374(.A1(KEYINPUT7), .A2(G85gat), .A3(G92gat), .ZN(new_n576));
  INV_X1    g375(.A(G106gat), .ZN(new_n577));
  OR3_X1    g376(.A1(new_n285), .A2(new_n577), .A3(KEYINPUT96), .ZN(new_n578));
  OAI21_X1  g377(.A(KEYINPUT96), .B1(new_n285), .B2(new_n577), .ZN(new_n579));
  NAND3_X1  g378(.A1(new_n578), .A2(KEYINPUT8), .A3(new_n579), .ZN(new_n580));
  NAND3_X1  g379(.A1(new_n575), .A2(new_n576), .A3(new_n580), .ZN(new_n581));
  XOR2_X1   g380(.A(G99gat), .B(G106gat), .Z(new_n582));
  NAND2_X1  g381(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  INV_X1    g382(.A(new_n582), .ZN(new_n584));
  NAND4_X1  g383(.A1(new_n575), .A2(new_n580), .A3(new_n584), .A4(new_n576), .ZN(new_n585));
  NAND2_X1  g384(.A1(new_n583), .A2(new_n585), .ZN(new_n586));
  INV_X1    g385(.A(new_n586), .ZN(new_n587));
  INV_X1    g386(.A(KEYINPUT100), .ZN(new_n588));
  NAND2_X1  g387(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  NOR2_X1   g388(.A1(new_n441), .A2(G57gat), .ZN(new_n590));
  AND2_X1   g389(.A1(new_n441), .A2(G57gat), .ZN(new_n591));
  INV_X1    g390(.A(G71gat), .ZN(new_n592));
  INV_X1    g391(.A(G78gat), .ZN(new_n593));
  NOR2_X1   g392(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  OAI22_X1  g393(.A1(new_n590), .A2(new_n591), .B1(new_n594), .B2(KEYINPUT9), .ZN(new_n595));
  XOR2_X1   g394(.A(G71gat), .B(G78gat), .Z(new_n596));
  XNOR2_X1  g395(.A(new_n595), .B(new_n596), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n586), .A2(KEYINPUT100), .ZN(new_n598));
  NAND3_X1  g397(.A1(new_n589), .A2(new_n597), .A3(new_n598), .ZN(new_n599));
  INV_X1    g398(.A(new_n598), .ZN(new_n600));
  OAI21_X1  g399(.A(new_n597), .B1(new_n586), .B2(KEYINPUT100), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  AOI21_X1  g401(.A(KEYINPUT10), .B1(new_n599), .B2(new_n602), .ZN(new_n603));
  XOR2_X1   g402(.A(new_n597), .B(KEYINPUT94), .Z(new_n604));
  INV_X1    g403(.A(KEYINPUT10), .ZN(new_n605));
  NOR3_X1   g404(.A1(new_n604), .A2(new_n605), .A3(new_n586), .ZN(new_n606));
  INV_X1    g405(.A(G230gat), .ZN(new_n607));
  OAI22_X1  g406(.A1(new_n603), .A2(new_n606), .B1(new_n607), .B2(new_n275), .ZN(new_n608));
  NOR2_X1   g407(.A1(new_n607), .A2(new_n275), .ZN(new_n609));
  NAND3_X1  g408(.A1(new_n599), .A2(new_n609), .A3(new_n602), .ZN(new_n610));
  AND2_X1   g409(.A1(new_n608), .A2(new_n610), .ZN(new_n611));
  XNOR2_X1  g410(.A(G120gat), .B(G148gat), .ZN(new_n612));
  XNOR2_X1  g411(.A(new_n612), .B(KEYINPUT101), .ZN(new_n613));
  XNOR2_X1  g412(.A(new_n613), .B(new_n211), .ZN(new_n614));
  XNOR2_X1  g413(.A(new_n614), .B(new_n346), .ZN(new_n615));
  OR2_X1    g414(.A1(new_n611), .A2(new_n615), .ZN(new_n616));
  NAND3_X1  g415(.A1(new_n608), .A2(new_n610), .A3(new_n615), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  NOR2_X1   g417(.A1(new_n572), .A2(new_n618), .ZN(new_n619));
  INV_X1    g418(.A(new_n619), .ZN(new_n620));
  NOR3_X1   g419(.A1(new_n509), .A2(new_n510), .A3(new_n620), .ZN(new_n621));
  INV_X1    g420(.A(KEYINPUT21), .ZN(new_n622));
  OAI21_X1  g421(.A(new_n543), .B1(new_n604), .B2(new_n622), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n597), .A2(new_n622), .ZN(new_n624));
  XNOR2_X1  g423(.A(new_n624), .B(new_n257), .ZN(new_n625));
  XNOR2_X1  g424(.A(new_n623), .B(new_n625), .ZN(new_n626));
  XNOR2_X1  g425(.A(G183gat), .B(G211gat), .ZN(new_n627));
  XNOR2_X1  g426(.A(KEYINPUT95), .B(G155gat), .ZN(new_n628));
  XNOR2_X1  g427(.A(new_n627), .B(new_n628), .ZN(new_n629));
  XNOR2_X1  g428(.A(new_n626), .B(new_n629), .ZN(new_n630));
  XNOR2_X1  g429(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n631));
  NAND2_X1  g430(.A1(G231gat), .A2(G233gat), .ZN(new_n632));
  XOR2_X1   g431(.A(new_n631), .B(new_n632), .Z(new_n633));
  XNOR2_X1  g432(.A(new_n630), .B(new_n633), .ZN(new_n634));
  INV_X1    g433(.A(new_n634), .ZN(new_n635));
  NAND3_X1  g434(.A1(new_n551), .A2(new_n586), .A3(new_n552), .ZN(new_n636));
  NAND3_X1  g435(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n525), .A2(new_n587), .ZN(new_n638));
  NAND3_X1  g437(.A1(new_n636), .A2(new_n637), .A3(new_n638), .ZN(new_n639));
  XOR2_X1   g438(.A(G190gat), .B(G218gat), .Z(new_n640));
  INV_X1    g439(.A(new_n640), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n639), .A2(new_n641), .ZN(new_n642));
  NAND4_X1  g441(.A1(new_n636), .A2(new_n640), .A3(new_n637), .A4(new_n638), .ZN(new_n643));
  AND2_X1   g442(.A1(new_n643), .A2(KEYINPUT98), .ZN(new_n644));
  NOR2_X1   g443(.A1(new_n643), .A2(KEYINPUT98), .ZN(new_n645));
  OAI21_X1  g444(.A(new_n642), .B1(new_n644), .B2(new_n645), .ZN(new_n646));
  OAI21_X1  g445(.A(KEYINPUT99), .B1(new_n644), .B2(new_n645), .ZN(new_n647));
  XNOR2_X1  g446(.A(G134gat), .B(G162gat), .ZN(new_n648));
  AOI21_X1  g447(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n649));
  XNOR2_X1  g448(.A(new_n648), .B(new_n649), .ZN(new_n650));
  NAND3_X1  g449(.A1(new_n646), .A2(new_n647), .A3(new_n650), .ZN(new_n651));
  INV_X1    g450(.A(new_n650), .ZN(new_n652));
  OAI221_X1 g451(.A(new_n642), .B1(KEYINPUT99), .B2(new_n652), .C1(new_n644), .C2(new_n645), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n651), .A2(new_n653), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n635), .A2(new_n654), .ZN(new_n655));
  INV_X1    g454(.A(new_n655), .ZN(new_n656));
  AND2_X1   g455(.A1(new_n621), .A2(new_n656), .ZN(new_n657));
  INV_X1    g456(.A(new_n430), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  XNOR2_X1  g458(.A(new_n659), .B(G1gat), .ZN(G1324gat));
  NOR2_X1   g459(.A1(new_n528), .A2(new_n530), .ZN(new_n661));
  INV_X1    g460(.A(new_n661), .ZN(new_n662));
  NAND4_X1  g461(.A1(new_n621), .A2(new_n656), .A3(new_n470), .A4(new_n662), .ZN(new_n663));
  NOR2_X1   g462(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n664));
  NOR2_X1   g463(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n657), .A2(new_n470), .ZN(new_n666));
  AOI22_X1  g465(.A1(new_n665), .A2(KEYINPUT42), .B1(new_n666), .B2(G8gat), .ZN(new_n667));
  INV_X1    g466(.A(KEYINPUT103), .ZN(new_n668));
  XOR2_X1   g467(.A(KEYINPUT102), .B(KEYINPUT42), .Z(new_n669));
  OAI21_X1  g468(.A(new_n668), .B1(new_n665), .B2(new_n669), .ZN(new_n670));
  INV_X1    g469(.A(new_n669), .ZN(new_n671));
  OAI211_X1 g470(.A(KEYINPUT103), .B(new_n671), .C1(new_n663), .C2(new_n664), .ZN(new_n672));
  NAND3_X1  g471(.A1(new_n667), .A2(new_n670), .A3(new_n672), .ZN(new_n673));
  INV_X1    g472(.A(KEYINPUT104), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  NAND4_X1  g474(.A1(new_n667), .A2(new_n670), .A3(new_n672), .A4(KEYINPUT104), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n675), .A2(new_n676), .ZN(G1325gat));
  NAND2_X1  g476(.A1(new_n621), .A2(new_n656), .ZN(new_n678));
  AOI21_X1  g477(.A(KEYINPUT36), .B1(new_n459), .B2(new_n460), .ZN(new_n679));
  OAI21_X1  g478(.A(KEYINPUT105), .B1(new_n679), .B2(new_n475), .ZN(new_n680));
  INV_X1    g479(.A(new_n680), .ZN(new_n681));
  NOR3_X1   g480(.A1(new_n679), .A2(KEYINPUT105), .A3(new_n475), .ZN(new_n682));
  NOR2_X1   g481(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  INV_X1    g482(.A(new_n683), .ZN(new_n684));
  OAI21_X1  g483(.A(G15gat), .B1(new_n678), .B2(new_n684), .ZN(new_n685));
  INV_X1    g484(.A(new_n461), .ZN(new_n686));
  OR2_X1    g485(.A1(new_n686), .A2(G15gat), .ZN(new_n687));
  OAI21_X1  g486(.A(new_n685), .B1(new_n678), .B2(new_n687), .ZN(new_n688));
  XOR2_X1   g487(.A(new_n688), .B(KEYINPUT106), .Z(G1326gat));
  NOR2_X1   g488(.A1(new_n678), .A2(new_n466), .ZN(new_n690));
  XOR2_X1   g489(.A(KEYINPUT43), .B(G22gat), .Z(new_n691));
  XNOR2_X1  g490(.A(new_n690), .B(new_n691), .ZN(G1327gat));
  NOR2_X1   g491(.A1(new_n509), .A2(new_n510), .ZN(new_n693));
  INV_X1    g492(.A(new_n654), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  NOR2_X1   g494(.A1(new_n620), .A2(new_n635), .ZN(new_n696));
  INV_X1    g495(.A(new_n696), .ZN(new_n697));
  NOR2_X1   g496(.A1(new_n695), .A2(new_n697), .ZN(new_n698));
  NAND3_X1  g497(.A1(new_n698), .A2(new_n514), .A3(new_n658), .ZN(new_n699));
  XNOR2_X1  g498(.A(new_n699), .B(KEYINPUT45), .ZN(new_n700));
  AND2_X1   g499(.A1(new_n504), .A2(new_n506), .ZN(new_n701));
  OAI21_X1  g500(.A(new_n701), .B1(new_n681), .B2(new_n682), .ZN(new_n702));
  AOI21_X1  g501(.A(new_n654), .B1(new_n702), .B2(new_n473), .ZN(new_n703));
  INV_X1    g502(.A(KEYINPUT44), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  NOR3_X1   g504(.A1(new_n509), .A2(new_n510), .A3(new_n654), .ZN(new_n706));
  OAI21_X1  g505(.A(new_n705), .B1(new_n706), .B2(new_n704), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n707), .A2(new_n696), .ZN(new_n708));
  OAI21_X1  g507(.A(G29gat), .B1(new_n708), .B2(new_n430), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n700), .A2(new_n709), .ZN(G1328gat));
  NAND3_X1  g509(.A1(new_n698), .A2(new_n517), .A3(new_n470), .ZN(new_n711));
  XOR2_X1   g510(.A(new_n711), .B(KEYINPUT46), .Z(new_n712));
  NOR2_X1   g511(.A1(new_n708), .A2(new_n450), .ZN(new_n713));
  OAI21_X1  g512(.A(new_n712), .B1(new_n713), .B2(new_n517), .ZN(G1329gat));
  OAI21_X1  g513(.A(G43gat), .B1(new_n708), .B2(new_n684), .ZN(new_n715));
  NOR3_X1   g514(.A1(new_n695), .A2(G43gat), .A3(new_n697), .ZN(new_n716));
  AND3_X1   g515(.A1(new_n716), .A2(KEYINPUT107), .A3(new_n461), .ZN(new_n717));
  AOI21_X1  g516(.A(KEYINPUT107), .B1(new_n716), .B2(new_n461), .ZN(new_n718));
  OAI21_X1  g517(.A(new_n715), .B1(new_n717), .B2(new_n718), .ZN(new_n719));
  INV_X1    g518(.A(KEYINPUT47), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  OAI211_X1 g520(.A(new_n715), .B(KEYINPUT47), .C1(new_n717), .C2(new_n718), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n721), .A2(new_n722), .ZN(G1330gat));
  NAND2_X1  g522(.A1(new_n695), .A2(KEYINPUT44), .ZN(new_n724));
  AOI21_X1  g523(.A(new_n697), .B1(new_n724), .B2(new_n705), .ZN(new_n725));
  NAND3_X1  g524(.A1(new_n725), .A2(KEYINPUT108), .A3(new_n505), .ZN(new_n726));
  INV_X1    g525(.A(KEYINPUT108), .ZN(new_n727));
  OAI21_X1  g526(.A(new_n727), .B1(new_n708), .B2(new_n466), .ZN(new_n728));
  NAND3_X1  g527(.A1(new_n726), .A2(new_n728), .A3(G50gat), .ZN(new_n729));
  NAND3_X1  g528(.A1(new_n698), .A2(new_n312), .A3(new_n505), .ZN(new_n730));
  NAND3_X1  g529(.A1(new_n729), .A2(KEYINPUT48), .A3(new_n730), .ZN(new_n731));
  INV_X1    g530(.A(KEYINPUT48), .ZN(new_n732));
  AOI21_X1  g531(.A(new_n312), .B1(new_n725), .B2(new_n505), .ZN(new_n733));
  INV_X1    g532(.A(new_n730), .ZN(new_n734));
  OAI21_X1  g533(.A(new_n732), .B1(new_n733), .B2(new_n734), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n731), .A2(new_n735), .ZN(G1331gat));
  AND2_X1   g535(.A1(new_n616), .A2(new_n617), .ZN(new_n737));
  AOI21_X1  g536(.A(new_n737), .B1(new_n702), .B2(new_n473), .ZN(new_n738));
  AOI22_X1  g537(.A1(new_n546), .A2(new_n548), .B1(new_n555), .B2(KEYINPUT18), .ZN(new_n739));
  NAND3_X1  g538(.A1(new_n569), .A2(new_n739), .A3(new_n562), .ZN(new_n740));
  NAND2_X1  g539(.A1(new_n570), .A2(new_n571), .ZN(new_n741));
  NAND2_X1  g540(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  NOR2_X1   g541(.A1(new_n655), .A2(new_n742), .ZN(new_n743));
  NAND2_X1  g542(.A1(new_n738), .A2(new_n743), .ZN(new_n744));
  INV_X1    g543(.A(new_n744), .ZN(new_n745));
  NAND2_X1  g544(.A1(new_n745), .A2(new_n658), .ZN(new_n746));
  XNOR2_X1  g545(.A(new_n746), .B(G57gat), .ZN(G1332gat));
  XNOR2_X1  g546(.A(new_n450), .B(KEYINPUT109), .ZN(new_n748));
  INV_X1    g547(.A(new_n748), .ZN(new_n749));
  NOR2_X1   g548(.A1(new_n744), .A2(new_n749), .ZN(new_n750));
  NOR2_X1   g549(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n751));
  AND2_X1   g550(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n752));
  OAI21_X1  g551(.A(new_n750), .B1(new_n751), .B2(new_n752), .ZN(new_n753));
  OAI21_X1  g552(.A(new_n753), .B1(new_n750), .B2(new_n751), .ZN(G1333gat));
  AOI21_X1  g553(.A(new_n592), .B1(new_n745), .B2(new_n683), .ZN(new_n755));
  NAND3_X1  g554(.A1(new_n745), .A2(KEYINPUT110), .A3(new_n461), .ZN(new_n756));
  INV_X1    g555(.A(KEYINPUT110), .ZN(new_n757));
  OAI21_X1  g556(.A(new_n757), .B1(new_n744), .B2(new_n686), .ZN(new_n758));
  NAND2_X1  g557(.A1(new_n756), .A2(new_n758), .ZN(new_n759));
  AOI21_X1  g558(.A(new_n755), .B1(new_n759), .B2(new_n592), .ZN(new_n760));
  XNOR2_X1  g559(.A(new_n760), .B(KEYINPUT50), .ZN(G1334gat));
  NOR2_X1   g560(.A1(new_n744), .A2(new_n466), .ZN(new_n762));
  XNOR2_X1  g561(.A(new_n762), .B(new_n593), .ZN(G1335gat));
  INV_X1    g562(.A(new_n707), .ZN(new_n764));
  NAND2_X1  g563(.A1(new_n634), .A2(new_n572), .ZN(new_n765));
  INV_X1    g564(.A(KEYINPUT111), .ZN(new_n766));
  XNOR2_X1  g565(.A(new_n765), .B(new_n766), .ZN(new_n767));
  INV_X1    g566(.A(new_n767), .ZN(new_n768));
  NOR2_X1   g567(.A1(new_n768), .A2(new_n737), .ZN(new_n769));
  INV_X1    g568(.A(new_n769), .ZN(new_n770));
  NOR3_X1   g569(.A1(new_n764), .A2(new_n430), .A3(new_n770), .ZN(new_n771));
  INV_X1    g570(.A(KEYINPUT51), .ZN(new_n772));
  AOI21_X1  g571(.A(new_n772), .B1(new_n703), .B2(new_n767), .ZN(new_n773));
  NAND2_X1  g572(.A1(new_n504), .A2(new_n506), .ZN(new_n774));
  INV_X1    g573(.A(KEYINPUT105), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n476), .A2(new_n775), .ZN(new_n776));
  AOI21_X1  g575(.A(new_n774), .B1(new_n776), .B2(new_n680), .ZN(new_n777));
  INV_X1    g576(.A(new_n473), .ZN(new_n778));
  OAI211_X1 g577(.A(new_n694), .B(new_n767), .C1(new_n777), .C2(new_n778), .ZN(new_n779));
  NOR2_X1   g578(.A1(new_n779), .A2(KEYINPUT51), .ZN(new_n780));
  NOR2_X1   g579(.A1(new_n773), .A2(new_n780), .ZN(new_n781));
  NAND2_X1  g580(.A1(new_n781), .A2(new_n618), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n658), .A2(new_n398), .ZN(new_n783));
  OAI22_X1  g582(.A1(new_n771), .A2(new_n398), .B1(new_n782), .B2(new_n783), .ZN(G1336gat));
  INV_X1    g583(.A(KEYINPUT52), .ZN(new_n785));
  NOR3_X1   g584(.A1(new_n749), .A2(new_n737), .A3(G92gat), .ZN(new_n786));
  NAND2_X1  g585(.A1(new_n781), .A2(new_n786), .ZN(new_n787));
  NOR3_X1   g586(.A1(new_n764), .A2(new_n749), .A3(new_n770), .ZN(new_n788));
  OAI211_X1 g587(.A(new_n785), .B(new_n787), .C1(new_n788), .C2(new_n574), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n779), .A2(KEYINPUT112), .ZN(new_n790));
  OAI21_X1  g589(.A(new_n790), .B1(new_n773), .B2(new_n780), .ZN(new_n791));
  NAND3_X1  g590(.A1(new_n779), .A2(KEYINPUT112), .A3(new_n772), .ZN(new_n792));
  NAND3_X1  g591(.A1(new_n791), .A2(new_n792), .A3(new_n786), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n793), .A2(KEYINPUT113), .ZN(new_n794));
  NAND3_X1  g593(.A1(new_n707), .A2(new_n470), .A3(new_n769), .ZN(new_n795));
  INV_X1    g594(.A(new_n574), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  INV_X1    g596(.A(KEYINPUT113), .ZN(new_n798));
  NAND4_X1  g597(.A1(new_n791), .A2(new_n798), .A3(new_n792), .A4(new_n786), .ZN(new_n799));
  AND3_X1   g598(.A1(new_n794), .A2(new_n797), .A3(new_n799), .ZN(new_n800));
  OAI21_X1  g599(.A(new_n789), .B1(new_n800), .B2(new_n785), .ZN(G1337gat));
  AOI21_X1  g600(.A(new_n704), .B1(new_n693), .B2(new_n694), .ZN(new_n802));
  AOI211_X1 g601(.A(KEYINPUT44), .B(new_n654), .C1(new_n702), .C2(new_n473), .ZN(new_n803));
  OAI211_X1 g602(.A(new_n683), .B(new_n769), .C1(new_n802), .C2(new_n803), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n804), .A2(KEYINPUT114), .ZN(new_n805));
  XOR2_X1   g604(.A(KEYINPUT115), .B(G99gat), .Z(new_n806));
  INV_X1    g605(.A(KEYINPUT114), .ZN(new_n807));
  NAND4_X1  g606(.A1(new_n707), .A2(new_n807), .A3(new_n683), .A4(new_n769), .ZN(new_n808));
  NAND3_X1  g607(.A1(new_n805), .A2(new_n806), .A3(new_n808), .ZN(new_n809));
  NOR2_X1   g608(.A1(new_n686), .A2(new_n806), .ZN(new_n810));
  NAND3_X1  g609(.A1(new_n781), .A2(new_n618), .A3(new_n810), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n809), .A2(new_n811), .ZN(new_n812));
  NAND2_X1  g611(.A1(new_n812), .A2(KEYINPUT116), .ZN(new_n813));
  INV_X1    g612(.A(KEYINPUT116), .ZN(new_n814));
  NAND3_X1  g613(.A1(new_n809), .A2(new_n814), .A3(new_n811), .ZN(new_n815));
  NAND2_X1  g614(.A1(new_n813), .A2(new_n815), .ZN(G1338gat));
  OAI211_X1 g615(.A(new_n505), .B(new_n769), .C1(new_n802), .C2(new_n803), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n817), .A2(G106gat), .ZN(new_n818));
  NOR3_X1   g617(.A1(new_n737), .A2(new_n466), .A3(G106gat), .ZN(new_n819));
  AOI21_X1  g618(.A(KEYINPUT53), .B1(new_n781), .B2(new_n819), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n818), .A2(new_n820), .ZN(new_n821));
  INV_X1    g620(.A(KEYINPUT117), .ZN(new_n822));
  NAND3_X1  g621(.A1(new_n791), .A2(new_n792), .A3(new_n819), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n818), .A2(new_n823), .ZN(new_n824));
  AOI21_X1  g623(.A(new_n822), .B1(new_n824), .B2(KEYINPUT53), .ZN(new_n825));
  INV_X1    g624(.A(KEYINPUT53), .ZN(new_n826));
  AOI211_X1 g625(.A(KEYINPUT117), .B(new_n826), .C1(new_n818), .C2(new_n823), .ZN(new_n827));
  OAI21_X1  g626(.A(new_n821), .B1(new_n825), .B2(new_n827), .ZN(G1339gat));
  NOR2_X1   g627(.A1(new_n748), .A2(new_n430), .ZN(new_n829));
  INV_X1    g628(.A(new_n829), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n599), .A2(new_n602), .ZN(new_n831));
  NAND2_X1  g630(.A1(new_n831), .A2(new_n605), .ZN(new_n832));
  INV_X1    g631(.A(new_n606), .ZN(new_n833));
  AOI21_X1  g632(.A(new_n609), .B1(new_n832), .B2(new_n833), .ZN(new_n834));
  INV_X1    g633(.A(KEYINPUT54), .ZN(new_n835));
  AOI21_X1  g634(.A(new_n615), .B1(new_n834), .B2(new_n835), .ZN(new_n836));
  NAND3_X1  g635(.A1(new_n832), .A2(new_n609), .A3(new_n833), .ZN(new_n837));
  NAND3_X1  g636(.A1(new_n837), .A2(new_n608), .A3(KEYINPUT54), .ZN(new_n838));
  AOI21_X1  g637(.A(KEYINPUT55), .B1(new_n836), .B2(new_n838), .ZN(new_n839));
  INV_X1    g638(.A(new_n839), .ZN(new_n840));
  INV_X1    g639(.A(KEYINPUT118), .ZN(new_n841));
  NAND2_X1  g640(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  NAND3_X1  g641(.A1(new_n836), .A2(KEYINPUT55), .A3(new_n838), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n843), .A2(new_n617), .ZN(new_n844));
  INV_X1    g643(.A(new_n844), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n839), .A2(KEYINPUT118), .ZN(new_n846));
  NAND4_X1  g645(.A1(new_n842), .A2(new_n845), .A3(new_n742), .A4(new_n846), .ZN(new_n847));
  OAI21_X1  g646(.A(new_n553), .B1(new_n538), .B2(new_n539), .ZN(new_n848));
  NAND3_X1  g647(.A1(new_n848), .A2(G229gat), .A3(G233gat), .ZN(new_n849));
  OAI21_X1  g648(.A(new_n849), .B1(new_n546), .B2(new_n548), .ZN(new_n850));
  INV_X1    g649(.A(new_n560), .ZN(new_n851));
  NAND2_X1  g650(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  NAND3_X1  g651(.A1(new_n618), .A2(new_n740), .A3(new_n852), .ZN(new_n853));
  AOI21_X1  g652(.A(new_n694), .B1(new_n847), .B2(new_n853), .ZN(new_n854));
  NAND4_X1  g653(.A1(new_n651), .A2(new_n653), .A3(new_n617), .A4(new_n843), .ZN(new_n855));
  NAND2_X1  g654(.A1(new_n740), .A2(new_n852), .ZN(new_n856));
  NOR2_X1   g655(.A1(new_n839), .A2(KEYINPUT118), .ZN(new_n857));
  AOI211_X1 g656(.A(new_n841), .B(KEYINPUT55), .C1(new_n836), .C2(new_n838), .ZN(new_n858));
  NOR4_X1   g657(.A1(new_n855), .A2(new_n856), .A3(new_n857), .A4(new_n858), .ZN(new_n859));
  OAI21_X1  g658(.A(new_n634), .B1(new_n854), .B2(new_n859), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n743), .A2(new_n737), .ZN(new_n861));
  AOI21_X1  g660(.A(new_n830), .B1(new_n860), .B2(new_n861), .ZN(new_n862));
  NOR2_X1   g661(.A1(new_n686), .A2(new_n505), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  OAI21_X1  g663(.A(G113gat), .B1(new_n864), .B2(new_n572), .ZN(new_n865));
  INV_X1    g664(.A(new_n394), .ZN(new_n866));
  NAND2_X1  g665(.A1(new_n862), .A2(new_n866), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n742), .A2(new_n253), .ZN(new_n868));
  OAI21_X1  g667(.A(new_n865), .B1(new_n867), .B2(new_n868), .ZN(G1340gat));
  OAI21_X1  g668(.A(G120gat), .B1(new_n864), .B2(new_n737), .ZN(new_n870));
  OR2_X1    g669(.A1(new_n737), .A2(new_n265), .ZN(new_n871));
  OAI21_X1  g670(.A(new_n870), .B1(new_n867), .B2(new_n871), .ZN(G1341gat));
  NOR3_X1   g671(.A1(new_n864), .A2(new_n257), .A3(new_n634), .ZN(new_n873));
  NAND3_X1  g672(.A1(new_n862), .A2(new_n635), .A3(new_n866), .ZN(new_n874));
  AOI21_X1  g673(.A(new_n873), .B1(new_n257), .B2(new_n874), .ZN(G1342gat));
  NAND2_X1  g674(.A1(new_n860), .A2(new_n861), .ZN(new_n876));
  AND4_X1   g675(.A1(new_n658), .A2(new_n876), .A3(new_n694), .A4(new_n450), .ZN(new_n877));
  NAND3_X1  g676(.A1(new_n877), .A2(new_n258), .A3(new_n866), .ZN(new_n878));
  NAND2_X1  g677(.A1(new_n878), .A2(KEYINPUT56), .ZN(new_n879));
  OAI21_X1  g678(.A(G134gat), .B1(new_n864), .B2(new_n654), .ZN(new_n880));
  NOR2_X1   g679(.A1(new_n878), .A2(KEYINPUT56), .ZN(new_n881));
  INV_X1    g680(.A(KEYINPUT119), .ZN(new_n882));
  NOR2_X1   g681(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  NOR3_X1   g682(.A1(new_n878), .A2(KEYINPUT119), .A3(KEYINPUT56), .ZN(new_n884));
  OAI211_X1 g683(.A(new_n879), .B(new_n880), .C1(new_n883), .C2(new_n884), .ZN(G1343gat));
  AOI21_X1  g684(.A(new_n466), .B1(new_n860), .B2(new_n861), .ZN(new_n886));
  INV_X1    g685(.A(KEYINPUT57), .ZN(new_n887));
  NAND2_X1  g686(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  NOR3_X1   g687(.A1(new_n572), .A2(new_n839), .A3(new_n844), .ZN(new_n889));
  INV_X1    g688(.A(new_n853), .ZN(new_n890));
  OAI21_X1  g689(.A(new_n654), .B1(new_n889), .B2(new_n890), .ZN(new_n891));
  NOR3_X1   g690(.A1(new_n855), .A2(new_n857), .A3(new_n858), .ZN(new_n892));
  INV_X1    g691(.A(new_n856), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  AOI21_X1  g693(.A(new_n635), .B1(new_n891), .B2(new_n894), .ZN(new_n895));
  NOR3_X1   g694(.A1(new_n655), .A2(new_n618), .A3(new_n742), .ZN(new_n896));
  OAI21_X1  g695(.A(new_n505), .B1(new_n895), .B2(new_n896), .ZN(new_n897));
  NAND2_X1  g696(.A1(new_n897), .A2(KEYINPUT57), .ZN(new_n898));
  NOR2_X1   g697(.A1(new_n683), .A2(new_n830), .ZN(new_n899));
  NAND3_X1  g698(.A1(new_n888), .A2(new_n898), .A3(new_n899), .ZN(new_n900));
  INV_X1    g699(.A(new_n900), .ZN(new_n901));
  NAND2_X1  g700(.A1(new_n901), .A2(new_n742), .ZN(new_n902));
  NAND2_X1  g701(.A1(new_n902), .A2(G141gat), .ZN(new_n903));
  NAND2_X1  g702(.A1(new_n886), .A2(new_n899), .ZN(new_n904));
  NOR3_X1   g703(.A1(new_n904), .A2(G141gat), .A3(new_n572), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n905), .A2(KEYINPUT120), .ZN(new_n906));
  INV_X1    g705(.A(KEYINPUT121), .ZN(new_n907));
  NAND3_X1  g706(.A1(new_n903), .A2(new_n906), .A3(new_n907), .ZN(new_n908));
  INV_X1    g707(.A(KEYINPUT58), .ZN(new_n909));
  OAI21_X1  g708(.A(KEYINPUT120), .B1(new_n909), .B2(KEYINPUT121), .ZN(new_n910));
  AOI21_X1  g709(.A(new_n905), .B1(new_n902), .B2(G141gat), .ZN(new_n911));
  AOI22_X1  g710(.A1(new_n908), .A2(new_n909), .B1(new_n910), .B2(new_n911), .ZN(G1344gat));
  INV_X1    g711(.A(new_n904), .ZN(new_n913));
  INV_X1    g712(.A(G148gat), .ZN(new_n914));
  NAND3_X1  g713(.A1(new_n913), .A2(new_n914), .A3(new_n618), .ZN(new_n915));
  AOI211_X1 g714(.A(KEYINPUT59), .B(new_n914), .C1(new_n901), .C2(new_n618), .ZN(new_n916));
  INV_X1    g715(.A(KEYINPUT59), .ZN(new_n917));
  NAND2_X1  g716(.A1(new_n897), .A2(new_n887), .ZN(new_n918));
  NAND3_X1  g717(.A1(new_n876), .A2(KEYINPUT57), .A3(new_n505), .ZN(new_n919));
  AOI21_X1  g718(.A(new_n737), .B1(new_n918), .B2(new_n919), .ZN(new_n920));
  NAND2_X1  g719(.A1(new_n920), .A2(new_n899), .ZN(new_n921));
  AOI21_X1  g720(.A(new_n917), .B1(new_n921), .B2(G148gat), .ZN(new_n922));
  OAI21_X1  g721(.A(new_n915), .B1(new_n916), .B2(new_n922), .ZN(G1345gat));
  INV_X1    g722(.A(G155gat), .ZN(new_n924));
  NOR3_X1   g723(.A1(new_n900), .A2(new_n924), .A3(new_n634), .ZN(new_n925));
  NAND2_X1  g724(.A1(new_n913), .A2(new_n635), .ZN(new_n926));
  XNOR2_X1  g725(.A(new_n926), .B(KEYINPUT122), .ZN(new_n927));
  AOI21_X1  g726(.A(new_n925), .B1(new_n927), .B2(new_n924), .ZN(G1346gat));
  OAI21_X1  g727(.A(new_n326), .B1(new_n900), .B2(new_n654), .ZN(new_n929));
  NOR3_X1   g728(.A1(new_n683), .A2(new_n326), .A3(new_n466), .ZN(new_n930));
  NAND2_X1  g729(.A1(new_n877), .A2(new_n930), .ZN(new_n931));
  NAND2_X1  g730(.A1(new_n929), .A2(new_n931), .ZN(G1347gat));
  AOI21_X1  g731(.A(new_n658), .B1(new_n860), .B2(new_n861), .ZN(new_n933));
  AND3_X1   g732(.A1(new_n933), .A2(new_n866), .A3(new_n748), .ZN(new_n934));
  NAND3_X1  g733(.A1(new_n934), .A2(new_n247), .A3(new_n742), .ZN(new_n935));
  XNOR2_X1  g734(.A(new_n935), .B(KEYINPUT123), .ZN(new_n936));
  NAND3_X1  g735(.A1(new_n933), .A2(new_n470), .A3(new_n863), .ZN(new_n937));
  OAI21_X1  g736(.A(G169gat), .B1(new_n937), .B2(new_n572), .ZN(new_n938));
  NAND2_X1  g737(.A1(new_n936), .A2(new_n938), .ZN(G1348gat));
  NAND2_X1  g738(.A1(new_n934), .A2(new_n618), .ZN(new_n940));
  NAND2_X1  g739(.A1(new_n940), .A2(new_n211), .ZN(new_n941));
  OR3_X1    g740(.A1(new_n937), .A2(new_n248), .A3(new_n737), .ZN(new_n942));
  NAND2_X1  g741(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  XOR2_X1   g742(.A(new_n943), .B(KEYINPUT124), .Z(G1349gat));
  NAND3_X1  g743(.A1(new_n934), .A2(new_n635), .A3(new_n227), .ZN(new_n945));
  OAI21_X1  g744(.A(G183gat), .B1(new_n937), .B2(new_n634), .ZN(new_n946));
  NAND2_X1  g745(.A1(new_n945), .A2(new_n946), .ZN(new_n947));
  XNOR2_X1  g746(.A(new_n947), .B(KEYINPUT60), .ZN(G1350gat));
  NAND3_X1  g747(.A1(new_n934), .A2(new_n221), .A3(new_n694), .ZN(new_n949));
  OAI21_X1  g748(.A(G190gat), .B1(new_n937), .B2(new_n654), .ZN(new_n950));
  AND2_X1   g749(.A1(new_n950), .A2(KEYINPUT61), .ZN(new_n951));
  NOR2_X1   g750(.A1(new_n950), .A2(KEYINPUT61), .ZN(new_n952));
  OAI21_X1  g751(.A(new_n949), .B1(new_n951), .B2(new_n952), .ZN(G1351gat));
  NOR3_X1   g752(.A1(new_n683), .A2(new_n466), .A3(new_n749), .ZN(new_n954));
  OR2_X1    g753(.A1(new_n954), .A2(KEYINPUT125), .ZN(new_n955));
  NAND2_X1  g754(.A1(new_n954), .A2(KEYINPUT125), .ZN(new_n956));
  AND3_X1   g755(.A1(new_n955), .A2(new_n933), .A3(new_n956), .ZN(new_n957));
  AND2_X1   g756(.A1(new_n957), .A2(new_n341), .ZN(new_n958));
  AND3_X1   g757(.A1(new_n958), .A2(KEYINPUT126), .A3(new_n742), .ZN(new_n959));
  AOI21_X1  g758(.A(KEYINPUT126), .B1(new_n958), .B2(new_n742), .ZN(new_n960));
  NAND2_X1  g759(.A1(new_n918), .A2(new_n919), .ZN(new_n961));
  NOR3_X1   g760(.A1(new_n683), .A2(new_n658), .A3(new_n450), .ZN(new_n962));
  AND2_X1   g761(.A1(new_n961), .A2(new_n962), .ZN(new_n963));
  AND2_X1   g762(.A1(new_n963), .A2(new_n742), .ZN(new_n964));
  OAI22_X1  g763(.A1(new_n959), .A2(new_n960), .B1(new_n341), .B2(new_n964), .ZN(G1352gat));
  NAND3_X1  g764(.A1(new_n957), .A2(new_n346), .A3(new_n618), .ZN(new_n966));
  OR2_X1    g765(.A1(new_n966), .A2(KEYINPUT62), .ZN(new_n967));
  NAND2_X1  g766(.A1(new_n966), .A2(KEYINPUT62), .ZN(new_n968));
  AND2_X1   g767(.A1(new_n920), .A2(new_n962), .ZN(new_n969));
  OAI211_X1 g768(.A(new_n967), .B(new_n968), .C1(new_n346), .C2(new_n969), .ZN(G1353gat));
  INV_X1    g769(.A(new_n339), .ZN(new_n971));
  NAND3_X1  g770(.A1(new_n957), .A2(new_n635), .A3(new_n971), .ZN(new_n972));
  AOI211_X1 g771(.A(new_n887), .B(new_n466), .C1(new_n860), .C2(new_n861), .ZN(new_n973));
  NAND3_X1  g772(.A1(new_n845), .A2(new_n742), .A3(new_n840), .ZN(new_n974));
  AOI21_X1  g773(.A(new_n694), .B1(new_n974), .B2(new_n853), .ZN(new_n975));
  OAI21_X1  g774(.A(new_n634), .B1(new_n975), .B2(new_n859), .ZN(new_n976));
  NAND2_X1  g775(.A1(new_n976), .A2(new_n861), .ZN(new_n977));
  AOI21_X1  g776(.A(KEYINPUT57), .B1(new_n977), .B2(new_n505), .ZN(new_n978));
  OAI211_X1 g777(.A(new_n635), .B(new_n962), .C1(new_n973), .C2(new_n978), .ZN(new_n979));
  INV_X1    g778(.A(KEYINPUT127), .ZN(new_n980));
  NAND2_X1  g779(.A1(new_n979), .A2(new_n980), .ZN(new_n981));
  NAND4_X1  g780(.A1(new_n961), .A2(KEYINPUT127), .A3(new_n635), .A4(new_n962), .ZN(new_n982));
  NAND3_X1  g781(.A1(new_n981), .A2(new_n982), .A3(G211gat), .ZN(new_n983));
  INV_X1    g782(.A(KEYINPUT63), .ZN(new_n984));
  AND2_X1   g783(.A1(new_n983), .A2(new_n984), .ZN(new_n985));
  NOR2_X1   g784(.A1(new_n983), .A2(new_n984), .ZN(new_n986));
  OAI21_X1  g785(.A(new_n972), .B1(new_n985), .B2(new_n986), .ZN(G1354gat));
  AOI21_X1  g786(.A(G218gat), .B1(new_n957), .B2(new_n694), .ZN(new_n988));
  AND2_X1   g787(.A1(new_n694), .A2(G218gat), .ZN(new_n989));
  AOI21_X1  g788(.A(new_n988), .B1(new_n963), .B2(new_n989), .ZN(G1355gat));
endmodule


