

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
         n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706,
         n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717,
         n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
         n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739,
         n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750,
         n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761,
         n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772,
         n773, n774, n775, n776, n777, n778, n779, n780, n781, n782;

  AND2_X1 U377 ( .A1(n614), .A2(n613), .ZN(n773) );
  XNOR2_X1 U378 ( .A(KEYINPUT72), .B(KEYINPUT73), .ZN(n431) );
  NOR2_X1 U379 ( .A1(G237), .A2(G953), .ZN(n436) );
  XNOR2_X1 U380 ( .A(G146), .B(G125), .ZN(n455) );
  AND2_X2 U381 ( .A1(n566), .A2(n565), .ZN(n575) );
  XNOR2_X2 U382 ( .A(G137), .B(G140), .ZN(n770) );
  BUF_X2 U383 ( .A(n373), .Z(n548) );
  NOR2_X1 U384 ( .A1(n720), .A2(n525), .ZN(n380) );
  NOR2_X1 U385 ( .A1(n700), .A2(n692), .ZN(n535) );
  XNOR2_X1 U386 ( .A(n451), .B(KEYINPUT91), .ZN(n453) );
  NAND2_X1 U387 ( .A1(n450), .A2(G224), .ZN(n451) );
  INV_X1 U388 ( .A(G953), .ZN(n450) );
  INV_X2 U389 ( .A(G953), .ZN(n371) );
  XNOR2_X1 U390 ( .A(n630), .B(n629), .ZN(n633) );
  AND2_X1 U391 ( .A1(n734), .A2(n358), .ZN(n357) );
  AND2_X1 U392 ( .A1(n573), .A2(n572), .ZN(n574) );
  NOR2_X1 U393 ( .A1(n570), .A2(KEYINPUT69), .ZN(n544) );
  NAND2_X1 U394 ( .A1(n356), .A2(n670), .ZN(n383) );
  INV_X1 U395 ( .A(n538), .ZN(n355) );
  NAND2_X1 U396 ( .A1(n397), .A2(n691), .ZN(n699) );
  XNOR2_X1 U397 ( .A(n356), .B(G119), .ZN(G21) );
  NAND2_X2 U398 ( .A1(n385), .A2(n387), .ZN(n356) );
  AND2_X2 U399 ( .A1(n633), .A2(n734), .ZN(n372) );
  AND2_X1 U400 ( .A1(n633), .A2(n357), .ZN(n637) );
  INV_X1 U401 ( .A(n372), .ZN(n741) );
  INV_X1 U402 ( .A(n634), .ZN(n358) );
  XNOR2_X1 U403 ( .A(n383), .B(KEYINPUT88), .ZN(n359) );
  XNOR2_X1 U404 ( .A(n383), .B(KEYINPUT88), .ZN(n570) );
  XNOR2_X1 U405 ( .A(n523), .B(n362), .ZN(n360) );
  XNOR2_X1 U406 ( .A(n523), .B(n362), .ZN(n361) );
  INV_X1 U407 ( .A(n360), .ZN(n545) );
  XOR2_X1 U408 ( .A(n522), .B(KEYINPUT35), .Z(n362) );
  XNOR2_X1 U409 ( .A(n506), .B(KEYINPUT33), .ZN(n720) );
  INV_X1 U410 ( .A(G237), .ZN(n444) );
  INV_X1 U411 ( .A(KEYINPUT0), .ZN(n384) );
  AND2_X1 U412 ( .A1(n393), .A2(n604), .ZN(n392) );
  XNOR2_X1 U413 ( .A(n689), .B(KEYINPUT86), .ZN(n393) );
  XNOR2_X1 U414 ( .A(n406), .B(n405), .ZN(n490) );
  XNOR2_X1 U415 ( .A(KEYINPUT71), .B(G134), .ZN(n421) );
  XNOR2_X1 U416 ( .A(n412), .B(n411), .ZN(n531) );
  XNOR2_X1 U417 ( .A(n410), .B(n409), .ZN(n411) );
  XNOR2_X1 U418 ( .A(n530), .B(KEYINPUT22), .ZN(n538) );
  XNOR2_X1 U419 ( .A(G110), .B(n770), .ZN(n425) );
  XNOR2_X1 U420 ( .A(n578), .B(n382), .ZN(n730) );
  INV_X1 U421 ( .A(KEYINPUT41), .ZN(n382) );
  NOR2_X1 U422 ( .A1(n684), .A2(n378), .ZN(n606) );
  NAND2_X1 U423 ( .A1(n536), .A2(n368), .ZN(n388) );
  BUF_X1 U424 ( .A(n531), .Z(n579) );
  INV_X1 U425 ( .A(n700), .ZN(n394) );
  XNOR2_X1 U426 ( .A(KEYINPUT92), .B(KEYINPUT17), .ZN(n454) );
  XNOR2_X1 U427 ( .A(G902), .B(KEYINPUT15), .ZN(n622) );
  BUF_X1 U428 ( .A(n461), .Z(n435) );
  XNOR2_X1 U429 ( .A(KEYINPUT5), .B(G137), .ZN(n437) );
  XNOR2_X1 U430 ( .A(G143), .B(G140), .ZN(n467) );
  XOR2_X1 U431 ( .A(KEYINPUT12), .B(KEYINPUT98), .Z(n468) );
  AND2_X1 U432 ( .A1(n505), .A2(n601), .ZN(n506) );
  NAND2_X1 U433 ( .A1(G234), .A2(G237), .ZN(n416) );
  NOR2_X1 U434 ( .A1(n714), .A2(n528), .ZN(n529) );
  NOR2_X1 U435 ( .A1(n546), .A2(n695), .ZN(n547) );
  XNOR2_X1 U436 ( .A(G116), .B(G107), .ZN(n487) );
  INV_X1 U437 ( .A(G146), .ZN(n422) );
  INV_X1 U438 ( .A(KEYINPUT19), .ZN(n400) );
  BUF_X1 U439 ( .A(n539), .Z(n695) );
  INV_X1 U440 ( .A(n531), .ZN(n397) );
  XNOR2_X1 U441 ( .A(n398), .B(n365), .ZN(n753) );
  XNOR2_X1 U442 ( .A(n407), .B(n399), .ZN(n398) );
  XNOR2_X1 U443 ( .A(n403), .B(n404), .ZN(n399) );
  XNOR2_X1 U444 ( .A(G134), .B(G122), .ZN(n483) );
  XNOR2_X1 U445 ( .A(n656), .B(n655), .ZN(n657) );
  XNOR2_X1 U446 ( .A(n642), .B(n643), .ZN(n644) );
  NOR2_X1 U447 ( .A1(n371), .A2(G952), .ZN(n755) );
  XNOR2_X1 U448 ( .A(n586), .B(n585), .ZN(n781) );
  NAND2_X1 U449 ( .A1(n730), .A2(n671), .ZN(n586) );
  NAND2_X1 U450 ( .A1(n395), .A2(n394), .ZN(n689) );
  XNOR2_X1 U451 ( .A(n603), .B(n369), .ZN(n395) );
  NOR2_X1 U452 ( .A1(n536), .A2(n368), .ZN(n386) );
  BUF_X1 U453 ( .A(n683), .Z(n686) );
  BUF_X1 U454 ( .A(G128), .Z(n677) );
  NAND2_X1 U455 ( .A1(n355), .A2(n364), .ZN(n651) );
  XNOR2_X1 U456 ( .A(n455), .B(KEYINPUT10), .ZN(n474) );
  NOR2_X1 U457 ( .A1(n541), .A2(n394), .ZN(n363) );
  NOR2_X1 U458 ( .A1(n558), .A2(n601), .ZN(n364) );
  XOR2_X1 U459 ( .A(n425), .B(n474), .Z(n365) );
  NAND2_X1 U460 ( .A1(n466), .A2(G210), .ZN(n366) );
  AND2_X1 U461 ( .A1(n600), .A2(n599), .ZN(n367) );
  XNOR2_X1 U462 ( .A(n537), .B(KEYINPUT65), .ZN(n368) );
  XOR2_X1 U463 ( .A(KEYINPUT108), .B(KEYINPUT36), .Z(n369) );
  NAND2_X1 U464 ( .A1(n355), .A2(n363), .ZN(n670) );
  OR2_X2 U465 ( .A1(n587), .A2(n684), .ZN(n588) );
  NAND2_X1 U466 ( .A1(n355), .A2(n386), .ZN(n385) );
  NAND2_X1 U467 ( .A1(n521), .A2(n520), .ZN(n523) );
  XNOR2_X1 U468 ( .A(n380), .B(KEYINPUT34), .ZN(n521) );
  XNOR2_X1 U469 ( .A(n530), .B(KEYINPUT22), .ZN(n370) );
  NAND2_X2 U470 ( .A1(n373), .A2(n529), .ZN(n530) );
  XNOR2_X2 U471 ( .A(n519), .B(n384), .ZN(n373) );
  NAND2_X1 U472 ( .A1(n582), .A2(n598), .ZN(n396) );
  NAND2_X1 U473 ( .A1(n465), .A2(n763), .ZN(n376) );
  NAND2_X1 U474 ( .A1(n374), .A2(n375), .ZN(n377) );
  NAND2_X1 U475 ( .A1(n377), .A2(n376), .ZN(n641) );
  INV_X1 U476 ( .A(n465), .ZN(n374) );
  INV_X1 U477 ( .A(n763), .ZN(n375) );
  XNOR2_X2 U478 ( .A(n768), .B(G101), .ZN(n458) );
  XNOR2_X1 U479 ( .A(n402), .B(n366), .ZN(n507) );
  NAND2_X1 U480 ( .A1(n367), .A2(n601), .ZN(n378) );
  NOR2_X2 U481 ( .A1(n507), .A2(n577), .ZN(n401) );
  XNOR2_X1 U482 ( .A(n401), .B(n400), .ZN(n590) );
  NAND2_X1 U483 ( .A1(n518), .A2(n590), .ZN(n519) );
  NAND2_X1 U484 ( .A1(n379), .A2(KEYINPUT44), .ZN(n566) );
  NAND2_X1 U485 ( .A1(n544), .A2(n543), .ZN(n379) );
  XNOR2_X1 U486 ( .A(n381), .B(n605), .ZN(n614) );
  NAND2_X1 U487 ( .A1(n390), .A2(n392), .ZN(n381) );
  INV_X1 U488 ( .A(n548), .ZN(n525) );
  AND2_X2 U489 ( .A1(n389), .A2(n388), .ZN(n387) );
  NAND2_X1 U490 ( .A1(n370), .A2(n368), .ZN(n389) );
  XNOR2_X1 U491 ( .A(n391), .B(n589), .ZN(n390) );
  NAND2_X1 U492 ( .A1(n650), .A2(n781), .ZN(n391) );
  XNOR2_X2 U493 ( .A(n588), .B(KEYINPUT40), .ZN(n650) );
  NOR2_X1 U494 ( .A1(n699), .A2(n396), .ZN(n448) );
  NAND2_X1 U495 ( .A1(n641), .A2(n622), .ZN(n402) );
  INV_X2 U496 ( .A(n741), .ZN(n751) );
  OR2_X1 U497 ( .A1(n562), .A2(KEYINPUT87), .ZN(n563) );
  XNOR2_X1 U498 ( .A(n769), .B(n422), .ZN(n423) );
  XNOR2_X1 U499 ( .A(n550), .B(n549), .ZN(n683) );
  XOR2_X1 U500 ( .A(KEYINPUT24), .B(KEYINPUT23), .Z(n404) );
  XNOR2_X1 U501 ( .A(n677), .B(G119), .ZN(n403) );
  XOR2_X1 U502 ( .A(KEYINPUT8), .B(KEYINPUT70), .Z(n406) );
  NAND2_X1 U503 ( .A1(G234), .A2(n371), .ZN(n405) );
  NAND2_X1 U504 ( .A1(n490), .A2(G221), .ZN(n407) );
  NOR2_X1 U505 ( .A1(G902), .A2(n753), .ZN(n412) );
  NAND2_X1 U506 ( .A1(G234), .A2(n622), .ZN(n408) );
  XNOR2_X1 U507 ( .A(KEYINPUT20), .B(n408), .ZN(n413) );
  NAND2_X1 U508 ( .A1(G217), .A2(n413), .ZN(n410) );
  INV_X1 U509 ( .A(KEYINPUT25), .ZN(n409) );
  AND2_X1 U510 ( .A1(n413), .A2(G221), .ZN(n414) );
  XNOR2_X1 U511 ( .A(n414), .B(KEYINPUT21), .ZN(n691) );
  INV_X1 U512 ( .A(n691), .ZN(n528) );
  INV_X1 U513 ( .A(KEYINPUT14), .ZN(n415) );
  XNOR2_X1 U514 ( .A(n416), .B(n415), .ZN(n727) );
  INV_X1 U515 ( .A(n371), .ZN(n777) );
  NAND2_X1 U516 ( .A1(G902), .A2(n777), .ZN(n417) );
  NOR2_X1 U517 ( .A1(G900), .A2(n417), .ZN(n419) );
  NAND2_X1 U518 ( .A1(n371), .A2(G952), .ZN(n513) );
  INV_X1 U519 ( .A(n513), .ZN(n418) );
  NOR2_X1 U520 ( .A1(n419), .A2(n418), .ZN(n420) );
  NOR2_X1 U521 ( .A1(n727), .A2(n420), .ZN(n598) );
  XNOR2_X2 U522 ( .A(G143), .B(G128), .ZN(n485) );
  XNOR2_X2 U523 ( .A(n485), .B(KEYINPUT4), .ZN(n768) );
  XNOR2_X1 U524 ( .A(n421), .B(G131), .ZN(n769) );
  XNOR2_X1 U525 ( .A(n458), .B(n423), .ZN(n442) );
  XNOR2_X1 U526 ( .A(G107), .B(G104), .ZN(n424) );
  XNOR2_X1 U527 ( .A(n425), .B(n424), .ZN(n428) );
  NAND2_X1 U528 ( .A1(n371), .A2(G227), .ZN(n426) );
  XNOR2_X1 U529 ( .A(n426), .B(KEYINPUT95), .ZN(n427) );
  XNOR2_X1 U530 ( .A(n428), .B(n427), .ZN(n429) );
  XNOR2_X1 U531 ( .A(n442), .B(n429), .ZN(n744) );
  OR2_X2 U532 ( .A1(n744), .A2(G902), .ZN(n430) );
  XNOR2_X2 U533 ( .A(n430), .B(G469), .ZN(n582) );
  XNOR2_X1 U534 ( .A(KEYINPUT3), .B(G119), .ZN(n432) );
  XNOR2_X1 U535 ( .A(n432), .B(n431), .ZN(n461) );
  XNOR2_X1 U536 ( .A(G116), .B(G113), .ZN(n433) );
  XNOR2_X1 U537 ( .A(n433), .B(KEYINPUT75), .ZN(n434) );
  XNOR2_X1 U538 ( .A(n435), .B(n434), .ZN(n440) );
  XNOR2_X1 U539 ( .A(KEYINPUT76), .B(n436), .ZN(n470) );
  NAND2_X1 U540 ( .A1(n470), .A2(G210), .ZN(n438) );
  XNOR2_X1 U541 ( .A(n438), .B(n437), .ZN(n439) );
  XNOR2_X1 U542 ( .A(n440), .B(n439), .ZN(n441) );
  XNOR2_X1 U543 ( .A(n442), .B(n441), .ZN(n635) );
  OR2_X2 U544 ( .A1(n635), .A2(G902), .ZN(n443) );
  INV_X1 U545 ( .A(G472), .ZN(n634) );
  XNOR2_X2 U546 ( .A(n443), .B(n634), .ZN(n539) );
  INV_X1 U547 ( .A(G902), .ZN(n478) );
  NAND2_X1 U548 ( .A1(n478), .A2(n444), .ZN(n466) );
  AND2_X1 U549 ( .A1(n466), .A2(G214), .ZN(n577) );
  OR2_X1 U550 ( .A1(n539), .A2(n577), .ZN(n446) );
  INV_X1 U551 ( .A(KEYINPUT30), .ZN(n445) );
  XNOR2_X1 U552 ( .A(n446), .B(n445), .ZN(n447) );
  NAND2_X1 U553 ( .A1(n448), .A2(n447), .ZN(n449) );
  XNOR2_X1 U554 ( .A(n449), .B(KEYINPUT77), .ZN(n499) );
  XOR2_X1 U555 ( .A(KEYINPUT78), .B(KEYINPUT18), .Z(n452) );
  XNOR2_X1 U556 ( .A(n453), .B(n452), .ZN(n457) );
  XNOR2_X1 U557 ( .A(n455), .B(n454), .ZN(n456) );
  XNOR2_X1 U558 ( .A(n457), .B(n456), .ZN(n459) );
  XNOR2_X1 U559 ( .A(n459), .B(n458), .ZN(n465) );
  XNOR2_X2 U560 ( .A(G122), .B(G113), .ZN(n460) );
  XNOR2_X2 U561 ( .A(n460), .B(G104), .ZN(n475) );
  XNOR2_X1 U562 ( .A(n461), .B(n475), .ZN(n464) );
  XNOR2_X1 U563 ( .A(KEYINPUT16), .B(G110), .ZN(n462) );
  XNOR2_X1 U564 ( .A(n487), .B(n462), .ZN(n463) );
  XNOR2_X1 U565 ( .A(n464), .B(n463), .ZN(n763) );
  BUF_X1 U566 ( .A(n507), .Z(n610) );
  XNOR2_X1 U567 ( .A(n468), .B(n467), .ZN(n469) );
  XOR2_X1 U568 ( .A(KEYINPUT11), .B(n469), .Z(n473) );
  NAND2_X1 U569 ( .A1(n470), .A2(G214), .ZN(n471) );
  XNOR2_X1 U570 ( .A(n471), .B(G131), .ZN(n472) );
  XNOR2_X1 U571 ( .A(n473), .B(n472), .ZN(n477) );
  XNOR2_X1 U572 ( .A(n474), .B(n475), .ZN(n476) );
  XNOR2_X1 U573 ( .A(n477), .B(n476), .ZN(n656) );
  NAND2_X1 U574 ( .A1(n656), .A2(n478), .ZN(n482) );
  XOR2_X1 U575 ( .A(KEYINPUT99), .B(KEYINPUT13), .Z(n480) );
  XNOR2_X1 U576 ( .A(KEYINPUT100), .B(G475), .ZN(n479) );
  XNOR2_X1 U577 ( .A(n480), .B(n479), .ZN(n481) );
  XNOR2_X1 U578 ( .A(n482), .B(n481), .ZN(n527) );
  XOR2_X1 U579 ( .A(KEYINPUT103), .B(KEYINPUT9), .Z(n484) );
  XNOR2_X1 U580 ( .A(n484), .B(n483), .ZN(n494) );
  BUF_X1 U581 ( .A(n485), .Z(n486) );
  XNOR2_X1 U582 ( .A(n486), .B(n487), .ZN(n489) );
  XOR2_X1 U583 ( .A(KEYINPUT7), .B(KEYINPUT102), .Z(n488) );
  XNOR2_X1 U584 ( .A(n489), .B(n488), .ZN(n492) );
  NAND2_X1 U585 ( .A1(G217), .A2(n490), .ZN(n491) );
  XOR2_X1 U586 ( .A(n492), .B(n491), .Z(n493) );
  XNOR2_X1 U587 ( .A(n494), .B(n493), .ZN(n748) );
  NOR2_X1 U588 ( .A1(G902), .A2(n748), .ZN(n495) );
  XNOR2_X1 U589 ( .A(G478), .B(n495), .ZN(n526) );
  NOR2_X1 U590 ( .A1(n527), .A2(n526), .ZN(n520) );
  INV_X1 U591 ( .A(n520), .ZN(n496) );
  NOR2_X1 U592 ( .A1(n610), .A2(n496), .ZN(n497) );
  NAND2_X1 U593 ( .A1(n499), .A2(n497), .ZN(n596) );
  XNOR2_X1 U594 ( .A(n596), .B(G143), .ZN(G45) );
  XNOR2_X1 U595 ( .A(KEYINPUT74), .B(KEYINPUT38), .ZN(n498) );
  XNOR2_X1 U596 ( .A(n610), .B(n498), .ZN(n712) );
  NAND2_X1 U597 ( .A1(n499), .A2(n712), .ZN(n501) );
  INV_X1 U598 ( .A(KEYINPUT39), .ZN(n500) );
  XNOR2_X1 U599 ( .A(n501), .B(n500), .ZN(n587) );
  INV_X1 U600 ( .A(KEYINPUT101), .ZN(n502) );
  XNOR2_X1 U601 ( .A(n527), .B(n502), .ZN(n555) );
  INV_X1 U602 ( .A(n526), .ZN(n554) );
  NAND2_X1 U603 ( .A1(n555), .A2(n554), .ZN(n687) );
  OR2_X1 U604 ( .A1(n587), .A2(n687), .ZN(n612) );
  XNOR2_X1 U605 ( .A(n612), .B(G134), .ZN(G36) );
  INV_X1 U606 ( .A(n699), .ZN(n504) );
  XNOR2_X1 U607 ( .A(KEYINPUT66), .B(KEYINPUT1), .ZN(n503) );
  XNOR2_X1 U608 ( .A(n582), .B(n503), .ZN(n540) );
  NAND2_X1 U609 ( .A1(n504), .A2(n540), .ZN(n546) );
  INV_X1 U610 ( .A(n546), .ZN(n505) );
  XNOR2_X1 U611 ( .A(n539), .B(KEYINPUT6), .ZN(n601) );
  NOR2_X1 U612 ( .A1(G898), .A2(n371), .ZN(n508) );
  XOR2_X1 U613 ( .A(KEYINPUT93), .B(n508), .Z(n764) );
  NAND2_X1 U614 ( .A1(G902), .A2(n764), .ZN(n511) );
  OR2_X1 U615 ( .A1(n727), .A2(n511), .ZN(n510) );
  INV_X1 U616 ( .A(KEYINPUT94), .ZN(n509) );
  NAND2_X1 U617 ( .A1(n510), .A2(n509), .ZN(n517) );
  INV_X1 U618 ( .A(n511), .ZN(n512) );
  NAND2_X1 U619 ( .A1(KEYINPUT94), .A2(n512), .ZN(n514) );
  AND2_X1 U620 ( .A1(n514), .A2(n513), .ZN(n515) );
  OR2_X1 U621 ( .A1(n727), .A2(n515), .ZN(n516) );
  NAND2_X1 U622 ( .A1(n517), .A2(n516), .ZN(n518) );
  INV_X1 U623 ( .A(KEYINPUT84), .ZN(n522) );
  XNOR2_X1 U624 ( .A(G122), .B(KEYINPUT126), .ZN(n524) );
  XNOR2_X1 U625 ( .A(n545), .B(n524), .ZN(G24) );
  NAND2_X1 U626 ( .A1(n527), .A2(n526), .ZN(n714) );
  INV_X1 U627 ( .A(KEYINPUT104), .ZN(n532) );
  XNOR2_X1 U628 ( .A(n579), .B(n532), .ZN(n692) );
  INV_X1 U629 ( .A(n540), .ZN(n700) );
  INV_X1 U630 ( .A(KEYINPUT80), .ZN(n533) );
  XNOR2_X1 U631 ( .A(n601), .B(n533), .ZN(n534) );
  NAND2_X1 U632 ( .A1(n535), .A2(n534), .ZN(n536) );
  XNOR2_X1 U633 ( .A(KEYINPUT79), .B(KEYINPUT32), .ZN(n537) );
  NAND2_X1 U634 ( .A1(n579), .A2(n695), .ZN(n541) );
  INV_X1 U635 ( .A(KEYINPUT87), .ZN(n542) );
  NAND2_X1 U636 ( .A1(n361), .A2(n542), .ZN(n543) );
  XNOR2_X1 U637 ( .A(n547), .B(KEYINPUT96), .ZN(n705) );
  NAND2_X1 U638 ( .A1(n705), .A2(n548), .ZN(n550) );
  XNOR2_X1 U639 ( .A(KEYINPUT97), .B(KEYINPUT31), .ZN(n549) );
  INV_X1 U640 ( .A(n582), .ZN(n551) );
  NOR2_X1 U641 ( .A1(n699), .A2(n551), .ZN(n552) );
  NAND2_X1 U642 ( .A1(n552), .A2(n695), .ZN(n553) );
  OR2_X1 U643 ( .A1(n525), .A2(n553), .ZN(n666) );
  NAND2_X1 U644 ( .A1(n683), .A2(n666), .ZN(n557) );
  OR2_X1 U645 ( .A1(n555), .A2(n554), .ZN(n684) );
  AND2_X1 U646 ( .A1(n687), .A2(n684), .ZN(n716) );
  INV_X1 U647 ( .A(n716), .ZN(n556) );
  NAND2_X1 U648 ( .A1(n557), .A2(n556), .ZN(n559) );
  NAND2_X1 U649 ( .A1(n692), .A2(n700), .ZN(n558) );
  NAND2_X1 U650 ( .A1(n559), .A2(n651), .ZN(n562) );
  INV_X1 U651 ( .A(n562), .ZN(n560) );
  AND2_X1 U652 ( .A1(KEYINPUT44), .A2(n560), .ZN(n561) );
  NAND2_X1 U653 ( .A1(n360), .A2(n561), .ZN(n564) );
  NAND2_X1 U654 ( .A1(n564), .A2(n563), .ZN(n565) );
  INV_X1 U655 ( .A(KEYINPUT69), .ZN(n567) );
  NOR2_X1 U656 ( .A1(n359), .A2(n567), .ZN(n568) );
  NAND2_X1 U657 ( .A1(n568), .A2(n360), .ZN(n573) );
  OR2_X1 U658 ( .A1(KEYINPUT69), .A2(KEYINPUT44), .ZN(n569) );
  NOR2_X1 U659 ( .A1(n359), .A2(n569), .ZN(n571) );
  NAND2_X1 U660 ( .A1(n571), .A2(n545), .ZN(n572) );
  NAND2_X1 U661 ( .A1(n575), .A2(n574), .ZN(n576) );
  XNOR2_X1 U662 ( .A(n576), .B(KEYINPUT45), .ZN(n756) );
  INV_X1 U663 ( .A(n577), .ZN(n711) );
  NAND2_X1 U664 ( .A1(n712), .A2(n711), .ZN(n715) );
  NOR2_X1 U665 ( .A1(n715), .A2(n714), .ZN(n578) );
  AND2_X1 U666 ( .A1(n579), .A2(n691), .ZN(n600) );
  NAND2_X1 U667 ( .A1(n600), .A2(n598), .ZN(n580) );
  NOR2_X1 U668 ( .A1(n580), .A2(n695), .ZN(n581) );
  XNOR2_X1 U669 ( .A(n581), .B(KEYINPUT28), .ZN(n583) );
  AND2_X1 U670 ( .A1(n582), .A2(n583), .ZN(n671) );
  INV_X1 U671 ( .A(KEYINPUT107), .ZN(n584) );
  XNOR2_X1 U672 ( .A(n584), .B(KEYINPUT42), .ZN(n585) );
  INV_X1 U673 ( .A(KEYINPUT46), .ZN(n589) );
  BUF_X1 U674 ( .A(n590), .Z(n591) );
  INV_X1 U675 ( .A(n591), .ZN(n592) );
  NOR2_X1 U676 ( .A1(n592), .A2(n716), .ZN(n593) );
  NAND2_X1 U677 ( .A1(n671), .A2(n593), .ZN(n595) );
  INV_X1 U678 ( .A(KEYINPUT47), .ZN(n594) );
  XNOR2_X1 U679 ( .A(n595), .B(n594), .ZN(n597) );
  AND2_X1 U680 ( .A1(n597), .A2(n596), .ZN(n604) );
  AND2_X1 U681 ( .A1(n598), .A2(n711), .ZN(n599) );
  INV_X1 U682 ( .A(n610), .ZN(n602) );
  NAND2_X1 U683 ( .A1(n606), .A2(n602), .ZN(n603) );
  INV_X1 U684 ( .A(KEYINPUT48), .ZN(n605) );
  XOR2_X1 U685 ( .A(KEYINPUT105), .B(n606), .Z(n607) );
  NAND2_X1 U686 ( .A1(n607), .A2(n700), .ZN(n609) );
  XNOR2_X1 U687 ( .A(KEYINPUT106), .B(KEYINPUT43), .ZN(n608) );
  XNOR2_X1 U688 ( .A(n609), .B(n608), .ZN(n611) );
  NAND2_X1 U689 ( .A1(n611), .A2(n610), .ZN(n652) );
  AND2_X1 U690 ( .A1(n652), .A2(n612), .ZN(n613) );
  AND2_X2 U691 ( .A1(n756), .A2(n773), .ZN(n631) );
  INV_X1 U692 ( .A(n622), .ZN(n617) );
  NAND2_X1 U693 ( .A1(KEYINPUT2), .A2(KEYINPUT83), .ZN(n615) );
  NAND2_X1 U694 ( .A1(n615), .A2(KEYINPUT82), .ZN(n616) );
  OR2_X1 U695 ( .A1(n617), .A2(n616), .ZN(n619) );
  AND2_X1 U696 ( .A1(KEYINPUT82), .A2(n619), .ZN(n618) );
  NAND2_X1 U697 ( .A1(n631), .A2(n618), .ZN(n626) );
  INV_X1 U698 ( .A(n619), .ZN(n624) );
  INV_X1 U699 ( .A(KEYINPUT2), .ZN(n620) );
  NOR2_X1 U700 ( .A1(n620), .A2(KEYINPUT83), .ZN(n621) );
  NOR2_X1 U701 ( .A1(n622), .A2(n621), .ZN(n623) );
  OR2_X1 U702 ( .A1(n624), .A2(n623), .ZN(n625) );
  NAND2_X1 U703 ( .A1(n626), .A2(n625), .ZN(n628) );
  NOR2_X1 U704 ( .A1(n631), .A2(KEYINPUT82), .ZN(n627) );
  NOR2_X2 U705 ( .A1(n628), .A2(n627), .ZN(n630) );
  INV_X1 U706 ( .A(KEYINPUT64), .ZN(n629) );
  BUF_X1 U707 ( .A(n631), .Z(n632) );
  NAND2_X1 U708 ( .A1(n632), .A2(KEYINPUT2), .ZN(n734) );
  XOR2_X1 U709 ( .A(KEYINPUT62), .B(n635), .Z(n636) );
  XNOR2_X1 U710 ( .A(n637), .B(n636), .ZN(n638) );
  NOR2_X1 U711 ( .A1(n638), .A2(n755), .ZN(n640) );
  XOR2_X1 U712 ( .A(KEYINPUT90), .B(KEYINPUT63), .Z(n639) );
  XNOR2_X1 U713 ( .A(n640), .B(n639), .ZN(G57) );
  NAND2_X1 U714 ( .A1(n372), .A2(G210), .ZN(n645) );
  BUF_X1 U715 ( .A(n641), .Z(n642) );
  XNOR2_X1 U716 ( .A(KEYINPUT54), .B(KEYINPUT55), .ZN(n643) );
  XNOR2_X1 U717 ( .A(n645), .B(n644), .ZN(n646) );
  NOR2_X2 U718 ( .A1(n646), .A2(n755), .ZN(n649) );
  XNOR2_X1 U719 ( .A(KEYINPUT121), .B(KEYINPUT56), .ZN(n647) );
  XNOR2_X1 U720 ( .A(n647), .B(KEYINPUT85), .ZN(n648) );
  XNOR2_X1 U721 ( .A(n649), .B(n648), .ZN(G51) );
  XNOR2_X1 U722 ( .A(n650), .B(G131), .ZN(G33) );
  XNOR2_X1 U723 ( .A(n651), .B(G101), .ZN(G3) );
  XNOR2_X1 U724 ( .A(n652), .B(G140), .ZN(G42) );
  NAND2_X1 U725 ( .A1(n372), .A2(G475), .ZN(n658) );
  XOR2_X1 U726 ( .A(KEYINPUT89), .B(KEYINPUT67), .Z(n654) );
  XNOR2_X1 U727 ( .A(KEYINPUT59), .B(KEYINPUT123), .ZN(n653) );
  XNOR2_X1 U728 ( .A(n654), .B(n653), .ZN(n655) );
  XNOR2_X1 U729 ( .A(n658), .B(n657), .ZN(n659) );
  NOR2_X2 U730 ( .A1(n659), .A2(n755), .ZN(n662) );
  XNOR2_X1 U731 ( .A(KEYINPUT124), .B(KEYINPUT60), .ZN(n660) );
  XNOR2_X1 U732 ( .A(n660), .B(KEYINPUT68), .ZN(n661) );
  XNOR2_X1 U733 ( .A(n662), .B(n661), .ZN(G60) );
  NOR2_X1 U734 ( .A1(n684), .A2(n666), .ZN(n664) );
  XNOR2_X1 U735 ( .A(KEYINPUT109), .B(KEYINPUT110), .ZN(n663) );
  XNOR2_X1 U736 ( .A(n664), .B(n663), .ZN(n665) );
  XNOR2_X1 U737 ( .A(G104), .B(n665), .ZN(G6) );
  NOR2_X1 U738 ( .A1(n687), .A2(n666), .ZN(n668) );
  XNOR2_X1 U739 ( .A(KEYINPUT27), .B(KEYINPUT26), .ZN(n667) );
  XNOR2_X1 U740 ( .A(n668), .B(n667), .ZN(n669) );
  XNOR2_X1 U741 ( .A(G107), .B(n669), .ZN(G9) );
  XNOR2_X1 U742 ( .A(n670), .B(G110), .ZN(G12) );
  INV_X1 U743 ( .A(n671), .ZN(n680) );
  INV_X1 U744 ( .A(n687), .ZN(n672) );
  NAND2_X1 U745 ( .A1(n672), .A2(n591), .ZN(n673) );
  NOR2_X1 U746 ( .A1(n680), .A2(n673), .ZN(n675) );
  XNOR2_X1 U747 ( .A(KEYINPUT29), .B(KEYINPUT111), .ZN(n674) );
  XNOR2_X1 U748 ( .A(n675), .B(n674), .ZN(n676) );
  XOR2_X1 U749 ( .A(n677), .B(n676), .Z(G30) );
  INV_X1 U750 ( .A(n684), .ZN(n678) );
  NAND2_X1 U751 ( .A1(n591), .A2(n678), .ZN(n679) );
  NOR2_X1 U752 ( .A1(n680), .A2(n679), .ZN(n681) );
  XOR2_X1 U753 ( .A(KEYINPUT112), .B(n681), .Z(n682) );
  XNOR2_X1 U754 ( .A(G146), .B(n682), .ZN(G48) );
  NOR2_X1 U755 ( .A1(n684), .A2(n686), .ZN(n685) );
  XOR2_X1 U756 ( .A(G113), .B(n685), .Z(G15) );
  NOR2_X1 U757 ( .A1(n687), .A2(n686), .ZN(n688) );
  XOR2_X1 U758 ( .A(G116), .B(n688), .Z(G18) );
  XOR2_X1 U759 ( .A(G125), .B(n689), .Z(n690) );
  XNOR2_X1 U760 ( .A(n690), .B(KEYINPUT37), .ZN(G27) );
  XOR2_X1 U761 ( .A(KEYINPUT120), .B(KEYINPUT53), .Z(n740) );
  NOR2_X1 U762 ( .A1(n692), .A2(n691), .ZN(n694) );
  XNOR2_X1 U763 ( .A(KEYINPUT113), .B(KEYINPUT49), .ZN(n693) );
  XNOR2_X1 U764 ( .A(n694), .B(n693), .ZN(n697) );
  INV_X1 U765 ( .A(n695), .ZN(n696) );
  NOR2_X1 U766 ( .A1(n697), .A2(n696), .ZN(n698) );
  XOR2_X1 U767 ( .A(KEYINPUT114), .B(n698), .Z(n704) );
  NAND2_X1 U768 ( .A1(n700), .A2(n699), .ZN(n701) );
  XNOR2_X1 U769 ( .A(n701), .B(KEYINPUT115), .ZN(n702) );
  XNOR2_X1 U770 ( .A(KEYINPUT50), .B(n702), .ZN(n703) );
  NOR2_X1 U771 ( .A1(n704), .A2(n703), .ZN(n706) );
  NOR2_X1 U772 ( .A1(n706), .A2(n705), .ZN(n708) );
  XNOR2_X1 U773 ( .A(KEYINPUT116), .B(KEYINPUT51), .ZN(n707) );
  XNOR2_X1 U774 ( .A(n708), .B(n707), .ZN(n709) );
  NAND2_X1 U775 ( .A1(n730), .A2(n709), .ZN(n710) );
  XNOR2_X1 U776 ( .A(n710), .B(KEYINPUT117), .ZN(n723) );
  NOR2_X1 U777 ( .A1(n712), .A2(n711), .ZN(n713) );
  NOR2_X1 U778 ( .A1(n714), .A2(n713), .ZN(n718) );
  NOR2_X1 U779 ( .A1(n716), .A2(n715), .ZN(n717) );
  NOR2_X1 U780 ( .A1(n718), .A2(n717), .ZN(n719) );
  XNOR2_X1 U781 ( .A(KEYINPUT118), .B(n719), .ZN(n721) );
  NOR2_X1 U782 ( .A1(n721), .A2(n720), .ZN(n722) );
  NOR2_X1 U783 ( .A1(n723), .A2(n722), .ZN(n724) );
  XOR2_X1 U784 ( .A(n724), .B(KEYINPUT119), .Z(n725) );
  XNOR2_X1 U785 ( .A(KEYINPUT52), .B(n725), .ZN(n726) );
  NOR2_X1 U786 ( .A1(n727), .A2(n726), .ZN(n728) );
  NAND2_X1 U787 ( .A1(n728), .A2(G952), .ZN(n732) );
  INV_X1 U788 ( .A(n720), .ZN(n729) );
  NAND2_X1 U789 ( .A1(n730), .A2(n729), .ZN(n731) );
  NAND2_X1 U790 ( .A1(n732), .A2(n731), .ZN(n737) );
  NOR2_X1 U791 ( .A1(n632), .A2(KEYINPUT2), .ZN(n733) );
  XNOR2_X1 U792 ( .A(n733), .B(KEYINPUT81), .ZN(n735) );
  AND2_X1 U793 ( .A1(n735), .A2(n734), .ZN(n736) );
  NOR2_X1 U794 ( .A1(n737), .A2(n736), .ZN(n738) );
  NAND2_X1 U795 ( .A1(n738), .A2(n371), .ZN(n739) );
  XNOR2_X1 U796 ( .A(n740), .B(n739), .ZN(G75) );
  NAND2_X1 U797 ( .A1(n751), .A2(G469), .ZN(n746) );
  XOR2_X1 U798 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n742) );
  XNOR2_X1 U799 ( .A(n742), .B(KEYINPUT122), .ZN(n743) );
  XNOR2_X1 U800 ( .A(n744), .B(n743), .ZN(n745) );
  XNOR2_X1 U801 ( .A(n746), .B(n745), .ZN(n747) );
  NOR2_X1 U802 ( .A1(n755), .A2(n747), .ZN(G54) );
  NAND2_X1 U803 ( .A1(n751), .A2(G478), .ZN(n749) );
  XNOR2_X1 U804 ( .A(n749), .B(n748), .ZN(n750) );
  NOR2_X1 U805 ( .A1(n755), .A2(n750), .ZN(G63) );
  NAND2_X1 U806 ( .A1(n751), .A2(G217), .ZN(n752) );
  XNOR2_X1 U807 ( .A(n753), .B(n752), .ZN(n754) );
  NOR2_X1 U808 ( .A1(n755), .A2(n754), .ZN(G66) );
  BUF_X1 U809 ( .A(n756), .Z(n757) );
  NAND2_X1 U810 ( .A1(n757), .A2(n371), .ZN(n762) );
  NAND2_X1 U811 ( .A1(n777), .A2(G224), .ZN(n758) );
  XNOR2_X1 U812 ( .A(KEYINPUT61), .B(n758), .ZN(n759) );
  NAND2_X1 U813 ( .A1(n759), .A2(G898), .ZN(n760) );
  XOR2_X1 U814 ( .A(KEYINPUT125), .B(n760), .Z(n761) );
  NAND2_X1 U815 ( .A1(n762), .A2(n761), .ZN(n767) );
  XOR2_X1 U816 ( .A(n763), .B(G101), .Z(n765) );
  NOR2_X1 U817 ( .A1(n765), .A2(n764), .ZN(n766) );
  XNOR2_X1 U818 ( .A(n767), .B(n766), .ZN(G69) );
  XNOR2_X1 U819 ( .A(n768), .B(n474), .ZN(n772) );
  XOR2_X1 U820 ( .A(n770), .B(n769), .Z(n771) );
  XNOR2_X1 U821 ( .A(n772), .B(n771), .ZN(n775) );
  XNOR2_X1 U822 ( .A(n773), .B(n775), .ZN(n774) );
  NAND2_X1 U823 ( .A1(n774), .A2(n371), .ZN(n780) );
  XOR2_X1 U824 ( .A(G227), .B(n775), .Z(n776) );
  NAND2_X1 U825 ( .A1(n776), .A2(G900), .ZN(n778) );
  NAND2_X1 U826 ( .A1(n778), .A2(n777), .ZN(n779) );
  NAND2_X1 U827 ( .A1(n780), .A2(n779), .ZN(G72) );
  XOR2_X1 U828 ( .A(G137), .B(n781), .Z(n782) );
  XNOR2_X1 U829 ( .A(KEYINPUT127), .B(n782), .ZN(G39) );
endmodule

