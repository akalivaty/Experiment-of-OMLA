

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579;

  XNOR2_X1 U320 ( .A(n494), .B(n493), .ZN(n495) );
  XNOR2_X1 U321 ( .A(n496), .B(n495), .ZN(n497) );
  XNOR2_X1 U322 ( .A(n410), .B(n409), .ZN(n418) );
  XNOR2_X1 U323 ( .A(n418), .B(n417), .ZN(n422) );
  XNOR2_X1 U324 ( .A(n508), .B(KEYINPUT48), .ZN(n509) );
  XNOR2_X1 U325 ( .A(n510), .B(n509), .ZN(n538) );
  XNOR2_X1 U326 ( .A(n547), .B(n546), .ZN(n557) );
  XOR2_X1 U327 ( .A(KEYINPUT93), .B(KEYINPUT6), .Z(n289) );
  XNOR2_X1 U328 ( .A(G1GAT), .B(G57GAT), .ZN(n288) );
  XNOR2_X1 U329 ( .A(n289), .B(n288), .ZN(n293) );
  XOR2_X1 U330 ( .A(KEYINPUT4), .B(KEYINPUT5), .Z(n291) );
  XNOR2_X1 U331 ( .A(KEYINPUT1), .B(KEYINPUT89), .ZN(n290) );
  XNOR2_X1 U332 ( .A(n291), .B(n290), .ZN(n292) );
  XOR2_X1 U333 ( .A(n293), .B(n292), .Z(n298) );
  XOR2_X1 U334 ( .A(KEYINPUT90), .B(KEYINPUT91), .Z(n295) );
  NAND2_X1 U335 ( .A1(G225GAT), .A2(G233GAT), .ZN(n294) );
  XNOR2_X1 U336 ( .A(n295), .B(n294), .ZN(n296) );
  XNOR2_X1 U337 ( .A(KEYINPUT92), .B(n296), .ZN(n297) );
  XNOR2_X1 U338 ( .A(n298), .B(n297), .ZN(n310) );
  XOR2_X1 U339 ( .A(G85GAT), .B(G162GAT), .Z(n300) );
  XNOR2_X1 U340 ( .A(G29GAT), .B(G134GAT), .ZN(n299) );
  XNOR2_X1 U341 ( .A(n300), .B(n299), .ZN(n304) );
  XOR2_X1 U342 ( .A(G155GAT), .B(G148GAT), .Z(n302) );
  XNOR2_X1 U343 ( .A(G127GAT), .B(G120GAT), .ZN(n301) );
  XNOR2_X1 U344 ( .A(n302), .B(n301), .ZN(n303) );
  XOR2_X1 U345 ( .A(n304), .B(n303), .Z(n308) );
  XNOR2_X1 U346 ( .A(G113GAT), .B(KEYINPUT0), .ZN(n305) );
  XNOR2_X1 U347 ( .A(n305), .B(KEYINPUT80), .ZN(n364) );
  XNOR2_X1 U348 ( .A(G141GAT), .B(KEYINPUT3), .ZN(n306) );
  XNOR2_X1 U349 ( .A(n306), .B(KEYINPUT2), .ZN(n344) );
  XNOR2_X1 U350 ( .A(n364), .B(n344), .ZN(n307) );
  XNOR2_X1 U351 ( .A(n308), .B(n307), .ZN(n309) );
  XOR2_X1 U352 ( .A(n310), .B(n309), .Z(n563) );
  XOR2_X1 U353 ( .A(KEYINPUT79), .B(G106GAT), .Z(n312) );
  XNOR2_X1 U354 ( .A(G190GAT), .B(G99GAT), .ZN(n311) );
  XNOR2_X1 U355 ( .A(n312), .B(n311), .ZN(n328) );
  XOR2_X1 U356 ( .A(KEYINPUT66), .B(KEYINPUT9), .Z(n314) );
  NAND2_X1 U357 ( .A1(G232GAT), .A2(G233GAT), .ZN(n313) );
  XNOR2_X1 U358 ( .A(n314), .B(n313), .ZN(n315) );
  XOR2_X1 U359 ( .A(n315), .B(KEYINPUT10), .Z(n320) );
  XOR2_X1 U360 ( .A(G29GAT), .B(G36GAT), .Z(n317) );
  XNOR2_X1 U361 ( .A(KEYINPUT8), .B(KEYINPUT7), .ZN(n316) );
  XNOR2_X1 U362 ( .A(n317), .B(n316), .ZN(n408) );
  XNOR2_X1 U363 ( .A(G85GAT), .B(KEYINPUT77), .ZN(n318) );
  XNOR2_X1 U364 ( .A(n318), .B(G92GAT), .ZN(n431) );
  XNOR2_X1 U365 ( .A(n408), .B(n431), .ZN(n319) );
  XNOR2_X1 U366 ( .A(n320), .B(n319), .ZN(n324) );
  XOR2_X1 U367 ( .A(KEYINPUT78), .B(KEYINPUT11), .Z(n322) );
  XNOR2_X1 U368 ( .A(G218GAT), .B(KEYINPUT65), .ZN(n321) );
  XNOR2_X1 U369 ( .A(n322), .B(n321), .ZN(n323) );
  XOR2_X1 U370 ( .A(n324), .B(n323), .Z(n326) );
  XOR2_X1 U371 ( .A(G43GAT), .B(G134GAT), .Z(n361) );
  XOR2_X1 U372 ( .A(G50GAT), .B(G162GAT), .Z(n343) );
  XNOR2_X1 U373 ( .A(n361), .B(n343), .ZN(n325) );
  XNOR2_X1 U374 ( .A(n326), .B(n325), .ZN(n327) );
  XNOR2_X1 U375 ( .A(n328), .B(n327), .ZN(n498) );
  XOR2_X1 U376 ( .A(G211GAT), .B(G78GAT), .Z(n330) );
  XNOR2_X1 U377 ( .A(G183GAT), .B(G71GAT), .ZN(n329) );
  XNOR2_X1 U378 ( .A(n330), .B(n329), .ZN(n341) );
  XNOR2_X1 U379 ( .A(G57GAT), .B(KEYINPUT13), .ZN(n331) );
  XNOR2_X1 U380 ( .A(n331), .B(KEYINPUT76), .ZN(n432) );
  XOR2_X1 U381 ( .A(G15GAT), .B(G127GAT), .Z(n360) );
  XOR2_X1 U382 ( .A(n432), .B(n360), .Z(n333) );
  NAND2_X1 U383 ( .A1(G231GAT), .A2(G233GAT), .ZN(n332) );
  XNOR2_X1 U384 ( .A(n333), .B(n332), .ZN(n337) );
  XOR2_X1 U385 ( .A(KEYINPUT15), .B(KEYINPUT12), .Z(n335) );
  XNOR2_X1 U386 ( .A(G64GAT), .B(KEYINPUT14), .ZN(n334) );
  XNOR2_X1 U387 ( .A(n335), .B(n334), .ZN(n336) );
  XOR2_X1 U388 ( .A(n337), .B(n336), .Z(n339) );
  XOR2_X1 U389 ( .A(G8GAT), .B(G1GAT), .Z(n414) );
  XOR2_X1 U390 ( .A(G22GAT), .B(G155GAT), .Z(n348) );
  XNOR2_X1 U391 ( .A(n414), .B(n348), .ZN(n338) );
  XNOR2_X1 U392 ( .A(n339), .B(n338), .ZN(n340) );
  XNOR2_X1 U393 ( .A(n341), .B(n340), .ZN(n574) );
  NAND2_X1 U394 ( .A1(n498), .A2(n574), .ZN(n342) );
  XOR2_X1 U395 ( .A(KEYINPUT16), .B(n342), .Z(n407) );
  XOR2_X1 U396 ( .A(n344), .B(n343), .Z(n346) );
  NAND2_X1 U397 ( .A1(G228GAT), .A2(G233GAT), .ZN(n345) );
  XNOR2_X1 U398 ( .A(n346), .B(n345), .ZN(n347) );
  XOR2_X1 U399 ( .A(n347), .B(KEYINPUT87), .Z(n350) );
  XNOR2_X1 U400 ( .A(n348), .B(KEYINPUT88), .ZN(n349) );
  XNOR2_X1 U401 ( .A(n350), .B(n349), .ZN(n354) );
  XOR2_X1 U402 ( .A(G204GAT), .B(KEYINPUT22), .Z(n352) );
  XNOR2_X1 U403 ( .A(KEYINPUT23), .B(KEYINPUT24), .ZN(n351) );
  XNOR2_X1 U404 ( .A(n352), .B(n351), .ZN(n353) );
  XOR2_X1 U405 ( .A(n354), .B(n353), .Z(n359) );
  XNOR2_X1 U406 ( .A(G106GAT), .B(G78GAT), .ZN(n355) );
  XNOR2_X1 U407 ( .A(n355), .B(G148GAT), .ZN(n433) );
  XOR2_X1 U408 ( .A(G211GAT), .B(KEYINPUT21), .Z(n357) );
  XNOR2_X1 U409 ( .A(G197GAT), .B(G218GAT), .ZN(n356) );
  XNOR2_X1 U410 ( .A(n357), .B(n356), .ZN(n385) );
  XNOR2_X1 U411 ( .A(n433), .B(n385), .ZN(n358) );
  XNOR2_X1 U412 ( .A(n359), .B(n358), .ZN(n540) );
  XNOR2_X1 U413 ( .A(n361), .B(n360), .ZN(n363) );
  XNOR2_X1 U414 ( .A(G99GAT), .B(G71GAT), .ZN(n362) );
  XNOR2_X1 U415 ( .A(n362), .B(G120GAT), .ZN(n434) );
  XNOR2_X1 U416 ( .A(n363), .B(n434), .ZN(n368) );
  XOR2_X1 U417 ( .A(n364), .B(KEYINPUT84), .Z(n366) );
  NAND2_X1 U418 ( .A1(G227GAT), .A2(G233GAT), .ZN(n365) );
  XNOR2_X1 U419 ( .A(n366), .B(n365), .ZN(n367) );
  XOR2_X1 U420 ( .A(n368), .B(n367), .Z(n379) );
  XOR2_X1 U421 ( .A(G176GAT), .B(G183GAT), .Z(n370) );
  XNOR2_X1 U422 ( .A(G169GAT), .B(KEYINPUT83), .ZN(n369) );
  XNOR2_X1 U423 ( .A(n370), .B(n369), .ZN(n374) );
  XOR2_X1 U424 ( .A(KEYINPUT19), .B(KEYINPUT18), .Z(n372) );
  XNOR2_X1 U425 ( .A(G190GAT), .B(KEYINPUT17), .ZN(n371) );
  XNOR2_X1 U426 ( .A(n372), .B(n371), .ZN(n373) );
  XOR2_X1 U427 ( .A(n374), .B(n373), .Z(n384) );
  XOR2_X1 U428 ( .A(KEYINPUT85), .B(KEYINPUT82), .Z(n376) );
  XNOR2_X1 U429 ( .A(KEYINPUT20), .B(KEYINPUT81), .ZN(n375) );
  XNOR2_X1 U430 ( .A(n376), .B(n375), .ZN(n377) );
  XNOR2_X1 U431 ( .A(n384), .B(n377), .ZN(n378) );
  XNOR2_X1 U432 ( .A(n379), .B(n378), .ZN(n544) );
  INV_X1 U433 ( .A(n544), .ZN(n487) );
  NAND2_X1 U434 ( .A1(n540), .A2(n487), .ZN(n380) );
  XNOR2_X1 U435 ( .A(KEYINPUT26), .B(n380), .ZN(n566) );
  XOR2_X1 U436 ( .A(KEYINPUT96), .B(KEYINPUT95), .Z(n382) );
  XNOR2_X1 U437 ( .A(G8GAT), .B(KEYINPUT94), .ZN(n381) );
  XNOR2_X1 U438 ( .A(n382), .B(n381), .ZN(n383) );
  XNOR2_X1 U439 ( .A(n384), .B(n383), .ZN(n392) );
  XOR2_X1 U440 ( .A(KEYINPUT97), .B(n385), .Z(n387) );
  NAND2_X1 U441 ( .A1(G226GAT), .A2(G233GAT), .ZN(n386) );
  XNOR2_X1 U442 ( .A(n387), .B(n386), .ZN(n388) );
  XOR2_X1 U443 ( .A(n388), .B(G92GAT), .Z(n390) );
  XOR2_X1 U444 ( .A(G204GAT), .B(G64GAT), .Z(n440) );
  XNOR2_X1 U445 ( .A(G36GAT), .B(n440), .ZN(n389) );
  XNOR2_X1 U446 ( .A(n390), .B(n389), .ZN(n391) );
  XNOR2_X1 U447 ( .A(n392), .B(n391), .ZN(n537) );
  XNOR2_X1 U448 ( .A(n537), .B(KEYINPUT27), .ZN(n399) );
  NOR2_X1 U449 ( .A1(n566), .A2(n399), .ZN(n524) );
  NOR2_X1 U450 ( .A1(n537), .A2(n487), .ZN(n393) );
  NOR2_X1 U451 ( .A1(n540), .A2(n393), .ZN(n394) );
  XNOR2_X1 U452 ( .A(n394), .B(KEYINPUT25), .ZN(n395) );
  XNOR2_X1 U453 ( .A(KEYINPUT99), .B(n395), .ZN(n396) );
  NOR2_X1 U454 ( .A1(n524), .A2(n396), .ZN(n397) );
  XOR2_X1 U455 ( .A(KEYINPUT100), .B(n397), .Z(n398) );
  NAND2_X1 U456 ( .A1(n563), .A2(n398), .ZN(n406) );
  INV_X1 U457 ( .A(n399), .ZN(n401) );
  XNOR2_X1 U458 ( .A(n540), .B(KEYINPUT67), .ZN(n400) );
  XNOR2_X1 U459 ( .A(n400), .B(KEYINPUT28), .ZN(n490) );
  NAND2_X1 U460 ( .A1(n401), .A2(n490), .ZN(n402) );
  NOR2_X1 U461 ( .A1(n563), .A2(n402), .ZN(n511) );
  XNOR2_X1 U462 ( .A(KEYINPUT98), .B(n511), .ZN(n404) );
  XNOR2_X1 U463 ( .A(n487), .B(KEYINPUT86), .ZN(n403) );
  NAND2_X1 U464 ( .A1(n404), .A2(n403), .ZN(n405) );
  NAND2_X1 U465 ( .A1(n406), .A2(n405), .ZN(n458) );
  NAND2_X1 U466 ( .A1(n407), .A2(n458), .ZN(n472) );
  XNOR2_X1 U467 ( .A(n408), .B(KEYINPUT72), .ZN(n410) );
  INV_X1 U468 ( .A(KEYINPUT69), .ZN(n409) );
  XOR2_X1 U469 ( .A(G113GAT), .B(G43GAT), .Z(n412) );
  XNOR2_X1 U470 ( .A(G169GAT), .B(G50GAT), .ZN(n411) );
  XNOR2_X1 U471 ( .A(n412), .B(n411), .ZN(n413) );
  XNOR2_X1 U472 ( .A(n414), .B(n413), .ZN(n416) );
  AND2_X1 U473 ( .A1(G229GAT), .A2(G233GAT), .ZN(n415) );
  XNOR2_X1 U474 ( .A(n416), .B(n415), .ZN(n417) );
  XOR2_X1 U475 ( .A(G141GAT), .B(G22GAT), .Z(n420) );
  XNOR2_X1 U476 ( .A(G15GAT), .B(G197GAT), .ZN(n419) );
  XOR2_X1 U477 ( .A(n420), .B(n419), .Z(n421) );
  XNOR2_X1 U478 ( .A(n422), .B(n421), .ZN(n430) );
  XOR2_X1 U479 ( .A(KEYINPUT73), .B(KEYINPUT71), .Z(n424) );
  XNOR2_X1 U480 ( .A(KEYINPUT70), .B(KEYINPUT68), .ZN(n423) );
  XNOR2_X1 U481 ( .A(n424), .B(n423), .ZN(n428) );
  XOR2_X1 U482 ( .A(KEYINPUT74), .B(KEYINPUT29), .Z(n426) );
  XNOR2_X1 U483 ( .A(KEYINPUT75), .B(KEYINPUT30), .ZN(n425) );
  XNOR2_X1 U484 ( .A(n426), .B(n425), .ZN(n427) );
  XNOR2_X1 U485 ( .A(n428), .B(n427), .ZN(n429) );
  XNOR2_X1 U486 ( .A(n430), .B(n429), .ZN(n504) );
  XOR2_X1 U487 ( .A(n432), .B(n431), .Z(n436) );
  XNOR2_X1 U488 ( .A(n434), .B(n433), .ZN(n435) );
  XNOR2_X1 U489 ( .A(n436), .B(n435), .ZN(n444) );
  XOR2_X1 U490 ( .A(KEYINPUT32), .B(KEYINPUT33), .Z(n438) );
  XNOR2_X1 U491 ( .A(G176GAT), .B(KEYINPUT31), .ZN(n437) );
  XNOR2_X1 U492 ( .A(n438), .B(n437), .ZN(n439) );
  XOR2_X1 U493 ( .A(n440), .B(n439), .Z(n442) );
  NAND2_X1 U494 ( .A1(G230GAT), .A2(G233GAT), .ZN(n441) );
  XNOR2_X1 U495 ( .A(n442), .B(n441), .ZN(n443) );
  XNOR2_X1 U496 ( .A(n444), .B(n443), .ZN(n569) );
  NAND2_X1 U497 ( .A1(n504), .A2(n569), .ZN(n461) );
  NOR2_X1 U498 ( .A1(n472), .A2(n461), .ZN(n445) );
  XNOR2_X1 U499 ( .A(n445), .B(KEYINPUT101), .ZN(n456) );
  NOR2_X1 U500 ( .A1(n563), .A2(n456), .ZN(n447) );
  XNOR2_X1 U501 ( .A(KEYINPUT34), .B(KEYINPUT102), .ZN(n446) );
  XNOR2_X1 U502 ( .A(n447), .B(n446), .ZN(n448) );
  XOR2_X1 U503 ( .A(G1GAT), .B(n448), .Z(G1324GAT) );
  NOR2_X1 U504 ( .A1(n537), .A2(n456), .ZN(n450) );
  XNOR2_X1 U505 ( .A(KEYINPUT103), .B(KEYINPUT104), .ZN(n449) );
  XNOR2_X1 U506 ( .A(n450), .B(n449), .ZN(n451) );
  XNOR2_X1 U507 ( .A(G8GAT), .B(n451), .ZN(G1325GAT) );
  NOR2_X1 U508 ( .A1(n456), .A2(n487), .ZN(n455) );
  XOR2_X1 U509 ( .A(KEYINPUT105), .B(KEYINPUT35), .Z(n453) );
  XNOR2_X1 U510 ( .A(G15GAT), .B(KEYINPUT106), .ZN(n452) );
  XNOR2_X1 U511 ( .A(n453), .B(n452), .ZN(n454) );
  XNOR2_X1 U512 ( .A(n455), .B(n454), .ZN(G1326GAT) );
  NOR2_X1 U513 ( .A1(n490), .A2(n456), .ZN(n457) );
  XOR2_X1 U514 ( .A(G22GAT), .B(n457), .Z(G1327GAT) );
  INV_X1 U515 ( .A(n498), .ZN(n556) );
  XNOR2_X1 U516 ( .A(KEYINPUT36), .B(n556), .ZN(n577) );
  NAND2_X1 U517 ( .A1(n577), .A2(n458), .ZN(n459) );
  NOR2_X1 U518 ( .A1(n459), .A2(n574), .ZN(n460) );
  XNOR2_X1 U519 ( .A(n460), .B(KEYINPUT37), .ZN(n482) );
  NOR2_X1 U520 ( .A1(n482), .A2(n461), .ZN(n462) );
  XOR2_X1 U521 ( .A(KEYINPUT38), .B(n462), .Z(n468) );
  NOR2_X1 U522 ( .A1(n468), .A2(n563), .ZN(n463) );
  XNOR2_X1 U523 ( .A(n463), .B(KEYINPUT39), .ZN(n464) );
  XNOR2_X1 U524 ( .A(G29GAT), .B(n464), .ZN(G1328GAT) );
  NOR2_X1 U525 ( .A1(n537), .A2(n468), .ZN(n465) );
  XOR2_X1 U526 ( .A(G36GAT), .B(n465), .Z(G1329GAT) );
  NOR2_X1 U527 ( .A1(n468), .A2(n487), .ZN(n466) );
  XOR2_X1 U528 ( .A(KEYINPUT40), .B(n466), .Z(n467) );
  XNOR2_X1 U529 ( .A(G43GAT), .B(n467), .ZN(G1330GAT) );
  XNOR2_X1 U530 ( .A(G50GAT), .B(KEYINPUT107), .ZN(n470) );
  NOR2_X1 U531 ( .A1(n490), .A2(n468), .ZN(n469) );
  XNOR2_X1 U532 ( .A(n470), .B(n469), .ZN(G1331GAT) );
  INV_X1 U533 ( .A(n504), .ZN(n513) );
  XNOR2_X1 U534 ( .A(KEYINPUT41), .B(n569), .ZN(n549) );
  NAND2_X1 U535 ( .A1(n513), .A2(n549), .ZN(n471) );
  XNOR2_X1 U536 ( .A(n471), .B(KEYINPUT108), .ZN(n483) );
  NOR2_X1 U537 ( .A1(n472), .A2(n483), .ZN(n473) );
  XNOR2_X1 U538 ( .A(n473), .B(KEYINPUT109), .ZN(n479) );
  NOR2_X1 U539 ( .A1(n563), .A2(n479), .ZN(n474) );
  XOR2_X1 U540 ( .A(G57GAT), .B(n474), .Z(n475) );
  XNOR2_X1 U541 ( .A(KEYINPUT42), .B(n475), .ZN(G1332GAT) );
  NOR2_X1 U542 ( .A1(n537), .A2(n479), .ZN(n476) );
  XOR2_X1 U543 ( .A(KEYINPUT110), .B(n476), .Z(n477) );
  XNOR2_X1 U544 ( .A(G64GAT), .B(n477), .ZN(G1333GAT) );
  NOR2_X1 U545 ( .A1(n487), .A2(n479), .ZN(n478) );
  XOR2_X1 U546 ( .A(G71GAT), .B(n478), .Z(G1334GAT) );
  NOR2_X1 U547 ( .A1(n490), .A2(n479), .ZN(n481) );
  XNOR2_X1 U548 ( .A(G78GAT), .B(KEYINPUT43), .ZN(n480) );
  XNOR2_X1 U549 ( .A(n481), .B(n480), .ZN(G1335GAT) );
  OR2_X1 U550 ( .A1(n483), .A2(n482), .ZN(n489) );
  NOR2_X1 U551 ( .A1(n563), .A2(n489), .ZN(n484) );
  XOR2_X1 U552 ( .A(G85GAT), .B(n484), .Z(G1336GAT) );
  NOR2_X1 U553 ( .A1(n537), .A2(n489), .ZN(n486) );
  XNOR2_X1 U554 ( .A(G92GAT), .B(KEYINPUT111), .ZN(n485) );
  XNOR2_X1 U555 ( .A(n486), .B(n485), .ZN(G1337GAT) );
  NOR2_X1 U556 ( .A1(n487), .A2(n489), .ZN(n488) );
  XOR2_X1 U557 ( .A(G99GAT), .B(n488), .Z(G1338GAT) );
  NOR2_X1 U558 ( .A1(n490), .A2(n489), .ZN(n491) );
  XOR2_X1 U559 ( .A(KEYINPUT44), .B(n491), .Z(n492) );
  XNOR2_X1 U560 ( .A(G106GAT), .B(n492), .ZN(G1339GAT) );
  NAND2_X1 U561 ( .A1(n549), .A2(n504), .ZN(n496) );
  XOR2_X1 U562 ( .A(KEYINPUT46), .B(KEYINPUT113), .Z(n494) );
  INV_X1 U563 ( .A(KEYINPUT112), .ZN(n493) );
  NOR2_X1 U564 ( .A1(n497), .A2(n574), .ZN(n499) );
  NAND2_X1 U565 ( .A1(n499), .A2(n498), .ZN(n500) );
  XNOR2_X1 U566 ( .A(n500), .B(KEYINPUT47), .ZN(n507) );
  XOR2_X1 U567 ( .A(KEYINPUT45), .B(KEYINPUT114), .Z(n502) );
  NAND2_X1 U568 ( .A1(n574), .A2(n577), .ZN(n501) );
  XNOR2_X1 U569 ( .A(n502), .B(n501), .ZN(n503) );
  NAND2_X1 U570 ( .A1(n503), .A2(n569), .ZN(n505) );
  NOR2_X1 U571 ( .A1(n505), .A2(n504), .ZN(n506) );
  NOR2_X1 U572 ( .A1(n507), .A2(n506), .ZN(n510) );
  XOR2_X1 U573 ( .A(KEYINPUT64), .B(KEYINPUT115), .Z(n508) );
  NAND2_X1 U574 ( .A1(n544), .A2(n511), .ZN(n512) );
  NOR2_X1 U575 ( .A1(n538), .A2(n512), .ZN(n520) );
  NAND2_X1 U576 ( .A1(n520), .A2(n504), .ZN(n514) );
  XNOR2_X1 U577 ( .A(n514), .B(G113GAT), .ZN(G1340GAT) );
  XOR2_X1 U578 ( .A(G120GAT), .B(KEYINPUT49), .Z(n516) );
  NAND2_X1 U579 ( .A1(n520), .A2(n549), .ZN(n515) );
  XNOR2_X1 U580 ( .A(n516), .B(n515), .ZN(G1341GAT) );
  XOR2_X1 U581 ( .A(KEYINPUT50), .B(KEYINPUT116), .Z(n518) );
  NAND2_X1 U582 ( .A1(n520), .A2(n574), .ZN(n517) );
  XNOR2_X1 U583 ( .A(n518), .B(n517), .ZN(n519) );
  XOR2_X1 U584 ( .A(G127GAT), .B(n519), .Z(G1342GAT) );
  XOR2_X1 U585 ( .A(KEYINPUT51), .B(KEYINPUT117), .Z(n522) );
  NAND2_X1 U586 ( .A1(n520), .A2(n556), .ZN(n521) );
  XNOR2_X1 U587 ( .A(n522), .B(n521), .ZN(n523) );
  XOR2_X1 U588 ( .A(G134GAT), .B(n523), .Z(G1343GAT) );
  XOR2_X1 U589 ( .A(G141GAT), .B(KEYINPUT119), .Z(n528) );
  NOR2_X1 U590 ( .A1(n563), .A2(n538), .ZN(n525) );
  NAND2_X1 U591 ( .A1(n525), .A2(n524), .ZN(n526) );
  XOR2_X1 U592 ( .A(KEYINPUT118), .B(n526), .Z(n535) );
  NAND2_X1 U593 ( .A1(n504), .A2(n535), .ZN(n527) );
  XNOR2_X1 U594 ( .A(n528), .B(n527), .ZN(G1344GAT) );
  XOR2_X1 U595 ( .A(KEYINPUT121), .B(KEYINPUT53), .Z(n530) );
  XNOR2_X1 U596 ( .A(G148GAT), .B(KEYINPUT52), .ZN(n529) );
  XNOR2_X1 U597 ( .A(n530), .B(n529), .ZN(n531) );
  XOR2_X1 U598 ( .A(KEYINPUT120), .B(n531), .Z(n533) );
  NAND2_X1 U599 ( .A1(n549), .A2(n535), .ZN(n532) );
  XNOR2_X1 U600 ( .A(n533), .B(n532), .ZN(G1345GAT) );
  NAND2_X1 U601 ( .A1(n535), .A2(n574), .ZN(n534) );
  XNOR2_X1 U602 ( .A(n534), .B(G155GAT), .ZN(G1346GAT) );
  NAND2_X1 U603 ( .A1(n535), .A2(n556), .ZN(n536) );
  XNOR2_X1 U604 ( .A(n536), .B(G162GAT), .ZN(G1347GAT) );
  NOR2_X1 U605 ( .A1(n538), .A2(n537), .ZN(n539) );
  XNOR2_X1 U606 ( .A(KEYINPUT54), .B(n539), .ZN(n564) );
  INV_X1 U607 ( .A(n540), .ZN(n541) );
  AND2_X1 U608 ( .A1(n563), .A2(n541), .ZN(n542) );
  AND2_X1 U609 ( .A1(n564), .A2(n542), .ZN(n543) );
  XOR2_X1 U610 ( .A(KEYINPUT55), .B(n543), .Z(n545) );
  NAND2_X1 U611 ( .A1(n545), .A2(n544), .ZN(n547) );
  INV_X1 U612 ( .A(KEYINPUT122), .ZN(n546) );
  NAND2_X1 U613 ( .A1(n557), .A2(n504), .ZN(n548) );
  XNOR2_X1 U614 ( .A(n548), .B(G169GAT), .ZN(G1348GAT) );
  XOR2_X1 U615 ( .A(KEYINPUT57), .B(KEYINPUT123), .Z(n551) );
  NAND2_X1 U616 ( .A1(n549), .A2(n557), .ZN(n550) );
  XNOR2_X1 U617 ( .A(n551), .B(n550), .ZN(n553) );
  XOR2_X1 U618 ( .A(G176GAT), .B(KEYINPUT56), .Z(n552) );
  XNOR2_X1 U619 ( .A(n553), .B(n552), .ZN(G1349GAT) );
  NAND2_X1 U620 ( .A1(n557), .A2(n574), .ZN(n554) );
  XNOR2_X1 U621 ( .A(n554), .B(KEYINPUT124), .ZN(n555) );
  XNOR2_X1 U622 ( .A(G183GAT), .B(n555), .ZN(G1350GAT) );
  NAND2_X1 U623 ( .A1(n557), .A2(n556), .ZN(n558) );
  XNOR2_X1 U624 ( .A(n558), .B(KEYINPUT58), .ZN(n559) );
  XNOR2_X1 U625 ( .A(G190GAT), .B(n559), .ZN(G1351GAT) );
  XOR2_X1 U626 ( .A(KEYINPUT60), .B(KEYINPUT126), .Z(n561) );
  XNOR2_X1 U627 ( .A(G197GAT), .B(KEYINPUT59), .ZN(n560) );
  XNOR2_X1 U628 ( .A(n561), .B(n560), .ZN(n562) );
  XOR2_X1 U629 ( .A(KEYINPUT125), .B(n562), .Z(n568) );
  NAND2_X1 U630 ( .A1(n564), .A2(n563), .ZN(n565) );
  NOR2_X1 U631 ( .A1(n566), .A2(n565), .ZN(n576) );
  NAND2_X1 U632 ( .A1(n576), .A2(n504), .ZN(n567) );
  XNOR2_X1 U633 ( .A(n568), .B(n567), .ZN(G1352GAT) );
  XOR2_X1 U634 ( .A(KEYINPUT127), .B(KEYINPUT61), .Z(n572) );
  INV_X1 U635 ( .A(n569), .ZN(n570) );
  NAND2_X1 U636 ( .A1(n576), .A2(n570), .ZN(n571) );
  XNOR2_X1 U637 ( .A(n572), .B(n571), .ZN(n573) );
  XOR2_X1 U638 ( .A(G204GAT), .B(n573), .Z(G1353GAT) );
  NAND2_X1 U639 ( .A1(n574), .A2(n576), .ZN(n575) );
  XNOR2_X1 U640 ( .A(n575), .B(G211GAT), .ZN(G1354GAT) );
  NAND2_X1 U641 ( .A1(n577), .A2(n576), .ZN(n578) );
  XNOR2_X1 U642 ( .A(n578), .B(KEYINPUT62), .ZN(n579) );
  XNOR2_X1 U643 ( .A(G218GAT), .B(n579), .ZN(G1355GAT) );
endmodule

