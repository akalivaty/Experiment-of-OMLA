

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362,
         n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373,
         n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, n384,
         n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395,
         n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406,
         n407, n408, n409, n410, n411, n412, n413, n414, n415, n416, n417,
         n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, n428,
         n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, n439,
         n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450,
         n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461,
         n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472,
         n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483,
         n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494,
         n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505,
         n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516,
         n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527,
         n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538,
         n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549,
         n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560,
         n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571,
         n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582,
         n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593,
         n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604,
         n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615,
         n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626,
         n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637,
         n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648,
         n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659,
         n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670,
         n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681,
         n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692,
         n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703,
         n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714,
         n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725,
         n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736,
         n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747,
         n748, n749, n750, n751, n752, n753, n754, n755, n756, n757, n758,
         n759, n760, n761, n762, n763, n764, n765, n766, n767, n768, n769,
         n770, n771, n772, n773, n774, n775;

  AND2_X1 U373 ( .A1(n650), .A2(n774), .ZN(n370) );
  NOR2_X1 U374 ( .A1(n772), .A2(n773), .ZN(n612) );
  NOR2_X1 U375 ( .A1(n702), .A2(n701), .ZN(n611) );
  XNOR2_X1 U376 ( .A(n609), .B(n401), .ZN(n622) );
  XNOR2_X1 U377 ( .A(n519), .B(KEYINPUT16), .ZN(n460) );
  XNOR2_X1 U378 ( .A(n396), .B(KEYINPUT42), .ZN(n772) );
  NOR2_X2 U379 ( .A1(n641), .A2(n413), .ZN(n642) );
  NOR2_X1 U380 ( .A1(n623), .A2(n534), .ZN(n536) );
  XNOR2_X1 U381 ( .A(n537), .B(KEYINPUT4), .ZN(n473) );
  INV_X1 U382 ( .A(G953), .ZN(n761) );
  AND2_X1 U383 ( .A1(n434), .A2(n433), .ZN(n352) );
  XNOR2_X2 U384 ( .A(n560), .B(n559), .ZN(n583) );
  BUF_X2 U385 ( .A(n580), .Z(n404) );
  XNOR2_X2 U386 ( .A(n507), .B(n438), .ZN(n759) );
  XNOR2_X2 U387 ( .A(n473), .B(n472), .ZN(n758) );
  XNOR2_X2 U388 ( .A(n371), .B(G119), .ZN(n519) );
  XNOR2_X2 U389 ( .A(n460), .B(n357), .ZN(n753) );
  XNOR2_X2 U390 ( .A(n544), .B(n543), .ZN(n584) );
  NOR2_X1 U391 ( .A1(n687), .A2(n575), .ZN(n407) );
  AND2_X1 U392 ( .A1(n660), .A2(n592), .ZN(n593) );
  NOR2_X1 U393 ( .A1(n771), .A2(n775), .ZN(n570) );
  XNOR2_X1 U394 ( .A(n407), .B(n406), .ZN(n579) );
  NAND2_X1 U395 ( .A1(n573), .A2(n444), .ZN(n391) );
  AND2_X1 U396 ( .A1(n572), .A2(n593), .ZN(n444) );
  NAND2_X1 U397 ( .A1(n352), .A2(n431), .ZN(n562) );
  XNOR2_X1 U398 ( .A(n589), .B(KEYINPUT84), .ZN(n591) );
  XNOR2_X1 U399 ( .A(n453), .B(KEYINPUT109), .ZN(n771) );
  AND2_X1 U400 ( .A1(n616), .A2(n588), .ZN(n589) );
  NAND2_X1 U401 ( .A1(n432), .A2(n436), .ZN(n431) );
  AND2_X1 U402 ( .A1(n435), .A2(n561), .ZN(n434) );
  NOR2_X1 U403 ( .A1(n622), .A2(n716), .ZN(n396) );
  XNOR2_X1 U404 ( .A(n536), .B(n535), .ZN(n580) );
  AND2_X1 U405 ( .A1(n574), .A2(n455), .ZN(n454) );
  INV_X1 U406 ( .A(n411), .ZN(n455) );
  XNOR2_X1 U407 ( .A(n437), .B(n359), .ZN(n605) );
  NAND2_X1 U408 ( .A1(n467), .A2(n466), .ZN(n469) );
  XNOR2_X1 U409 ( .A(n392), .B(G146), .ZN(n507) );
  XNOR2_X1 U410 ( .A(G137), .B(G110), .ZN(n486) );
  INV_X1 U411 ( .A(KEYINPUT76), .ZN(n465) );
  XNOR2_X2 U412 ( .A(n481), .B(n480), .ZN(n608) );
  INV_X1 U413 ( .A(G469), .ZN(n480) );
  INV_X1 U414 ( .A(G146), .ZN(n498) );
  NAND2_X1 U415 ( .A1(n387), .A2(n354), .ZN(n385) );
  NAND2_X1 U416 ( .A1(n741), .A2(n388), .ZN(n387) );
  OR2_X1 U417 ( .A1(n736), .A2(G475), .ZN(n386) );
  BUF_X1 U418 ( .A(n507), .Z(n509) );
  NAND2_X1 U419 ( .A1(n681), .A2(KEYINPUT73), .ZN(n451) );
  XNOR2_X1 U420 ( .A(n632), .B(n395), .ZN(n698) );
  INV_X1 U421 ( .A(KEYINPUT38), .ZN(n395) );
  OR2_X1 U422 ( .A1(G237), .A2(G902), .ZN(n526) );
  XNOR2_X1 U423 ( .A(G140), .B(KEYINPUT10), .ZN(n438) );
  XNOR2_X1 U424 ( .A(G902), .B(KEYINPUT15), .ZN(n653) );
  XNOR2_X1 U425 ( .A(n608), .B(n482), .ZN(n687) );
  NAND2_X1 U426 ( .A1(n698), .A2(n699), .ZN(n702) );
  OR2_X1 U427 ( .A1(n743), .A2(G902), .ZN(n437) );
  XOR2_X1 U428 ( .A(KEYINPUT86), .B(KEYINPUT0), .Z(n535) );
  XNOR2_X1 U429 ( .A(n430), .B(n429), .ZN(n428) );
  XNOR2_X1 U430 ( .A(G101), .B(G116), .ZN(n430) );
  XNOR2_X1 U431 ( .A(KEYINPUT72), .B(KEYINPUT5), .ZN(n429) );
  XNOR2_X1 U432 ( .A(n488), .B(KEYINPUT24), .ZN(n489) );
  XNOR2_X1 U433 ( .A(n408), .B(n487), .ZN(n488) );
  XOR2_X1 U434 ( .A(KEYINPUT23), .B(KEYINPUT96), .Z(n487) );
  XNOR2_X1 U435 ( .A(n486), .B(KEYINPUT81), .ZN(n408) );
  INV_X1 U436 ( .A(G134), .ZN(n470) );
  XNOR2_X1 U437 ( .A(G122), .B(G116), .ZN(n459) );
  XNOR2_X1 U438 ( .A(KEYINPUT87), .B(KEYINPUT33), .ZN(n502) );
  NAND2_X1 U439 ( .A1(n374), .A2(n373), .ZN(n419) );
  NAND2_X1 U440 ( .A1(n601), .A2(n602), .ZN(n424) );
  INV_X1 U441 ( .A(KEYINPUT106), .ZN(n412) );
  OR2_X1 U442 ( .A1(n659), .A2(G902), .ZN(n442) );
  NAND2_X1 U443 ( .A1(n385), .A2(n389), .ZN(n383) );
  NOR2_X1 U444 ( .A1(n736), .A2(KEYINPUT60), .ZN(n382) );
  AND2_X1 U445 ( .A1(n378), .A2(KEYINPUT60), .ZN(n377) );
  XNOR2_X1 U446 ( .A(n758), .B(n479), .ZN(n729) );
  XNOR2_X1 U447 ( .A(n476), .B(n498), .ZN(n478) );
  NAND2_X1 U448 ( .A1(n741), .A2(G210), .ZN(n441) );
  INV_X1 U449 ( .A(G125), .ZN(n392) );
  XNOR2_X1 U450 ( .A(G104), .B(G122), .ZN(n549) );
  XNOR2_X1 U451 ( .A(G143), .B(G113), .ZN(n545) );
  NOR2_X1 U452 ( .A1(KEYINPUT73), .A2(n447), .ZN(n446) );
  INV_X1 U453 ( .A(n451), .ZN(n447) );
  NOR2_X1 U454 ( .A1(n353), .A2(n653), .ZN(n449) );
  NAND2_X1 U455 ( .A1(G234), .A2(G237), .ZN(n528) );
  INV_X1 U456 ( .A(KEYINPUT71), .ZN(n406) );
  XNOR2_X1 U457 ( .A(n525), .B(n523), .ZN(n461) );
  XNOR2_X1 U458 ( .A(n594), .B(KEYINPUT113), .ZN(n375) );
  XNOR2_X1 U459 ( .A(G101), .B(G110), .ZN(n477) );
  XOR2_X1 U460 ( .A(G107), .B(G140), .Z(n475) );
  INV_X1 U461 ( .A(n681), .ZN(n415) );
  INV_X1 U462 ( .A(KEYINPUT116), .ZN(n403) );
  NOR2_X1 U463 ( .A1(n404), .A2(KEYINPUT34), .ZN(n436) );
  XNOR2_X1 U464 ( .A(n410), .B(KEYINPUT22), .ZN(n372) );
  NOR2_X1 U465 ( .A1(n580), .A2(n567), .ZN(n410) );
  AND2_X1 U466 ( .A1(n590), .A2(n399), .ZN(n398) );
  INV_X1 U467 ( .A(n699), .ZN(n417) );
  NAND2_X1 U468 ( .A1(n375), .A2(n603), .ZN(n631) );
  INV_X1 U469 ( .A(KEYINPUT115), .ZN(n401) );
  BUF_X1 U470 ( .A(n605), .Z(n411) );
  XNOR2_X1 U471 ( .A(n558), .B(n557), .ZN(n559) );
  INV_X1 U472 ( .A(G475), .ZN(n557) );
  BUF_X1 U473 ( .A(n691), .Z(n400) );
  AND2_X1 U474 ( .A1(n372), .A2(n397), .ZN(n588) );
  INV_X1 U475 ( .A(KEYINPUT6), .ZN(n402) );
  XNOR2_X1 U476 ( .A(n758), .B(n443), .ZN(n659) );
  XNOR2_X1 U477 ( .A(n499), .B(n498), .ZN(n443) );
  XNOR2_X1 U478 ( .A(n428), .B(n497), .ZN(n427) );
  NAND2_X1 U479 ( .A1(n741), .A2(G472), .ZN(n458) );
  XNOR2_X1 U480 ( .A(n409), .B(n494), .ZN(n743) );
  XNOR2_X1 U481 ( .A(n489), .B(n490), .ZN(n409) );
  XOR2_X1 U482 ( .A(G128), .B(G119), .Z(n492) );
  XOR2_X1 U483 ( .A(KEYINPUT7), .B(KEYINPUT9), .Z(n540) );
  XNOR2_X1 U484 ( .A(n426), .B(n425), .ZN(n773) );
  INV_X1 U485 ( .A(KEYINPUT40), .ZN(n425) );
  NAND2_X1 U486 ( .A1(n379), .A2(n377), .ZN(n376) );
  AND2_X1 U487 ( .A1(n383), .A2(n381), .ZN(n380) );
  INV_X1 U488 ( .A(n385), .ZN(n379) );
  XNOR2_X1 U489 ( .A(n731), .B(n730), .ZN(n732) );
  XNOR2_X1 U490 ( .A(n729), .B(n463), .ZN(n730) );
  INV_X1 U491 ( .A(KEYINPUT56), .ZN(n439) );
  OR2_X1 U492 ( .A1(n681), .A2(KEYINPUT73), .ZN(n353) );
  AND2_X1 U493 ( .A1(n386), .A2(n390), .ZN(n354) );
  XOR2_X1 U494 ( .A(KEYINPUT75), .B(n616), .Z(n355) );
  AND2_X1 U495 ( .A1(n774), .A2(n451), .ZN(n356) );
  XOR2_X1 U496 ( .A(n459), .B(G107), .Z(n357) );
  AND2_X1 U497 ( .A1(n419), .A2(n424), .ZN(n358) );
  XOR2_X1 U498 ( .A(n496), .B(KEYINPUT25), .Z(n359) );
  XOR2_X1 U499 ( .A(n514), .B(KEYINPUT91), .Z(n360) );
  AND2_X1 U500 ( .A1(n420), .A2(n603), .ZN(n361) );
  NOR2_X1 U501 ( .A1(n616), .A2(n394), .ZN(n362) );
  BUF_X1 U502 ( .A(n687), .Z(n397) );
  AND2_X1 U503 ( .A1(n424), .A2(n423), .ZN(n363) );
  AND2_X1 U504 ( .A1(n355), .A2(n398), .ZN(n364) );
  XOR2_X1 U505 ( .A(KEYINPUT45), .B(KEYINPUT65), .Z(n365) );
  XNOR2_X1 U506 ( .A(n726), .B(n725), .ZN(n366) );
  XOR2_X1 U507 ( .A(n659), .B(KEYINPUT62), .Z(n367) );
  INV_X1 U508 ( .A(n736), .ZN(n737) );
  INV_X1 U509 ( .A(KEYINPUT60), .ZN(n389) );
  NOR2_X1 U510 ( .A1(G952), .A2(n761), .ZN(n745) );
  INV_X1 U511 ( .A(n745), .ZN(n390) );
  NAND2_X1 U512 ( .A1(n368), .A2(n608), .ZN(n609) );
  XNOR2_X1 U513 ( .A(n606), .B(n607), .ZN(n368) );
  NAND2_X1 U514 ( .A1(n450), .A2(n369), .ZN(n452) );
  NAND2_X1 U515 ( .A1(n370), .A2(n449), .ZN(n369) );
  XNOR2_X1 U516 ( .A(n416), .B(KEYINPUT30), .ZN(n600) );
  XNOR2_X1 U517 ( .A(n441), .B(n366), .ZN(n440) );
  XNOR2_X1 U518 ( .A(n458), .B(n367), .ZN(n457) );
  NAND2_X1 U519 ( .A1(n691), .A2(n615), .ZN(n606) );
  NAND2_X1 U520 ( .A1(n650), .A2(n356), .ZN(n448) );
  AND2_X1 U521 ( .A1(n370), .A2(n415), .ZN(n760) );
  XNOR2_X2 U522 ( .A(G113), .B(KEYINPUT3), .ZN(n371) );
  AND2_X1 U523 ( .A1(n372), .A2(n364), .ZN(n568) );
  NAND2_X1 U524 ( .A1(n420), .A2(KEYINPUT39), .ZN(n373) );
  NAND2_X1 U525 ( .A1(n375), .A2(n361), .ZN(n374) );
  NAND2_X1 U526 ( .A1(n631), .A2(n602), .ZN(n423) );
  NAND2_X1 U527 ( .A1(n380), .A2(n376), .ZN(G60) );
  NAND2_X1 U528 ( .A1(n384), .A2(n737), .ZN(n378) );
  NAND2_X1 U529 ( .A1(n384), .A2(n382), .ZN(n381) );
  INV_X1 U530 ( .A(n741), .ZN(n384) );
  AND2_X1 U531 ( .A1(n736), .A2(G475), .ZN(n388) );
  NOR2_X1 U532 ( .A1(n446), .A2(n653), .ZN(n445) );
  NAND2_X1 U533 ( .A1(n421), .A2(n422), .ZN(n418) );
  INV_X1 U534 ( .A(n574), .ZN(n691) );
  XNOR2_X2 U535 ( .A(n391), .B(n365), .ZN(n748) );
  NAND2_X1 U536 ( .A1(n576), .A2(n608), .ZN(n594) );
  XNOR2_X1 U537 ( .A(n393), .B(n555), .ZN(n733) );
  XNOR2_X1 U538 ( .A(n554), .B(n556), .ZN(n393) );
  NAND2_X1 U539 ( .A1(n358), .A2(n418), .ZN(n426) );
  AND2_X1 U540 ( .A1(n670), .A2(n362), .ZN(n643) );
  INV_X1 U541 ( .A(n615), .ZN(n394) );
  NAND2_X1 U542 ( .A1(n591), .A2(n684), .ZN(n660) );
  NAND2_X1 U543 ( .A1(n656), .A2(n655), .ZN(n658) );
  NOR2_X1 U544 ( .A1(KEYINPUT44), .A2(n564), .ZN(n569) );
  NAND2_X1 U545 ( .A1(n588), .A2(n454), .ZN(n453) );
  INV_X1 U546 ( .A(n397), .ZN(n399) );
  XNOR2_X1 U547 ( .A(n574), .B(n402), .ZN(n616) );
  XNOR2_X2 U548 ( .A(n442), .B(n500), .ZN(n574) );
  XNOR2_X1 U549 ( .A(n643), .B(n403), .ZN(n617) );
  XNOR2_X1 U550 ( .A(n515), .B(n360), .ZN(n518) );
  NAND2_X1 U551 ( .A1(n405), .A2(KEYINPUT44), .ZN(n572) );
  NAND2_X1 U552 ( .A1(n570), .A2(n571), .ZN(n405) );
  XNOR2_X2 U553 ( .A(n585), .B(n412), .ZN(n614) );
  NAND2_X1 U554 ( .A1(n457), .A2(n390), .ZN(n456) );
  NAND2_X1 U555 ( .A1(n639), .A2(n640), .ZN(n413) );
  XNOR2_X1 U556 ( .A(n414), .B(n439), .ZN(G51) );
  NAND2_X1 U557 ( .A1(n440), .A2(n390), .ZN(n414) );
  NOR2_X2 U558 ( .A1(n623), .A2(n622), .ZN(n671) );
  NAND2_X1 U559 ( .A1(n632), .A2(n699), .ZN(n613) );
  INV_X1 U560 ( .A(n600), .ZN(n630) );
  NOR2_X1 U561 ( .A1(n574), .A2(n417), .ZN(n416) );
  NAND2_X1 U562 ( .A1(n418), .A2(n363), .ZN(n651) );
  INV_X1 U563 ( .A(n614), .ZN(n420) );
  NOR2_X1 U564 ( .A1(n631), .A2(n602), .ZN(n421) );
  INV_X1 U565 ( .A(n601), .ZN(n422) );
  XNOR2_X1 U566 ( .A(n519), .B(n427), .ZN(n499) );
  INV_X1 U567 ( .A(n707), .ZN(n432) );
  NAND2_X1 U568 ( .A1(n707), .A2(KEYINPUT34), .ZN(n433) );
  NAND2_X1 U569 ( .A1(n404), .A2(KEYINPUT34), .ZN(n435) );
  XNOR2_X2 U570 ( .A(n503), .B(n502), .ZN(n707) );
  NOR2_X2 U571 ( .A1(n584), .A2(n583), .ZN(n585) );
  NAND2_X1 U572 ( .A1(n448), .A2(n445), .ZN(n450) );
  NAND2_X1 U573 ( .A1(n452), .A2(n748), .ZN(n652) );
  XNOR2_X1 U574 ( .A(n456), .B(KEYINPUT63), .ZN(G57) );
  XNOR2_X2 U575 ( .A(n613), .B(n527), .ZN(n623) );
  XNOR2_X2 U576 ( .A(n524), .B(n461), .ZN(n632) );
  AND2_X4 U577 ( .A1(n658), .A2(n657), .ZN(n741) );
  INV_X1 U578 ( .A(n404), .ZN(n578) );
  XNOR2_X1 U579 ( .A(KEYINPUT64), .B(KEYINPUT46), .ZN(n462) );
  XOR2_X1 U580 ( .A(n728), .B(n727), .Z(n463) );
  INV_X1 U581 ( .A(KEYINPUT67), .ZN(n563) );
  INV_X1 U582 ( .A(G143), .ZN(n468) );
  XNOR2_X1 U583 ( .A(n753), .B(n520), .ZN(n521) );
  INV_X1 U584 ( .A(KEYINPUT1), .ZN(n482) );
  INV_X1 U585 ( .A(KEYINPUT19), .ZN(n527) );
  XNOR2_X1 U586 ( .A(n493), .B(n492), .ZN(n494) );
  INV_X1 U587 ( .A(KEYINPUT39), .ZN(n602) );
  INV_X1 U588 ( .A(G128), .ZN(n464) );
  NAND2_X1 U589 ( .A1(n464), .A2(KEYINPUT76), .ZN(n467) );
  NAND2_X1 U590 ( .A1(n465), .A2(G128), .ZN(n466) );
  XNOR2_X2 U591 ( .A(n469), .B(n468), .ZN(n516) );
  XNOR2_X2 U592 ( .A(n516), .B(n470), .ZN(n537) );
  XNOR2_X1 U593 ( .A(G131), .B(KEYINPUT69), .ZN(n471) );
  XNOR2_X1 U594 ( .A(n471), .B(KEYINPUT68), .ZN(n553) );
  XOR2_X1 U595 ( .A(n553), .B(G137), .Z(n472) );
  NAND2_X1 U596 ( .A1(G227), .A2(n761), .ZN(n474) );
  XNOR2_X1 U597 ( .A(n475), .B(n474), .ZN(n476) );
  XNOR2_X1 U598 ( .A(n477), .B(G104), .ZN(n751) );
  XNOR2_X1 U599 ( .A(KEYINPUT70), .B(n751), .ZN(n520) );
  XNOR2_X1 U600 ( .A(n478), .B(n520), .ZN(n479) );
  NOR2_X1 U601 ( .A1(n729), .A2(G902), .ZN(n481) );
  NAND2_X1 U602 ( .A1(G234), .A2(n653), .ZN(n483) );
  XNOR2_X1 U603 ( .A(KEYINPUT20), .B(n483), .ZN(n495) );
  NAND2_X1 U604 ( .A1(n495), .A2(G221), .ZN(n484) );
  XOR2_X1 U605 ( .A(KEYINPUT21), .B(n484), .Z(n683) );
  XNOR2_X1 U606 ( .A(KEYINPUT98), .B(n683), .ZN(n566) );
  INV_X1 U607 ( .A(KEYINPUT97), .ZN(n485) );
  XNOR2_X1 U608 ( .A(n759), .B(n485), .ZN(n490) );
  NAND2_X1 U609 ( .A1(G234), .A2(n761), .ZN(n491) );
  XOR2_X1 U610 ( .A(KEYINPUT8), .B(n491), .Z(n538) );
  NAND2_X1 U611 ( .A1(n538), .A2(G221), .ZN(n493) );
  NAND2_X1 U612 ( .A1(G217), .A2(n495), .ZN(n496) );
  NAND2_X1 U613 ( .A1(n566), .A2(n605), .ZN(n575) );
  NOR2_X1 U614 ( .A1(G953), .A2(G237), .ZN(n546) );
  NAND2_X1 U615 ( .A1(n546), .A2(G210), .ZN(n497) );
  XNOR2_X1 U616 ( .A(G472), .B(KEYINPUT99), .ZN(n500) );
  INV_X1 U617 ( .A(n616), .ZN(n501) );
  NAND2_X1 U618 ( .A1(n579), .A2(n501), .ZN(n503) );
  XNOR2_X1 U619 ( .A(KEYINPUT92), .B(KEYINPUT93), .ZN(n504) );
  XNOR2_X1 U620 ( .A(n504), .B(KEYINPUT77), .ZN(n525) );
  XOR2_X1 U621 ( .A(KEYINPUT90), .B(KEYINPUT17), .Z(n506) );
  XNOR2_X1 U622 ( .A(KEYINPUT4), .B(KEYINPUT89), .ZN(n505) );
  XNOR2_X1 U623 ( .A(n506), .B(n505), .ZN(n510) );
  INV_X1 U624 ( .A(n510), .ZN(n508) );
  NAND2_X1 U625 ( .A1(n508), .A2(n509), .ZN(n513) );
  INV_X1 U626 ( .A(n509), .ZN(n511) );
  NAND2_X1 U627 ( .A1(n511), .A2(n510), .ZN(n512) );
  NAND2_X1 U628 ( .A1(n513), .A2(n512), .ZN(n515) );
  NAND2_X1 U629 ( .A1(G224), .A2(n761), .ZN(n514) );
  XNOR2_X1 U630 ( .A(n516), .B(KEYINPUT18), .ZN(n517) );
  XNOR2_X1 U631 ( .A(n518), .B(n517), .ZN(n522) );
  XNOR2_X1 U632 ( .A(n521), .B(n522), .ZN(n726) );
  NAND2_X1 U633 ( .A1(n726), .A2(n653), .ZN(n524) );
  AND2_X1 U634 ( .A1(G210), .A2(n526), .ZN(n523) );
  NAND2_X1 U635 ( .A1(G214), .A2(n526), .ZN(n699) );
  XNOR2_X1 U636 ( .A(n528), .B(KEYINPUT14), .ZN(n531) );
  NAND2_X1 U637 ( .A1(G952), .A2(n531), .ZN(n714) );
  NOR2_X1 U638 ( .A1(n714), .A2(G953), .ZN(n529) );
  XOR2_X1 U639 ( .A(n529), .B(KEYINPUT94), .Z(n597) );
  INV_X1 U640 ( .A(n597), .ZN(n533) );
  NOR2_X1 U641 ( .A1(G898), .A2(n761), .ZN(n530) );
  XNOR2_X1 U642 ( .A(KEYINPUT95), .B(n530), .ZN(n755) );
  NAND2_X1 U643 ( .A1(G902), .A2(n531), .ZN(n595) );
  NOR2_X1 U644 ( .A1(n755), .A2(n595), .ZN(n532) );
  NOR2_X1 U645 ( .A1(n533), .A2(n532), .ZN(n534) );
  XNOR2_X1 U646 ( .A(KEYINPUT105), .B(G478), .ZN(n544) );
  XOR2_X1 U647 ( .A(n537), .B(n357), .Z(n542) );
  NAND2_X1 U648 ( .A1(G217), .A2(n538), .ZN(n539) );
  XNOR2_X1 U649 ( .A(n540), .B(n539), .ZN(n541) );
  XNOR2_X1 U650 ( .A(n542), .B(n541), .ZN(n739) );
  NOR2_X1 U651 ( .A1(G902), .A2(n739), .ZN(n543) );
  XNOR2_X1 U652 ( .A(n545), .B(KEYINPUT11), .ZN(n556) );
  XOR2_X1 U653 ( .A(KEYINPUT12), .B(KEYINPUT103), .Z(n548) );
  NAND2_X1 U654 ( .A1(G214), .A2(n546), .ZN(n547) );
  XNOR2_X1 U655 ( .A(n547), .B(n548), .ZN(n552) );
  XOR2_X1 U656 ( .A(KEYINPUT101), .B(KEYINPUT102), .Z(n550) );
  XNOR2_X1 U657 ( .A(n550), .B(n549), .ZN(n551) );
  XOR2_X1 U658 ( .A(n552), .B(n551), .Z(n555) );
  XNOR2_X1 U659 ( .A(n553), .B(n759), .ZN(n554) );
  NOR2_X1 U660 ( .A1(G902), .A2(n733), .ZN(n560) );
  XNOR2_X1 U661 ( .A(KEYINPUT104), .B(KEYINPUT13), .ZN(n558) );
  INV_X1 U662 ( .A(n583), .ZN(n565) );
  NAND2_X1 U663 ( .A1(n584), .A2(n565), .ZN(n633) );
  XOR2_X1 U664 ( .A(KEYINPUT74), .B(n633), .Z(n561) );
  XNOR2_X2 U665 ( .A(n562), .B(KEYINPUT35), .ZN(n769) );
  XNOR2_X1 U666 ( .A(n769), .B(n563), .ZN(n564) );
  NOR2_X1 U667 ( .A1(n584), .A2(n565), .ZN(n610) );
  NAND2_X1 U668 ( .A1(n566), .A2(n610), .ZN(n567) );
  XOR2_X1 U669 ( .A(KEYINPUT108), .B(n411), .Z(n590) );
  XNOR2_X1 U670 ( .A(n568), .B(KEYINPUT32), .ZN(n775) );
  NAND2_X1 U671 ( .A1(n569), .A2(n570), .ZN(n573) );
  NOR2_X1 U672 ( .A1(n769), .A2(KEYINPUT67), .ZN(n571) );
  INV_X1 U673 ( .A(n575), .ZN(n576) );
  NOR2_X1 U674 ( .A1(n400), .A2(n594), .ZN(n577) );
  NAND2_X1 U675 ( .A1(n578), .A2(n577), .ZN(n662) );
  NAND2_X1 U676 ( .A1(n400), .A2(n579), .ZN(n695) );
  NOR2_X1 U677 ( .A1(n404), .A2(n695), .ZN(n582) );
  XNOR2_X1 U678 ( .A(KEYINPUT31), .B(KEYINPUT100), .ZN(n581) );
  XNOR2_X1 U679 ( .A(n582), .B(n581), .ZN(n677) );
  NAND2_X1 U680 ( .A1(n662), .A2(n677), .ZN(n587) );
  NAND2_X1 U681 ( .A1(n584), .A2(n583), .ZN(n676) );
  NAND2_X1 U682 ( .A1(n676), .A2(n614), .ZN(n586) );
  XNOR2_X1 U683 ( .A(KEYINPUT107), .B(n586), .ZN(n703) );
  INV_X1 U684 ( .A(n703), .ZN(n626) );
  NAND2_X1 U685 ( .A1(n587), .A2(n626), .ZN(n592) );
  INV_X1 U686 ( .A(n590), .ZN(n684) );
  NOR2_X1 U687 ( .A1(G900), .A2(n595), .ZN(n596) );
  NAND2_X1 U688 ( .A1(n596), .A2(G953), .ZN(n598) );
  NAND2_X1 U689 ( .A1(n598), .A2(n597), .ZN(n599) );
  XNOR2_X1 U690 ( .A(n599), .B(KEYINPUT78), .ZN(n603) );
  NAND2_X1 U691 ( .A1(n698), .A2(n600), .ZN(n601) );
  XOR2_X1 U692 ( .A(KEYINPUT114), .B(KEYINPUT28), .Z(n607) );
  NAND2_X1 U693 ( .A1(n603), .A2(n683), .ZN(n604) );
  NOR2_X1 U694 ( .A1(n605), .A2(n604), .ZN(n615) );
  INV_X1 U695 ( .A(n610), .ZN(n701) );
  XNOR2_X1 U696 ( .A(n611), .B(KEYINPUT41), .ZN(n716) );
  XNOR2_X1 U697 ( .A(n612), .B(n462), .ZN(n621) );
  BUF_X1 U698 ( .A(n613), .Z(n618) );
  XOR2_X1 U699 ( .A(KEYINPUT110), .B(n614), .Z(n670) );
  NOR2_X1 U700 ( .A1(n618), .A2(n617), .ZN(n619) );
  XNOR2_X1 U701 ( .A(n619), .B(KEYINPUT36), .ZN(n620) );
  NAND2_X1 U702 ( .A1(n620), .A2(n399), .ZN(n680) );
  NAND2_X1 U703 ( .A1(n621), .A2(n680), .ZN(n641) );
  INV_X1 U704 ( .A(KEYINPUT47), .ZN(n624) );
  NAND2_X1 U705 ( .A1(n671), .A2(n624), .ZN(n625) );
  NAND2_X1 U706 ( .A1(n625), .A2(KEYINPUT80), .ZN(n627) );
  NAND2_X1 U707 ( .A1(n627), .A2(n626), .ZN(n640) );
  NAND2_X1 U708 ( .A1(n703), .A2(KEYINPUT80), .ZN(n628) );
  NAND2_X1 U709 ( .A1(n628), .A2(n671), .ZN(n629) );
  NAND2_X1 U710 ( .A1(n629), .A2(KEYINPUT47), .ZN(n636) );
  NOR2_X1 U711 ( .A1(n631), .A2(n630), .ZN(n635) );
  INV_X1 U712 ( .A(n632), .ZN(n647) );
  NOR2_X1 U713 ( .A1(n647), .A2(n633), .ZN(n634) );
  NAND2_X1 U714 ( .A1(n635), .A2(n634), .ZN(n669) );
  NAND2_X1 U715 ( .A1(n636), .A2(n669), .ZN(n638) );
  NOR2_X1 U716 ( .A1(KEYINPUT47), .A2(KEYINPUT80), .ZN(n637) );
  NOR2_X1 U717 ( .A1(n638), .A2(n637), .ZN(n639) );
  XNOR2_X1 U718 ( .A(n642), .B(KEYINPUT48), .ZN(n650) );
  NAND2_X1 U719 ( .A1(n643), .A2(n699), .ZN(n644) );
  XNOR2_X1 U720 ( .A(KEYINPUT111), .B(n644), .ZN(n645) );
  NAND2_X1 U721 ( .A1(n645), .A2(n397), .ZN(n646) );
  XNOR2_X1 U722 ( .A(KEYINPUT43), .B(n646), .ZN(n648) );
  NAND2_X1 U723 ( .A1(n648), .A2(n647), .ZN(n649) );
  XNOR2_X1 U724 ( .A(KEYINPUT112), .B(n649), .ZN(n774) );
  NOR2_X1 U725 ( .A1(n676), .A2(n651), .ZN(n681) );
  XNOR2_X1 U726 ( .A(n652), .B(KEYINPUT82), .ZN(n656) );
  XNOR2_X1 U727 ( .A(KEYINPUT83), .B(n653), .ZN(n654) );
  NAND2_X1 U728 ( .A1(n654), .A2(KEYINPUT2), .ZN(n655) );
  AND2_X1 U729 ( .A1(n748), .A2(n760), .ZN(n682) );
  NAND2_X1 U730 ( .A1(KEYINPUT2), .A2(n682), .ZN(n657) );
  XNOR2_X1 U731 ( .A(G101), .B(n660), .ZN(G3) );
  INV_X1 U732 ( .A(n670), .ZN(n674) );
  NOR2_X1 U733 ( .A1(n662), .A2(n674), .ZN(n661) );
  XOR2_X1 U734 ( .A(G104), .B(n661), .Z(G6) );
  NOR2_X1 U735 ( .A1(n676), .A2(n662), .ZN(n664) );
  XNOR2_X1 U736 ( .A(KEYINPUT27), .B(KEYINPUT26), .ZN(n663) );
  XNOR2_X1 U737 ( .A(n664), .B(n663), .ZN(n665) );
  XNOR2_X1 U738 ( .A(G107), .B(n665), .ZN(G9) );
  XOR2_X1 U739 ( .A(G128), .B(KEYINPUT29), .Z(n668) );
  INV_X1 U740 ( .A(n676), .ZN(n666) );
  NAND2_X1 U741 ( .A1(n671), .A2(n666), .ZN(n667) );
  XNOR2_X1 U742 ( .A(n668), .B(n667), .ZN(G30) );
  XNOR2_X1 U743 ( .A(G143), .B(n669), .ZN(G45) );
  XOR2_X1 U744 ( .A(G146), .B(KEYINPUT117), .Z(n673) );
  NAND2_X1 U745 ( .A1(n671), .A2(n670), .ZN(n672) );
  XNOR2_X1 U746 ( .A(n673), .B(n672), .ZN(G48) );
  NOR2_X1 U747 ( .A1(n677), .A2(n674), .ZN(n675) );
  XOR2_X1 U748 ( .A(G113), .B(n675), .Z(G15) );
  NOR2_X1 U749 ( .A1(n677), .A2(n676), .ZN(n678) );
  XOR2_X1 U750 ( .A(G116), .B(n678), .Z(G18) );
  XOR2_X1 U751 ( .A(G125), .B(KEYINPUT37), .Z(n679) );
  XNOR2_X1 U752 ( .A(n680), .B(n679), .ZN(G27) );
  XOR2_X1 U753 ( .A(G134), .B(n681), .Z(G36) );
  XNOR2_X1 U754 ( .A(KEYINPUT2), .B(n682), .ZN(n720) );
  NOR2_X1 U755 ( .A1(n684), .A2(n683), .ZN(n686) );
  XNOR2_X1 U756 ( .A(KEYINPUT49), .B(KEYINPUT118), .ZN(n685) );
  XNOR2_X1 U757 ( .A(n686), .B(n685), .ZN(n693) );
  NAND2_X1 U758 ( .A1(n575), .A2(n397), .ZN(n688) );
  XNOR2_X1 U759 ( .A(n688), .B(KEYINPUT119), .ZN(n689) );
  XNOR2_X1 U760 ( .A(KEYINPUT50), .B(n689), .ZN(n690) );
  NOR2_X1 U761 ( .A1(n400), .A2(n690), .ZN(n692) );
  NAND2_X1 U762 ( .A1(n693), .A2(n692), .ZN(n694) );
  NAND2_X1 U763 ( .A1(n695), .A2(n694), .ZN(n696) );
  XNOR2_X1 U764 ( .A(KEYINPUT51), .B(n696), .ZN(n697) );
  NOR2_X1 U765 ( .A1(n716), .A2(n697), .ZN(n710) );
  NOR2_X1 U766 ( .A1(n699), .A2(n698), .ZN(n700) );
  NOR2_X1 U767 ( .A1(n701), .A2(n700), .ZN(n706) );
  NOR2_X1 U768 ( .A1(n703), .A2(n702), .ZN(n704) );
  XNOR2_X1 U769 ( .A(n704), .B(KEYINPUT120), .ZN(n705) );
  NOR2_X1 U770 ( .A1(n706), .A2(n705), .ZN(n708) );
  NOR2_X1 U771 ( .A1(n708), .A2(n707), .ZN(n709) );
  NOR2_X1 U772 ( .A1(n710), .A2(n709), .ZN(n711) );
  XOR2_X1 U773 ( .A(n711), .B(KEYINPUT121), .Z(n712) );
  XNOR2_X1 U774 ( .A(KEYINPUT52), .B(n712), .ZN(n713) );
  NOR2_X1 U775 ( .A1(n714), .A2(n713), .ZN(n715) );
  XNOR2_X1 U776 ( .A(n715), .B(KEYINPUT122), .ZN(n718) );
  NOR2_X1 U777 ( .A1(n707), .A2(n716), .ZN(n717) );
  NOR2_X1 U778 ( .A1(n718), .A2(n717), .ZN(n719) );
  NAND2_X1 U779 ( .A1(n720), .A2(n719), .ZN(n721) );
  NOR2_X1 U780 ( .A1(n721), .A2(G953), .ZN(n722) );
  XNOR2_X1 U781 ( .A(n722), .B(KEYINPUT53), .ZN(G75) );
  XOR2_X1 U782 ( .A(KEYINPUT79), .B(KEYINPUT85), .Z(n724) );
  XNOR2_X1 U783 ( .A(KEYINPUT55), .B(KEYINPUT54), .ZN(n723) );
  XNOR2_X1 U784 ( .A(n724), .B(n723), .ZN(n725) );
  NAND2_X1 U785 ( .A1(n741), .A2(G469), .ZN(n731) );
  XOR2_X1 U786 ( .A(KEYINPUT123), .B(KEYINPUT124), .Z(n728) );
  XNOR2_X1 U787 ( .A(KEYINPUT58), .B(KEYINPUT57), .ZN(n727) );
  NOR2_X1 U788 ( .A1(n745), .A2(n732), .ZN(G54) );
  XNOR2_X1 U789 ( .A(KEYINPUT66), .B(KEYINPUT59), .ZN(n735) );
  XNOR2_X1 U790 ( .A(n733), .B(KEYINPUT88), .ZN(n734) );
  XNOR2_X1 U791 ( .A(n735), .B(n734), .ZN(n736) );
  NAND2_X1 U792 ( .A1(G478), .A2(n741), .ZN(n738) );
  XNOR2_X1 U793 ( .A(n739), .B(n738), .ZN(n740) );
  NOR2_X1 U794 ( .A1(n745), .A2(n740), .ZN(G63) );
  NAND2_X1 U795 ( .A1(G217), .A2(n741), .ZN(n742) );
  XNOR2_X1 U796 ( .A(n743), .B(n742), .ZN(n744) );
  NOR2_X1 U797 ( .A1(n745), .A2(n744), .ZN(G66) );
  NAND2_X1 U798 ( .A1(G953), .A2(G224), .ZN(n746) );
  XNOR2_X1 U799 ( .A(KEYINPUT61), .B(n746), .ZN(n747) );
  NAND2_X1 U800 ( .A1(n747), .A2(G898), .ZN(n750) );
  NAND2_X1 U801 ( .A1(n748), .A2(n761), .ZN(n749) );
  NAND2_X1 U802 ( .A1(n750), .A2(n749), .ZN(n757) );
  XOR2_X1 U803 ( .A(n751), .B(KEYINPUT125), .Z(n752) );
  XNOR2_X1 U804 ( .A(n753), .B(n752), .ZN(n754) );
  NAND2_X1 U805 ( .A1(n755), .A2(n754), .ZN(n756) );
  XOR2_X1 U806 ( .A(n757), .B(n756), .Z(G69) );
  XOR2_X1 U807 ( .A(n758), .B(n759), .Z(n764) );
  XOR2_X1 U808 ( .A(n764), .B(n760), .Z(n762) );
  NAND2_X1 U809 ( .A1(n762), .A2(n761), .ZN(n763) );
  XNOR2_X1 U810 ( .A(n763), .B(KEYINPUT126), .ZN(n768) );
  XNOR2_X1 U811 ( .A(G227), .B(n764), .ZN(n765) );
  NAND2_X1 U812 ( .A1(n765), .A2(G900), .ZN(n766) );
  NAND2_X1 U813 ( .A1(n766), .A2(G953), .ZN(n767) );
  NAND2_X1 U814 ( .A1(n768), .A2(n767), .ZN(G72) );
  XNOR2_X1 U815 ( .A(n769), .B(G122), .ZN(n770) );
  XNOR2_X1 U816 ( .A(n770), .B(KEYINPUT127), .ZN(G24) );
  XOR2_X1 U817 ( .A(n771), .B(G110), .Z(G12) );
  XOR2_X1 U818 ( .A(n772), .B(G137), .Z(G39) );
  XOR2_X1 U819 ( .A(n773), .B(G131), .Z(G33) );
  XNOR2_X1 U820 ( .A(G140), .B(n774), .ZN(G42) );
  XOR2_X1 U821 ( .A(G119), .B(n775), .Z(G21) );
endmodule

