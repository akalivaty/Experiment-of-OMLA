//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 0 0 1 0 1 0 0 0 1 1 0 1 1 1 0 1 0 0 1 0 1 1 0 1 0 1 1 0 1 0 1 1 1 1 0 1 0 1 0 1 1 0 1 0 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:15:14 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n684, new_n686,
    new_n687, new_n688, new_n690, new_n691, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n710,
    new_n711, new_n712, new_n713, new_n714, new_n715, new_n716, new_n717,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n729, new_n730, new_n731, new_n732, new_n734,
    new_n735, new_n736, new_n737, new_n739, new_n740, new_n741, new_n743,
    new_n744, new_n745, new_n746, new_n748, new_n750, new_n751, new_n752,
    new_n753, new_n754, new_n755, new_n756, new_n757, new_n758, new_n759,
    new_n760, new_n761, new_n762, new_n763, new_n764, new_n765, new_n766,
    new_n767, new_n768, new_n769, new_n770, new_n771, new_n772, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n816, new_n817,
    new_n818, new_n819, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n860, new_n862, new_n864,
    new_n865, new_n866, new_n867, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n921, new_n922, new_n923,
    new_n925, new_n926, new_n927, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n936, new_n937, new_n939, new_n940, new_n941,
    new_n943, new_n944, new_n945, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n952, new_n953, new_n954, new_n955, new_n956, new_n957,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n972, new_n973,
    new_n974, new_n975, new_n976, new_n977, new_n978, new_n979, new_n981,
    new_n982, new_n983, new_n984, new_n985;
  INV_X1    g000(.A(G148gat), .ZN(new_n202));
  NAND2_X1  g001(.A1(new_n202), .A2(KEYINPUT72), .ZN(new_n203));
  INV_X1    g002(.A(KEYINPUT72), .ZN(new_n204));
  NAND2_X1  g003(.A1(new_n204), .A2(G148gat), .ZN(new_n205));
  NAND3_X1  g004(.A1(new_n203), .A2(new_n205), .A3(G141gat), .ZN(new_n206));
  INV_X1    g005(.A(G141gat), .ZN(new_n207));
  NAND2_X1  g006(.A1(new_n207), .A2(G148gat), .ZN(new_n208));
  AND2_X1   g007(.A1(G155gat), .A2(G162gat), .ZN(new_n209));
  INV_X1    g008(.A(new_n209), .ZN(new_n210));
  NOR2_X1   g009(.A1(G155gat), .A2(G162gat), .ZN(new_n211));
  INV_X1    g010(.A(KEYINPUT2), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  AOI22_X1  g012(.A1(new_n206), .A2(new_n208), .B1(new_n210), .B2(new_n213), .ZN(new_n214));
  XNOR2_X1  g013(.A(G155gat), .B(G162gat), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n202), .A2(G141gat), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n208), .A2(new_n216), .ZN(new_n217));
  AOI21_X1  g016(.A(new_n215), .B1(new_n212), .B2(new_n217), .ZN(new_n218));
  OAI21_X1  g017(.A(KEYINPUT3), .B1(new_n214), .B2(new_n218), .ZN(new_n219));
  AND2_X1   g018(.A1(G228gat), .A2(G233gat), .ZN(new_n220));
  AND2_X1   g019(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n206), .A2(new_n208), .ZN(new_n222));
  AOI21_X1  g021(.A(new_n209), .B1(new_n212), .B2(new_n211), .ZN(new_n223));
  INV_X1    g022(.A(new_n223), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n217), .A2(new_n212), .ZN(new_n225));
  NOR2_X1   g024(.A1(new_n209), .A2(new_n211), .ZN(new_n226));
  AOI22_X1  g025(.A1(new_n222), .A2(new_n224), .B1(new_n225), .B2(new_n226), .ZN(new_n227));
  OR2_X1    g026(.A1(G197gat), .A2(G204gat), .ZN(new_n228));
  NAND2_X1  g027(.A1(G197gat), .A2(G204gat), .ZN(new_n229));
  INV_X1    g028(.A(KEYINPUT22), .ZN(new_n230));
  NAND2_X1  g029(.A1(G211gat), .A2(G218gat), .ZN(new_n231));
  AOI22_X1  g030(.A1(new_n228), .A2(new_n229), .B1(new_n230), .B2(new_n231), .ZN(new_n232));
  INV_X1    g031(.A(new_n232), .ZN(new_n233));
  OR2_X1    g032(.A1(G211gat), .A2(G218gat), .ZN(new_n234));
  INV_X1    g033(.A(KEYINPUT68), .ZN(new_n235));
  NAND3_X1  g034(.A1(new_n234), .A2(new_n235), .A3(new_n231), .ZN(new_n236));
  INV_X1    g035(.A(new_n236), .ZN(new_n237));
  AOI21_X1  g036(.A(new_n235), .B1(new_n234), .B2(new_n231), .ZN(new_n238));
  OAI21_X1  g037(.A(new_n233), .B1(new_n237), .B2(new_n238), .ZN(new_n239));
  INV_X1    g038(.A(new_n238), .ZN(new_n240));
  NAND3_X1  g039(.A1(new_n240), .A2(new_n232), .A3(new_n236), .ZN(new_n241));
  INV_X1    g040(.A(KEYINPUT29), .ZN(new_n242));
  NAND3_X1  g041(.A1(new_n239), .A2(new_n241), .A3(new_n242), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n239), .A2(new_n241), .ZN(new_n244));
  INV_X1    g043(.A(new_n244), .ZN(new_n245));
  INV_X1    g044(.A(KEYINPUT3), .ZN(new_n246));
  AOI21_X1  g045(.A(KEYINPUT29), .B1(new_n227), .B2(new_n246), .ZN(new_n247));
  OAI221_X1 g046(.A(new_n221), .B1(new_n227), .B2(new_n243), .C1(new_n245), .C2(new_n247), .ZN(new_n248));
  NOR2_X1   g047(.A1(new_n247), .A2(new_n245), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n243), .A2(KEYINPUT76), .ZN(new_n250));
  INV_X1    g049(.A(KEYINPUT76), .ZN(new_n251));
  NAND4_X1  g050(.A1(new_n239), .A2(new_n241), .A3(new_n251), .A4(new_n242), .ZN(new_n252));
  NAND3_X1  g051(.A1(new_n250), .A2(new_n246), .A3(new_n252), .ZN(new_n253));
  XNOR2_X1  g052(.A(G141gat), .B(G148gat), .ZN(new_n254));
  OAI21_X1  g053(.A(new_n226), .B1(new_n254), .B2(KEYINPUT2), .ZN(new_n255));
  INV_X1    g054(.A(new_n208), .ZN(new_n256));
  XNOR2_X1  g055(.A(KEYINPUT72), .B(G148gat), .ZN(new_n257));
  AOI21_X1  g056(.A(new_n256), .B1(new_n257), .B2(G141gat), .ZN(new_n258));
  OAI21_X1  g057(.A(new_n255), .B1(new_n258), .B2(new_n223), .ZN(new_n259));
  AOI21_X1  g058(.A(new_n249), .B1(new_n253), .B2(new_n259), .ZN(new_n260));
  OAI21_X1  g059(.A(new_n248), .B1(new_n260), .B2(new_n220), .ZN(new_n261));
  XOR2_X1   g060(.A(KEYINPUT77), .B(G22gat), .Z(new_n262));
  INV_X1    g061(.A(new_n262), .ZN(new_n263));
  NAND2_X1  g062(.A1(new_n261), .A2(new_n263), .ZN(new_n264));
  OAI211_X1 g063(.A(new_n262), .B(new_n248), .C1(new_n260), .C2(new_n220), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  XNOR2_X1  g065(.A(G78gat), .B(G106gat), .ZN(new_n267));
  XNOR2_X1  g066(.A(KEYINPUT31), .B(G50gat), .ZN(new_n268));
  XNOR2_X1  g067(.A(new_n267), .B(new_n268), .ZN(new_n269));
  XOR2_X1   g068(.A(new_n269), .B(KEYINPUT75), .Z(new_n270));
  AND2_X1   g069(.A1(new_n265), .A2(new_n269), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n261), .A2(G22gat), .ZN(new_n272));
  AOI22_X1  g071(.A1(new_n266), .A2(new_n270), .B1(new_n271), .B2(new_n272), .ZN(new_n273));
  INV_X1    g072(.A(KEYINPUT66), .ZN(new_n274));
  INV_X1    g073(.A(KEYINPUT25), .ZN(new_n275));
  AND2_X1   g074(.A1(G169gat), .A2(G176gat), .ZN(new_n276));
  INV_X1    g075(.A(G169gat), .ZN(new_n277));
  INV_X1    g076(.A(G176gat), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  INV_X1    g078(.A(KEYINPUT23), .ZN(new_n280));
  AOI21_X1  g079(.A(new_n276), .B1(new_n279), .B2(new_n280), .ZN(new_n281));
  NAND2_X1  g080(.A1(G183gat), .A2(G190gat), .ZN(new_n282));
  INV_X1    g081(.A(KEYINPUT24), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  INV_X1    g083(.A(G183gat), .ZN(new_n285));
  INV_X1    g084(.A(G190gat), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  NAND3_X1  g086(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n288));
  NAND3_X1  g087(.A1(new_n284), .A2(new_n287), .A3(new_n288), .ZN(new_n289));
  NAND3_X1  g088(.A1(new_n277), .A2(new_n278), .A3(KEYINPUT23), .ZN(new_n290));
  NAND3_X1  g089(.A1(new_n281), .A2(new_n289), .A3(new_n290), .ZN(new_n291));
  AND3_X1   g090(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n292));
  NOR2_X1   g091(.A1(G183gat), .A2(G190gat), .ZN(new_n293));
  NOR2_X1   g092(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  NAND2_X1  g093(.A1(new_n284), .A2(KEYINPUT64), .ZN(new_n295));
  AOI21_X1  g094(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n296));
  INV_X1    g095(.A(KEYINPUT64), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n296), .A2(new_n297), .ZN(new_n298));
  NAND3_X1  g097(.A1(new_n294), .A2(new_n295), .A3(new_n298), .ZN(new_n299));
  OAI21_X1  g098(.A(new_n280), .B1(G169gat), .B2(G176gat), .ZN(new_n300));
  NAND2_X1  g099(.A1(G169gat), .A2(G176gat), .ZN(new_n301));
  AND4_X1   g100(.A1(KEYINPUT25), .A2(new_n290), .A3(new_n300), .A4(new_n301), .ZN(new_n302));
  AOI22_X1  g101(.A1(new_n275), .A2(new_n291), .B1(new_n299), .B2(new_n302), .ZN(new_n303));
  NAND3_X1  g102(.A1(new_n277), .A2(new_n278), .A3(KEYINPUT26), .ZN(new_n304));
  INV_X1    g103(.A(KEYINPUT26), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n301), .A2(new_n305), .ZN(new_n306));
  NOR2_X1   g105(.A1(G169gat), .A2(G176gat), .ZN(new_n307));
  OAI211_X1 g106(.A(new_n282), .B(new_n304), .C1(new_n306), .C2(new_n307), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n285), .A2(KEYINPUT27), .ZN(new_n309));
  INV_X1    g108(.A(KEYINPUT27), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n310), .A2(G183gat), .ZN(new_n311));
  NAND3_X1  g110(.A1(new_n309), .A2(new_n311), .A3(new_n286), .ZN(new_n312));
  INV_X1    g111(.A(KEYINPUT28), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  XNOR2_X1  g113(.A(KEYINPUT27), .B(G183gat), .ZN(new_n315));
  NAND3_X1  g114(.A1(new_n315), .A2(KEYINPUT28), .A3(new_n286), .ZN(new_n316));
  AOI21_X1  g115(.A(new_n308), .B1(new_n314), .B2(new_n316), .ZN(new_n317));
  OAI21_X1  g116(.A(new_n274), .B1(new_n303), .B2(new_n317), .ZN(new_n318));
  INV_X1    g117(.A(G120gat), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n319), .A2(G113gat), .ZN(new_n320));
  INV_X1    g119(.A(G113gat), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n321), .A2(G120gat), .ZN(new_n322));
  AOI21_X1  g121(.A(KEYINPUT1), .B1(new_n320), .B2(new_n322), .ZN(new_n323));
  XNOR2_X1  g122(.A(G127gat), .B(G134gat), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n323), .A2(new_n324), .ZN(new_n325));
  XNOR2_X1  g124(.A(G113gat), .B(G120gat), .ZN(new_n326));
  OAI22_X1  g125(.A1(new_n326), .A2(KEYINPUT1), .B1(G127gat), .B2(G134gat), .ZN(new_n327));
  XNOR2_X1  g126(.A(KEYINPUT65), .B(G134gat), .ZN(new_n328));
  INV_X1    g127(.A(G127gat), .ZN(new_n329));
  NOR2_X1   g128(.A1(new_n328), .A2(new_n329), .ZN(new_n330));
  OAI21_X1  g129(.A(new_n325), .B1(new_n327), .B2(new_n330), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n299), .A2(new_n302), .ZN(new_n332));
  NOR3_X1   g131(.A1(new_n292), .A2(new_n296), .A3(new_n293), .ZN(new_n333));
  NAND3_X1  g132(.A1(new_n290), .A2(new_n300), .A3(new_n301), .ZN(new_n334));
  OAI21_X1  g133(.A(new_n275), .B1(new_n333), .B2(new_n334), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n332), .A2(new_n335), .ZN(new_n336));
  INV_X1    g135(.A(new_n308), .ZN(new_n337));
  AOI21_X1  g136(.A(KEYINPUT28), .B1(new_n315), .B2(new_n286), .ZN(new_n338));
  AND4_X1   g137(.A1(KEYINPUT28), .A2(new_n309), .A3(new_n311), .A4(new_n286), .ZN(new_n339));
  OAI21_X1  g138(.A(new_n337), .B1(new_n338), .B2(new_n339), .ZN(new_n340));
  NAND3_X1  g139(.A1(new_n336), .A2(KEYINPUT66), .A3(new_n340), .ZN(new_n341));
  NAND3_X1  g140(.A1(new_n318), .A2(new_n331), .A3(new_n341), .ZN(new_n342));
  INV_X1    g141(.A(G227gat), .ZN(new_n343));
  INV_X1    g142(.A(G233gat), .ZN(new_n344));
  NOR2_X1   g143(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  NAND4_X1  g144(.A1(new_n290), .A2(new_n300), .A3(KEYINPUT25), .A4(new_n301), .ZN(new_n346));
  AOI21_X1  g145(.A(new_n297), .B1(new_n282), .B2(new_n283), .ZN(new_n347));
  NOR3_X1   g146(.A1(new_n347), .A2(new_n293), .A3(new_n292), .ZN(new_n348));
  AOI21_X1  g147(.A(new_n346), .B1(new_n348), .B2(new_n298), .ZN(new_n349));
  AND3_X1   g148(.A1(new_n290), .A2(new_n300), .A3(new_n301), .ZN(new_n350));
  AOI21_X1  g149(.A(KEYINPUT25), .B1(new_n350), .B2(new_n289), .ZN(new_n351));
  OAI21_X1  g150(.A(new_n340), .B1(new_n349), .B2(new_n351), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n320), .A2(new_n322), .ZN(new_n353));
  INV_X1    g152(.A(KEYINPUT1), .ZN(new_n354));
  INV_X1    g153(.A(G134gat), .ZN(new_n355));
  AOI22_X1  g154(.A1(new_n353), .A2(new_n354), .B1(new_n329), .B2(new_n355), .ZN(new_n356));
  AND2_X1   g155(.A1(new_n355), .A2(KEYINPUT65), .ZN(new_n357));
  NOR2_X1   g156(.A1(new_n355), .A2(KEYINPUT65), .ZN(new_n358));
  OAI21_X1  g157(.A(G127gat), .B1(new_n357), .B2(new_n358), .ZN(new_n359));
  AOI22_X1  g158(.A1(new_n356), .A2(new_n359), .B1(new_n324), .B2(new_n323), .ZN(new_n360));
  NAND3_X1  g159(.A1(new_n352), .A2(new_n274), .A3(new_n360), .ZN(new_n361));
  NAND3_X1  g160(.A1(new_n342), .A2(new_n345), .A3(new_n361), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n362), .A2(KEYINPUT32), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n363), .A2(KEYINPUT67), .ZN(new_n364));
  INV_X1    g163(.A(KEYINPUT67), .ZN(new_n365));
  NAND3_X1  g164(.A1(new_n362), .A2(new_n365), .A3(KEYINPUT32), .ZN(new_n366));
  XNOR2_X1  g165(.A(G15gat), .B(G43gat), .ZN(new_n367));
  XNOR2_X1  g166(.A(G71gat), .B(G99gat), .ZN(new_n368));
  XNOR2_X1  g167(.A(new_n367), .B(new_n368), .ZN(new_n369));
  INV_X1    g168(.A(KEYINPUT33), .ZN(new_n370));
  AOI21_X1  g169(.A(new_n369), .B1(new_n362), .B2(new_n370), .ZN(new_n371));
  NAND3_X1  g170(.A1(new_n364), .A2(new_n366), .A3(new_n371), .ZN(new_n372));
  AOI21_X1  g171(.A(new_n345), .B1(new_n342), .B2(new_n361), .ZN(new_n373));
  INV_X1    g172(.A(KEYINPUT34), .ZN(new_n374));
  NOR2_X1   g173(.A1(new_n373), .A2(new_n374), .ZN(new_n375));
  AOI211_X1 g174(.A(KEYINPUT34), .B(new_n345), .C1(new_n342), .C2(new_n361), .ZN(new_n376));
  NOR2_X1   g175(.A1(new_n375), .A2(new_n376), .ZN(new_n377));
  OAI211_X1 g176(.A(new_n362), .B(KEYINPUT32), .C1(new_n370), .C2(new_n369), .ZN(new_n378));
  AND3_X1   g177(.A1(new_n372), .A2(new_n377), .A3(new_n378), .ZN(new_n379));
  AOI21_X1  g178(.A(new_n377), .B1(new_n372), .B2(new_n378), .ZN(new_n380));
  NOR3_X1   g179(.A1(new_n273), .A2(new_n379), .A3(new_n380), .ZN(new_n381));
  NAND2_X1  g180(.A1(G226gat), .A2(G233gat), .ZN(new_n382));
  INV_X1    g181(.A(new_n382), .ZN(new_n383));
  AOI21_X1  g182(.A(new_n383), .B1(new_n352), .B2(new_n242), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n314), .A2(new_n316), .ZN(new_n385));
  AOI22_X1  g184(.A1(new_n332), .A2(new_n335), .B1(new_n385), .B2(new_n337), .ZN(new_n386));
  NOR2_X1   g185(.A1(new_n386), .A2(new_n382), .ZN(new_n387));
  NOR3_X1   g186(.A1(new_n384), .A2(new_n387), .A3(new_n244), .ZN(new_n388));
  INV_X1    g187(.A(new_n388), .ZN(new_n389));
  XNOR2_X1  g188(.A(G8gat), .B(G36gat), .ZN(new_n390));
  XNOR2_X1  g189(.A(G64gat), .B(G92gat), .ZN(new_n391));
  XOR2_X1   g190(.A(new_n390), .B(new_n391), .Z(new_n392));
  INV_X1    g191(.A(KEYINPUT70), .ZN(new_n393));
  OAI21_X1  g192(.A(new_n393), .B1(new_n386), .B2(new_n382), .ZN(new_n394));
  NAND3_X1  g193(.A1(new_n352), .A2(KEYINPUT70), .A3(new_n383), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n394), .A2(new_n395), .ZN(new_n396));
  INV_X1    g195(.A(KEYINPUT69), .ZN(new_n397));
  AOI21_X1  g196(.A(KEYINPUT29), .B1(new_n336), .B2(new_n340), .ZN(new_n398));
  OAI21_X1  g197(.A(new_n397), .B1(new_n398), .B2(new_n383), .ZN(new_n399));
  OAI211_X1 g198(.A(KEYINPUT69), .B(new_n382), .C1(new_n386), .C2(KEYINPUT29), .ZN(new_n400));
  AOI21_X1  g199(.A(new_n396), .B1(new_n399), .B2(new_n400), .ZN(new_n401));
  OAI211_X1 g200(.A(new_n389), .B(new_n392), .C1(new_n401), .C2(new_n245), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n402), .A2(KEYINPUT30), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n399), .A2(new_n400), .ZN(new_n404));
  AND2_X1   g203(.A1(new_n394), .A2(new_n395), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n404), .A2(new_n405), .ZN(new_n406));
  NAND2_X1  g205(.A1(new_n406), .A2(new_n244), .ZN(new_n407));
  INV_X1    g206(.A(KEYINPUT30), .ZN(new_n408));
  NAND4_X1  g207(.A1(new_n407), .A2(new_n408), .A3(new_n389), .A4(new_n392), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n403), .A2(new_n409), .ZN(new_n410));
  XOR2_X1   g209(.A(G1gat), .B(G29gat), .Z(new_n411));
  XNOR2_X1  g210(.A(new_n411), .B(KEYINPUT0), .ZN(new_n412));
  XNOR2_X1  g211(.A(G57gat), .B(G85gat), .ZN(new_n413));
  XNOR2_X1  g212(.A(new_n412), .B(new_n413), .ZN(new_n414));
  NAND2_X1  g213(.A1(G225gat), .A2(G233gat), .ZN(new_n415));
  OAI211_X1 g214(.A(new_n246), .B(new_n255), .C1(new_n258), .C2(new_n223), .ZN(new_n416));
  NAND3_X1  g215(.A1(new_n219), .A2(new_n416), .A3(new_n331), .ZN(new_n417));
  INV_X1    g216(.A(KEYINPUT4), .ZN(new_n418));
  OAI21_X1  g217(.A(new_n418), .B1(new_n331), .B2(new_n259), .ZN(new_n419));
  NAND3_X1  g218(.A1(new_n360), .A2(new_n227), .A3(KEYINPUT4), .ZN(new_n420));
  AND4_X1   g219(.A1(new_n415), .A2(new_n417), .A3(new_n419), .A4(new_n420), .ZN(new_n421));
  INV_X1    g220(.A(KEYINPUT5), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n360), .A2(new_n227), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n331), .A2(new_n259), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n423), .A2(new_n424), .ZN(new_n425));
  INV_X1    g224(.A(new_n415), .ZN(new_n426));
  AOI21_X1  g225(.A(new_n422), .B1(new_n425), .B2(new_n426), .ZN(new_n427));
  NOR2_X1   g226(.A1(new_n421), .A2(new_n427), .ZN(new_n428));
  NAND4_X1  g227(.A1(new_n417), .A2(new_n419), .A3(new_n420), .A4(new_n415), .ZN(new_n429));
  NOR2_X1   g228(.A1(new_n429), .A2(new_n422), .ZN(new_n430));
  OAI21_X1  g229(.A(new_n414), .B1(new_n428), .B2(new_n430), .ZN(new_n431));
  INV_X1    g230(.A(KEYINPUT6), .ZN(new_n432));
  AND2_X1   g231(.A1(new_n419), .A2(new_n420), .ZN(new_n433));
  NAND4_X1  g232(.A1(new_n433), .A2(KEYINPUT5), .A3(new_n415), .A4(new_n417), .ZN(new_n434));
  AOI21_X1  g233(.A(new_n415), .B1(new_n423), .B2(new_n424), .ZN(new_n435));
  OAI21_X1  g234(.A(new_n429), .B1(new_n422), .B2(new_n435), .ZN(new_n436));
  INV_X1    g235(.A(new_n414), .ZN(new_n437));
  NAND3_X1  g236(.A1(new_n434), .A2(new_n436), .A3(new_n437), .ZN(new_n438));
  NAND3_X1  g237(.A1(new_n431), .A2(new_n432), .A3(new_n438), .ZN(new_n439));
  AND2_X1   g238(.A1(new_n434), .A2(new_n436), .ZN(new_n440));
  INV_X1    g239(.A(KEYINPUT73), .ZN(new_n441));
  NAND4_X1  g240(.A1(new_n440), .A2(new_n441), .A3(KEYINPUT6), .A4(new_n437), .ZN(new_n442));
  NAND4_X1  g241(.A1(new_n434), .A2(new_n436), .A3(KEYINPUT6), .A4(new_n437), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n443), .A2(KEYINPUT73), .ZN(new_n444));
  NAND3_X1  g243(.A1(new_n439), .A2(new_n442), .A3(new_n444), .ZN(new_n445));
  AOI21_X1  g244(.A(new_n245), .B1(new_n404), .B2(new_n405), .ZN(new_n446));
  OAI21_X1  g245(.A(KEYINPUT71), .B1(new_n446), .B2(new_n388), .ZN(new_n447));
  INV_X1    g246(.A(KEYINPUT71), .ZN(new_n448));
  OAI211_X1 g247(.A(new_n448), .B(new_n389), .C1(new_n401), .C2(new_n245), .ZN(new_n449));
  INV_X1    g248(.A(new_n392), .ZN(new_n450));
  NAND3_X1  g249(.A1(new_n447), .A2(new_n449), .A3(new_n450), .ZN(new_n451));
  NAND3_X1  g250(.A1(new_n410), .A2(new_n445), .A3(new_n451), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n452), .A2(KEYINPUT74), .ZN(new_n453));
  INV_X1    g252(.A(KEYINPUT74), .ZN(new_n454));
  NAND4_X1  g253(.A1(new_n410), .A2(new_n445), .A3(new_n454), .A4(new_n451), .ZN(new_n455));
  NAND3_X1  g254(.A1(new_n381), .A2(new_n453), .A3(new_n455), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n456), .A2(KEYINPUT35), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n372), .A2(new_n378), .ZN(new_n458));
  INV_X1    g257(.A(new_n377), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  NAND3_X1  g259(.A1(new_n372), .A2(new_n377), .A3(new_n378), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  XNOR2_X1  g261(.A(KEYINPUT81), .B(KEYINPUT35), .ZN(new_n463));
  NOR3_X1   g262(.A1(new_n462), .A2(new_n273), .A3(new_n463), .ZN(new_n464));
  INV_X1    g263(.A(KEYINPUT80), .ZN(new_n465));
  AOI21_X1  g264(.A(new_n388), .B1(new_n406), .B2(new_n244), .ZN(new_n466));
  AOI21_X1  g265(.A(new_n408), .B1(new_n466), .B2(new_n392), .ZN(new_n467));
  NOR4_X1   g266(.A1(new_n446), .A2(KEYINPUT30), .A3(new_n388), .A4(new_n450), .ZN(new_n468));
  OAI21_X1  g267(.A(new_n451), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  INV_X1    g268(.A(new_n469), .ZN(new_n470));
  OAI21_X1  g269(.A(KEYINPUT79), .B1(new_n428), .B2(new_n430), .ZN(new_n471));
  INV_X1    g270(.A(KEYINPUT79), .ZN(new_n472));
  NAND3_X1  g271(.A1(new_n434), .A2(new_n436), .A3(new_n472), .ZN(new_n473));
  NAND3_X1  g272(.A1(new_n471), .A2(new_n437), .A3(new_n473), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n434), .A2(new_n436), .ZN(new_n475));
  AOI21_X1  g274(.A(KEYINPUT6), .B1(new_n475), .B2(new_n414), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n474), .A2(new_n476), .ZN(new_n477));
  XNOR2_X1  g276(.A(new_n443), .B(new_n441), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  AOI21_X1  g278(.A(new_n465), .B1(new_n470), .B2(new_n479), .ZN(new_n480));
  NAND4_X1  g279(.A1(new_n479), .A2(new_n465), .A3(new_n451), .A4(new_n410), .ZN(new_n481));
  INV_X1    g280(.A(new_n481), .ZN(new_n482));
  OAI21_X1  g281(.A(new_n464), .B1(new_n480), .B2(new_n482), .ZN(new_n483));
  INV_X1    g282(.A(KEYINPUT37), .ZN(new_n484));
  OAI211_X1 g283(.A(new_n484), .B(new_n389), .C1(new_n401), .C2(new_n245), .ZN(new_n485));
  NOR2_X1   g284(.A1(new_n384), .A2(new_n387), .ZN(new_n486));
  AOI21_X1  g285(.A(new_n484), .B1(new_n486), .B2(new_n244), .ZN(new_n487));
  OAI21_X1  g286(.A(new_n487), .B1(new_n401), .B2(new_n244), .ZN(new_n488));
  INV_X1    g287(.A(KEYINPUT38), .ZN(new_n489));
  NAND4_X1  g288(.A1(new_n485), .A2(new_n488), .A3(new_n489), .A4(new_n450), .ZN(new_n490));
  AND4_X1   g289(.A1(new_n478), .A2(new_n477), .A3(new_n490), .A4(new_n402), .ZN(new_n491));
  NAND3_X1  g290(.A1(new_n447), .A2(KEYINPUT37), .A3(new_n449), .ZN(new_n492));
  AOI21_X1  g291(.A(new_n392), .B1(new_n466), .B2(new_n484), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n494), .A2(KEYINPUT38), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n491), .A2(new_n495), .ZN(new_n496));
  OAI21_X1  g295(.A(KEYINPUT78), .B1(new_n425), .B2(new_n426), .ZN(new_n497));
  INV_X1    g296(.A(KEYINPUT78), .ZN(new_n498));
  NAND4_X1  g297(.A1(new_n423), .A2(new_n424), .A3(new_n498), .A4(new_n415), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n497), .A2(new_n499), .ZN(new_n500));
  NAND3_X1  g299(.A1(new_n417), .A2(new_n419), .A3(new_n420), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n501), .A2(new_n426), .ZN(new_n502));
  NAND3_X1  g301(.A1(new_n500), .A2(KEYINPUT39), .A3(new_n502), .ZN(new_n503));
  OR2_X1    g302(.A1(new_n502), .A2(KEYINPUT39), .ZN(new_n504));
  NAND3_X1  g303(.A1(new_n503), .A2(new_n504), .A3(new_n414), .ZN(new_n505));
  INV_X1    g304(.A(KEYINPUT40), .ZN(new_n506));
  NAND2_X1  g305(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  NAND4_X1  g306(.A1(new_n503), .A2(new_n504), .A3(KEYINPUT40), .A4(new_n414), .ZN(new_n508));
  AND3_X1   g307(.A1(new_n507), .A2(new_n474), .A3(new_n508), .ZN(new_n509));
  AOI21_X1  g308(.A(new_n273), .B1(new_n469), .B2(new_n509), .ZN(new_n510));
  NAND3_X1  g309(.A1(new_n460), .A2(KEYINPUT36), .A3(new_n461), .ZN(new_n511));
  INV_X1    g310(.A(KEYINPUT36), .ZN(new_n512));
  OAI21_X1  g311(.A(new_n512), .B1(new_n379), .B2(new_n380), .ZN(new_n513));
  AOI22_X1  g312(.A1(new_n496), .A2(new_n510), .B1(new_n511), .B2(new_n513), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n453), .A2(new_n455), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n515), .A2(new_n273), .ZN(new_n516));
  AOI22_X1  g315(.A1(new_n457), .A2(new_n483), .B1(new_n514), .B2(new_n516), .ZN(new_n517));
  XNOR2_X1  g316(.A(G15gat), .B(G22gat), .ZN(new_n518));
  OR2_X1    g317(.A1(new_n518), .A2(G1gat), .ZN(new_n519));
  INV_X1    g318(.A(G8gat), .ZN(new_n520));
  INV_X1    g319(.A(KEYINPUT16), .ZN(new_n521));
  OAI21_X1  g320(.A(new_n518), .B1(new_n521), .B2(G1gat), .ZN(new_n522));
  NAND3_X1  g321(.A1(new_n519), .A2(new_n520), .A3(new_n522), .ZN(new_n523));
  INV_X1    g322(.A(new_n523), .ZN(new_n524));
  INV_X1    g323(.A(KEYINPUT84), .ZN(new_n525));
  AOI21_X1  g324(.A(new_n520), .B1(new_n519), .B2(new_n522), .ZN(new_n526));
  NOR3_X1   g325(.A1(new_n524), .A2(new_n525), .A3(new_n526), .ZN(new_n527));
  INV_X1    g326(.A(new_n527), .ZN(new_n528));
  INV_X1    g327(.A(G36gat), .ZN(new_n529));
  AND2_X1   g328(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n530));
  NOR2_X1   g329(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n531));
  OAI21_X1  g330(.A(new_n529), .B1(new_n530), .B2(new_n531), .ZN(new_n532));
  INV_X1    g331(.A(G29gat), .ZN(new_n533));
  NAND3_X1  g332(.A1(new_n533), .A2(KEYINPUT14), .A3(G36gat), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n532), .A2(new_n534), .ZN(new_n535));
  OR2_X1    g334(.A1(new_n535), .A2(KEYINPUT15), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n535), .A2(KEYINPUT15), .ZN(new_n537));
  XNOR2_X1  g336(.A(G43gat), .B(G50gat), .ZN(new_n538));
  NAND3_X1  g337(.A1(new_n536), .A2(new_n537), .A3(new_n538), .ZN(new_n539));
  OR2_X1    g338(.A1(new_n537), .A2(new_n538), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  OAI21_X1  g340(.A(new_n525), .B1(new_n524), .B2(new_n526), .ZN(new_n542));
  NAND3_X1  g341(.A1(new_n528), .A2(new_n541), .A3(new_n542), .ZN(new_n543));
  AND2_X1   g342(.A1(new_n539), .A2(new_n540), .ZN(new_n544));
  INV_X1    g343(.A(new_n526), .ZN(new_n545));
  AOI21_X1  g344(.A(KEYINPUT84), .B1(new_n545), .B2(new_n523), .ZN(new_n546));
  OAI21_X1  g345(.A(new_n544), .B1(new_n527), .B2(new_n546), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n543), .A2(new_n547), .ZN(new_n548));
  NAND2_X1  g347(.A1(G229gat), .A2(G233gat), .ZN(new_n549));
  XOR2_X1   g348(.A(new_n549), .B(KEYINPUT13), .Z(new_n550));
  NAND2_X1  g349(.A1(new_n548), .A2(new_n550), .ZN(new_n551));
  INV_X1    g350(.A(KEYINPUT86), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  XNOR2_X1  g352(.A(KEYINPUT82), .B(KEYINPUT17), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n541), .A2(new_n554), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n555), .A2(KEYINPUT83), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n544), .A2(KEYINPUT17), .ZN(new_n557));
  NOR2_X1   g356(.A1(new_n524), .A2(new_n526), .ZN(new_n558));
  INV_X1    g357(.A(KEYINPUT83), .ZN(new_n559));
  NAND3_X1  g358(.A1(new_n541), .A2(new_n559), .A3(new_n554), .ZN(new_n560));
  NAND4_X1  g359(.A1(new_n556), .A2(new_n557), .A3(new_n558), .A4(new_n560), .ZN(new_n561));
  NAND4_X1  g360(.A1(new_n561), .A2(KEYINPUT18), .A3(new_n549), .A4(new_n543), .ZN(new_n562));
  NAND3_X1  g361(.A1(new_n548), .A2(KEYINPUT86), .A3(new_n550), .ZN(new_n563));
  AND3_X1   g362(.A1(new_n553), .A2(new_n562), .A3(new_n563), .ZN(new_n564));
  NAND3_X1  g363(.A1(new_n561), .A2(new_n549), .A3(new_n543), .ZN(new_n565));
  INV_X1    g364(.A(KEYINPUT18), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  XNOR2_X1  g366(.A(G113gat), .B(G141gat), .ZN(new_n568));
  XNOR2_X1  g367(.A(new_n568), .B(G197gat), .ZN(new_n569));
  XOR2_X1   g368(.A(KEYINPUT11), .B(G169gat), .Z(new_n570));
  XNOR2_X1  g369(.A(new_n569), .B(new_n570), .ZN(new_n571));
  XOR2_X1   g370(.A(new_n571), .B(KEYINPUT12), .Z(new_n572));
  INV_X1    g371(.A(new_n572), .ZN(new_n573));
  OAI211_X1 g372(.A(new_n564), .B(new_n567), .C1(KEYINPUT85), .C2(new_n573), .ZN(new_n574));
  NAND4_X1  g373(.A1(new_n553), .A2(new_n562), .A3(KEYINPUT85), .A4(new_n563), .ZN(new_n575));
  INV_X1    g374(.A(new_n567), .ZN(new_n576));
  NAND3_X1  g375(.A1(new_n553), .A2(new_n562), .A3(new_n563), .ZN(new_n577));
  OAI211_X1 g376(.A(new_n575), .B(new_n572), .C1(new_n576), .C2(new_n577), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n574), .A2(new_n578), .ZN(new_n579));
  INV_X1    g378(.A(KEYINPUT87), .ZN(new_n580));
  NAND2_X1  g379(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  NAND3_X1  g380(.A1(new_n574), .A2(new_n578), .A3(KEYINPUT87), .ZN(new_n582));
  NAND2_X1  g381(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  NOR2_X1   g382(.A1(new_n517), .A2(new_n583), .ZN(new_n584));
  INV_X1    g383(.A(KEYINPUT21), .ZN(new_n585));
  XNOR2_X1  g384(.A(G57gat), .B(G64gat), .ZN(new_n586));
  INV_X1    g385(.A(KEYINPUT9), .ZN(new_n587));
  NAND2_X1  g386(.A1(G71gat), .A2(G78gat), .ZN(new_n588));
  AOI21_X1  g387(.A(new_n586), .B1(new_n587), .B2(new_n588), .ZN(new_n589));
  XNOR2_X1  g388(.A(G71gat), .B(G78gat), .ZN(new_n590));
  OR2_X1    g389(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n589), .A2(new_n590), .ZN(new_n592));
  NAND2_X1  g391(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  OAI22_X1  g392(.A1(new_n546), .A2(new_n527), .B1(new_n585), .B2(new_n593), .ZN(new_n594));
  XOR2_X1   g393(.A(new_n594), .B(KEYINPUT90), .Z(new_n595));
  NAND2_X1  g394(.A1(G231gat), .A2(G233gat), .ZN(new_n596));
  XNOR2_X1  g395(.A(new_n596), .B(KEYINPUT89), .ZN(new_n597));
  XNOR2_X1  g396(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n598));
  XNOR2_X1  g397(.A(new_n597), .B(new_n598), .ZN(new_n599));
  INV_X1    g398(.A(new_n599), .ZN(new_n600));
  OR2_X1    g399(.A1(new_n595), .A2(new_n600), .ZN(new_n601));
  XNOR2_X1  g400(.A(KEYINPUT88), .B(KEYINPUT21), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n593), .A2(new_n602), .ZN(new_n603));
  XOR2_X1   g402(.A(G127gat), .B(G155gat), .Z(new_n604));
  XNOR2_X1  g403(.A(new_n603), .B(new_n604), .ZN(new_n605));
  XOR2_X1   g404(.A(G183gat), .B(G211gat), .Z(new_n606));
  XNOR2_X1  g405(.A(new_n605), .B(new_n606), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n595), .A2(new_n600), .ZN(new_n608));
  AND3_X1   g407(.A1(new_n601), .A2(new_n607), .A3(new_n608), .ZN(new_n609));
  AOI21_X1  g408(.A(new_n607), .B1(new_n601), .B2(new_n608), .ZN(new_n610));
  NOR2_X1   g409(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  AND2_X1   g410(.A1(G232gat), .A2(G233gat), .ZN(new_n612));
  NOR2_X1   g411(.A1(new_n612), .A2(KEYINPUT41), .ZN(new_n613));
  XNOR2_X1  g412(.A(G134gat), .B(G162gat), .ZN(new_n614));
  XNOR2_X1  g413(.A(new_n613), .B(new_n614), .ZN(new_n615));
  INV_X1    g414(.A(new_n615), .ZN(new_n616));
  NAND3_X1  g415(.A1(new_n556), .A2(new_n557), .A3(new_n560), .ZN(new_n617));
  INV_X1    g416(.A(G85gat), .ZN(new_n618));
  INV_X1    g417(.A(G92gat), .ZN(new_n619));
  INV_X1    g418(.A(KEYINPUT7), .ZN(new_n620));
  AOI211_X1 g419(.A(new_n618), .B(new_n619), .C1(KEYINPUT91), .C2(new_n620), .ZN(new_n621));
  OAI21_X1  g420(.A(new_n621), .B1(KEYINPUT91), .B2(new_n620), .ZN(new_n622));
  INV_X1    g421(.A(KEYINPUT8), .ZN(new_n623));
  NAND2_X1  g422(.A1(G99gat), .A2(G106gat), .ZN(new_n624));
  INV_X1    g423(.A(KEYINPUT92), .ZN(new_n625));
  AOI21_X1  g424(.A(new_n623), .B1(new_n624), .B2(new_n625), .ZN(new_n626));
  OAI21_X1  g425(.A(new_n626), .B1(new_n625), .B2(new_n624), .ZN(new_n627));
  INV_X1    g426(.A(KEYINPUT91), .ZN(new_n628));
  OAI22_X1  g427(.A1(new_n628), .A2(KEYINPUT7), .B1(G85gat), .B2(G92gat), .ZN(new_n629));
  OAI21_X1  g428(.A(new_n629), .B1(new_n618), .B2(new_n619), .ZN(new_n630));
  NAND3_X1  g429(.A1(new_n622), .A2(new_n627), .A3(new_n630), .ZN(new_n631));
  XNOR2_X1  g430(.A(G99gat), .B(G106gat), .ZN(new_n632));
  INV_X1    g431(.A(new_n632), .ZN(new_n633));
  NAND2_X1  g432(.A1(new_n631), .A2(new_n633), .ZN(new_n634));
  NAND4_X1  g433(.A1(new_n622), .A2(new_n632), .A3(new_n627), .A4(new_n630), .ZN(new_n635));
  AND3_X1   g434(.A1(new_n634), .A2(KEYINPUT93), .A3(new_n635), .ZN(new_n636));
  AOI21_X1  g435(.A(KEYINPUT93), .B1(new_n634), .B2(new_n635), .ZN(new_n637));
  NOR2_X1   g436(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  OR2_X1    g437(.A1(new_n617), .A2(new_n638), .ZN(new_n639));
  AOI22_X1  g438(.A1(new_n638), .A2(new_n541), .B1(KEYINPUT41), .B2(new_n612), .ZN(new_n640));
  XOR2_X1   g439(.A(G190gat), .B(G218gat), .Z(new_n641));
  INV_X1    g440(.A(new_n641), .ZN(new_n642));
  NAND3_X1  g441(.A1(new_n639), .A2(new_n640), .A3(new_n642), .ZN(new_n643));
  INV_X1    g442(.A(new_n643), .ZN(new_n644));
  AOI21_X1  g443(.A(new_n642), .B1(new_n639), .B2(new_n640), .ZN(new_n645));
  OAI21_X1  g444(.A(new_n616), .B1(new_n644), .B2(new_n645), .ZN(new_n646));
  INV_X1    g445(.A(new_n645), .ZN(new_n647));
  NAND3_X1  g446(.A1(new_n647), .A2(new_n615), .A3(new_n643), .ZN(new_n648));
  NAND2_X1  g447(.A1(new_n646), .A2(new_n648), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n611), .A2(new_n649), .ZN(new_n650));
  NAND2_X1  g449(.A1(G230gat), .A2(G233gat), .ZN(new_n651));
  XNOR2_X1  g450(.A(new_n651), .B(KEYINPUT95), .ZN(new_n652));
  INV_X1    g451(.A(new_n652), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n634), .A2(new_n635), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n654), .A2(KEYINPUT94), .ZN(new_n655));
  INV_X1    g454(.A(KEYINPUT94), .ZN(new_n656));
  NAND3_X1  g455(.A1(new_n634), .A2(new_n656), .A3(new_n635), .ZN(new_n657));
  NAND3_X1  g456(.A1(new_n655), .A2(new_n593), .A3(new_n657), .ZN(new_n658));
  NAND4_X1  g457(.A1(new_n654), .A2(KEYINPUT94), .A3(new_n591), .A4(new_n592), .ZN(new_n659));
  AOI21_X1  g458(.A(KEYINPUT10), .B1(new_n658), .B2(new_n659), .ZN(new_n660));
  INV_X1    g459(.A(KEYINPUT10), .ZN(new_n661));
  NOR4_X1   g460(.A1(new_n636), .A2(new_n637), .A3(new_n661), .A4(new_n593), .ZN(new_n662));
  OAI21_X1  g461(.A(new_n653), .B1(new_n660), .B2(new_n662), .ZN(new_n663));
  NAND3_X1  g462(.A1(new_n658), .A2(new_n652), .A3(new_n659), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  XNOR2_X1  g464(.A(G120gat), .B(G148gat), .ZN(new_n666));
  XNOR2_X1  g465(.A(G176gat), .B(G204gat), .ZN(new_n667));
  XOR2_X1   g466(.A(new_n666), .B(new_n667), .Z(new_n668));
  INV_X1    g467(.A(new_n668), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n665), .A2(new_n669), .ZN(new_n670));
  NAND3_X1  g469(.A1(new_n663), .A2(new_n664), .A3(new_n668), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  NOR2_X1   g471(.A1(new_n650), .A2(new_n672), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n584), .A2(new_n673), .ZN(new_n674));
  INV_X1    g473(.A(new_n674), .ZN(new_n675));
  INV_X1    g474(.A(new_n445), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  XNOR2_X1  g476(.A(new_n677), .B(G1gat), .ZN(G1324gat));
  INV_X1    g477(.A(KEYINPUT42), .ZN(new_n679));
  XOR2_X1   g478(.A(KEYINPUT16), .B(G8gat), .Z(new_n680));
  NAND3_X1  g479(.A1(new_n675), .A2(new_n469), .A3(new_n680), .ZN(new_n681));
  OAI21_X1  g480(.A(G8gat), .B1(new_n674), .B2(new_n470), .ZN(new_n682));
  AOI21_X1  g481(.A(new_n679), .B1(new_n681), .B2(new_n682), .ZN(new_n683));
  AOI21_X1  g482(.A(new_n683), .B1(new_n679), .B2(new_n681), .ZN(new_n684));
  XOR2_X1   g483(.A(new_n684), .B(KEYINPUT96), .Z(G1325gat));
  NAND2_X1  g484(.A1(new_n513), .A2(new_n511), .ZN(new_n686));
  OAI21_X1  g485(.A(G15gat), .B1(new_n674), .B2(new_n686), .ZN(new_n687));
  OR2_X1    g486(.A1(new_n462), .A2(G15gat), .ZN(new_n688));
  OAI21_X1  g487(.A(new_n687), .B1(new_n674), .B2(new_n688), .ZN(G1326gat));
  NAND3_X1  g488(.A1(new_n584), .A2(new_n273), .A3(new_n673), .ZN(new_n690));
  XNOR2_X1  g489(.A(KEYINPUT43), .B(G22gat), .ZN(new_n691));
  XNOR2_X1  g490(.A(new_n690), .B(new_n691), .ZN(G1327gat));
  INV_X1    g491(.A(new_n611), .ZN(new_n693));
  INV_X1    g492(.A(new_n672), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  NOR2_X1   g494(.A1(new_n695), .A2(new_n649), .ZN(new_n696));
  NAND2_X1  g495(.A1(new_n584), .A2(new_n696), .ZN(new_n697));
  NOR3_X1   g496(.A1(new_n697), .A2(G29gat), .A3(new_n445), .ZN(new_n698));
  XOR2_X1   g497(.A(new_n698), .B(KEYINPUT45), .Z(new_n699));
  NAND2_X1  g498(.A1(new_n457), .A2(new_n483), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n514), .A2(new_n516), .ZN(new_n701));
  AOI21_X1  g500(.A(new_n649), .B1(new_n700), .B2(new_n701), .ZN(new_n702));
  NAND2_X1  g501(.A1(new_n702), .A2(KEYINPUT97), .ZN(new_n703));
  XNOR2_X1  g502(.A(new_n703), .B(KEYINPUT44), .ZN(new_n704));
  AND2_X1   g503(.A1(new_n574), .A2(new_n578), .ZN(new_n705));
  NOR2_X1   g504(.A1(new_n695), .A2(new_n705), .ZN(new_n706));
  NAND2_X1  g505(.A1(new_n704), .A2(new_n706), .ZN(new_n707));
  OAI21_X1  g506(.A(G29gat), .B1(new_n707), .B2(new_n445), .ZN(new_n708));
  NAND2_X1  g507(.A1(new_n699), .A2(new_n708), .ZN(G1328gat));
  AND2_X1   g508(.A1(KEYINPUT98), .A2(KEYINPUT46), .ZN(new_n710));
  NOR2_X1   g509(.A1(KEYINPUT98), .A2(KEYINPUT46), .ZN(new_n711));
  NOR2_X1   g510(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  NOR3_X1   g511(.A1(new_n697), .A2(G36gat), .A3(new_n470), .ZN(new_n713));
  MUX2_X1   g512(.A(new_n712), .B(new_n710), .S(new_n713), .Z(new_n714));
  NOR2_X1   g513(.A1(new_n707), .A2(new_n470), .ZN(new_n715));
  AND2_X1   g514(.A1(new_n715), .A2(KEYINPUT99), .ZN(new_n716));
  OAI21_X1  g515(.A(G36gat), .B1(new_n715), .B2(KEYINPUT99), .ZN(new_n717));
  OAI21_X1  g516(.A(new_n714), .B1(new_n716), .B2(new_n717), .ZN(G1329gat));
  OR3_X1    g517(.A1(new_n697), .A2(G43gat), .A3(new_n462), .ZN(new_n719));
  AND2_X1   g518(.A1(new_n513), .A2(new_n511), .ZN(new_n720));
  NAND3_X1  g519(.A1(new_n704), .A2(new_n720), .A3(new_n706), .ZN(new_n721));
  NAND2_X1  g520(.A1(new_n721), .A2(KEYINPUT100), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n722), .A2(G43gat), .ZN(new_n723));
  NOR2_X1   g522(.A1(new_n721), .A2(KEYINPUT100), .ZN(new_n724));
  OAI211_X1 g523(.A(KEYINPUT47), .B(new_n719), .C1(new_n723), .C2(new_n724), .ZN(new_n725));
  NAND2_X1  g524(.A1(new_n721), .A2(G43gat), .ZN(new_n726));
  AND2_X1   g525(.A1(new_n726), .A2(new_n719), .ZN(new_n727));
  OAI21_X1  g526(.A(new_n725), .B1(KEYINPUT47), .B2(new_n727), .ZN(G1330gat));
  INV_X1    g527(.A(new_n273), .ZN(new_n729));
  OAI21_X1  g528(.A(G50gat), .B1(new_n707), .B2(new_n729), .ZN(new_n730));
  OR2_X1    g529(.A1(new_n729), .A2(G50gat), .ZN(new_n731));
  OAI21_X1  g530(.A(new_n730), .B1(new_n697), .B2(new_n731), .ZN(new_n732));
  XOR2_X1   g531(.A(new_n732), .B(KEYINPUT48), .Z(G1331gat));
  NOR4_X1   g532(.A1(new_n517), .A2(new_n579), .A3(new_n650), .A4(new_n694), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n734), .A2(new_n676), .ZN(new_n735));
  XNOR2_X1  g534(.A(new_n735), .B(KEYINPUT102), .ZN(new_n736));
  XOR2_X1   g535(.A(KEYINPUT101), .B(G57gat), .Z(new_n737));
  XNOR2_X1  g536(.A(new_n736), .B(new_n737), .ZN(G1332gat));
  AOI21_X1  g537(.A(new_n470), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n734), .A2(new_n739), .ZN(new_n740));
  NOR2_X1   g539(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n741));
  XOR2_X1   g540(.A(new_n740), .B(new_n741), .Z(G1333gat));
  NAND3_X1  g541(.A1(new_n734), .A2(G71gat), .A3(new_n720), .ZN(new_n743));
  XOR2_X1   g542(.A(new_n462), .B(KEYINPUT103), .Z(new_n744));
  AND2_X1   g543(.A1(new_n734), .A2(new_n744), .ZN(new_n745));
  OAI21_X1  g544(.A(new_n743), .B1(new_n745), .B2(G71gat), .ZN(new_n746));
  XNOR2_X1  g545(.A(new_n746), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g546(.A1(new_n734), .A2(new_n273), .ZN(new_n748));
  XNOR2_X1  g547(.A(new_n748), .B(G78gat), .ZN(G1335gat));
  INV_X1    g548(.A(KEYINPUT105), .ZN(new_n750));
  NOR2_X1   g549(.A1(new_n611), .A2(new_n579), .ZN(new_n751));
  INV_X1    g550(.A(new_n751), .ZN(new_n752));
  AOI21_X1  g551(.A(new_n752), .B1(new_n702), .B2(KEYINPUT104), .ZN(new_n753));
  INV_X1    g552(.A(KEYINPUT104), .ZN(new_n754));
  OAI21_X1  g553(.A(new_n754), .B1(new_n517), .B2(new_n649), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n753), .A2(new_n755), .ZN(new_n756));
  INV_X1    g555(.A(KEYINPUT51), .ZN(new_n757));
  OAI21_X1  g556(.A(new_n750), .B1(new_n756), .B2(new_n757), .ZN(new_n758));
  NAND4_X1  g557(.A1(new_n753), .A2(KEYINPUT105), .A3(KEYINPUT51), .A4(new_n755), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n756), .A2(new_n757), .ZN(new_n760));
  NAND3_X1  g559(.A1(new_n758), .A2(new_n759), .A3(new_n760), .ZN(new_n761));
  INV_X1    g560(.A(KEYINPUT106), .ZN(new_n762));
  AOI21_X1  g561(.A(new_n694), .B1(new_n761), .B2(new_n762), .ZN(new_n763));
  NAND4_X1  g562(.A1(new_n758), .A2(new_n759), .A3(KEYINPUT106), .A4(new_n760), .ZN(new_n764));
  NAND4_X1  g563(.A1(new_n763), .A2(new_n618), .A3(new_n676), .A4(new_n764), .ZN(new_n765));
  NOR2_X1   g564(.A1(new_n752), .A2(new_n694), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n704), .A2(new_n766), .ZN(new_n767));
  OAI21_X1  g566(.A(G85gat), .B1(new_n767), .B2(new_n445), .ZN(new_n768));
  NAND2_X1  g567(.A1(new_n765), .A2(new_n768), .ZN(new_n769));
  INV_X1    g568(.A(KEYINPUT107), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  NAND3_X1  g570(.A1(new_n765), .A2(KEYINPUT107), .A3(new_n768), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n771), .A2(new_n772), .ZN(G1336gat));
  OAI21_X1  g572(.A(G92gat), .B1(new_n767), .B2(new_n470), .ZN(new_n774));
  NOR3_X1   g573(.A1(new_n694), .A2(G92gat), .A3(new_n470), .ZN(new_n775));
  XOR2_X1   g574(.A(new_n775), .B(KEYINPUT108), .Z(new_n776));
  NOR2_X1   g575(.A1(new_n756), .A2(new_n757), .ZN(new_n777));
  XOR2_X1   g576(.A(KEYINPUT110), .B(KEYINPUT51), .Z(new_n778));
  INV_X1    g577(.A(new_n778), .ZN(new_n779));
  INV_X1    g578(.A(KEYINPUT109), .ZN(new_n780));
  INV_X1    g579(.A(new_n649), .ZN(new_n781));
  AND2_X1   g580(.A1(new_n477), .A2(new_n478), .ZN(new_n782));
  OAI21_X1  g581(.A(KEYINPUT80), .B1(new_n782), .B2(new_n469), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n783), .A2(new_n481), .ZN(new_n784));
  AOI22_X1  g583(.A1(KEYINPUT35), .A2(new_n456), .B1(new_n784), .B2(new_n464), .ZN(new_n785));
  NAND2_X1  g584(.A1(new_n469), .A2(new_n509), .ZN(new_n786));
  NAND2_X1  g585(.A1(new_n786), .A2(new_n729), .ZN(new_n787));
  NAND4_X1  g586(.A1(new_n477), .A2(new_n478), .A3(new_n490), .A4(new_n402), .ZN(new_n788));
  AOI21_X1  g587(.A(new_n489), .B1(new_n492), .B2(new_n493), .ZN(new_n789));
  NOR2_X1   g588(.A1(new_n788), .A2(new_n789), .ZN(new_n790));
  OAI21_X1  g589(.A(new_n686), .B1(new_n787), .B2(new_n790), .ZN(new_n791));
  AOI21_X1  g590(.A(new_n729), .B1(new_n453), .B2(new_n455), .ZN(new_n792));
  NOR2_X1   g591(.A1(new_n791), .A2(new_n792), .ZN(new_n793));
  OAI211_X1 g592(.A(KEYINPUT104), .B(new_n781), .C1(new_n785), .C2(new_n793), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n794), .A2(new_n751), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n700), .A2(new_n701), .ZN(new_n796));
  AOI21_X1  g595(.A(KEYINPUT104), .B1(new_n796), .B2(new_n781), .ZN(new_n797));
  OAI21_X1  g596(.A(new_n780), .B1(new_n795), .B2(new_n797), .ZN(new_n798));
  NAND4_X1  g597(.A1(new_n755), .A2(KEYINPUT109), .A3(new_n794), .A4(new_n751), .ZN(new_n799));
  AOI21_X1  g598(.A(new_n779), .B1(new_n798), .B2(new_n799), .ZN(new_n800));
  AOI21_X1  g599(.A(new_n777), .B1(new_n800), .B2(KEYINPUT111), .ZN(new_n801));
  AOI21_X1  g600(.A(KEYINPUT109), .B1(new_n753), .B2(new_n755), .ZN(new_n802));
  AND4_X1   g601(.A1(KEYINPUT109), .A2(new_n755), .A3(new_n751), .A4(new_n794), .ZN(new_n803));
  OAI21_X1  g602(.A(new_n778), .B1(new_n802), .B2(new_n803), .ZN(new_n804));
  INV_X1    g603(.A(KEYINPUT111), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  AOI21_X1  g605(.A(new_n776), .B1(new_n801), .B2(new_n806), .ZN(new_n807));
  OAI21_X1  g606(.A(new_n774), .B1(new_n807), .B2(KEYINPUT112), .ZN(new_n808));
  INV_X1    g607(.A(KEYINPUT112), .ZN(new_n809));
  AOI211_X1 g608(.A(new_n809), .B(new_n776), .C1(new_n801), .C2(new_n806), .ZN(new_n810));
  OAI21_X1  g609(.A(KEYINPUT52), .B1(new_n808), .B2(new_n810), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n761), .A2(new_n775), .ZN(new_n812));
  INV_X1    g611(.A(KEYINPUT52), .ZN(new_n813));
  NAND3_X1  g612(.A1(new_n812), .A2(new_n774), .A3(new_n813), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n811), .A2(new_n814), .ZN(G1337gat));
  XOR2_X1   g614(.A(KEYINPUT113), .B(G99gat), .Z(new_n816));
  NOR2_X1   g615(.A1(new_n462), .A2(new_n816), .ZN(new_n817));
  NAND3_X1  g616(.A1(new_n763), .A2(new_n764), .A3(new_n817), .ZN(new_n818));
  OAI21_X1  g617(.A(new_n816), .B1(new_n767), .B2(new_n686), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n818), .A2(new_n819), .ZN(G1338gat));
  NAND3_X1  g619(.A1(new_n704), .A2(new_n273), .A3(new_n766), .ZN(new_n821));
  AOI21_X1  g620(.A(KEYINPUT53), .B1(new_n821), .B2(G106gat), .ZN(new_n822));
  NOR3_X1   g621(.A1(new_n694), .A2(G106gat), .A3(new_n729), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n761), .A2(new_n823), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n822), .A2(new_n824), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n801), .A2(new_n806), .ZN(new_n826));
  AOI22_X1  g625(.A1(new_n826), .A2(new_n823), .B1(G106gat), .B2(new_n821), .ZN(new_n827));
  INV_X1    g626(.A(KEYINPUT53), .ZN(new_n828));
  OAI21_X1  g627(.A(new_n825), .B1(new_n827), .B2(new_n828), .ZN(G1339gat));
  NAND2_X1  g628(.A1(new_n673), .A2(new_n705), .ZN(new_n830));
  INV_X1    g629(.A(KEYINPUT55), .ZN(new_n831));
  INV_X1    g630(.A(new_n662), .ZN(new_n832));
  AND2_X1   g631(.A1(new_n658), .A2(new_n659), .ZN(new_n833));
  OAI211_X1 g632(.A(new_n832), .B(new_n652), .C1(new_n833), .C2(KEYINPUT10), .ZN(new_n834));
  AND3_X1   g633(.A1(new_n834), .A2(KEYINPUT54), .A3(new_n663), .ZN(new_n835));
  INV_X1    g634(.A(KEYINPUT54), .ZN(new_n836));
  OAI211_X1 g635(.A(new_n836), .B(new_n653), .C1(new_n660), .C2(new_n662), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n837), .A2(new_n669), .ZN(new_n838));
  OAI21_X1  g637(.A(new_n831), .B1(new_n835), .B2(new_n838), .ZN(new_n839));
  INV_X1    g638(.A(new_n838), .ZN(new_n840));
  NAND3_X1  g639(.A1(new_n834), .A2(KEYINPUT54), .A3(new_n663), .ZN(new_n841));
  NAND3_X1  g640(.A1(new_n840), .A2(KEYINPUT55), .A3(new_n841), .ZN(new_n842));
  NAND3_X1  g641(.A1(new_n839), .A2(new_n671), .A3(new_n842), .ZN(new_n843));
  AOI21_X1  g642(.A(new_n549), .B1(new_n561), .B2(new_n543), .ZN(new_n844));
  NOR2_X1   g643(.A1(new_n548), .A2(new_n550), .ZN(new_n845));
  OAI21_X1  g644(.A(new_n571), .B1(new_n844), .B2(new_n845), .ZN(new_n846));
  NAND3_X1  g645(.A1(new_n564), .A2(new_n573), .A3(new_n567), .ZN(new_n847));
  NAND4_X1  g646(.A1(new_n646), .A2(new_n648), .A3(new_n846), .A4(new_n847), .ZN(new_n848));
  NOR2_X1   g647(.A1(new_n843), .A2(new_n848), .ZN(new_n849));
  NAND2_X1  g648(.A1(new_n847), .A2(new_n846), .ZN(new_n850));
  OAI22_X1  g649(.A1(new_n843), .A2(new_n705), .B1(new_n694), .B2(new_n850), .ZN(new_n851));
  AOI21_X1  g650(.A(new_n849), .B1(new_n851), .B2(new_n649), .ZN(new_n852));
  OAI21_X1  g651(.A(new_n830), .B1(new_n852), .B2(new_n611), .ZN(new_n853));
  AND2_X1   g652(.A1(new_n853), .A2(new_n381), .ZN(new_n854));
  NOR2_X1   g653(.A1(new_n469), .A2(new_n445), .ZN(new_n855));
  AND2_X1   g654(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  AOI21_X1  g655(.A(G113gat), .B1(new_n856), .B2(new_n579), .ZN(new_n857));
  NOR2_X1   g656(.A1(new_n583), .A2(new_n321), .ZN(new_n858));
  AOI21_X1  g657(.A(new_n857), .B1(new_n856), .B2(new_n858), .ZN(G1340gat));
  NAND2_X1  g658(.A1(new_n856), .A2(new_n672), .ZN(new_n860));
  XNOR2_X1  g659(.A(new_n860), .B(G120gat), .ZN(G1341gat));
  NAND2_X1  g660(.A1(new_n856), .A2(new_n611), .ZN(new_n862));
  XNOR2_X1  g661(.A(new_n862), .B(G127gat), .ZN(G1342gat));
  AND2_X1   g662(.A1(new_n856), .A2(new_n781), .ZN(new_n864));
  NOR2_X1   g663(.A1(new_n864), .A2(new_n355), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n864), .A2(new_n328), .ZN(new_n866));
  AOI21_X1  g665(.A(new_n865), .B1(KEYINPUT56), .B2(new_n866), .ZN(new_n867));
  OAI21_X1  g666(.A(new_n867), .B1(KEYINPUT56), .B2(new_n866), .ZN(G1343gat));
  NAND2_X1  g667(.A1(new_n853), .A2(new_n273), .ZN(new_n869));
  INV_X1    g668(.A(new_n869), .ZN(new_n870));
  OAI21_X1  g669(.A(KEYINPUT114), .B1(new_n870), .B2(KEYINPUT57), .ZN(new_n871));
  INV_X1    g670(.A(KEYINPUT114), .ZN(new_n872));
  INV_X1    g671(.A(KEYINPUT57), .ZN(new_n873));
  NAND3_X1  g672(.A1(new_n869), .A2(new_n872), .A3(new_n873), .ZN(new_n874));
  INV_X1    g673(.A(KEYINPUT116), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n842), .A2(new_n671), .ZN(new_n876));
  AOI21_X1  g675(.A(KEYINPUT55), .B1(new_n840), .B2(new_n841), .ZN(new_n877));
  OAI21_X1  g676(.A(new_n875), .B1(new_n876), .B2(new_n877), .ZN(new_n878));
  NAND4_X1  g677(.A1(new_n839), .A2(KEYINPUT116), .A3(new_n671), .A4(new_n842), .ZN(new_n879));
  NAND4_X1  g678(.A1(new_n878), .A2(new_n581), .A3(new_n582), .A4(new_n879), .ZN(new_n880));
  NAND3_X1  g679(.A1(new_n672), .A2(new_n846), .A3(new_n847), .ZN(new_n881));
  XNOR2_X1  g680(.A(new_n881), .B(KEYINPUT115), .ZN(new_n882));
  AOI21_X1  g681(.A(new_n781), .B1(new_n880), .B2(new_n882), .ZN(new_n883));
  OAI21_X1  g682(.A(new_n693), .B1(new_n883), .B2(new_n849), .ZN(new_n884));
  AND2_X1   g683(.A1(new_n884), .A2(new_n830), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n273), .A2(KEYINPUT57), .ZN(new_n886));
  OAI211_X1 g685(.A(new_n871), .B(new_n874), .C1(new_n885), .C2(new_n886), .ZN(new_n887));
  NAND2_X1  g686(.A1(new_n686), .A2(new_n855), .ZN(new_n888));
  INV_X1    g687(.A(new_n888), .ZN(new_n889));
  AND2_X1   g688(.A1(new_n887), .A2(new_n889), .ZN(new_n890));
  AOI21_X1  g689(.A(new_n207), .B1(new_n890), .B2(new_n579), .ZN(new_n891));
  NOR2_X1   g690(.A1(new_n869), .A2(new_n888), .ZN(new_n892));
  INV_X1    g691(.A(new_n583), .ZN(new_n893));
  NAND3_X1  g692(.A1(new_n892), .A2(new_n207), .A3(new_n893), .ZN(new_n894));
  XOR2_X1   g693(.A(new_n894), .B(KEYINPUT117), .Z(new_n895));
  OAI21_X1  g694(.A(KEYINPUT58), .B1(new_n891), .B2(new_n895), .ZN(new_n896));
  NAND2_X1  g695(.A1(new_n887), .A2(new_n889), .ZN(new_n897));
  OAI21_X1  g696(.A(G141gat), .B1(new_n897), .B2(new_n583), .ZN(new_n898));
  XOR2_X1   g697(.A(KEYINPUT118), .B(KEYINPUT58), .Z(new_n899));
  NAND3_X1  g698(.A1(new_n898), .A2(new_n894), .A3(new_n899), .ZN(new_n900));
  NAND2_X1  g699(.A1(new_n896), .A2(new_n900), .ZN(G1344gat));
  OAI21_X1  g700(.A(KEYINPUT120), .B1(new_n869), .B2(new_n873), .ZN(new_n902));
  INV_X1    g701(.A(KEYINPUT120), .ZN(new_n903));
  NAND4_X1  g702(.A1(new_n853), .A2(new_n903), .A3(KEYINPUT57), .A4(new_n273), .ZN(new_n904));
  NAND2_X1  g703(.A1(new_n902), .A2(new_n904), .ZN(new_n905));
  INV_X1    g704(.A(new_n905), .ZN(new_n906));
  NAND2_X1  g705(.A1(new_n673), .A2(new_n583), .ZN(new_n907));
  NAND2_X1  g706(.A1(new_n884), .A2(new_n907), .ZN(new_n908));
  AOI21_X1  g707(.A(KEYINPUT57), .B1(new_n908), .B2(new_n273), .ZN(new_n909));
  INV_X1    g708(.A(new_n909), .ZN(new_n910));
  AOI211_X1 g709(.A(new_n694), .B(new_n888), .C1(new_n906), .C2(new_n910), .ZN(new_n911));
  OAI21_X1  g710(.A(KEYINPUT59), .B1(new_n911), .B2(new_n202), .ZN(new_n912));
  NAND3_X1  g711(.A1(new_n887), .A2(new_n672), .A3(new_n889), .ZN(new_n913));
  INV_X1    g712(.A(KEYINPUT119), .ZN(new_n914));
  NOR2_X1   g713(.A1(new_n257), .A2(KEYINPUT59), .ZN(new_n915));
  AND3_X1   g714(.A1(new_n913), .A2(new_n914), .A3(new_n915), .ZN(new_n916));
  AOI21_X1  g715(.A(new_n914), .B1(new_n913), .B2(new_n915), .ZN(new_n917));
  OAI21_X1  g716(.A(new_n912), .B1(new_n916), .B2(new_n917), .ZN(new_n918));
  NAND3_X1  g717(.A1(new_n892), .A2(new_n257), .A3(new_n672), .ZN(new_n919));
  NAND2_X1  g718(.A1(new_n918), .A2(new_n919), .ZN(G1345gat));
  OAI21_X1  g719(.A(G155gat), .B1(new_n897), .B2(new_n693), .ZN(new_n921));
  INV_X1    g720(.A(G155gat), .ZN(new_n922));
  NAND3_X1  g721(.A1(new_n892), .A2(new_n922), .A3(new_n611), .ZN(new_n923));
  NAND2_X1  g722(.A1(new_n921), .A2(new_n923), .ZN(G1346gat));
  OAI21_X1  g723(.A(G162gat), .B1(new_n897), .B2(new_n649), .ZN(new_n925));
  INV_X1    g724(.A(G162gat), .ZN(new_n926));
  NAND3_X1  g725(.A1(new_n892), .A2(new_n926), .A3(new_n781), .ZN(new_n927));
  NAND2_X1  g726(.A1(new_n925), .A2(new_n927), .ZN(G1347gat));
  NOR2_X1   g727(.A1(new_n470), .A2(new_n676), .ZN(new_n929));
  AND2_X1   g728(.A1(new_n854), .A2(new_n929), .ZN(new_n930));
  AOI21_X1  g729(.A(G169gat), .B1(new_n930), .B2(new_n579), .ZN(new_n931));
  NAND4_X1  g730(.A1(new_n853), .A2(new_n729), .A3(new_n744), .A4(new_n929), .ZN(new_n932));
  XOR2_X1   g731(.A(new_n932), .B(KEYINPUT121), .Z(new_n933));
  NOR2_X1   g732(.A1(new_n583), .A2(new_n277), .ZN(new_n934));
  AOI21_X1  g733(.A(new_n931), .B1(new_n933), .B2(new_n934), .ZN(G1348gat));
  NAND3_X1  g734(.A1(new_n930), .A2(new_n278), .A3(new_n672), .ZN(new_n936));
  AND2_X1   g735(.A1(new_n933), .A2(new_n672), .ZN(new_n937));
  OAI21_X1  g736(.A(new_n936), .B1(new_n937), .B2(new_n278), .ZN(G1349gat));
  NAND3_X1  g737(.A1(new_n930), .A2(new_n315), .A3(new_n611), .ZN(new_n939));
  AND2_X1   g738(.A1(new_n933), .A2(new_n611), .ZN(new_n940));
  OAI21_X1  g739(.A(new_n939), .B1(new_n940), .B2(new_n285), .ZN(new_n941));
  XNOR2_X1  g740(.A(new_n941), .B(KEYINPUT60), .ZN(G1350gat));
  AOI21_X1  g741(.A(new_n286), .B1(new_n933), .B2(new_n781), .ZN(new_n943));
  XOR2_X1   g742(.A(new_n943), .B(KEYINPUT61), .Z(new_n944));
  NAND3_X1  g743(.A1(new_n930), .A2(new_n286), .A3(new_n781), .ZN(new_n945));
  NAND2_X1  g744(.A1(new_n944), .A2(new_n945), .ZN(G1351gat));
  NAND2_X1  g745(.A1(new_n906), .A2(new_n910), .ZN(new_n947));
  AND2_X1   g746(.A1(new_n686), .A2(new_n929), .ZN(new_n948));
  NAND2_X1  g747(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  NAND2_X1  g748(.A1(new_n893), .A2(G197gat), .ZN(new_n950));
  NOR3_X1   g749(.A1(new_n720), .A2(new_n470), .A3(new_n729), .ZN(new_n951));
  AND2_X1   g750(.A1(new_n951), .A2(KEYINPUT122), .ZN(new_n952));
  NOR2_X1   g751(.A1(new_n951), .A2(KEYINPUT122), .ZN(new_n953));
  NOR3_X1   g752(.A1(new_n952), .A2(new_n953), .A3(new_n676), .ZN(new_n954));
  NAND2_X1  g753(.A1(new_n954), .A2(new_n853), .ZN(new_n955));
  NOR2_X1   g754(.A1(new_n955), .A2(new_n705), .ZN(new_n956));
  OAI22_X1  g755(.A1(new_n949), .A2(new_n950), .B1(G197gat), .B2(new_n956), .ZN(new_n957));
  XNOR2_X1  g756(.A(new_n957), .B(KEYINPUT123), .ZN(G1352gat));
  NAND3_X1  g757(.A1(new_n947), .A2(new_n672), .A3(new_n948), .ZN(new_n959));
  NAND2_X1  g758(.A1(new_n959), .A2(G204gat), .ZN(new_n960));
  NOR2_X1   g759(.A1(new_n694), .A2(G204gat), .ZN(new_n961));
  INV_X1    g760(.A(new_n961), .ZN(new_n962));
  OR3_X1    g761(.A1(new_n955), .A2(KEYINPUT124), .A3(new_n962), .ZN(new_n963));
  OAI21_X1  g762(.A(KEYINPUT124), .B1(new_n955), .B2(new_n962), .ZN(new_n964));
  NAND2_X1  g763(.A1(new_n963), .A2(new_n964), .ZN(new_n965));
  XNOR2_X1  g764(.A(new_n965), .B(KEYINPUT62), .ZN(new_n966));
  NAND2_X1  g765(.A1(new_n960), .A2(new_n966), .ZN(new_n967));
  INV_X1    g766(.A(KEYINPUT125), .ZN(new_n968));
  NAND2_X1  g767(.A1(new_n967), .A2(new_n968), .ZN(new_n969));
  NAND3_X1  g768(.A1(new_n960), .A2(new_n966), .A3(KEYINPUT125), .ZN(new_n970));
  NAND2_X1  g769(.A1(new_n969), .A2(new_n970), .ZN(G1353gat));
  OR3_X1    g770(.A1(new_n955), .A2(G211gat), .A3(new_n693), .ZN(new_n972));
  OAI211_X1 g771(.A(new_n611), .B(new_n948), .C1(new_n905), .C2(new_n909), .ZN(new_n973));
  AND3_X1   g772(.A1(new_n973), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n974));
  AOI21_X1  g773(.A(KEYINPUT63), .B1(new_n973), .B2(G211gat), .ZN(new_n975));
  OAI21_X1  g774(.A(new_n972), .B1(new_n974), .B2(new_n975), .ZN(new_n976));
  NAND2_X1  g775(.A1(new_n976), .A2(KEYINPUT126), .ZN(new_n977));
  INV_X1    g776(.A(KEYINPUT126), .ZN(new_n978));
  OAI211_X1 g777(.A(new_n978), .B(new_n972), .C1(new_n974), .C2(new_n975), .ZN(new_n979));
  NAND2_X1  g778(.A1(new_n977), .A2(new_n979), .ZN(G1354gat));
  INV_X1    g779(.A(new_n955), .ZN(new_n981));
  AOI21_X1  g780(.A(G218gat), .B1(new_n981), .B2(new_n781), .ZN(new_n982));
  INV_X1    g781(.A(new_n949), .ZN(new_n983));
  NAND2_X1  g782(.A1(new_n781), .A2(G218gat), .ZN(new_n984));
  XNOR2_X1  g783(.A(new_n984), .B(KEYINPUT127), .ZN(new_n985));
  AOI21_X1  g784(.A(new_n982), .B1(new_n983), .B2(new_n985), .ZN(G1355gat));
endmodule


