

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n340, n341, n342, n343, n344, n345, n346, n347, n348, n349, n350,
         n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361,
         n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372,
         n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383,
         n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394,
         n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405,
         n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416,
         n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427,
         n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438,
         n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449,
         n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460,
         n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471,
         n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482,
         n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493,
         n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504,
         n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515,
         n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526,
         n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537,
         n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
         n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559,
         n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570,
         n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581,
         n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592,
         n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603,
         n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614,
         n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625,
         n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636,
         n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647,
         n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658,
         n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669,
         n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680,
         n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691,
         n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702,
         n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713,
         n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724,
         n725, n726;

  XNOR2_X1 U363 ( .A(n533), .B(n400), .ZN(n665) );
  NOR2_X2 U364 ( .A1(G953), .A2(G237), .ZN(n479) );
  INV_X2 U365 ( .A(G953), .ZN(n715) );
  INV_X1 U366 ( .A(KEYINPUT23), .ZN(n378) );
  OR2_X1 U367 ( .A1(n698), .A2(n473), .ZN(n477) );
  AND2_X2 U368 ( .A1(n565), .A2(n663), .ZN(n617) );
  XNOR2_X2 U369 ( .A(n568), .B(KEYINPUT33), .ZN(n694) );
  AND2_X1 U370 ( .A1(n401), .A2(n402), .ZN(n603) );
  XNOR2_X1 U371 ( .A(n424), .B(G472), .ZN(n598) );
  NOR2_X1 U372 ( .A1(n607), .A2(n606), .ZN(n608) );
  AND2_X1 U373 ( .A1(n353), .A2(n352), .ZN(n351) );
  AND2_X1 U374 ( .A1(n356), .A2(n341), .ZN(n354) );
  XNOR2_X1 U375 ( .A(KEYINPUT77), .B(KEYINPUT8), .ZN(n435) );
  XNOR2_X1 U376 ( .A(n396), .B(G104), .ZN(n395) );
  XNOR2_X1 U377 ( .A(G110), .B(G107), .ZN(n396) );
  XNOR2_X1 U378 ( .A(G101), .B(G146), .ZN(n452) );
  XNOR2_X1 U379 ( .A(n348), .B(n451), .ZN(n713) );
  XNOR2_X1 U380 ( .A(n429), .B(G146), .ZN(n464) );
  INV_X1 U381 ( .A(G125), .ZN(n429) );
  XNOR2_X1 U382 ( .A(n500), .B(KEYINPUT4), .ZN(n397) );
  XNOR2_X1 U383 ( .A(n399), .B(KEYINPUT111), .ZN(n668) );
  OR2_X1 U384 ( .A1(n665), .A2(n664), .ZN(n399) );
  XNOR2_X1 U385 ( .A(n397), .B(n411), .ZN(n348) );
  XNOR2_X1 U386 ( .A(G131), .B(G134), .ZN(n411) );
  XOR2_X1 U387 ( .A(KEYINPUT93), .B(KEYINPUT5), .Z(n419) );
  XNOR2_X1 U388 ( .A(G146), .B(G116), .ZN(n421) );
  XNOR2_X1 U389 ( .A(n377), .B(G137), .ZN(n376) );
  INV_X1 U390 ( .A(KEYINPUT68), .ZN(n377) );
  INV_X1 U391 ( .A(G116), .ZN(n468) );
  XNOR2_X1 U392 ( .A(n409), .B(n416), .ZN(n470) );
  XNOR2_X1 U393 ( .A(G119), .B(G113), .ZN(n416) );
  XNOR2_X1 U394 ( .A(n417), .B(KEYINPUT3), .ZN(n409) );
  XNOR2_X1 U395 ( .A(G101), .B(KEYINPUT66), .ZN(n417) );
  XNOR2_X1 U396 ( .A(n406), .B(G140), .ZN(n451) );
  INV_X1 U397 ( .A(G137), .ZN(n406) );
  XOR2_X1 U398 ( .A(KEYINPUT24), .B(KEYINPUT88), .Z(n432) );
  XNOR2_X1 U399 ( .A(G119), .B(G128), .ZN(n430) );
  XNOR2_X1 U400 ( .A(n464), .B(n408), .ZN(n712) );
  XNOR2_X1 U401 ( .A(KEYINPUT10), .B(KEYINPUT65), .ZN(n408) );
  XNOR2_X1 U402 ( .A(n556), .B(n388), .ZN(n387) );
  INV_X1 U403 ( .A(KEYINPUT107), .ZN(n388) );
  INV_X1 U404 ( .A(KEYINPUT43), .ZN(n385) );
  AND2_X1 U405 ( .A1(n364), .A2(n362), .ZN(n361) );
  AND2_X1 U406 ( .A1(n360), .A2(n577), .ZN(n359) );
  BUF_X1 U407 ( .A(n533), .Z(n559) );
  NAND2_X1 U408 ( .A1(n707), .A2(G469), .ZN(n370) );
  NAND2_X1 U409 ( .A1(n707), .A2(G210), .ZN(n394) );
  XNOR2_X1 U410 ( .A(n693), .B(n413), .ZN(n412) );
  XNOR2_X1 U411 ( .A(KEYINPUT78), .B(KEYINPUT2), .ZN(n413) );
  NAND2_X1 U412 ( .A1(n593), .A2(n592), .ZN(n596) );
  INV_X1 U413 ( .A(G237), .ZN(n474) );
  INV_X1 U414 ( .A(G902), .ZN(n475) );
  XOR2_X1 U415 ( .A(KEYINPUT20), .B(KEYINPUT89), .Z(n426) );
  NAND2_X1 U416 ( .A1(n350), .A2(n355), .ZN(n349) );
  XNOR2_X1 U417 ( .A(n378), .B(G110), .ZN(n431) );
  XOR2_X1 U418 ( .A(KEYINPUT96), .B(KEYINPUT11), .Z(n481) );
  XNOR2_X1 U419 ( .A(G131), .B(G143), .ZN(n487) );
  XNOR2_X1 U420 ( .A(G113), .B(G140), .ZN(n482) );
  XOR2_X1 U421 ( .A(KEYINPUT12), .B(KEYINPUT97), .Z(n483) );
  XNOR2_X1 U422 ( .A(KEYINPUT83), .B(KEYINPUT84), .ZN(n459) );
  XNOR2_X1 U423 ( .A(KEYINPUT17), .B(KEYINPUT70), .ZN(n458) );
  XNOR2_X1 U424 ( .A(KEYINPUT18), .B(KEYINPUT71), .ZN(n462) );
  NAND2_X1 U425 ( .A1(G234), .A2(G237), .ZN(n444) );
  INV_X1 U426 ( .A(KEYINPUT38), .ZN(n400) );
  XNOR2_X1 U427 ( .A(KEYINPUT73), .B(KEYINPUT34), .ZN(n576) );
  INV_X1 U428 ( .A(n576), .ZN(n365) );
  XNOR2_X1 U429 ( .A(n379), .B(KEYINPUT9), .ZN(n496) );
  INV_X1 U430 ( .A(KEYINPUT99), .ZN(n379) );
  XNOR2_X1 U431 ( .A(G134), .B(G122), .ZN(n495) );
  XNOR2_X1 U432 ( .A(KEYINPUT101), .B(KEYINPUT7), .ZN(n493) );
  XOR2_X1 U433 ( .A(KEYINPUT100), .B(KEYINPUT98), .Z(n494) );
  XNOR2_X1 U434 ( .A(n395), .B(n452), .ZN(n454) );
  OR2_X1 U435 ( .A1(n566), .A2(n609), .ZN(n588) );
  NOR2_X1 U436 ( .A1(G902), .A2(n702), .ZN(n492) );
  INV_X1 U437 ( .A(G478), .ZN(n383) );
  NAND2_X1 U438 ( .A1(n382), .A2(n381), .ZN(n543) );
  XNOR2_X1 U439 ( .A(n410), .B(n470), .ZN(n423) );
  XNOR2_X1 U440 ( .A(n617), .B(n398), .ZN(n716) );
  INV_X1 U441 ( .A(n717), .ZN(n398) );
  XNOR2_X1 U442 ( .A(KEYINPUT16), .B(G110), .ZN(n467) );
  AND2_X1 U443 ( .A1(n616), .A2(n715), .ZN(n638) );
  XNOR2_X1 U444 ( .A(n437), .B(n405), .ZN(n404) );
  XNOR2_X1 U445 ( .A(n451), .B(KEYINPUT87), .ZN(n405) );
  XNOR2_X1 U446 ( .A(n386), .B(n384), .ZN(n560) );
  XNOR2_X1 U447 ( .A(n558), .B(n385), .ZN(n384) );
  NOR2_X1 U448 ( .A1(n387), .A2(n557), .ZN(n386) );
  XNOR2_X1 U449 ( .A(n510), .B(n511), .ZN(n722) );
  XNOR2_X1 U450 ( .A(n578), .B(KEYINPUT35), .ZN(n579) );
  NAND2_X1 U451 ( .A1(n361), .A2(n359), .ZN(n580) );
  XNOR2_X1 U452 ( .A(n602), .B(n601), .ZN(n659) );
  XNOR2_X1 U453 ( .A(n543), .B(n380), .ZN(n655) );
  INV_X1 U454 ( .A(KEYINPUT106), .ZN(n380) );
  INV_X1 U455 ( .A(KEYINPUT60), .ZN(n371) );
  INV_X1 U456 ( .A(KEYINPUT124), .ZN(n367) );
  NAND2_X1 U457 ( .A1(n369), .A2(n391), .ZN(n368) );
  XNOR2_X1 U458 ( .A(n370), .B(n345), .ZN(n369) );
  INV_X1 U459 ( .A(KEYINPUT56), .ZN(n389) );
  NAND2_X1 U460 ( .A1(n392), .A2(n391), .ZN(n390) );
  XNOR2_X1 U461 ( .A(n394), .B(n393), .ZN(n392) );
  AND2_X1 U462 ( .A1(n412), .A2(n340), .ZN(n696) );
  XNOR2_X1 U463 ( .A(n492), .B(n491), .ZN(n529) );
  INV_X1 U464 ( .A(n529), .ZN(n381) );
  NOR2_X1 U465 ( .A1(n695), .A2(n344), .ZN(n340) );
  AND2_X1 U466 ( .A1(n357), .A2(KEYINPUT82), .ZN(n341) );
  NOR2_X1 U467 ( .A1(n605), .A2(n604), .ZN(n342) );
  XNOR2_X1 U468 ( .A(n506), .B(n383), .ZN(n528) );
  INV_X1 U469 ( .A(n528), .ZN(n382) );
  OR2_X1 U470 ( .A1(n594), .A2(n596), .ZN(n343) );
  AND2_X1 U471 ( .A1(n694), .A2(n685), .ZN(n344) );
  INV_X1 U472 ( .A(KEYINPUT82), .ZN(n355) );
  XNOR2_X1 U473 ( .A(n628), .B(n627), .ZN(n345) );
  XNOR2_X1 U474 ( .A(KEYINPUT62), .B(n623), .ZN(n346) );
  XNOR2_X1 U475 ( .A(n702), .B(KEYINPUT59), .ZN(n347) );
  INV_X1 U476 ( .A(n711), .ZN(n391) );
  XNOR2_X1 U477 ( .A(n423), .B(n348), .ZN(n623) );
  XNOR2_X1 U478 ( .A(n608), .B(KEYINPUT103), .ZN(n356) );
  NAND2_X1 U479 ( .A1(n351), .A2(n349), .ZN(n613) );
  NAND2_X1 U480 ( .A1(n358), .A2(n357), .ZN(n350) );
  OR2_X1 U481 ( .A1(n356), .A2(KEYINPUT82), .ZN(n352) );
  NAND2_X1 U482 ( .A1(n354), .A2(n358), .ZN(n353) );
  INV_X1 U483 ( .A(n643), .ZN(n357) );
  NAND2_X1 U484 ( .A1(n724), .A2(KEYINPUT44), .ZN(n358) );
  NAND2_X1 U485 ( .A1(n605), .A2(n365), .ZN(n360) );
  NAND2_X1 U486 ( .A1(n363), .A2(n694), .ZN(n362) );
  AND2_X1 U487 ( .A1(n581), .A2(n576), .ZN(n363) );
  NAND2_X1 U488 ( .A1(n366), .A2(n365), .ZN(n364) );
  INV_X1 U489 ( .A(n694), .ZN(n366) );
  XNOR2_X1 U490 ( .A(n368), .B(n367), .ZN(G54) );
  NOR2_X1 U491 ( .A1(n518), .A2(n517), .ZN(n519) );
  XNOR2_X1 U492 ( .A(n372), .B(n371), .ZN(G60) );
  NAND2_X1 U493 ( .A1(n375), .A2(n391), .ZN(n372) );
  XNOR2_X1 U494 ( .A(n373), .B(KEYINPUT63), .ZN(G57) );
  NAND2_X1 U495 ( .A1(n374), .A2(n391), .ZN(n373) );
  NOR2_X1 U496 ( .A1(n525), .A2(n665), .ZN(n520) );
  XNOR2_X1 U497 ( .A(n624), .B(n346), .ZN(n374) );
  XNOR2_X1 U498 ( .A(n703), .B(n347), .ZN(n375) );
  INV_X1 U499 ( .A(n692), .ZN(n620) );
  XNOR2_X1 U500 ( .A(n376), .B(n421), .ZN(n422) );
  NAND2_X1 U501 ( .A1(n516), .A2(n603), .ZN(n518) );
  XNOR2_X1 U502 ( .A(n519), .B(KEYINPUT69), .ZN(n525) );
  NAND2_X1 U503 ( .A1(n692), .A2(KEYINPUT79), .ZN(n619) );
  NAND2_X2 U504 ( .A1(n617), .A2(n616), .ZN(n692) );
  NOR2_X2 U505 ( .A1(n566), .A2(n403), .ZN(n599) );
  XNOR2_X1 U506 ( .A(n397), .B(n460), .ZN(n466) );
  NOR2_X1 U507 ( .A1(n726), .A2(n722), .ZN(n522) );
  XNOR2_X1 U508 ( .A(n521), .B(KEYINPUT40), .ZN(n726) );
  XNOR2_X2 U509 ( .A(n620), .B(KEYINPUT2), .ZN(n621) );
  XNOR2_X1 U510 ( .A(n420), .B(n422), .ZN(n410) );
  INV_X1 U511 ( .A(n598), .ZN(n512) );
  NAND2_X1 U512 ( .A1(n598), .A2(n546), .ZN(n514) );
  INV_X1 U513 ( .A(n403), .ZN(n402) );
  XNOR2_X1 U514 ( .A(n434), .B(n712), .ZN(n407) );
  XNOR2_X1 U515 ( .A(n407), .B(n404), .ZN(n708) );
  XNOR2_X2 U516 ( .A(n542), .B(KEYINPUT1), .ZN(n566) );
  XNOR2_X2 U517 ( .A(n456), .B(G469), .ZN(n542) );
  XNOR2_X2 U518 ( .A(n615), .B(KEYINPUT45), .ZN(n616) );
  XNOR2_X1 U519 ( .A(n390), .B(n389), .ZN(G51) );
  INV_X1 U520 ( .A(n701), .ZN(n393) );
  XNOR2_X2 U521 ( .A(n619), .B(n618), .ZN(n622) );
  INV_X1 U522 ( .A(n542), .ZN(n401) );
  NAND2_X1 U523 ( .A1(n566), .A2(n403), .ZN(n674) );
  NAND2_X1 U524 ( .A1(n515), .A2(n675), .ZN(n403) );
  XNOR2_X2 U525 ( .A(G143), .B(G128), .ZN(n500) );
  AND2_X1 U526 ( .A1(n566), .A2(n512), .ZN(n414) );
  AND2_X1 U527 ( .A1(n666), .A2(n675), .ZN(n415) );
  AND2_X1 U528 ( .A1(n551), .A2(n550), .ZN(n552) );
  INV_X1 U529 ( .A(n725), .ZN(n592) );
  INV_X1 U530 ( .A(KEYINPUT48), .ZN(n554) );
  INV_X1 U531 ( .A(KEYINPUT30), .ZN(n513) );
  XNOR2_X1 U532 ( .A(n713), .B(n455), .ZN(n626) );
  XNOR2_X1 U533 ( .A(n514), .B(n513), .ZN(n516) );
  XNOR2_X1 U534 ( .A(n433), .B(n432), .ZN(n434) );
  NAND2_X1 U535 ( .A1(n583), .A2(n414), .ZN(n585) );
  XOR2_X1 U536 ( .A(KEYINPUT114), .B(KEYINPUT42), .Z(n511) );
  NAND2_X1 U537 ( .A1(n479), .A2(G210), .ZN(n418) );
  XNOR2_X1 U538 ( .A(n419), .B(n418), .ZN(n420) );
  NAND2_X1 U539 ( .A1(n623), .A2(n475), .ZN(n424) );
  XNOR2_X2 U540 ( .A(KEYINPUT15), .B(G902), .ZN(n618) );
  NAND2_X1 U541 ( .A1(G234), .A2(n618), .ZN(n425) );
  XNOR2_X1 U542 ( .A(n426), .B(n425), .ZN(n438) );
  AND2_X1 U543 ( .A1(n438), .A2(G221), .ZN(n428) );
  XNOR2_X1 U544 ( .A(KEYINPUT92), .B(KEYINPUT21), .ZN(n427) );
  XNOR2_X1 U545 ( .A(n428), .B(n427), .ZN(n675) );
  XNOR2_X1 U546 ( .A(n431), .B(n430), .ZN(n433) );
  NAND2_X1 U547 ( .A1(n715), .A2(G234), .ZN(n436) );
  XNOR2_X1 U548 ( .A(n436), .B(n435), .ZN(n499) );
  NAND2_X1 U549 ( .A1(G221), .A2(n499), .ZN(n437) );
  NOR2_X1 U550 ( .A1(n708), .A2(G902), .ZN(n443) );
  XOR2_X1 U551 ( .A(KEYINPUT25), .B(KEYINPUT91), .Z(n440) );
  NAND2_X1 U552 ( .A1(G217), .A2(n438), .ZN(n439) );
  XNOR2_X1 U553 ( .A(n440), .B(n439), .ZN(n441) );
  XNOR2_X1 U554 ( .A(n441), .B(KEYINPUT90), .ZN(n442) );
  XNOR2_X1 U555 ( .A(n443), .B(n442), .ZN(n515) );
  INV_X1 U556 ( .A(n515), .ZN(n586) );
  INV_X1 U557 ( .A(n586), .ZN(n676) );
  XNOR2_X1 U558 ( .A(KEYINPUT14), .B(n444), .ZN(n446) );
  NAND2_X1 U559 ( .A1(G902), .A2(n446), .ZN(n569) );
  OR2_X1 U560 ( .A1(n715), .A2(n569), .ZN(n445) );
  NOR2_X1 U561 ( .A1(G900), .A2(n445), .ZN(n447) );
  NAND2_X1 U562 ( .A1(G952), .A2(n446), .ZN(n691) );
  NOR2_X1 U563 ( .A1(G953), .A2(n691), .ZN(n571) );
  NOR2_X1 U564 ( .A1(n447), .A2(n571), .ZN(n517) );
  NOR2_X1 U565 ( .A1(n676), .A2(n517), .ZN(n448) );
  NAND2_X1 U566 ( .A1(n675), .A2(n448), .ZN(n545) );
  NOR2_X1 U567 ( .A1(n512), .A2(n545), .ZN(n450) );
  XNOR2_X1 U568 ( .A(KEYINPUT110), .B(KEYINPUT28), .ZN(n449) );
  XOR2_X1 U569 ( .A(n450), .B(n449), .Z(n457) );
  NAND2_X1 U570 ( .A1(G227), .A2(n715), .ZN(n453) );
  XNOR2_X1 U571 ( .A(n454), .B(n453), .ZN(n455) );
  NOR2_X1 U572 ( .A1(n626), .A2(G902), .ZN(n456) );
  NOR2_X1 U573 ( .A1(n457), .A2(n542), .ZN(n535) );
  XNOR2_X1 U574 ( .A(n459), .B(n458), .ZN(n460) );
  NAND2_X1 U575 ( .A1(n715), .A2(G224), .ZN(n461) );
  XNOR2_X1 U576 ( .A(n462), .B(n461), .ZN(n463) );
  XNOR2_X1 U577 ( .A(n464), .B(n463), .ZN(n465) );
  XNOR2_X1 U578 ( .A(n466), .B(n465), .ZN(n472) );
  XNOR2_X2 U579 ( .A(G122), .B(G104), .ZN(n486) );
  XNOR2_X1 U580 ( .A(n486), .B(n467), .ZN(n469) );
  XNOR2_X1 U581 ( .A(n468), .B(G107), .ZN(n501) );
  XNOR2_X1 U582 ( .A(n469), .B(n501), .ZN(n471) );
  XNOR2_X1 U583 ( .A(n471), .B(n470), .ZN(n640) );
  XNOR2_X1 U584 ( .A(n472), .B(n640), .ZN(n698) );
  INV_X1 U585 ( .A(n618), .ZN(n473) );
  NAND2_X1 U586 ( .A1(n475), .A2(n474), .ZN(n478) );
  NAND2_X1 U587 ( .A1(n478), .A2(G210), .ZN(n476) );
  XNOR2_X2 U588 ( .A(n477), .B(n476), .ZN(n533) );
  NAND2_X1 U589 ( .A1(n478), .A2(G214), .ZN(n546) );
  NAND2_X1 U590 ( .A1(G214), .A2(n479), .ZN(n480) );
  XNOR2_X1 U591 ( .A(n481), .B(n480), .ZN(n485) );
  XNOR2_X1 U592 ( .A(n483), .B(n482), .ZN(n484) );
  XOR2_X1 U593 ( .A(n485), .B(n484), .Z(n490) );
  XOR2_X1 U594 ( .A(n487), .B(n486), .Z(n488) );
  XNOR2_X1 U595 ( .A(n712), .B(n488), .ZN(n489) );
  XNOR2_X1 U596 ( .A(n490), .B(n489), .ZN(n702) );
  XOR2_X1 U597 ( .A(KEYINPUT13), .B(G475), .Z(n491) );
  XNOR2_X1 U598 ( .A(n494), .B(n493), .ZN(n498) );
  XNOR2_X1 U599 ( .A(n496), .B(n495), .ZN(n497) );
  XOR2_X1 U600 ( .A(n498), .B(n497), .Z(n505) );
  NAND2_X1 U601 ( .A1(n499), .A2(G217), .ZN(n503) );
  XNOR2_X1 U602 ( .A(n500), .B(n501), .ZN(n502) );
  XNOR2_X1 U603 ( .A(n503), .B(n502), .ZN(n504) );
  XNOR2_X1 U604 ( .A(n505), .B(n504), .ZN(n704) );
  NOR2_X1 U605 ( .A1(n704), .A2(G902), .ZN(n506) );
  AND2_X1 U606 ( .A1(n529), .A2(n382), .ZN(n666) );
  NAND2_X1 U607 ( .A1(n668), .A2(n666), .ZN(n509) );
  XOR2_X1 U608 ( .A(KEYINPUT112), .B(KEYINPUT113), .Z(n507) );
  XNOR2_X1 U609 ( .A(KEYINPUT41), .B(n507), .ZN(n508) );
  XNOR2_X2 U610 ( .A(n509), .B(n508), .ZN(n685) );
  NAND2_X1 U611 ( .A1(n535), .A2(n685), .ZN(n510) );
  XNOR2_X1 U612 ( .A(n520), .B(KEYINPUT39), .ZN(n564) );
  NOR2_X1 U613 ( .A1(n564), .A2(n543), .ZN(n521) );
  XNOR2_X1 U614 ( .A(n522), .B(KEYINPUT46), .ZN(n553) );
  NAND2_X1 U615 ( .A1(n381), .A2(n528), .ZN(n523) );
  XNOR2_X1 U616 ( .A(KEYINPUT105), .B(n523), .ZN(n577) );
  INV_X1 U617 ( .A(n577), .ZN(n524) );
  NOR2_X1 U618 ( .A1(n525), .A2(n524), .ZN(n527) );
  INV_X1 U619 ( .A(n559), .ZN(n526) );
  NAND2_X1 U620 ( .A1(n527), .A2(n526), .ZN(n630) );
  AND2_X1 U621 ( .A1(n529), .A2(n528), .ZN(n658) );
  INV_X1 U622 ( .A(n658), .ZN(n563) );
  NAND2_X1 U623 ( .A1(n563), .A2(n543), .ZN(n530) );
  XNOR2_X1 U624 ( .A(KEYINPUT102), .B(n530), .ZN(n669) );
  INV_X1 U625 ( .A(n669), .ZN(n606) );
  NAND2_X1 U626 ( .A1(KEYINPUT47), .A2(n606), .ZN(n531) );
  NAND2_X1 U627 ( .A1(n630), .A2(n531), .ZN(n532) );
  XNOR2_X1 U628 ( .A(n532), .B(KEYINPUT75), .ZN(n540) );
  INV_X1 U629 ( .A(n546), .ZN(n664) );
  OR2_X1 U630 ( .A1(n533), .A2(n664), .ZN(n534) );
  XNOR2_X2 U631 ( .A(n534), .B(KEYINPUT19), .ZN(n574) );
  NAND2_X1 U632 ( .A1(n535), .A2(n574), .ZN(n536) );
  XNOR2_X1 U633 ( .A(n536), .B(KEYINPUT47), .ZN(n538) );
  INV_X1 U634 ( .A(n536), .ZN(n651) );
  NAND2_X1 U635 ( .A1(n651), .A2(n606), .ZN(n537) );
  NAND2_X1 U636 ( .A1(n538), .A2(n537), .ZN(n539) );
  NAND2_X1 U637 ( .A1(n540), .A2(n539), .ZN(n541) );
  XNOR2_X1 U638 ( .A(n541), .B(KEYINPUT67), .ZN(n551) );
  INV_X1 U639 ( .A(n566), .ZN(n557) );
  XNOR2_X1 U640 ( .A(n512), .B(KEYINPUT6), .ZN(n609) );
  NAND2_X1 U641 ( .A1(n609), .A2(n655), .ZN(n544) );
  NOR2_X1 U642 ( .A1(n545), .A2(n544), .ZN(n547) );
  NAND2_X1 U643 ( .A1(n547), .A2(n546), .ZN(n556) );
  NOR2_X1 U644 ( .A1(n556), .A2(n559), .ZN(n548) );
  XOR2_X1 U645 ( .A(KEYINPUT36), .B(n548), .Z(n549) );
  NOR2_X1 U646 ( .A1(n566), .A2(n549), .ZN(n661) );
  INV_X1 U647 ( .A(n661), .ZN(n550) );
  NAND2_X1 U648 ( .A1(n553), .A2(n552), .ZN(n555) );
  XNOR2_X1 U649 ( .A(n555), .B(n554), .ZN(n561) );
  XOR2_X1 U650 ( .A(KEYINPUT108), .B(KEYINPUT109), .Z(n558) );
  NAND2_X1 U651 ( .A1(n560), .A2(n559), .ZN(n632) );
  NAND2_X1 U652 ( .A1(n561), .A2(n632), .ZN(n562) );
  XNOR2_X1 U653 ( .A(n562), .B(KEYINPUT81), .ZN(n565) );
  OR2_X1 U654 ( .A1(n564), .A2(n563), .ZN(n663) );
  XNOR2_X1 U655 ( .A(n599), .B(KEYINPUT104), .ZN(n567) );
  NAND2_X1 U656 ( .A1(n567), .A2(n609), .ZN(n568) );
  XNOR2_X1 U657 ( .A(KEYINPUT85), .B(G898), .ZN(n635) );
  NAND2_X1 U658 ( .A1(G953), .A2(n635), .ZN(n639) );
  NOR2_X1 U659 ( .A1(n569), .A2(n639), .ZN(n570) );
  OR2_X1 U660 ( .A1(n571), .A2(n570), .ZN(n572) );
  XNOR2_X1 U661 ( .A(n572), .B(KEYINPUT86), .ZN(n573) );
  NAND2_X1 U662 ( .A1(n574), .A2(n573), .ZN(n575) );
  XNOR2_X2 U663 ( .A(n575), .B(KEYINPUT0), .ZN(n605) );
  XNOR2_X1 U664 ( .A(KEYINPUT80), .B(KEYINPUT72), .ZN(n578) );
  XNOR2_X2 U665 ( .A(n580), .B(n579), .ZN(n724) );
  NOR2_X1 U666 ( .A1(n724), .A2(KEYINPUT44), .ZN(n594) );
  INV_X1 U667 ( .A(n605), .ZN(n581) );
  NAND2_X1 U668 ( .A1(n581), .A2(n415), .ZN(n582) );
  XNOR2_X1 U669 ( .A(n582), .B(KEYINPUT22), .ZN(n612) );
  INV_X1 U670 ( .A(n612), .ZN(n583) );
  INV_X1 U671 ( .A(KEYINPUT64), .ZN(n584) );
  XNOR2_X1 U672 ( .A(n585), .B(n584), .ZN(n587) );
  AND2_X1 U673 ( .A1(n587), .A2(n586), .ZN(n631) );
  INV_X1 U674 ( .A(n631), .ZN(n593) );
  NOR2_X1 U675 ( .A1(n676), .A2(n588), .ZN(n589) );
  XOR2_X1 U676 ( .A(KEYINPUT74), .B(n589), .Z(n590) );
  NOR2_X1 U677 ( .A1(n590), .A2(n612), .ZN(n591) );
  XNOR2_X1 U678 ( .A(n591), .B(KEYINPUT32), .ZN(n725) );
  INV_X1 U679 ( .A(KEYINPUT44), .ZN(n595) );
  NAND2_X1 U680 ( .A1(n596), .A2(n595), .ZN(n597) );
  NAND2_X1 U681 ( .A1(n343), .A2(n597), .ZN(n614) );
  NAND2_X1 U682 ( .A1(n599), .A2(n598), .ZN(n600) );
  XNOR2_X1 U683 ( .A(n600), .B(KEYINPUT94), .ZN(n673) );
  NOR2_X1 U684 ( .A1(n673), .A2(n605), .ZN(n602) );
  XNOR2_X1 U685 ( .A(KEYINPUT31), .B(KEYINPUT95), .ZN(n601) );
  NAND2_X1 U686 ( .A1(n603), .A2(n512), .ZN(n604) );
  NOR2_X1 U687 ( .A1(n659), .A2(n342), .ZN(n607) );
  NAND2_X1 U688 ( .A1(n566), .A2(n676), .ZN(n610) );
  OR2_X1 U689 ( .A1(n610), .A2(n609), .ZN(n611) );
  NOR2_X1 U690 ( .A1(n612), .A2(n611), .ZN(n643) );
  NAND2_X1 U691 ( .A1(n614), .A2(n613), .ZN(n615) );
  NOR2_X4 U692 ( .A1(n622), .A2(n621), .ZN(n707) );
  NAND2_X1 U693 ( .A1(n707), .A2(G472), .ZN(n624) );
  INV_X1 U694 ( .A(G952), .ZN(n625) );
  AND2_X1 U695 ( .A1(n625), .A2(G953), .ZN(n711) );
  XOR2_X1 U696 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n628) );
  XNOR2_X1 U697 ( .A(n626), .B(KEYINPUT123), .ZN(n627) );
  XNOR2_X1 U698 ( .A(G143), .B(KEYINPUT116), .ZN(n629) );
  XNOR2_X1 U699 ( .A(n630), .B(n629), .ZN(G45) );
  XOR2_X1 U700 ( .A(n631), .B(G110), .Z(G12) );
  XNOR2_X1 U701 ( .A(n632), .B(G140), .ZN(G42) );
  NAND2_X1 U702 ( .A1(G953), .A2(G224), .ZN(n633) );
  XOR2_X1 U703 ( .A(KEYINPUT61), .B(n633), .Z(n634) );
  NOR2_X1 U704 ( .A1(n635), .A2(n634), .ZN(n636) );
  XOR2_X1 U705 ( .A(KEYINPUT125), .B(n636), .Z(n637) );
  NOR2_X1 U706 ( .A1(n638), .A2(n637), .ZN(n642) );
  NAND2_X1 U707 ( .A1(n640), .A2(n639), .ZN(n641) );
  XNOR2_X1 U708 ( .A(n642), .B(n641), .ZN(G69) );
  XOR2_X1 U709 ( .A(G101), .B(n643), .Z(G3) );
  NAND2_X1 U710 ( .A1(n655), .A2(n342), .ZN(n644) );
  XNOR2_X1 U711 ( .A(n644), .B(G104), .ZN(G6) );
  XOR2_X1 U712 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n646) );
  NAND2_X1 U713 ( .A1(n342), .A2(n658), .ZN(n645) );
  XNOR2_X1 U714 ( .A(n646), .B(n645), .ZN(n647) );
  XNOR2_X1 U715 ( .A(G107), .B(n647), .ZN(G9) );
  XOR2_X1 U716 ( .A(KEYINPUT115), .B(KEYINPUT29), .Z(n649) );
  NAND2_X1 U717 ( .A1(n651), .A2(n658), .ZN(n648) );
  XNOR2_X1 U718 ( .A(n649), .B(n648), .ZN(n650) );
  XOR2_X1 U719 ( .A(G128), .B(n650), .Z(G30) );
  XOR2_X1 U720 ( .A(KEYINPUT117), .B(KEYINPUT118), .Z(n653) );
  NAND2_X1 U721 ( .A1(n651), .A2(n655), .ZN(n652) );
  XNOR2_X1 U722 ( .A(n653), .B(n652), .ZN(n654) );
  XNOR2_X1 U723 ( .A(G146), .B(n654), .ZN(G48) );
  XOR2_X1 U724 ( .A(G113), .B(KEYINPUT119), .Z(n657) );
  NAND2_X1 U725 ( .A1(n659), .A2(n655), .ZN(n656) );
  XNOR2_X1 U726 ( .A(n657), .B(n656), .ZN(G15) );
  NAND2_X1 U727 ( .A1(n659), .A2(n658), .ZN(n660) );
  XNOR2_X1 U728 ( .A(n660), .B(G116), .ZN(G18) );
  XNOR2_X1 U729 ( .A(G125), .B(n661), .ZN(n662) );
  XNOR2_X1 U730 ( .A(n662), .B(KEYINPUT37), .ZN(G27) );
  XNOR2_X1 U731 ( .A(G134), .B(n663), .ZN(G36) );
  NAND2_X1 U732 ( .A1(n665), .A2(n664), .ZN(n667) );
  NAND2_X1 U733 ( .A1(n667), .A2(n666), .ZN(n671) );
  NAND2_X1 U734 ( .A1(n669), .A2(n668), .ZN(n670) );
  NAND2_X1 U735 ( .A1(n671), .A2(n670), .ZN(n672) );
  NAND2_X1 U736 ( .A1(n694), .A2(n672), .ZN(n688) );
  XNOR2_X1 U737 ( .A(KEYINPUT50), .B(n674), .ZN(n682) );
  XNOR2_X1 U738 ( .A(KEYINPUT120), .B(KEYINPUT49), .ZN(n678) );
  NOR2_X1 U739 ( .A1(n676), .A2(n675), .ZN(n677) );
  XNOR2_X1 U740 ( .A(n678), .B(n677), .ZN(n679) );
  NAND2_X1 U741 ( .A1(n679), .A2(n512), .ZN(n680) );
  XNOR2_X1 U742 ( .A(KEYINPUT121), .B(n680), .ZN(n681) );
  NAND2_X1 U743 ( .A1(n682), .A2(n681), .ZN(n683) );
  NAND2_X1 U744 ( .A1(n673), .A2(n683), .ZN(n684) );
  XOR2_X1 U745 ( .A(KEYINPUT51), .B(n684), .Z(n686) );
  NAND2_X1 U746 ( .A1(n686), .A2(n685), .ZN(n687) );
  NAND2_X1 U747 ( .A1(n688), .A2(n687), .ZN(n689) );
  XOR2_X1 U748 ( .A(KEYINPUT52), .B(n689), .Z(n690) );
  NOR2_X1 U749 ( .A1(n691), .A2(n690), .ZN(n695) );
  NAND2_X1 U750 ( .A1(n692), .A2(KEYINPUT76), .ZN(n693) );
  NAND2_X1 U751 ( .A1(n715), .A2(n696), .ZN(n697) );
  XOR2_X1 U752 ( .A(KEYINPUT53), .B(n697), .Z(G75) );
  XNOR2_X1 U753 ( .A(KEYINPUT54), .B(KEYINPUT122), .ZN(n699) );
  XOR2_X1 U754 ( .A(n699), .B(KEYINPUT55), .Z(n700) );
  XNOR2_X1 U755 ( .A(n698), .B(n700), .ZN(n701) );
  NAND2_X1 U756 ( .A1(n707), .A2(G475), .ZN(n703) );
  NAND2_X1 U757 ( .A1(n707), .A2(G478), .ZN(n705) );
  XNOR2_X1 U758 ( .A(n705), .B(n704), .ZN(n706) );
  NOR2_X1 U759 ( .A1(n711), .A2(n706), .ZN(G63) );
  NAND2_X1 U760 ( .A1(n707), .A2(G217), .ZN(n709) );
  XNOR2_X1 U761 ( .A(n709), .B(n708), .ZN(n710) );
  NOR2_X1 U762 ( .A1(n711), .A2(n710), .ZN(G66) );
  XNOR2_X1 U763 ( .A(n712), .B(KEYINPUT126), .ZN(n714) );
  XNOR2_X1 U764 ( .A(n714), .B(n713), .ZN(n717) );
  NAND2_X1 U765 ( .A1(n716), .A2(n715), .ZN(n721) );
  XNOR2_X1 U766 ( .A(G227), .B(n717), .ZN(n718) );
  NAND2_X1 U767 ( .A1(n718), .A2(G900), .ZN(n719) );
  NAND2_X1 U768 ( .A1(G953), .A2(n719), .ZN(n720) );
  NAND2_X1 U769 ( .A1(n721), .A2(n720), .ZN(G72) );
  XNOR2_X1 U770 ( .A(n722), .B(G137), .ZN(n723) );
  XNOR2_X1 U771 ( .A(n723), .B(KEYINPUT127), .ZN(G39) );
  XOR2_X1 U772 ( .A(n724), .B(G122), .Z(G24) );
  XOR2_X1 U773 ( .A(n725), .B(G119), .Z(G21) );
  XOR2_X1 U774 ( .A(n726), .B(G131), .Z(G33) );
endmodule

