//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 1 1 0 0 0 0 1 1 1 0 1 0 1 1 0 0 1 0 0 0 0 0 0 1 1 1 1 1 0 0 1 0 1 0 1 1 0 0 1 1 0 0 1 0 0 1 1 1 1 1 1 0 0 0 0 1 0 1 0 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:16:03 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n686, new_n687, new_n688, new_n689, new_n690, new_n691, new_n692,
    new_n693, new_n694, new_n696, new_n697, new_n698, new_n699, new_n700,
    new_n701, new_n702, new_n703, new_n705, new_n706, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n730, new_n731,
    new_n732, new_n733, new_n734, new_n735, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n771,
    new_n772, new_n773, new_n774, new_n776, new_n777, new_n779, new_n780,
    new_n781, new_n782, new_n783, new_n784, new_n785, new_n786, new_n787,
    new_n788, new_n789, new_n790, new_n791, new_n792, new_n793, new_n794,
    new_n795, new_n796, new_n797, new_n798, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n810,
    new_n811, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n866, new_n867, new_n868, new_n870,
    new_n871, new_n872, new_n873, new_n875, new_n876, new_n877, new_n878,
    new_n879, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n924, new_n925, new_n927, new_n928, new_n929, new_n930, new_n931,
    new_n932, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n942, new_n943, new_n945, new_n946, new_n947, new_n949,
    new_n950, new_n951, new_n953, new_n954, new_n955, new_n956, new_n957,
    new_n958, new_n959, new_n960, new_n962, new_n963, new_n964, new_n965,
    new_n967, new_n968, new_n969, new_n970, new_n971, new_n972, new_n973,
    new_n974, new_n975, new_n976, new_n978, new_n979, new_n980;
  XNOR2_X1  g000(.A(G1gat), .B(G29gat), .ZN(new_n202));
  XNOR2_X1  g001(.A(new_n202), .B(KEYINPUT0), .ZN(new_n203));
  XNOR2_X1  g002(.A(G57gat), .B(G85gat), .ZN(new_n204));
  XNOR2_X1  g003(.A(new_n203), .B(new_n204), .ZN(new_n205));
  NAND2_X1  g004(.A1(G155gat), .A2(G162gat), .ZN(new_n206));
  NAND2_X1  g005(.A1(new_n206), .A2(KEYINPUT2), .ZN(new_n207));
  INV_X1    g006(.A(G141gat), .ZN(new_n208));
  NOR2_X1   g007(.A1(new_n208), .A2(G148gat), .ZN(new_n209));
  INV_X1    g008(.A(G148gat), .ZN(new_n210));
  NOR2_X1   g009(.A1(new_n210), .A2(G141gat), .ZN(new_n211));
  OAI211_X1 g010(.A(KEYINPUT74), .B(new_n207), .C1(new_n209), .C2(new_n211), .ZN(new_n212));
  XNOR2_X1  g011(.A(G155gat), .B(G162gat), .ZN(new_n213));
  INV_X1    g012(.A(new_n213), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n212), .A2(new_n214), .ZN(new_n215));
  AND2_X1   g014(.A1(KEYINPUT66), .A2(G127gat), .ZN(new_n216));
  NOR2_X1   g015(.A1(KEYINPUT66), .A2(G127gat), .ZN(new_n217));
  OAI21_X1  g016(.A(G134gat), .B1(new_n216), .B2(new_n217), .ZN(new_n218));
  NOR2_X1   g017(.A1(G127gat), .A2(G134gat), .ZN(new_n219));
  INV_X1    g018(.A(new_n219), .ZN(new_n220));
  XNOR2_X1  g019(.A(G113gat), .B(G120gat), .ZN(new_n221));
  OAI211_X1 g020(.A(new_n218), .B(new_n220), .C1(KEYINPUT1), .C2(new_n221), .ZN(new_n222));
  INV_X1    g021(.A(KEYINPUT74), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n210), .A2(G141gat), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n208), .A2(G148gat), .ZN(new_n225));
  AOI21_X1  g024(.A(new_n223), .B1(new_n224), .B2(new_n225), .ZN(new_n226));
  NAND3_X1  g025(.A1(new_n226), .A2(new_n213), .A3(new_n207), .ZN(new_n227));
  INV_X1    g026(.A(G120gat), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n228), .A2(G113gat), .ZN(new_n229));
  INV_X1    g028(.A(G113gat), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n230), .A2(G120gat), .ZN(new_n231));
  AOI21_X1  g030(.A(KEYINPUT1), .B1(new_n229), .B2(new_n231), .ZN(new_n232));
  XNOR2_X1  g031(.A(G127gat), .B(G134gat), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n232), .A2(new_n233), .ZN(new_n234));
  NAND4_X1  g033(.A1(new_n215), .A2(new_n222), .A3(new_n227), .A4(new_n234), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n235), .A2(KEYINPUT77), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n229), .A2(new_n231), .ZN(new_n237));
  INV_X1    g036(.A(KEYINPUT1), .ZN(new_n238));
  AOI21_X1  g037(.A(new_n219), .B1(new_n237), .B2(new_n238), .ZN(new_n239));
  AOI22_X1  g038(.A1(new_n239), .A2(new_n218), .B1(new_n233), .B2(new_n232), .ZN(new_n240));
  INV_X1    g039(.A(KEYINPUT77), .ZN(new_n241));
  NAND4_X1  g040(.A1(new_n240), .A2(new_n241), .A3(new_n227), .A4(new_n215), .ZN(new_n242));
  AOI21_X1  g041(.A(KEYINPUT4), .B1(new_n236), .B2(new_n242), .ZN(new_n243));
  AND3_X1   g042(.A1(new_n235), .A2(KEYINPUT76), .A3(KEYINPUT4), .ZN(new_n244));
  AOI21_X1  g043(.A(KEYINPUT76), .B1(new_n235), .B2(KEYINPUT4), .ZN(new_n245));
  NOR3_X1   g044(.A1(new_n243), .A2(new_n244), .A3(new_n245), .ZN(new_n246));
  NAND2_X1  g045(.A1(G225gat), .A2(G233gat), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n215), .A2(new_n227), .ZN(new_n248));
  AOI22_X1  g047(.A1(new_n248), .A2(KEYINPUT3), .B1(new_n234), .B2(new_n222), .ZN(new_n249));
  INV_X1    g048(.A(KEYINPUT3), .ZN(new_n250));
  NAND3_X1  g049(.A1(new_n215), .A2(new_n250), .A3(new_n227), .ZN(new_n251));
  AOI21_X1  g050(.A(KEYINPUT75), .B1(new_n249), .B2(new_n251), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n224), .A2(new_n225), .ZN(new_n253));
  AND4_X1   g052(.A1(KEYINPUT74), .A2(new_n253), .A3(new_n213), .A4(new_n207), .ZN(new_n254));
  AOI21_X1  g053(.A(new_n213), .B1(new_n226), .B2(new_n207), .ZN(new_n255));
  OAI21_X1  g054(.A(KEYINPUT3), .B1(new_n254), .B2(new_n255), .ZN(new_n256));
  NAND2_X1  g055(.A1(new_n222), .A2(new_n234), .ZN(new_n257));
  NAND4_X1  g056(.A1(new_n256), .A2(KEYINPUT75), .A3(new_n251), .A4(new_n257), .ZN(new_n258));
  INV_X1    g057(.A(new_n258), .ZN(new_n259));
  OAI21_X1  g058(.A(new_n247), .B1(new_n252), .B2(new_n259), .ZN(new_n260));
  OAI21_X1  g059(.A(KEYINPUT78), .B1(new_n246), .B2(new_n260), .ZN(new_n261));
  NOR2_X1   g060(.A1(new_n244), .A2(new_n245), .ZN(new_n262));
  INV_X1    g061(.A(KEYINPUT4), .ZN(new_n263));
  NOR2_X1   g062(.A1(new_n254), .A2(new_n255), .ZN(new_n264));
  AOI21_X1  g063(.A(new_n241), .B1(new_n264), .B2(new_n240), .ZN(new_n265));
  NOR2_X1   g064(.A1(new_n235), .A2(KEYINPUT77), .ZN(new_n266));
  OAI21_X1  g065(.A(new_n263), .B1(new_n265), .B2(new_n266), .ZN(new_n267));
  NAND2_X1  g066(.A1(new_n262), .A2(new_n267), .ZN(new_n268));
  INV_X1    g067(.A(new_n247), .ZN(new_n269));
  NAND3_X1  g068(.A1(new_n256), .A2(new_n251), .A3(new_n257), .ZN(new_n270));
  INV_X1    g069(.A(KEYINPUT75), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  AOI21_X1  g071(.A(new_n269), .B1(new_n272), .B2(new_n258), .ZN(new_n273));
  INV_X1    g072(.A(KEYINPUT78), .ZN(new_n274));
  NAND3_X1  g073(.A1(new_n268), .A2(new_n273), .A3(new_n274), .ZN(new_n275));
  NAND2_X1  g074(.A1(new_n248), .A2(new_n257), .ZN(new_n276));
  NAND3_X1  g075(.A1(new_n236), .A2(new_n242), .A3(new_n276), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n277), .A2(new_n269), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n278), .A2(KEYINPUT5), .ZN(new_n279));
  INV_X1    g078(.A(KEYINPUT79), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  NAND3_X1  g080(.A1(new_n278), .A2(KEYINPUT79), .A3(KEYINPUT5), .ZN(new_n282));
  AOI22_X1  g081(.A1(new_n261), .A2(new_n275), .B1(new_n281), .B2(new_n282), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n235), .A2(new_n263), .ZN(new_n284));
  INV_X1    g083(.A(new_n284), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n236), .A2(new_n242), .ZN(new_n286));
  AOI21_X1  g085(.A(new_n285), .B1(new_n286), .B2(KEYINPUT4), .ZN(new_n287));
  INV_X1    g086(.A(KEYINPUT5), .ZN(new_n288));
  NAND2_X1  g087(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  NOR2_X1   g088(.A1(new_n289), .A2(new_n260), .ZN(new_n290));
  OAI21_X1  g089(.A(new_n205), .B1(new_n283), .B2(new_n290), .ZN(new_n291));
  AND3_X1   g090(.A1(new_n268), .A2(new_n274), .A3(new_n273), .ZN(new_n292));
  AOI21_X1  g091(.A(new_n274), .B1(new_n268), .B2(new_n273), .ZN(new_n293));
  AOI21_X1  g092(.A(KEYINPUT79), .B1(new_n278), .B2(KEYINPUT5), .ZN(new_n294));
  AOI211_X1 g093(.A(new_n280), .B(new_n288), .C1(new_n277), .C2(new_n269), .ZN(new_n295));
  OAI22_X1  g094(.A1(new_n292), .A2(new_n293), .B1(new_n294), .B2(new_n295), .ZN(new_n296));
  INV_X1    g095(.A(new_n205), .ZN(new_n297));
  OAI21_X1  g096(.A(new_n297), .B1(new_n289), .B2(new_n260), .ZN(new_n298));
  INV_X1    g097(.A(new_n298), .ZN(new_n299));
  AOI21_X1  g098(.A(KEYINPUT6), .B1(new_n296), .B2(new_n299), .ZN(new_n300));
  OAI21_X1  g099(.A(new_n291), .B1(new_n300), .B2(KEYINPUT80), .ZN(new_n301));
  INV_X1    g100(.A(KEYINPUT6), .ZN(new_n302));
  OAI211_X1 g101(.A(KEYINPUT80), .B(new_n302), .C1(new_n283), .C2(new_n298), .ZN(new_n303));
  INV_X1    g102(.A(new_n303), .ZN(new_n304));
  OAI21_X1  g103(.A(KEYINPUT81), .B1(new_n301), .B2(new_n304), .ZN(new_n305));
  OAI21_X1  g104(.A(new_n302), .B1(new_n283), .B2(new_n298), .ZN(new_n306));
  INV_X1    g105(.A(KEYINPUT80), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n306), .A2(new_n307), .ZN(new_n308));
  INV_X1    g107(.A(KEYINPUT81), .ZN(new_n309));
  NAND4_X1  g108(.A1(new_n308), .A2(new_n309), .A3(new_n303), .A4(new_n291), .ZN(new_n310));
  OAI211_X1 g109(.A(KEYINPUT6), .B(new_n205), .C1(new_n283), .C2(new_n290), .ZN(new_n311));
  NAND3_X1  g110(.A1(new_n305), .A2(new_n310), .A3(new_n311), .ZN(new_n312));
  XNOR2_X1  g111(.A(G197gat), .B(G204gat), .ZN(new_n313));
  INV_X1    g112(.A(G211gat), .ZN(new_n314));
  INV_X1    g113(.A(G218gat), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n315), .A2(KEYINPUT71), .ZN(new_n316));
  INV_X1    g115(.A(KEYINPUT71), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n317), .A2(G218gat), .ZN(new_n318));
  AOI21_X1  g117(.A(new_n314), .B1(new_n316), .B2(new_n318), .ZN(new_n319));
  XOR2_X1   g118(.A(KEYINPUT70), .B(KEYINPUT22), .Z(new_n320));
  OAI21_X1  g119(.A(new_n313), .B1(new_n319), .B2(new_n320), .ZN(new_n321));
  XNOR2_X1  g120(.A(G211gat), .B(G218gat), .ZN(new_n322));
  INV_X1    g121(.A(new_n322), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n321), .A2(new_n323), .ZN(new_n324));
  OAI211_X1 g123(.A(new_n322), .B(new_n313), .C1(new_n319), .C2(new_n320), .ZN(new_n325));
  NAND3_X1  g124(.A1(new_n324), .A2(KEYINPUT72), .A3(new_n325), .ZN(new_n326));
  XNOR2_X1  g125(.A(KEYINPUT70), .B(KEYINPUT22), .ZN(new_n327));
  XNOR2_X1  g126(.A(KEYINPUT71), .B(G218gat), .ZN(new_n328));
  OAI21_X1  g127(.A(new_n327), .B1(new_n328), .B2(new_n314), .ZN(new_n329));
  AOI21_X1  g128(.A(new_n322), .B1(new_n329), .B2(new_n313), .ZN(new_n330));
  INV_X1    g129(.A(KEYINPUT72), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n330), .A2(new_n331), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n326), .A2(new_n332), .ZN(new_n333));
  INV_X1    g132(.A(new_n333), .ZN(new_n334));
  NAND2_X1  g133(.A1(G226gat), .A2(G233gat), .ZN(new_n335));
  INV_X1    g134(.A(new_n335), .ZN(new_n336));
  INV_X1    g135(.A(G169gat), .ZN(new_n337));
  INV_X1    g136(.A(G176gat), .ZN(new_n338));
  NOR2_X1   g137(.A1(new_n337), .A2(new_n338), .ZN(new_n339));
  INV_X1    g138(.A(new_n339), .ZN(new_n340));
  INV_X1    g139(.A(KEYINPUT26), .ZN(new_n341));
  NOR2_X1   g140(.A1(G169gat), .A2(G176gat), .ZN(new_n342));
  AND3_X1   g141(.A1(new_n342), .A2(KEYINPUT65), .A3(new_n341), .ZN(new_n343));
  AOI21_X1  g142(.A(KEYINPUT65), .B1(new_n342), .B2(new_n341), .ZN(new_n344));
  OAI221_X1 g143(.A(new_n340), .B1(new_n341), .B2(new_n342), .C1(new_n343), .C2(new_n344), .ZN(new_n345));
  NAND2_X1  g144(.A1(G183gat), .A2(G190gat), .ZN(new_n346));
  XNOR2_X1  g145(.A(KEYINPUT27), .B(G183gat), .ZN(new_n347));
  XNOR2_X1  g146(.A(KEYINPUT64), .B(KEYINPUT28), .ZN(new_n348));
  INV_X1    g147(.A(G190gat), .ZN(new_n349));
  NAND3_X1  g148(.A1(new_n347), .A2(new_n348), .A3(new_n349), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n347), .A2(new_n349), .ZN(new_n351));
  INV_X1    g150(.A(KEYINPUT64), .ZN(new_n352));
  NAND3_X1  g151(.A1(new_n351), .A2(new_n352), .A3(KEYINPUT28), .ZN(new_n353));
  NAND4_X1  g152(.A1(new_n345), .A2(new_n346), .A3(new_n350), .A4(new_n353), .ZN(new_n354));
  INV_X1    g153(.A(KEYINPUT23), .ZN(new_n355));
  XNOR2_X1  g154(.A(new_n342), .B(new_n355), .ZN(new_n356));
  NOR2_X1   g155(.A1(new_n346), .A2(KEYINPUT24), .ZN(new_n357));
  NOR2_X1   g156(.A1(new_n357), .A2(new_n339), .ZN(new_n358));
  OR2_X1    g157(.A1(G183gat), .A2(G190gat), .ZN(new_n359));
  NAND3_X1  g158(.A1(new_n359), .A2(KEYINPUT24), .A3(new_n346), .ZN(new_n360));
  NAND3_X1  g159(.A1(new_n356), .A2(new_n358), .A3(new_n360), .ZN(new_n361));
  INV_X1    g160(.A(KEYINPUT25), .ZN(new_n362));
  AND2_X1   g161(.A1(new_n361), .A2(new_n362), .ZN(new_n363));
  NOR2_X1   g162(.A1(new_n361), .A2(new_n362), .ZN(new_n364));
  OAI21_X1  g163(.A(new_n354), .B1(new_n363), .B2(new_n364), .ZN(new_n365));
  INV_X1    g164(.A(KEYINPUT29), .ZN(new_n366));
  AOI21_X1  g165(.A(new_n336), .B1(new_n365), .B2(new_n366), .ZN(new_n367));
  XNOR2_X1  g166(.A(new_n361), .B(new_n362), .ZN(new_n368));
  AOI21_X1  g167(.A(new_n335), .B1(new_n368), .B2(new_n354), .ZN(new_n369));
  OAI21_X1  g168(.A(new_n334), .B1(new_n367), .B2(new_n369), .ZN(new_n370));
  XNOR2_X1  g169(.A(G8gat), .B(G36gat), .ZN(new_n371));
  XNOR2_X1  g170(.A(new_n371), .B(KEYINPUT73), .ZN(new_n372));
  XNOR2_X1  g171(.A(G64gat), .B(G92gat), .ZN(new_n373));
  XNOR2_X1  g172(.A(new_n372), .B(new_n373), .ZN(new_n374));
  NAND2_X1  g173(.A1(new_n365), .A2(new_n336), .ZN(new_n375));
  AOI21_X1  g174(.A(KEYINPUT29), .B1(new_n368), .B2(new_n354), .ZN(new_n376));
  OAI211_X1 g175(.A(new_n333), .B(new_n375), .C1(new_n376), .C2(new_n336), .ZN(new_n377));
  NAND3_X1  g176(.A1(new_n370), .A2(new_n374), .A3(new_n377), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n378), .A2(KEYINPUT30), .ZN(new_n379));
  AOI21_X1  g178(.A(new_n374), .B1(new_n370), .B2(new_n377), .ZN(new_n380));
  NOR2_X1   g179(.A1(new_n379), .A2(new_n380), .ZN(new_n381));
  AOI211_X1 g180(.A(KEYINPUT30), .B(new_n374), .C1(new_n370), .C2(new_n377), .ZN(new_n382));
  NOR2_X1   g181(.A1(new_n381), .A2(new_n382), .ZN(new_n383));
  INV_X1    g182(.A(new_n383), .ZN(new_n384));
  INV_X1    g183(.A(KEYINPUT83), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n251), .A2(new_n366), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n333), .A2(new_n386), .ZN(new_n387));
  NAND2_X1  g186(.A1(G228gat), .A2(G233gat), .ZN(new_n388));
  INV_X1    g187(.A(new_n388), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n387), .A2(new_n389), .ZN(new_n390));
  NAND3_X1  g189(.A1(new_n326), .A2(new_n366), .A3(new_n332), .ZN(new_n391));
  AOI21_X1  g190(.A(new_n264), .B1(new_n391), .B2(new_n250), .ZN(new_n392));
  NOR2_X1   g191(.A1(new_n390), .A2(new_n392), .ZN(new_n393));
  INV_X1    g192(.A(new_n325), .ZN(new_n394));
  OAI21_X1  g193(.A(new_n366), .B1(new_n394), .B2(new_n330), .ZN(new_n395));
  AOI21_X1  g194(.A(new_n264), .B1(new_n395), .B2(new_n250), .ZN(new_n396));
  AOI22_X1  g195(.A1(new_n326), .A2(new_n332), .B1(new_n366), .B2(new_n251), .ZN(new_n397));
  OAI21_X1  g196(.A(new_n388), .B1(new_n396), .B2(new_n397), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n398), .A2(KEYINPUT82), .ZN(new_n399));
  INV_X1    g198(.A(KEYINPUT82), .ZN(new_n400));
  OAI211_X1 g199(.A(new_n400), .B(new_n388), .C1(new_n396), .C2(new_n397), .ZN(new_n401));
  AOI21_X1  g200(.A(new_n393), .B1(new_n399), .B2(new_n401), .ZN(new_n402));
  INV_X1    g201(.A(G22gat), .ZN(new_n403));
  AOI21_X1  g202(.A(new_n385), .B1(new_n402), .B2(new_n403), .ZN(new_n404));
  XNOR2_X1  g203(.A(G78gat), .B(G106gat), .ZN(new_n405));
  XNOR2_X1  g204(.A(KEYINPUT31), .B(G50gat), .ZN(new_n406));
  XNOR2_X1  g205(.A(new_n405), .B(new_n406), .ZN(new_n407));
  INV_X1    g206(.A(new_n407), .ZN(new_n408));
  INV_X1    g207(.A(new_n390), .ZN(new_n409));
  INV_X1    g208(.A(new_n392), .ZN(new_n410));
  AOI221_X4 g209(.A(G22gat), .B1(new_n409), .B2(new_n410), .C1(new_n399), .C2(new_n401), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n399), .A2(new_n401), .ZN(new_n412));
  INV_X1    g211(.A(new_n393), .ZN(new_n413));
  AOI21_X1  g212(.A(new_n403), .B1(new_n412), .B2(new_n413), .ZN(new_n414));
  OAI22_X1  g213(.A1(new_n404), .A2(new_n408), .B1(new_n411), .B2(new_n414), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n412), .A2(new_n413), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n416), .A2(G22gat), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n402), .A2(new_n403), .ZN(new_n418));
  NAND4_X1  g217(.A1(new_n417), .A2(new_n385), .A3(new_n418), .A4(new_n407), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n415), .A2(new_n419), .ZN(new_n420));
  XNOR2_X1  g219(.A(G15gat), .B(G43gat), .ZN(new_n421));
  XNOR2_X1  g220(.A(G71gat), .B(G99gat), .ZN(new_n422));
  XNOR2_X1  g221(.A(new_n421), .B(new_n422), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n365), .A2(new_n240), .ZN(new_n424));
  INV_X1    g223(.A(G227gat), .ZN(new_n425));
  INV_X1    g224(.A(G233gat), .ZN(new_n426));
  NOR2_X1   g225(.A1(new_n425), .A2(new_n426), .ZN(new_n427));
  NAND3_X1  g226(.A1(new_n368), .A2(new_n257), .A3(new_n354), .ZN(new_n428));
  NAND3_X1  g227(.A1(new_n424), .A2(new_n427), .A3(new_n428), .ZN(new_n429));
  AOI21_X1  g228(.A(new_n423), .B1(new_n429), .B2(KEYINPUT32), .ZN(new_n430));
  INV_X1    g229(.A(KEYINPUT33), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n429), .A2(new_n431), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n430), .A2(new_n432), .ZN(new_n433));
  OR2_X1    g232(.A1(new_n423), .A2(KEYINPUT67), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n423), .A2(KEYINPUT67), .ZN(new_n435));
  NAND3_X1  g234(.A1(new_n434), .A2(KEYINPUT33), .A3(new_n435), .ZN(new_n436));
  NAND3_X1  g235(.A1(new_n429), .A2(KEYINPUT32), .A3(new_n436), .ZN(new_n437));
  INV_X1    g236(.A(KEYINPUT34), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n424), .A2(new_n428), .ZN(new_n439));
  INV_X1    g238(.A(new_n427), .ZN(new_n440));
  AOI21_X1  g239(.A(new_n438), .B1(new_n439), .B2(new_n440), .ZN(new_n441));
  AOI211_X1 g240(.A(KEYINPUT34), .B(new_n427), .C1(new_n424), .C2(new_n428), .ZN(new_n442));
  NOR2_X1   g241(.A1(new_n441), .A2(new_n442), .ZN(new_n443));
  OAI211_X1 g242(.A(new_n433), .B(new_n437), .C1(new_n443), .C2(KEYINPUT68), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n433), .A2(new_n437), .ZN(new_n445));
  INV_X1    g244(.A(KEYINPUT68), .ZN(new_n446));
  INV_X1    g245(.A(new_n443), .ZN(new_n447));
  NAND3_X1  g246(.A1(new_n445), .A2(new_n446), .A3(new_n447), .ZN(new_n448));
  AND3_X1   g247(.A1(new_n420), .A2(new_n444), .A3(new_n448), .ZN(new_n449));
  NAND3_X1  g248(.A1(new_n312), .A2(new_n384), .A3(new_n449), .ZN(new_n450));
  INV_X1    g249(.A(new_n290), .ZN(new_n451));
  AOI21_X1  g250(.A(new_n297), .B1(new_n296), .B2(new_n451), .ZN(new_n452));
  OAI21_X1  g251(.A(new_n311), .B1(new_n452), .B2(new_n306), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n453), .A2(new_n384), .ZN(new_n454));
  XNOR2_X1  g253(.A(new_n454), .B(KEYINPUT87), .ZN(new_n455));
  INV_X1    g254(.A(new_n420), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n445), .A2(new_n447), .ZN(new_n457));
  NAND3_X1  g256(.A1(new_n443), .A2(new_n433), .A3(new_n437), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  NOR3_X1   g258(.A1(new_n456), .A2(KEYINPUT35), .A3(new_n459), .ZN(new_n460));
  AOI22_X1  g259(.A1(new_n450), .A2(KEYINPUT35), .B1(new_n455), .B2(new_n460), .ZN(new_n461));
  INV_X1    g260(.A(KEYINPUT84), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n420), .A2(new_n462), .ZN(new_n463));
  NAND3_X1  g262(.A1(new_n415), .A2(KEYINPUT84), .A3(new_n419), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  AOI21_X1  g264(.A(new_n465), .B1(new_n312), .B2(new_n384), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n272), .A2(new_n258), .ZN(new_n467));
  AOI21_X1  g266(.A(new_n247), .B1(new_n287), .B2(new_n467), .ZN(new_n468));
  INV_X1    g267(.A(new_n468), .ZN(new_n469));
  INV_X1    g268(.A(KEYINPUT39), .ZN(new_n470));
  INV_X1    g269(.A(new_n277), .ZN(new_n471));
  AOI21_X1  g270(.A(new_n470), .B1(new_n471), .B2(new_n247), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n469), .A2(new_n472), .ZN(new_n473));
  AOI211_X1 g272(.A(KEYINPUT39), .B(new_n247), .C1(new_n287), .C2(new_n467), .ZN(new_n474));
  NOR3_X1   g273(.A1(new_n474), .A2(KEYINPUT85), .A3(new_n205), .ZN(new_n475));
  INV_X1    g274(.A(KEYINPUT85), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n468), .A2(new_n470), .ZN(new_n477));
  AOI21_X1  g276(.A(new_n476), .B1(new_n477), .B2(new_n297), .ZN(new_n478));
  OAI211_X1 g277(.A(KEYINPUT40), .B(new_n473), .C1(new_n475), .C2(new_n478), .ZN(new_n479));
  NAND3_X1  g278(.A1(new_n383), .A2(new_n479), .A3(new_n291), .ZN(new_n480));
  INV_X1    g279(.A(KEYINPUT86), .ZN(new_n481));
  OAI21_X1  g280(.A(KEYINPUT85), .B1(new_n474), .B2(new_n205), .ZN(new_n482));
  NAND3_X1  g281(.A1(new_n477), .A2(new_n476), .A3(new_n297), .ZN(new_n483));
  AOI22_X1  g282(.A1(new_n482), .A2(new_n483), .B1(new_n469), .B2(new_n472), .ZN(new_n484));
  OAI21_X1  g283(.A(new_n481), .B1(new_n484), .B2(KEYINPUT40), .ZN(new_n485));
  OAI21_X1  g284(.A(new_n473), .B1(new_n475), .B2(new_n478), .ZN(new_n486));
  INV_X1    g285(.A(KEYINPUT40), .ZN(new_n487));
  NAND3_X1  g286(.A1(new_n486), .A2(KEYINPUT86), .A3(new_n487), .ZN(new_n488));
  AOI21_X1  g287(.A(new_n480), .B1(new_n485), .B2(new_n488), .ZN(new_n489));
  INV_X1    g288(.A(KEYINPUT37), .ZN(new_n490));
  AND3_X1   g289(.A1(new_n370), .A2(new_n490), .A3(new_n377), .ZN(new_n491));
  AOI21_X1  g290(.A(new_n490), .B1(new_n370), .B2(new_n377), .ZN(new_n492));
  OAI21_X1  g291(.A(new_n374), .B1(new_n491), .B2(new_n492), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n493), .A2(KEYINPUT38), .ZN(new_n494));
  INV_X1    g293(.A(new_n380), .ZN(new_n495));
  INV_X1    g294(.A(KEYINPUT38), .ZN(new_n496));
  OAI211_X1 g295(.A(new_n496), .B(new_n374), .C1(new_n491), .C2(new_n492), .ZN(new_n497));
  NAND3_X1  g296(.A1(new_n494), .A2(new_n495), .A3(new_n497), .ZN(new_n498));
  OAI21_X1  g297(.A(new_n420), .B1(new_n453), .B2(new_n498), .ZN(new_n499));
  INV_X1    g298(.A(KEYINPUT69), .ZN(new_n500));
  INV_X1    g299(.A(KEYINPUT36), .ZN(new_n501));
  AOI21_X1  g300(.A(new_n500), .B1(new_n459), .B2(new_n501), .ZN(new_n502));
  AND3_X1   g301(.A1(new_n443), .A2(new_n433), .A3(new_n437), .ZN(new_n503));
  AOI21_X1  g302(.A(new_n443), .B1(new_n433), .B2(new_n437), .ZN(new_n504));
  OAI211_X1 g303(.A(new_n500), .B(new_n501), .C1(new_n503), .C2(new_n504), .ZN(new_n505));
  NAND3_X1  g304(.A1(new_n448), .A2(KEYINPUT36), .A3(new_n444), .ZN(new_n506));
  NAND2_X1  g305(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  OAI22_X1  g306(.A1(new_n489), .A2(new_n499), .B1(new_n502), .B2(new_n507), .ZN(new_n508));
  NOR2_X1   g307(.A1(new_n466), .A2(new_n508), .ZN(new_n509));
  OAI21_X1  g308(.A(KEYINPUT88), .B1(new_n461), .B2(new_n509), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n450), .A2(KEYINPUT35), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n455), .A2(new_n460), .ZN(new_n512));
  NAND2_X1  g311(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  INV_X1    g312(.A(KEYINPUT88), .ZN(new_n514));
  NOR2_X1   g313(.A1(new_n507), .A2(new_n502), .ZN(new_n515));
  INV_X1    g314(.A(new_n499), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n485), .A2(new_n488), .ZN(new_n517));
  AND3_X1   g316(.A1(new_n383), .A2(new_n479), .A3(new_n291), .ZN(new_n518));
  NAND2_X1  g317(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  AOI21_X1  g318(.A(new_n515), .B1(new_n516), .B2(new_n519), .ZN(new_n520));
  NAND3_X1  g319(.A1(new_n308), .A2(new_n303), .A3(new_n291), .ZN(new_n521));
  AOI22_X1  g320(.A1(new_n521), .A2(KEYINPUT81), .B1(KEYINPUT6), .B2(new_n452), .ZN(new_n522));
  AOI21_X1  g321(.A(new_n383), .B1(new_n522), .B2(new_n310), .ZN(new_n523));
  OAI21_X1  g322(.A(new_n520), .B1(new_n523), .B2(new_n465), .ZN(new_n524));
  NAND3_X1  g323(.A1(new_n513), .A2(new_n514), .A3(new_n524), .ZN(new_n525));
  AND2_X1   g324(.A1(new_n510), .A2(new_n525), .ZN(new_n526));
  INV_X1    g325(.A(G36gat), .ZN(new_n527));
  AND2_X1   g326(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n528));
  NOR2_X1   g327(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n529));
  OAI21_X1  g328(.A(new_n527), .B1(new_n528), .B2(new_n529), .ZN(new_n530));
  INV_X1    g329(.A(G29gat), .ZN(new_n531));
  NAND3_X1  g330(.A1(new_n531), .A2(KEYINPUT14), .A3(G36gat), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n530), .A2(new_n532), .ZN(new_n533));
  OR2_X1    g332(.A1(new_n533), .A2(KEYINPUT15), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n533), .A2(KEYINPUT15), .ZN(new_n535));
  XNOR2_X1  g334(.A(G43gat), .B(G50gat), .ZN(new_n536));
  NAND3_X1  g335(.A1(new_n534), .A2(new_n535), .A3(new_n536), .ZN(new_n537));
  OR2_X1    g336(.A1(new_n535), .A2(new_n536), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  XNOR2_X1  g338(.A(new_n539), .B(KEYINPUT17), .ZN(new_n540));
  INV_X1    g339(.A(G99gat), .ZN(new_n541));
  INV_X1    g340(.A(G106gat), .ZN(new_n542));
  OAI21_X1  g341(.A(KEYINPUT8), .B1(new_n541), .B2(new_n542), .ZN(new_n543));
  OAI21_X1  g342(.A(new_n543), .B1(G85gat), .B2(G92gat), .ZN(new_n544));
  XOR2_X1   g343(.A(G99gat), .B(G106gat), .Z(new_n545));
  AOI21_X1  g344(.A(new_n544), .B1(KEYINPUT97), .B2(new_n545), .ZN(new_n546));
  OR2_X1    g345(.A1(new_n545), .A2(KEYINPUT97), .ZN(new_n547));
  NAND2_X1  g346(.A1(G85gat), .A2(G92gat), .ZN(new_n548));
  INV_X1    g347(.A(KEYINPUT96), .ZN(new_n549));
  OR3_X1    g348(.A1(new_n548), .A2(new_n549), .A3(KEYINPUT7), .ZN(new_n550));
  OAI21_X1  g349(.A(new_n549), .B1(new_n548), .B2(KEYINPUT7), .ZN(new_n551));
  AOI21_X1  g350(.A(KEYINPUT95), .B1(new_n548), .B2(KEYINPUT7), .ZN(new_n552));
  AND3_X1   g351(.A1(new_n548), .A2(KEYINPUT95), .A3(KEYINPUT7), .ZN(new_n553));
  OAI211_X1 g352(.A(new_n550), .B(new_n551), .C1(new_n552), .C2(new_n553), .ZN(new_n554));
  AND3_X1   g353(.A1(new_n546), .A2(new_n547), .A3(new_n554), .ZN(new_n555));
  AOI21_X1  g354(.A(new_n547), .B1(new_n546), .B2(new_n554), .ZN(new_n556));
  NOR2_X1   g355(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n557), .A2(KEYINPUT98), .ZN(new_n558));
  INV_X1    g357(.A(KEYINPUT98), .ZN(new_n559));
  OAI21_X1  g358(.A(new_n559), .B1(new_n555), .B2(new_n556), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n558), .A2(new_n560), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n540), .A2(new_n561), .ZN(new_n562));
  NAND3_X1  g361(.A1(new_n558), .A2(new_n539), .A3(new_n560), .ZN(new_n563));
  NAND3_X1  g362(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n564));
  NAND3_X1  g363(.A1(new_n562), .A2(new_n563), .A3(new_n564), .ZN(new_n565));
  XOR2_X1   g364(.A(G190gat), .B(G218gat), .Z(new_n566));
  OR2_X1    g365(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n565), .A2(new_n566), .ZN(new_n568));
  NAND2_X1  g367(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  AOI21_X1  g368(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n570));
  XNOR2_X1  g369(.A(new_n570), .B(KEYINPUT94), .ZN(new_n571));
  XNOR2_X1  g370(.A(G134gat), .B(G162gat), .ZN(new_n572));
  XNOR2_X1  g371(.A(new_n571), .B(new_n572), .ZN(new_n573));
  INV_X1    g372(.A(new_n573), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n569), .A2(new_n574), .ZN(new_n575));
  NAND3_X1  g374(.A1(new_n567), .A2(new_n573), .A3(new_n568), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  INV_X1    g376(.A(new_n577), .ZN(new_n578));
  XOR2_X1   g377(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n579));
  XNOR2_X1  g378(.A(new_n579), .B(G155gat), .ZN(new_n580));
  XNOR2_X1  g379(.A(G183gat), .B(G211gat), .ZN(new_n581));
  XOR2_X1   g380(.A(new_n580), .B(new_n581), .Z(new_n582));
  INV_X1    g381(.A(new_n582), .ZN(new_n583));
  XOR2_X1   g382(.A(G57gat), .B(G64gat), .Z(new_n584));
  INV_X1    g383(.A(KEYINPUT93), .ZN(new_n585));
  INV_X1    g384(.A(KEYINPUT9), .ZN(new_n586));
  INV_X1    g385(.A(G71gat), .ZN(new_n587));
  INV_X1    g386(.A(G78gat), .ZN(new_n588));
  OAI21_X1  g387(.A(new_n586), .B1(new_n587), .B2(new_n588), .ZN(new_n589));
  OAI21_X1  g388(.A(new_n584), .B1(new_n585), .B2(new_n589), .ZN(new_n590));
  XOR2_X1   g389(.A(G71gat), .B(G78gat), .Z(new_n591));
  AND2_X1   g390(.A1(new_n589), .A2(new_n585), .ZN(new_n592));
  OR3_X1    g391(.A1(new_n590), .A2(new_n591), .A3(new_n592), .ZN(new_n593));
  OAI21_X1  g392(.A(new_n591), .B1(new_n590), .B2(new_n592), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  INV_X1    g394(.A(KEYINPUT21), .ZN(new_n596));
  NAND2_X1  g395(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  INV_X1    g396(.A(G231gat), .ZN(new_n598));
  NOR2_X1   g397(.A1(new_n598), .A2(new_n426), .ZN(new_n599));
  AND2_X1   g398(.A1(new_n597), .A2(new_n599), .ZN(new_n600));
  NOR2_X1   g399(.A1(new_n597), .A2(new_n599), .ZN(new_n601));
  NOR3_X1   g400(.A1(new_n600), .A2(new_n601), .A3(G127gat), .ZN(new_n602));
  INV_X1    g401(.A(new_n602), .ZN(new_n603));
  XNOR2_X1  g402(.A(G15gat), .B(G22gat), .ZN(new_n604));
  OR2_X1    g403(.A1(new_n604), .A2(G1gat), .ZN(new_n605));
  INV_X1    g404(.A(KEYINPUT16), .ZN(new_n606));
  OAI21_X1  g405(.A(new_n604), .B1(new_n606), .B2(G1gat), .ZN(new_n607));
  INV_X1    g406(.A(G8gat), .ZN(new_n608));
  NAND3_X1  g407(.A1(new_n605), .A2(new_n607), .A3(new_n608), .ZN(new_n609));
  XNOR2_X1  g408(.A(new_n609), .B(KEYINPUT91), .ZN(new_n610));
  NAND3_X1  g409(.A1(new_n605), .A2(new_n607), .A3(KEYINPUT90), .ZN(new_n611));
  OAI211_X1 g410(.A(new_n611), .B(G8gat), .C1(KEYINPUT90), .C2(new_n605), .ZN(new_n612));
  NAND2_X1  g411(.A1(new_n610), .A2(new_n612), .ZN(new_n613));
  INV_X1    g412(.A(new_n613), .ZN(new_n614));
  OAI21_X1  g413(.A(new_n614), .B1(new_n596), .B2(new_n595), .ZN(new_n615));
  OAI21_X1  g414(.A(G127gat), .B1(new_n600), .B2(new_n601), .ZN(new_n616));
  NAND3_X1  g415(.A1(new_n603), .A2(new_n615), .A3(new_n616), .ZN(new_n617));
  INV_X1    g416(.A(new_n617), .ZN(new_n618));
  AOI21_X1  g417(.A(new_n615), .B1(new_n603), .B2(new_n616), .ZN(new_n619));
  OAI21_X1  g418(.A(new_n583), .B1(new_n618), .B2(new_n619), .ZN(new_n620));
  INV_X1    g419(.A(new_n619), .ZN(new_n621));
  NAND3_X1  g420(.A1(new_n621), .A2(new_n617), .A3(new_n582), .ZN(new_n622));
  NAND2_X1  g421(.A1(new_n620), .A2(new_n622), .ZN(new_n623));
  INV_X1    g422(.A(G230gat), .ZN(new_n624));
  NOR2_X1   g423(.A1(new_n624), .A2(new_n426), .ZN(new_n625));
  INV_X1    g424(.A(KEYINPUT10), .ZN(new_n626));
  INV_X1    g425(.A(new_n595), .ZN(new_n627));
  NOR2_X1   g426(.A1(new_n557), .A2(new_n627), .ZN(new_n628));
  NOR3_X1   g427(.A1(new_n595), .A2(new_n555), .A3(new_n556), .ZN(new_n629));
  OAI21_X1  g428(.A(new_n626), .B1(new_n628), .B2(new_n629), .ZN(new_n630));
  NAND4_X1  g429(.A1(new_n558), .A2(KEYINPUT10), .A3(new_n627), .A4(new_n560), .ZN(new_n631));
  AOI21_X1  g430(.A(new_n625), .B1(new_n630), .B2(new_n631), .ZN(new_n632));
  NOR2_X1   g431(.A1(new_n628), .A2(new_n629), .ZN(new_n633));
  AOI21_X1  g432(.A(new_n632), .B1(new_n625), .B2(new_n633), .ZN(new_n634));
  XOR2_X1   g433(.A(G120gat), .B(G148gat), .Z(new_n635));
  XNOR2_X1  g434(.A(new_n635), .B(KEYINPUT99), .ZN(new_n636));
  XNOR2_X1  g435(.A(G176gat), .B(G204gat), .ZN(new_n637));
  XOR2_X1   g436(.A(new_n636), .B(new_n637), .Z(new_n638));
  OR2_X1    g437(.A1(new_n634), .A2(new_n638), .ZN(new_n639));
  INV_X1    g438(.A(new_n632), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n633), .A2(new_n625), .ZN(new_n641));
  NAND3_X1  g440(.A1(new_n640), .A2(new_n641), .A3(new_n638), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n639), .A2(new_n642), .ZN(new_n643));
  INV_X1    g442(.A(new_n643), .ZN(new_n644));
  NAND3_X1  g443(.A1(new_n578), .A2(new_n623), .A3(new_n644), .ZN(new_n645));
  XOR2_X1   g444(.A(G113gat), .B(G141gat), .Z(new_n646));
  XNOR2_X1  g445(.A(KEYINPUT89), .B(G197gat), .ZN(new_n647));
  XNOR2_X1  g446(.A(new_n646), .B(new_n647), .ZN(new_n648));
  XOR2_X1   g447(.A(KEYINPUT11), .B(G169gat), .Z(new_n649));
  XNOR2_X1  g448(.A(new_n648), .B(new_n649), .ZN(new_n650));
  XOR2_X1   g449(.A(new_n650), .B(KEYINPUT12), .Z(new_n651));
  INV_X1    g450(.A(new_n651), .ZN(new_n652));
  NAND2_X1  g451(.A1(G229gat), .A2(G233gat), .ZN(new_n653));
  INV_X1    g452(.A(new_n653), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n613), .A2(new_n539), .ZN(new_n655));
  NOR2_X1   g454(.A1(new_n539), .A2(KEYINPUT17), .ZN(new_n656));
  INV_X1    g455(.A(KEYINPUT17), .ZN(new_n657));
  AOI21_X1  g456(.A(new_n657), .B1(new_n537), .B2(new_n538), .ZN(new_n658));
  NOR2_X1   g457(.A1(new_n656), .A2(new_n658), .ZN(new_n659));
  OAI211_X1 g458(.A(KEYINPUT92), .B(new_n655), .C1(new_n659), .C2(new_n613), .ZN(new_n660));
  INV_X1    g459(.A(KEYINPUT92), .ZN(new_n661));
  NAND3_X1  g460(.A1(new_n540), .A2(new_n661), .A3(new_n614), .ZN(new_n662));
  AOI21_X1  g461(.A(new_n654), .B1(new_n660), .B2(new_n662), .ZN(new_n663));
  OR2_X1    g462(.A1(new_n613), .A2(new_n539), .ZN(new_n664));
  AND2_X1   g463(.A1(new_n664), .A2(new_n655), .ZN(new_n665));
  XOR2_X1   g464(.A(new_n653), .B(KEYINPUT13), .Z(new_n666));
  INV_X1    g465(.A(new_n666), .ZN(new_n667));
  OAI22_X1  g466(.A1(new_n663), .A2(KEYINPUT18), .B1(new_n665), .B2(new_n667), .ZN(new_n668));
  AND2_X1   g467(.A1(new_n663), .A2(KEYINPUT18), .ZN(new_n669));
  OAI21_X1  g468(.A(new_n652), .B1(new_n668), .B2(new_n669), .ZN(new_n670));
  NOR2_X1   g469(.A1(new_n665), .A2(new_n667), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n660), .A2(new_n662), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n672), .A2(new_n653), .ZN(new_n673));
  INV_X1    g472(.A(KEYINPUT18), .ZN(new_n674));
  AOI21_X1  g473(.A(new_n671), .B1(new_n673), .B2(new_n674), .ZN(new_n675));
  NAND2_X1  g474(.A1(new_n663), .A2(KEYINPUT18), .ZN(new_n676));
  NAND3_X1  g475(.A1(new_n675), .A2(new_n676), .A3(new_n651), .ZN(new_n677));
  NAND2_X1  g476(.A1(new_n670), .A2(new_n677), .ZN(new_n678));
  INV_X1    g477(.A(new_n678), .ZN(new_n679));
  NOR2_X1   g478(.A1(new_n645), .A2(new_n679), .ZN(new_n680));
  NAND2_X1  g479(.A1(new_n526), .A2(new_n680), .ZN(new_n681));
  INV_X1    g480(.A(new_n681), .ZN(new_n682));
  INV_X1    g481(.A(new_n312), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  XNOR2_X1  g483(.A(new_n684), .B(G1gat), .ZN(G1324gat));
  OAI21_X1  g484(.A(G8gat), .B1(new_n681), .B2(new_n384), .ZN(new_n686));
  INV_X1    g485(.A(KEYINPUT42), .ZN(new_n687));
  XOR2_X1   g486(.A(KEYINPUT16), .B(G8gat), .Z(new_n688));
  NAND3_X1  g487(.A1(new_n682), .A2(new_n383), .A3(new_n688), .ZN(new_n689));
  INV_X1    g488(.A(KEYINPUT101), .ZN(new_n690));
  XOR2_X1   g489(.A(KEYINPUT100), .B(KEYINPUT42), .Z(new_n691));
  NAND3_X1  g490(.A1(new_n689), .A2(new_n690), .A3(new_n691), .ZN(new_n692));
  INV_X1    g491(.A(new_n692), .ZN(new_n693));
  AOI21_X1  g492(.A(new_n690), .B1(new_n689), .B2(new_n691), .ZN(new_n694));
  OAI221_X1 g493(.A(new_n686), .B1(new_n687), .B2(new_n689), .C1(new_n693), .C2(new_n694), .ZN(G1325gat));
  INV_X1    g494(.A(new_n459), .ZN(new_n696));
  AOI21_X1  g495(.A(G15gat), .B1(new_n682), .B2(new_n696), .ZN(new_n697));
  OR2_X1    g496(.A1(new_n515), .A2(KEYINPUT102), .ZN(new_n698));
  NAND2_X1  g497(.A1(new_n515), .A2(KEYINPUT102), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  INV_X1    g499(.A(new_n700), .ZN(new_n701));
  NAND2_X1  g500(.A1(new_n701), .A2(G15gat), .ZN(new_n702));
  XNOR2_X1  g501(.A(new_n702), .B(KEYINPUT103), .ZN(new_n703));
  AOI21_X1  g502(.A(new_n697), .B1(new_n682), .B2(new_n703), .ZN(G1326gat));
  NOR2_X1   g503(.A1(new_n681), .A2(new_n465), .ZN(new_n705));
  XOR2_X1   g504(.A(KEYINPUT43), .B(G22gat), .Z(new_n706));
  XNOR2_X1  g505(.A(new_n705), .B(new_n706), .ZN(G1327gat));
  NAND3_X1  g506(.A1(new_n510), .A2(new_n525), .A3(new_n577), .ZN(new_n708));
  INV_X1    g507(.A(new_n708), .ZN(new_n709));
  NOR3_X1   g508(.A1(new_n679), .A2(new_n623), .A3(new_n643), .ZN(new_n710));
  NAND2_X1  g509(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  NOR3_X1   g510(.A1(new_n711), .A2(G29gat), .A3(new_n312), .ZN(new_n712));
  XOR2_X1   g511(.A(new_n712), .B(KEYINPUT45), .Z(new_n713));
  XOR2_X1   g512(.A(new_n710), .B(KEYINPUT104), .Z(new_n714));
  OAI21_X1  g513(.A(KEYINPUT105), .B1(new_n466), .B2(new_n508), .ZN(new_n715));
  INV_X1    g514(.A(KEYINPUT105), .ZN(new_n716));
  OAI211_X1 g515(.A(new_n520), .B(new_n716), .C1(new_n523), .C2(new_n465), .ZN(new_n717));
  NAND2_X1  g516(.A1(new_n715), .A2(new_n717), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n718), .A2(new_n513), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n719), .A2(KEYINPUT106), .ZN(new_n720));
  AOI21_X1  g519(.A(new_n461), .B1(new_n715), .B2(new_n717), .ZN(new_n721));
  INV_X1    g520(.A(KEYINPUT106), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  NOR2_X1   g522(.A1(new_n578), .A2(KEYINPUT44), .ZN(new_n724));
  NAND3_X1  g523(.A1(new_n720), .A2(new_n723), .A3(new_n724), .ZN(new_n725));
  NAND2_X1  g524(.A1(new_n708), .A2(KEYINPUT44), .ZN(new_n726));
  AOI21_X1  g525(.A(new_n714), .B1(new_n725), .B2(new_n726), .ZN(new_n727));
  AND2_X1   g526(.A1(new_n727), .A2(new_n683), .ZN(new_n728));
  OAI21_X1  g527(.A(new_n713), .B1(new_n728), .B2(new_n531), .ZN(G1328gat));
  NAND4_X1  g528(.A1(new_n709), .A2(new_n527), .A3(new_n383), .A4(new_n710), .ZN(new_n730));
  XNOR2_X1  g529(.A(new_n730), .B(KEYINPUT46), .ZN(new_n731));
  AOI21_X1  g530(.A(new_n527), .B1(new_n727), .B2(new_n383), .ZN(new_n732));
  INV_X1    g531(.A(KEYINPUT107), .ZN(new_n733));
  OR3_X1    g532(.A1(new_n731), .A2(new_n732), .A3(new_n733), .ZN(new_n734));
  OAI21_X1  g533(.A(new_n733), .B1(new_n731), .B2(new_n732), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n734), .A2(new_n735), .ZN(G1329gat));
  NOR3_X1   g535(.A1(new_n711), .A2(G43gat), .A3(new_n459), .ZN(new_n737));
  NAND2_X1  g536(.A1(new_n727), .A2(new_n701), .ZN(new_n738));
  AOI21_X1  g537(.A(new_n737), .B1(new_n738), .B2(G43gat), .ZN(new_n739));
  INV_X1    g538(.A(KEYINPUT47), .ZN(new_n740));
  OR2_X1    g539(.A1(new_n737), .A2(new_n740), .ZN(new_n741));
  INV_X1    g540(.A(G43gat), .ZN(new_n742));
  AOI21_X1  g541(.A(new_n742), .B1(new_n727), .B2(new_n515), .ZN(new_n743));
  OAI22_X1  g542(.A1(new_n739), .A2(KEYINPUT47), .B1(new_n741), .B2(new_n743), .ZN(G1330gat));
  NOR3_X1   g543(.A1(new_n711), .A2(G50gat), .A3(new_n465), .ZN(new_n745));
  INV_X1    g544(.A(new_n465), .ZN(new_n746));
  NAND2_X1  g545(.A1(new_n727), .A2(new_n746), .ZN(new_n747));
  AOI21_X1  g546(.A(new_n745), .B1(new_n747), .B2(G50gat), .ZN(new_n748));
  INV_X1    g547(.A(KEYINPUT48), .ZN(new_n749));
  OR2_X1    g548(.A1(new_n745), .A2(new_n749), .ZN(new_n750));
  INV_X1    g549(.A(G50gat), .ZN(new_n751));
  AOI21_X1  g550(.A(new_n751), .B1(new_n727), .B2(new_n456), .ZN(new_n752));
  OAI22_X1  g551(.A1(new_n748), .A2(KEYINPUT48), .B1(new_n750), .B2(new_n752), .ZN(G1331gat));
  AND2_X1   g552(.A1(new_n720), .A2(new_n723), .ZN(new_n754));
  NAND3_X1  g553(.A1(new_n623), .A2(new_n576), .A3(new_n575), .ZN(new_n755));
  NOR3_X1   g554(.A1(new_n755), .A2(new_n644), .A3(new_n678), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n754), .A2(new_n756), .ZN(new_n757));
  NOR2_X1   g556(.A1(new_n757), .A2(new_n312), .ZN(new_n758));
  XOR2_X1   g557(.A(KEYINPUT108), .B(G57gat), .Z(new_n759));
  XNOR2_X1  g558(.A(new_n758), .B(new_n759), .ZN(G1332gat));
  AND2_X1   g559(.A1(new_n754), .A2(new_n756), .ZN(new_n761));
  AOI21_X1  g560(.A(new_n384), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  NAND2_X1  g562(.A1(new_n763), .A2(KEYINPUT109), .ZN(new_n764));
  NOR2_X1   g563(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n765));
  INV_X1    g564(.A(KEYINPUT109), .ZN(new_n766));
  NAND3_X1  g565(.A1(new_n761), .A2(new_n766), .A3(new_n762), .ZN(new_n767));
  AND3_X1   g566(.A1(new_n764), .A2(new_n765), .A3(new_n767), .ZN(new_n768));
  AOI21_X1  g567(.A(new_n765), .B1(new_n764), .B2(new_n767), .ZN(new_n769));
  NOR2_X1   g568(.A1(new_n768), .A2(new_n769), .ZN(G1333gat));
  NAND3_X1  g569(.A1(new_n761), .A2(new_n587), .A3(new_n696), .ZN(new_n771));
  OAI21_X1  g570(.A(G71gat), .B1(new_n757), .B2(new_n700), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  INV_X1    g572(.A(KEYINPUT50), .ZN(new_n774));
  XNOR2_X1  g573(.A(new_n773), .B(new_n774), .ZN(G1334gat));
  NOR2_X1   g574(.A1(new_n757), .A2(new_n465), .ZN(new_n776));
  XNOR2_X1  g575(.A(KEYINPUT110), .B(G78gat), .ZN(new_n777));
  XNOR2_X1  g576(.A(new_n776), .B(new_n777), .ZN(G1335gat));
  NAND2_X1  g577(.A1(new_n725), .A2(new_n726), .ZN(new_n779));
  NOR2_X1   g578(.A1(new_n644), .A2(new_n678), .ZN(new_n780));
  INV_X1    g579(.A(new_n623), .ZN(new_n781));
  NAND2_X1  g580(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  INV_X1    g581(.A(new_n782), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n779), .A2(new_n783), .ZN(new_n784));
  OAI21_X1  g583(.A(G85gat), .B1(new_n784), .B2(new_n312), .ZN(new_n785));
  INV_X1    g584(.A(KEYINPUT51), .ZN(new_n786));
  NOR2_X1   g585(.A1(new_n678), .A2(new_n623), .ZN(new_n787));
  AOI21_X1  g586(.A(new_n578), .B1(new_n718), .B2(new_n513), .ZN(new_n788));
  INV_X1    g587(.A(KEYINPUT111), .ZN(new_n789));
  OAI21_X1  g588(.A(new_n787), .B1(new_n788), .B2(new_n789), .ZN(new_n790));
  NOR3_X1   g589(.A1(new_n721), .A2(KEYINPUT111), .A3(new_n578), .ZN(new_n791));
  OAI21_X1  g590(.A(new_n786), .B1(new_n790), .B2(new_n791), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n788), .A2(new_n789), .ZN(new_n793));
  OAI21_X1  g592(.A(KEYINPUT111), .B1(new_n721), .B2(new_n578), .ZN(new_n794));
  NAND4_X1  g593(.A1(new_n793), .A2(new_n794), .A3(KEYINPUT51), .A4(new_n787), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n792), .A2(new_n795), .ZN(new_n796));
  INV_X1    g595(.A(new_n796), .ZN(new_n797));
  OR3_X1    g596(.A1(new_n312), .A2(G85gat), .A3(new_n644), .ZN(new_n798));
  OAI21_X1  g597(.A(new_n785), .B1(new_n797), .B2(new_n798), .ZN(G1336gat));
  INV_X1    g598(.A(G92gat), .ZN(new_n800));
  AOI21_X1  g599(.A(new_n782), .B1(new_n725), .B2(new_n726), .ZN(new_n801));
  AOI21_X1  g600(.A(new_n800), .B1(new_n801), .B2(new_n383), .ZN(new_n802));
  NOR3_X1   g601(.A1(new_n644), .A2(G92gat), .A3(new_n384), .ZN(new_n803));
  AOI21_X1  g602(.A(new_n802), .B1(new_n796), .B2(new_n803), .ZN(new_n804));
  INV_X1    g603(.A(KEYINPUT52), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  AND2_X1   g605(.A1(new_n796), .A2(new_n803), .ZN(new_n807));
  OAI21_X1  g606(.A(KEYINPUT52), .B1(new_n807), .B2(new_n802), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n806), .A2(new_n808), .ZN(G1337gat));
  OAI21_X1  g608(.A(G99gat), .B1(new_n784), .B2(new_n700), .ZN(new_n810));
  NAND3_X1  g609(.A1(new_n643), .A2(new_n696), .A3(new_n541), .ZN(new_n811));
  OAI21_X1  g610(.A(new_n810), .B1(new_n797), .B2(new_n811), .ZN(G1338gat));
  AOI21_X1  g611(.A(new_n542), .B1(new_n801), .B2(new_n746), .ZN(new_n813));
  NOR3_X1   g612(.A1(new_n644), .A2(G106gat), .A3(new_n420), .ZN(new_n814));
  INV_X1    g613(.A(new_n814), .ZN(new_n815));
  AOI21_X1  g614(.A(new_n815), .B1(new_n792), .B2(new_n795), .ZN(new_n816));
  OAI21_X1  g615(.A(KEYINPUT53), .B1(new_n813), .B2(new_n816), .ZN(new_n817));
  AOI21_X1  g616(.A(new_n542), .B1(new_n801), .B2(new_n456), .ZN(new_n818));
  NOR4_X1   g617(.A1(new_n818), .A2(new_n816), .A3(KEYINPUT112), .A4(KEYINPUT53), .ZN(new_n819));
  INV_X1    g618(.A(KEYINPUT112), .ZN(new_n820));
  AOI21_X1  g619(.A(KEYINPUT53), .B1(new_n796), .B2(new_n814), .ZN(new_n821));
  OAI21_X1  g620(.A(G106gat), .B1(new_n784), .B2(new_n420), .ZN(new_n822));
  AOI21_X1  g621(.A(new_n820), .B1(new_n821), .B2(new_n822), .ZN(new_n823));
  OAI21_X1  g622(.A(new_n817), .B1(new_n819), .B2(new_n823), .ZN(G1339gat));
  INV_X1    g623(.A(KEYINPUT115), .ZN(new_n825));
  NAND3_X1  g624(.A1(new_n630), .A2(new_n625), .A3(new_n631), .ZN(new_n826));
  NAND3_X1  g625(.A1(new_n640), .A2(new_n826), .A3(KEYINPUT54), .ZN(new_n827));
  XOR2_X1   g626(.A(KEYINPUT114), .B(KEYINPUT54), .Z(new_n828));
  AOI21_X1  g627(.A(new_n638), .B1(new_n632), .B2(new_n828), .ZN(new_n829));
  NAND3_X1  g628(.A1(new_n827), .A2(KEYINPUT55), .A3(new_n829), .ZN(new_n830));
  AND2_X1   g629(.A1(new_n830), .A2(new_n642), .ZN(new_n831));
  NAND2_X1  g630(.A1(new_n827), .A2(new_n829), .ZN(new_n832));
  INV_X1    g631(.A(KEYINPUT55), .ZN(new_n833));
  NAND2_X1  g632(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  NAND3_X1  g633(.A1(new_n678), .A2(new_n831), .A3(new_n834), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n665), .A2(new_n667), .ZN(new_n836));
  NAND3_X1  g635(.A1(new_n660), .A2(new_n662), .A3(new_n654), .ZN(new_n837));
  AND2_X1   g636(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  NOR2_X1   g637(.A1(new_n838), .A2(new_n650), .ZN(new_n839));
  NOR2_X1   g638(.A1(new_n668), .A2(new_n669), .ZN(new_n840));
  AOI21_X1  g639(.A(new_n839), .B1(new_n840), .B2(new_n651), .ZN(new_n841));
  NAND2_X1  g640(.A1(new_n841), .A2(new_n643), .ZN(new_n842));
  AOI21_X1  g641(.A(new_n577), .B1(new_n835), .B2(new_n842), .ZN(new_n843));
  AND3_X1   g642(.A1(new_n834), .A2(new_n642), .A3(new_n830), .ZN(new_n844));
  AND3_X1   g643(.A1(new_n844), .A2(new_n577), .A3(new_n841), .ZN(new_n845));
  OAI21_X1  g644(.A(new_n825), .B1(new_n843), .B2(new_n845), .ZN(new_n846));
  NAND3_X1  g645(.A1(new_n844), .A2(new_n577), .A3(new_n841), .ZN(new_n847));
  AOI22_X1  g646(.A1(new_n844), .A2(new_n678), .B1(new_n841), .B2(new_n643), .ZN(new_n848));
  OAI211_X1 g647(.A(new_n847), .B(KEYINPUT115), .C1(new_n848), .C2(new_n577), .ZN(new_n849));
  NAND3_X1  g648(.A1(new_n846), .A2(new_n849), .A3(new_n781), .ZN(new_n850));
  OAI21_X1  g649(.A(KEYINPUT113), .B1(new_n645), .B2(new_n678), .ZN(new_n851));
  INV_X1    g650(.A(new_n755), .ZN(new_n852));
  INV_X1    g651(.A(KEYINPUT113), .ZN(new_n853));
  NAND4_X1  g652(.A1(new_n852), .A2(new_n853), .A3(new_n679), .A4(new_n644), .ZN(new_n854));
  NAND2_X1  g653(.A1(new_n851), .A2(new_n854), .ZN(new_n855));
  AOI21_X1  g654(.A(new_n312), .B1(new_n850), .B2(new_n855), .ZN(new_n856));
  INV_X1    g655(.A(new_n449), .ZN(new_n857));
  NOR2_X1   g656(.A1(new_n857), .A2(new_n383), .ZN(new_n858));
  NAND2_X1  g657(.A1(new_n856), .A2(new_n858), .ZN(new_n859));
  NOR3_X1   g658(.A1(new_n859), .A2(G113gat), .A3(new_n679), .ZN(new_n860));
  AOI21_X1  g659(.A(new_n746), .B1(new_n850), .B2(new_n855), .ZN(new_n861));
  AND4_X1   g660(.A1(new_n683), .A2(new_n861), .A3(new_n384), .A4(new_n696), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n862), .A2(new_n678), .ZN(new_n863));
  AOI21_X1  g662(.A(new_n860), .B1(G113gat), .B2(new_n863), .ZN(new_n864));
  XOR2_X1   g663(.A(new_n864), .B(KEYINPUT116), .Z(G1340gat));
  INV_X1    g664(.A(new_n859), .ZN(new_n866));
  AOI21_X1  g665(.A(G120gat), .B1(new_n866), .B2(new_n643), .ZN(new_n867));
  NOR2_X1   g666(.A1(new_n644), .A2(new_n228), .ZN(new_n868));
  AOI21_X1  g667(.A(new_n867), .B1(new_n862), .B2(new_n868), .ZN(G1341gat));
  NAND2_X1  g668(.A1(new_n866), .A2(new_n623), .ZN(new_n870));
  NOR2_X1   g669(.A1(new_n216), .A2(new_n217), .ZN(new_n871));
  NOR2_X1   g670(.A1(new_n781), .A2(new_n871), .ZN(new_n872));
  AOI22_X1  g671(.A1(new_n870), .A2(new_n871), .B1(new_n862), .B2(new_n872), .ZN(new_n873));
  XOR2_X1   g672(.A(new_n873), .B(KEYINPUT117), .Z(G1342gat));
  INV_X1    g673(.A(G134gat), .ZN(new_n875));
  NAND3_X1  g674(.A1(new_n866), .A2(new_n875), .A3(new_n577), .ZN(new_n876));
  AND2_X1   g675(.A1(new_n876), .A2(KEYINPUT56), .ZN(new_n877));
  AOI21_X1  g676(.A(new_n875), .B1(new_n862), .B2(new_n577), .ZN(new_n878));
  NOR2_X1   g677(.A1(new_n877), .A2(new_n878), .ZN(new_n879));
  OAI21_X1  g678(.A(new_n879), .B1(KEYINPUT56), .B2(new_n876), .ZN(G1343gat));
  XOR2_X1   g679(.A(KEYINPUT121), .B(KEYINPUT58), .Z(new_n881));
  NAND2_X1  g680(.A1(new_n700), .A2(new_n456), .ZN(new_n882));
  NOR2_X1   g681(.A1(new_n882), .A2(new_n383), .ZN(new_n883));
  AND2_X1   g682(.A1(new_n856), .A2(new_n883), .ZN(new_n884));
  INV_X1    g683(.A(new_n884), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n678), .A2(new_n208), .ZN(new_n886));
  XOR2_X1   g685(.A(new_n886), .B(KEYINPUT120), .Z(new_n887));
  AOI211_X1 g686(.A(KEYINPUT57), .B(new_n420), .C1(new_n850), .C2(new_n855), .ZN(new_n888));
  NOR2_X1   g687(.A1(new_n515), .A2(new_n383), .ZN(new_n889));
  NAND2_X1  g688(.A1(new_n683), .A2(new_n889), .ZN(new_n890));
  INV_X1    g689(.A(new_n890), .ZN(new_n891));
  OAI21_X1  g690(.A(new_n781), .B1(new_n843), .B2(new_n845), .ZN(new_n892));
  AOI21_X1  g691(.A(new_n465), .B1(new_n892), .B2(new_n855), .ZN(new_n893));
  INV_X1    g692(.A(KEYINPUT57), .ZN(new_n894));
  OAI21_X1  g693(.A(new_n891), .B1(new_n893), .B2(new_n894), .ZN(new_n895));
  NOR3_X1   g694(.A1(new_n888), .A2(new_n679), .A3(new_n895), .ZN(new_n896));
  OAI221_X1 g695(.A(new_n881), .B1(new_n885), .B2(new_n887), .C1(new_n208), .C2(new_n896), .ZN(new_n897));
  INV_X1    g696(.A(KEYINPUT118), .ZN(new_n898));
  OAI21_X1  g697(.A(new_n898), .B1(new_n888), .B2(new_n895), .ZN(new_n899));
  AOI21_X1  g698(.A(new_n420), .B1(new_n850), .B2(new_n855), .ZN(new_n900));
  NAND2_X1  g699(.A1(new_n900), .A2(new_n894), .ZN(new_n901));
  NAND2_X1  g700(.A1(new_n892), .A2(new_n855), .ZN(new_n902));
  NAND2_X1  g701(.A1(new_n902), .A2(new_n746), .ZN(new_n903));
  AOI21_X1  g702(.A(new_n890), .B1(new_n903), .B2(KEYINPUT57), .ZN(new_n904));
  NAND3_X1  g703(.A1(new_n901), .A2(new_n904), .A3(KEYINPUT118), .ZN(new_n905));
  NAND3_X1  g704(.A1(new_n899), .A2(new_n905), .A3(new_n678), .ZN(new_n906));
  INV_X1    g705(.A(KEYINPUT119), .ZN(new_n907));
  AND3_X1   g706(.A1(new_n906), .A2(new_n907), .A3(G141gat), .ZN(new_n908));
  AOI21_X1  g707(.A(new_n907), .B1(new_n906), .B2(G141gat), .ZN(new_n909));
  NOR2_X1   g708(.A1(new_n885), .A2(new_n887), .ZN(new_n910));
  NOR3_X1   g709(.A1(new_n908), .A2(new_n909), .A3(new_n910), .ZN(new_n911));
  INV_X1    g710(.A(KEYINPUT58), .ZN(new_n912));
  OAI21_X1  g711(.A(new_n897), .B1(new_n911), .B2(new_n912), .ZN(G1344gat));
  INV_X1    g712(.A(KEYINPUT59), .ZN(new_n914));
  AOI211_X1 g713(.A(new_n914), .B(G148gat), .C1(new_n884), .C2(new_n643), .ZN(new_n915));
  NAND2_X1  g714(.A1(new_n899), .A2(new_n905), .ZN(new_n916));
  OAI21_X1  g715(.A(new_n914), .B1(new_n916), .B2(new_n644), .ZN(new_n917));
  OAI21_X1  g716(.A(new_n892), .B1(new_n678), .B2(new_n645), .ZN(new_n918));
  NAND3_X1  g717(.A1(new_n918), .A2(new_n894), .A3(new_n746), .ZN(new_n919));
  OAI21_X1  g718(.A(new_n919), .B1(new_n900), .B2(new_n894), .ZN(new_n920));
  NAND3_X1  g719(.A1(new_n891), .A2(KEYINPUT59), .A3(new_n643), .ZN(new_n921));
  OAI21_X1  g720(.A(new_n917), .B1(new_n920), .B2(new_n921), .ZN(new_n922));
  AOI21_X1  g721(.A(new_n915), .B1(new_n922), .B2(G148gat), .ZN(G1345gat));
  OAI21_X1  g722(.A(G155gat), .B1(new_n916), .B2(new_n781), .ZN(new_n924));
  OR2_X1    g723(.A1(new_n781), .A2(G155gat), .ZN(new_n925));
  OAI21_X1  g724(.A(new_n924), .B1(new_n885), .B2(new_n925), .ZN(G1346gat));
  NOR3_X1   g725(.A1(new_n885), .A2(G162gat), .A3(new_n578), .ZN(new_n927));
  XNOR2_X1  g726(.A(new_n927), .B(KEYINPUT122), .ZN(new_n928));
  INV_X1    g727(.A(KEYINPUT123), .ZN(new_n929));
  NOR3_X1   g728(.A1(new_n916), .A2(new_n929), .A3(new_n578), .ZN(new_n930));
  OAI21_X1  g729(.A(new_n929), .B1(new_n916), .B2(new_n578), .ZN(new_n931));
  NAND2_X1  g730(.A1(new_n931), .A2(G162gat), .ZN(new_n932));
  OAI21_X1  g731(.A(new_n928), .B1(new_n930), .B2(new_n932), .ZN(G1347gat));
  AOI21_X1  g732(.A(new_n683), .B1(new_n850), .B2(new_n855), .ZN(new_n934));
  NOR2_X1   g733(.A1(new_n857), .A2(new_n384), .ZN(new_n935));
  NAND2_X1  g734(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  INV_X1    g735(.A(new_n936), .ZN(new_n937));
  AOI21_X1  g736(.A(G169gat), .B1(new_n937), .B2(new_n678), .ZN(new_n938));
  NAND4_X1  g737(.A1(new_n861), .A2(new_n312), .A3(new_n383), .A4(new_n696), .ZN(new_n939));
  NOR3_X1   g738(.A1(new_n939), .A2(new_n337), .A3(new_n679), .ZN(new_n940));
  NOR2_X1   g739(.A1(new_n938), .A2(new_n940), .ZN(G1348gat));
  OAI21_X1  g740(.A(G176gat), .B1(new_n939), .B2(new_n644), .ZN(new_n942));
  NAND2_X1  g741(.A1(new_n643), .A2(new_n338), .ZN(new_n943));
  OAI21_X1  g742(.A(new_n942), .B1(new_n936), .B2(new_n943), .ZN(G1349gat));
  OAI21_X1  g743(.A(G183gat), .B1(new_n939), .B2(new_n781), .ZN(new_n945));
  NAND2_X1  g744(.A1(new_n623), .A2(new_n347), .ZN(new_n946));
  OAI21_X1  g745(.A(new_n945), .B1(new_n936), .B2(new_n946), .ZN(new_n947));
  XNOR2_X1  g746(.A(new_n947), .B(KEYINPUT60), .ZN(G1350gat));
  OAI21_X1  g747(.A(G190gat), .B1(new_n939), .B2(new_n578), .ZN(new_n949));
  XNOR2_X1  g748(.A(new_n949), .B(KEYINPUT61), .ZN(new_n950));
  NAND3_X1  g749(.A1(new_n937), .A2(new_n349), .A3(new_n577), .ZN(new_n951));
  NAND2_X1  g750(.A1(new_n950), .A2(new_n951), .ZN(G1351gat));
  NOR2_X1   g751(.A1(new_n882), .A2(new_n384), .ZN(new_n953));
  NAND2_X1  g752(.A1(new_n934), .A2(new_n953), .ZN(new_n954));
  OR3_X1    g753(.A1(new_n954), .A2(G197gat), .A3(new_n679), .ZN(new_n955));
  NAND3_X1  g754(.A1(new_n700), .A2(new_n312), .A3(new_n383), .ZN(new_n956));
  OR2_X1    g755(.A1(new_n920), .A2(new_n956), .ZN(new_n957));
  OAI21_X1  g756(.A(KEYINPUT124), .B1(new_n957), .B2(new_n679), .ZN(new_n958));
  NAND2_X1  g757(.A1(new_n958), .A2(G197gat), .ZN(new_n959));
  NOR3_X1   g758(.A1(new_n957), .A2(KEYINPUT124), .A3(new_n679), .ZN(new_n960));
  OAI21_X1  g759(.A(new_n955), .B1(new_n959), .B2(new_n960), .ZN(G1352gat));
  XNOR2_X1  g760(.A(KEYINPUT125), .B(G204gat), .ZN(new_n962));
  NOR3_X1   g761(.A1(new_n954), .A2(new_n644), .A3(new_n962), .ZN(new_n963));
  XNOR2_X1  g762(.A(new_n963), .B(KEYINPUT62), .ZN(new_n964));
  OAI21_X1  g763(.A(new_n962), .B1(new_n957), .B2(new_n644), .ZN(new_n965));
  NAND2_X1  g764(.A1(new_n964), .A2(new_n965), .ZN(G1353gat));
  INV_X1    g765(.A(new_n954), .ZN(new_n967));
  NAND3_X1  g766(.A1(new_n967), .A2(new_n314), .A3(new_n623), .ZN(new_n968));
  INV_X1    g767(.A(new_n957), .ZN(new_n969));
  NAND2_X1  g768(.A1(new_n969), .A2(new_n623), .ZN(new_n970));
  INV_X1    g769(.A(KEYINPUT63), .ZN(new_n971));
  NOR2_X1   g770(.A1(new_n971), .A2(KEYINPUT126), .ZN(new_n972));
  AOI21_X1  g771(.A(new_n314), .B1(KEYINPUT126), .B2(new_n971), .ZN(new_n973));
  NAND3_X1  g772(.A1(new_n970), .A2(new_n972), .A3(new_n973), .ZN(new_n974));
  INV_X1    g773(.A(new_n974), .ZN(new_n975));
  AOI21_X1  g774(.A(new_n972), .B1(new_n970), .B2(new_n973), .ZN(new_n976));
  OAI21_X1  g775(.A(new_n968), .B1(new_n975), .B2(new_n976), .ZN(G1354gat));
  AOI21_X1  g776(.A(G218gat), .B1(new_n967), .B2(new_n577), .ZN(new_n978));
  AOI211_X1 g777(.A(new_n328), .B(new_n578), .C1(new_n969), .C2(KEYINPUT127), .ZN(new_n979));
  OR2_X1    g778(.A1(new_n969), .A2(KEYINPUT127), .ZN(new_n980));
  AOI21_X1  g779(.A(new_n978), .B1(new_n979), .B2(new_n980), .ZN(G1355gat));
endmodule


