//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 1 0 1 1 1 0 0 0 1 1 1 1 1 0 0 1 1 1 1 0 0 0 0 0 0 0 1 0 1 0 0 0 1 0 1 0 1 0 0 0 1 1 1 0 1 0 1 1 0 0 1 0 1 1 0 0 0 0 1 0 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:38:31 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n245, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1091, new_n1092, new_n1093,
    new_n1094, new_n1095, new_n1096, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1113, new_n1114, new_n1115, new_n1116, new_n1117, new_n1118,
    new_n1119, new_n1120, new_n1121, new_n1122, new_n1123, new_n1124,
    new_n1125, new_n1126, new_n1127, new_n1128, new_n1129, new_n1130,
    new_n1131, new_n1132, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1255, new_n1256, new_n1257, new_n1258,
    new_n1260, new_n1261, new_n1262, new_n1263, new_n1264, new_n1265,
    new_n1266, new_n1267, new_n1268, new_n1269, new_n1270, new_n1271,
    new_n1272, new_n1273, new_n1274, new_n1275, new_n1276, new_n1277,
    new_n1278, new_n1279, new_n1280, new_n1281, new_n1283, new_n1284,
    new_n1285, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1349, new_n1350, new_n1351, new_n1352, new_n1353,
    new_n1354, new_n1355, new_n1356, new_n1357, new_n1358, new_n1359,
    new_n1360, new_n1361, new_n1362, new_n1363, new_n1364, new_n1365,
    new_n1366, new_n1367;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(new_n201), .ZN(new_n202));
  NOR3_X1   g0002(.A1(new_n202), .A2(G50), .A3(G77), .ZN(G353));
  OAI21_X1  g0003(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0004(.A(G1), .ZN(new_n205));
  INV_X1    g0005(.A(G20), .ZN(new_n206));
  NOR2_X1   g0006(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  INV_X1    g0007(.A(new_n207), .ZN(new_n208));
  AOI22_X1  g0008(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n209));
  XNOR2_X1  g0009(.A(new_n209), .B(KEYINPUT65), .ZN(new_n210));
  AOI22_X1  g0010(.A1(G87), .A2(G250), .B1(G116), .B2(G270), .ZN(new_n211));
  AOI22_X1  g0011(.A1(G50), .A2(G226), .B1(G68), .B2(G238), .ZN(new_n212));
  AOI22_X1  g0012(.A1(G77), .A2(G244), .B1(G97), .B2(G257), .ZN(new_n213));
  NAND3_X1  g0013(.A1(new_n211), .A2(new_n212), .A3(new_n213), .ZN(new_n214));
  OAI21_X1  g0014(.A(new_n208), .B1(new_n210), .B2(new_n214), .ZN(new_n215));
  XOR2_X1   g0015(.A(new_n215), .B(KEYINPUT66), .Z(new_n216));
  INV_X1    g0016(.A(KEYINPUT1), .ZN(new_n217));
  OR2_X1    g0017(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  NAND2_X1  g0018(.A1(new_n216), .A2(new_n217), .ZN(new_n219));
  NOR2_X1   g0019(.A1(new_n208), .A2(G13), .ZN(new_n220));
  OAI211_X1 g0020(.A(new_n220), .B(G250), .C1(G257), .C2(G264), .ZN(new_n221));
  XNOR2_X1  g0021(.A(KEYINPUT64), .B(KEYINPUT0), .ZN(new_n222));
  XNOR2_X1  g0022(.A(new_n221), .B(new_n222), .ZN(new_n223));
  NAND2_X1  g0023(.A1(G1), .A2(G13), .ZN(new_n224));
  NOR2_X1   g0024(.A1(new_n224), .A2(new_n206), .ZN(new_n225));
  NAND2_X1  g0025(.A1(new_n202), .A2(G50), .ZN(new_n226));
  INV_X1    g0026(.A(new_n226), .ZN(new_n227));
  AOI21_X1  g0027(.A(new_n223), .B1(new_n225), .B2(new_n227), .ZN(new_n228));
  AND3_X1   g0028(.A1(new_n218), .A2(new_n219), .A3(new_n228), .ZN(G361));
  XNOR2_X1  g0029(.A(G238), .B(G244), .ZN(new_n230));
  INV_X1    g0030(.A(G232), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n230), .B(new_n231), .ZN(new_n232));
  XOR2_X1   g0032(.A(KEYINPUT2), .B(G226), .Z(new_n233));
  XNOR2_X1  g0033(.A(new_n232), .B(new_n233), .ZN(new_n234));
  XOR2_X1   g0034(.A(G264), .B(G270), .Z(new_n235));
  XNOR2_X1  g0035(.A(G250), .B(G257), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n234), .B(new_n237), .ZN(G358));
  XOR2_X1   g0038(.A(G87), .B(G97), .Z(new_n239));
  XNOR2_X1  g0039(.A(new_n239), .B(KEYINPUT67), .ZN(new_n240));
  XOR2_X1   g0040(.A(G107), .B(G116), .Z(new_n241));
  XOR2_X1   g0041(.A(new_n240), .B(new_n241), .Z(new_n242));
  XNOR2_X1  g0042(.A(G50), .B(G68), .ZN(new_n243));
  XNOR2_X1  g0043(.A(G58), .B(G77), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n242), .B(new_n245), .ZN(G351));
  INV_X1    g0046(.A(KEYINPUT10), .ZN(new_n247));
  NOR2_X1   g0047(.A1(new_n247), .A2(KEYINPUT74), .ZN(new_n248));
  AOI21_X1  g0048(.A(new_n224), .B1(G33), .B2(G41), .ZN(new_n249));
  NOR2_X1   g0049(.A1(KEYINPUT68), .A2(G1698), .ZN(new_n250));
  INV_X1    g0050(.A(new_n250), .ZN(new_n251));
  INV_X1    g0051(.A(G33), .ZN(new_n252));
  NAND2_X1  g0052(.A1(new_n252), .A2(KEYINPUT3), .ZN(new_n253));
  INV_X1    g0053(.A(KEYINPUT3), .ZN(new_n254));
  NAND2_X1  g0054(.A1(new_n254), .A2(G33), .ZN(new_n255));
  NAND2_X1  g0055(.A1(KEYINPUT68), .A2(G1698), .ZN(new_n256));
  NAND4_X1  g0056(.A1(new_n251), .A2(new_n253), .A3(new_n255), .A4(new_n256), .ZN(new_n257));
  INV_X1    g0057(.A(G222), .ZN(new_n258));
  INV_X1    g0058(.A(G77), .ZN(new_n259));
  XNOR2_X1  g0059(.A(KEYINPUT3), .B(G33), .ZN(new_n260));
  OAI22_X1  g0060(.A1(new_n257), .A2(new_n258), .B1(new_n259), .B2(new_n260), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n253), .A2(new_n255), .ZN(new_n262));
  INV_X1    g0062(.A(G223), .ZN(new_n263));
  INV_X1    g0063(.A(G1698), .ZN(new_n264));
  NOR3_X1   g0064(.A1(new_n262), .A2(new_n263), .A3(new_n264), .ZN(new_n265));
  OAI21_X1  g0065(.A(new_n249), .B1(new_n261), .B2(new_n265), .ZN(new_n266));
  INV_X1    g0066(.A(G274), .ZN(new_n267));
  OAI21_X1  g0067(.A(new_n205), .B1(G41), .B2(G45), .ZN(new_n268));
  NOR3_X1   g0068(.A1(new_n249), .A2(new_n267), .A3(new_n268), .ZN(new_n269));
  AND2_X1   g0069(.A1(G1), .A2(G13), .ZN(new_n270));
  NAND2_X1  g0070(.A1(G33), .A2(G41), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n272), .A2(new_n268), .ZN(new_n273));
  INV_X1    g0073(.A(new_n273), .ZN(new_n274));
  AOI21_X1  g0074(.A(new_n269), .B1(G226), .B2(new_n274), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n266), .A2(new_n275), .ZN(new_n276));
  INV_X1    g0076(.A(new_n276), .ZN(new_n277));
  AOI21_X1  g0077(.A(new_n248), .B1(new_n277), .B2(G190), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n276), .A2(G200), .ZN(new_n279));
  AND2_X1   g0079(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  NAND3_X1  g0080(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n281), .A2(new_n224), .ZN(new_n282));
  XNOR2_X1  g0082(.A(KEYINPUT8), .B(G58), .ZN(new_n283));
  XNOR2_X1  g0083(.A(new_n283), .B(KEYINPUT69), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n206), .A2(G33), .ZN(new_n285));
  XNOR2_X1  g0085(.A(new_n285), .B(KEYINPUT70), .ZN(new_n286));
  NOR2_X1   g0086(.A1(new_n284), .A2(new_n286), .ZN(new_n287));
  NOR2_X1   g0087(.A1(new_n202), .A2(G50), .ZN(new_n288));
  OR3_X1    g0088(.A1(new_n288), .A2(KEYINPUT71), .A3(new_n206), .ZN(new_n289));
  NOR2_X1   g0089(.A1(G20), .A2(G33), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n290), .A2(G150), .ZN(new_n291));
  OAI21_X1  g0091(.A(KEYINPUT71), .B1(new_n288), .B2(new_n206), .ZN(new_n292));
  NAND3_X1  g0092(.A1(new_n289), .A2(new_n291), .A3(new_n292), .ZN(new_n293));
  OAI21_X1  g0093(.A(new_n282), .B1(new_n287), .B2(new_n293), .ZN(new_n294));
  NAND3_X1  g0094(.A1(new_n205), .A2(G13), .A3(G20), .ZN(new_n295));
  INV_X1    g0095(.A(new_n295), .ZN(new_n296));
  NOR2_X1   g0096(.A1(new_n296), .A2(new_n282), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n297), .A2(KEYINPUT72), .ZN(new_n298));
  INV_X1    g0098(.A(KEYINPUT72), .ZN(new_n299));
  OAI21_X1  g0099(.A(new_n299), .B1(new_n296), .B2(new_n282), .ZN(new_n300));
  OAI211_X1 g0100(.A(new_n298), .B(new_n300), .C1(G1), .C2(new_n206), .ZN(new_n301));
  INV_X1    g0101(.A(G50), .ZN(new_n302));
  OR2_X1    g0102(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n296), .A2(new_n302), .ZN(new_n304));
  NAND3_X1  g0104(.A1(new_n294), .A2(new_n303), .A3(new_n304), .ZN(new_n305));
  INV_X1    g0105(.A(KEYINPUT9), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n305), .A2(new_n306), .ZN(new_n307));
  NAND4_X1  g0107(.A1(new_n294), .A2(new_n303), .A3(KEYINPUT9), .A4(new_n304), .ZN(new_n308));
  NAND3_X1  g0108(.A1(new_n280), .A2(new_n307), .A3(new_n308), .ZN(new_n309));
  NAND3_X1  g0109(.A1(new_n309), .A2(KEYINPUT74), .A3(new_n247), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n247), .A2(KEYINPUT74), .ZN(new_n311));
  NAND4_X1  g0111(.A1(new_n280), .A2(new_n311), .A3(new_n307), .A4(new_n308), .ZN(new_n312));
  NOR2_X1   g0112(.A1(new_n276), .A2(G179), .ZN(new_n313));
  INV_X1    g0113(.A(G169), .ZN(new_n314));
  AOI21_X1  g0114(.A(new_n313), .B1(new_n314), .B2(new_n276), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n315), .A2(new_n305), .ZN(new_n316));
  NAND3_X1  g0116(.A1(new_n310), .A2(new_n312), .A3(new_n316), .ZN(new_n317));
  INV_X1    g0117(.A(new_n317), .ZN(new_n318));
  INV_X1    g0118(.A(KEYINPUT69), .ZN(new_n319));
  XNOR2_X1  g0119(.A(new_n283), .B(new_n319), .ZN(new_n320));
  NOR2_X1   g0120(.A1(new_n320), .A2(new_n296), .ZN(new_n321));
  AOI21_X1  g0121(.A(new_n321), .B1(new_n301), .B2(new_n320), .ZN(new_n322));
  INV_X1    g0122(.A(new_n282), .ZN(new_n323));
  INV_X1    g0123(.A(G58), .ZN(new_n324));
  INV_X1    g0124(.A(G68), .ZN(new_n325));
  NOR2_X1   g0125(.A1(new_n324), .A2(new_n325), .ZN(new_n326));
  OAI21_X1  g0126(.A(G20), .B1(new_n326), .B2(new_n201), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n290), .A2(G159), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n327), .A2(new_n328), .ZN(new_n329));
  INV_X1    g0129(.A(KEYINPUT78), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n330), .A2(new_n254), .ZN(new_n331));
  NAND2_X1  g0131(.A1(KEYINPUT78), .A2(KEYINPUT3), .ZN(new_n332));
  NAND3_X1  g0132(.A1(new_n331), .A2(G33), .A3(new_n332), .ZN(new_n333));
  AOI21_X1  g0133(.A(G20), .B1(new_n333), .B2(new_n253), .ZN(new_n334));
  INV_X1    g0134(.A(KEYINPUT7), .ZN(new_n335));
  AOI21_X1  g0135(.A(new_n325), .B1(new_n334), .B2(new_n335), .ZN(new_n336));
  INV_X1    g0136(.A(new_n253), .ZN(new_n337));
  AND2_X1   g0137(.A1(KEYINPUT78), .A2(KEYINPUT3), .ZN(new_n338));
  NOR2_X1   g0138(.A1(KEYINPUT78), .A2(KEYINPUT3), .ZN(new_n339));
  NOR2_X1   g0139(.A1(new_n338), .A2(new_n339), .ZN(new_n340));
  AOI21_X1  g0140(.A(new_n337), .B1(new_n340), .B2(G33), .ZN(new_n341));
  OAI21_X1  g0141(.A(KEYINPUT7), .B1(new_n341), .B2(G20), .ZN(new_n342));
  AOI21_X1  g0142(.A(new_n329), .B1(new_n336), .B2(new_n342), .ZN(new_n343));
  AOI21_X1  g0143(.A(new_n323), .B1(new_n343), .B2(KEYINPUT16), .ZN(new_n344));
  INV_X1    g0144(.A(KEYINPUT16), .ZN(new_n345));
  NOR2_X1   g0145(.A1(new_n335), .A2(G20), .ZN(new_n346));
  AOI21_X1  g0146(.A(G33), .B1(new_n331), .B2(new_n332), .ZN(new_n347));
  INV_X1    g0147(.A(new_n255), .ZN(new_n348));
  OAI21_X1  g0148(.A(new_n346), .B1(new_n347), .B2(new_n348), .ZN(new_n349));
  OAI21_X1  g0149(.A(new_n335), .B1(new_n260), .B2(G20), .ZN(new_n350));
  AOI21_X1  g0150(.A(new_n325), .B1(new_n349), .B2(new_n350), .ZN(new_n351));
  OAI21_X1  g0151(.A(new_n345), .B1(new_n351), .B2(new_n329), .ZN(new_n352));
  AOI21_X1  g0152(.A(new_n322), .B1(new_n344), .B2(new_n352), .ZN(new_n353));
  AOI21_X1  g0153(.A(new_n267), .B1(new_n270), .B2(new_n271), .ZN(new_n354));
  INV_X1    g0154(.A(new_n268), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  OAI21_X1  g0156(.A(new_n356), .B1(new_n273), .B2(new_n231), .ZN(new_n357));
  AND2_X1   g0157(.A1(KEYINPUT68), .A2(G1698), .ZN(new_n358));
  NOR2_X1   g0158(.A1(new_n358), .A2(new_n250), .ZN(new_n359));
  AOI22_X1  g0159(.A1(new_n359), .A2(G223), .B1(G226), .B2(G1698), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n333), .A2(new_n253), .ZN(new_n361));
  INV_X1    g0161(.A(G87), .ZN(new_n362));
  OAI22_X1  g0162(.A1(new_n360), .A2(new_n361), .B1(new_n252), .B2(new_n362), .ZN(new_n363));
  AOI21_X1  g0163(.A(new_n357), .B1(new_n363), .B2(new_n249), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n364), .A2(G179), .ZN(new_n365));
  AOI22_X1  g0165(.A1(new_n274), .A2(G232), .B1(new_n354), .B2(new_n355), .ZN(new_n366));
  NOR2_X1   g0166(.A1(new_n252), .A2(new_n362), .ZN(new_n367));
  XNOR2_X1  g0167(.A(KEYINPUT68), .B(G1698), .ZN(new_n368));
  INV_X1    g0168(.A(G226), .ZN(new_n369));
  OAI22_X1  g0169(.A1(new_n368), .A2(new_n263), .B1(new_n369), .B2(new_n264), .ZN(new_n370));
  AOI21_X1  g0170(.A(new_n367), .B1(new_n370), .B2(new_n341), .ZN(new_n371));
  OAI21_X1  g0171(.A(new_n366), .B1(new_n371), .B2(new_n272), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n372), .A2(G169), .ZN(new_n373));
  AND2_X1   g0173(.A1(new_n365), .A2(new_n373), .ZN(new_n374));
  OAI21_X1  g0174(.A(KEYINPUT18), .B1(new_n353), .B2(new_n374), .ZN(new_n375));
  INV_X1    g0175(.A(new_n329), .ZN(new_n376));
  NOR3_X1   g0176(.A1(new_n338), .A2(new_n339), .A3(new_n252), .ZN(new_n377));
  OAI211_X1 g0177(.A(new_n335), .B(new_n206), .C1(new_n377), .C2(new_n337), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n378), .A2(G68), .ZN(new_n379));
  NOR2_X1   g0179(.A1(new_n334), .A2(new_n335), .ZN(new_n380));
  OAI211_X1 g0180(.A(KEYINPUT16), .B(new_n376), .C1(new_n379), .C2(new_n380), .ZN(new_n381));
  NAND3_X1  g0181(.A1(new_n381), .A2(new_n352), .A3(new_n282), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n301), .A2(new_n320), .ZN(new_n383));
  OAI21_X1  g0183(.A(new_n383), .B1(new_n296), .B2(new_n320), .ZN(new_n384));
  AOI22_X1  g0184(.A1(new_n382), .A2(new_n384), .B1(new_n373), .B2(new_n365), .ZN(new_n385));
  INV_X1    g0185(.A(KEYINPUT18), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n385), .A2(new_n386), .ZN(new_n387));
  INV_X1    g0187(.A(G190), .ZN(new_n388));
  OAI211_X1 g0188(.A(new_n388), .B(new_n366), .C1(new_n371), .C2(new_n272), .ZN(new_n389));
  OAI21_X1  g0189(.A(new_n389), .B1(new_n364), .B2(G200), .ZN(new_n390));
  NAND3_X1  g0190(.A1(new_n382), .A2(new_n390), .A3(new_n384), .ZN(new_n391));
  INV_X1    g0191(.A(KEYINPUT17), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n391), .A2(new_n392), .ZN(new_n393));
  NAND4_X1  g0193(.A1(new_n382), .A2(new_n390), .A3(new_n384), .A4(KEYINPUT17), .ZN(new_n394));
  NAND4_X1  g0194(.A1(new_n375), .A2(new_n387), .A3(new_n393), .A4(new_n394), .ZN(new_n395));
  INV_X1    g0195(.A(new_n395), .ZN(new_n396));
  NAND3_X1  g0196(.A1(new_n272), .A2(G238), .A3(new_n268), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n356), .A2(new_n397), .ZN(new_n398));
  NAND3_X1  g0198(.A1(new_n260), .A2(G232), .A3(G1698), .ZN(new_n399));
  NAND2_X1  g0199(.A1(G33), .A2(G97), .ZN(new_n400));
  OAI211_X1 g0200(.A(new_n399), .B(new_n400), .C1(new_n369), .C2(new_n257), .ZN(new_n401));
  AOI21_X1  g0201(.A(new_n398), .B1(new_n401), .B2(new_n249), .ZN(new_n402));
  XNOR2_X1  g0202(.A(KEYINPUT75), .B(KEYINPUT13), .ZN(new_n403));
  INV_X1    g0203(.A(new_n403), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n402), .A2(new_n404), .ZN(new_n405));
  INV_X1    g0205(.A(KEYINPUT13), .ZN(new_n406));
  OAI211_X1 g0206(.A(new_n405), .B(G190), .C1(new_n406), .C2(new_n402), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n401), .A2(new_n249), .ZN(new_n408));
  INV_X1    g0208(.A(new_n398), .ZN(new_n409));
  AOI21_X1  g0209(.A(new_n404), .B1(new_n408), .B2(new_n409), .ZN(new_n410));
  AOI211_X1 g0210(.A(new_n403), .B(new_n398), .C1(new_n401), .C2(new_n249), .ZN(new_n411));
  OAI21_X1  g0211(.A(G200), .B1(new_n410), .B2(new_n411), .ZN(new_n412));
  AOI22_X1  g0212(.A1(new_n290), .A2(G50), .B1(G20), .B2(new_n325), .ZN(new_n413));
  OAI21_X1  g0213(.A(new_n413), .B1(new_n286), .B2(new_n259), .ZN(new_n414));
  NAND3_X1  g0214(.A1(new_n414), .A2(KEYINPUT11), .A3(new_n282), .ZN(new_n415));
  OAI21_X1  g0215(.A(KEYINPUT12), .B1(new_n295), .B2(G68), .ZN(new_n416));
  OR3_X1    g0216(.A1(new_n295), .A2(KEYINPUT12), .A3(G68), .ZN(new_n417));
  AOI21_X1  g0217(.A(new_n325), .B1(new_n205), .B2(G20), .ZN(new_n418));
  AOI22_X1  g0218(.A1(new_n416), .A2(new_n417), .B1(new_n297), .B2(new_n418), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n415), .A2(new_n419), .ZN(new_n420));
  AOI21_X1  g0220(.A(KEYINPUT11), .B1(new_n414), .B2(new_n282), .ZN(new_n421));
  NOR2_X1   g0221(.A1(new_n420), .A2(new_n421), .ZN(new_n422));
  NAND3_X1  g0222(.A1(new_n407), .A2(new_n412), .A3(new_n422), .ZN(new_n423));
  INV_X1    g0223(.A(new_n423), .ZN(new_n424));
  OAI21_X1  g0224(.A(G169), .B1(new_n410), .B2(new_n411), .ZN(new_n425));
  NAND2_X1  g0225(.A1(KEYINPUT76), .A2(KEYINPUT14), .ZN(new_n426));
  INV_X1    g0226(.A(new_n426), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n425), .A2(new_n427), .ZN(new_n428));
  OAI211_X1 g0228(.A(new_n405), .B(G179), .C1(new_n406), .C2(new_n402), .ZN(new_n429));
  OAI211_X1 g0229(.A(G169), .B(new_n426), .C1(new_n410), .C2(new_n411), .ZN(new_n430));
  NAND3_X1  g0230(.A1(new_n428), .A2(new_n429), .A3(new_n430), .ZN(new_n431));
  INV_X1    g0231(.A(KEYINPUT77), .ZN(new_n432));
  OAI21_X1  g0232(.A(new_n432), .B1(new_n420), .B2(new_n421), .ZN(new_n433));
  INV_X1    g0233(.A(new_n421), .ZN(new_n434));
  NAND4_X1  g0234(.A1(new_n434), .A2(KEYINPUT77), .A3(new_n415), .A4(new_n419), .ZN(new_n435));
  AND2_X1   g0235(.A1(new_n433), .A2(new_n435), .ZN(new_n436));
  AOI21_X1  g0236(.A(new_n424), .B1(new_n431), .B2(new_n436), .ZN(new_n437));
  INV_X1    g0237(.A(new_n290), .ZN(new_n438));
  OAI22_X1  g0238(.A1(new_n283), .A2(new_n438), .B1(new_n206), .B2(new_n259), .ZN(new_n439));
  XNOR2_X1  g0239(.A(KEYINPUT15), .B(G87), .ZN(new_n440));
  NOR2_X1   g0240(.A1(new_n440), .A2(new_n285), .ZN(new_n441));
  OAI21_X1  g0241(.A(new_n282), .B1(new_n439), .B2(new_n441), .ZN(new_n442));
  AOI21_X1  g0242(.A(new_n259), .B1(new_n205), .B2(G20), .ZN(new_n443));
  AOI22_X1  g0243(.A1(new_n297), .A2(new_n443), .B1(new_n259), .B2(new_n296), .ZN(new_n444));
  AND2_X1   g0244(.A1(new_n442), .A2(new_n444), .ZN(new_n445));
  NAND3_X1  g0245(.A1(new_n359), .A2(new_n260), .A3(G232), .ZN(new_n446));
  NAND3_X1  g0246(.A1(new_n260), .A2(G238), .A3(G1698), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n262), .A2(G107), .ZN(new_n448));
  NAND3_X1  g0248(.A1(new_n446), .A2(new_n447), .A3(new_n448), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n449), .A2(new_n249), .ZN(new_n450));
  AOI21_X1  g0250(.A(new_n269), .B1(G244), .B2(new_n274), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n452), .A2(KEYINPUT73), .ZN(new_n453));
  INV_X1    g0253(.A(KEYINPUT73), .ZN(new_n454));
  NAND3_X1  g0254(.A1(new_n450), .A2(new_n451), .A3(new_n454), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n453), .A2(new_n455), .ZN(new_n456));
  INV_X1    g0256(.A(G179), .ZN(new_n457));
  AOI21_X1  g0257(.A(new_n445), .B1(new_n456), .B2(new_n457), .ZN(new_n458));
  NAND3_X1  g0258(.A1(new_n453), .A2(new_n314), .A3(new_n455), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  INV_X1    g0260(.A(new_n455), .ZN(new_n461));
  AOI21_X1  g0261(.A(new_n454), .B1(new_n450), .B2(new_n451), .ZN(new_n462));
  OAI21_X1  g0262(.A(G190), .B1(new_n461), .B2(new_n462), .ZN(new_n463));
  NAND3_X1  g0263(.A1(new_n453), .A2(G200), .A3(new_n455), .ZN(new_n464));
  NAND3_X1  g0264(.A1(new_n463), .A2(new_n464), .A3(new_n445), .ZN(new_n465));
  AND2_X1   g0265(.A1(new_n460), .A2(new_n465), .ZN(new_n466));
  NAND4_X1  g0266(.A1(new_n318), .A2(new_n396), .A3(new_n437), .A4(new_n466), .ZN(new_n467));
  INV_X1    g0267(.A(new_n467), .ZN(new_n468));
  INV_X1    g0268(.A(KEYINPUT80), .ZN(new_n469));
  INV_X1    g0269(.A(G41), .ZN(new_n470));
  NAND3_X1  g0270(.A1(new_n469), .A2(new_n470), .A3(KEYINPUT5), .ZN(new_n471));
  INV_X1    g0271(.A(KEYINPUT5), .ZN(new_n472));
  OAI21_X1  g0272(.A(new_n472), .B1(KEYINPUT80), .B2(G41), .ZN(new_n473));
  INV_X1    g0273(.A(G45), .ZN(new_n474));
  NOR2_X1   g0274(.A1(new_n474), .A2(G1), .ZN(new_n475));
  NAND3_X1  g0275(.A1(new_n471), .A2(new_n473), .A3(new_n475), .ZN(new_n476));
  NAND3_X1  g0276(.A1(new_n476), .A2(G264), .A3(new_n272), .ZN(new_n477));
  INV_X1    g0277(.A(KEYINPUT91), .ZN(new_n478));
  OR2_X1    g0278(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n477), .A2(new_n478), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  NAND4_X1  g0281(.A1(new_n354), .A2(new_n471), .A3(new_n473), .A4(new_n475), .ZN(new_n482));
  NAND4_X1  g0282(.A1(new_n333), .A2(new_n359), .A3(G250), .A4(new_n253), .ZN(new_n483));
  NAND2_X1  g0283(.A1(G33), .A2(G294), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  INV_X1    g0285(.A(G257), .ZN(new_n486));
  NOR2_X1   g0286(.A1(new_n486), .A2(new_n264), .ZN(new_n487));
  NAND3_X1  g0287(.A1(new_n333), .A2(new_n253), .A3(new_n487), .ZN(new_n488));
  INV_X1    g0288(.A(KEYINPUT90), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  NAND4_X1  g0290(.A1(new_n333), .A2(KEYINPUT90), .A3(new_n253), .A4(new_n487), .ZN(new_n491));
  AOI21_X1  g0291(.A(new_n485), .B1(new_n490), .B2(new_n491), .ZN(new_n492));
  OAI211_X1 g0292(.A(new_n481), .B(new_n482), .C1(new_n492), .C2(new_n272), .ZN(new_n493));
  INV_X1    g0293(.A(new_n493), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n494), .A2(G190), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n493), .A2(G200), .ZN(new_n496));
  INV_X1    g0296(.A(KEYINPUT22), .ZN(new_n497));
  NOR2_X1   g0297(.A1(new_n497), .A2(new_n362), .ZN(new_n498));
  NAND4_X1  g0298(.A1(new_n333), .A2(new_n206), .A3(new_n253), .A4(new_n498), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n206), .A2(G87), .ZN(new_n500));
  OAI21_X1  g0300(.A(new_n497), .B1(new_n262), .B2(new_n500), .ZN(new_n501));
  INV_X1    g0301(.A(KEYINPUT23), .ZN(new_n502));
  OAI21_X1  g0302(.A(new_n502), .B1(new_n206), .B2(G107), .ZN(new_n503));
  INV_X1    g0303(.A(G107), .ZN(new_n504));
  NAND3_X1  g0304(.A1(new_n504), .A2(KEYINPUT23), .A3(G20), .ZN(new_n505));
  INV_X1    g0305(.A(G116), .ZN(new_n506));
  NOR2_X1   g0306(.A1(new_n252), .A2(new_n506), .ZN(new_n507));
  AOI22_X1  g0307(.A1(new_n503), .A2(new_n505), .B1(new_n507), .B2(new_n206), .ZN(new_n508));
  NAND3_X1  g0308(.A1(new_n499), .A2(new_n501), .A3(new_n508), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n509), .A2(KEYINPUT24), .ZN(new_n510));
  INV_X1    g0310(.A(KEYINPUT24), .ZN(new_n511));
  NAND4_X1  g0311(.A1(new_n499), .A2(new_n501), .A3(new_n511), .A4(new_n508), .ZN(new_n512));
  AOI21_X1  g0312(.A(new_n323), .B1(new_n510), .B2(new_n512), .ZN(new_n513));
  INV_X1    g0313(.A(KEYINPUT25), .ZN(new_n514));
  AOI211_X1 g0314(.A(G107), .B(new_n295), .C1(KEYINPUT88), .C2(new_n514), .ZN(new_n515));
  NOR2_X1   g0315(.A1(new_n514), .A2(KEYINPUT88), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  INV_X1    g0317(.A(new_n517), .ZN(new_n518));
  NOR2_X1   g0318(.A1(new_n515), .A2(new_n516), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n205), .A2(G33), .ZN(new_n520));
  NAND4_X1  g0320(.A1(new_n295), .A2(new_n520), .A3(new_n224), .A4(new_n281), .ZN(new_n521));
  OAI22_X1  g0321(.A1(new_n518), .A2(new_n519), .B1(new_n504), .B2(new_n521), .ZN(new_n522));
  NOR2_X1   g0322(.A1(new_n513), .A2(new_n522), .ZN(new_n523));
  NAND3_X1  g0323(.A1(new_n495), .A2(new_n496), .A3(new_n523), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n354), .A2(new_n475), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n205), .A2(G45), .ZN(new_n526));
  NAND3_X1  g0326(.A1(new_n272), .A2(G250), .A3(new_n526), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n525), .A2(new_n527), .ZN(new_n528));
  AOI22_X1  g0328(.A1(new_n359), .A2(G238), .B1(G244), .B2(G1698), .ZN(new_n529));
  OAI22_X1  g0329(.A1(new_n529), .A2(new_n361), .B1(new_n252), .B2(new_n506), .ZN(new_n530));
  AOI21_X1  g0330(.A(new_n528), .B1(new_n530), .B2(new_n249), .ZN(new_n531));
  NOR2_X1   g0331(.A1(new_n531), .A2(G169), .ZN(new_n532));
  AOI21_X1  g0332(.A(new_n532), .B1(new_n457), .B2(new_n531), .ZN(new_n533));
  INV_X1    g0333(.A(KEYINPUT83), .ZN(new_n534));
  INV_X1    g0334(.A(new_n440), .ZN(new_n535));
  NOR2_X1   g0335(.A1(new_n535), .A2(new_n295), .ZN(new_n536));
  INV_X1    g0336(.A(new_n536), .ZN(new_n537));
  INV_X1    g0337(.A(KEYINPUT19), .ZN(new_n538));
  NAND4_X1  g0338(.A1(new_n538), .A2(new_n206), .A3(G33), .A4(G97), .ZN(new_n539));
  NOR2_X1   g0339(.A1(G97), .A2(G107), .ZN(new_n540));
  AOI22_X1  g0340(.A1(new_n540), .A2(new_n362), .B1(new_n400), .B2(new_n206), .ZN(new_n541));
  OAI21_X1  g0341(.A(new_n539), .B1(new_n541), .B2(new_n538), .ZN(new_n542));
  NAND4_X1  g0342(.A1(new_n333), .A2(new_n206), .A3(G68), .A4(new_n253), .ZN(new_n543));
  AND2_X1   g0343(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  OAI211_X1 g0344(.A(KEYINPUT82), .B(new_n537), .C1(new_n544), .C2(new_n323), .ZN(new_n545));
  INV_X1    g0345(.A(KEYINPUT82), .ZN(new_n546));
  AOI21_X1  g0346(.A(new_n323), .B1(new_n542), .B2(new_n543), .ZN(new_n547));
  OAI21_X1  g0347(.A(new_n546), .B1(new_n547), .B2(new_n536), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n545), .A2(new_n548), .ZN(new_n549));
  NOR2_X1   g0349(.A1(new_n521), .A2(new_n440), .ZN(new_n550));
  INV_X1    g0350(.A(new_n550), .ZN(new_n551));
  AOI21_X1  g0351(.A(new_n534), .B1(new_n549), .B2(new_n551), .ZN(new_n552));
  AOI211_X1 g0352(.A(KEYINPUT83), .B(new_n550), .C1(new_n545), .C2(new_n548), .ZN(new_n553));
  OAI21_X1  g0353(.A(new_n533), .B1(new_n552), .B2(new_n553), .ZN(new_n554));
  INV_X1    g0354(.A(new_n521), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n555), .A2(G87), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n549), .A2(new_n556), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n531), .A2(G190), .ZN(new_n558));
  INV_X1    g0358(.A(G200), .ZN(new_n559));
  OAI21_X1  g0359(.A(new_n558), .B1(new_n559), .B2(new_n531), .ZN(new_n560));
  OR2_X1    g0360(.A1(new_n557), .A2(new_n560), .ZN(new_n561));
  NAND3_X1  g0361(.A1(new_n524), .A2(new_n554), .A3(new_n561), .ZN(new_n562));
  NAND2_X1  g0362(.A1(G33), .A2(G283), .ZN(new_n563));
  NAND4_X1  g0363(.A1(new_n253), .A2(new_n255), .A3(G250), .A4(G1698), .ZN(new_n564));
  NAND2_X1  g0364(.A1(KEYINPUT4), .A2(G244), .ZN(new_n565));
  OAI211_X1 g0365(.A(new_n563), .B(new_n564), .C1(new_n257), .C2(new_n565), .ZN(new_n566));
  INV_X1    g0366(.A(new_n566), .ZN(new_n567));
  NAND4_X1  g0367(.A1(new_n333), .A2(new_n359), .A3(G244), .A4(new_n253), .ZN(new_n568));
  INV_X1    g0368(.A(KEYINPUT4), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  AOI21_X1  g0370(.A(new_n272), .B1(new_n567), .B2(new_n570), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n476), .A2(new_n272), .ZN(new_n572));
  OAI21_X1  g0372(.A(new_n482), .B1(new_n572), .B2(new_n486), .ZN(new_n573));
  OAI21_X1  g0373(.A(new_n314), .B1(new_n571), .B2(new_n573), .ZN(new_n574));
  AOI21_X1  g0374(.A(new_n504), .B1(new_n349), .B2(new_n350), .ZN(new_n575));
  INV_X1    g0375(.A(KEYINPUT6), .ZN(new_n576));
  INV_X1    g0376(.A(G97), .ZN(new_n577));
  NOR3_X1   g0377(.A1(new_n576), .A2(new_n577), .A3(G107), .ZN(new_n578));
  XNOR2_X1  g0378(.A(G97), .B(G107), .ZN(new_n579));
  AOI21_X1  g0379(.A(new_n578), .B1(new_n576), .B2(new_n579), .ZN(new_n580));
  OAI22_X1  g0380(.A1(new_n580), .A2(new_n206), .B1(new_n259), .B2(new_n438), .ZN(new_n581));
  OAI21_X1  g0381(.A(new_n282), .B1(new_n575), .B2(new_n581), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n521), .A2(G97), .ZN(new_n583));
  OAI21_X1  g0383(.A(new_n583), .B1(G97), .B2(new_n296), .ZN(new_n584));
  INV_X1    g0384(.A(KEYINPUT79), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  OAI211_X1 g0386(.A(new_n583), .B(KEYINPUT79), .C1(G97), .C2(new_n296), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n582), .A2(new_n588), .ZN(new_n589));
  INV_X1    g0389(.A(new_n573), .ZN(new_n590));
  AOI21_X1  g0390(.A(new_n566), .B1(new_n569), .B2(new_n568), .ZN(new_n591));
  OAI211_X1 g0391(.A(new_n457), .B(new_n590), .C1(new_n591), .C2(new_n272), .ZN(new_n592));
  NAND3_X1  g0392(.A1(new_n574), .A2(new_n589), .A3(new_n592), .ZN(new_n593));
  INV_X1    g0393(.A(KEYINPUT81), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  NOR2_X1   g0395(.A1(new_n571), .A2(new_n573), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n596), .A2(G190), .ZN(new_n597));
  OAI21_X1  g0397(.A(new_n590), .B1(new_n591), .B2(new_n272), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n598), .A2(G200), .ZN(new_n599));
  NAND4_X1  g0399(.A1(new_n597), .A2(new_n599), .A3(new_n582), .A4(new_n588), .ZN(new_n600));
  NAND4_X1  g0400(.A1(new_n574), .A2(new_n589), .A3(new_n592), .A4(KEYINPUT81), .ZN(new_n601));
  NAND3_X1  g0401(.A1(new_n595), .A2(new_n600), .A3(new_n601), .ZN(new_n602));
  NOR2_X1   g0402(.A1(new_n562), .A2(new_n602), .ZN(new_n603));
  INV_X1    g0403(.A(KEYINPUT84), .ZN(new_n604));
  NOR3_X1   g0404(.A1(new_n358), .A2(new_n250), .A3(new_n486), .ZN(new_n605));
  NAND2_X1  g0405(.A1(G264), .A2(G1698), .ZN(new_n606));
  INV_X1    g0406(.A(new_n606), .ZN(new_n607));
  OAI211_X1 g0407(.A(new_n253), .B(new_n333), .C1(new_n605), .C2(new_n607), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n262), .A2(G303), .ZN(new_n609));
  AOI21_X1  g0409(.A(new_n272), .B1(new_n608), .B2(new_n609), .ZN(new_n610));
  NAND3_X1  g0410(.A1(new_n476), .A2(G270), .A3(new_n272), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n611), .A2(new_n482), .ZN(new_n612));
  OAI21_X1  g0412(.A(new_n604), .B1(new_n610), .B2(new_n612), .ZN(new_n613));
  AND2_X1   g0413(.A1(new_n611), .A2(new_n482), .ZN(new_n614));
  INV_X1    g0414(.A(G303), .ZN(new_n615));
  NOR2_X1   g0415(.A1(new_n260), .A2(new_n615), .ZN(new_n616));
  OAI21_X1  g0416(.A(new_n606), .B1(new_n368), .B2(new_n486), .ZN(new_n617));
  AOI21_X1  g0417(.A(new_n616), .B1(new_n341), .B2(new_n617), .ZN(new_n618));
  OAI211_X1 g0418(.A(new_n614), .B(KEYINPUT84), .C1(new_n272), .C2(new_n618), .ZN(new_n619));
  NAND3_X1  g0419(.A1(new_n613), .A2(new_n619), .A3(G200), .ZN(new_n620));
  NOR2_X1   g0420(.A1(new_n295), .A2(G116), .ZN(new_n621));
  AOI21_X1  g0421(.A(new_n621), .B1(new_n555), .B2(G116), .ZN(new_n622));
  AOI22_X1  g0422(.A1(new_n281), .A2(new_n224), .B1(G20), .B2(new_n506), .ZN(new_n623));
  OAI211_X1 g0423(.A(new_n563), .B(new_n206), .C1(G33), .C2(new_n577), .ZN(new_n624));
  AOI21_X1  g0424(.A(KEYINPUT20), .B1(new_n623), .B2(new_n624), .ZN(new_n625));
  AND3_X1   g0425(.A1(new_n623), .A2(KEYINPUT20), .A3(new_n624), .ZN(new_n626));
  OAI21_X1  g0426(.A(new_n622), .B1(new_n625), .B2(new_n626), .ZN(new_n627));
  INV_X1    g0427(.A(new_n627), .ZN(new_n628));
  NAND3_X1  g0428(.A1(new_n620), .A2(KEYINPUT87), .A3(new_n628), .ZN(new_n629));
  AND2_X1   g0429(.A1(new_n613), .A2(new_n619), .ZN(new_n630));
  OAI21_X1  g0430(.A(new_n629), .B1(new_n388), .B2(new_n630), .ZN(new_n631));
  AOI21_X1  g0431(.A(KEYINPUT87), .B1(new_n620), .B2(new_n628), .ZN(new_n632));
  NOR2_X1   g0432(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n510), .A2(new_n512), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n634), .A2(new_n282), .ZN(new_n635));
  INV_X1    g0435(.A(KEYINPUT89), .ZN(new_n636));
  INV_X1    g0436(.A(new_n519), .ZN(new_n637));
  AOI22_X1  g0437(.A1(new_n637), .A2(new_n517), .B1(G107), .B2(new_n555), .ZN(new_n638));
  NAND3_X1  g0438(.A1(new_n635), .A2(new_n636), .A3(new_n638), .ZN(new_n639));
  OAI21_X1  g0439(.A(KEYINPUT89), .B1(new_n513), .B2(new_n522), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n493), .A2(G169), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n494), .A2(G179), .ZN(new_n643));
  AOI21_X1  g0443(.A(new_n641), .B1(new_n642), .B2(new_n643), .ZN(new_n644));
  INV_X1    g0444(.A(KEYINPUT85), .ZN(new_n645));
  OR2_X1    g0445(.A1(new_n626), .A2(new_n625), .ZN(new_n646));
  AOI21_X1  g0446(.A(new_n314), .B1(new_n646), .B2(new_n622), .ZN(new_n647));
  NAND4_X1  g0447(.A1(new_n630), .A2(new_n645), .A3(KEYINPUT21), .A4(new_n647), .ZN(new_n648));
  NAND3_X1  g0448(.A1(new_n613), .A2(new_n647), .A3(new_n619), .ZN(new_n649));
  INV_X1    g0449(.A(KEYINPUT21), .ZN(new_n650));
  OAI21_X1  g0450(.A(KEYINPUT85), .B1(new_n649), .B2(new_n650), .ZN(new_n651));
  OAI211_X1 g0451(.A(new_n614), .B(G179), .C1(new_n272), .C2(new_n618), .ZN(new_n652));
  NOR2_X1   g0452(.A1(new_n652), .A2(new_n628), .ZN(new_n653));
  XNOR2_X1  g0453(.A(KEYINPUT86), .B(KEYINPUT21), .ZN(new_n654));
  AOI21_X1  g0454(.A(new_n653), .B1(new_n649), .B2(new_n654), .ZN(new_n655));
  NAND3_X1  g0455(.A1(new_n648), .A2(new_n651), .A3(new_n655), .ZN(new_n656));
  NOR3_X1   g0456(.A1(new_n633), .A2(new_n644), .A3(new_n656), .ZN(new_n657));
  AND3_X1   g0457(.A1(new_n468), .A2(new_n603), .A3(new_n657), .ZN(G372));
  NAND2_X1  g0458(.A1(new_n382), .A2(new_n384), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n365), .A2(new_n373), .ZN(new_n660));
  AND3_X1   g0460(.A1(new_n659), .A2(new_n386), .A3(new_n660), .ZN(new_n661));
  AOI21_X1  g0461(.A(new_n386), .B1(new_n659), .B2(new_n660), .ZN(new_n662));
  NOR2_X1   g0462(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  INV_X1    g0463(.A(new_n460), .ZN(new_n664));
  AOI22_X1  g0464(.A1(new_n664), .A2(new_n423), .B1(new_n431), .B2(new_n436), .ZN(new_n665));
  AND2_X1   g0465(.A1(new_n393), .A2(new_n394), .ZN(new_n666));
  INV_X1    g0466(.A(new_n666), .ZN(new_n667));
  OAI21_X1  g0467(.A(new_n663), .B1(new_n665), .B2(new_n667), .ZN(new_n668));
  AND2_X1   g0468(.A1(new_n310), .A2(new_n312), .ZN(new_n669));
  AOI22_X1  g0469(.A1(new_n668), .A2(new_n669), .B1(new_n305), .B2(new_n315), .ZN(new_n670));
  INV_X1    g0470(.A(new_n554), .ZN(new_n671));
  INV_X1    g0471(.A(KEYINPUT93), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n593), .A2(new_n672), .ZN(new_n673));
  NAND4_X1  g0473(.A1(new_n574), .A2(new_n589), .A3(new_n592), .A4(KEYINPUT93), .ZN(new_n674));
  AND4_X1   g0474(.A1(new_n554), .A2(new_n561), .A3(new_n673), .A4(new_n674), .ZN(new_n675));
  INV_X1    g0475(.A(KEYINPUT26), .ZN(new_n676));
  AOI21_X1  g0476(.A(new_n671), .B1(new_n675), .B2(new_n676), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n595), .A2(new_n601), .ZN(new_n678));
  NAND3_X1  g0478(.A1(new_n678), .A2(new_n554), .A3(new_n561), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n679), .A2(KEYINPUT26), .ZN(new_n680));
  AND3_X1   g0480(.A1(new_n595), .A2(new_n600), .A3(new_n601), .ZN(new_n681));
  NAND4_X1  g0481(.A1(new_n681), .A2(new_n554), .A3(new_n561), .A4(new_n524), .ZN(new_n682));
  AOI21_X1  g0482(.A(new_n523), .B1(new_n643), .B2(new_n642), .ZN(new_n683));
  INV_X1    g0483(.A(KEYINPUT92), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n656), .A2(new_n684), .ZN(new_n685));
  NAND4_X1  g0485(.A1(new_n648), .A2(new_n651), .A3(new_n655), .A4(KEYINPUT92), .ZN(new_n686));
  AOI21_X1  g0486(.A(new_n683), .B1(new_n685), .B2(new_n686), .ZN(new_n687));
  OAI211_X1 g0487(.A(new_n677), .B(new_n680), .C1(new_n682), .C2(new_n687), .ZN(new_n688));
  INV_X1    g0488(.A(new_n688), .ZN(new_n689));
  OAI21_X1  g0489(.A(new_n670), .B1(new_n689), .B2(new_n467), .ZN(G369));
  INV_X1    g0490(.A(G330), .ZN(new_n691));
  NOR2_X1   g0491(.A1(new_n633), .A2(new_n656), .ZN(new_n692));
  NAND3_X1  g0492(.A1(new_n205), .A2(new_n206), .A3(G13), .ZN(new_n693));
  OR2_X1    g0493(.A1(new_n693), .A2(KEYINPUT27), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n693), .A2(KEYINPUT27), .ZN(new_n695));
  NAND3_X1  g0495(.A1(new_n694), .A2(G213), .A3(new_n695), .ZN(new_n696));
  INV_X1    g0496(.A(G343), .ZN(new_n697));
  NOR2_X1   g0497(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  INV_X1    g0498(.A(new_n698), .ZN(new_n699));
  OAI21_X1  g0499(.A(new_n692), .B1(new_n628), .B2(new_n699), .ZN(new_n700));
  NAND4_X1  g0500(.A1(new_n685), .A2(new_n627), .A3(new_n686), .A4(new_n698), .ZN(new_n701));
  AOI21_X1  g0501(.A(new_n691), .B1(new_n700), .B2(new_n701), .ZN(new_n702));
  INV_X1    g0502(.A(new_n702), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n643), .A2(new_n642), .ZN(new_n704));
  NAND3_X1  g0504(.A1(new_n704), .A2(new_n640), .A3(new_n639), .ZN(new_n705));
  OAI211_X1 g0505(.A(new_n705), .B(new_n524), .C1(new_n641), .C2(new_n699), .ZN(new_n706));
  OAI21_X1  g0506(.A(new_n706), .B1(new_n705), .B2(new_n699), .ZN(new_n707));
  INV_X1    g0507(.A(new_n707), .ZN(new_n708));
  NOR2_X1   g0508(.A1(new_n703), .A2(new_n708), .ZN(new_n709));
  INV_X1    g0509(.A(new_n709), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n656), .A2(new_n699), .ZN(new_n711));
  NOR2_X1   g0511(.A1(new_n706), .A2(new_n711), .ZN(new_n712));
  INV_X1    g0512(.A(new_n712), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n683), .A2(new_n699), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  INV_X1    g0515(.A(new_n715), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n710), .A2(new_n716), .ZN(G399));
  NAND2_X1  g0517(.A1(new_n220), .A2(new_n470), .ZN(new_n718));
  NAND3_X1  g0518(.A1(new_n540), .A2(new_n362), .A3(new_n506), .ZN(new_n719));
  INV_X1    g0519(.A(new_n719), .ZN(new_n720));
  NAND3_X1  g0520(.A1(new_n718), .A2(G1), .A3(new_n720), .ZN(new_n721));
  OAI21_X1  g0521(.A(new_n721), .B1(new_n226), .B2(new_n718), .ZN(new_n722));
  XNOR2_X1  g0522(.A(new_n722), .B(KEYINPUT28), .ZN(new_n723));
  NOR2_X1   g0523(.A1(new_n644), .A2(new_n656), .ZN(new_n724));
  NOR2_X1   g0524(.A1(new_n682), .A2(new_n724), .ZN(new_n725));
  NAND4_X1  g0525(.A1(new_n678), .A2(new_n554), .A3(new_n676), .A4(new_n561), .ZN(new_n726));
  OAI211_X1 g0526(.A(new_n554), .B(new_n726), .C1(new_n675), .C2(new_n676), .ZN(new_n727));
  OAI21_X1  g0527(.A(new_n699), .B1(new_n725), .B2(new_n727), .ZN(new_n728));
  NAND2_X1  g0528(.A1(new_n728), .A2(KEYINPUT29), .ZN(new_n729));
  INV_X1    g0529(.A(KEYINPUT29), .ZN(new_n730));
  NOR2_X1   g0530(.A1(new_n687), .A2(new_n682), .ZN(new_n731));
  AND2_X1   g0531(.A1(new_n673), .A2(new_n674), .ZN(new_n732));
  NAND4_X1  g0532(.A1(new_n732), .A2(new_n676), .A3(new_n554), .A4(new_n561), .ZN(new_n733));
  NAND3_X1  g0533(.A1(new_n680), .A2(new_n733), .A3(new_n554), .ZN(new_n734));
  OAI211_X1 g0534(.A(new_n730), .B(new_n699), .C1(new_n731), .C2(new_n734), .ZN(new_n735));
  NAND2_X1  g0535(.A1(new_n729), .A2(new_n735), .ZN(new_n736));
  INV_X1    g0536(.A(new_n736), .ZN(new_n737));
  NAND2_X1  g0537(.A1(G244), .A2(G1698), .ZN(new_n738));
  INV_X1    g0538(.A(G238), .ZN(new_n739));
  OAI21_X1  g0539(.A(new_n738), .B1(new_n368), .B2(new_n739), .ZN(new_n740));
  AOI21_X1  g0540(.A(new_n507), .B1(new_n341), .B2(new_n740), .ZN(new_n741));
  OAI211_X1 g0541(.A(new_n525), .B(new_n527), .C1(new_n741), .C2(new_n272), .ZN(new_n742));
  NOR2_X1   g0542(.A1(new_n652), .A2(new_n742), .ZN(new_n743));
  NAND2_X1  g0543(.A1(new_n490), .A2(new_n491), .ZN(new_n744));
  AND2_X1   g0544(.A1(new_n483), .A2(new_n484), .ZN(new_n745));
  NAND2_X1  g0545(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  AOI22_X1  g0546(.A1(new_n746), .A2(new_n249), .B1(new_n480), .B2(new_n479), .ZN(new_n747));
  NAND3_X1  g0547(.A1(new_n743), .A2(new_n747), .A3(new_n596), .ZN(new_n748));
  INV_X1    g0548(.A(KEYINPUT30), .ZN(new_n749));
  NAND2_X1  g0549(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  NOR2_X1   g0550(.A1(new_n531), .A2(G179), .ZN(new_n751));
  NAND4_X1  g0551(.A1(new_n630), .A2(new_n598), .A3(new_n493), .A4(new_n751), .ZN(new_n752));
  NAND2_X1  g0552(.A1(new_n750), .A2(new_n752), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n753), .A2(KEYINPUT94), .ZN(new_n754));
  NAND4_X1  g0554(.A1(new_n743), .A2(new_n747), .A3(new_n596), .A4(KEYINPUT30), .ZN(new_n755));
  INV_X1    g0555(.A(KEYINPUT94), .ZN(new_n756));
  NAND3_X1  g0556(.A1(new_n750), .A2(new_n756), .A3(new_n752), .ZN(new_n757));
  NAND3_X1  g0557(.A1(new_n754), .A2(new_n755), .A3(new_n757), .ZN(new_n758));
  INV_X1    g0558(.A(KEYINPUT31), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n699), .A2(new_n759), .ZN(new_n760));
  NAND3_X1  g0560(.A1(new_n750), .A2(new_n755), .A3(new_n752), .ZN(new_n761));
  NAND2_X1  g0561(.A1(new_n761), .A2(new_n698), .ZN(new_n762));
  AOI22_X1  g0562(.A1(new_n758), .A2(new_n760), .B1(new_n759), .B2(new_n762), .ZN(new_n763));
  NAND3_X1  g0563(.A1(new_n657), .A2(new_n603), .A3(new_n699), .ZN(new_n764));
  NAND2_X1  g0564(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  NAND2_X1  g0565(.A1(new_n765), .A2(G330), .ZN(new_n766));
  NAND2_X1  g0566(.A1(new_n737), .A2(new_n766), .ZN(new_n767));
  INV_X1    g0567(.A(new_n767), .ZN(new_n768));
  OAI21_X1  g0568(.A(new_n723), .B1(new_n768), .B2(G1), .ZN(G364));
  NAND3_X1  g0569(.A1(new_n700), .A2(new_n691), .A3(new_n701), .ZN(new_n770));
  INV_X1    g0570(.A(new_n718), .ZN(new_n771));
  AND2_X1   g0571(.A1(new_n206), .A2(G13), .ZN(new_n772));
  AOI21_X1  g0572(.A(new_n205), .B1(new_n772), .B2(G45), .ZN(new_n773));
  INV_X1    g0573(.A(new_n773), .ZN(new_n774));
  OAI211_X1 g0574(.A(new_n703), .B(new_n770), .C1(new_n771), .C2(new_n774), .ZN(new_n775));
  NOR2_X1   g0575(.A1(G13), .A2(G33), .ZN(new_n776));
  INV_X1    g0576(.A(new_n776), .ZN(new_n777));
  NOR2_X1   g0577(.A1(new_n777), .A2(G20), .ZN(new_n778));
  NAND3_X1  g0578(.A1(new_n700), .A2(new_n701), .A3(new_n778), .ZN(new_n779));
  NOR2_X1   g0579(.A1(new_n771), .A2(new_n774), .ZN(new_n780));
  NAND2_X1  g0580(.A1(new_n220), .A2(new_n260), .ZN(new_n781));
  INV_X1    g0581(.A(G355), .ZN(new_n782));
  OAI22_X1  g0582(.A1(new_n781), .A2(new_n782), .B1(G116), .B2(new_n220), .ZN(new_n783));
  NAND2_X1  g0583(.A1(new_n220), .A2(new_n361), .ZN(new_n784));
  AOI21_X1  g0584(.A(new_n784), .B1(new_n474), .B2(new_n227), .ZN(new_n785));
  NAND2_X1  g0585(.A1(new_n245), .A2(G45), .ZN(new_n786));
  AOI21_X1  g0586(.A(new_n783), .B1(new_n785), .B2(new_n786), .ZN(new_n787));
  AOI21_X1  g0587(.A(new_n224), .B1(G20), .B2(new_n314), .ZN(new_n788));
  NOR2_X1   g0588(.A1(new_n778), .A2(new_n788), .ZN(new_n789));
  INV_X1    g0589(.A(new_n789), .ZN(new_n790));
  OAI21_X1  g0590(.A(new_n780), .B1(new_n787), .B2(new_n790), .ZN(new_n791));
  NOR2_X1   g0591(.A1(new_n206), .A2(G179), .ZN(new_n792));
  NAND3_X1  g0592(.A1(new_n792), .A2(new_n388), .A3(G200), .ZN(new_n793));
  NOR2_X1   g0593(.A1(new_n793), .A2(new_n504), .ZN(new_n794));
  NOR2_X1   g0594(.A1(new_n206), .A2(new_n457), .ZN(new_n795));
  NAND2_X1  g0595(.A1(new_n795), .A2(G200), .ZN(new_n796));
  NOR2_X1   g0596(.A1(new_n796), .A2(G190), .ZN(new_n797));
  INV_X1    g0597(.A(new_n797), .ZN(new_n798));
  NAND3_X1  g0598(.A1(new_n457), .A2(new_n559), .A3(G190), .ZN(new_n799));
  NAND2_X1  g0599(.A1(new_n799), .A2(G20), .ZN(new_n800));
  INV_X1    g0600(.A(new_n800), .ZN(new_n801));
  OAI22_X1  g0601(.A1(new_n798), .A2(new_n325), .B1(new_n577), .B2(new_n801), .ZN(new_n802));
  NOR2_X1   g0602(.A1(new_n796), .A2(new_n388), .ZN(new_n803));
  AOI211_X1 g0603(.A(new_n794), .B(new_n802), .C1(G50), .C2(new_n803), .ZN(new_n804));
  NOR2_X1   g0604(.A1(G190), .A2(G200), .ZN(new_n805));
  NAND2_X1  g0605(.A1(new_n792), .A2(new_n805), .ZN(new_n806));
  INV_X1    g0606(.A(new_n806), .ZN(new_n807));
  NAND2_X1  g0607(.A1(new_n807), .A2(G159), .ZN(new_n808));
  OR2_X1    g0608(.A1(new_n808), .A2(KEYINPUT32), .ZN(new_n809));
  NAND3_X1  g0609(.A1(new_n792), .A2(G190), .A3(G200), .ZN(new_n810));
  INV_X1    g0610(.A(new_n810), .ZN(new_n811));
  AOI22_X1  g0611(.A1(new_n808), .A2(KEYINPUT32), .B1(new_n811), .B2(G87), .ZN(new_n812));
  NAND2_X1  g0612(.A1(new_n795), .A2(new_n805), .ZN(new_n813));
  OAI21_X1  g0613(.A(new_n260), .B1(new_n813), .B2(new_n259), .ZN(new_n814));
  NAND3_X1  g0614(.A1(new_n795), .A2(G190), .A3(new_n559), .ZN(new_n815));
  INV_X1    g0615(.A(new_n815), .ZN(new_n816));
  AOI21_X1  g0616(.A(new_n814), .B1(G58), .B2(new_n816), .ZN(new_n817));
  NAND4_X1  g0617(.A1(new_n804), .A2(new_n809), .A3(new_n812), .A4(new_n817), .ZN(new_n818));
  INV_X1    g0618(.A(G322), .ZN(new_n819));
  NOR2_X1   g0619(.A1(new_n815), .A2(new_n819), .ZN(new_n820));
  INV_X1    g0620(.A(G311), .ZN(new_n821));
  OAI21_X1  g0621(.A(new_n262), .B1(new_n813), .B2(new_n821), .ZN(new_n822));
  AOI211_X1 g0622(.A(new_n820), .B(new_n822), .C1(G329), .C2(new_n807), .ZN(new_n823));
  NAND2_X1  g0623(.A1(new_n803), .A2(G326), .ZN(new_n824));
  XNOR2_X1  g0624(.A(KEYINPUT33), .B(G317), .ZN(new_n825));
  AOI22_X1  g0625(.A1(new_n797), .A2(new_n825), .B1(new_n811), .B2(G303), .ZN(new_n826));
  INV_X1    g0626(.A(new_n793), .ZN(new_n827));
  AOI22_X1  g0627(.A1(new_n827), .A2(G283), .B1(new_n800), .B2(G294), .ZN(new_n828));
  NAND4_X1  g0628(.A1(new_n823), .A2(new_n824), .A3(new_n826), .A4(new_n828), .ZN(new_n829));
  NAND2_X1  g0629(.A1(new_n818), .A2(new_n829), .ZN(new_n830));
  AOI21_X1  g0630(.A(new_n791), .B1(new_n830), .B2(new_n788), .ZN(new_n831));
  NAND2_X1  g0631(.A1(new_n779), .A2(new_n831), .ZN(new_n832));
  AND2_X1   g0632(.A1(new_n775), .A2(new_n832), .ZN(new_n833));
  INV_X1    g0633(.A(new_n833), .ZN(G396));
  NOR2_X1   g0634(.A1(new_n788), .A2(new_n776), .ZN(new_n835));
  INV_X1    g0635(.A(new_n835), .ZN(new_n836));
  OAI21_X1  g0636(.A(new_n780), .B1(G77), .B2(new_n836), .ZN(new_n837));
  INV_X1    g0637(.A(G283), .ZN(new_n838));
  INV_X1    g0638(.A(new_n803), .ZN(new_n839));
  OAI22_X1  g0639(.A1(new_n838), .A2(new_n798), .B1(new_n839), .B2(new_n615), .ZN(new_n840));
  AOI21_X1  g0640(.A(new_n840), .B1(G107), .B2(new_n811), .ZN(new_n841));
  INV_X1    g0641(.A(G294), .ZN(new_n842));
  OAI22_X1  g0642(.A1(new_n815), .A2(new_n842), .B1(new_n806), .B2(new_n821), .ZN(new_n843));
  INV_X1    g0643(.A(new_n813), .ZN(new_n844));
  AOI211_X1 g0644(.A(new_n260), .B(new_n843), .C1(G116), .C2(new_n844), .ZN(new_n845));
  AOI22_X1  g0645(.A1(new_n827), .A2(G87), .B1(new_n800), .B2(G97), .ZN(new_n846));
  NAND3_X1  g0646(.A1(new_n841), .A2(new_n845), .A3(new_n846), .ZN(new_n847));
  AOI22_X1  g0647(.A1(new_n816), .A2(G143), .B1(new_n844), .B2(G159), .ZN(new_n848));
  INV_X1    g0648(.A(G137), .ZN(new_n849));
  INV_X1    g0649(.A(G150), .ZN(new_n850));
  OAI221_X1 g0650(.A(new_n848), .B1(new_n839), .B2(new_n849), .C1(new_n850), .C2(new_n798), .ZN(new_n851));
  INV_X1    g0651(.A(KEYINPUT34), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  AOI21_X1  g0653(.A(new_n361), .B1(G132), .B2(new_n807), .ZN(new_n854));
  NOR2_X1   g0654(.A1(new_n810), .A2(new_n302), .ZN(new_n855));
  NOR2_X1   g0655(.A1(new_n793), .A2(new_n325), .ZN(new_n856));
  AOI211_X1 g0656(.A(new_n855), .B(new_n856), .C1(G58), .C2(new_n800), .ZN(new_n857));
  NAND3_X1  g0657(.A1(new_n853), .A2(new_n854), .A3(new_n857), .ZN(new_n858));
  NOR2_X1   g0658(.A1(new_n851), .A2(new_n852), .ZN(new_n859));
  OAI21_X1  g0659(.A(new_n847), .B1(new_n858), .B2(new_n859), .ZN(new_n860));
  AOI21_X1  g0660(.A(new_n837), .B1(new_n860), .B2(new_n788), .ZN(new_n861));
  OR2_X1    g0661(.A1(new_n445), .A2(new_n699), .ZN(new_n862));
  AOI22_X1  g0662(.A1(new_n465), .A2(new_n862), .B1(new_n458), .B2(new_n459), .ZN(new_n863));
  AND3_X1   g0663(.A1(new_n458), .A2(new_n459), .A3(new_n699), .ZN(new_n864));
  OAI21_X1  g0664(.A(KEYINPUT95), .B1(new_n863), .B2(new_n864), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n465), .A2(new_n862), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n866), .A2(new_n460), .ZN(new_n867));
  INV_X1    g0667(.A(KEYINPUT95), .ZN(new_n868));
  NAND3_X1  g0668(.A1(new_n458), .A2(new_n459), .A3(new_n699), .ZN(new_n869));
  NAND3_X1  g0669(.A1(new_n867), .A2(new_n868), .A3(new_n869), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n865), .A2(new_n870), .ZN(new_n871));
  OAI21_X1  g0671(.A(new_n861), .B1(new_n871), .B2(new_n777), .ZN(new_n872));
  XNOR2_X1  g0672(.A(new_n872), .B(KEYINPUT96), .ZN(new_n873));
  OAI211_X1 g0673(.A(new_n699), .B(new_n871), .C1(new_n731), .C2(new_n734), .ZN(new_n874));
  INV_X1    g0674(.A(KEYINPUT97), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  NAND4_X1  g0676(.A1(new_n688), .A2(KEYINPUT97), .A3(new_n699), .A4(new_n871), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  NOR3_X1   g0678(.A1(new_n863), .A2(new_n864), .A3(KEYINPUT95), .ZN(new_n879));
  AOI21_X1  g0679(.A(new_n868), .B1(new_n867), .B2(new_n869), .ZN(new_n880));
  NOR2_X1   g0680(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  OAI21_X1  g0681(.A(new_n881), .B1(new_n689), .B2(new_n698), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n878), .A2(new_n882), .ZN(new_n883));
  NOR2_X1   g0683(.A1(new_n883), .A2(new_n766), .ZN(new_n884));
  INV_X1    g0684(.A(new_n884), .ZN(new_n885));
  AOI21_X1  g0685(.A(new_n780), .B1(new_n883), .B2(new_n766), .ZN(new_n886));
  AOI21_X1  g0686(.A(new_n873), .B1(new_n885), .B2(new_n886), .ZN(new_n887));
  INV_X1    g0687(.A(new_n887), .ZN(G384));
  INV_X1    g0688(.A(new_n580), .ZN(new_n889));
  OR2_X1    g0689(.A1(new_n889), .A2(KEYINPUT35), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n889), .A2(KEYINPUT35), .ZN(new_n891));
  NAND4_X1  g0691(.A1(new_n890), .A2(G116), .A3(new_n225), .A4(new_n891), .ZN(new_n892));
  XOR2_X1   g0692(.A(new_n892), .B(KEYINPUT36), .Z(new_n893));
  OR3_X1    g0693(.A1(new_n226), .A2(new_n259), .A3(new_n326), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n302), .A2(G68), .ZN(new_n895));
  AOI211_X1 g0695(.A(new_n205), .B(G13), .C1(new_n894), .C2(new_n895), .ZN(new_n896));
  NOR2_X1   g0696(.A1(new_n893), .A2(new_n896), .ZN(new_n897));
  INV_X1    g0697(.A(new_n696), .ZN(new_n898));
  NOR2_X1   g0698(.A1(new_n663), .A2(new_n898), .ZN(new_n899));
  AND3_X1   g0699(.A1(new_n382), .A2(new_n390), .A3(new_n384), .ZN(new_n900));
  NOR2_X1   g0700(.A1(new_n900), .A2(new_n385), .ZN(new_n901));
  INV_X1    g0701(.A(KEYINPUT37), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n659), .A2(new_n898), .ZN(new_n903));
  NAND3_X1  g0703(.A1(new_n901), .A2(new_n902), .A3(new_n903), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n659), .A2(new_n660), .ZN(new_n905));
  NAND3_X1  g0705(.A1(new_n905), .A2(new_n903), .A3(new_n391), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n906), .A2(KEYINPUT37), .ZN(new_n907));
  INV_X1    g0707(.A(new_n903), .ZN(new_n908));
  AOI22_X1  g0708(.A1(new_n904), .A2(new_n907), .B1(new_n395), .B2(new_n908), .ZN(new_n909));
  OAI21_X1  g0709(.A(KEYINPUT99), .B1(new_n909), .B2(KEYINPUT38), .ZN(new_n910));
  OR2_X1    g0710(.A1(new_n343), .A2(KEYINPUT16), .ZN(new_n911));
  AOI21_X1  g0711(.A(new_n322), .B1(new_n911), .B2(new_n344), .ZN(new_n912));
  OAI21_X1  g0712(.A(new_n391), .B1(new_n912), .B2(new_n374), .ZN(new_n913));
  NOR2_X1   g0713(.A1(new_n912), .A2(new_n696), .ZN(new_n914));
  OAI21_X1  g0714(.A(KEYINPUT37), .B1(new_n913), .B2(new_n914), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n915), .A2(new_n904), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n395), .A2(new_n914), .ZN(new_n917));
  NAND3_X1  g0717(.A1(new_n916), .A2(KEYINPUT38), .A3(new_n917), .ZN(new_n918));
  INV_X1    g0718(.A(KEYINPUT99), .ZN(new_n919));
  INV_X1    g0719(.A(KEYINPUT38), .ZN(new_n920));
  AOI21_X1  g0720(.A(new_n902), .B1(new_n901), .B2(new_n903), .ZN(new_n921));
  AND4_X1   g0721(.A1(new_n902), .A2(new_n905), .A3(new_n903), .A4(new_n391), .ZN(new_n922));
  NOR2_X1   g0722(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  AOI21_X1  g0723(.A(new_n903), .B1(new_n663), .B2(new_n666), .ZN(new_n924));
  OAI211_X1 g0724(.A(new_n919), .B(new_n920), .C1(new_n923), .C2(new_n924), .ZN(new_n925));
  NAND3_X1  g0725(.A1(new_n910), .A2(new_n918), .A3(new_n925), .ZN(new_n926));
  INV_X1    g0726(.A(KEYINPUT39), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  AND3_X1   g0728(.A1(new_n916), .A2(KEYINPUT38), .A3(new_n917), .ZN(new_n929));
  AOI21_X1  g0729(.A(KEYINPUT38), .B1(new_n916), .B2(new_n917), .ZN(new_n930));
  OR2_X1    g0730(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  OAI21_X1  g0731(.A(new_n928), .B1(new_n927), .B2(new_n931), .ZN(new_n932));
  INV_X1    g0732(.A(new_n932), .ZN(new_n933));
  NAND3_X1  g0733(.A1(new_n431), .A2(new_n436), .A3(new_n699), .ZN(new_n934));
  INV_X1    g0734(.A(new_n934), .ZN(new_n935));
  AOI21_X1  g0735(.A(new_n899), .B1(new_n933), .B2(new_n935), .ZN(new_n936));
  AOI21_X1  g0736(.A(new_n864), .B1(new_n876), .B2(new_n877), .ZN(new_n937));
  AND2_X1   g0737(.A1(new_n425), .A2(new_n427), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n430), .A2(new_n429), .ZN(new_n939));
  OAI21_X1  g0739(.A(new_n436), .B1(new_n938), .B2(new_n939), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n436), .A2(new_n698), .ZN(new_n941));
  NAND3_X1  g0741(.A1(new_n940), .A2(new_n423), .A3(new_n941), .ZN(new_n942));
  OAI211_X1 g0742(.A(new_n436), .B(new_n698), .C1(new_n431), .C2(new_n424), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  INV_X1    g0744(.A(new_n944), .ZN(new_n945));
  OAI21_X1  g0745(.A(KEYINPUT98), .B1(new_n937), .B2(new_n945), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n946), .A2(new_n931), .ZN(new_n947));
  NOR3_X1   g0747(.A1(new_n937), .A2(KEYINPUT98), .A3(new_n945), .ZN(new_n948));
  OAI21_X1  g0748(.A(new_n936), .B1(new_n947), .B2(new_n948), .ZN(new_n949));
  INV_X1    g0749(.A(KEYINPUT100), .ZN(new_n950));
  AOI21_X1  g0750(.A(new_n950), .B1(new_n736), .B2(new_n468), .ZN(new_n951));
  AOI211_X1 g0751(.A(KEYINPUT100), .B(new_n467), .C1(new_n729), .C2(new_n735), .ZN(new_n952));
  OAI21_X1  g0752(.A(new_n670), .B1(new_n951), .B2(new_n952), .ZN(new_n953));
  XNOR2_X1  g0753(.A(new_n949), .B(new_n953), .ZN(new_n954));
  OAI21_X1  g0754(.A(new_n944), .B1(new_n879), .B2(new_n880), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n761), .A2(new_n760), .ZN(new_n956));
  INV_X1    g0756(.A(new_n956), .ZN(new_n957));
  AOI21_X1  g0757(.A(KEYINPUT31), .B1(new_n762), .B2(KEYINPUT101), .ZN(new_n958));
  INV_X1    g0758(.A(KEYINPUT101), .ZN(new_n959));
  NAND3_X1  g0759(.A1(new_n761), .A2(new_n959), .A3(new_n698), .ZN(new_n960));
  AOI21_X1  g0760(.A(new_n957), .B1(new_n958), .B2(new_n960), .ZN(new_n961));
  AOI21_X1  g0761(.A(new_n955), .B1(new_n961), .B2(new_n764), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n926), .A2(new_n962), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n963), .A2(KEYINPUT40), .ZN(new_n964));
  INV_X1    g0764(.A(KEYINPUT40), .ZN(new_n965));
  NAND3_X1  g0765(.A1(new_n931), .A2(new_n962), .A3(new_n965), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n964), .A2(new_n966), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n762), .A2(KEYINPUT101), .ZN(new_n968));
  NAND3_X1  g0768(.A1(new_n968), .A2(new_n759), .A3(new_n960), .ZN(new_n969));
  NAND3_X1  g0769(.A1(new_n764), .A2(new_n956), .A3(new_n969), .ZN(new_n970));
  NAND3_X1  g0770(.A1(new_n967), .A2(new_n468), .A3(new_n970), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n468), .A2(new_n970), .ZN(new_n972));
  NAND3_X1  g0772(.A1(new_n964), .A2(new_n972), .A3(new_n966), .ZN(new_n973));
  NAND3_X1  g0773(.A1(new_n971), .A2(G330), .A3(new_n973), .ZN(new_n974));
  AND2_X1   g0774(.A1(new_n954), .A2(new_n974), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n975), .A2(KEYINPUT102), .ZN(new_n976));
  OAI221_X1 g0776(.A(new_n976), .B1(new_n205), .B2(new_n772), .C1(new_n954), .C2(new_n974), .ZN(new_n977));
  NOR2_X1   g0777(.A1(new_n975), .A2(KEYINPUT102), .ZN(new_n978));
  OAI21_X1  g0778(.A(new_n897), .B1(new_n977), .B2(new_n978), .ZN(G367));
  NAND2_X1  g0779(.A1(new_n557), .A2(new_n698), .ZN(new_n980));
  XOR2_X1   g0780(.A(new_n980), .B(KEYINPUT103), .Z(new_n981));
  NAND2_X1  g0781(.A1(new_n554), .A2(new_n561), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n981), .A2(new_n982), .ZN(new_n983));
  OAI21_X1  g0783(.A(new_n983), .B1(new_n671), .B2(new_n981), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n984), .A2(new_n778), .ZN(new_n985));
  INV_X1    g0785(.A(G159), .ZN(new_n986));
  OAI22_X1  g0786(.A1(new_n798), .A2(new_n986), .B1(new_n810), .B2(new_n324), .ZN(new_n987));
  AOI21_X1  g0787(.A(new_n987), .B1(G68), .B2(new_n800), .ZN(new_n988));
  OAI22_X1  g0788(.A1(new_n815), .A2(new_n850), .B1(new_n806), .B2(new_n849), .ZN(new_n989));
  AOI211_X1 g0789(.A(new_n262), .B(new_n989), .C1(G50), .C2(new_n844), .ZN(new_n990));
  AOI22_X1  g0790(.A1(new_n803), .A2(G143), .B1(new_n827), .B2(G77), .ZN(new_n991));
  NAND3_X1  g0791(.A1(new_n988), .A2(new_n990), .A3(new_n991), .ZN(new_n992));
  OAI22_X1  g0792(.A1(new_n801), .A2(new_n504), .B1(new_n793), .B2(new_n577), .ZN(new_n993));
  AOI21_X1  g0793(.A(new_n993), .B1(G311), .B2(new_n803), .ZN(new_n994));
  NAND3_X1  g0794(.A1(new_n811), .A2(KEYINPUT46), .A3(G116), .ZN(new_n995));
  INV_X1    g0795(.A(G317), .ZN(new_n996));
  OAI22_X1  g0796(.A1(new_n815), .A2(new_n615), .B1(new_n806), .B2(new_n996), .ZN(new_n997));
  AOI21_X1  g0797(.A(new_n997), .B1(G283), .B2(new_n844), .ZN(new_n998));
  AOI21_X1  g0798(.A(new_n341), .B1(G294), .B2(new_n797), .ZN(new_n999));
  NAND4_X1  g0799(.A1(new_n994), .A2(new_n995), .A3(new_n998), .A4(new_n999), .ZN(new_n1000));
  AOI21_X1  g0800(.A(KEYINPUT46), .B1(new_n811), .B2(G116), .ZN(new_n1001));
  XNOR2_X1  g0801(.A(new_n1001), .B(KEYINPUT110), .ZN(new_n1002));
  OAI21_X1  g0802(.A(new_n992), .B1(new_n1000), .B2(new_n1002), .ZN(new_n1003));
  XNOR2_X1  g0803(.A(new_n1003), .B(KEYINPUT47), .ZN(new_n1004));
  NAND2_X1  g0804(.A1(new_n1004), .A2(new_n788), .ZN(new_n1005));
  OAI221_X1 g0805(.A(new_n789), .B1(new_n220), .B2(new_n440), .C1(new_n237), .C2(new_n784), .ZN(new_n1006));
  NAND4_X1  g0806(.A1(new_n985), .A2(new_n780), .A3(new_n1005), .A4(new_n1006), .ZN(new_n1007));
  XOR2_X1   g0807(.A(KEYINPUT106), .B(KEYINPUT44), .Z(new_n1008));
  INV_X1    g0808(.A(new_n1008), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n589), .A2(new_n698), .ZN(new_n1010));
  NAND2_X1  g0810(.A1(new_n681), .A2(new_n1010), .ZN(new_n1011));
  OAI22_X1  g0811(.A1(new_n1011), .A2(KEYINPUT104), .B1(new_n593), .B2(new_n699), .ZN(new_n1012));
  AND2_X1   g0812(.A1(new_n1011), .A2(KEYINPUT104), .ZN(new_n1013));
  NOR2_X1   g0813(.A1(new_n1012), .A2(new_n1013), .ZN(new_n1014));
  INV_X1    g0814(.A(new_n1014), .ZN(new_n1015));
  OAI21_X1  g0815(.A(new_n1009), .B1(new_n716), .B2(new_n1015), .ZN(new_n1016));
  NAND3_X1  g0816(.A1(new_n715), .A2(new_n1014), .A3(new_n1008), .ZN(new_n1017));
  AND2_X1   g0817(.A1(new_n1016), .A2(new_n1017), .ZN(new_n1018));
  NAND3_X1  g0818(.A1(new_n716), .A2(KEYINPUT45), .A3(new_n1015), .ZN(new_n1019));
  INV_X1    g0819(.A(KEYINPUT45), .ZN(new_n1020));
  OAI21_X1  g0820(.A(new_n1020), .B1(new_n715), .B2(new_n1014), .ZN(new_n1021));
  NAND2_X1  g0821(.A1(new_n1019), .A2(new_n1021), .ZN(new_n1022));
  NAND4_X1  g0822(.A1(new_n1018), .A2(KEYINPUT107), .A3(new_n709), .A4(new_n1022), .ZN(new_n1023));
  NAND2_X1  g0823(.A1(new_n709), .A2(KEYINPUT107), .ZN(new_n1024));
  INV_X1    g0824(.A(new_n1022), .ZN(new_n1025));
  NAND2_X1  g0825(.A1(new_n1016), .A2(new_n1017), .ZN(new_n1026));
  OAI21_X1  g0826(.A(new_n1024), .B1(new_n1025), .B2(new_n1026), .ZN(new_n1027));
  NAND2_X1  g0827(.A1(new_n1023), .A2(new_n1027), .ZN(new_n1028));
  NAND2_X1  g0828(.A1(new_n708), .A2(new_n711), .ZN(new_n1029));
  NAND2_X1  g0829(.A1(new_n1029), .A2(new_n713), .ZN(new_n1030));
  XNOR2_X1  g0830(.A(new_n1030), .B(new_n702), .ZN(new_n1031));
  NAND3_X1  g0831(.A1(new_n1031), .A2(new_n737), .A3(new_n766), .ZN(new_n1032));
  NAND2_X1  g0832(.A1(new_n1032), .A2(KEYINPUT108), .ZN(new_n1033));
  XNOR2_X1  g0833(.A(new_n1030), .B(new_n703), .ZN(new_n1034));
  NOR2_X1   g0834(.A1(new_n1034), .A2(new_n767), .ZN(new_n1035));
  INV_X1    g0835(.A(KEYINPUT108), .ZN(new_n1036));
  NAND2_X1  g0836(.A1(new_n1035), .A2(new_n1036), .ZN(new_n1037));
  AND4_X1   g0837(.A1(KEYINPUT109), .A2(new_n1028), .A3(new_n1033), .A4(new_n1037), .ZN(new_n1038));
  AOI22_X1  g0838(.A1(new_n1023), .A2(new_n1027), .B1(new_n1032), .B2(KEYINPUT108), .ZN(new_n1039));
  AOI21_X1  g0839(.A(KEYINPUT109), .B1(new_n1039), .B2(new_n1037), .ZN(new_n1040));
  OAI21_X1  g0840(.A(new_n768), .B1(new_n1038), .B2(new_n1040), .ZN(new_n1041));
  XNOR2_X1  g0841(.A(new_n718), .B(KEYINPUT41), .ZN(new_n1042));
  INV_X1    g0842(.A(new_n1042), .ZN(new_n1043));
  AOI21_X1  g0843(.A(new_n774), .B1(new_n1041), .B2(new_n1043), .ZN(new_n1044));
  NAND2_X1  g0844(.A1(new_n1015), .A2(new_n712), .ZN(new_n1045));
  XNOR2_X1  g0845(.A(new_n1045), .B(KEYINPUT42), .ZN(new_n1046));
  AOI21_X1  g0846(.A(new_n678), .B1(new_n1015), .B2(new_n644), .ZN(new_n1047));
  NOR2_X1   g0847(.A1(new_n1047), .A2(new_n698), .ZN(new_n1048));
  INV_X1    g0848(.A(KEYINPUT43), .ZN(new_n1049));
  OAI22_X1  g0849(.A1(new_n1046), .A2(new_n1048), .B1(new_n1049), .B2(new_n984), .ZN(new_n1050));
  NAND2_X1  g0850(.A1(new_n984), .A2(new_n1049), .ZN(new_n1051));
  INV_X1    g0851(.A(new_n1051), .ZN(new_n1052));
  XNOR2_X1  g0852(.A(new_n1050), .B(new_n1052), .ZN(new_n1053));
  NOR2_X1   g0853(.A1(new_n710), .A2(new_n1014), .ZN(new_n1054));
  INV_X1    g0854(.A(new_n1054), .ZN(new_n1055));
  OAI21_X1  g0855(.A(KEYINPUT105), .B1(new_n1053), .B2(new_n1055), .ZN(new_n1056));
  XNOR2_X1  g0856(.A(new_n1050), .B(new_n1051), .ZN(new_n1057));
  INV_X1    g0857(.A(KEYINPUT105), .ZN(new_n1058));
  NAND3_X1  g0858(.A1(new_n1057), .A2(new_n1058), .A3(new_n1054), .ZN(new_n1059));
  NAND2_X1  g0859(.A1(new_n1053), .A2(new_n1055), .ZN(new_n1060));
  NAND3_X1  g0860(.A1(new_n1056), .A2(new_n1059), .A3(new_n1060), .ZN(new_n1061));
  OAI21_X1  g0861(.A(new_n1007), .B1(new_n1044), .B2(new_n1061), .ZN(G387));
  NAND2_X1  g0862(.A1(new_n1034), .A2(new_n767), .ZN(new_n1063));
  NAND3_X1  g0863(.A1(new_n1032), .A2(new_n771), .A3(new_n1063), .ZN(new_n1064));
  NAND2_X1  g0864(.A1(new_n708), .A2(new_n778), .ZN(new_n1065));
  OAI22_X1  g0865(.A1(new_n781), .A2(new_n720), .B1(G107), .B2(new_n220), .ZN(new_n1066));
  OR2_X1    g0866(.A1(new_n234), .A2(new_n474), .ZN(new_n1067));
  NOR2_X1   g0867(.A1(new_n283), .A2(G50), .ZN(new_n1068));
  XNOR2_X1  g0868(.A(new_n1068), .B(KEYINPUT50), .ZN(new_n1069));
  AOI211_X1 g0869(.A(G45), .B(new_n719), .C1(G68), .C2(G77), .ZN(new_n1070));
  AOI21_X1  g0870(.A(new_n784), .B1(new_n1069), .B2(new_n1070), .ZN(new_n1071));
  AOI21_X1  g0871(.A(new_n1066), .B1(new_n1067), .B2(new_n1071), .ZN(new_n1072));
  OAI21_X1  g0872(.A(new_n780), .B1(new_n1072), .B2(new_n790), .ZN(new_n1073));
  XOR2_X1   g0873(.A(new_n1073), .B(KEYINPUT111), .Z(new_n1074));
  OAI22_X1  g0874(.A1(new_n259), .A2(new_n810), .B1(new_n793), .B2(new_n577), .ZN(new_n1075));
  XNOR2_X1  g0875(.A(KEYINPUT112), .B(G150), .ZN(new_n1076));
  AOI211_X1 g0876(.A(new_n361), .B(new_n1075), .C1(new_n807), .C2(new_n1076), .ZN(new_n1077));
  XNOR2_X1  g0877(.A(new_n1077), .B(KEYINPUT113), .ZN(new_n1078));
  AOI22_X1  g0878(.A1(new_n816), .A2(G50), .B1(new_n844), .B2(G68), .ZN(new_n1079));
  NAND2_X1  g0879(.A1(new_n535), .A2(new_n800), .ZN(new_n1080));
  OAI211_X1 g0880(.A(new_n1079), .B(new_n1080), .C1(new_n986), .C2(new_n839), .ZN(new_n1081));
  AOI21_X1  g0881(.A(new_n1081), .B1(new_n320), .B2(new_n797), .ZN(new_n1082));
  NAND2_X1  g0882(.A1(new_n1078), .A2(new_n1082), .ZN(new_n1083));
  AOI21_X1  g0883(.A(new_n341), .B1(G326), .B2(new_n807), .ZN(new_n1084));
  OAI22_X1  g0884(.A1(new_n801), .A2(new_n838), .B1(new_n810), .B2(new_n842), .ZN(new_n1085));
  AOI22_X1  g0885(.A1(new_n816), .A2(G317), .B1(new_n844), .B2(G303), .ZN(new_n1086));
  OAI221_X1 g0886(.A(new_n1086), .B1(new_n839), .B2(new_n819), .C1(new_n821), .C2(new_n798), .ZN(new_n1087));
  INV_X1    g0887(.A(KEYINPUT48), .ZN(new_n1088));
  AOI21_X1  g0888(.A(new_n1085), .B1(new_n1087), .B2(new_n1088), .ZN(new_n1089));
  OAI21_X1  g0889(.A(new_n1089), .B1(new_n1088), .B2(new_n1087), .ZN(new_n1090));
  INV_X1    g0890(.A(KEYINPUT49), .ZN(new_n1091));
  OAI221_X1 g0891(.A(new_n1084), .B1(new_n506), .B2(new_n793), .C1(new_n1090), .C2(new_n1091), .ZN(new_n1092));
  AND2_X1   g0892(.A1(new_n1090), .A2(new_n1091), .ZN(new_n1093));
  OAI21_X1  g0893(.A(new_n1083), .B1(new_n1092), .B2(new_n1093), .ZN(new_n1094));
  AOI21_X1  g0894(.A(new_n1074), .B1(new_n788), .B2(new_n1094), .ZN(new_n1095));
  AOI22_X1  g0895(.A1(new_n1031), .A2(new_n774), .B1(new_n1065), .B2(new_n1095), .ZN(new_n1096));
  NAND2_X1  g0896(.A1(new_n1064), .A2(new_n1096), .ZN(G393));
  NAND2_X1  g0897(.A1(new_n1018), .A2(new_n1022), .ZN(new_n1098));
  XNOR2_X1  g0898(.A(new_n1098), .B(new_n710), .ZN(new_n1099));
  OAI21_X1  g0899(.A(new_n771), .B1(new_n1099), .B2(new_n1035), .ZN(new_n1100));
  NAND3_X1  g0900(.A1(new_n1028), .A2(new_n1033), .A3(new_n1037), .ZN(new_n1101));
  INV_X1    g0901(.A(KEYINPUT109), .ZN(new_n1102));
  NAND2_X1  g0902(.A1(new_n1101), .A2(new_n1102), .ZN(new_n1103));
  NAND3_X1  g0903(.A1(new_n1039), .A2(KEYINPUT109), .A3(new_n1037), .ZN(new_n1104));
  AOI21_X1  g0904(.A(new_n1100), .B1(new_n1103), .B2(new_n1104), .ZN(new_n1105));
  NAND2_X1  g0905(.A1(new_n1099), .A2(new_n774), .ZN(new_n1106));
  NAND2_X1  g0906(.A1(new_n1014), .A2(new_n778), .ZN(new_n1107));
  AOI22_X1  g0907(.A1(G150), .A2(new_n803), .B1(new_n816), .B2(G159), .ZN(new_n1108));
  XNOR2_X1  g0908(.A(KEYINPUT114), .B(KEYINPUT51), .ZN(new_n1109));
  XNOR2_X1  g0909(.A(new_n1108), .B(new_n1109), .ZN(new_n1110));
  NOR2_X1   g0910(.A1(new_n813), .A2(new_n283), .ZN(new_n1111));
  AOI211_X1 g0911(.A(new_n361), .B(new_n1111), .C1(G143), .C2(new_n807), .ZN(new_n1112));
  NOR2_X1   g0912(.A1(new_n801), .A2(new_n259), .ZN(new_n1113));
  OAI22_X1  g0913(.A1(new_n325), .A2(new_n810), .B1(new_n793), .B2(new_n362), .ZN(new_n1114));
  AOI211_X1 g0914(.A(new_n1113), .B(new_n1114), .C1(G50), .C2(new_n797), .ZN(new_n1115));
  NAND3_X1  g0915(.A1(new_n1110), .A2(new_n1112), .A3(new_n1115), .ZN(new_n1116));
  OAI22_X1  g0916(.A1(new_n839), .A2(new_n996), .B1(new_n821), .B2(new_n815), .ZN(new_n1117));
  XNOR2_X1  g0917(.A(new_n1117), .B(KEYINPUT52), .ZN(new_n1118));
  OAI22_X1  g0918(.A1(new_n810), .A2(new_n838), .B1(new_n806), .B2(new_n819), .ZN(new_n1119));
  INV_X1    g0919(.A(KEYINPUT115), .ZN(new_n1120));
  AOI211_X1 g0920(.A(new_n260), .B(new_n794), .C1(new_n1119), .C2(new_n1120), .ZN(new_n1121));
  OAI211_X1 g0921(.A(new_n1118), .B(new_n1121), .C1(new_n1120), .C2(new_n1119), .ZN(new_n1122));
  AOI22_X1  g0922(.A1(new_n844), .A2(G294), .B1(G116), .B2(new_n800), .ZN(new_n1123));
  OAI21_X1  g0923(.A(new_n1123), .B1(new_n615), .B2(new_n798), .ZN(new_n1124));
  XNOR2_X1  g0924(.A(new_n1124), .B(KEYINPUT116), .ZN(new_n1125));
  OAI21_X1  g0925(.A(new_n1116), .B1(new_n1122), .B2(new_n1125), .ZN(new_n1126));
  NAND2_X1  g0926(.A1(new_n1126), .A2(new_n788), .ZN(new_n1127));
  INV_X1    g0927(.A(new_n242), .ZN(new_n1128));
  OAI221_X1 g0928(.A(new_n789), .B1(new_n577), .B2(new_n220), .C1(new_n1128), .C2(new_n784), .ZN(new_n1129));
  NAND4_X1  g0929(.A1(new_n1107), .A2(new_n780), .A3(new_n1127), .A4(new_n1129), .ZN(new_n1130));
  NAND2_X1  g0930(.A1(new_n1106), .A2(new_n1130), .ZN(new_n1131));
  NOR2_X1   g0931(.A1(new_n1105), .A2(new_n1131), .ZN(new_n1132));
  INV_X1    g0932(.A(new_n1132), .ZN(G390));
  AOI211_X1 g0933(.A(new_n774), .B(new_n771), .C1(new_n284), .C2(new_n835), .ZN(new_n1134));
  INV_X1    g0934(.A(new_n788), .ZN(new_n1135));
  AOI22_X1  g0935(.A1(G97), .A2(new_n844), .B1(new_n807), .B2(G294), .ZN(new_n1136));
  OAI211_X1 g0936(.A(new_n1136), .B(new_n262), .C1(new_n506), .C2(new_n815), .ZN(new_n1137));
  AOI211_X1 g0937(.A(new_n856), .B(new_n1137), .C1(G87), .C2(new_n811), .ZN(new_n1138));
  NOR2_X1   g0938(.A1(new_n798), .A2(new_n504), .ZN(new_n1139));
  AOI211_X1 g0939(.A(new_n1113), .B(new_n1139), .C1(G283), .C2(new_n803), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n811), .A2(new_n1076), .ZN(new_n1141));
  XOR2_X1   g0941(.A(new_n1141), .B(KEYINPUT53), .Z(new_n1142));
  OAI22_X1  g0942(.A1(new_n798), .A2(new_n849), .B1(new_n793), .B2(new_n302), .ZN(new_n1143));
  INV_X1    g0943(.A(G128), .ZN(new_n1144));
  OAI22_X1  g0944(.A1(new_n839), .A2(new_n1144), .B1(new_n986), .B2(new_n801), .ZN(new_n1145));
  INV_X1    g0945(.A(G125), .ZN(new_n1146));
  OAI21_X1  g0946(.A(new_n260), .B1(new_n806), .B2(new_n1146), .ZN(new_n1147));
  INV_X1    g0947(.A(G132), .ZN(new_n1148));
  XNOR2_X1  g0948(.A(KEYINPUT54), .B(G143), .ZN(new_n1149));
  OAI22_X1  g0949(.A1(new_n815), .A2(new_n1148), .B1(new_n813), .B2(new_n1149), .ZN(new_n1150));
  NOR4_X1   g0950(.A1(new_n1143), .A2(new_n1145), .A3(new_n1147), .A4(new_n1150), .ZN(new_n1151));
  AOI22_X1  g0951(.A1(new_n1138), .A2(new_n1140), .B1(new_n1142), .B2(new_n1151), .ZN(new_n1152));
  OAI221_X1 g0952(.A(new_n1134), .B1(new_n1135), .B2(new_n1152), .C1(new_n933), .C2(new_n777), .ZN(new_n1153));
  OAI21_X1  g0953(.A(new_n934), .B1(new_n937), .B2(new_n945), .ZN(new_n1154));
  NAND2_X1  g0954(.A1(new_n1154), .A2(new_n932), .ZN(new_n1155));
  OAI211_X1 g0955(.A(new_n699), .B(new_n871), .C1(new_n725), .C2(new_n727), .ZN(new_n1156));
  AND2_X1   g0956(.A1(new_n1156), .A2(new_n869), .ZN(new_n1157));
  NOR2_X1   g0957(.A1(new_n1157), .A2(new_n945), .ZN(new_n1158));
  NAND2_X1  g0958(.A1(new_n926), .A2(new_n934), .ZN(new_n1159));
  NOR2_X1   g0959(.A1(new_n1158), .A2(new_n1159), .ZN(new_n1160));
  INV_X1    g0960(.A(new_n1160), .ZN(new_n1161));
  NAND4_X1  g0961(.A1(new_n765), .A2(G330), .A3(new_n871), .A4(new_n944), .ZN(new_n1162));
  NAND3_X1  g0962(.A1(new_n1155), .A2(new_n1161), .A3(new_n1162), .ZN(new_n1163));
  AOI21_X1  g0963(.A(new_n1160), .B1(new_n1154), .B2(new_n932), .ZN(new_n1164));
  AOI21_X1  g0964(.A(new_n691), .B1(new_n961), .B2(new_n764), .ZN(new_n1165));
  INV_X1    g0965(.A(new_n955), .ZN(new_n1166));
  NAND2_X1  g0966(.A1(new_n1165), .A2(new_n1166), .ZN(new_n1167));
  OAI21_X1  g0967(.A(new_n1163), .B1(new_n1164), .B2(new_n1167), .ZN(new_n1168));
  OAI21_X1  g0968(.A(new_n1153), .B1(new_n1168), .B2(new_n773), .ZN(new_n1169));
  INV_X1    g0969(.A(KEYINPUT117), .ZN(new_n1170));
  NAND3_X1  g0970(.A1(new_n1162), .A2(new_n869), .A3(new_n1156), .ZN(new_n1171));
  AOI21_X1  g0971(.A(new_n944), .B1(new_n1165), .B2(new_n871), .ZN(new_n1172));
  OAI21_X1  g0972(.A(new_n1170), .B1(new_n1171), .B2(new_n1172), .ZN(new_n1173));
  NAND3_X1  g0973(.A1(new_n970), .A2(G330), .A3(new_n871), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n1174), .A2(new_n945), .ZN(new_n1175));
  NAND4_X1  g0975(.A1(new_n1175), .A2(new_n1157), .A3(KEYINPUT117), .A4(new_n1162), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n878), .A2(new_n869), .ZN(new_n1177));
  OAI21_X1  g0977(.A(new_n945), .B1(new_n766), .B2(new_n881), .ZN(new_n1178));
  NAND2_X1  g0978(.A1(new_n1178), .A2(new_n1167), .ZN(new_n1179));
  AOI22_X1  g0979(.A1(new_n1173), .A2(new_n1176), .B1(new_n1177), .B2(new_n1179), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n468), .A2(new_n1165), .ZN(new_n1181));
  OAI211_X1 g0981(.A(new_n670), .B(new_n1181), .C1(new_n951), .C2(new_n952), .ZN(new_n1182));
  NOR2_X1   g0982(.A1(new_n1180), .A2(new_n1182), .ZN(new_n1183));
  INV_X1    g0983(.A(new_n1183), .ZN(new_n1184));
  AOI21_X1  g0984(.A(new_n718), .B1(new_n1168), .B2(new_n1184), .ZN(new_n1185));
  OAI211_X1 g0985(.A(new_n1183), .B(new_n1163), .C1(new_n1164), .C2(new_n1167), .ZN(new_n1186));
  AOI21_X1  g0986(.A(new_n1169), .B1(new_n1185), .B2(new_n1186), .ZN(new_n1187));
  INV_X1    g0987(.A(new_n1187), .ZN(G378));
  NAND2_X1  g0988(.A1(new_n305), .A2(new_n898), .ZN(new_n1189));
  XOR2_X1   g0989(.A(new_n1189), .B(KEYINPUT55), .Z(new_n1190));
  INV_X1    g0990(.A(new_n1190), .ZN(new_n1191));
  NAND3_X1  g0991(.A1(new_n669), .A2(new_n316), .A3(new_n1191), .ZN(new_n1192));
  XOR2_X1   g0992(.A(KEYINPUT119), .B(KEYINPUT56), .Z(new_n1193));
  NAND2_X1  g0993(.A1(new_n317), .A2(new_n1190), .ZN(new_n1194));
  AND3_X1   g0994(.A1(new_n1192), .A2(new_n1193), .A3(new_n1194), .ZN(new_n1195));
  AOI21_X1  g0995(.A(new_n1193), .B1(new_n1192), .B2(new_n1194), .ZN(new_n1196));
  NOR2_X1   g0996(.A1(new_n1195), .A2(new_n1196), .ZN(new_n1197));
  AOI21_X1  g0997(.A(new_n1197), .B1(new_n967), .B2(G330), .ZN(new_n1198));
  AOI21_X1  g0998(.A(new_n965), .B1(new_n926), .B2(new_n962), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n970), .A2(new_n1166), .ZN(new_n1200));
  OAI21_X1  g1000(.A(new_n965), .B1(new_n929), .B2(new_n930), .ZN(new_n1201));
  NOR2_X1   g1001(.A1(new_n1200), .A2(new_n1201), .ZN(new_n1202));
  OAI211_X1 g1002(.A(G330), .B(new_n1197), .C1(new_n1199), .C2(new_n1202), .ZN(new_n1203));
  INV_X1    g1003(.A(new_n1203), .ZN(new_n1204));
  OAI21_X1  g1004(.A(KEYINPUT120), .B1(new_n1198), .B2(new_n1204), .ZN(new_n1205));
  OAI21_X1  g1005(.A(G330), .B1(new_n1199), .B2(new_n1202), .ZN(new_n1206));
  OAI21_X1  g1006(.A(new_n1206), .B1(new_n1195), .B2(new_n1196), .ZN(new_n1207));
  INV_X1    g1007(.A(KEYINPUT120), .ZN(new_n1208));
  NAND3_X1  g1008(.A1(new_n1207), .A2(new_n1208), .A3(new_n1203), .ZN(new_n1209));
  NAND3_X1  g1009(.A1(new_n949), .A2(new_n1205), .A3(new_n1209), .ZN(new_n1210));
  INV_X1    g1010(.A(KEYINPUT98), .ZN(new_n1211));
  NAND3_X1  g1011(.A1(new_n1177), .A2(new_n1211), .A3(new_n944), .ZN(new_n1212));
  NAND3_X1  g1012(.A1(new_n1212), .A2(new_n931), .A3(new_n946), .ZN(new_n1213));
  NAND4_X1  g1013(.A1(new_n1213), .A2(new_n936), .A3(new_n1203), .A4(new_n1207), .ZN(new_n1214));
  NAND2_X1  g1014(.A1(new_n1210), .A2(new_n1214), .ZN(new_n1215));
  NAND2_X1  g1015(.A1(new_n1215), .A2(new_n774), .ZN(new_n1216));
  INV_X1    g1016(.A(KEYINPUT121), .ZN(new_n1217));
  NOR2_X1   g1017(.A1(new_n1197), .A2(new_n777), .ZN(new_n1218));
  NOR2_X1   g1018(.A1(new_n341), .A2(G41), .ZN(new_n1219));
  AOI211_X1 g1019(.A(G50), .B(new_n1219), .C1(new_n252), .C2(new_n470), .ZN(new_n1220));
  AOI22_X1  g1020(.A1(new_n816), .A2(G107), .B1(new_n844), .B2(new_n535), .ZN(new_n1221));
  OAI21_X1  g1021(.A(new_n1221), .B1(new_n838), .B2(new_n806), .ZN(new_n1222));
  OAI22_X1  g1022(.A1(new_n577), .A2(new_n798), .B1(new_n839), .B2(new_n506), .ZN(new_n1223));
  OAI22_X1  g1023(.A1(new_n801), .A2(new_n325), .B1(new_n810), .B2(new_n259), .ZN(new_n1224));
  INV_X1    g1024(.A(new_n1219), .ZN(new_n1225));
  NOR4_X1   g1025(.A1(new_n1222), .A2(new_n1223), .A3(new_n1224), .A4(new_n1225), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n827), .A2(G58), .ZN(new_n1227));
  XNOR2_X1  g1027(.A(new_n1227), .B(KEYINPUT118), .ZN(new_n1228));
  AND2_X1   g1028(.A1(new_n1226), .A2(new_n1228), .ZN(new_n1229));
  AOI21_X1  g1029(.A(new_n1220), .B1(new_n1229), .B2(KEYINPUT58), .ZN(new_n1230));
  OAI22_X1  g1030(.A1(new_n1146), .A2(new_n839), .B1(new_n798), .B2(new_n1148), .ZN(new_n1231));
  AOI22_X1  g1031(.A1(new_n816), .A2(G128), .B1(new_n844), .B2(G137), .ZN(new_n1232));
  OAI21_X1  g1032(.A(new_n1232), .B1(new_n810), .B2(new_n1149), .ZN(new_n1233));
  AOI211_X1 g1033(.A(new_n1231), .B(new_n1233), .C1(G150), .C2(new_n800), .ZN(new_n1234));
  INV_X1    g1034(.A(new_n1234), .ZN(new_n1235));
  NAND2_X1  g1035(.A1(new_n1235), .A2(KEYINPUT59), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n827), .A2(G159), .ZN(new_n1237));
  AOI211_X1 g1037(.A(G33), .B(G41), .C1(new_n807), .C2(G124), .ZN(new_n1238));
  NAND3_X1  g1038(.A1(new_n1236), .A2(new_n1237), .A3(new_n1238), .ZN(new_n1239));
  NOR2_X1   g1039(.A1(new_n1235), .A2(KEYINPUT59), .ZN(new_n1240));
  OAI221_X1 g1040(.A(new_n1230), .B1(KEYINPUT58), .B2(new_n1229), .C1(new_n1239), .C2(new_n1240), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(new_n1241), .A2(new_n788), .ZN(new_n1242));
  OAI211_X1 g1042(.A(new_n1242), .B(new_n780), .C1(G50), .C2(new_n836), .ZN(new_n1243));
  NOR2_X1   g1043(.A1(new_n1218), .A2(new_n1243), .ZN(new_n1244));
  INV_X1    g1044(.A(new_n1244), .ZN(new_n1245));
  NAND3_X1  g1045(.A1(new_n1216), .A2(new_n1217), .A3(new_n1245), .ZN(new_n1246));
  AOI21_X1  g1046(.A(new_n773), .B1(new_n1210), .B2(new_n1214), .ZN(new_n1247));
  OAI21_X1  g1047(.A(KEYINPUT121), .B1(new_n1247), .B2(new_n1244), .ZN(new_n1248));
  NAND2_X1  g1048(.A1(new_n1246), .A2(new_n1248), .ZN(new_n1249));
  INV_X1    g1049(.A(new_n1182), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(new_n1186), .A2(new_n1250), .ZN(new_n1251));
  INV_X1    g1051(.A(KEYINPUT57), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(new_n1207), .A2(new_n1203), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(new_n949), .A2(new_n1253), .ZN(new_n1254));
  AOI21_X1  g1054(.A(new_n1252), .B1(new_n1254), .B2(new_n1214), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(new_n1251), .A2(new_n1255), .ZN(new_n1256));
  AOI22_X1  g1056(.A1(new_n1186), .A2(new_n1250), .B1(new_n1210), .B2(new_n1214), .ZN(new_n1257));
  OAI211_X1 g1057(.A(new_n1256), .B(new_n771), .C1(new_n1257), .C2(KEYINPUT57), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(new_n1249), .A2(new_n1258), .ZN(G375));
  NAND2_X1  g1059(.A1(new_n1173), .A2(new_n1176), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(new_n1177), .A2(new_n1179), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(new_n1260), .A2(new_n1261), .ZN(new_n1262));
  NAND2_X1  g1062(.A1(new_n945), .A2(new_n776), .ZN(new_n1263));
  OAI21_X1  g1063(.A(new_n780), .B1(G68), .B2(new_n836), .ZN(new_n1264));
  OAI22_X1  g1064(.A1(new_n1148), .A2(new_n839), .B1(new_n798), .B2(new_n1149), .ZN(new_n1265));
  AOI21_X1  g1065(.A(new_n1265), .B1(G50), .B2(new_n800), .ZN(new_n1266));
  OAI22_X1  g1066(.A1(new_n813), .A2(new_n850), .B1(new_n806), .B2(new_n1144), .ZN(new_n1267));
  OAI21_X1  g1067(.A(new_n341), .B1(new_n986), .B2(new_n810), .ZN(new_n1268));
  AOI211_X1 g1068(.A(new_n1267), .B(new_n1268), .C1(G137), .C2(new_n816), .ZN(new_n1269));
  NAND3_X1  g1069(.A1(new_n1266), .A2(new_n1269), .A3(new_n1228), .ZN(new_n1270));
  AOI22_X1  g1070(.A1(new_n803), .A2(G294), .B1(new_n844), .B2(G107), .ZN(new_n1271));
  OAI21_X1  g1071(.A(new_n1271), .B1(new_n506), .B2(new_n798), .ZN(new_n1272));
  XOR2_X1   g1072(.A(new_n1272), .B(KEYINPUT122), .Z(new_n1273));
  OAI221_X1 g1073(.A(new_n1080), .B1(new_n259), .B2(new_n793), .C1(new_n577), .C2(new_n810), .ZN(new_n1274));
  OAI221_X1 g1074(.A(new_n262), .B1(new_n806), .B2(new_n615), .C1(new_n815), .C2(new_n838), .ZN(new_n1275));
  OR2_X1    g1075(.A1(new_n1274), .A2(new_n1275), .ZN(new_n1276));
  OAI21_X1  g1076(.A(new_n1270), .B1(new_n1273), .B2(new_n1276), .ZN(new_n1277));
  AOI21_X1  g1077(.A(new_n1264), .B1(new_n1277), .B2(new_n788), .ZN(new_n1278));
  AOI22_X1  g1078(.A1(new_n1262), .A2(new_n774), .B1(new_n1263), .B2(new_n1278), .ZN(new_n1279));
  NAND2_X1  g1079(.A1(new_n1184), .A2(new_n1043), .ZN(new_n1280));
  NOR2_X1   g1080(.A1(new_n1250), .A2(new_n1262), .ZN(new_n1281));
  OAI21_X1  g1081(.A(new_n1279), .B1(new_n1280), .B2(new_n1281), .ZN(G381));
  NAND3_X1  g1082(.A1(new_n1249), .A2(new_n1187), .A3(new_n1258), .ZN(new_n1283));
  NOR3_X1   g1083(.A1(G384), .A2(G393), .A3(G396), .ZN(new_n1284));
  NAND2_X1  g1084(.A1(new_n1132), .A2(new_n1284), .ZN(new_n1285));
  OR4_X1    g1085(.A1(G387), .A2(new_n1283), .A3(G381), .A4(new_n1285), .ZN(G407));
  OAI211_X1 g1086(.A(G407), .B(G213), .C1(G343), .C2(new_n1283), .ZN(G409));
  NAND3_X1  g1087(.A1(new_n1249), .A2(G378), .A3(new_n1258), .ZN(new_n1288));
  NAND2_X1  g1088(.A1(new_n1257), .A2(new_n1043), .ZN(new_n1289));
  NAND2_X1  g1089(.A1(new_n1254), .A2(new_n1214), .ZN(new_n1290));
  AOI21_X1  g1090(.A(new_n1244), .B1(new_n1290), .B2(new_n774), .ZN(new_n1291));
  NAND2_X1  g1091(.A1(new_n1289), .A2(new_n1291), .ZN(new_n1292));
  NAND2_X1  g1092(.A1(new_n1292), .A2(new_n1187), .ZN(new_n1293));
  NAND2_X1  g1093(.A1(new_n1288), .A2(new_n1293), .ZN(new_n1294));
  NAND2_X1  g1094(.A1(new_n1294), .A2(KEYINPUT123), .ZN(new_n1295));
  NAND2_X1  g1095(.A1(new_n697), .A2(G213), .ZN(new_n1296));
  INV_X1    g1096(.A(KEYINPUT123), .ZN(new_n1297));
  NAND3_X1  g1097(.A1(new_n1288), .A2(new_n1297), .A3(new_n1293), .ZN(new_n1298));
  NAND3_X1  g1098(.A1(new_n1295), .A2(new_n1296), .A3(new_n1298), .ZN(new_n1299));
  AOI21_X1  g1099(.A(new_n1281), .B1(new_n1184), .B2(KEYINPUT60), .ZN(new_n1300));
  NAND3_X1  g1100(.A1(new_n1180), .A2(KEYINPUT60), .A3(new_n1182), .ZN(new_n1301));
  NAND2_X1  g1101(.A1(new_n1301), .A2(new_n771), .ZN(new_n1302));
  OAI21_X1  g1102(.A(new_n1279), .B1(new_n1300), .B2(new_n1302), .ZN(new_n1303));
  NOR2_X1   g1103(.A1(new_n1303), .A2(new_n887), .ZN(new_n1304));
  INV_X1    g1104(.A(new_n1304), .ZN(new_n1305));
  NAND2_X1  g1105(.A1(new_n1303), .A2(new_n887), .ZN(new_n1306));
  NAND2_X1  g1106(.A1(new_n1305), .A2(new_n1306), .ZN(new_n1307));
  INV_X1    g1107(.A(new_n1296), .ZN(new_n1308));
  NAND2_X1  g1108(.A1(new_n1308), .A2(G2897), .ZN(new_n1309));
  NOR2_X1   g1109(.A1(new_n1307), .A2(new_n1309), .ZN(new_n1310));
  AOI22_X1  g1110(.A1(new_n1305), .A2(new_n1306), .B1(G2897), .B2(new_n1308), .ZN(new_n1311));
  OR2_X1    g1111(.A1(new_n1310), .A2(new_n1311), .ZN(new_n1312));
  NAND2_X1  g1112(.A1(new_n1299), .A2(new_n1312), .ZN(new_n1313));
  XNOR2_X1  g1113(.A(G393), .B(G396), .ZN(new_n1314));
  INV_X1    g1114(.A(new_n1314), .ZN(new_n1315));
  OAI21_X1  g1115(.A(new_n1315), .B1(new_n1105), .B2(new_n1131), .ZN(new_n1316));
  NAND2_X1  g1116(.A1(new_n1103), .A2(new_n1104), .ZN(new_n1317));
  XNOR2_X1  g1117(.A(new_n1098), .B(new_n709), .ZN(new_n1318));
  AOI21_X1  g1118(.A(new_n718), .B1(new_n1318), .B2(new_n1032), .ZN(new_n1319));
  NAND2_X1  g1119(.A1(new_n1317), .A2(new_n1319), .ZN(new_n1320));
  NAND4_X1  g1120(.A1(new_n1320), .A2(new_n1106), .A3(new_n1130), .A4(new_n1314), .ZN(new_n1321));
  NAND2_X1  g1121(.A1(new_n1316), .A2(new_n1321), .ZN(new_n1322));
  NAND2_X1  g1122(.A1(G387), .A2(new_n1322), .ZN(new_n1323));
  AND3_X1   g1123(.A1(new_n1056), .A2(new_n1059), .A3(new_n1060), .ZN(new_n1324));
  AOI21_X1  g1124(.A(new_n1042), .B1(new_n1317), .B2(new_n768), .ZN(new_n1325));
  OAI21_X1  g1125(.A(new_n1324), .B1(new_n1325), .B2(new_n774), .ZN(new_n1326));
  NAND4_X1  g1126(.A1(new_n1326), .A2(new_n1007), .A3(new_n1316), .A4(new_n1321), .ZN(new_n1327));
  INV_X1    g1127(.A(KEYINPUT61), .ZN(new_n1328));
  NAND3_X1  g1128(.A1(new_n1323), .A2(new_n1327), .A3(new_n1328), .ZN(new_n1329));
  AOI21_X1  g1129(.A(new_n1308), .B1(new_n1288), .B2(new_n1293), .ZN(new_n1330));
  INV_X1    g1130(.A(new_n1306), .ZN(new_n1331));
  NOR2_X1   g1131(.A1(new_n1331), .A2(new_n1304), .ZN(new_n1332));
  AND2_X1   g1132(.A1(new_n1332), .A2(KEYINPUT63), .ZN(new_n1333));
  AOI21_X1  g1133(.A(new_n1329), .B1(new_n1330), .B2(new_n1333), .ZN(new_n1334));
  NAND4_X1  g1134(.A1(new_n1295), .A2(new_n1296), .A3(new_n1332), .A4(new_n1298), .ZN(new_n1335));
  INV_X1    g1135(.A(new_n1335), .ZN(new_n1336));
  OAI211_X1 g1136(.A(new_n1313), .B(new_n1334), .C1(new_n1336), .C2(KEYINPUT63), .ZN(new_n1337));
  XOR2_X1   g1137(.A(KEYINPUT124), .B(KEYINPUT61), .Z(new_n1338));
  NOR2_X1   g1138(.A1(new_n1310), .A2(new_n1311), .ZN(new_n1339));
  OAI21_X1  g1139(.A(new_n1338), .B1(new_n1339), .B2(new_n1330), .ZN(new_n1340));
  INV_X1    g1140(.A(KEYINPUT62), .ZN(new_n1341));
  NAND2_X1  g1141(.A1(new_n1335), .A2(new_n1341), .ZN(new_n1342));
  NAND3_X1  g1142(.A1(new_n1330), .A2(KEYINPUT62), .A3(new_n1332), .ZN(new_n1343));
  AOI21_X1  g1143(.A(new_n1340), .B1(new_n1342), .B2(new_n1343), .ZN(new_n1344));
  AND3_X1   g1144(.A1(new_n1323), .A2(new_n1327), .A3(KEYINPUT125), .ZN(new_n1345));
  AOI21_X1  g1145(.A(KEYINPUT125), .B1(new_n1323), .B2(new_n1327), .ZN(new_n1346));
  NOR2_X1   g1146(.A1(new_n1345), .A2(new_n1346), .ZN(new_n1347));
  OAI21_X1  g1147(.A(new_n1337), .B1(new_n1344), .B2(new_n1347), .ZN(G405));
  INV_X1    g1148(.A(new_n1288), .ZN(new_n1349));
  AOI21_X1  g1149(.A(G378), .B1(new_n1249), .B2(new_n1258), .ZN(new_n1350));
  NOR3_X1   g1150(.A1(new_n1349), .A2(new_n1350), .A3(new_n1332), .ZN(new_n1351));
  NAND2_X1  g1151(.A1(G375), .A2(new_n1187), .ZN(new_n1352));
  AOI21_X1  g1152(.A(new_n1307), .B1(new_n1352), .B2(new_n1288), .ZN(new_n1353));
  OAI21_X1  g1153(.A(KEYINPUT126), .B1(new_n1351), .B2(new_n1353), .ZN(new_n1354));
  NAND2_X1  g1154(.A1(new_n1354), .A2(KEYINPUT127), .ZN(new_n1355));
  OAI21_X1  g1155(.A(new_n1332), .B1(new_n1349), .B2(new_n1350), .ZN(new_n1356));
  NAND3_X1  g1156(.A1(new_n1352), .A2(new_n1307), .A3(new_n1288), .ZN(new_n1357));
  NAND2_X1  g1157(.A1(new_n1356), .A2(new_n1357), .ZN(new_n1358));
  INV_X1    g1158(.A(KEYINPUT127), .ZN(new_n1359));
  NAND3_X1  g1159(.A1(new_n1358), .A2(KEYINPUT126), .A3(new_n1359), .ZN(new_n1360));
  INV_X1    g1160(.A(KEYINPUT126), .ZN(new_n1361));
  NAND3_X1  g1161(.A1(new_n1356), .A2(new_n1357), .A3(new_n1361), .ZN(new_n1362));
  NAND4_X1  g1162(.A1(new_n1355), .A2(new_n1347), .A3(new_n1360), .A4(new_n1362), .ZN(new_n1363));
  NAND2_X1  g1163(.A1(new_n1347), .A2(new_n1362), .ZN(new_n1364));
  AOI21_X1  g1164(.A(new_n1359), .B1(new_n1358), .B2(KEYINPUT126), .ZN(new_n1365));
  AOI211_X1 g1165(.A(new_n1361), .B(KEYINPUT127), .C1(new_n1356), .C2(new_n1357), .ZN(new_n1366));
  OAI21_X1  g1166(.A(new_n1364), .B1(new_n1365), .B2(new_n1366), .ZN(new_n1367));
  NAND2_X1  g1167(.A1(new_n1363), .A2(new_n1367), .ZN(G402));
endmodule


