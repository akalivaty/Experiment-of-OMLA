

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302,
         n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313,
         n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324,
         n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335,
         n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346,
         n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590, n591;

  XNOR2_X1 U324 ( .A(n342), .B(n341), .ZN(n343) );
  XNOR2_X1 U325 ( .A(n339), .B(n338), .ZN(n344) );
  XNOR2_X1 U326 ( .A(n337), .B(n336), .ZN(n338) );
  XNOR2_X1 U327 ( .A(n569), .B(n345), .ZN(n554) );
  XNOR2_X1 U328 ( .A(KEYINPUT7), .B(G50GAT), .ZN(n329) );
  XNOR2_X1 U329 ( .A(n327), .B(n326), .ZN(n331) );
  INV_X1 U330 ( .A(n572), .ZN(n367) );
  XNOR2_X1 U331 ( .A(n331), .B(n330), .ZN(n333) );
  XNOR2_X1 U332 ( .A(KEYINPUT55), .B(KEYINPUT124), .ZN(n441) );
  XNOR2_X1 U333 ( .A(n442), .B(n441), .ZN(n462) );
  AND2_X1 U334 ( .A1(n462), .A2(n542), .ZN(n571) );
  XNOR2_X1 U335 ( .A(n344), .B(n343), .ZN(n569) );
  XNOR2_X1 U336 ( .A(n459), .B(G176GAT), .ZN(n460) );
  XNOR2_X1 U337 ( .A(n461), .B(n460), .ZN(G1349GAT) );
  XOR2_X1 U338 ( .A(KEYINPUT33), .B(KEYINPUT31), .Z(n293) );
  NAND2_X1 U339 ( .A1(G230GAT), .A2(G233GAT), .ZN(n292) );
  XNOR2_X1 U340 ( .A(n293), .B(n292), .ZN(n294) );
  XOR2_X1 U341 ( .A(n294), .B(KEYINPUT32), .Z(n300) );
  XOR2_X1 U342 ( .A(G92GAT), .B(G85GAT), .Z(n296) );
  XNOR2_X1 U343 ( .A(G99GAT), .B(G106GAT), .ZN(n295) );
  XNOR2_X1 U344 ( .A(n296), .B(n295), .ZN(n337) );
  XOR2_X1 U345 ( .A(KEYINPUT74), .B(KEYINPUT13), .Z(n298) );
  XNOR2_X1 U346 ( .A(G71GAT), .B(G78GAT), .ZN(n297) );
  XNOR2_X1 U347 ( .A(n298), .B(n297), .ZN(n323) );
  XNOR2_X1 U348 ( .A(n337), .B(n323), .ZN(n299) );
  XNOR2_X1 U349 ( .A(n300), .B(n299), .ZN(n304) );
  XOR2_X1 U350 ( .A(KEYINPUT75), .B(KEYINPUT76), .Z(n302) );
  XNOR2_X1 U351 ( .A(G148GAT), .B(G204GAT), .ZN(n301) );
  XNOR2_X1 U352 ( .A(n302), .B(n301), .ZN(n303) );
  XOR2_X1 U353 ( .A(n304), .B(n303), .Z(n306) );
  XOR2_X1 U354 ( .A(G120GAT), .B(G57GAT), .Z(n404) );
  XOR2_X1 U355 ( .A(G176GAT), .B(G64GAT), .Z(n378) );
  XNOR2_X1 U356 ( .A(n404), .B(n378), .ZN(n305) );
  XNOR2_X1 U357 ( .A(n306), .B(n305), .ZN(n583) );
  XOR2_X1 U358 ( .A(KEYINPUT41), .B(n583), .Z(n562) );
  INV_X1 U359 ( .A(n583), .ZN(n350) );
  INV_X1 U360 ( .A(KEYINPUT45), .ZN(n348) );
  XOR2_X1 U361 ( .A(G211GAT), .B(G155GAT), .Z(n308) );
  XNOR2_X1 U362 ( .A(G183GAT), .B(G127GAT), .ZN(n307) );
  XNOR2_X1 U363 ( .A(n308), .B(n307), .ZN(n312) );
  XOR2_X1 U364 ( .A(G64GAT), .B(G57GAT), .Z(n310) );
  XNOR2_X1 U365 ( .A(G1GAT), .B(G8GAT), .ZN(n309) );
  XNOR2_X1 U366 ( .A(n310), .B(n309), .ZN(n311) );
  XOR2_X1 U367 ( .A(n312), .B(n311), .Z(n317) );
  XOR2_X1 U368 ( .A(KEYINPUT81), .B(KEYINPUT82), .Z(n314) );
  NAND2_X1 U369 ( .A1(G231GAT), .A2(G233GAT), .ZN(n313) );
  XNOR2_X1 U370 ( .A(n314), .B(n313), .ZN(n315) );
  XNOR2_X1 U371 ( .A(KEYINPUT79), .B(n315), .ZN(n316) );
  XNOR2_X1 U372 ( .A(n317), .B(n316), .ZN(n321) );
  XOR2_X1 U373 ( .A(KEYINPUT80), .B(KEYINPUT15), .Z(n319) );
  XNOR2_X1 U374 ( .A(KEYINPUT12), .B(KEYINPUT14), .ZN(n318) );
  XNOR2_X1 U375 ( .A(n319), .B(n318), .ZN(n320) );
  XOR2_X1 U376 ( .A(n321), .B(n320), .Z(n325) );
  XNOR2_X1 U377 ( .A(G15GAT), .B(G22GAT), .ZN(n322) );
  XNOR2_X1 U378 ( .A(n322), .B(KEYINPUT70), .ZN(n359) );
  XNOR2_X1 U379 ( .A(n359), .B(n323), .ZN(n324) );
  XNOR2_X1 U380 ( .A(n325), .B(n324), .ZN(n550) );
  INV_X1 U381 ( .A(n550), .ZN(n587) );
  XNOR2_X1 U382 ( .A(KEYINPUT36), .B(KEYINPUT107), .ZN(n346) );
  XOR2_X1 U383 ( .A(G43GAT), .B(G29GAT), .Z(n327) );
  XNOR2_X1 U384 ( .A(G36GAT), .B(KEYINPUT8), .ZN(n326) );
  INV_X1 U385 ( .A(KEYINPUT69), .ZN(n328) );
  XNOR2_X1 U386 ( .A(n329), .B(n328), .ZN(n330) );
  INV_X1 U387 ( .A(n333), .ZN(n352) );
  XOR2_X1 U388 ( .A(G190GAT), .B(G218GAT), .Z(n390) );
  INV_X1 U389 ( .A(n390), .ZN(n332) );
  NAND2_X1 U390 ( .A1(n352), .A2(n332), .ZN(n335) );
  NAND2_X1 U391 ( .A1(n333), .A2(n390), .ZN(n334) );
  NAND2_X1 U392 ( .A1(n335), .A2(n334), .ZN(n339) );
  NAND2_X1 U393 ( .A1(G232GAT), .A2(G233GAT), .ZN(n336) );
  XOR2_X1 U394 ( .A(G134GAT), .B(G162GAT), .Z(n407) );
  XNOR2_X1 U395 ( .A(n407), .B(KEYINPUT9), .ZN(n340) );
  XNOR2_X1 U396 ( .A(n340), .B(KEYINPUT11), .ZN(n342) );
  XNOR2_X1 U397 ( .A(KEYINPUT77), .B(KEYINPUT10), .ZN(n341) );
  INV_X1 U398 ( .A(KEYINPUT78), .ZN(n345) );
  XNOR2_X1 U399 ( .A(n346), .B(n554), .ZN(n498) );
  NOR2_X1 U400 ( .A1(n587), .A2(n498), .ZN(n347) );
  XNOR2_X1 U401 ( .A(n348), .B(n347), .ZN(n349) );
  NOR2_X1 U402 ( .A1(n350), .A2(n349), .ZN(n351) );
  XNOR2_X1 U403 ( .A(n351), .B(KEYINPUT118), .ZN(n368) );
  XOR2_X1 U404 ( .A(KEYINPUT72), .B(KEYINPUT71), .Z(n354) );
  XNOR2_X1 U405 ( .A(KEYINPUT30), .B(KEYINPUT29), .ZN(n353) );
  XNOR2_X1 U406 ( .A(n354), .B(n353), .ZN(n355) );
  XNOR2_X1 U407 ( .A(n333), .B(n355), .ZN(n366) );
  XOR2_X1 U408 ( .A(KEYINPUT66), .B(KEYINPUT67), .Z(n357) );
  XOR2_X1 U409 ( .A(G113GAT), .B(G1GAT), .Z(n417) );
  XOR2_X1 U410 ( .A(G169GAT), .B(G8GAT), .Z(n381) );
  XNOR2_X1 U411 ( .A(n417), .B(n381), .ZN(n356) );
  XNOR2_X1 U412 ( .A(n357), .B(n356), .ZN(n358) );
  XOR2_X1 U413 ( .A(n358), .B(G197GAT), .Z(n364) );
  XOR2_X1 U414 ( .A(n359), .B(KEYINPUT68), .Z(n361) );
  NAND2_X1 U415 ( .A1(G229GAT), .A2(G233GAT), .ZN(n360) );
  XNOR2_X1 U416 ( .A(n361), .B(n360), .ZN(n362) );
  XNOR2_X1 U417 ( .A(n362), .B(G141GAT), .ZN(n363) );
  XNOR2_X1 U418 ( .A(n364), .B(n363), .ZN(n365) );
  XOR2_X1 U419 ( .A(n366), .B(n365), .Z(n579) );
  XNOR2_X1 U420 ( .A(n579), .B(KEYINPUT73), .ZN(n572) );
  AND2_X1 U421 ( .A1(n368), .A2(n367), .ZN(n375) );
  XOR2_X1 U422 ( .A(KEYINPUT117), .B(KEYINPUT47), .Z(n373) );
  NOR2_X1 U423 ( .A1(n562), .A2(n579), .ZN(n369) );
  XNOR2_X1 U424 ( .A(n369), .B(KEYINPUT46), .ZN(n370) );
  NOR2_X1 U425 ( .A1(n550), .A2(n370), .ZN(n371) );
  NAND2_X1 U426 ( .A1(n371), .A2(n569), .ZN(n372) );
  XNOR2_X1 U427 ( .A(n373), .B(n372), .ZN(n374) );
  NOR2_X1 U428 ( .A1(n375), .A2(n374), .ZN(n377) );
  XNOR2_X1 U429 ( .A(KEYINPUT48), .B(KEYINPUT64), .ZN(n376) );
  XNOR2_X1 U430 ( .A(n377), .B(n376), .ZN(n540) );
  XOR2_X1 U431 ( .A(n378), .B(KEYINPUT99), .Z(n380) );
  NAND2_X1 U432 ( .A1(G226GAT), .A2(G233GAT), .ZN(n379) );
  XNOR2_X1 U433 ( .A(n380), .B(n379), .ZN(n384) );
  XNOR2_X1 U434 ( .A(G36GAT), .B(n381), .ZN(n382) );
  XNOR2_X1 U435 ( .A(n382), .B(G92GAT), .ZN(n383) );
  XOR2_X1 U436 ( .A(n384), .B(n383), .Z(n392) );
  XOR2_X1 U437 ( .A(KEYINPUT87), .B(KEYINPUT88), .Z(n386) );
  XNOR2_X1 U438 ( .A(KEYINPUT89), .B(KEYINPUT21), .ZN(n385) );
  XNOR2_X1 U439 ( .A(n386), .B(n385), .ZN(n387) );
  XOR2_X1 U440 ( .A(n387), .B(G211GAT), .Z(n389) );
  XNOR2_X1 U441 ( .A(G197GAT), .B(G204GAT), .ZN(n388) );
  XNOR2_X1 U442 ( .A(n389), .B(n388), .ZN(n436) );
  XNOR2_X1 U443 ( .A(n436), .B(n390), .ZN(n391) );
  XNOR2_X1 U444 ( .A(n392), .B(n391), .ZN(n397) );
  XOR2_X1 U445 ( .A(KEYINPUT84), .B(KEYINPUT17), .Z(n394) );
  XNOR2_X1 U446 ( .A(KEYINPUT18), .B(G183GAT), .ZN(n393) );
  XNOR2_X1 U447 ( .A(n394), .B(n393), .ZN(n395) );
  XOR2_X1 U448 ( .A(KEYINPUT19), .B(n395), .Z(n456) );
  INV_X1 U449 ( .A(n456), .ZN(n396) );
  XOR2_X1 U450 ( .A(n397), .B(n396), .Z(n473) );
  INV_X1 U451 ( .A(n473), .ZN(n530) );
  NOR2_X1 U452 ( .A1(n540), .A2(n530), .ZN(n398) );
  XNOR2_X1 U453 ( .A(n398), .B(KEYINPUT54), .ZN(n422) );
  XOR2_X1 U454 ( .A(KEYINPUT6), .B(KEYINPUT96), .Z(n400) );
  XNOR2_X1 U455 ( .A(KEYINPUT94), .B(KEYINPUT4), .ZN(n399) );
  XNOR2_X1 U456 ( .A(n400), .B(n399), .ZN(n421) );
  XOR2_X1 U457 ( .A(KEYINPUT1), .B(KEYINPUT97), .Z(n402) );
  XNOR2_X1 U458 ( .A(KEYINPUT95), .B(KEYINPUT5), .ZN(n401) );
  XNOR2_X1 U459 ( .A(n402), .B(n401), .ZN(n403) );
  XOR2_X1 U460 ( .A(n403), .B(G85GAT), .Z(n406) );
  XNOR2_X1 U461 ( .A(G29GAT), .B(n404), .ZN(n405) );
  XNOR2_X1 U462 ( .A(n406), .B(n405), .ZN(n411) );
  XOR2_X1 U463 ( .A(KEYINPUT0), .B(G127GAT), .Z(n446) );
  XOR2_X1 U464 ( .A(n407), .B(n446), .Z(n409) );
  NAND2_X1 U465 ( .A1(G225GAT), .A2(G233GAT), .ZN(n408) );
  XNOR2_X1 U466 ( .A(n409), .B(n408), .ZN(n410) );
  XOR2_X1 U467 ( .A(n411), .B(n410), .Z(n419) );
  XOR2_X1 U468 ( .A(KEYINPUT3), .B(G148GAT), .Z(n413) );
  XNOR2_X1 U469 ( .A(G141GAT), .B(G155GAT), .ZN(n412) );
  XNOR2_X1 U470 ( .A(n413), .B(n412), .ZN(n415) );
  XOR2_X1 U471 ( .A(KEYINPUT2), .B(KEYINPUT90), .Z(n414) );
  XNOR2_X1 U472 ( .A(n415), .B(n414), .ZN(n440) );
  INV_X1 U473 ( .A(n440), .ZN(n416) );
  XNOR2_X1 U474 ( .A(n417), .B(n416), .ZN(n418) );
  XNOR2_X1 U475 ( .A(n419), .B(n418), .ZN(n420) );
  XOR2_X1 U476 ( .A(n421), .B(n420), .Z(n483) );
  XNOR2_X1 U477 ( .A(KEYINPUT98), .B(n483), .ZN(n528) );
  NAND2_X1 U478 ( .A1(n422), .A2(n528), .ZN(n423) );
  XNOR2_X1 U479 ( .A(n423), .B(KEYINPUT65), .ZN(n577) );
  XOR2_X1 U480 ( .A(G78GAT), .B(KEYINPUT86), .Z(n425) );
  XNOR2_X1 U481 ( .A(KEYINPUT24), .B(KEYINPUT23), .ZN(n424) );
  XNOR2_X1 U482 ( .A(n425), .B(n424), .ZN(n429) );
  XOR2_X1 U483 ( .A(KEYINPUT92), .B(KEYINPUT93), .Z(n427) );
  XNOR2_X1 U484 ( .A(G22GAT), .B(KEYINPUT22), .ZN(n426) );
  XNOR2_X1 U485 ( .A(n427), .B(n426), .ZN(n428) );
  XOR2_X1 U486 ( .A(n429), .B(n428), .Z(n438) );
  XOR2_X1 U487 ( .A(G106GAT), .B(G162GAT), .Z(n431) );
  XNOR2_X1 U488 ( .A(G50GAT), .B(G218GAT), .ZN(n430) );
  XNOR2_X1 U489 ( .A(n431), .B(n430), .ZN(n432) );
  XOR2_X1 U490 ( .A(KEYINPUT91), .B(n432), .Z(n434) );
  NAND2_X1 U491 ( .A1(G228GAT), .A2(G233GAT), .ZN(n433) );
  XNOR2_X1 U492 ( .A(n434), .B(n433), .ZN(n435) );
  XNOR2_X1 U493 ( .A(n436), .B(n435), .ZN(n437) );
  XNOR2_X1 U494 ( .A(n438), .B(n437), .ZN(n439) );
  XNOR2_X1 U495 ( .A(n440), .B(n439), .ZN(n477) );
  NAND2_X1 U496 ( .A1(n577), .A2(n477), .ZN(n442) );
  XOR2_X1 U497 ( .A(G99GAT), .B(G134GAT), .Z(n444) );
  XNOR2_X1 U498 ( .A(G43GAT), .B(G190GAT), .ZN(n443) );
  XNOR2_X1 U499 ( .A(n444), .B(n443), .ZN(n445) );
  XOR2_X1 U500 ( .A(n446), .B(n445), .Z(n448) );
  NAND2_X1 U501 ( .A1(G227GAT), .A2(G233GAT), .ZN(n447) );
  XNOR2_X1 U502 ( .A(n448), .B(n447), .ZN(n452) );
  XOR2_X1 U503 ( .A(KEYINPUT20), .B(G176GAT), .Z(n450) );
  XNOR2_X1 U504 ( .A(G169GAT), .B(G120GAT), .ZN(n449) );
  XNOR2_X1 U505 ( .A(n450), .B(n449), .ZN(n451) );
  XOR2_X1 U506 ( .A(n452), .B(n451), .Z(n458) );
  XOR2_X1 U507 ( .A(KEYINPUT85), .B(G71GAT), .Z(n454) );
  XNOR2_X1 U508 ( .A(G15GAT), .B(G113GAT), .ZN(n453) );
  XNOR2_X1 U509 ( .A(n454), .B(n453), .ZN(n455) );
  XNOR2_X1 U510 ( .A(n456), .B(n455), .ZN(n457) );
  XNOR2_X1 U511 ( .A(n458), .B(n457), .ZN(n542) );
  NAND2_X1 U512 ( .A1(n462), .A2(n542), .ZN(n574) );
  NOR2_X1 U513 ( .A1(n562), .A2(n574), .ZN(n461) );
  XNOR2_X1 U514 ( .A(KEYINPUT56), .B(KEYINPUT57), .ZN(n459) );
  INV_X1 U515 ( .A(G190GAT), .ZN(n466) );
  XOR2_X1 U516 ( .A(KEYINPUT58), .B(KEYINPUT126), .Z(n464) );
  NAND2_X1 U517 ( .A1(n571), .A2(n554), .ZN(n463) );
  XNOR2_X1 U518 ( .A(n464), .B(n463), .ZN(n465) );
  XNOR2_X1 U519 ( .A(n466), .B(n465), .ZN(G1351GAT) );
  XOR2_X1 U520 ( .A(KEYINPUT103), .B(KEYINPUT34), .Z(n468) );
  XNOR2_X1 U521 ( .A(G1GAT), .B(KEYINPUT102), .ZN(n467) );
  XNOR2_X1 U522 ( .A(n468), .B(n467), .ZN(n488) );
  NAND2_X1 U523 ( .A1(n572), .A2(n583), .ZN(n503) );
  NOR2_X1 U524 ( .A1(n587), .A2(n554), .ZN(n469) );
  XOR2_X1 U525 ( .A(KEYINPUT83), .B(n469), .Z(n470) );
  XNOR2_X1 U526 ( .A(n470), .B(KEYINPUT16), .ZN(n486) );
  XOR2_X1 U527 ( .A(n530), .B(KEYINPUT27), .Z(n479) );
  INV_X1 U528 ( .A(n479), .ZN(n471) );
  NOR2_X1 U529 ( .A1(n528), .A2(n471), .ZN(n472) );
  XOR2_X1 U530 ( .A(KEYINPUT100), .B(n472), .Z(n558) );
  XOR2_X1 U531 ( .A(n477), .B(KEYINPUT28), .Z(n495) );
  NOR2_X1 U532 ( .A1(n558), .A2(n495), .ZN(n541) );
  INV_X1 U533 ( .A(n542), .ZN(n532) );
  NAND2_X1 U534 ( .A1(n541), .A2(n532), .ZN(n485) );
  NAND2_X1 U535 ( .A1(n473), .A2(n542), .ZN(n474) );
  NAND2_X1 U536 ( .A1(n474), .A2(n477), .ZN(n475) );
  XNOR2_X1 U537 ( .A(n475), .B(KEYINPUT25), .ZN(n476) );
  XNOR2_X1 U538 ( .A(n476), .B(KEYINPUT101), .ZN(n481) );
  NOR2_X1 U539 ( .A1(n477), .A2(n542), .ZN(n478) );
  XNOR2_X1 U540 ( .A(n478), .B(KEYINPUT26), .ZN(n578) );
  NAND2_X1 U541 ( .A1(n479), .A2(n578), .ZN(n480) );
  NAND2_X1 U542 ( .A1(n481), .A2(n480), .ZN(n482) );
  NAND2_X1 U543 ( .A1(n483), .A2(n482), .ZN(n484) );
  NAND2_X1 U544 ( .A1(n485), .A2(n484), .ZN(n499) );
  NAND2_X1 U545 ( .A1(n486), .A2(n499), .ZN(n516) );
  OR2_X1 U546 ( .A1(n503), .A2(n516), .ZN(n496) );
  NOR2_X1 U547 ( .A1(n528), .A2(n496), .ZN(n487) );
  XOR2_X1 U548 ( .A(n488), .B(n487), .Z(G1324GAT) );
  NOR2_X1 U549 ( .A1(n530), .A2(n496), .ZN(n490) );
  XNOR2_X1 U550 ( .A(KEYINPUT104), .B(KEYINPUT105), .ZN(n489) );
  XNOR2_X1 U551 ( .A(n490), .B(n489), .ZN(n491) );
  XNOR2_X1 U552 ( .A(G8GAT), .B(n491), .ZN(G1325GAT) );
  NOR2_X1 U553 ( .A1(n532), .A2(n496), .ZN(n493) );
  XNOR2_X1 U554 ( .A(KEYINPUT106), .B(KEYINPUT35), .ZN(n492) );
  XNOR2_X1 U555 ( .A(n493), .B(n492), .ZN(n494) );
  XNOR2_X1 U556 ( .A(G15GAT), .B(n494), .ZN(G1326GAT) );
  INV_X1 U557 ( .A(n495), .ZN(n535) );
  NOR2_X1 U558 ( .A1(n535), .A2(n496), .ZN(n497) );
  XOR2_X1 U559 ( .A(G22GAT), .B(n497), .Z(G1327GAT) );
  NAND2_X1 U560 ( .A1(n587), .A2(n499), .ZN(n500) );
  NOR2_X1 U561 ( .A1(n498), .A2(n500), .ZN(n502) );
  XNOR2_X1 U562 ( .A(KEYINPUT108), .B(KEYINPUT37), .ZN(n501) );
  XNOR2_X1 U563 ( .A(n502), .B(n501), .ZN(n526) );
  NOR2_X1 U564 ( .A1(n503), .A2(n526), .ZN(n504) );
  XOR2_X1 U565 ( .A(KEYINPUT38), .B(n504), .Z(n512) );
  NOR2_X1 U566 ( .A1(n512), .A2(n528), .ZN(n506) );
  XNOR2_X1 U567 ( .A(G29GAT), .B(KEYINPUT39), .ZN(n505) );
  XNOR2_X1 U568 ( .A(n506), .B(n505), .ZN(G1328GAT) );
  NOR2_X1 U569 ( .A1(n530), .A2(n512), .ZN(n507) );
  XOR2_X1 U570 ( .A(G36GAT), .B(n507), .Z(G1329GAT) );
  XOR2_X1 U571 ( .A(KEYINPUT110), .B(KEYINPUT40), .Z(n509) );
  XNOR2_X1 U572 ( .A(G43GAT), .B(KEYINPUT109), .ZN(n508) );
  XNOR2_X1 U573 ( .A(n509), .B(n508), .ZN(n511) );
  NOR2_X1 U574 ( .A1(n512), .A2(n532), .ZN(n510) );
  XOR2_X1 U575 ( .A(n511), .B(n510), .Z(G1330GAT) );
  NOR2_X1 U576 ( .A1(n512), .A2(n535), .ZN(n513) );
  XOR2_X1 U577 ( .A(G50GAT), .B(n513), .Z(G1331GAT) );
  XOR2_X1 U578 ( .A(KEYINPUT112), .B(KEYINPUT42), .Z(n515) );
  XNOR2_X1 U579 ( .A(G57GAT), .B(KEYINPUT111), .ZN(n514) );
  XNOR2_X1 U580 ( .A(n515), .B(n514), .ZN(n518) );
  INV_X1 U581 ( .A(n562), .ZN(n545) );
  NAND2_X1 U582 ( .A1(n579), .A2(n545), .ZN(n525) );
  OR2_X1 U583 ( .A1(n525), .A2(n516), .ZN(n521) );
  NOR2_X1 U584 ( .A1(n528), .A2(n521), .ZN(n517) );
  XOR2_X1 U585 ( .A(n518), .B(n517), .Z(G1332GAT) );
  NOR2_X1 U586 ( .A1(n530), .A2(n521), .ZN(n519) );
  XOR2_X1 U587 ( .A(G64GAT), .B(n519), .Z(G1333GAT) );
  NOR2_X1 U588 ( .A1(n532), .A2(n521), .ZN(n520) );
  XOR2_X1 U589 ( .A(G71GAT), .B(n520), .Z(G1334GAT) );
  NOR2_X1 U590 ( .A1(n535), .A2(n521), .ZN(n523) );
  XNOR2_X1 U591 ( .A(KEYINPUT113), .B(KEYINPUT43), .ZN(n522) );
  XNOR2_X1 U592 ( .A(n523), .B(n522), .ZN(n524) );
  XOR2_X1 U593 ( .A(G78GAT), .B(n524), .Z(G1335GAT) );
  NOR2_X1 U594 ( .A1(n526), .A2(n525), .ZN(n527) );
  XOR2_X1 U595 ( .A(KEYINPUT114), .B(n527), .Z(n536) );
  NOR2_X1 U596 ( .A1(n536), .A2(n528), .ZN(n529) );
  XOR2_X1 U597 ( .A(G85GAT), .B(n529), .Z(G1336GAT) );
  NOR2_X1 U598 ( .A1(n530), .A2(n536), .ZN(n531) );
  XOR2_X1 U599 ( .A(G92GAT), .B(n531), .Z(G1337GAT) );
  NOR2_X1 U600 ( .A1(n536), .A2(n532), .ZN(n534) );
  XNOR2_X1 U601 ( .A(G99GAT), .B(KEYINPUT115), .ZN(n533) );
  XNOR2_X1 U602 ( .A(n534), .B(n533), .ZN(G1338GAT) );
  NOR2_X1 U603 ( .A1(n536), .A2(n535), .ZN(n538) );
  XNOR2_X1 U604 ( .A(KEYINPUT44), .B(KEYINPUT116), .ZN(n537) );
  XNOR2_X1 U605 ( .A(n538), .B(n537), .ZN(n539) );
  XOR2_X1 U606 ( .A(G106GAT), .B(n539), .Z(G1339GAT) );
  NAND2_X1 U607 ( .A1(n542), .A2(n541), .ZN(n543) );
  NOR2_X1 U608 ( .A1(n540), .A2(n543), .ZN(n555) );
  NAND2_X1 U609 ( .A1(n572), .A2(n555), .ZN(n544) );
  XNOR2_X1 U610 ( .A(G113GAT), .B(n544), .ZN(G1340GAT) );
  XOR2_X1 U611 ( .A(G120GAT), .B(KEYINPUT120), .Z(n547) );
  NAND2_X1 U612 ( .A1(n555), .A2(n545), .ZN(n546) );
  XNOR2_X1 U613 ( .A(n547), .B(n546), .ZN(n549) );
  XOR2_X1 U614 ( .A(KEYINPUT119), .B(KEYINPUT49), .Z(n548) );
  XNOR2_X1 U615 ( .A(n549), .B(n548), .ZN(G1341GAT) );
  XOR2_X1 U616 ( .A(KEYINPUT50), .B(KEYINPUT121), .Z(n552) );
  NAND2_X1 U617 ( .A1(n555), .A2(n550), .ZN(n551) );
  XNOR2_X1 U618 ( .A(n552), .B(n551), .ZN(n553) );
  XNOR2_X1 U619 ( .A(G127GAT), .B(n553), .ZN(G1342GAT) );
  XOR2_X1 U620 ( .A(G134GAT), .B(KEYINPUT51), .Z(n557) );
  NAND2_X1 U621 ( .A1(n555), .A2(n554), .ZN(n556) );
  XNOR2_X1 U622 ( .A(n557), .B(n556), .ZN(G1343GAT) );
  NOR2_X1 U623 ( .A1(n540), .A2(n558), .ZN(n559) );
  NAND2_X1 U624 ( .A1(n559), .A2(n578), .ZN(n568) );
  NOR2_X1 U625 ( .A1(n579), .A2(n568), .ZN(n560) );
  XOR2_X1 U626 ( .A(KEYINPUT122), .B(n560), .Z(n561) );
  XNOR2_X1 U627 ( .A(G141GAT), .B(n561), .ZN(G1344GAT) );
  NOR2_X1 U628 ( .A1(n568), .A2(n562), .ZN(n566) );
  XOR2_X1 U629 ( .A(KEYINPUT53), .B(KEYINPUT52), .Z(n564) );
  XNOR2_X1 U630 ( .A(G148GAT), .B(KEYINPUT123), .ZN(n563) );
  XNOR2_X1 U631 ( .A(n564), .B(n563), .ZN(n565) );
  XNOR2_X1 U632 ( .A(n566), .B(n565), .ZN(G1345GAT) );
  NOR2_X1 U633 ( .A1(n587), .A2(n568), .ZN(n567) );
  XOR2_X1 U634 ( .A(G155GAT), .B(n567), .Z(G1346GAT) );
  NOR2_X1 U635 ( .A1(n569), .A2(n568), .ZN(n570) );
  XOR2_X1 U636 ( .A(G162GAT), .B(n570), .Z(G1347GAT) );
  AND2_X1 U637 ( .A1(n572), .A2(n571), .ZN(n573) );
  XOR2_X1 U638 ( .A(G169GAT), .B(n573), .Z(G1348GAT) );
  NOR2_X1 U639 ( .A1(n587), .A2(n574), .ZN(n576) );
  XNOR2_X1 U640 ( .A(G183GAT), .B(KEYINPUT125), .ZN(n575) );
  XNOR2_X1 U641 ( .A(n576), .B(n575), .ZN(G1350GAT) );
  NAND2_X1 U642 ( .A1(n577), .A2(n578), .ZN(n589) );
  NOR2_X1 U643 ( .A1(n579), .A2(n589), .ZN(n581) );
  XNOR2_X1 U644 ( .A(KEYINPUT60), .B(KEYINPUT59), .ZN(n580) );
  XNOR2_X1 U645 ( .A(n581), .B(n580), .ZN(n582) );
  XNOR2_X1 U646 ( .A(G197GAT), .B(n582), .ZN(G1352GAT) );
  NOR2_X1 U647 ( .A1(n583), .A2(n589), .ZN(n585) );
  XNOR2_X1 U648 ( .A(KEYINPUT61), .B(KEYINPUT127), .ZN(n584) );
  XNOR2_X1 U649 ( .A(n585), .B(n584), .ZN(n586) );
  XOR2_X1 U650 ( .A(G204GAT), .B(n586), .Z(G1353GAT) );
  NOR2_X1 U651 ( .A1(n587), .A2(n589), .ZN(n588) );
  XOR2_X1 U652 ( .A(G211GAT), .B(n588), .Z(G1354GAT) );
  NOR2_X1 U653 ( .A1(n498), .A2(n589), .ZN(n590) );
  XOR2_X1 U654 ( .A(KEYINPUT62), .B(n590), .Z(n591) );
  XNOR2_X1 U655 ( .A(G218GAT), .B(n591), .ZN(G1355GAT) );
endmodule

