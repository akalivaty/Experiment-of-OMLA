//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 1 0 0 0 1 0 0 0 1 1 1 1 0 0 0 0 1 1 0 1 1 0 1 0 0 1 1 0 1 1 1 0 0 1 0 1 0 1 1 0 0 0 0 0 1 1 0 0 0 1 0 1 0 1 0 1 1 0 1 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:22:34 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n695, new_n696,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n705,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n714,
    new_n715, new_n716, new_n717, new_n718, new_n719, new_n720, new_n721,
    new_n722, new_n723, new_n724, new_n725, new_n726, new_n727, new_n728,
    new_n729, new_n730, new_n731, new_n733, new_n734, new_n735, new_n736,
    new_n737, new_n738, new_n739, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n760, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n782,
    new_n783, new_n784, new_n785, new_n786, new_n787, new_n788, new_n789,
    new_n790, new_n791, new_n792, new_n793, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n914, new_n915, new_n916, new_n917,
    new_n918, new_n919, new_n920, new_n921, new_n922, new_n924, new_n925,
    new_n926, new_n927, new_n929, new_n930, new_n931, new_n933, new_n934,
    new_n935, new_n936, new_n937, new_n938, new_n939, new_n940, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n951, new_n952, new_n953, new_n954, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007;
  INV_X1    g000(.A(G217), .ZN(new_n187));
  INV_X1    g001(.A(G902), .ZN(new_n188));
  AOI21_X1  g002(.A(new_n187), .B1(G234), .B2(new_n188), .ZN(new_n189));
  INV_X1    g003(.A(G140), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n190), .A2(G125), .ZN(new_n191));
  INV_X1    g005(.A(G125), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n192), .A2(G140), .ZN(new_n193));
  INV_X1    g007(.A(KEYINPUT75), .ZN(new_n194));
  NAND4_X1  g008(.A1(new_n191), .A2(new_n193), .A3(new_n194), .A4(KEYINPUT16), .ZN(new_n195));
  AND3_X1   g009(.A1(new_n191), .A2(new_n193), .A3(KEYINPUT16), .ZN(new_n196));
  OAI21_X1  g010(.A(KEYINPUT75), .B1(new_n191), .B2(KEYINPUT16), .ZN(new_n197));
  OAI21_X1  g011(.A(new_n195), .B1(new_n196), .B2(new_n197), .ZN(new_n198));
  OR2_X1    g012(.A1(new_n198), .A2(G146), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n198), .A2(G146), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n199), .A2(new_n200), .ZN(new_n201));
  XOR2_X1   g015(.A(G119), .B(G128), .Z(new_n202));
  XNOR2_X1  g016(.A(KEYINPUT24), .B(G110), .ZN(new_n203));
  NOR2_X1   g017(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  INV_X1    g018(.A(G119), .ZN(new_n205));
  OAI21_X1  g019(.A(KEYINPUT74), .B1(new_n205), .B2(G128), .ZN(new_n206));
  AOI22_X1  g020(.A1(new_n206), .A2(KEYINPUT23), .B1(new_n205), .B2(G128), .ZN(new_n207));
  OAI21_X1  g021(.A(new_n207), .B1(KEYINPUT23), .B2(new_n206), .ZN(new_n208));
  AOI21_X1  g022(.A(new_n204), .B1(new_n208), .B2(G110), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n201), .A2(new_n209), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n202), .A2(new_n203), .ZN(new_n211));
  OAI21_X1  g025(.A(new_n211), .B1(new_n208), .B2(G110), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n191), .A2(new_n193), .ZN(new_n213));
  NOR2_X1   g027(.A1(new_n213), .A2(G146), .ZN(new_n214));
  AOI21_X1  g028(.A(new_n214), .B1(new_n198), .B2(G146), .ZN(new_n215));
  INV_X1    g029(.A(KEYINPUT76), .ZN(new_n216));
  NAND3_X1  g030(.A1(new_n212), .A2(new_n215), .A3(new_n216), .ZN(new_n217));
  INV_X1    g031(.A(new_n217), .ZN(new_n218));
  AOI21_X1  g032(.A(new_n216), .B1(new_n212), .B2(new_n215), .ZN(new_n219));
  OAI21_X1  g033(.A(new_n210), .B1(new_n218), .B2(new_n219), .ZN(new_n220));
  XNOR2_X1  g034(.A(KEYINPUT22), .B(G137), .ZN(new_n221));
  INV_X1    g035(.A(G953), .ZN(new_n222));
  AND3_X1   g036(.A1(new_n222), .A2(G221), .A3(G234), .ZN(new_n223));
  XOR2_X1   g037(.A(new_n221), .B(new_n223), .Z(new_n224));
  NAND2_X1  g038(.A1(new_n220), .A2(new_n224), .ZN(new_n225));
  INV_X1    g039(.A(new_n219), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n226), .A2(new_n217), .ZN(new_n227));
  AOI21_X1  g041(.A(KEYINPUT77), .B1(new_n227), .B2(new_n210), .ZN(new_n228));
  OAI211_X1 g042(.A(new_n210), .B(KEYINPUT77), .C1(new_n218), .C2(new_n219), .ZN(new_n229));
  INV_X1    g043(.A(new_n229), .ZN(new_n230));
  NOR2_X1   g044(.A1(new_n228), .A2(new_n230), .ZN(new_n231));
  OAI21_X1  g045(.A(new_n225), .B1(new_n231), .B2(new_n224), .ZN(new_n232));
  AOI21_X1  g046(.A(KEYINPUT25), .B1(new_n232), .B2(new_n188), .ZN(new_n233));
  INV_X1    g047(.A(KEYINPUT77), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n220), .A2(new_n234), .ZN(new_n235));
  AOI21_X1  g049(.A(new_n224), .B1(new_n235), .B2(new_n229), .ZN(new_n236));
  INV_X1    g050(.A(new_n225), .ZN(new_n237));
  OAI211_X1 g051(.A(KEYINPUT25), .B(new_n188), .C1(new_n236), .C2(new_n237), .ZN(new_n238));
  INV_X1    g052(.A(new_n238), .ZN(new_n239));
  OAI21_X1  g053(.A(new_n189), .B1(new_n233), .B2(new_n239), .ZN(new_n240));
  NOR2_X1   g054(.A1(new_n189), .A2(G902), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n232), .A2(new_n241), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n240), .A2(new_n242), .ZN(new_n243));
  NOR2_X1   g057(.A1(G472), .A2(G902), .ZN(new_n244));
  INV_X1    g058(.A(G137), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n245), .A2(KEYINPUT65), .ZN(new_n246));
  INV_X1    g060(.A(KEYINPUT65), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n247), .A2(G137), .ZN(new_n248));
  AOI21_X1  g062(.A(G134), .B1(new_n246), .B2(new_n248), .ZN(new_n249));
  INV_X1    g063(.A(KEYINPUT66), .ZN(new_n250));
  INV_X1    g064(.A(G134), .ZN(new_n251));
  OAI21_X1  g065(.A(new_n250), .B1(new_n251), .B2(G137), .ZN(new_n252));
  NAND3_X1  g066(.A1(new_n245), .A2(KEYINPUT66), .A3(G134), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n252), .A2(new_n253), .ZN(new_n254));
  OAI21_X1  g068(.A(G131), .B1(new_n249), .B2(new_n254), .ZN(new_n255));
  INV_X1    g069(.A(G146), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n256), .A2(G143), .ZN(new_n257));
  INV_X1    g071(.A(G143), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n258), .A2(G146), .ZN(new_n259));
  INV_X1    g073(.A(G128), .ZN(new_n260));
  OAI211_X1 g074(.A(new_n257), .B(new_n259), .C1(KEYINPUT1), .C2(new_n260), .ZN(new_n261));
  OAI21_X1  g075(.A(KEYINPUT1), .B1(new_n258), .B2(G146), .ZN(new_n262));
  NOR2_X1   g076(.A1(new_n258), .A2(G146), .ZN(new_n263));
  NOR2_X1   g077(.A1(new_n256), .A2(G143), .ZN(new_n264));
  OAI211_X1 g078(.A(G128), .B(new_n262), .C1(new_n263), .C2(new_n264), .ZN(new_n265));
  AND2_X1   g079(.A1(KEYINPUT11), .A2(G134), .ZN(new_n266));
  NAND3_X1  g080(.A1(new_n246), .A2(new_n248), .A3(new_n266), .ZN(new_n267));
  AOI21_X1  g081(.A(KEYINPUT11), .B1(new_n245), .B2(G134), .ZN(new_n268));
  INV_X1    g082(.A(new_n268), .ZN(new_n269));
  AOI21_X1  g083(.A(G131), .B1(new_n251), .B2(G137), .ZN(new_n270));
  NAND3_X1  g084(.A1(new_n267), .A2(new_n269), .A3(new_n270), .ZN(new_n271));
  NAND4_X1  g085(.A1(new_n255), .A2(new_n261), .A3(new_n265), .A4(new_n271), .ZN(new_n272));
  AND2_X1   g086(.A1(KEYINPUT0), .A2(G128), .ZN(new_n273));
  NAND3_X1  g087(.A1(new_n257), .A2(new_n259), .A3(new_n273), .ZN(new_n274));
  XNOR2_X1  g088(.A(G143), .B(G146), .ZN(new_n275));
  XNOR2_X1  g089(.A(KEYINPUT0), .B(G128), .ZN(new_n276));
  OAI21_X1  g090(.A(new_n274), .B1(new_n275), .B2(new_n276), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n277), .A2(KEYINPUT64), .ZN(new_n278));
  INV_X1    g092(.A(KEYINPUT64), .ZN(new_n279));
  OAI211_X1 g093(.A(new_n274), .B(new_n279), .C1(new_n275), .C2(new_n276), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n278), .A2(new_n280), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n251), .A2(G137), .ZN(new_n282));
  NAND3_X1  g096(.A1(new_n267), .A2(new_n269), .A3(new_n282), .ZN(new_n283));
  XNOR2_X1  g097(.A(KEYINPUT65), .B(G137), .ZN(new_n284));
  AOI21_X1  g098(.A(new_n268), .B1(new_n284), .B2(new_n266), .ZN(new_n285));
  AOI22_X1  g099(.A1(G131), .A2(new_n283), .B1(new_n285), .B2(new_n270), .ZN(new_n286));
  OAI21_X1  g100(.A(new_n272), .B1(new_n281), .B2(new_n286), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n205), .A2(G116), .ZN(new_n288));
  INV_X1    g102(.A(G116), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n289), .A2(G119), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n288), .A2(new_n290), .ZN(new_n291));
  XNOR2_X1  g105(.A(KEYINPUT2), .B(G113), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  INV_X1    g107(.A(G113), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n294), .A2(KEYINPUT2), .ZN(new_n295));
  INV_X1    g109(.A(KEYINPUT2), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n296), .A2(G113), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n295), .A2(new_n297), .ZN(new_n298));
  XNOR2_X1  g112(.A(G116), .B(G119), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n298), .A2(new_n299), .ZN(new_n300));
  INV_X1    g114(.A(KEYINPUT67), .ZN(new_n301));
  NAND3_X1  g115(.A1(new_n293), .A2(new_n300), .A3(new_n301), .ZN(new_n302));
  NAND3_X1  g116(.A1(new_n291), .A2(new_n292), .A3(KEYINPUT67), .ZN(new_n303));
  AND2_X1   g117(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n287), .A2(new_n304), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n302), .A2(new_n303), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n272), .A2(new_n306), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n283), .A2(G131), .ZN(new_n308));
  AOI21_X1  g122(.A(new_n277), .B1(new_n308), .B2(new_n271), .ZN(new_n309));
  OAI21_X1  g123(.A(KEYINPUT68), .B1(new_n307), .B2(new_n309), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n308), .A2(new_n271), .ZN(new_n311));
  INV_X1    g125(.A(new_n277), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  INV_X1    g127(.A(KEYINPUT68), .ZN(new_n314));
  NAND4_X1  g128(.A1(new_n313), .A2(new_n314), .A3(new_n272), .A4(new_n306), .ZN(new_n315));
  NAND3_X1  g129(.A1(new_n305), .A2(new_n310), .A3(new_n315), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n316), .A2(KEYINPUT28), .ZN(new_n317));
  NOR2_X1   g131(.A1(new_n307), .A2(new_n309), .ZN(new_n318));
  NOR2_X1   g132(.A1(new_n318), .A2(KEYINPUT28), .ZN(new_n319));
  INV_X1    g133(.A(new_n319), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n317), .A2(new_n320), .ZN(new_n321));
  XOR2_X1   g135(.A(KEYINPUT69), .B(KEYINPUT27), .Z(new_n322));
  INV_X1    g136(.A(G237), .ZN(new_n323));
  NAND3_X1  g137(.A1(new_n323), .A2(new_n222), .A3(G210), .ZN(new_n324));
  XNOR2_X1  g138(.A(new_n322), .B(new_n324), .ZN(new_n325));
  XNOR2_X1  g139(.A(KEYINPUT26), .B(G101), .ZN(new_n326));
  XNOR2_X1  g140(.A(new_n325), .B(new_n326), .ZN(new_n327));
  INV_X1    g141(.A(new_n327), .ZN(new_n328));
  AOI21_X1  g142(.A(KEYINPUT71), .B1(new_n321), .B2(new_n328), .ZN(new_n329));
  AOI21_X1  g143(.A(new_n319), .B1(new_n316), .B2(KEYINPUT28), .ZN(new_n330));
  INV_X1    g144(.A(KEYINPUT71), .ZN(new_n331));
  NOR3_X1   g145(.A1(new_n330), .A2(new_n331), .A3(new_n327), .ZN(new_n332));
  NOR2_X1   g146(.A1(new_n329), .A2(new_n332), .ZN(new_n333));
  NAND3_X1  g147(.A1(new_n310), .A2(new_n315), .A3(new_n327), .ZN(new_n334));
  INV_X1    g148(.A(new_n272), .ZN(new_n335));
  OAI21_X1  g149(.A(KEYINPUT30), .B1(new_n335), .B2(new_n309), .ZN(new_n336));
  INV_X1    g150(.A(KEYINPUT30), .ZN(new_n337));
  OAI211_X1 g151(.A(new_n337), .B(new_n272), .C1(new_n281), .C2(new_n286), .ZN(new_n338));
  AOI21_X1  g152(.A(new_n306), .B1(new_n336), .B2(new_n338), .ZN(new_n339));
  OAI21_X1  g153(.A(KEYINPUT31), .B1(new_n334), .B2(new_n339), .ZN(new_n340));
  NOR3_X1   g154(.A1(new_n334), .A2(new_n339), .A3(KEYINPUT31), .ZN(new_n341));
  INV_X1    g155(.A(KEYINPUT70), .ZN(new_n342));
  OAI21_X1  g156(.A(new_n340), .B1(new_n341), .B2(new_n342), .ZN(new_n343));
  INV_X1    g157(.A(new_n334), .ZN(new_n344));
  INV_X1    g158(.A(new_n339), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n344), .A2(new_n345), .ZN(new_n346));
  NAND3_X1  g160(.A1(new_n346), .A2(KEYINPUT70), .A3(KEYINPUT31), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n343), .A2(new_n347), .ZN(new_n348));
  OAI21_X1  g162(.A(new_n244), .B1(new_n333), .B2(new_n348), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n349), .A2(KEYINPUT72), .ZN(new_n350));
  INV_X1    g164(.A(KEYINPUT32), .ZN(new_n351));
  OAI211_X1 g165(.A(new_n343), .B(new_n347), .C1(new_n329), .C2(new_n332), .ZN(new_n352));
  INV_X1    g166(.A(KEYINPUT72), .ZN(new_n353));
  NAND3_X1  g167(.A1(new_n352), .A2(new_n353), .A3(new_n244), .ZN(new_n354));
  NAND3_X1  g168(.A1(new_n350), .A2(new_n351), .A3(new_n354), .ZN(new_n355));
  INV_X1    g169(.A(new_n244), .ZN(new_n356));
  AND2_X1   g170(.A1(new_n343), .A2(new_n347), .ZN(new_n357));
  INV_X1    g171(.A(new_n332), .ZN(new_n358));
  OAI21_X1  g172(.A(new_n331), .B1(new_n330), .B2(new_n327), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n358), .A2(new_n359), .ZN(new_n360));
  AOI21_X1  g174(.A(new_n356), .B1(new_n357), .B2(new_n360), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n310), .A2(new_n315), .ZN(new_n362));
  OAI21_X1  g176(.A(new_n328), .B1(new_n339), .B2(new_n362), .ZN(new_n363));
  INV_X1    g177(.A(KEYINPUT73), .ZN(new_n364));
  XNOR2_X1  g178(.A(new_n363), .B(new_n364), .ZN(new_n365));
  AOI21_X1  g179(.A(KEYINPUT29), .B1(new_n330), .B2(new_n327), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n365), .A2(new_n366), .ZN(new_n367));
  OAI21_X1  g181(.A(new_n304), .B1(new_n335), .B2(new_n309), .ZN(new_n368));
  NAND3_X1  g182(.A1(new_n310), .A2(new_n315), .A3(new_n368), .ZN(new_n369));
  AOI21_X1  g183(.A(new_n319), .B1(new_n369), .B2(KEYINPUT28), .ZN(new_n370));
  AND2_X1   g184(.A1(new_n327), .A2(KEYINPUT29), .ZN(new_n371));
  AOI21_X1  g185(.A(G902), .B1(new_n370), .B2(new_n371), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n367), .A2(new_n372), .ZN(new_n373));
  AOI22_X1  g187(.A1(new_n361), .A2(KEYINPUT32), .B1(new_n373), .B2(G472), .ZN(new_n374));
  AOI21_X1  g188(.A(new_n243), .B1(new_n355), .B2(new_n374), .ZN(new_n375));
  OAI21_X1  g189(.A(G214), .B1(G237), .B2(G902), .ZN(new_n376));
  INV_X1    g190(.A(new_n376), .ZN(new_n377));
  OAI21_X1  g191(.A(G210), .B1(G237), .B2(G902), .ZN(new_n378));
  XOR2_X1   g192(.A(new_n378), .B(KEYINPUT85), .Z(new_n379));
  INV_X1    g193(.A(new_n379), .ZN(new_n380));
  INV_X1    g194(.A(KEYINPUT4), .ZN(new_n381));
  INV_X1    g195(.A(G107), .ZN(new_n382));
  NOR2_X1   g196(.A1(new_n382), .A2(G104), .ZN(new_n383));
  INV_X1    g197(.A(KEYINPUT3), .ZN(new_n384));
  INV_X1    g198(.A(G104), .ZN(new_n385));
  OAI21_X1  g199(.A(new_n384), .B1(new_n385), .B2(G107), .ZN(new_n386));
  NAND3_X1  g200(.A1(new_n382), .A2(KEYINPUT3), .A3(G104), .ZN(new_n387));
  AOI21_X1  g201(.A(new_n383), .B1(new_n386), .B2(new_n387), .ZN(new_n388));
  INV_X1    g202(.A(G101), .ZN(new_n389));
  AOI21_X1  g203(.A(new_n381), .B1(new_n388), .B2(new_n389), .ZN(new_n390));
  INV_X1    g204(.A(KEYINPUT78), .ZN(new_n391));
  OAI21_X1  g205(.A(G101), .B1(new_n388), .B2(new_n391), .ZN(new_n392));
  AOI211_X1 g206(.A(KEYINPUT78), .B(new_n383), .C1(new_n386), .C2(new_n387), .ZN(new_n393));
  OAI21_X1  g207(.A(new_n390), .B1(new_n392), .B2(new_n393), .ZN(new_n394));
  AND3_X1   g208(.A1(new_n382), .A2(KEYINPUT3), .A3(G104), .ZN(new_n395));
  AOI21_X1  g209(.A(KEYINPUT3), .B1(new_n382), .B2(G104), .ZN(new_n396));
  OAI22_X1  g210(.A1(new_n395), .A2(new_n396), .B1(G104), .B2(new_n382), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n397), .A2(KEYINPUT78), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n388), .A2(new_n391), .ZN(new_n399));
  NAND4_X1  g213(.A1(new_n398), .A2(new_n381), .A3(new_n399), .A4(G101), .ZN(new_n400));
  NAND3_X1  g214(.A1(new_n304), .A2(new_n394), .A3(new_n400), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n382), .A2(G104), .ZN(new_n402));
  INV_X1    g216(.A(KEYINPUT79), .ZN(new_n403));
  OAI21_X1  g217(.A(new_n402), .B1(new_n383), .B2(new_n403), .ZN(new_n404));
  NOR3_X1   g218(.A1(new_n382), .A2(KEYINPUT79), .A3(G104), .ZN(new_n405));
  OAI21_X1  g219(.A(G101), .B1(new_n404), .B2(new_n405), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n388), .A2(new_n389), .ZN(new_n407));
  INV_X1    g221(.A(KEYINPUT5), .ZN(new_n408));
  NAND3_X1  g222(.A1(new_n408), .A2(new_n205), .A3(G116), .ZN(new_n409));
  OAI211_X1 g223(.A(G113), .B(new_n409), .C1(new_n291), .C2(new_n408), .ZN(new_n410));
  NAND4_X1  g224(.A1(new_n406), .A2(new_n407), .A3(new_n410), .A4(new_n300), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n401), .A2(new_n411), .ZN(new_n412));
  XNOR2_X1  g226(.A(G110), .B(G122), .ZN(new_n413));
  INV_X1    g227(.A(new_n413), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n412), .A2(new_n414), .ZN(new_n415));
  NAND3_X1  g229(.A1(new_n401), .A2(new_n413), .A3(new_n411), .ZN(new_n416));
  NAND3_X1  g230(.A1(new_n415), .A2(KEYINPUT6), .A3(new_n416), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n265), .A2(new_n261), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n418), .A2(new_n192), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n277), .A2(G125), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  INV_X1    g235(.A(G224), .ZN(new_n422));
  NOR2_X1   g236(.A1(new_n422), .A2(G953), .ZN(new_n423));
  XNOR2_X1  g237(.A(new_n421), .B(new_n423), .ZN(new_n424));
  INV_X1    g238(.A(KEYINPUT6), .ZN(new_n425));
  NAND3_X1  g239(.A1(new_n412), .A2(new_n425), .A3(new_n414), .ZN(new_n426));
  NAND3_X1  g240(.A1(new_n417), .A2(new_n424), .A3(new_n426), .ZN(new_n427));
  INV_X1    g241(.A(KEYINPUT80), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n427), .A2(new_n428), .ZN(new_n429));
  NAND4_X1  g243(.A1(new_n417), .A2(KEYINPUT80), .A3(new_n424), .A4(new_n426), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n429), .A2(new_n430), .ZN(new_n431));
  XNOR2_X1  g245(.A(KEYINPUT81), .B(KEYINPUT8), .ZN(new_n432));
  XNOR2_X1  g246(.A(new_n413), .B(new_n432), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n406), .A2(new_n407), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n410), .A2(new_n300), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  AOI21_X1  g250(.A(new_n433), .B1(new_n436), .B2(new_n411), .ZN(new_n437));
  OAI21_X1  g251(.A(KEYINPUT7), .B1(new_n422), .B2(G953), .ZN(new_n438));
  INV_X1    g252(.A(new_n438), .ZN(new_n439));
  AND4_X1   g253(.A1(KEYINPUT83), .A2(new_n419), .A3(new_n420), .A4(new_n439), .ZN(new_n440));
  NOR2_X1   g254(.A1(new_n437), .A2(new_n440), .ZN(new_n441));
  INV_X1    g255(.A(KEYINPUT83), .ZN(new_n442));
  INV_X1    g256(.A(KEYINPUT82), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n419), .A2(new_n443), .ZN(new_n444));
  NAND3_X1  g258(.A1(new_n418), .A2(KEYINPUT82), .A3(new_n192), .ZN(new_n445));
  NAND3_X1  g259(.A1(new_n444), .A2(new_n420), .A3(new_n445), .ZN(new_n446));
  AOI21_X1  g260(.A(new_n442), .B1(new_n446), .B2(new_n438), .ZN(new_n447));
  NOR2_X1   g261(.A1(new_n421), .A2(new_n438), .ZN(new_n448));
  OAI211_X1 g262(.A(new_n416), .B(new_n441), .C1(new_n447), .C2(new_n448), .ZN(new_n449));
  AND3_X1   g263(.A1(new_n449), .A2(KEYINPUT84), .A3(new_n188), .ZN(new_n450));
  AOI21_X1  g264(.A(KEYINPUT84), .B1(new_n449), .B2(new_n188), .ZN(new_n451));
  NOR2_X1   g265(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  AOI21_X1  g266(.A(new_n380), .B1(new_n431), .B2(new_n452), .ZN(new_n453));
  INV_X1    g267(.A(KEYINPUT86), .ZN(new_n454));
  XNOR2_X1  g268(.A(new_n453), .B(new_n454), .ZN(new_n455));
  NAND3_X1  g269(.A1(new_n431), .A2(new_n452), .A3(new_n380), .ZN(new_n456));
  INV_X1    g270(.A(KEYINPUT87), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  NAND4_X1  g272(.A1(new_n431), .A2(new_n452), .A3(KEYINPUT87), .A4(new_n380), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  AOI21_X1  g274(.A(new_n377), .B1(new_n455), .B2(new_n460), .ZN(new_n461));
  INV_X1    g275(.A(KEYINPUT13), .ZN(new_n462));
  INV_X1    g276(.A(KEYINPUT94), .ZN(new_n463));
  AOI21_X1  g277(.A(new_n463), .B1(G128), .B2(new_n258), .ZN(new_n464));
  NOR3_X1   g278(.A1(new_n260), .A2(KEYINPUT94), .A3(G143), .ZN(new_n465));
  OAI21_X1  g279(.A(new_n462), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  OAI21_X1  g280(.A(KEYINPUT94), .B1(new_n260), .B2(G143), .ZN(new_n467));
  NAND3_X1  g281(.A1(new_n463), .A2(new_n258), .A3(G128), .ZN(new_n468));
  NAND3_X1  g282(.A1(new_n467), .A2(new_n468), .A3(KEYINPUT13), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n260), .A2(G143), .ZN(new_n470));
  NAND3_X1  g284(.A1(new_n466), .A2(new_n469), .A3(new_n470), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n471), .A2(G134), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n467), .A2(new_n468), .ZN(new_n473));
  NAND3_X1  g287(.A1(new_n473), .A2(new_n251), .A3(new_n470), .ZN(new_n474));
  XNOR2_X1  g288(.A(G116), .B(G122), .ZN(new_n475));
  INV_X1    g289(.A(KEYINPUT93), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  INV_X1    g291(.A(new_n477), .ZN(new_n478));
  NOR2_X1   g292(.A1(new_n475), .A2(new_n476), .ZN(new_n479));
  NOR3_X1   g293(.A1(new_n478), .A2(new_n479), .A3(new_n382), .ZN(new_n480));
  XOR2_X1   g294(.A(G116), .B(G122), .Z(new_n481));
  NAND2_X1  g295(.A1(new_n481), .A2(KEYINPUT93), .ZN(new_n482));
  AOI21_X1  g296(.A(G107), .B1(new_n482), .B2(new_n477), .ZN(new_n483));
  OAI211_X1 g297(.A(new_n472), .B(new_n474), .C1(new_n480), .C2(new_n483), .ZN(new_n484));
  OAI21_X1  g298(.A(new_n382), .B1(new_n478), .B2(new_n479), .ZN(new_n485));
  NAND3_X1  g299(.A1(new_n289), .A2(KEYINPUT14), .A3(G122), .ZN(new_n486));
  OAI211_X1 g300(.A(G107), .B(new_n486), .C1(new_n481), .C2(KEYINPUT14), .ZN(new_n487));
  INV_X1    g301(.A(new_n474), .ZN(new_n488));
  AOI21_X1  g302(.A(new_n251), .B1(new_n473), .B2(new_n470), .ZN(new_n489));
  OAI211_X1 g303(.A(new_n485), .B(new_n487), .C1(new_n488), .C2(new_n489), .ZN(new_n490));
  XNOR2_X1  g304(.A(KEYINPUT9), .B(G234), .ZN(new_n491));
  NOR3_X1   g305(.A1(new_n491), .A2(new_n187), .A3(G953), .ZN(new_n492));
  NAND3_X1  g306(.A1(new_n484), .A2(new_n490), .A3(new_n492), .ZN(new_n493));
  INV_X1    g307(.A(new_n493), .ZN(new_n494));
  AOI21_X1  g308(.A(new_n492), .B1(new_n484), .B2(new_n490), .ZN(new_n495));
  OAI21_X1  g309(.A(new_n188), .B1(new_n494), .B2(new_n495), .ZN(new_n496));
  INV_X1    g310(.A(KEYINPUT95), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n484), .A2(new_n490), .ZN(new_n499));
  INV_X1    g313(.A(new_n492), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  AOI21_X1  g315(.A(G902), .B1(new_n501), .B2(new_n493), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n502), .A2(KEYINPUT95), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n498), .A2(new_n503), .ZN(new_n504));
  INV_X1    g318(.A(KEYINPUT15), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n505), .A2(G478), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n504), .A2(new_n506), .ZN(new_n507));
  AOI21_X1  g321(.A(new_n506), .B1(new_n502), .B2(KEYINPUT95), .ZN(new_n508));
  INV_X1    g322(.A(new_n508), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n507), .A2(new_n509), .ZN(new_n510));
  AND3_X1   g324(.A1(new_n323), .A2(new_n222), .A3(G214), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n258), .A2(KEYINPUT88), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  XNOR2_X1  g327(.A(KEYINPUT88), .B(G143), .ZN(new_n514));
  OAI21_X1  g328(.A(new_n513), .B1(new_n511), .B2(new_n514), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n515), .A2(G131), .ZN(new_n516));
  INV_X1    g330(.A(KEYINPUT17), .ZN(new_n517));
  INV_X1    g331(.A(G131), .ZN(new_n518));
  OAI211_X1 g332(.A(new_n513), .B(new_n518), .C1(new_n511), .C2(new_n514), .ZN(new_n519));
  NAND3_X1  g333(.A1(new_n516), .A2(new_n517), .A3(new_n519), .ZN(new_n520));
  NAND3_X1  g334(.A1(new_n515), .A2(KEYINPUT17), .A3(G131), .ZN(new_n521));
  NAND4_X1  g335(.A1(new_n520), .A2(new_n200), .A3(new_n199), .A4(new_n521), .ZN(new_n522));
  AND2_X1   g336(.A1(new_n511), .A2(new_n512), .ZN(new_n523));
  NOR2_X1   g337(.A1(new_n514), .A2(new_n511), .ZN(new_n524));
  NOR2_X1   g338(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  NAND2_X1  g339(.A1(KEYINPUT18), .A2(G131), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n213), .A2(KEYINPUT90), .ZN(new_n527));
  INV_X1    g341(.A(KEYINPUT90), .ZN(new_n528));
  NAND3_X1  g342(.A1(new_n191), .A2(new_n193), .A3(new_n528), .ZN(new_n529));
  NAND3_X1  g343(.A1(new_n527), .A2(G146), .A3(new_n529), .ZN(new_n530));
  INV_X1    g344(.A(new_n214), .ZN(new_n531));
  AOI22_X1  g345(.A1(new_n525), .A2(new_n526), .B1(new_n530), .B2(new_n531), .ZN(new_n532));
  INV_X1    g346(.A(new_n526), .ZN(new_n533));
  NAND3_X1  g347(.A1(new_n515), .A2(KEYINPUT89), .A3(new_n533), .ZN(new_n534));
  INV_X1    g348(.A(new_n534), .ZN(new_n535));
  AOI21_X1  g349(.A(KEYINPUT89), .B1(new_n515), .B2(new_n533), .ZN(new_n536));
  OAI21_X1  g350(.A(new_n532), .B1(new_n535), .B2(new_n536), .ZN(new_n537));
  XNOR2_X1  g351(.A(G113), .B(G122), .ZN(new_n538));
  XNOR2_X1  g352(.A(new_n538), .B(new_n385), .ZN(new_n539));
  AND3_X1   g353(.A1(new_n522), .A2(new_n537), .A3(new_n539), .ZN(new_n540));
  AOI21_X1  g354(.A(new_n539), .B1(new_n522), .B2(new_n537), .ZN(new_n541));
  OAI21_X1  g355(.A(new_n188), .B1(new_n540), .B2(new_n541), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n542), .A2(G475), .ZN(new_n543));
  NAND3_X1  g357(.A1(new_n522), .A2(new_n537), .A3(new_n539), .ZN(new_n544));
  INV_X1    g358(.A(new_n536), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n545), .A2(new_n534), .ZN(new_n546));
  AOI22_X1  g360(.A1(new_n516), .A2(new_n519), .B1(G146), .B2(new_n198), .ZN(new_n547));
  NAND3_X1  g361(.A1(new_n527), .A2(KEYINPUT19), .A3(new_n529), .ZN(new_n548));
  INV_X1    g362(.A(KEYINPUT91), .ZN(new_n549));
  OR3_X1    g363(.A1(new_n213), .A2(new_n549), .A3(KEYINPUT19), .ZN(new_n550));
  OAI21_X1  g364(.A(new_n549), .B1(new_n213), .B2(KEYINPUT19), .ZN(new_n551));
  NAND4_X1  g365(.A1(new_n548), .A2(new_n550), .A3(new_n256), .A4(new_n551), .ZN(new_n552));
  AOI22_X1  g366(.A1(new_n546), .A2(new_n532), .B1(new_n547), .B2(new_n552), .ZN(new_n553));
  OAI21_X1  g367(.A(new_n544), .B1(new_n553), .B2(new_n539), .ZN(new_n554));
  INV_X1    g368(.A(KEYINPUT92), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  INV_X1    g370(.A(KEYINPUT20), .ZN(new_n557));
  NOR2_X1   g371(.A1(G475), .A2(G902), .ZN(new_n558));
  AOI22_X1  g372(.A1(new_n556), .A2(new_n557), .B1(new_n554), .B2(new_n558), .ZN(new_n559));
  NAND4_X1  g373(.A1(new_n554), .A2(KEYINPUT92), .A3(new_n557), .A4(new_n558), .ZN(new_n560));
  INV_X1    g374(.A(new_n560), .ZN(new_n561));
  OAI21_X1  g375(.A(new_n543), .B1(new_n559), .B2(new_n561), .ZN(new_n562));
  INV_X1    g376(.A(G952), .ZN(new_n563));
  AOI211_X1 g377(.A(G953), .B(new_n563), .C1(G234), .C2(G237), .ZN(new_n564));
  AOI211_X1 g378(.A(new_n188), .B(new_n222), .C1(G234), .C2(G237), .ZN(new_n565));
  XNOR2_X1  g379(.A(KEYINPUT21), .B(G898), .ZN(new_n566));
  AOI21_X1  g380(.A(new_n564), .B1(new_n565), .B2(new_n566), .ZN(new_n567));
  NOR3_X1   g381(.A1(new_n510), .A2(new_n562), .A3(new_n567), .ZN(new_n568));
  OAI21_X1  g382(.A(G221), .B1(new_n491), .B2(G902), .ZN(new_n569));
  INV_X1    g383(.A(new_n569), .ZN(new_n570));
  NOR2_X1   g384(.A1(new_n434), .A2(new_n418), .ZN(new_n571));
  INV_X1    g385(.A(KEYINPUT10), .ZN(new_n572));
  XNOR2_X1  g386(.A(new_n571), .B(new_n572), .ZN(new_n573));
  NAND3_X1  g387(.A1(new_n394), .A2(new_n400), .A3(new_n312), .ZN(new_n574));
  AOI21_X1  g388(.A(new_n286), .B1(new_n573), .B2(new_n574), .ZN(new_n575));
  INV_X1    g389(.A(new_n575), .ZN(new_n576));
  NAND3_X1  g390(.A1(new_n573), .A2(new_n286), .A3(new_n574), .ZN(new_n577));
  XNOR2_X1  g391(.A(G110), .B(G140), .ZN(new_n578));
  AND2_X1   g392(.A1(new_n222), .A2(G227), .ZN(new_n579));
  XNOR2_X1  g393(.A(new_n578), .B(new_n579), .ZN(new_n580));
  INV_X1    g394(.A(new_n580), .ZN(new_n581));
  AND2_X1   g395(.A1(new_n577), .A2(new_n581), .ZN(new_n582));
  XNOR2_X1  g396(.A(new_n434), .B(new_n418), .ZN(new_n583));
  AND3_X1   g397(.A1(new_n583), .A2(KEYINPUT12), .A3(new_n311), .ZN(new_n584));
  AOI21_X1  g398(.A(KEYINPUT12), .B1(new_n583), .B2(new_n311), .ZN(new_n585));
  OAI21_X1  g399(.A(new_n577), .B1(new_n584), .B2(new_n585), .ZN(new_n586));
  AOI22_X1  g400(.A1(new_n576), .A2(new_n582), .B1(new_n586), .B2(new_n580), .ZN(new_n587));
  OAI21_X1  g401(.A(G469), .B1(new_n587), .B2(G902), .ZN(new_n588));
  AND3_X1   g402(.A1(new_n573), .A2(new_n286), .A3(new_n574), .ZN(new_n589));
  OAI21_X1  g403(.A(new_n580), .B1(new_n589), .B2(new_n575), .ZN(new_n590));
  OAI211_X1 g404(.A(new_n577), .B(new_n581), .C1(new_n584), .C2(new_n585), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  INV_X1    g406(.A(G469), .ZN(new_n593));
  NAND3_X1  g407(.A1(new_n592), .A2(new_n593), .A3(new_n188), .ZN(new_n594));
  AOI21_X1  g408(.A(new_n570), .B1(new_n588), .B2(new_n594), .ZN(new_n595));
  AND2_X1   g409(.A1(new_n568), .A2(new_n595), .ZN(new_n596));
  NAND3_X1  g410(.A1(new_n375), .A2(new_n461), .A3(new_n596), .ZN(new_n597));
  XNOR2_X1  g411(.A(KEYINPUT96), .B(G101), .ZN(new_n598));
  XNOR2_X1  g412(.A(new_n597), .B(new_n598), .ZN(G3));
  NAND2_X1  g413(.A1(new_n352), .A2(new_n188), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n600), .A2(G472), .ZN(new_n601));
  NAND3_X1  g415(.A1(new_n601), .A2(new_n350), .A3(new_n354), .ZN(new_n602));
  NAND3_X1  g416(.A1(new_n595), .A2(new_n240), .A3(new_n242), .ZN(new_n603));
  NOR2_X1   g417(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n547), .A2(new_n552), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n605), .A2(new_n537), .ZN(new_n606));
  INV_X1    g420(.A(new_n539), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  AOI21_X1  g422(.A(KEYINPUT92), .B1(new_n608), .B2(new_n544), .ZN(new_n609));
  AOI21_X1  g423(.A(new_n539), .B1(new_n605), .B2(new_n537), .ZN(new_n610));
  NOR2_X1   g424(.A1(new_n540), .A2(new_n610), .ZN(new_n611));
  INV_X1    g425(.A(new_n558), .ZN(new_n612));
  OAI22_X1  g426(.A1(new_n609), .A2(KEYINPUT20), .B1(new_n611), .B2(new_n612), .ZN(new_n613));
  AOI22_X1  g427(.A1(new_n613), .A2(new_n560), .B1(G475), .B2(new_n542), .ZN(new_n614));
  OR3_X1    g428(.A1(new_n494), .A2(KEYINPUT33), .A3(new_n495), .ZN(new_n615));
  OAI21_X1  g429(.A(KEYINPUT33), .B1(new_n494), .B2(new_n495), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n615), .A2(new_n616), .ZN(new_n617));
  AND2_X1   g431(.A1(new_n188), .A2(G478), .ZN(new_n618));
  INV_X1    g432(.A(KEYINPUT98), .ZN(new_n619));
  XOR2_X1   g433(.A(KEYINPUT97), .B(G478), .Z(new_n620));
  OAI21_X1  g434(.A(new_n619), .B1(new_n502), .B2(new_n620), .ZN(new_n621));
  INV_X1    g435(.A(new_n620), .ZN(new_n622));
  NAND3_X1  g436(.A1(new_n496), .A2(KEYINPUT98), .A3(new_n622), .ZN(new_n623));
  AOI22_X1  g437(.A1(new_n617), .A2(new_n618), .B1(new_n621), .B2(new_n623), .ZN(new_n624));
  NOR3_X1   g438(.A1(new_n614), .A2(new_n624), .A3(new_n567), .ZN(new_n625));
  AND3_X1   g439(.A1(new_n431), .A2(new_n452), .A3(new_n380), .ZN(new_n626));
  OAI211_X1 g440(.A(new_n625), .B(new_n376), .C1(new_n626), .C2(new_n453), .ZN(new_n627));
  INV_X1    g441(.A(new_n627), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n604), .A2(new_n628), .ZN(new_n629));
  XOR2_X1   g443(.A(KEYINPUT34), .B(G104), .Z(new_n630));
  XNOR2_X1  g444(.A(new_n629), .B(new_n630), .ZN(G6));
  AOI21_X1  g445(.A(new_n508), .B1(new_n504), .B2(new_n506), .ZN(new_n632));
  NOR3_X1   g446(.A1(new_n611), .A2(KEYINPUT20), .A3(new_n612), .ZN(new_n633));
  AOI21_X1  g447(.A(new_n557), .B1(new_n554), .B2(new_n558), .ZN(new_n634));
  OAI21_X1  g448(.A(new_n543), .B1(new_n633), .B2(new_n634), .ZN(new_n635));
  NOR3_X1   g449(.A1(new_n632), .A2(new_n635), .A3(new_n567), .ZN(new_n636));
  OAI211_X1 g450(.A(new_n636), .B(new_n376), .C1(new_n626), .C2(new_n453), .ZN(new_n637));
  INV_X1    g451(.A(new_n637), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n604), .A2(new_n638), .ZN(new_n639));
  XOR2_X1   g453(.A(KEYINPUT35), .B(G107), .Z(new_n640));
  XNOR2_X1  g454(.A(new_n639), .B(new_n640), .ZN(G9));
  INV_X1    g455(.A(KEYINPUT25), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n235), .A2(new_n229), .ZN(new_n643));
  INV_X1    g457(.A(new_n224), .ZN(new_n644));
  AOI21_X1  g458(.A(new_n237), .B1(new_n643), .B2(new_n644), .ZN(new_n645));
  OAI21_X1  g459(.A(new_n642), .B1(new_n645), .B2(G902), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n646), .A2(new_n238), .ZN(new_n647));
  NOR2_X1   g461(.A1(new_n644), .A2(KEYINPUT36), .ZN(new_n648));
  XNOR2_X1  g462(.A(new_n648), .B(KEYINPUT99), .ZN(new_n649));
  XNOR2_X1  g463(.A(new_n231), .B(new_n649), .ZN(new_n650));
  AOI22_X1  g464(.A1(new_n647), .A2(new_n189), .B1(new_n241), .B2(new_n650), .ZN(new_n651));
  NOR2_X1   g465(.A1(new_n602), .A2(new_n651), .ZN(new_n652));
  NAND3_X1  g466(.A1(new_n461), .A2(new_n652), .A3(new_n596), .ZN(new_n653));
  XNOR2_X1  g467(.A(new_n653), .B(KEYINPUT100), .ZN(new_n654));
  XNOR2_X1  g468(.A(KEYINPUT37), .B(G110), .ZN(new_n655));
  XNOR2_X1  g469(.A(new_n654), .B(new_n655), .ZN(G12));
  NAND2_X1  g470(.A1(new_n355), .A2(new_n374), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n431), .A2(new_n452), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n658), .A2(new_n379), .ZN(new_n659));
  AOI21_X1  g473(.A(new_n377), .B1(new_n659), .B2(new_n456), .ZN(new_n660));
  INV_X1    g474(.A(new_n564), .ZN(new_n661));
  INV_X1    g475(.A(new_n565), .ZN(new_n662));
  OAI21_X1  g476(.A(new_n661), .B1(new_n662), .B2(G900), .ZN(new_n663));
  OAI211_X1 g477(.A(new_n543), .B(new_n663), .C1(new_n633), .C2(new_n634), .ZN(new_n664));
  NOR2_X1   g478(.A1(new_n664), .A2(new_n632), .ZN(new_n665));
  INV_X1    g479(.A(new_n595), .ZN(new_n666));
  NOR2_X1   g480(.A1(new_n666), .A2(new_n651), .ZN(new_n667));
  NAND4_X1  g481(.A1(new_n657), .A2(new_n660), .A3(new_n665), .A4(new_n667), .ZN(new_n668));
  XNOR2_X1  g482(.A(new_n668), .B(G128), .ZN(G30));
  NAND2_X1  g483(.A1(new_n659), .A2(new_n454), .ZN(new_n670));
  NAND2_X1  g484(.A1(new_n453), .A2(KEYINPUT86), .ZN(new_n671));
  NAND3_X1  g485(.A1(new_n460), .A2(new_n670), .A3(new_n671), .ZN(new_n672));
  XNOR2_X1  g486(.A(new_n672), .B(KEYINPUT38), .ZN(new_n673));
  XNOR2_X1  g487(.A(KEYINPUT101), .B(KEYINPUT39), .ZN(new_n674));
  XNOR2_X1  g488(.A(new_n663), .B(new_n674), .ZN(new_n675));
  NAND2_X1  g489(.A1(new_n595), .A2(new_n675), .ZN(new_n676));
  XOR2_X1   g490(.A(new_n676), .B(KEYINPUT40), .Z(new_n677));
  NAND3_X1  g491(.A1(new_n352), .A2(KEYINPUT32), .A3(new_n244), .ZN(new_n678));
  INV_X1    g492(.A(G472), .ZN(new_n679));
  INV_X1    g493(.A(new_n369), .ZN(new_n680));
  OAI21_X1  g494(.A(new_n346), .B1(new_n327), .B2(new_n680), .ZN(new_n681));
  AND2_X1   g495(.A1(new_n681), .A2(new_n188), .ZN(new_n682));
  OAI211_X1 g496(.A(new_n355), .B(new_n678), .C1(new_n679), .C2(new_n682), .ZN(new_n683));
  NOR2_X1   g497(.A1(new_n614), .A2(new_n632), .ZN(new_n684));
  AND3_X1   g498(.A1(new_n651), .A2(new_n376), .A3(new_n684), .ZN(new_n685));
  NAND4_X1  g499(.A1(new_n673), .A2(new_n677), .A3(new_n683), .A4(new_n685), .ZN(new_n686));
  XNOR2_X1  g500(.A(new_n686), .B(G143), .ZN(G45));
  NAND2_X1  g501(.A1(new_n617), .A2(new_n618), .ZN(new_n688));
  NAND2_X1  g502(.A1(new_n621), .A2(new_n623), .ZN(new_n689));
  NAND2_X1  g503(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  NAND3_X1  g504(.A1(new_n562), .A2(new_n690), .A3(new_n663), .ZN(new_n691));
  INV_X1    g505(.A(KEYINPUT102), .ZN(new_n692));
  NAND2_X1  g506(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  NAND4_X1  g507(.A1(new_n562), .A2(new_n690), .A3(KEYINPUT102), .A4(new_n663), .ZN(new_n694));
  AND2_X1   g508(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  NAND4_X1  g509(.A1(new_n657), .A2(new_n660), .A3(new_n667), .A4(new_n695), .ZN(new_n696));
  XNOR2_X1  g510(.A(new_n696), .B(G146), .ZN(G48));
  INV_X1    g511(.A(new_n243), .ZN(new_n698));
  AOI21_X1  g512(.A(new_n593), .B1(new_n592), .B2(new_n188), .ZN(new_n699));
  AOI211_X1 g513(.A(G469), .B(G902), .C1(new_n590), .C2(new_n591), .ZN(new_n700));
  NOR3_X1   g514(.A1(new_n699), .A2(new_n700), .A3(new_n570), .ZN(new_n701));
  NAND4_X1  g515(.A1(new_n657), .A2(new_n628), .A3(new_n698), .A4(new_n701), .ZN(new_n702));
  XNOR2_X1  g516(.A(KEYINPUT41), .B(G113), .ZN(new_n703));
  XNOR2_X1  g517(.A(new_n702), .B(new_n703), .ZN(G15));
  NAND4_X1  g518(.A1(new_n657), .A2(new_n698), .A3(new_n638), .A4(new_n701), .ZN(new_n705));
  XNOR2_X1  g519(.A(new_n705), .B(G116), .ZN(G18));
  NAND2_X1  g520(.A1(new_n660), .A2(new_n701), .ZN(new_n707));
  INV_X1    g521(.A(new_n707), .ZN(new_n708));
  NAND2_X1  g522(.A1(new_n650), .A2(new_n241), .ZN(new_n709));
  NAND2_X1  g523(.A1(new_n240), .A2(new_n709), .ZN(new_n710));
  AND2_X1   g524(.A1(new_n710), .A2(new_n568), .ZN(new_n711));
  NAND3_X1  g525(.A1(new_n708), .A2(new_n711), .A3(new_n657), .ZN(new_n712));
  XNOR2_X1  g526(.A(new_n712), .B(G119), .ZN(G21));
  OAI211_X1 g527(.A(new_n684), .B(new_n376), .C1(new_n626), .C2(new_n453), .ZN(new_n714));
  XNOR2_X1  g528(.A(new_n714), .B(KEYINPUT105), .ZN(new_n715));
  INV_X1    g529(.A(KEYINPUT103), .ZN(new_n716));
  OAI211_X1 g530(.A(new_n340), .B(new_n716), .C1(new_n370), .C2(new_n327), .ZN(new_n717));
  INV_X1    g531(.A(new_n717), .ZN(new_n718));
  NOR2_X1   g532(.A1(new_n718), .A2(new_n341), .ZN(new_n719));
  OAI21_X1  g533(.A(new_n340), .B1(new_n370), .B2(new_n327), .ZN(new_n720));
  NAND2_X1  g534(.A1(new_n720), .A2(KEYINPUT103), .ZN(new_n721));
  AOI21_X1  g535(.A(new_n356), .B1(new_n719), .B2(new_n721), .ZN(new_n722));
  AOI21_X1  g536(.A(G902), .B1(new_n357), .B2(new_n360), .ZN(new_n723));
  OAI21_X1  g537(.A(KEYINPUT104), .B1(new_n723), .B2(new_n679), .ZN(new_n724));
  AOI21_X1  g538(.A(new_n679), .B1(new_n352), .B2(new_n188), .ZN(new_n725));
  INV_X1    g539(.A(KEYINPUT104), .ZN(new_n726));
  NAND2_X1  g540(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  AOI21_X1  g541(.A(new_n722), .B1(new_n724), .B2(new_n727), .ZN(new_n728));
  INV_X1    g542(.A(new_n567), .ZN(new_n729));
  AND2_X1   g543(.A1(new_n701), .A2(new_n729), .ZN(new_n730));
  NAND4_X1  g544(.A1(new_n715), .A2(new_n698), .A3(new_n728), .A4(new_n730), .ZN(new_n731));
  XNOR2_X1  g545(.A(new_n731), .B(G122), .ZN(G24));
  INV_X1    g546(.A(new_n722), .ZN(new_n733));
  NOR2_X1   g547(.A1(new_n725), .A2(new_n726), .ZN(new_n734));
  AOI211_X1 g548(.A(KEYINPUT104), .B(new_n679), .C1(new_n352), .C2(new_n188), .ZN(new_n735));
  OAI211_X1 g549(.A(new_n710), .B(new_n733), .C1(new_n734), .C2(new_n735), .ZN(new_n736));
  INV_X1    g550(.A(new_n736), .ZN(new_n737));
  NAND3_X1  g551(.A1(new_n737), .A2(new_n695), .A3(new_n708), .ZN(new_n738));
  XOR2_X1   g552(.A(KEYINPUT106), .B(G125), .Z(new_n739));
  XNOR2_X1  g553(.A(new_n738), .B(new_n739), .ZN(G27));
  NAND4_X1  g554(.A1(new_n460), .A2(new_n670), .A3(new_n376), .A4(new_n671), .ZN(new_n741));
  NAND2_X1  g555(.A1(new_n693), .A2(new_n694), .ZN(new_n742));
  NOR3_X1   g556(.A1(new_n741), .A2(new_n666), .A3(new_n742), .ZN(new_n743));
  NAND2_X1  g557(.A1(new_n678), .A2(KEYINPUT107), .ZN(new_n744));
  NAND2_X1  g558(.A1(new_n349), .A2(new_n351), .ZN(new_n745));
  NAND2_X1  g559(.A1(new_n373), .A2(G472), .ZN(new_n746));
  INV_X1    g560(.A(KEYINPUT107), .ZN(new_n747));
  NAND4_X1  g561(.A1(new_n352), .A2(new_n747), .A3(KEYINPUT32), .A4(new_n244), .ZN(new_n748));
  NAND4_X1  g562(.A1(new_n744), .A2(new_n745), .A3(new_n746), .A4(new_n748), .ZN(new_n749));
  INV_X1    g563(.A(KEYINPUT108), .ZN(new_n750));
  AND3_X1   g564(.A1(new_n749), .A2(new_n750), .A3(new_n698), .ZN(new_n751));
  AOI21_X1  g565(.A(new_n750), .B1(new_n749), .B2(new_n698), .ZN(new_n752));
  OAI211_X1 g566(.A(KEYINPUT42), .B(new_n743), .C1(new_n751), .C2(new_n752), .ZN(new_n753));
  NOR2_X1   g567(.A1(new_n741), .A2(new_n666), .ZN(new_n754));
  NAND3_X1  g568(.A1(new_n754), .A2(new_n375), .A3(new_n695), .ZN(new_n755));
  INV_X1    g569(.A(KEYINPUT42), .ZN(new_n756));
  NAND2_X1  g570(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  NAND2_X1  g571(.A1(new_n753), .A2(new_n757), .ZN(new_n758));
  XNOR2_X1  g572(.A(new_n758), .B(G131), .ZN(G33));
  NAND3_X1  g573(.A1(new_n754), .A2(new_n375), .A3(new_n665), .ZN(new_n760));
  XNOR2_X1  g574(.A(new_n760), .B(G134), .ZN(G36));
  NOR2_X1   g575(.A1(new_n562), .A2(new_n624), .ZN(new_n762));
  XOR2_X1   g576(.A(new_n762), .B(KEYINPUT43), .Z(new_n763));
  INV_X1    g577(.A(new_n602), .ZN(new_n764));
  NOR3_X1   g578(.A1(new_n763), .A2(new_n764), .A3(new_n651), .ZN(new_n765));
  NAND2_X1  g579(.A1(new_n765), .A2(KEYINPUT44), .ZN(new_n766));
  XOR2_X1   g580(.A(new_n766), .B(KEYINPUT109), .Z(new_n767));
  INV_X1    g581(.A(new_n741), .ZN(new_n768));
  OAI21_X1  g582(.A(new_n768), .B1(new_n765), .B2(KEYINPUT44), .ZN(new_n769));
  OR2_X1    g583(.A1(new_n587), .A2(KEYINPUT45), .ZN(new_n770));
  NAND2_X1  g584(.A1(new_n587), .A2(KEYINPUT45), .ZN(new_n771));
  NAND3_X1  g585(.A1(new_n770), .A2(G469), .A3(new_n771), .ZN(new_n772));
  NAND2_X1  g586(.A1(G469), .A2(G902), .ZN(new_n773));
  AOI21_X1  g587(.A(KEYINPUT46), .B1(new_n772), .B2(new_n773), .ZN(new_n774));
  NOR2_X1   g588(.A1(new_n774), .A2(new_n700), .ZN(new_n775));
  NAND3_X1  g589(.A1(new_n772), .A2(KEYINPUT46), .A3(new_n773), .ZN(new_n776));
  AOI21_X1  g590(.A(new_n570), .B1(new_n775), .B2(new_n776), .ZN(new_n777));
  NAND2_X1  g591(.A1(new_n777), .A2(new_n675), .ZN(new_n778));
  NOR2_X1   g592(.A1(new_n769), .A2(new_n778), .ZN(new_n779));
  NAND2_X1  g593(.A1(new_n767), .A2(new_n779), .ZN(new_n780));
  XNOR2_X1  g594(.A(new_n780), .B(G137), .ZN(G39));
  INV_X1    g595(.A(KEYINPUT110), .ZN(new_n782));
  NAND2_X1  g596(.A1(new_n777), .A2(new_n782), .ZN(new_n783));
  INV_X1    g597(.A(KEYINPUT111), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n784), .A2(KEYINPUT47), .ZN(new_n785));
  NAND2_X1  g599(.A1(new_n783), .A2(new_n785), .ZN(new_n786));
  NOR2_X1   g600(.A1(new_n784), .A2(KEYINPUT47), .ZN(new_n787));
  NOR2_X1   g601(.A1(new_n777), .A2(new_n782), .ZN(new_n788));
  OR3_X1    g602(.A1(new_n786), .A2(new_n787), .A3(new_n788), .ZN(new_n789));
  OAI21_X1  g603(.A(new_n787), .B1(new_n786), .B2(new_n788), .ZN(new_n790));
  NAND2_X1  g604(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  NOR4_X1   g605(.A1(new_n657), .A2(new_n741), .A3(new_n698), .A4(new_n742), .ZN(new_n792));
  NAND2_X1  g606(.A1(new_n791), .A2(new_n792), .ZN(new_n793));
  XNOR2_X1  g607(.A(new_n793), .B(G140), .ZN(G42));
  NOR2_X1   g608(.A1(new_n699), .A2(new_n700), .ZN(new_n795));
  INV_X1    g609(.A(new_n795), .ZN(new_n796));
  OR2_X1    g610(.A1(new_n796), .A2(KEYINPUT49), .ZN(new_n797));
  NAND2_X1  g611(.A1(new_n796), .A2(KEYINPUT49), .ZN(new_n798));
  NOR2_X1   g612(.A1(new_n570), .A2(new_n377), .ZN(new_n799));
  NAND4_X1  g613(.A1(new_n797), .A2(new_n762), .A3(new_n798), .A4(new_n799), .ZN(new_n800));
  OR4_X1    g614(.A1(new_n243), .A2(new_n673), .A3(new_n683), .A4(new_n800), .ZN(new_n801));
  NOR2_X1   g615(.A1(new_n763), .A2(new_n661), .ZN(new_n802));
  NAND3_X1  g616(.A1(new_n802), .A2(new_n698), .A3(new_n728), .ZN(new_n803));
  INV_X1    g617(.A(new_n803), .ZN(new_n804));
  NOR2_X1   g618(.A1(new_n796), .A2(new_n569), .ZN(new_n805));
  OAI211_X1 g619(.A(new_n768), .B(new_n804), .C1(new_n791), .C2(new_n805), .ZN(new_n806));
  INV_X1    g620(.A(new_n701), .ZN(new_n807));
  NOR4_X1   g621(.A1(new_n803), .A2(new_n673), .A3(new_n376), .A4(new_n807), .ZN(new_n808));
  XNOR2_X1  g622(.A(new_n808), .B(KEYINPUT50), .ZN(new_n809));
  NOR2_X1   g623(.A1(new_n741), .A2(new_n807), .ZN(new_n810));
  NAND2_X1  g624(.A1(new_n802), .A2(new_n810), .ZN(new_n811));
  NOR2_X1   g625(.A1(new_n811), .A2(new_n736), .ZN(new_n812));
  XOR2_X1   g626(.A(new_n812), .B(KEYINPUT120), .Z(new_n813));
  INV_X1    g627(.A(new_n810), .ZN(new_n814));
  NOR4_X1   g628(.A1(new_n814), .A2(new_n243), .A3(new_n683), .A4(new_n661), .ZN(new_n815));
  NOR2_X1   g629(.A1(new_n562), .A2(new_n690), .ZN(new_n816));
  AOI21_X1  g630(.A(new_n813), .B1(new_n815), .B2(new_n816), .ZN(new_n817));
  NAND3_X1  g631(.A1(new_n806), .A2(new_n809), .A3(new_n817), .ZN(new_n818));
  INV_X1    g632(.A(KEYINPUT51), .ZN(new_n819));
  NOR2_X1   g633(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  NAND2_X1  g634(.A1(new_n818), .A2(new_n819), .ZN(new_n821));
  NOR2_X1   g635(.A1(new_n751), .A2(new_n752), .ZN(new_n822));
  NOR2_X1   g636(.A1(new_n822), .A2(new_n811), .ZN(new_n823));
  XOR2_X1   g637(.A(new_n823), .B(KEYINPUT48), .Z(new_n824));
  NAND2_X1  g638(.A1(new_n804), .A2(new_n708), .ZN(new_n825));
  XNOR2_X1  g639(.A(new_n825), .B(KEYINPUT121), .ZN(new_n826));
  NOR2_X1   g640(.A1(new_n614), .A2(new_n624), .ZN(new_n827));
  AOI211_X1 g641(.A(new_n563), .B(G953), .C1(new_n815), .C2(new_n827), .ZN(new_n828));
  NAND4_X1  g642(.A1(new_n821), .A2(new_n824), .A3(new_n826), .A4(new_n828), .ZN(new_n829));
  NAND2_X1  g643(.A1(new_n651), .A2(new_n663), .ZN(new_n830));
  XNOR2_X1  g644(.A(new_n830), .B(KEYINPUT116), .ZN(new_n831));
  NAND4_X1  g645(.A1(new_n831), .A2(new_n595), .A3(new_n683), .A4(new_n715), .ZN(new_n832));
  NAND4_X1  g646(.A1(new_n832), .A2(new_n668), .A3(new_n696), .A4(new_n738), .ZN(new_n833));
  NAND2_X1  g647(.A1(new_n833), .A2(KEYINPUT52), .ZN(new_n834));
  NAND2_X1  g648(.A1(new_n738), .A2(new_n668), .ZN(new_n835));
  INV_X1    g649(.A(new_n835), .ZN(new_n836));
  INV_X1    g650(.A(KEYINPUT52), .ZN(new_n837));
  NAND4_X1  g651(.A1(new_n836), .A2(new_n837), .A3(new_n696), .A4(new_n832), .ZN(new_n838));
  NAND2_X1  g652(.A1(new_n834), .A2(new_n838), .ZN(new_n839));
  NAND2_X1  g653(.A1(new_n510), .A2(KEYINPUT112), .ZN(new_n840));
  INV_X1    g654(.A(KEYINPUT112), .ZN(new_n841));
  NAND2_X1  g655(.A1(new_n632), .A2(new_n841), .ZN(new_n842));
  AND4_X1   g656(.A1(new_n614), .A2(new_n840), .A3(new_n729), .A4(new_n842), .ZN(new_n843));
  NAND3_X1  g657(.A1(new_n672), .A2(new_n376), .A3(new_n843), .ZN(new_n844));
  INV_X1    g658(.A(KEYINPUT113), .ZN(new_n845));
  NAND2_X1  g659(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  NAND4_X1  g660(.A1(new_n672), .A2(new_n843), .A3(KEYINPUT113), .A4(new_n376), .ZN(new_n847));
  NAND3_X1  g661(.A1(new_n846), .A2(new_n604), .A3(new_n847), .ZN(new_n848));
  NAND3_X1  g662(.A1(new_n461), .A2(new_n604), .A3(new_n625), .ZN(new_n849));
  NAND4_X1  g663(.A1(new_n848), .A2(new_n597), .A3(new_n653), .A4(new_n849), .ZN(new_n850));
  NAND4_X1  g664(.A1(new_n455), .A2(new_n376), .A3(new_n460), .A4(new_n595), .ZN(new_n851));
  INV_X1    g665(.A(KEYINPUT114), .ZN(new_n852));
  NOR4_X1   g666(.A1(new_n851), .A2(new_n736), .A3(new_n852), .A4(new_n742), .ZN(new_n853));
  AOI21_X1  g667(.A(KEYINPUT114), .B1(new_n743), .B2(new_n737), .ZN(new_n854));
  NOR2_X1   g668(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  NOR2_X1   g669(.A1(new_n850), .A2(new_n855), .ZN(new_n856));
  NAND4_X1  g670(.A1(new_n731), .A2(new_n702), .A3(new_n705), .A4(new_n712), .ZN(new_n857));
  AND2_X1   g671(.A1(new_n840), .A2(new_n842), .ZN(new_n858));
  NOR2_X1   g672(.A1(new_n858), .A2(new_n664), .ZN(new_n859));
  NAND4_X1  g673(.A1(new_n768), .A2(new_n657), .A3(new_n667), .A4(new_n859), .ZN(new_n860));
  NAND2_X1  g674(.A1(new_n760), .A2(new_n860), .ZN(new_n861));
  NOR2_X1   g675(.A1(new_n857), .A2(new_n861), .ZN(new_n862));
  NAND4_X1  g676(.A1(new_n856), .A2(KEYINPUT115), .A3(new_n758), .A4(new_n862), .ZN(new_n863));
  INV_X1    g677(.A(KEYINPUT115), .ZN(new_n864));
  INV_X1    g678(.A(KEYINPUT105), .ZN(new_n865));
  XNOR2_X1  g679(.A(new_n714), .B(new_n865), .ZN(new_n866));
  NAND2_X1  g680(.A1(new_n724), .A2(new_n727), .ZN(new_n867));
  NAND4_X1  g681(.A1(new_n867), .A2(new_n698), .A3(new_n730), .A4(new_n733), .ZN(new_n868));
  OAI21_X1  g682(.A(new_n705), .B1(new_n866), .B2(new_n868), .ZN(new_n869));
  NAND2_X1  g683(.A1(new_n702), .A2(new_n712), .ZN(new_n870));
  NOR2_X1   g684(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  INV_X1    g685(.A(new_n861), .ZN(new_n872));
  NAND3_X1  g686(.A1(new_n758), .A2(new_n871), .A3(new_n872), .ZN(new_n873));
  AND3_X1   g687(.A1(new_n460), .A2(new_n670), .A3(new_n671), .ZN(new_n874));
  NAND4_X1  g688(.A1(new_n874), .A2(new_n376), .A3(new_n595), .A4(new_n695), .ZN(new_n875));
  OAI21_X1  g689(.A(new_n852), .B1(new_n875), .B2(new_n736), .ZN(new_n876));
  NAND3_X1  g690(.A1(new_n743), .A2(KEYINPUT114), .A3(new_n737), .ZN(new_n877));
  NAND2_X1  g691(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  AND3_X1   g692(.A1(new_n597), .A2(new_n849), .A3(new_n653), .ZN(new_n879));
  NAND3_X1  g693(.A1(new_n878), .A2(new_n879), .A3(new_n848), .ZN(new_n880));
  OAI21_X1  g694(.A(new_n864), .B1(new_n873), .B2(new_n880), .ZN(new_n881));
  AOI21_X1  g695(.A(new_n839), .B1(new_n863), .B2(new_n881), .ZN(new_n882));
  INV_X1    g696(.A(KEYINPUT53), .ZN(new_n883));
  OAI21_X1  g697(.A(new_n883), .B1(new_n836), .B2(new_n837), .ZN(new_n884));
  AND2_X1   g698(.A1(new_n882), .A2(new_n884), .ZN(new_n885));
  NAND2_X1  g699(.A1(new_n863), .A2(new_n881), .ZN(new_n886));
  INV_X1    g700(.A(new_n839), .ZN(new_n887));
  AOI21_X1  g701(.A(KEYINPUT53), .B1(new_n886), .B2(new_n887), .ZN(new_n888));
  OAI21_X1  g702(.A(KEYINPUT54), .B1(new_n885), .B2(new_n888), .ZN(new_n889));
  AND3_X1   g703(.A1(new_n758), .A2(new_n871), .A3(new_n872), .ZN(new_n890));
  AOI21_X1  g704(.A(KEYINPUT115), .B1(new_n890), .B2(new_n856), .ZN(new_n891));
  NOR3_X1   g705(.A1(new_n873), .A2(new_n880), .A3(new_n864), .ZN(new_n892));
  OAI21_X1  g706(.A(new_n887), .B1(new_n891), .B2(new_n892), .ZN(new_n893));
  NAND3_X1  g707(.A1(new_n893), .A2(KEYINPUT117), .A3(new_n883), .ZN(new_n894));
  INV_X1    g708(.A(KEYINPUT117), .ZN(new_n895));
  OAI21_X1  g709(.A(new_n895), .B1(new_n882), .B2(KEYINPUT53), .ZN(new_n896));
  INV_X1    g710(.A(KEYINPUT118), .ZN(new_n897));
  NOR2_X1   g711(.A1(new_n873), .A2(new_n880), .ZN(new_n898));
  INV_X1    g712(.A(new_n898), .ZN(new_n899));
  AOI21_X1  g713(.A(new_n883), .B1(new_n835), .B2(KEYINPUT52), .ZN(new_n900));
  NAND3_X1  g714(.A1(new_n834), .A2(new_n838), .A3(new_n900), .ZN(new_n901));
  OAI21_X1  g715(.A(new_n897), .B1(new_n899), .B2(new_n901), .ZN(new_n902));
  NAND4_X1  g716(.A1(new_n887), .A2(new_n898), .A3(KEYINPUT118), .A4(new_n900), .ZN(new_n903));
  NAND2_X1  g717(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  NAND3_X1  g718(.A1(new_n894), .A2(new_n896), .A3(new_n904), .ZN(new_n905));
  OAI211_X1 g719(.A(new_n889), .B(KEYINPUT119), .C1(new_n905), .C2(KEYINPUT54), .ZN(new_n906));
  AOI22_X1  g720(.A1(new_n888), .A2(KEYINPUT117), .B1(new_n902), .B2(new_n903), .ZN(new_n907));
  INV_X1    g721(.A(KEYINPUT119), .ZN(new_n908));
  INV_X1    g722(.A(KEYINPUT54), .ZN(new_n909));
  NAND4_X1  g723(.A1(new_n907), .A2(new_n908), .A3(new_n909), .A4(new_n896), .ZN(new_n910));
  AOI211_X1 g724(.A(new_n820), .B(new_n829), .C1(new_n906), .C2(new_n910), .ZN(new_n911));
  NOR2_X1   g725(.A1(G952), .A2(G953), .ZN(new_n912));
  OAI21_X1  g726(.A(new_n801), .B1(new_n911), .B2(new_n912), .ZN(G75));
  NOR2_X1   g727(.A1(new_n222), .A2(G952), .ZN(new_n914));
  INV_X1    g728(.A(new_n914), .ZN(new_n915));
  AOI21_X1  g729(.A(new_n188), .B1(new_n907), .B2(new_n896), .ZN(new_n916));
  AOI21_X1  g730(.A(KEYINPUT56), .B1(new_n916), .B2(new_n379), .ZN(new_n917));
  NAND2_X1  g731(.A1(new_n417), .A2(new_n426), .ZN(new_n918));
  XOR2_X1   g732(.A(new_n918), .B(new_n424), .Z(new_n919));
  XNOR2_X1  g733(.A(new_n919), .B(KEYINPUT55), .ZN(new_n920));
  INV_X1    g734(.A(new_n920), .ZN(new_n921));
  OAI21_X1  g735(.A(new_n915), .B1(new_n917), .B2(new_n921), .ZN(new_n922));
  AOI21_X1  g736(.A(new_n922), .B1(new_n917), .B2(new_n921), .ZN(G51));
  XNOR2_X1  g737(.A(new_n905), .B(new_n909), .ZN(new_n924));
  XNOR2_X1  g738(.A(new_n773), .B(KEYINPUT57), .ZN(new_n925));
  OAI21_X1  g739(.A(new_n592), .B1(new_n924), .B2(new_n925), .ZN(new_n926));
  NAND4_X1  g740(.A1(new_n916), .A2(G469), .A3(new_n771), .A4(new_n770), .ZN(new_n927));
  AOI21_X1  g741(.A(new_n914), .B1(new_n926), .B2(new_n927), .ZN(G54));
  NAND3_X1  g742(.A1(new_n916), .A2(KEYINPUT58), .A3(G475), .ZN(new_n929));
  AND2_X1   g743(.A1(new_n929), .A2(new_n611), .ZN(new_n930));
  NOR2_X1   g744(.A1(new_n929), .A2(new_n611), .ZN(new_n931));
  NOR3_X1   g745(.A1(new_n930), .A2(new_n931), .A3(new_n914), .ZN(G60));
  INV_X1    g746(.A(new_n617), .ZN(new_n933));
  NAND2_X1  g747(.A1(new_n906), .A2(new_n910), .ZN(new_n934));
  NAND2_X1  g748(.A1(G478), .A2(G902), .ZN(new_n935));
  XOR2_X1   g749(.A(new_n935), .B(KEYINPUT59), .Z(new_n936));
  OAI21_X1  g750(.A(new_n933), .B1(new_n934), .B2(new_n936), .ZN(new_n937));
  XNOR2_X1  g751(.A(new_n905), .B(KEYINPUT54), .ZN(new_n938));
  NOR2_X1   g752(.A1(new_n933), .A2(new_n936), .ZN(new_n939));
  AOI21_X1  g753(.A(new_n914), .B1(new_n938), .B2(new_n939), .ZN(new_n940));
  AND2_X1   g754(.A1(new_n937), .A2(new_n940), .ZN(G63));
  NAND2_X1  g755(.A1(G217), .A2(G902), .ZN(new_n942));
  XNOR2_X1  g756(.A(new_n942), .B(KEYINPUT60), .ZN(new_n943));
  INV_X1    g757(.A(new_n943), .ZN(new_n944));
  NAND3_X1  g758(.A1(new_n905), .A2(new_n650), .A3(new_n944), .ZN(new_n945));
  AOI21_X1  g759(.A(new_n943), .B1(new_n907), .B2(new_n896), .ZN(new_n946));
  OAI211_X1 g760(.A(new_n945), .B(new_n915), .C1(new_n946), .C2(new_n232), .ZN(new_n947));
  AND3_X1   g761(.A1(new_n947), .A2(KEYINPUT122), .A3(KEYINPUT61), .ZN(new_n948));
  AOI21_X1  g762(.A(KEYINPUT61), .B1(new_n947), .B2(KEYINPUT122), .ZN(new_n949));
  NOR2_X1   g763(.A1(new_n948), .A2(new_n949), .ZN(G66));
  OAI21_X1  g764(.A(G953), .B1(new_n566), .B2(new_n422), .ZN(new_n951));
  NOR2_X1   g765(.A1(new_n850), .A2(new_n857), .ZN(new_n952));
  OAI21_X1  g766(.A(new_n951), .B1(new_n952), .B2(G953), .ZN(new_n953));
  OAI21_X1  g767(.A(new_n918), .B1(G898), .B2(new_n222), .ZN(new_n954));
  XNOR2_X1  g768(.A(new_n953), .B(new_n954), .ZN(G69));
  AOI21_X1  g769(.A(new_n827), .B1(new_n858), .B2(new_n614), .ZN(new_n956));
  NOR2_X1   g770(.A1(new_n956), .A2(new_n676), .ZN(new_n957));
  NAND3_X1  g771(.A1(new_n957), .A2(new_n375), .A3(new_n768), .ZN(new_n958));
  NAND2_X1  g772(.A1(new_n780), .A2(new_n958), .ZN(new_n959));
  INV_X1    g773(.A(KEYINPUT124), .ZN(new_n960));
  NAND2_X1  g774(.A1(new_n959), .A2(new_n960), .ZN(new_n961));
  NAND3_X1  g775(.A1(new_n780), .A2(KEYINPUT124), .A3(new_n958), .ZN(new_n962));
  AOI22_X1  g776(.A1(new_n961), .A2(new_n962), .B1(new_n791), .B2(new_n792), .ZN(new_n963));
  NAND2_X1  g777(.A1(new_n836), .A2(new_n696), .ZN(new_n964));
  XNOR2_X1  g778(.A(new_n964), .B(KEYINPUT123), .ZN(new_n965));
  NAND2_X1  g779(.A1(new_n965), .A2(new_n686), .ZN(new_n966));
  OR2_X1    g780(.A1(new_n966), .A2(KEYINPUT62), .ZN(new_n967));
  NAND2_X1  g781(.A1(new_n966), .A2(KEYINPUT62), .ZN(new_n968));
  NAND3_X1  g782(.A1(new_n963), .A2(new_n967), .A3(new_n968), .ZN(new_n969));
  INV_X1    g783(.A(new_n336), .ZN(new_n970));
  INV_X1    g784(.A(new_n338), .ZN(new_n971));
  NOR2_X1   g785(.A1(new_n970), .A2(new_n971), .ZN(new_n972));
  NAND3_X1  g786(.A1(new_n548), .A2(new_n550), .A3(new_n551), .ZN(new_n973));
  XOR2_X1   g787(.A(new_n972), .B(new_n973), .Z(new_n974));
  AND2_X1   g788(.A1(new_n974), .A2(new_n222), .ZN(new_n975));
  AOI21_X1  g789(.A(new_n222), .B1(G227), .B2(G900), .ZN(new_n976));
  INV_X1    g790(.A(new_n976), .ZN(new_n977));
  AOI22_X1  g791(.A1(new_n969), .A2(new_n975), .B1(KEYINPUT126), .B2(new_n977), .ZN(new_n978));
  INV_X1    g792(.A(new_n978), .ZN(new_n979));
  INV_X1    g793(.A(KEYINPUT125), .ZN(new_n980));
  INV_X1    g794(.A(new_n760), .ZN(new_n981));
  AOI21_X1  g795(.A(new_n981), .B1(new_n767), .B2(new_n779), .ZN(new_n982));
  OR3_X1    g796(.A1(new_n778), .A2(new_n822), .A3(new_n866), .ZN(new_n983));
  NAND4_X1  g797(.A1(new_n793), .A2(new_n758), .A3(new_n982), .A4(new_n983), .ZN(new_n984));
  INV_X1    g798(.A(new_n965), .ZN(new_n985));
  OAI21_X1  g799(.A(new_n980), .B1(new_n984), .B2(new_n985), .ZN(new_n986));
  AND3_X1   g800(.A1(new_n982), .A2(new_n758), .A3(new_n983), .ZN(new_n987));
  NAND4_X1  g801(.A1(new_n987), .A2(KEYINPUT125), .A3(new_n793), .A4(new_n965), .ZN(new_n988));
  NAND3_X1  g802(.A1(new_n986), .A2(new_n988), .A3(new_n222), .ZN(new_n989));
  NAND2_X1  g803(.A1(G900), .A2(G953), .ZN(new_n990));
  AOI21_X1  g804(.A(new_n974), .B1(new_n989), .B2(new_n990), .ZN(new_n991));
  NOR2_X1   g805(.A1(new_n977), .A2(KEYINPUT126), .ZN(new_n992));
  NOR3_X1   g806(.A1(new_n979), .A2(new_n991), .A3(new_n992), .ZN(new_n993));
  INV_X1    g807(.A(new_n992), .ZN(new_n994));
  INV_X1    g808(.A(new_n991), .ZN(new_n995));
  AOI21_X1  g809(.A(new_n994), .B1(new_n995), .B2(new_n978), .ZN(new_n996));
  NOR2_X1   g810(.A1(new_n993), .A2(new_n996), .ZN(G72));
  NAND3_X1  g811(.A1(new_n986), .A2(new_n988), .A3(new_n952), .ZN(new_n998));
  NAND2_X1  g812(.A1(G472), .A2(G902), .ZN(new_n999));
  XOR2_X1   g813(.A(new_n999), .B(KEYINPUT63), .Z(new_n1000));
  AOI21_X1  g814(.A(new_n327), .B1(new_n998), .B2(new_n1000), .ZN(new_n1001));
  NOR2_X1   g815(.A1(new_n339), .A2(new_n362), .ZN(new_n1002));
  NAND4_X1  g816(.A1(new_n963), .A2(new_n968), .A3(new_n952), .A4(new_n967), .ZN(new_n1003));
  AOI21_X1  g817(.A(new_n1002), .B1(new_n1003), .B2(new_n1000), .ZN(new_n1004));
  OAI21_X1  g818(.A(new_n363), .B1(new_n1001), .B2(new_n1004), .ZN(new_n1005));
  NAND2_X1  g819(.A1(new_n365), .A2(new_n346), .ZN(new_n1006));
  OAI211_X1 g820(.A(new_n1000), .B(new_n1006), .C1(new_n885), .C2(new_n888), .ZN(new_n1007));
  AND3_X1   g821(.A1(new_n1005), .A2(new_n915), .A3(new_n1007), .ZN(G57));
endmodule


