//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 0 0 0 0 0 1 0 1 1 0 0 1 0 0 0 1 0 1 1 0 0 1 1 0 0 0 0 0 1 0 1 0 0 1 0 0 1 1 0 1 1 1 0 0 0 1 0 0 0 0 1 1 0 1 0 0 1 1 0 1 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:35:30 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n206, new_n207, new_n208,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n236, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n244, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n252, new_n253,
    new_n254, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n811, new_n812, new_n813,
    new_n814, new_n815, new_n816, new_n817, new_n818, new_n819, new_n820,
    new_n821, new_n822, new_n823, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n981, new_n982, new_n983,
    new_n984, new_n985, new_n986, new_n987, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1017, new_n1018, new_n1019, new_n1020, new_n1021, new_n1022,
    new_n1023, new_n1024, new_n1025, new_n1026, new_n1027, new_n1028,
    new_n1029, new_n1030, new_n1031, new_n1032, new_n1033, new_n1034,
    new_n1035, new_n1036, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1050, new_n1051, new_n1052, new_n1053,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1110, new_n1111, new_n1112, new_n1113, new_n1114,
    new_n1115, new_n1116, new_n1117, new_n1118, new_n1119, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1171, new_n1172, new_n1173, new_n1174, new_n1175,
    new_n1176, new_n1177, new_n1178, new_n1179, new_n1180, new_n1181,
    new_n1182, new_n1183, new_n1184, new_n1185, new_n1186, new_n1187,
    new_n1188, new_n1189, new_n1190, new_n1192, new_n1193, new_n1195,
    new_n1196, new_n1197, new_n1198, new_n1199, new_n1201, new_n1202,
    new_n1203, new_n1204, new_n1205, new_n1206, new_n1207, new_n1208,
    new_n1209, new_n1210, new_n1211, new_n1212, new_n1213, new_n1214,
    new_n1215, new_n1216, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1252, new_n1253, new_n1254, new_n1255, new_n1256, new_n1257,
    new_n1258, new_n1259, new_n1260, new_n1261, new_n1262, new_n1263,
    new_n1264;
  INV_X1    g0000(.A(G50), .ZN(new_n201));
  INV_X1    g0001(.A(G58), .ZN(new_n202));
  INV_X1    g0002(.A(G68), .ZN(new_n203));
  NAND3_X1  g0003(.A1(new_n201), .A2(new_n202), .A3(new_n203), .ZN(new_n204));
  NOR2_X1   g0004(.A1(new_n204), .A2(G77), .ZN(G353));
  INV_X1    g0005(.A(G97), .ZN(new_n206));
  INV_X1    g0006(.A(G107), .ZN(new_n207));
  NAND2_X1  g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  NAND2_X1  g0008(.A1(new_n208), .A2(G87), .ZN(G355));
  NAND2_X1  g0009(.A1(G1), .A2(G20), .ZN(new_n210));
  NOR2_X1   g0010(.A1(new_n210), .A2(G13), .ZN(new_n211));
  OAI211_X1 g0011(.A(new_n211), .B(G250), .C1(G257), .C2(G264), .ZN(new_n212));
  XNOR2_X1  g0012(.A(new_n212), .B(KEYINPUT0), .ZN(new_n213));
  NAND2_X1  g0013(.A1(G1), .A2(G13), .ZN(new_n214));
  NAND2_X1  g0014(.A1(new_n214), .A2(KEYINPUT64), .ZN(new_n215));
  INV_X1    g0015(.A(KEYINPUT64), .ZN(new_n216));
  NAND3_X1  g0016(.A1(new_n216), .A2(G1), .A3(G13), .ZN(new_n217));
  NAND2_X1  g0017(.A1(new_n215), .A2(new_n217), .ZN(new_n218));
  INV_X1    g0018(.A(new_n218), .ZN(new_n219));
  INV_X1    g0019(.A(G20), .ZN(new_n220));
  NOR2_X1   g0020(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  NAND2_X1  g0021(.A1(new_n202), .A2(new_n203), .ZN(new_n222));
  NAND2_X1  g0022(.A1(new_n222), .A2(G50), .ZN(new_n223));
  INV_X1    g0023(.A(new_n223), .ZN(new_n224));
  NAND2_X1  g0024(.A1(new_n221), .A2(new_n224), .ZN(new_n225));
  AOI22_X1  g0025(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n226));
  INV_X1    g0026(.A(G238), .ZN(new_n227));
  INV_X1    g0027(.A(G87), .ZN(new_n228));
  INV_X1    g0028(.A(G250), .ZN(new_n229));
  OAI221_X1 g0029(.A(new_n226), .B1(new_n203), .B2(new_n227), .C1(new_n228), .C2(new_n229), .ZN(new_n230));
  AOI22_X1  g0030(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n231));
  INV_X1    g0031(.A(G232), .ZN(new_n232));
  INV_X1    g0032(.A(G257), .ZN(new_n233));
  OAI221_X1 g0033(.A(new_n231), .B1(new_n202), .B2(new_n232), .C1(new_n206), .C2(new_n233), .ZN(new_n234));
  OAI21_X1  g0034(.A(new_n210), .B1(new_n230), .B2(new_n234), .ZN(new_n235));
  OAI211_X1 g0035(.A(new_n213), .B(new_n225), .C1(KEYINPUT1), .C2(new_n235), .ZN(new_n236));
  AOI21_X1  g0036(.A(new_n236), .B1(KEYINPUT1), .B2(new_n235), .ZN(G361));
  XNOR2_X1  g0037(.A(G238), .B(G244), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n238), .B(G232), .ZN(new_n239));
  XNOR2_X1  g0039(.A(KEYINPUT2), .B(G226), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XOR2_X1   g0041(.A(G264), .B(G270), .Z(new_n242));
  XNOR2_X1  g0042(.A(G250), .B(G257), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n241), .B(new_n244), .ZN(G358));
  XNOR2_X1  g0045(.A(G107), .B(G116), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n246), .B(KEYINPUT65), .ZN(new_n247));
  XOR2_X1   g0047(.A(G87), .B(G97), .Z(new_n248));
  XOR2_X1   g0048(.A(new_n247), .B(new_n248), .Z(new_n249));
  NAND2_X1  g0049(.A1(new_n201), .A2(G68), .ZN(new_n250));
  NAND2_X1  g0050(.A1(new_n203), .A2(G50), .ZN(new_n251));
  NAND2_X1  g0051(.A1(new_n250), .A2(new_n251), .ZN(new_n252));
  XNOR2_X1  g0052(.A(G58), .B(G77), .ZN(new_n253));
  XNOR2_X1  g0053(.A(new_n252), .B(new_n253), .ZN(new_n254));
  XOR2_X1   g0054(.A(new_n249), .B(new_n254), .Z(G351));
  INV_X1    g0055(.A(G33), .ZN(new_n256));
  OAI211_X1 g0056(.A(new_n215), .B(new_n217), .C1(new_n256), .C2(new_n210), .ZN(new_n257));
  OR2_X1    g0057(.A1(new_n257), .A2(KEYINPUT67), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n257), .A2(KEYINPUT67), .ZN(new_n259));
  AND2_X1   g0059(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  NOR2_X1   g0060(.A1(G20), .A2(G33), .ZN(new_n261));
  AOI22_X1  g0061(.A1(new_n204), .A2(G20), .B1(G150), .B2(new_n261), .ZN(new_n262));
  INV_X1    g0062(.A(KEYINPUT8), .ZN(new_n263));
  OR3_X1    g0063(.A1(new_n263), .A2(new_n202), .A3(KEYINPUT68), .ZN(new_n264));
  OAI21_X1  g0064(.A(new_n263), .B1(new_n202), .B2(KEYINPUT68), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n220), .A2(G33), .ZN(new_n267));
  OAI21_X1  g0067(.A(new_n262), .B1(new_n266), .B2(new_n267), .ZN(new_n268));
  INV_X1    g0068(.A(G13), .ZN(new_n269));
  NOR3_X1   g0069(.A1(new_n269), .A2(new_n220), .A3(G1), .ZN(new_n270));
  AOI22_X1  g0070(.A1(new_n260), .A2(new_n268), .B1(new_n201), .B2(new_n270), .ZN(new_n271));
  AOI21_X1  g0071(.A(new_n270), .B1(new_n258), .B2(new_n259), .ZN(new_n272));
  INV_X1    g0072(.A(new_n272), .ZN(new_n273));
  OAI21_X1  g0073(.A(G50), .B1(new_n220), .B2(G1), .ZN(new_n274));
  OAI21_X1  g0074(.A(new_n271), .B1(new_n273), .B2(new_n274), .ZN(new_n275));
  XNOR2_X1  g0075(.A(new_n275), .B(KEYINPUT9), .ZN(new_n276));
  AND2_X1   g0076(.A1(KEYINPUT3), .A2(G33), .ZN(new_n277));
  NOR2_X1   g0077(.A1(KEYINPUT3), .A2(G33), .ZN(new_n278));
  NOR2_X1   g0078(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  NOR2_X1   g0079(.A1(new_n279), .A2(G1698), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n280), .A2(G222), .ZN(new_n281));
  INV_X1    g0081(.A(G1698), .ZN(new_n282));
  OR2_X1    g0082(.A1(KEYINPUT3), .A2(G33), .ZN(new_n283));
  NAND2_X1  g0083(.A1(KEYINPUT3), .A2(G33), .ZN(new_n284));
  AOI21_X1  g0084(.A(new_n282), .B1(new_n283), .B2(new_n284), .ZN(new_n285));
  AOI22_X1  g0085(.A1(new_n285), .A2(G223), .B1(new_n279), .B2(G77), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n281), .A2(new_n286), .ZN(new_n287));
  NAND2_X1  g0087(.A1(G33), .A2(G41), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n218), .A2(new_n288), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n289), .A2(KEYINPUT66), .ZN(new_n290));
  INV_X1    g0090(.A(KEYINPUT66), .ZN(new_n291));
  NAND3_X1  g0091(.A1(new_n218), .A2(new_n291), .A3(new_n288), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n290), .A2(new_n292), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n287), .A2(new_n293), .ZN(new_n294));
  INV_X1    g0094(.A(G1), .ZN(new_n295));
  OAI21_X1  g0095(.A(new_n295), .B1(G41), .B2(G45), .ZN(new_n296));
  INV_X1    g0096(.A(new_n296), .ZN(new_n297));
  NAND3_X1  g0097(.A1(new_n288), .A2(G1), .A3(G13), .ZN(new_n298));
  NAND3_X1  g0098(.A1(new_n297), .A2(new_n298), .A3(G274), .ZN(new_n299));
  INV_X1    g0099(.A(G226), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n298), .A2(new_n296), .ZN(new_n301));
  OAI211_X1 g0101(.A(new_n294), .B(new_n299), .C1(new_n300), .C2(new_n301), .ZN(new_n302));
  INV_X1    g0102(.A(G190), .ZN(new_n303));
  NOR2_X1   g0103(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  AOI21_X1  g0104(.A(new_n304), .B1(G200), .B2(new_n302), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n276), .A2(new_n305), .ZN(new_n306));
  XNOR2_X1  g0106(.A(new_n306), .B(KEYINPUT10), .ZN(new_n307));
  INV_X1    g0107(.A(G169), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n302), .A2(new_n308), .ZN(new_n309));
  OAI211_X1 g0109(.A(new_n275), .B(new_n309), .C1(G179), .C2(new_n302), .ZN(new_n310));
  INV_X1    g0110(.A(G77), .ZN(new_n311));
  NOR2_X1   g0111(.A1(new_n220), .A2(G1), .ZN(new_n312));
  NOR3_X1   g0112(.A1(new_n273), .A2(new_n311), .A3(new_n312), .ZN(new_n313));
  NAND2_X1  g0113(.A1(G20), .A2(G77), .ZN(new_n314));
  XNOR2_X1  g0114(.A(KEYINPUT15), .B(G87), .ZN(new_n315));
  INV_X1    g0115(.A(new_n261), .ZN(new_n316));
  XNOR2_X1  g0116(.A(KEYINPUT8), .B(G58), .ZN(new_n317));
  OAI221_X1 g0117(.A(new_n314), .B1(new_n315), .B2(new_n267), .C1(new_n316), .C2(new_n317), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n260), .A2(new_n318), .ZN(new_n319));
  INV_X1    g0119(.A(new_n270), .ZN(new_n320));
  OAI21_X1  g0120(.A(new_n319), .B1(G77), .B2(new_n320), .ZN(new_n321));
  NOR2_X1   g0121(.A1(new_n313), .A2(new_n321), .ZN(new_n322));
  XNOR2_X1  g0122(.A(KEYINPUT69), .B(G107), .ZN(new_n323));
  INV_X1    g0123(.A(new_n323), .ZN(new_n324));
  AOI22_X1  g0124(.A1(new_n279), .A2(new_n324), .B1(new_n285), .B2(G238), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n280), .A2(G232), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n327), .A2(new_n293), .ZN(new_n328));
  INV_X1    g0128(.A(new_n301), .ZN(new_n329));
  AND2_X1   g0129(.A1(new_n298), .A2(G274), .ZN(new_n330));
  AOI22_X1  g0130(.A1(G244), .A2(new_n329), .B1(new_n330), .B2(new_n297), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n328), .A2(new_n331), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n332), .A2(G200), .ZN(new_n333));
  OAI211_X1 g0133(.A(new_n322), .B(new_n333), .C1(new_n303), .C2(new_n332), .ZN(new_n334));
  INV_X1    g0134(.A(new_n322), .ZN(new_n335));
  INV_X1    g0135(.A(G179), .ZN(new_n336));
  NAND3_X1  g0136(.A1(new_n328), .A2(new_n336), .A3(new_n331), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n332), .A2(new_n308), .ZN(new_n338));
  NAND3_X1  g0138(.A1(new_n335), .A2(new_n337), .A3(new_n338), .ZN(new_n339));
  NAND4_X1  g0139(.A1(new_n307), .A2(new_n310), .A3(new_n334), .A4(new_n339), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n283), .A2(new_n284), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n232), .A2(G1698), .ZN(new_n342));
  OAI211_X1 g0142(.A(new_n341), .B(new_n342), .C1(G226), .C2(G1698), .ZN(new_n343));
  NAND2_X1  g0143(.A1(G33), .A2(G97), .ZN(new_n344));
  AOI22_X1  g0144(.A1(new_n290), .A2(new_n292), .B1(new_n343), .B2(new_n344), .ZN(new_n345));
  OAI21_X1  g0145(.A(new_n299), .B1(new_n227), .B2(new_n301), .ZN(new_n346));
  OAI21_X1  g0146(.A(KEYINPUT13), .B1(new_n345), .B2(new_n346), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n343), .A2(new_n344), .ZN(new_n348));
  AND2_X1   g0148(.A1(G33), .A2(G41), .ZN(new_n349));
  AOI211_X1 g0149(.A(KEYINPUT66), .B(new_n349), .C1(new_n215), .C2(new_n217), .ZN(new_n350));
  AOI21_X1  g0150(.A(new_n291), .B1(new_n218), .B2(new_n288), .ZN(new_n351));
  OAI21_X1  g0151(.A(new_n348), .B1(new_n350), .B2(new_n351), .ZN(new_n352));
  INV_X1    g0152(.A(KEYINPUT13), .ZN(new_n353));
  INV_X1    g0153(.A(new_n346), .ZN(new_n354));
  NAND3_X1  g0154(.A1(new_n352), .A2(new_n353), .A3(new_n354), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n347), .A2(new_n355), .ZN(new_n356));
  INV_X1    g0156(.A(KEYINPUT14), .ZN(new_n357));
  NAND3_X1  g0157(.A1(new_n356), .A2(new_n357), .A3(G169), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n358), .A2(KEYINPUT70), .ZN(new_n359));
  AND2_X1   g0159(.A1(new_n347), .A2(new_n355), .ZN(new_n360));
  OAI21_X1  g0160(.A(KEYINPUT14), .B1(new_n360), .B2(new_n308), .ZN(new_n361));
  INV_X1    g0161(.A(KEYINPUT70), .ZN(new_n362));
  NAND4_X1  g0162(.A1(new_n356), .A2(new_n362), .A3(new_n357), .A4(G169), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n360), .A2(G179), .ZN(new_n364));
  NAND4_X1  g0164(.A1(new_n359), .A2(new_n361), .A3(new_n363), .A4(new_n364), .ZN(new_n365));
  AOI22_X1  g0165(.A1(new_n261), .A2(G50), .B1(G20), .B2(new_n203), .ZN(new_n366));
  OAI21_X1  g0166(.A(new_n366), .B1(new_n311), .B2(new_n267), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n260), .A2(new_n367), .ZN(new_n368));
  INV_X1    g0168(.A(KEYINPUT11), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n368), .A2(new_n369), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n270), .A2(new_n203), .ZN(new_n371));
  XNOR2_X1  g0171(.A(new_n371), .B(KEYINPUT12), .ZN(new_n372));
  NAND3_X1  g0172(.A1(new_n260), .A2(KEYINPUT11), .A3(new_n367), .ZN(new_n373));
  OAI211_X1 g0173(.A(new_n272), .B(G68), .C1(G1), .C2(new_n220), .ZN(new_n374));
  NAND4_X1  g0174(.A1(new_n370), .A2(new_n372), .A3(new_n373), .A4(new_n374), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n365), .A2(new_n375), .ZN(new_n376));
  AOI21_X1  g0176(.A(new_n375), .B1(G190), .B2(new_n360), .ZN(new_n377));
  INV_X1    g0177(.A(G200), .ZN(new_n378));
  OAI21_X1  g0178(.A(new_n377), .B1(new_n378), .B2(new_n360), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n376), .A2(new_n379), .ZN(new_n380));
  NOR2_X1   g0180(.A1(new_n266), .A2(new_n312), .ZN(new_n381));
  AOI22_X1  g0181(.A1(new_n272), .A2(new_n381), .B1(new_n270), .B2(new_n266), .ZN(new_n382));
  AOI21_X1  g0182(.A(KEYINPUT7), .B1(new_n279), .B2(new_n220), .ZN(new_n383));
  INV_X1    g0183(.A(KEYINPUT7), .ZN(new_n384));
  NOR4_X1   g0184(.A1(new_n277), .A2(new_n278), .A3(new_n384), .A4(G20), .ZN(new_n385));
  OAI21_X1  g0185(.A(G68), .B1(new_n383), .B2(new_n385), .ZN(new_n386));
  NAND2_X1  g0186(.A1(G58), .A2(G68), .ZN(new_n387));
  AOI21_X1  g0187(.A(new_n220), .B1(new_n222), .B2(new_n387), .ZN(new_n388));
  INV_X1    g0188(.A(new_n388), .ZN(new_n389));
  INV_X1    g0189(.A(KEYINPUT71), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n261), .A2(G159), .ZN(new_n391));
  NAND3_X1  g0191(.A1(new_n389), .A2(new_n390), .A3(new_n391), .ZN(new_n392));
  INV_X1    g0192(.A(new_n391), .ZN(new_n393));
  OAI21_X1  g0193(.A(KEYINPUT71), .B1(new_n388), .B2(new_n393), .ZN(new_n394));
  NAND4_X1  g0194(.A1(new_n386), .A2(KEYINPUT16), .A3(new_n392), .A4(new_n394), .ZN(new_n395));
  NOR2_X1   g0195(.A1(new_n388), .A2(new_n393), .ZN(new_n396));
  AOI21_X1  g0196(.A(KEYINPUT16), .B1(new_n386), .B2(new_n396), .ZN(new_n397));
  INV_X1    g0197(.A(KEYINPUT72), .ZN(new_n398));
  OAI211_X1 g0198(.A(new_n260), .B(new_n395), .C1(new_n397), .C2(new_n398), .ZN(new_n399));
  INV_X1    g0199(.A(KEYINPUT16), .ZN(new_n400));
  OAI21_X1  g0200(.A(new_n384), .B1(new_n341), .B2(G20), .ZN(new_n401));
  NAND3_X1  g0201(.A1(new_n279), .A2(KEYINPUT7), .A3(new_n220), .ZN(new_n402));
  AOI21_X1  g0202(.A(new_n203), .B1(new_n401), .B2(new_n402), .ZN(new_n403));
  INV_X1    g0203(.A(new_n396), .ZN(new_n404));
  OAI211_X1 g0204(.A(new_n398), .B(new_n400), .C1(new_n403), .C2(new_n404), .ZN(new_n405));
  INV_X1    g0205(.A(new_n405), .ZN(new_n406));
  OAI21_X1  g0206(.A(new_n382), .B1(new_n399), .B2(new_n406), .ZN(new_n407));
  NAND2_X1  g0207(.A1(G33), .A2(G87), .ZN(new_n408));
  NOR2_X1   g0208(.A1(G223), .A2(G1698), .ZN(new_n409));
  AOI21_X1  g0209(.A(new_n409), .B1(new_n300), .B2(G1698), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n410), .A2(new_n341), .ZN(new_n411));
  AOI22_X1  g0211(.A1(new_n290), .A2(new_n292), .B1(new_n408), .B2(new_n411), .ZN(new_n412));
  OAI21_X1  g0212(.A(new_n299), .B1(new_n232), .B2(new_n301), .ZN(new_n413));
  OR2_X1    g0213(.A1(new_n412), .A2(new_n413), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n413), .A2(KEYINPUT73), .ZN(new_n415));
  INV_X1    g0215(.A(KEYINPUT73), .ZN(new_n416));
  OAI211_X1 g0216(.A(new_n299), .B(new_n416), .C1(new_n232), .C2(new_n301), .ZN(new_n417));
  AND2_X1   g0217(.A1(new_n415), .A2(new_n417), .ZN(new_n418));
  NOR2_X1   g0218(.A1(new_n412), .A2(G179), .ZN(new_n419));
  AOI22_X1  g0219(.A1(new_n414), .A2(new_n308), .B1(new_n418), .B2(new_n419), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n407), .A2(new_n420), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n421), .A2(KEYINPUT18), .ZN(new_n422));
  INV_X1    g0222(.A(KEYINPUT18), .ZN(new_n423));
  NAND3_X1  g0223(.A1(new_n407), .A2(new_n423), .A3(new_n420), .ZN(new_n424));
  OAI21_X1  g0224(.A(new_n378), .B1(new_n412), .B2(new_n413), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n411), .A2(new_n408), .ZN(new_n426));
  OAI21_X1  g0226(.A(new_n426), .B1(new_n351), .B2(new_n350), .ZN(new_n427));
  NAND4_X1  g0227(.A1(new_n427), .A2(new_n415), .A3(new_n303), .A4(new_n417), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n425), .A2(new_n428), .ZN(new_n429));
  OAI211_X1 g0229(.A(new_n429), .B(new_n382), .C1(new_n399), .C2(new_n406), .ZN(new_n430));
  INV_X1    g0230(.A(KEYINPUT17), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  OR2_X1    g0232(.A1(new_n397), .A2(new_n398), .ZN(new_n433));
  NAND4_X1  g0233(.A1(new_n433), .A2(new_n260), .A3(new_n405), .A4(new_n395), .ZN(new_n434));
  NAND4_X1  g0234(.A1(new_n434), .A2(KEYINPUT17), .A3(new_n382), .A4(new_n429), .ZN(new_n435));
  NAND4_X1  g0235(.A1(new_n422), .A2(new_n424), .A3(new_n432), .A4(new_n435), .ZN(new_n436));
  NOR3_X1   g0236(.A1(new_n340), .A2(new_n380), .A3(new_n436), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n233), .A2(G1698), .ZN(new_n438));
  OAI21_X1  g0238(.A(new_n438), .B1(G250), .B2(G1698), .ZN(new_n439));
  INV_X1    g0239(.A(G294), .ZN(new_n440));
  OAI22_X1  g0240(.A1(new_n439), .A2(new_n279), .B1(new_n256), .B2(new_n440), .ZN(new_n441));
  OAI21_X1  g0241(.A(new_n441), .B1(new_n351), .B2(new_n350), .ZN(new_n442));
  INV_X1    g0242(.A(KEYINPUT79), .ZN(new_n443));
  INV_X1    g0243(.A(G41), .ZN(new_n444));
  OAI21_X1  g0244(.A(new_n443), .B1(new_n444), .B2(KEYINPUT5), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n444), .A2(KEYINPUT5), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  INV_X1    g0247(.A(KEYINPUT5), .ZN(new_n448));
  NOR2_X1   g0248(.A1(new_n448), .A2(G41), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n449), .A2(new_n443), .ZN(new_n450));
  INV_X1    g0250(.A(G45), .ZN(new_n451));
  NOR2_X1   g0251(.A1(new_n451), .A2(G1), .ZN(new_n452));
  NAND4_X1  g0252(.A1(new_n330), .A2(new_n447), .A3(new_n450), .A4(new_n452), .ZN(new_n453));
  AOI21_X1  g0253(.A(KEYINPUT79), .B1(new_n448), .B2(G41), .ZN(new_n454));
  NOR2_X1   g0254(.A1(new_n454), .A2(new_n449), .ZN(new_n455));
  OAI21_X1  g0255(.A(new_n452), .B1(new_n446), .B2(KEYINPUT79), .ZN(new_n456));
  OAI211_X1 g0256(.A(G264), .B(new_n298), .C1(new_n455), .C2(new_n456), .ZN(new_n457));
  NAND3_X1  g0257(.A1(new_n442), .A2(new_n453), .A3(new_n457), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n458), .A2(G169), .ZN(new_n459));
  INV_X1    g0259(.A(KEYINPUT88), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  NAND3_X1  g0261(.A1(new_n458), .A2(KEYINPUT88), .A3(G169), .ZN(new_n462));
  OAI211_X1 g0262(.A(new_n461), .B(new_n462), .C1(new_n336), .C2(new_n458), .ZN(new_n463));
  OAI211_X1 g0263(.A(new_n220), .B(G87), .C1(new_n277), .C2(new_n278), .ZN(new_n464));
  OAI21_X1  g0264(.A(new_n464), .B1(KEYINPUT85), .B2(KEYINPUT22), .ZN(new_n465));
  NOR2_X1   g0265(.A1(KEYINPUT85), .A2(KEYINPUT22), .ZN(new_n466));
  NAND4_X1  g0266(.A1(new_n341), .A2(new_n220), .A3(G87), .A4(new_n466), .ZN(new_n467));
  NAND2_X1  g0267(.A1(KEYINPUT85), .A2(KEYINPUT22), .ZN(new_n468));
  NAND3_X1  g0268(.A1(new_n465), .A2(new_n467), .A3(new_n468), .ZN(new_n469));
  INV_X1    g0269(.A(KEYINPUT23), .ZN(new_n470));
  AOI21_X1  g0270(.A(new_n470), .B1(new_n323), .B2(G20), .ZN(new_n471));
  NOR3_X1   g0271(.A1(new_n220), .A2(KEYINPUT23), .A3(G107), .ZN(new_n472));
  INV_X1    g0272(.A(G116), .ZN(new_n473));
  INV_X1    g0273(.A(KEYINPUT86), .ZN(new_n474));
  INV_X1    g0274(.A(KEYINPUT24), .ZN(new_n475));
  OAI22_X1  g0275(.A1(new_n267), .A2(new_n473), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  NOR3_X1   g0276(.A1(new_n471), .A2(new_n472), .A3(new_n476), .ZN(new_n477));
  NAND4_X1  g0277(.A1(new_n469), .A2(new_n477), .A3(new_n474), .A4(new_n475), .ZN(new_n478));
  INV_X1    g0278(.A(new_n478), .ZN(new_n479));
  AOI22_X1  g0279(.A1(new_n469), .A2(new_n477), .B1(new_n474), .B2(new_n475), .ZN(new_n480));
  OAI21_X1  g0280(.A(new_n260), .B1(new_n479), .B2(new_n480), .ZN(new_n481));
  NOR2_X1   g0281(.A1(new_n269), .A2(G1), .ZN(new_n482));
  NAND3_X1  g0282(.A1(new_n482), .A2(G20), .A3(new_n207), .ZN(new_n483));
  XNOR2_X1  g0283(.A(new_n483), .B(KEYINPUT25), .ZN(new_n484));
  NOR2_X1   g0284(.A1(new_n256), .A2(G1), .ZN(new_n485));
  AOI211_X1 g0285(.A(new_n270), .B(new_n485), .C1(new_n258), .C2(new_n259), .ZN(new_n486));
  AOI21_X1  g0286(.A(new_n484), .B1(new_n486), .B2(G107), .ZN(new_n487));
  NAND3_X1  g0287(.A1(new_n481), .A2(KEYINPUT87), .A3(new_n487), .ZN(new_n488));
  INV_X1    g0288(.A(KEYINPUT87), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n258), .A2(new_n259), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n469), .A2(new_n477), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n474), .A2(new_n475), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  AOI21_X1  g0293(.A(new_n490), .B1(new_n493), .B2(new_n478), .ZN(new_n494));
  INV_X1    g0294(.A(new_n485), .ZN(new_n495));
  NAND3_X1  g0295(.A1(new_n272), .A2(G107), .A3(new_n495), .ZN(new_n496));
  INV_X1    g0296(.A(new_n484), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  OAI21_X1  g0298(.A(new_n489), .B1(new_n494), .B2(new_n498), .ZN(new_n499));
  NAND3_X1  g0299(.A1(new_n463), .A2(new_n488), .A3(new_n499), .ZN(new_n500));
  NAND3_X1  g0300(.A1(new_n272), .A2(G116), .A3(new_n495), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n473), .A2(G20), .ZN(new_n502));
  AND3_X1   g0302(.A1(KEYINPUT76), .A2(G33), .A3(G283), .ZN(new_n503));
  AOI21_X1  g0303(.A(KEYINPUT76), .B1(G33), .B2(G283), .ZN(new_n504));
  NOR2_X1   g0304(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  OAI21_X1  g0305(.A(new_n220), .B1(new_n206), .B2(G33), .ZN(new_n506));
  OAI211_X1 g0306(.A(new_n257), .B(new_n502), .C1(new_n505), .C2(new_n506), .ZN(new_n507));
  INV_X1    g0307(.A(KEYINPUT20), .ZN(new_n508));
  XNOR2_X1  g0308(.A(new_n507), .B(new_n508), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n270), .A2(new_n473), .ZN(new_n510));
  NAND3_X1  g0310(.A1(new_n501), .A2(new_n509), .A3(new_n510), .ZN(new_n511));
  OAI211_X1 g0311(.A(G270), .B(new_n298), .C1(new_n455), .C2(new_n456), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n453), .A2(new_n512), .ZN(new_n513));
  OAI211_X1 g0313(.A(G257), .B(new_n282), .C1(new_n277), .C2(new_n278), .ZN(new_n514));
  INV_X1    g0314(.A(G303), .ZN(new_n515));
  NOR3_X1   g0315(.A1(new_n277), .A2(new_n278), .A3(new_n515), .ZN(new_n516));
  OAI21_X1  g0316(.A(new_n514), .B1(new_n516), .B2(KEYINPUT82), .ZN(new_n517));
  INV_X1    g0317(.A(KEYINPUT82), .ZN(new_n518));
  NAND4_X1  g0318(.A1(new_n341), .A2(new_n518), .A3(G257), .A4(new_n282), .ZN(new_n519));
  OAI211_X1 g0319(.A(G264), .B(G1698), .C1(new_n277), .C2(new_n278), .ZN(new_n520));
  AND2_X1   g0320(.A1(new_n520), .A2(KEYINPUT83), .ZN(new_n521));
  NOR2_X1   g0321(.A1(new_n520), .A2(KEYINPUT83), .ZN(new_n522));
  OAI211_X1 g0322(.A(new_n517), .B(new_n519), .C1(new_n521), .C2(new_n522), .ZN(new_n523));
  AOI21_X1  g0323(.A(new_n513), .B1(new_n523), .B2(new_n293), .ZN(new_n524));
  INV_X1    g0324(.A(KEYINPUT21), .ZN(new_n525));
  NOR3_X1   g0325(.A1(new_n524), .A2(new_n525), .A3(new_n308), .ZN(new_n526));
  AOI211_X1 g0326(.A(new_n336), .B(new_n513), .C1(new_n293), .C2(new_n523), .ZN(new_n527));
  OAI21_X1  g0327(.A(new_n511), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  INV_X1    g0328(.A(KEYINPUT84), .ZN(new_n529));
  NOR2_X1   g0329(.A1(new_n524), .A2(new_n308), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n511), .A2(new_n530), .ZN(new_n531));
  AOI21_X1  g0331(.A(new_n529), .B1(new_n531), .B2(new_n525), .ZN(new_n532));
  AOI211_X1 g0332(.A(KEYINPUT84), .B(KEYINPUT21), .C1(new_n511), .C2(new_n530), .ZN(new_n533));
  OAI211_X1 g0333(.A(new_n500), .B(new_n528), .C1(new_n532), .C2(new_n533), .ZN(new_n534));
  INV_X1    g0334(.A(KEYINPUT6), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n535), .A2(KEYINPUT74), .ZN(new_n536));
  INV_X1    g0336(.A(KEYINPUT74), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n537), .A2(KEYINPUT6), .ZN(new_n538));
  NAND4_X1  g0338(.A1(new_n536), .A2(new_n538), .A3(G97), .A4(new_n207), .ZN(new_n539));
  INV_X1    g0339(.A(new_n539), .ZN(new_n540));
  NAND2_X1  g0340(.A1(G97), .A2(G107), .ZN(new_n541));
  AOI22_X1  g0341(.A1(new_n536), .A2(new_n538), .B1(new_n208), .B2(new_n541), .ZN(new_n542));
  OAI21_X1  g0342(.A(G20), .B1(new_n540), .B2(new_n542), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n261), .A2(G77), .ZN(new_n544));
  NAND3_X1  g0344(.A1(new_n543), .A2(KEYINPUT75), .A3(new_n544), .ZN(new_n545));
  OAI21_X1  g0345(.A(new_n324), .B1(new_n383), .B2(new_n385), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  AOI21_X1  g0347(.A(KEYINPUT75), .B1(new_n543), .B2(new_n544), .ZN(new_n548));
  OAI21_X1  g0348(.A(new_n260), .B1(new_n547), .B2(new_n548), .ZN(new_n549));
  NOR2_X1   g0349(.A1(new_n320), .A2(G97), .ZN(new_n550));
  AOI21_X1  g0350(.A(new_n550), .B1(new_n486), .B2(G97), .ZN(new_n551));
  AND2_X1   g0351(.A1(new_n549), .A2(new_n551), .ZN(new_n552));
  NAND4_X1  g0352(.A1(new_n341), .A2(KEYINPUT4), .A3(G244), .A4(new_n282), .ZN(new_n553));
  OAI211_X1 g0353(.A(G244), .B(new_n282), .C1(new_n277), .C2(new_n278), .ZN(new_n554));
  INV_X1    g0354(.A(KEYINPUT4), .ZN(new_n555));
  AOI21_X1  g0355(.A(new_n505), .B1(new_n554), .B2(new_n555), .ZN(new_n556));
  OAI211_X1 g0356(.A(G250), .B(G1698), .C1(new_n277), .C2(new_n278), .ZN(new_n557));
  AND2_X1   g0357(.A1(new_n557), .A2(KEYINPUT77), .ZN(new_n558));
  NOR2_X1   g0358(.A1(new_n557), .A2(KEYINPUT77), .ZN(new_n559));
  OAI211_X1 g0359(.A(new_n553), .B(new_n556), .C1(new_n558), .C2(new_n559), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n560), .A2(new_n293), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n561), .A2(KEYINPUT78), .ZN(new_n562));
  OAI211_X1 g0362(.A(G257), .B(new_n298), .C1(new_n455), .C2(new_n456), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n453), .A2(new_n563), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n564), .A2(KEYINPUT80), .ZN(new_n565));
  INV_X1    g0365(.A(KEYINPUT80), .ZN(new_n566));
  NAND3_X1  g0366(.A1(new_n453), .A2(new_n563), .A3(new_n566), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n565), .A2(new_n567), .ZN(new_n568));
  INV_X1    g0368(.A(KEYINPUT78), .ZN(new_n569));
  NAND3_X1  g0369(.A1(new_n560), .A2(new_n569), .A3(new_n293), .ZN(new_n570));
  NAND3_X1  g0370(.A1(new_n562), .A2(new_n568), .A3(new_n570), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n571), .A2(G200), .ZN(new_n572));
  AOI21_X1  g0372(.A(new_n564), .B1(new_n560), .B2(new_n293), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n573), .A2(G190), .ZN(new_n574));
  NAND3_X1  g0374(.A1(new_n552), .A2(new_n572), .A3(new_n574), .ZN(new_n575));
  NOR2_X1   g0375(.A1(G87), .A2(G97), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n323), .A2(new_n576), .ZN(new_n577));
  INV_X1    g0377(.A(KEYINPUT19), .ZN(new_n578));
  OAI21_X1  g0378(.A(new_n220), .B1(new_n344), .B2(new_n578), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n577), .A2(new_n579), .ZN(new_n580));
  NAND3_X1  g0380(.A1(new_n341), .A2(new_n220), .A3(G68), .ZN(new_n581));
  OAI21_X1  g0381(.A(new_n578), .B1(new_n267), .B2(new_n206), .ZN(new_n582));
  NAND3_X1  g0382(.A1(new_n580), .A2(new_n581), .A3(new_n582), .ZN(new_n583));
  INV_X1    g0383(.A(KEYINPUT81), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  NAND4_X1  g0385(.A1(new_n580), .A2(KEYINPUT81), .A3(new_n581), .A4(new_n582), .ZN(new_n586));
  NAND3_X1  g0386(.A1(new_n260), .A2(new_n585), .A3(new_n586), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n315), .A2(new_n270), .ZN(new_n588));
  NAND3_X1  g0388(.A1(new_n272), .A2(G87), .A3(new_n495), .ZN(new_n589));
  AND3_X1   g0389(.A1(new_n587), .A2(new_n588), .A3(new_n589), .ZN(new_n590));
  OAI211_X1 g0390(.A(G238), .B(new_n282), .C1(new_n277), .C2(new_n278), .ZN(new_n591));
  OAI211_X1 g0391(.A(G244), .B(G1698), .C1(new_n277), .C2(new_n278), .ZN(new_n592));
  OAI211_X1 g0392(.A(new_n591), .B(new_n592), .C1(new_n256), .C2(new_n473), .ZN(new_n593));
  OAI21_X1  g0393(.A(new_n593), .B1(new_n350), .B2(new_n351), .ZN(new_n594));
  NOR2_X1   g0394(.A1(new_n452), .A2(new_n229), .ZN(new_n595));
  AOI22_X1  g0395(.A1(new_n330), .A2(new_n452), .B1(new_n298), .B2(new_n595), .ZN(new_n596));
  AOI21_X1  g0396(.A(new_n378), .B1(new_n594), .B2(new_n596), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n594), .A2(new_n596), .ZN(new_n598));
  INV_X1    g0398(.A(new_n598), .ZN(new_n599));
  AOI21_X1  g0399(.A(new_n597), .B1(new_n599), .B2(G190), .ZN(new_n600));
  INV_X1    g0400(.A(new_n315), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n486), .A2(new_n601), .ZN(new_n602));
  NAND3_X1  g0402(.A1(new_n602), .A2(new_n587), .A3(new_n588), .ZN(new_n603));
  AOI21_X1  g0403(.A(G169), .B1(new_n594), .B2(new_n596), .ZN(new_n604));
  AOI21_X1  g0404(.A(new_n604), .B1(new_n599), .B2(new_n336), .ZN(new_n605));
  AOI22_X1  g0405(.A1(new_n590), .A2(new_n600), .B1(new_n603), .B2(new_n605), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n549), .A2(new_n551), .ZN(new_n607));
  OR2_X1    g0407(.A1(new_n573), .A2(G169), .ZN(new_n608));
  OAI211_X1 g0408(.A(new_n607), .B(new_n608), .C1(G179), .C2(new_n571), .ZN(new_n609));
  AND2_X1   g0409(.A1(new_n458), .A2(new_n378), .ZN(new_n610));
  NOR2_X1   g0410(.A1(new_n458), .A2(G190), .ZN(new_n611));
  OAI211_X1 g0411(.A(new_n481), .B(new_n487), .C1(new_n610), .C2(new_n611), .ZN(new_n612));
  NAND4_X1  g0412(.A1(new_n575), .A2(new_n606), .A3(new_n609), .A4(new_n612), .ZN(new_n613));
  INV_X1    g0413(.A(new_n524), .ZN(new_n614));
  NOR2_X1   g0414(.A1(new_n614), .A2(new_n303), .ZN(new_n615));
  AOI211_X1 g0415(.A(new_n511), .B(new_n615), .C1(G200), .C2(new_n614), .ZN(new_n616));
  NOR3_X1   g0416(.A1(new_n534), .A2(new_n613), .A3(new_n616), .ZN(new_n617));
  AND2_X1   g0417(.A1(new_n437), .A2(new_n617), .ZN(G372));
  AND2_X1   g0418(.A1(new_n435), .A2(new_n432), .ZN(new_n619));
  INV_X1    g0419(.A(new_n619), .ZN(new_n620));
  INV_X1    g0420(.A(new_n339), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n379), .A2(new_n621), .ZN(new_n622));
  AOI21_X1  g0422(.A(new_n620), .B1(new_n622), .B2(new_n376), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n422), .A2(new_n424), .ZN(new_n624));
  INV_X1    g0424(.A(KEYINPUT89), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  NAND3_X1  g0426(.A1(new_n422), .A2(KEYINPUT89), .A3(new_n424), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  OAI21_X1  g0428(.A(new_n307), .B1(new_n623), .B2(new_n628), .ZN(new_n629));
  AND2_X1   g0429(.A1(new_n629), .A2(new_n310), .ZN(new_n630));
  INV_X1    g0430(.A(new_n437), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n590), .A2(new_n600), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n603), .A2(new_n605), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  INV_X1    g0434(.A(KEYINPUT26), .ZN(new_n635));
  OR3_X1    g0435(.A1(new_n634), .A2(new_n609), .A3(new_n635), .ZN(new_n636));
  OAI21_X1  g0436(.A(new_n635), .B1(new_n634), .B2(new_n609), .ZN(new_n637));
  AOI22_X1  g0437(.A1(new_n636), .A2(new_n637), .B1(new_n603), .B2(new_n605), .ZN(new_n638));
  INV_X1    g0438(.A(new_n613), .ZN(new_n639));
  OAI21_X1  g0439(.A(new_n528), .B1(new_n532), .B2(new_n533), .ZN(new_n640));
  OAI21_X1  g0440(.A(new_n463), .B1(new_n494), .B2(new_n498), .ZN(new_n641));
  INV_X1    g0441(.A(new_n641), .ZN(new_n642));
  OAI21_X1  g0442(.A(new_n639), .B1(new_n640), .B2(new_n642), .ZN(new_n643));
  AND2_X1   g0443(.A1(new_n638), .A2(new_n643), .ZN(new_n644));
  OAI21_X1  g0444(.A(new_n630), .B1(new_n631), .B2(new_n644), .ZN(G369));
  INV_X1    g0445(.A(KEYINPUT27), .ZN(new_n646));
  NAND3_X1  g0446(.A1(new_n482), .A2(new_n646), .A3(new_n220), .ZN(new_n647));
  XNOR2_X1  g0447(.A(new_n647), .B(KEYINPUT90), .ZN(new_n648));
  INV_X1    g0448(.A(G213), .ZN(new_n649));
  AOI21_X1  g0449(.A(new_n646), .B1(new_n482), .B2(new_n220), .ZN(new_n650));
  NOR3_X1   g0450(.A1(new_n648), .A2(new_n649), .A3(new_n650), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n651), .A2(G343), .ZN(new_n652));
  INV_X1    g0452(.A(new_n652), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n511), .A2(new_n653), .ZN(new_n654));
  XNOR2_X1  g0454(.A(new_n640), .B(new_n654), .ZN(new_n655));
  NOR2_X1   g0455(.A1(new_n655), .A2(new_n616), .ZN(new_n656));
  XNOR2_X1  g0456(.A(KEYINPUT91), .B(G330), .ZN(new_n657));
  INV_X1    g0457(.A(new_n657), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n656), .A2(new_n658), .ZN(new_n659));
  INV_X1    g0459(.A(new_n659), .ZN(new_n660));
  OR2_X1    g0460(.A1(new_n500), .A2(new_n652), .ZN(new_n661));
  NAND3_X1  g0461(.A1(new_n488), .A2(new_n499), .A3(new_n653), .ZN(new_n662));
  NAND3_X1  g0462(.A1(new_n500), .A2(new_n662), .A3(new_n612), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n661), .A2(new_n663), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n660), .A2(new_n664), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n640), .A2(new_n652), .ZN(new_n666));
  NOR2_X1   g0466(.A1(new_n666), .A2(new_n663), .ZN(new_n667));
  XNOR2_X1  g0467(.A(new_n652), .B(KEYINPUT92), .ZN(new_n668));
  INV_X1    g0468(.A(new_n668), .ZN(new_n669));
  AOI21_X1  g0469(.A(new_n667), .B1(new_n642), .B2(new_n669), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n665), .A2(new_n670), .ZN(G399));
  INV_X1    g0471(.A(new_n211), .ZN(new_n672));
  NOR2_X1   g0472(.A1(new_n672), .A2(G41), .ZN(new_n673));
  INV_X1    g0473(.A(new_n673), .ZN(new_n674));
  NOR2_X1   g0474(.A1(new_n577), .A2(G116), .ZN(new_n675));
  NAND3_X1  g0475(.A1(new_n674), .A2(new_n675), .A3(G1), .ZN(new_n676));
  OAI21_X1  g0476(.A(new_n676), .B1(new_n223), .B2(new_n674), .ZN(new_n677));
  XNOR2_X1  g0477(.A(new_n677), .B(KEYINPUT28), .ZN(new_n678));
  NOR3_X1   g0478(.A1(new_n644), .A2(KEYINPUT29), .A3(new_n668), .ZN(new_n679));
  AND2_X1   g0479(.A1(new_n638), .A2(KEYINPUT93), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n639), .A2(new_n534), .ZN(new_n681));
  OAI21_X1  g0481(.A(new_n681), .B1(new_n638), .B2(KEYINPUT93), .ZN(new_n682));
  OAI21_X1  g0482(.A(new_n652), .B1(new_n680), .B2(new_n682), .ZN(new_n683));
  AOI21_X1  g0483(.A(new_n679), .B1(new_n683), .B2(KEYINPUT29), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n617), .A2(new_n669), .ZN(new_n685));
  AND4_X1   g0485(.A1(new_n594), .A2(new_n442), .A3(new_n596), .A4(new_n457), .ZN(new_n686));
  NAND4_X1  g0486(.A1(new_n686), .A2(new_n573), .A3(new_n524), .A4(G179), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n687), .A2(KEYINPUT30), .ZN(new_n688));
  INV_X1    g0488(.A(KEYINPUT30), .ZN(new_n689));
  NAND4_X1  g0489(.A1(new_n527), .A2(new_n689), .A3(new_n573), .A4(new_n686), .ZN(new_n690));
  NAND3_X1  g0490(.A1(new_n458), .A2(new_n598), .A3(new_n336), .ZN(new_n691));
  NOR2_X1   g0491(.A1(new_n691), .A2(new_n524), .ZN(new_n692));
  AOI22_X1  g0492(.A1(new_n688), .A2(new_n690), .B1(new_n692), .B2(new_n571), .ZN(new_n693));
  INV_X1    g0493(.A(KEYINPUT31), .ZN(new_n694));
  NOR3_X1   g0494(.A1(new_n693), .A2(new_n694), .A3(new_n669), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n688), .A2(new_n690), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n692), .A2(new_n571), .ZN(new_n697));
  AOI21_X1  g0497(.A(new_n652), .B1(new_n696), .B2(new_n697), .ZN(new_n698));
  INV_X1    g0498(.A(new_n698), .ZN(new_n699));
  AOI21_X1  g0499(.A(new_n695), .B1(new_n694), .B2(new_n699), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n685), .A2(new_n700), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n701), .A2(new_n658), .ZN(new_n702));
  AND2_X1   g0502(.A1(new_n684), .A2(new_n702), .ZN(new_n703));
  OAI21_X1  g0503(.A(new_n678), .B1(new_n703), .B2(G1), .ZN(G364));
  NOR2_X1   g0504(.A1(new_n269), .A2(G20), .ZN(new_n705));
  AOI21_X1  g0505(.A(new_n295), .B1(new_n705), .B2(G45), .ZN(new_n706));
  INV_X1    g0506(.A(new_n706), .ZN(new_n707));
  NOR2_X1   g0507(.A1(new_n673), .A2(new_n707), .ZN(new_n708));
  NOR2_X1   g0508(.A1(new_n660), .A2(new_n708), .ZN(new_n709));
  NOR2_X1   g0509(.A1(new_n656), .A2(new_n658), .ZN(new_n710));
  INV_X1    g0510(.A(new_n710), .ZN(new_n711));
  NOR2_X1   g0511(.A1(G13), .A2(G33), .ZN(new_n712));
  INV_X1    g0512(.A(new_n712), .ZN(new_n713));
  NOR2_X1   g0513(.A1(new_n713), .A2(G20), .ZN(new_n714));
  OAI21_X1  g0514(.A(new_n714), .B1(new_n655), .B2(new_n616), .ZN(new_n715));
  AOI21_X1  g0515(.A(new_n219), .B1(G20), .B2(new_n308), .ZN(new_n716));
  NOR2_X1   g0516(.A1(new_n220), .A2(G179), .ZN(new_n717));
  NOR2_X1   g0517(.A1(G190), .A2(G200), .ZN(new_n718));
  AND2_X1   g0518(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  OR2_X1    g0519(.A1(new_n719), .A2(KEYINPUT95), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n719), .A2(KEYINPUT95), .ZN(new_n721));
  NAND2_X1  g0521(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  INV_X1    g0522(.A(new_n722), .ZN(new_n723));
  AND2_X1   g0523(.A1(new_n723), .A2(G329), .ZN(new_n724));
  NOR3_X1   g0524(.A1(new_n303), .A2(G179), .A3(G200), .ZN(new_n725));
  NOR2_X1   g0525(.A1(new_n725), .A2(new_n220), .ZN(new_n726));
  INV_X1    g0526(.A(new_n726), .ZN(new_n727));
  NAND3_X1  g0527(.A1(new_n717), .A2(G190), .A3(G200), .ZN(new_n728));
  INV_X1    g0528(.A(new_n728), .ZN(new_n729));
  AOI22_X1  g0529(.A1(new_n727), .A2(G294), .B1(new_n729), .B2(G303), .ZN(new_n730));
  INV_X1    g0530(.A(G283), .ZN(new_n731));
  NAND3_X1  g0531(.A1(new_n717), .A2(new_n303), .A3(G200), .ZN(new_n732));
  OAI21_X1  g0532(.A(new_n730), .B1(new_n731), .B2(new_n732), .ZN(new_n733));
  NAND2_X1  g0533(.A1(G20), .A2(G179), .ZN(new_n734));
  NOR3_X1   g0534(.A1(new_n734), .A2(new_n303), .A3(G200), .ZN(new_n735));
  NAND2_X1  g0535(.A1(new_n735), .A2(G322), .ZN(new_n736));
  INV_X1    g0536(.A(G311), .ZN(new_n737));
  INV_X1    g0537(.A(new_n734), .ZN(new_n738));
  NAND2_X1  g0538(.A1(new_n738), .A2(new_n718), .ZN(new_n739));
  OAI211_X1 g0539(.A(new_n736), .B(new_n279), .C1(new_n737), .C2(new_n739), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n738), .A2(G200), .ZN(new_n741));
  NOR2_X1   g0541(.A1(new_n741), .A2(G190), .ZN(new_n742));
  INV_X1    g0542(.A(new_n742), .ZN(new_n743));
  XOR2_X1   g0543(.A(KEYINPUT33), .B(G317), .Z(new_n744));
  NOR2_X1   g0544(.A1(new_n741), .A2(new_n303), .ZN(new_n745));
  INV_X1    g0545(.A(new_n745), .ZN(new_n746));
  INV_X1    g0546(.A(G326), .ZN(new_n747));
  OAI22_X1  g0547(.A1(new_n743), .A2(new_n744), .B1(new_n746), .B2(new_n747), .ZN(new_n748));
  NOR4_X1   g0548(.A1(new_n724), .A2(new_n733), .A3(new_n740), .A4(new_n748), .ZN(new_n749));
  XOR2_X1   g0549(.A(new_n749), .B(KEYINPUT97), .Z(new_n750));
  INV_X1    g0550(.A(G159), .ZN(new_n751));
  NOR2_X1   g0551(.A1(new_n722), .A2(new_n751), .ZN(new_n752));
  XNOR2_X1  g0552(.A(new_n752), .B(KEYINPUT32), .ZN(new_n753));
  XOR2_X1   g0553(.A(new_n726), .B(KEYINPUT96), .Z(new_n754));
  NAND2_X1  g0554(.A1(new_n754), .A2(G97), .ZN(new_n755));
  OAI21_X1  g0555(.A(new_n341), .B1(new_n739), .B2(new_n311), .ZN(new_n756));
  AOI21_X1  g0556(.A(new_n756), .B1(G58), .B2(new_n735), .ZN(new_n757));
  NOR2_X1   g0557(.A1(new_n732), .A2(new_n207), .ZN(new_n758));
  OAI22_X1  g0558(.A1(new_n201), .A2(new_n746), .B1(new_n743), .B2(new_n203), .ZN(new_n759));
  AOI211_X1 g0559(.A(new_n758), .B(new_n759), .C1(G87), .C2(new_n729), .ZN(new_n760));
  AND4_X1   g0560(.A1(new_n753), .A2(new_n755), .A3(new_n757), .A4(new_n760), .ZN(new_n761));
  OAI21_X1  g0561(.A(new_n716), .B1(new_n750), .B2(new_n761), .ZN(new_n762));
  NOR2_X1   g0562(.A1(new_n716), .A2(new_n714), .ZN(new_n763));
  NOR2_X1   g0563(.A1(new_n672), .A2(new_n341), .ZN(new_n764));
  INV_X1    g0564(.A(new_n764), .ZN(new_n765));
  NOR2_X1   g0565(.A1(new_n254), .A2(new_n451), .ZN(new_n766));
  XNOR2_X1  g0566(.A(new_n766), .B(KEYINPUT94), .ZN(new_n767));
  AOI211_X1 g0567(.A(new_n765), .B(new_n767), .C1(new_n451), .C2(new_n224), .ZN(new_n768));
  NAND2_X1  g0568(.A1(new_n341), .A2(new_n211), .ZN(new_n769));
  INV_X1    g0569(.A(G355), .ZN(new_n770));
  OAI22_X1  g0570(.A1(new_n769), .A2(new_n770), .B1(G116), .B2(new_n211), .ZN(new_n771));
  OAI21_X1  g0571(.A(new_n763), .B1(new_n768), .B2(new_n771), .ZN(new_n772));
  AND3_X1   g0572(.A1(new_n762), .A2(new_n708), .A3(new_n772), .ZN(new_n773));
  AOI22_X1  g0573(.A1(new_n709), .A2(new_n711), .B1(new_n715), .B2(new_n773), .ZN(new_n774));
  INV_X1    g0574(.A(new_n774), .ZN(G396));
  AOI21_X1  g0575(.A(new_n668), .B1(new_n638), .B2(new_n643), .ZN(new_n776));
  NOR2_X1   g0576(.A1(new_n339), .A2(new_n653), .ZN(new_n777));
  OAI21_X1  g0577(.A(new_n334), .B1(new_n322), .B2(new_n652), .ZN(new_n778));
  AOI21_X1  g0578(.A(new_n777), .B1(new_n778), .B2(new_n339), .ZN(new_n779));
  XNOR2_X1  g0579(.A(new_n776), .B(new_n779), .ZN(new_n780));
  AOI21_X1  g0580(.A(new_n708), .B1(new_n780), .B2(new_n702), .ZN(new_n781));
  OAI21_X1  g0581(.A(new_n781), .B1(new_n702), .B2(new_n780), .ZN(new_n782));
  INV_X1    g0582(.A(new_n708), .ZN(new_n783));
  NOR2_X1   g0583(.A1(new_n716), .A2(new_n712), .ZN(new_n784));
  AOI21_X1  g0584(.A(new_n783), .B1(new_n784), .B2(new_n311), .ZN(new_n785));
  INV_X1    g0585(.A(new_n716), .ZN(new_n786));
  INV_X1    g0586(.A(new_n739), .ZN(new_n787));
  AOI22_X1  g0587(.A1(new_n787), .A2(G159), .B1(G143), .B2(new_n735), .ZN(new_n788));
  INV_X1    g0588(.A(G137), .ZN(new_n789));
  INV_X1    g0589(.A(G150), .ZN(new_n790));
  OAI221_X1 g0590(.A(new_n788), .B1(new_n746), .B2(new_n789), .C1(new_n790), .C2(new_n743), .ZN(new_n791));
  INV_X1    g0591(.A(KEYINPUT34), .ZN(new_n792));
  OR2_X1    g0592(.A1(new_n791), .A2(new_n792), .ZN(new_n793));
  NAND2_X1  g0593(.A1(new_n791), .A2(new_n792), .ZN(new_n794));
  NAND2_X1  g0594(.A1(new_n723), .A2(G132), .ZN(new_n795));
  OAI22_X1  g0595(.A1(new_n726), .A2(new_n202), .B1(new_n728), .B2(new_n201), .ZN(new_n796));
  NOR2_X1   g0596(.A1(new_n732), .A2(new_n203), .ZN(new_n797));
  NOR3_X1   g0597(.A1(new_n796), .A2(new_n279), .A3(new_n797), .ZN(new_n798));
  NAND4_X1  g0598(.A1(new_n793), .A2(new_n794), .A3(new_n795), .A4(new_n798), .ZN(new_n799));
  NAND2_X1  g0599(.A1(new_n723), .A2(G311), .ZN(new_n800));
  OAI22_X1  g0600(.A1(new_n746), .A2(new_n515), .B1(new_n732), .B2(new_n228), .ZN(new_n801));
  OAI22_X1  g0601(.A1(new_n743), .A2(new_n731), .B1(new_n728), .B2(new_n207), .ZN(new_n802));
  NOR2_X1   g0602(.A1(new_n801), .A2(new_n802), .ZN(new_n803));
  OAI21_X1  g0603(.A(new_n279), .B1(new_n739), .B2(new_n473), .ZN(new_n804));
  AOI21_X1  g0604(.A(new_n804), .B1(G294), .B2(new_n735), .ZN(new_n805));
  NAND4_X1  g0605(.A1(new_n800), .A2(new_n803), .A3(new_n755), .A4(new_n805), .ZN(new_n806));
  AND2_X1   g0606(.A1(new_n799), .A2(new_n806), .ZN(new_n807));
  OAI221_X1 g0607(.A(new_n785), .B1(new_n786), .B2(new_n807), .C1(new_n779), .C2(new_n713), .ZN(new_n808));
  AND2_X1   g0608(.A1(new_n782), .A2(new_n808), .ZN(new_n809));
  INV_X1    g0609(.A(new_n809), .ZN(G384));
  NOR2_X1   g0610(.A1(new_n705), .A2(new_n295), .ZN(new_n811));
  INV_X1    g0611(.A(KEYINPUT106), .ZN(new_n812));
  NAND2_X1  g0612(.A1(new_n392), .A2(new_n394), .ZN(new_n813));
  OAI21_X1  g0613(.A(new_n400), .B1(new_n813), .B2(new_n403), .ZN(new_n814));
  NAND3_X1  g0614(.A1(new_n814), .A2(new_n260), .A3(new_n395), .ZN(new_n815));
  NAND2_X1  g0615(.A1(new_n815), .A2(new_n382), .ZN(new_n816));
  NAND2_X1  g0616(.A1(new_n420), .A2(new_n816), .ZN(new_n817));
  NAND3_X1  g0617(.A1(new_n817), .A2(new_n430), .A3(KEYINPUT101), .ZN(new_n818));
  NAND2_X1  g0618(.A1(new_n816), .A2(new_n651), .ZN(new_n819));
  NAND2_X1  g0619(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  AOI21_X1  g0620(.A(KEYINPUT101), .B1(new_n817), .B2(new_n430), .ZN(new_n821));
  OAI21_X1  g0621(.A(KEYINPUT37), .B1(new_n820), .B2(new_n821), .ZN(new_n822));
  XNOR2_X1  g0622(.A(new_n651), .B(KEYINPUT102), .ZN(new_n823));
  NAND2_X1  g0623(.A1(new_n407), .A2(new_n823), .ZN(new_n824));
  NAND3_X1  g0624(.A1(new_n824), .A2(new_n421), .A3(new_n430), .ZN(new_n825));
  XNOR2_X1  g0625(.A(KEYINPUT103), .B(KEYINPUT37), .ZN(new_n826));
  OR2_X1    g0626(.A1(new_n825), .A2(new_n826), .ZN(new_n827));
  NAND2_X1  g0627(.A1(new_n822), .A2(new_n827), .ZN(new_n828));
  INV_X1    g0628(.A(new_n819), .ZN(new_n829));
  AND3_X1   g0629(.A1(new_n436), .A2(KEYINPUT100), .A3(new_n829), .ZN(new_n830));
  AOI21_X1  g0630(.A(KEYINPUT100), .B1(new_n436), .B2(new_n829), .ZN(new_n831));
  OAI21_X1  g0631(.A(new_n828), .B1(new_n830), .B2(new_n831), .ZN(new_n832));
  INV_X1    g0632(.A(KEYINPUT38), .ZN(new_n833));
  NAND2_X1  g0633(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  OAI211_X1 g0634(.A(new_n828), .B(KEYINPUT38), .C1(new_n830), .C2(new_n831), .ZN(new_n835));
  NAND2_X1  g0635(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  NAND2_X1  g0636(.A1(new_n375), .A2(new_n653), .ZN(new_n837));
  INV_X1    g0637(.A(KEYINPUT99), .ZN(new_n838));
  XNOR2_X1  g0638(.A(new_n837), .B(new_n838), .ZN(new_n839));
  INV_X1    g0639(.A(new_n839), .ZN(new_n840));
  NAND2_X1  g0640(.A1(new_n380), .A2(new_n840), .ZN(new_n841));
  NAND3_X1  g0641(.A1(new_n839), .A2(new_n376), .A3(new_n379), .ZN(new_n842));
  NAND3_X1  g0642(.A1(new_n841), .A2(new_n779), .A3(new_n842), .ZN(new_n843));
  INV_X1    g0643(.A(KEYINPUT104), .ZN(new_n844));
  OAI21_X1  g0644(.A(new_n694), .B1(new_n698), .B2(new_n844), .ZN(new_n845));
  NOR3_X1   g0645(.A1(new_n693), .A2(KEYINPUT104), .A3(new_n652), .ZN(new_n846));
  OAI21_X1  g0646(.A(KEYINPUT105), .B1(new_n845), .B2(new_n846), .ZN(new_n847));
  NAND2_X1  g0647(.A1(new_n698), .A2(new_n844), .ZN(new_n848));
  OAI21_X1  g0648(.A(KEYINPUT104), .B1(new_n693), .B2(new_n652), .ZN(new_n849));
  INV_X1    g0649(.A(KEYINPUT105), .ZN(new_n850));
  NAND4_X1  g0650(.A1(new_n848), .A2(new_n849), .A3(new_n850), .A4(new_n694), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n847), .A2(new_n851), .ZN(new_n852));
  NOR2_X1   g0652(.A1(new_n699), .A2(new_n694), .ZN(new_n853));
  AOI21_X1  g0653(.A(new_n853), .B1(new_n617), .B2(new_n669), .ZN(new_n854));
  AOI21_X1  g0654(.A(new_n843), .B1(new_n852), .B2(new_n854), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n836), .A2(new_n855), .ZN(new_n856));
  INV_X1    g0656(.A(KEYINPUT40), .ZN(new_n857));
  AOI21_X1  g0657(.A(new_n812), .B1(new_n856), .B2(new_n857), .ZN(new_n858));
  AOI211_X1 g0658(.A(KEYINPUT106), .B(KEYINPUT40), .C1(new_n836), .C2(new_n855), .ZN(new_n859));
  OR2_X1    g0659(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  INV_X1    g0660(.A(new_n824), .ZN(new_n861));
  OAI21_X1  g0661(.A(new_n861), .B1(new_n628), .B2(new_n620), .ZN(new_n862));
  XNOR2_X1  g0662(.A(new_n825), .B(new_n826), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n864), .A2(new_n833), .ZN(new_n865));
  AOI21_X1  g0665(.A(new_n857), .B1(new_n865), .B2(new_n835), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n866), .A2(new_n855), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n860), .A2(new_n867), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n852), .A2(new_n854), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n437), .A2(new_n869), .ZN(new_n870));
  XNOR2_X1  g0670(.A(new_n870), .B(KEYINPUT107), .ZN(new_n871));
  OR2_X1    g0671(.A1(new_n868), .A2(new_n871), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n872), .A2(new_n658), .ZN(new_n873));
  AOI21_X1  g0673(.A(new_n873), .B1(new_n868), .B2(new_n871), .ZN(new_n874));
  INV_X1    g0674(.A(new_n874), .ZN(new_n875));
  NAND3_X1  g0675(.A1(new_n834), .A2(KEYINPUT39), .A3(new_n835), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n865), .A2(new_n835), .ZN(new_n877));
  INV_X1    g0677(.A(KEYINPUT39), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n877), .A2(new_n878), .ZN(new_n879));
  NOR2_X1   g0679(.A1(new_n376), .A2(new_n653), .ZN(new_n880));
  NAND3_X1  g0680(.A1(new_n876), .A2(new_n879), .A3(new_n880), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n778), .A2(new_n339), .ZN(new_n882));
  AOI21_X1  g0682(.A(new_n777), .B1(new_n776), .B2(new_n882), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n841), .A2(new_n842), .ZN(new_n884));
  NOR2_X1   g0684(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  INV_X1    g0685(.A(new_n823), .ZN(new_n886));
  AOI22_X1  g0686(.A1(new_n885), .A2(new_n836), .B1(new_n628), .B2(new_n886), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n881), .A2(new_n887), .ZN(new_n888));
  OAI21_X1  g0688(.A(new_n630), .B1(new_n684), .B2(new_n631), .ZN(new_n889));
  XNOR2_X1  g0689(.A(new_n888), .B(new_n889), .ZN(new_n890));
  AOI21_X1  g0690(.A(new_n811), .B1(new_n875), .B2(new_n890), .ZN(new_n891));
  OAI21_X1  g0691(.A(new_n891), .B1(new_n890), .B2(new_n875), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n536), .A2(new_n538), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n208), .A2(new_n541), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n895), .A2(new_n539), .ZN(new_n896));
  OR2_X1    g0696(.A1(new_n896), .A2(KEYINPUT35), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n896), .A2(KEYINPUT35), .ZN(new_n898));
  NAND4_X1  g0698(.A1(new_n897), .A2(G116), .A3(new_n221), .A4(new_n898), .ZN(new_n899));
  XOR2_X1   g0699(.A(KEYINPUT98), .B(KEYINPUT36), .Z(new_n900));
  XNOR2_X1  g0700(.A(new_n899), .B(new_n900), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n387), .A2(G77), .ZN(new_n902));
  OAI21_X1  g0702(.A(new_n250), .B1(new_n223), .B2(new_n902), .ZN(new_n903));
  NAND3_X1  g0703(.A1(new_n903), .A2(G1), .A3(new_n269), .ZN(new_n904));
  NAND3_X1  g0704(.A1(new_n892), .A2(new_n901), .A3(new_n904), .ZN(G367));
  XOR2_X1   g0705(.A(new_n673), .B(KEYINPUT41), .Z(new_n906));
  INV_X1    g0706(.A(new_n906), .ZN(new_n907));
  INV_X1    g0707(.A(new_n664), .ZN(new_n908));
  AOI21_X1  g0708(.A(new_n667), .B1(new_n908), .B2(new_n666), .ZN(new_n909));
  XNOR2_X1  g0709(.A(new_n659), .B(new_n909), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n703), .A2(new_n910), .ZN(new_n911));
  OAI211_X1 g0711(.A(new_n575), .B(new_n609), .C1(new_n552), .C2(new_n669), .ZN(new_n912));
  OR2_X1    g0712(.A1(new_n609), .A2(new_n669), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n670), .A2(new_n914), .ZN(new_n915));
  XOR2_X1   g0715(.A(new_n915), .B(KEYINPUT45), .Z(new_n916));
  NOR2_X1   g0716(.A1(new_n670), .A2(new_n914), .ZN(new_n917));
  XNOR2_X1  g0717(.A(new_n917), .B(KEYINPUT44), .ZN(new_n918));
  NAND3_X1  g0718(.A1(new_n660), .A2(KEYINPUT110), .A3(new_n664), .ZN(new_n919));
  NAND3_X1  g0719(.A1(new_n916), .A2(new_n918), .A3(new_n919), .ZN(new_n920));
  INV_X1    g0720(.A(KEYINPUT110), .ZN(new_n921));
  NAND3_X1  g0721(.A1(new_n920), .A2(new_n921), .A3(new_n665), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n665), .A2(new_n921), .ZN(new_n923));
  NAND4_X1  g0723(.A1(new_n916), .A2(new_n923), .A3(new_n918), .A4(new_n919), .ZN(new_n924));
  AOI21_X1  g0724(.A(new_n911), .B1(new_n922), .B2(new_n924), .ZN(new_n925));
  INV_X1    g0725(.A(new_n703), .ZN(new_n926));
  OAI21_X1  g0726(.A(new_n907), .B1(new_n925), .B2(new_n926), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n927), .A2(new_n706), .ZN(new_n928));
  OAI21_X1  g0728(.A(new_n606), .B1(new_n590), .B2(new_n652), .ZN(new_n929));
  OR3_X1    g0729(.A1(new_n633), .A2(new_n590), .A3(new_n652), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  INV_X1    g0731(.A(new_n931), .ZN(new_n932));
  INV_X1    g0732(.A(KEYINPUT43), .ZN(new_n933));
  NOR2_X1   g0733(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n667), .A2(new_n914), .ZN(new_n935));
  NOR2_X1   g0735(.A1(new_n935), .A2(KEYINPUT42), .ZN(new_n936));
  XNOR2_X1  g0736(.A(new_n936), .B(KEYINPUT109), .ZN(new_n937));
  OAI21_X1  g0737(.A(new_n609), .B1(new_n912), .B2(new_n500), .ZN(new_n938));
  OR2_X1    g0738(.A1(new_n938), .A2(KEYINPUT108), .ZN(new_n939));
  AOI21_X1  g0739(.A(new_n668), .B1(new_n938), .B2(KEYINPUT108), .ZN(new_n940));
  AOI22_X1  g0740(.A1(new_n939), .A2(new_n940), .B1(new_n935), .B2(KEYINPUT42), .ZN(new_n941));
  AOI21_X1  g0741(.A(new_n934), .B1(new_n937), .B2(new_n941), .ZN(new_n942));
  NOR3_X1   g0742(.A1(new_n942), .A2(KEYINPUT43), .A3(new_n931), .ZN(new_n943));
  INV_X1    g0743(.A(new_n943), .ZN(new_n944));
  INV_X1    g0744(.A(new_n914), .ZN(new_n945));
  NOR2_X1   g0745(.A1(new_n665), .A2(new_n945), .ZN(new_n946));
  OAI21_X1  g0746(.A(new_n942), .B1(KEYINPUT43), .B2(new_n931), .ZN(new_n947));
  AND3_X1   g0747(.A1(new_n944), .A2(new_n946), .A3(new_n947), .ZN(new_n948));
  AOI21_X1  g0748(.A(new_n946), .B1(new_n944), .B2(new_n947), .ZN(new_n949));
  NOR2_X1   g0749(.A1(new_n948), .A2(new_n949), .ZN(new_n950));
  AND2_X1   g0750(.A1(new_n928), .A2(new_n950), .ZN(new_n951));
  OAI21_X1  g0751(.A(new_n763), .B1(new_n211), .B2(new_n315), .ZN(new_n952));
  NOR2_X1   g0752(.A1(new_n244), .A2(new_n765), .ZN(new_n953));
  OAI21_X1  g0753(.A(new_n708), .B1(new_n952), .B2(new_n953), .ZN(new_n954));
  NOR2_X1   g0754(.A1(new_n732), .A2(new_n311), .ZN(new_n955));
  OAI22_X1  g0755(.A1(new_n743), .A2(new_n751), .B1(new_n728), .B2(new_n202), .ZN(new_n956));
  AOI211_X1 g0756(.A(new_n955), .B(new_n956), .C1(G143), .C2(new_n745), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n754), .A2(G68), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n723), .A2(G137), .ZN(new_n959));
  OAI21_X1  g0759(.A(new_n341), .B1(new_n739), .B2(new_n201), .ZN(new_n960));
  AOI21_X1  g0760(.A(new_n960), .B1(G150), .B2(new_n735), .ZN(new_n961));
  NAND4_X1  g0761(.A1(new_n957), .A2(new_n958), .A3(new_n959), .A4(new_n961), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n729), .A2(G116), .ZN(new_n963));
  XNOR2_X1  g0763(.A(new_n963), .B(KEYINPUT46), .ZN(new_n964));
  OAI21_X1  g0764(.A(new_n279), .B1(new_n739), .B2(new_n731), .ZN(new_n965));
  AOI21_X1  g0765(.A(new_n965), .B1(G303), .B2(new_n735), .ZN(new_n966));
  INV_X1    g0766(.A(G317), .ZN(new_n967));
  OAI211_X1 g0767(.A(new_n964), .B(new_n966), .C1(new_n967), .C2(new_n722), .ZN(new_n968));
  AOI22_X1  g0768(.A1(new_n742), .A2(G294), .B1(new_n745), .B2(G311), .ZN(new_n969));
  INV_X1    g0769(.A(new_n732), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n970), .A2(G97), .ZN(new_n971));
  OAI211_X1 g0771(.A(new_n969), .B(new_n971), .C1(new_n323), .C2(new_n726), .ZN(new_n972));
  OAI21_X1  g0772(.A(new_n962), .B1(new_n968), .B2(new_n972), .ZN(new_n973));
  XNOR2_X1  g0773(.A(new_n973), .B(KEYINPUT47), .ZN(new_n974));
  AOI21_X1  g0774(.A(new_n954), .B1(new_n974), .B2(new_n716), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n932), .A2(new_n714), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n975), .A2(new_n976), .ZN(new_n977));
  INV_X1    g0777(.A(new_n977), .ZN(new_n978));
  NOR2_X1   g0778(.A1(new_n951), .A2(new_n978), .ZN(new_n979));
  INV_X1    g0779(.A(new_n979), .ZN(G387));
  NAND2_X1  g0780(.A1(new_n908), .A2(new_n714), .ZN(new_n981));
  INV_X1    g0781(.A(new_n763), .ZN(new_n982));
  OAI21_X1  g0782(.A(new_n764), .B1(new_n241), .B2(new_n451), .ZN(new_n983));
  OAI21_X1  g0783(.A(new_n983), .B1(new_n675), .B2(new_n769), .ZN(new_n984));
  NOR2_X1   g0784(.A1(new_n317), .A2(G50), .ZN(new_n985));
  XNOR2_X1  g0785(.A(new_n985), .B(KEYINPUT50), .ZN(new_n986));
  AOI21_X1  g0786(.A(G45), .B1(G68), .B2(G77), .ZN(new_n987));
  NAND3_X1  g0787(.A1(new_n986), .A2(new_n675), .A3(new_n987), .ZN(new_n988));
  AOI22_X1  g0788(.A1(new_n984), .A2(new_n988), .B1(new_n207), .B2(new_n672), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n745), .A2(G159), .ZN(new_n990));
  AND2_X1   g0790(.A1(new_n990), .A2(new_n971), .ZN(new_n991));
  OAI221_X1 g0791(.A(new_n991), .B1(new_n311), .B2(new_n728), .C1(new_n266), .C2(new_n743), .ZN(new_n992));
  INV_X1    g0792(.A(new_n754), .ZN(new_n993));
  NOR2_X1   g0793(.A1(new_n993), .A2(new_n315), .ZN(new_n994));
  AOI21_X1  g0794(.A(new_n279), .B1(G50), .B2(new_n735), .ZN(new_n995));
  OAI221_X1 g0795(.A(new_n995), .B1(new_n203), .B2(new_n739), .C1(new_n722), .C2(new_n790), .ZN(new_n996));
  NOR3_X1   g0796(.A1(new_n992), .A2(new_n994), .A3(new_n996), .ZN(new_n997));
  AOI22_X1  g0797(.A1(new_n787), .A2(G303), .B1(G317), .B2(new_n735), .ZN(new_n998));
  XOR2_X1   g0798(.A(KEYINPUT111), .B(G322), .Z(new_n999));
  OAI221_X1 g0799(.A(new_n998), .B1(new_n746), .B2(new_n999), .C1(new_n737), .C2(new_n743), .ZN(new_n1000));
  INV_X1    g0800(.A(KEYINPUT48), .ZN(new_n1001));
  OR2_X1    g0801(.A1(new_n1000), .A2(new_n1001), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n1000), .A2(new_n1001), .ZN(new_n1003));
  AOI22_X1  g0803(.A1(new_n727), .A2(G283), .B1(new_n729), .B2(G294), .ZN(new_n1004));
  NAND3_X1  g0804(.A1(new_n1002), .A2(new_n1003), .A3(new_n1004), .ZN(new_n1005));
  XNOR2_X1  g0805(.A(new_n1005), .B(KEYINPUT112), .ZN(new_n1006));
  OR2_X1    g0806(.A1(new_n1006), .A2(KEYINPUT49), .ZN(new_n1007));
  OAI221_X1 g0807(.A(new_n279), .B1(new_n473), .B2(new_n732), .C1(new_n722), .C2(new_n747), .ZN(new_n1008));
  AOI21_X1  g0808(.A(new_n1008), .B1(new_n1006), .B2(KEYINPUT49), .ZN(new_n1009));
  AOI21_X1  g0809(.A(new_n997), .B1(new_n1007), .B2(new_n1009), .ZN(new_n1010));
  OAI221_X1 g0810(.A(new_n708), .B1(new_n982), .B2(new_n989), .C1(new_n1010), .C2(new_n786), .ZN(new_n1011));
  XNOR2_X1  g0811(.A(new_n1011), .B(KEYINPUT113), .ZN(new_n1012));
  AOI22_X1  g0812(.A1(new_n981), .A2(new_n1012), .B1(new_n910), .B2(new_n707), .ZN(new_n1013));
  NAND2_X1  g0813(.A1(new_n911), .A2(new_n673), .ZN(new_n1014));
  NOR2_X1   g0814(.A1(new_n703), .A2(new_n910), .ZN(new_n1015));
  OAI21_X1  g0815(.A(new_n1013), .B1(new_n1014), .B2(new_n1015), .ZN(G393));
  INV_X1    g0816(.A(KEYINPUT115), .ZN(new_n1017));
  NAND2_X1  g0817(.A1(new_n922), .A2(new_n924), .ZN(new_n1018));
  NAND2_X1  g0818(.A1(new_n1018), .A2(new_n707), .ZN(new_n1019));
  OAI22_X1  g0819(.A1(new_n743), .A2(new_n515), .B1(new_n728), .B2(new_n731), .ZN(new_n1020));
  AOI21_X1  g0820(.A(new_n1020), .B1(G116), .B2(new_n727), .ZN(new_n1021));
  AOI211_X1 g0821(.A(new_n341), .B(new_n758), .C1(G294), .C2(new_n787), .ZN(new_n1022));
  OAI211_X1 g0822(.A(new_n1021), .B(new_n1022), .C1(new_n722), .C2(new_n999), .ZN(new_n1023));
  AOI22_X1  g0823(.A1(new_n745), .A2(G317), .B1(G311), .B2(new_n735), .ZN(new_n1024));
  XNOR2_X1  g0824(.A(new_n1024), .B(KEYINPUT52), .ZN(new_n1025));
  OR2_X1    g0825(.A1(new_n1023), .A2(new_n1025), .ZN(new_n1026));
  AOI22_X1  g0826(.A1(new_n745), .A2(G150), .B1(G159), .B2(new_n735), .ZN(new_n1027));
  XNOR2_X1  g0827(.A(new_n1027), .B(KEYINPUT51), .ZN(new_n1028));
  INV_X1    g0828(.A(new_n1028), .ZN(new_n1029));
  NAND2_X1  g0829(.A1(new_n754), .A2(G77), .ZN(new_n1030));
  NAND2_X1  g0830(.A1(new_n723), .A2(G143), .ZN(new_n1031));
  OAI21_X1  g0831(.A(new_n341), .B1(new_n739), .B2(new_n317), .ZN(new_n1032));
  OAI22_X1  g0832(.A1(new_n743), .A2(new_n201), .B1(new_n728), .B2(new_n203), .ZN(new_n1033));
  AOI211_X1 g0833(.A(new_n1032), .B(new_n1033), .C1(G87), .C2(new_n970), .ZN(new_n1034));
  NAND4_X1  g0834(.A1(new_n1029), .A2(new_n1030), .A3(new_n1031), .A4(new_n1034), .ZN(new_n1035));
  AOI21_X1  g0835(.A(new_n786), .B1(new_n1026), .B2(new_n1035), .ZN(new_n1036));
  NAND2_X1  g0836(.A1(new_n249), .A2(new_n764), .ZN(new_n1037));
  OAI211_X1 g0837(.A(new_n1037), .B(new_n763), .C1(new_n206), .C2(new_n211), .ZN(new_n1038));
  NAND2_X1  g0838(.A1(new_n1038), .A2(new_n708), .ZN(new_n1039));
  XOR2_X1   g0839(.A(new_n1039), .B(KEYINPUT114), .Z(new_n1040));
  AOI211_X1 g0840(.A(new_n1036), .B(new_n1040), .C1(new_n945), .C2(new_n714), .ZN(new_n1041));
  INV_X1    g0841(.A(new_n1041), .ZN(new_n1042));
  AOI21_X1  g0842(.A(new_n1017), .B1(new_n1019), .B2(new_n1042), .ZN(new_n1043));
  INV_X1    g0843(.A(new_n1043), .ZN(new_n1044));
  NAND3_X1  g0844(.A1(new_n1019), .A2(new_n1017), .A3(new_n1042), .ZN(new_n1045));
  NAND3_X1  g0845(.A1(new_n922), .A2(new_n911), .A3(new_n924), .ZN(new_n1046));
  NOR2_X1   g0846(.A1(new_n925), .A2(new_n674), .ZN(new_n1047));
  AOI22_X1  g0847(.A1(new_n1044), .A2(new_n1045), .B1(new_n1046), .B2(new_n1047), .ZN(new_n1048));
  INV_X1    g0848(.A(new_n1048), .ZN(G390));
  NAND2_X1  g0849(.A1(new_n879), .A2(new_n876), .ZN(new_n1050));
  NAND2_X1  g0850(.A1(new_n1050), .A2(new_n712), .ZN(new_n1051));
  OAI22_X1  g0851(.A1(new_n731), .A2(new_n746), .B1(new_n743), .B2(new_n323), .ZN(new_n1052));
  AOI211_X1 g0852(.A(new_n797), .B(new_n1052), .C1(G87), .C2(new_n729), .ZN(new_n1053));
  NAND2_X1  g0853(.A1(new_n723), .A2(G294), .ZN(new_n1054));
  INV_X1    g0854(.A(new_n735), .ZN(new_n1055));
  OAI21_X1  g0855(.A(new_n279), .B1(new_n1055), .B2(new_n473), .ZN(new_n1056));
  AOI21_X1  g0856(.A(new_n1056), .B1(G97), .B2(new_n787), .ZN(new_n1057));
  NAND4_X1  g0857(.A1(new_n1053), .A2(new_n1030), .A3(new_n1054), .A4(new_n1057), .ZN(new_n1058));
  XNOR2_X1  g0858(.A(KEYINPUT54), .B(G143), .ZN(new_n1059));
  INV_X1    g0859(.A(new_n1059), .ZN(new_n1060));
  AOI22_X1  g0860(.A1(new_n742), .A2(G137), .B1(new_n787), .B2(new_n1060), .ZN(new_n1061));
  XOR2_X1   g0861(.A(new_n1061), .B(KEYINPUT117), .Z(new_n1062));
  NAND2_X1  g0862(.A1(new_n723), .A2(G125), .ZN(new_n1063));
  NOR2_X1   g0863(.A1(new_n732), .A2(new_n201), .ZN(new_n1064));
  INV_X1    g0864(.A(G132), .ZN(new_n1065));
  OAI21_X1  g0865(.A(new_n341), .B1(new_n1055), .B2(new_n1065), .ZN(new_n1066));
  AOI211_X1 g0866(.A(new_n1064), .B(new_n1066), .C1(G128), .C2(new_n745), .ZN(new_n1067));
  NOR2_X1   g0867(.A1(new_n728), .A2(new_n790), .ZN(new_n1068));
  XOR2_X1   g0868(.A(KEYINPUT118), .B(KEYINPUT53), .Z(new_n1069));
  XNOR2_X1  g0869(.A(new_n1068), .B(new_n1069), .ZN(new_n1070));
  NAND2_X1  g0870(.A1(new_n754), .A2(G159), .ZN(new_n1071));
  NAND4_X1  g0871(.A1(new_n1063), .A2(new_n1067), .A3(new_n1070), .A4(new_n1071), .ZN(new_n1072));
  OAI21_X1  g0872(.A(new_n1058), .B1(new_n1062), .B2(new_n1072), .ZN(new_n1073));
  NAND2_X1  g0873(.A1(new_n1073), .A2(new_n716), .ZN(new_n1074));
  AOI21_X1  g0874(.A(new_n783), .B1(new_n784), .B2(new_n266), .ZN(new_n1075));
  NAND3_X1  g0875(.A1(new_n1051), .A2(new_n1074), .A3(new_n1075), .ZN(new_n1076));
  OAI21_X1  g0876(.A(new_n1050), .B1(new_n885), .B2(new_n880), .ZN(new_n1077));
  INV_X1    g0877(.A(new_n880), .ZN(new_n1078));
  OAI211_X1 g0878(.A(new_n652), .B(new_n882), .C1(new_n680), .C2(new_n682), .ZN(new_n1079));
  INV_X1    g0879(.A(new_n777), .ZN(new_n1080));
  AND2_X1   g0880(.A1(new_n1079), .A2(new_n1080), .ZN(new_n1081));
  OAI211_X1 g0881(.A(new_n1078), .B(new_n877), .C1(new_n1081), .C2(new_n884), .ZN(new_n1082));
  NAND2_X1  g0882(.A1(new_n1077), .A2(new_n1082), .ZN(new_n1083));
  INV_X1    g0883(.A(G330), .ZN(new_n1084));
  AOI21_X1  g0884(.A(new_n1084), .B1(new_n852), .B2(new_n854), .ZN(new_n1085));
  INV_X1    g0885(.A(new_n884), .ZN(new_n1086));
  NAND3_X1  g0886(.A1(new_n1085), .A2(new_n779), .A3(new_n1086), .ZN(new_n1087));
  INV_X1    g0887(.A(new_n1087), .ZN(new_n1088));
  NAND2_X1  g0888(.A1(new_n1083), .A2(new_n1088), .ZN(new_n1089));
  NAND3_X1  g0889(.A1(new_n701), .A2(new_n658), .A3(new_n779), .ZN(new_n1090));
  OR2_X1    g0890(.A1(new_n1090), .A2(new_n884), .ZN(new_n1091));
  NAND3_X1  g0891(.A1(new_n1077), .A2(new_n1082), .A3(new_n1091), .ZN(new_n1092));
  NAND2_X1  g0892(.A1(new_n1089), .A2(new_n1092), .ZN(new_n1093));
  INV_X1    g0893(.A(new_n1085), .ZN(new_n1094));
  INV_X1    g0894(.A(new_n779), .ZN(new_n1095));
  OAI21_X1  g0895(.A(new_n884), .B1(new_n1094), .B2(new_n1095), .ZN(new_n1096));
  AND3_X1   g0896(.A1(new_n1081), .A2(new_n1096), .A3(new_n1091), .ZN(new_n1097));
  NAND2_X1  g0897(.A1(new_n1090), .A2(new_n884), .ZN(new_n1098));
  AOI21_X1  g0898(.A(new_n883), .B1(new_n1087), .B2(new_n1098), .ZN(new_n1099));
  NOR2_X1   g0899(.A1(new_n1097), .A2(new_n1099), .ZN(new_n1100));
  NAND2_X1  g0900(.A1(new_n437), .A2(new_n1085), .ZN(new_n1101));
  OAI211_X1 g0901(.A(new_n630), .B(new_n1101), .C1(new_n684), .C2(new_n631), .ZN(new_n1102));
  NOR2_X1   g0902(.A1(new_n1100), .A2(new_n1102), .ZN(new_n1103));
  OR2_X1    g0903(.A1(new_n1103), .A2(KEYINPUT116), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n1103), .A2(KEYINPUT116), .ZN(new_n1105));
  AND3_X1   g0905(.A1(new_n1104), .A2(new_n1093), .A3(new_n1105), .ZN(new_n1106));
  NAND3_X1  g0906(.A1(new_n1103), .A2(new_n1092), .A3(new_n1089), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n1107), .A2(new_n673), .ZN(new_n1108));
  OAI221_X1 g0908(.A(new_n1076), .B1(new_n706), .B2(new_n1093), .C1(new_n1106), .C2(new_n1108), .ZN(G378));
  AOI21_X1  g0909(.A(new_n1084), .B1(new_n866), .B2(new_n855), .ZN(new_n1110));
  OAI21_X1  g0910(.A(new_n1110), .B1(new_n858), .B2(new_n859), .ZN(new_n1111));
  NAND2_X1  g0911(.A1(new_n1111), .A2(KEYINPUT121), .ZN(new_n1112));
  INV_X1    g0912(.A(KEYINPUT121), .ZN(new_n1113));
  OAI211_X1 g0913(.A(new_n1110), .B(new_n1113), .C1(new_n858), .C2(new_n859), .ZN(new_n1114));
  NAND2_X1  g0914(.A1(new_n307), .A2(new_n310), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n275), .A2(new_n651), .ZN(new_n1116));
  XNOR2_X1  g0916(.A(new_n1116), .B(KEYINPUT120), .ZN(new_n1117));
  XNOR2_X1  g0917(.A(new_n1115), .B(new_n1117), .ZN(new_n1118));
  XOR2_X1   g0918(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1119));
  XOR2_X1   g0919(.A(new_n1118), .B(new_n1119), .Z(new_n1120));
  INV_X1    g0920(.A(new_n1120), .ZN(new_n1121));
  NAND3_X1  g0921(.A1(new_n1112), .A2(new_n1114), .A3(new_n1121), .ZN(new_n1122));
  INV_X1    g0922(.A(new_n888), .ZN(new_n1123));
  NAND4_X1  g0923(.A1(new_n860), .A2(new_n1113), .A3(new_n1110), .A4(new_n1120), .ZN(new_n1124));
  AND3_X1   g0924(.A1(new_n1122), .A2(new_n1123), .A3(new_n1124), .ZN(new_n1125));
  AOI21_X1  g0925(.A(new_n1123), .B1(new_n1122), .B2(new_n1124), .ZN(new_n1126));
  NOR2_X1   g0926(.A1(new_n1125), .A2(new_n1126), .ZN(new_n1127));
  INV_X1    g0927(.A(KEYINPUT57), .ZN(new_n1128));
  INV_X1    g0928(.A(new_n1102), .ZN(new_n1129));
  AOI21_X1  g0929(.A(new_n1128), .B1(new_n1107), .B2(new_n1129), .ZN(new_n1130));
  AOI21_X1  g0930(.A(new_n674), .B1(new_n1127), .B2(new_n1130), .ZN(new_n1131));
  AND2_X1   g0931(.A1(new_n1107), .A2(new_n1129), .ZN(new_n1132));
  INV_X1    g0932(.A(KEYINPUT122), .ZN(new_n1133));
  OAI21_X1  g0933(.A(new_n1133), .B1(new_n1125), .B2(new_n1126), .ZN(new_n1134));
  NAND2_X1  g0934(.A1(new_n1122), .A2(new_n1124), .ZN(new_n1135));
  NAND2_X1  g0935(.A1(new_n1135), .A2(new_n888), .ZN(new_n1136));
  NAND3_X1  g0936(.A1(new_n1122), .A2(new_n1123), .A3(new_n1124), .ZN(new_n1137));
  NAND3_X1  g0937(.A1(new_n1136), .A2(KEYINPUT122), .A3(new_n1137), .ZN(new_n1138));
  AOI21_X1  g0938(.A(new_n1132), .B1(new_n1134), .B2(new_n1138), .ZN(new_n1139));
  OAI21_X1  g0939(.A(new_n1131), .B1(new_n1139), .B2(KEYINPUT57), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n279), .A2(new_n444), .ZN(new_n1141));
  AOI21_X1  g0941(.A(new_n1141), .B1(new_n729), .B2(G77), .ZN(new_n1142));
  OAI221_X1 g0942(.A(new_n1142), .B1(new_n202), .B2(new_n732), .C1(new_n722), .C2(new_n731), .ZN(new_n1143));
  XOR2_X1   g0943(.A(new_n1143), .B(KEYINPUT119), .Z(new_n1144));
  AOI22_X1  g0944(.A1(new_n787), .A2(new_n601), .B1(G107), .B2(new_n735), .ZN(new_n1145));
  OAI21_X1  g0945(.A(new_n1145), .B1(new_n473), .B2(new_n746), .ZN(new_n1146));
  AOI21_X1  g0946(.A(new_n1146), .B1(G97), .B2(new_n742), .ZN(new_n1147));
  NAND3_X1  g0947(.A1(new_n1144), .A2(new_n958), .A3(new_n1147), .ZN(new_n1148));
  INV_X1    g0948(.A(KEYINPUT58), .ZN(new_n1149));
  OR2_X1    g0949(.A1(new_n1148), .A2(new_n1149), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n1148), .A2(new_n1149), .ZN(new_n1151));
  OAI211_X1 g0951(.A(new_n1141), .B(new_n201), .C1(G33), .C2(G41), .ZN(new_n1152));
  INV_X1    g0952(.A(G128), .ZN(new_n1153));
  OAI22_X1  g0953(.A1(new_n1055), .A2(new_n1153), .B1(new_n739), .B2(new_n789), .ZN(new_n1154));
  AOI21_X1  g0954(.A(new_n1154), .B1(G132), .B2(new_n742), .ZN(new_n1155));
  AOI22_X1  g0955(.A1(new_n745), .A2(G125), .B1(new_n729), .B2(new_n1060), .ZN(new_n1156));
  OAI211_X1 g0956(.A(new_n1155), .B(new_n1156), .C1(new_n993), .C2(new_n790), .ZN(new_n1157));
  OR2_X1    g0957(.A1(new_n1157), .A2(KEYINPUT59), .ZN(new_n1158));
  NAND2_X1  g0958(.A1(new_n1157), .A2(KEYINPUT59), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n723), .A2(G124), .ZN(new_n1160));
  AOI211_X1 g0960(.A(G33), .B(G41), .C1(new_n970), .C2(G159), .ZN(new_n1161));
  NAND4_X1  g0961(.A1(new_n1158), .A2(new_n1159), .A3(new_n1160), .A4(new_n1161), .ZN(new_n1162));
  NAND4_X1  g0962(.A1(new_n1150), .A2(new_n1151), .A3(new_n1152), .A4(new_n1162), .ZN(new_n1163));
  NAND2_X1  g0963(.A1(new_n1163), .A2(new_n716), .ZN(new_n1164));
  AOI21_X1  g0964(.A(new_n783), .B1(new_n784), .B2(new_n201), .ZN(new_n1165));
  OAI211_X1 g0965(.A(new_n1164), .B(new_n1165), .C1(new_n1121), .C2(new_n713), .ZN(new_n1166));
  INV_X1    g0966(.A(new_n1166), .ZN(new_n1167));
  NAND2_X1  g0967(.A1(new_n1134), .A2(new_n1138), .ZN(new_n1168));
  AOI21_X1  g0968(.A(new_n1167), .B1(new_n1168), .B2(new_n707), .ZN(new_n1169));
  NAND2_X1  g0969(.A1(new_n1140), .A2(new_n1169), .ZN(G375));
  NAND2_X1  g0970(.A1(new_n1100), .A2(new_n1102), .ZN(new_n1171));
  NAND4_X1  g0971(.A1(new_n1104), .A2(new_n907), .A3(new_n1105), .A4(new_n1171), .ZN(new_n1172));
  AOI21_X1  g0972(.A(new_n783), .B1(new_n784), .B2(new_n203), .ZN(new_n1173));
  OAI22_X1  g0973(.A1(new_n722), .A2(new_n1153), .B1(new_n751), .B2(new_n728), .ZN(new_n1174));
  XOR2_X1   g0974(.A(new_n1174), .B(KEYINPUT123), .Z(new_n1175));
  NOR2_X1   g0975(.A1(new_n993), .A2(new_n201), .ZN(new_n1176));
  OAI221_X1 g0976(.A(new_n341), .B1(new_n739), .B2(new_n790), .C1(new_n1055), .C2(new_n789), .ZN(new_n1177));
  NOR2_X1   g0977(.A1(new_n743), .A2(new_n1059), .ZN(new_n1178));
  OAI22_X1  g0978(.A1(new_n746), .A2(new_n1065), .B1(new_n732), .B2(new_n202), .ZN(new_n1179));
  NOR4_X1   g0979(.A1(new_n1176), .A2(new_n1177), .A3(new_n1178), .A4(new_n1179), .ZN(new_n1180));
  INV_X1    g0980(.A(new_n994), .ZN(new_n1181));
  NOR2_X1   g0981(.A1(new_n722), .A2(new_n515), .ZN(new_n1182));
  OAI221_X1 g0982(.A(new_n279), .B1(new_n739), .B2(new_n323), .C1(new_n1055), .C2(new_n731), .ZN(new_n1183));
  OAI22_X1  g0983(.A1(new_n743), .A2(new_n473), .B1(new_n732), .B2(new_n311), .ZN(new_n1184));
  OAI22_X1  g0984(.A1(new_n746), .A2(new_n440), .B1(new_n728), .B2(new_n206), .ZN(new_n1185));
  NOR4_X1   g0985(.A1(new_n1182), .A2(new_n1183), .A3(new_n1184), .A4(new_n1185), .ZN(new_n1186));
  AOI22_X1  g0986(.A1(new_n1175), .A2(new_n1180), .B1(new_n1181), .B2(new_n1186), .ZN(new_n1187));
  OAI221_X1 g0987(.A(new_n1173), .B1(new_n786), .B2(new_n1187), .C1(new_n1086), .C2(new_n713), .ZN(new_n1188));
  OAI21_X1  g0988(.A(new_n1188), .B1(new_n1100), .B2(new_n706), .ZN(new_n1189));
  INV_X1    g0989(.A(new_n1189), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n1172), .A2(new_n1190), .ZN(G381));
  NOR3_X1   g0991(.A1(G393), .A2(G396), .A3(G384), .ZN(new_n1192));
  NAND3_X1  g0992(.A1(new_n979), .A2(new_n1048), .A3(new_n1192), .ZN(new_n1193));
  OR4_X1    g0993(.A1(G378), .A2(G375), .A3(G381), .A4(new_n1193), .ZN(G407));
  NOR2_X1   g0994(.A1(new_n1106), .A2(new_n1108), .ZN(new_n1195));
  OAI21_X1  g0995(.A(new_n1076), .B1(new_n1093), .B2(new_n706), .ZN(new_n1196));
  NOR2_X1   g0996(.A1(new_n1195), .A2(new_n1196), .ZN(new_n1197));
  NOR2_X1   g0997(.A1(new_n649), .A2(G343), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(new_n1197), .A2(new_n1198), .ZN(new_n1199));
  OAI211_X1 g0999(.A(G407), .B(G213), .C1(G375), .C2(new_n1199), .ZN(G409));
  OAI21_X1  g1000(.A(KEYINPUT125), .B1(new_n951), .B2(new_n978), .ZN(new_n1201));
  INV_X1    g1001(.A(new_n1201), .ZN(new_n1202));
  NOR3_X1   g1002(.A1(new_n951), .A2(KEYINPUT125), .A3(new_n978), .ZN(new_n1203));
  XNOR2_X1  g1003(.A(G393), .B(new_n774), .ZN(new_n1204));
  INV_X1    g1004(.A(new_n1204), .ZN(new_n1205));
  NAND2_X1  g1005(.A1(new_n1048), .A2(new_n1205), .ZN(new_n1206));
  INV_X1    g1006(.A(new_n1206), .ZN(new_n1207));
  NOR2_X1   g1007(.A1(new_n1048), .A2(new_n1205), .ZN(new_n1208));
  OAI22_X1  g1008(.A1(new_n1202), .A2(new_n1203), .B1(new_n1207), .B2(new_n1208), .ZN(new_n1209));
  INV_X1    g1009(.A(new_n1203), .ZN(new_n1210));
  INV_X1    g1010(.A(new_n1208), .ZN(new_n1211));
  NAND4_X1  g1011(.A1(new_n1210), .A2(new_n1211), .A3(new_n1201), .A4(new_n1206), .ZN(new_n1212));
  NAND2_X1  g1012(.A1(new_n1209), .A2(new_n1212), .ZN(new_n1213));
  INV_X1    g1013(.A(new_n1132), .ZN(new_n1214));
  AOI21_X1  g1014(.A(KEYINPUT57), .B1(new_n1168), .B2(new_n1214), .ZN(new_n1215));
  INV_X1    g1015(.A(new_n1131), .ZN(new_n1216));
  OAI211_X1 g1016(.A(G378), .B(new_n1169), .C1(new_n1215), .C2(new_n1216), .ZN(new_n1217));
  AOI211_X1 g1017(.A(new_n906), .B(new_n1132), .C1(new_n1134), .C2(new_n1138), .ZN(new_n1218));
  INV_X1    g1018(.A(new_n1127), .ZN(new_n1219));
  OAI21_X1  g1019(.A(new_n1166), .B1(new_n1219), .B2(new_n706), .ZN(new_n1220));
  OAI21_X1  g1020(.A(new_n1197), .B1(new_n1218), .B2(new_n1220), .ZN(new_n1221));
  AOI21_X1  g1021(.A(new_n1198), .B1(new_n1217), .B2(new_n1221), .ZN(new_n1222));
  OAI21_X1  g1022(.A(KEYINPUT60), .B1(new_n1100), .B2(new_n1102), .ZN(new_n1223));
  NAND2_X1  g1023(.A1(new_n1223), .A2(new_n1171), .ZN(new_n1224));
  NAND3_X1  g1024(.A1(new_n1100), .A2(KEYINPUT60), .A3(new_n1102), .ZN(new_n1225));
  NAND3_X1  g1025(.A1(new_n1224), .A2(new_n673), .A3(new_n1225), .ZN(new_n1226));
  NAND3_X1  g1026(.A1(new_n1226), .A2(G384), .A3(new_n1190), .ZN(new_n1227));
  INV_X1    g1027(.A(new_n1227), .ZN(new_n1228));
  AOI21_X1  g1028(.A(G384), .B1(new_n1226), .B2(new_n1190), .ZN(new_n1229));
  NOR2_X1   g1029(.A1(new_n1228), .A2(new_n1229), .ZN(new_n1230));
  NAND2_X1  g1030(.A1(new_n1222), .A2(new_n1230), .ZN(new_n1231));
  INV_X1    g1031(.A(KEYINPUT63), .ZN(new_n1232));
  AOI21_X1  g1032(.A(new_n1213), .B1(new_n1231), .B2(new_n1232), .ZN(new_n1233));
  NAND3_X1  g1033(.A1(new_n1222), .A2(KEYINPUT63), .A3(new_n1230), .ZN(new_n1234));
  INV_X1    g1034(.A(KEYINPUT61), .ZN(new_n1235));
  INV_X1    g1035(.A(KEYINPUT124), .ZN(new_n1236));
  OAI21_X1  g1036(.A(new_n1236), .B1(new_n1228), .B2(new_n1229), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(new_n1198), .A2(G2897), .ZN(new_n1238));
  OR2_X1    g1038(.A1(new_n1237), .A2(new_n1238), .ZN(new_n1239));
  NOR3_X1   g1039(.A1(new_n1228), .A2(new_n1236), .A3(new_n1229), .ZN(new_n1240));
  OAI21_X1  g1040(.A(new_n1237), .B1(new_n1240), .B2(new_n1238), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(new_n1239), .A2(new_n1241), .ZN(new_n1242));
  OAI21_X1  g1042(.A(new_n1235), .B1(new_n1222), .B2(new_n1242), .ZN(new_n1243));
  INV_X1    g1043(.A(new_n1243), .ZN(new_n1244));
  NAND3_X1  g1044(.A1(new_n1233), .A2(new_n1234), .A3(new_n1244), .ZN(new_n1245));
  INV_X1    g1045(.A(KEYINPUT62), .ZN(new_n1246));
  AND3_X1   g1046(.A1(new_n1222), .A2(new_n1246), .A3(new_n1230), .ZN(new_n1247));
  AOI21_X1  g1047(.A(new_n1246), .B1(new_n1222), .B2(new_n1230), .ZN(new_n1248));
  NOR3_X1   g1048(.A1(new_n1247), .A2(new_n1243), .A3(new_n1248), .ZN(new_n1249));
  INV_X1    g1049(.A(new_n1213), .ZN(new_n1250));
  OAI21_X1  g1050(.A(new_n1245), .B1(new_n1249), .B2(new_n1250), .ZN(G405));
  AOI21_X1  g1051(.A(G378), .B1(new_n1140), .B2(new_n1169), .ZN(new_n1252));
  INV_X1    g1052(.A(new_n1252), .ZN(new_n1253));
  OR3_X1    g1053(.A1(new_n1228), .A2(new_n1229), .A3(KEYINPUT126), .ZN(new_n1254));
  NAND3_X1  g1054(.A1(new_n1253), .A2(new_n1217), .A3(new_n1254), .ZN(new_n1255));
  OAI21_X1  g1055(.A(KEYINPUT126), .B1(new_n1228), .B2(new_n1229), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(new_n1254), .A2(new_n1256), .ZN(new_n1257));
  INV_X1    g1057(.A(new_n1217), .ZN(new_n1258));
  OAI21_X1  g1058(.A(new_n1257), .B1(new_n1258), .B2(new_n1252), .ZN(new_n1259));
  NAND3_X1  g1059(.A1(new_n1255), .A2(new_n1259), .A3(new_n1213), .ZN(new_n1260));
  AOI21_X1  g1060(.A(new_n1213), .B1(new_n1255), .B2(new_n1259), .ZN(new_n1261));
  INV_X1    g1061(.A(KEYINPUT127), .ZN(new_n1262));
  OAI21_X1  g1062(.A(new_n1260), .B1(new_n1261), .B2(new_n1262), .ZN(new_n1263));
  AOI211_X1 g1063(.A(KEYINPUT127), .B(new_n1213), .C1(new_n1255), .C2(new_n1259), .ZN(new_n1264));
  NOR2_X1   g1064(.A1(new_n1263), .A2(new_n1264), .ZN(G402));
endmodule


