

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359,
         n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370,
         n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381,
         n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392,
         n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403,
         n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414,
         n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425,
         n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436,
         n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447,
         n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458,
         n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469,
         n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480,
         n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491,
         n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502,
         n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513,
         n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601,
         n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612,
         n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623,
         n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634,
         n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645,
         n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656,
         n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667,
         n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678,
         n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689,
         n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700,
         n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711,
         n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722,
         n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733,
         n734, n735, n736, n737, n738, n739, n740, n741, n742, n743;

  NOR2_X1 U373 ( .A1(n661), .A2(n579), .ZN(n594) );
  INV_X4 U374 ( .A(G953), .ZN(n457) );
  XNOR2_X2 U375 ( .A(n483), .B(KEYINPUT33), .ZN(n693) );
  XNOR2_X2 U376 ( .A(n421), .B(G143), .ZN(n485) );
  AND2_X1 U377 ( .A1(n375), .A2(n372), .ZN(n371) );
  AND2_X1 U378 ( .A1(n409), .A2(n408), .ZN(n555) );
  AND2_X1 U379 ( .A1(n360), .A2(n366), .ZN(n357) );
  NAND2_X1 U380 ( .A1(n614), .A2(n664), .ZN(n565) );
  XOR2_X1 U381 ( .A(G146), .B(KEYINPUT4), .Z(n484) );
  XNOR2_X2 U382 ( .A(n565), .B(KEYINPUT19), .ZN(n576) );
  XNOR2_X1 U383 ( .A(n444), .B(n530), .ZN(n727) );
  XNOR2_X2 U384 ( .A(n412), .B(n351), .ZN(n614) );
  INV_X1 U385 ( .A(G134), .ZN(n443) );
  NAND2_X1 U386 ( .A1(n399), .A2(n398), .ZN(n397) );
  NAND2_X1 U387 ( .A1(n706), .A2(G469), .ZN(n399) );
  INV_X1 U388 ( .A(n714), .ZN(n413) );
  NOR2_X1 U389 ( .A1(n706), .A2(n395), .ZN(n394) );
  NAND2_X1 U390 ( .A1(n453), .A2(n396), .ZN(n395) );
  INV_X1 U391 ( .A(G469), .ZN(n396) );
  XNOR2_X1 U392 ( .A(n442), .B(n441), .ZN(n444) );
  INV_X1 U393 ( .A(KEYINPUT78), .ZN(n404) );
  NAND2_X1 U394 ( .A1(n362), .A2(n361), .ZN(n360) );
  NOR2_X1 U395 ( .A1(n657), .A2(KEYINPUT99), .ZN(n361) );
  INV_X1 U396 ( .A(n669), .ZN(n367) );
  NAND2_X1 U397 ( .A1(n644), .A2(KEYINPUT99), .ZN(n366) );
  INV_X1 U398 ( .A(KEYINPUT104), .ZN(n364) );
  XNOR2_X1 U399 ( .A(KEYINPUT20), .B(KEYINPUT94), .ZN(n464) );
  NOR2_X1 U400 ( .A1(G953), .A2(G237), .ZN(n513) );
  XOR2_X1 U401 ( .A(KEYINPUT95), .B(KEYINPUT25), .Z(n467) );
  XNOR2_X1 U402 ( .A(G113), .B(KEYINPUT97), .ZN(n476) );
  XOR2_X1 U403 ( .A(KEYINPUT5), .B(KEYINPUT71), .Z(n477) );
  NOR2_X1 U404 ( .A1(n606), .A2(n607), .ZN(n417) );
  XNOR2_X1 U405 ( .A(n475), .B(n426), .ZN(n492) );
  XNOR2_X1 U406 ( .A(n427), .B(G119), .ZN(n426) );
  INV_X1 U407 ( .A(G101), .ZN(n427) );
  AND2_X1 U408 ( .A1(n729), .A2(n620), .ZN(n401) );
  OR2_X1 U409 ( .A1(G902), .A2(G237), .ZN(n495) );
  NOR2_X1 U410 ( .A1(n394), .A2(KEYINPUT1), .ZN(n389) );
  XNOR2_X1 U411 ( .A(n525), .B(n524), .ZN(n552) );
  XNOR2_X1 U412 ( .A(n523), .B(G475), .ZN(n524) );
  XNOR2_X1 U413 ( .A(n432), .B(n431), .ZN(n674) );
  INV_X1 U414 ( .A(KEYINPUT67), .ZN(n431) );
  NOR2_X1 U415 ( .A1(n678), .A2(n677), .ZN(n432) );
  OR2_X1 U416 ( .A1(G902), .A2(n635), .ZN(n481) );
  XOR2_X1 U417 ( .A(G122), .B(G107), .Z(n526) );
  XNOR2_X1 U418 ( .A(n528), .B(n381), .ZN(n380) );
  INV_X1 U419 ( .A(KEYINPUT9), .ZN(n381) );
  XNOR2_X1 U420 ( .A(n597), .B(KEYINPUT39), .ZN(n616) );
  AND2_X1 U421 ( .A1(n553), .A2(n554), .ZN(n598) );
  XNOR2_X1 U422 ( .A(n727), .B(n452), .ZN(n706) );
  XNOR2_X1 U423 ( .A(n449), .B(n448), .ZN(n450) );
  NOR2_X1 U424 ( .A1(G952), .A2(n457), .ZN(n713) );
  XNOR2_X1 U425 ( .A(n437), .B(n704), .ZN(n436) );
  AND2_X1 U426 ( .A1(n373), .A2(n457), .ZN(n372) );
  NAND2_X1 U427 ( .A1(n374), .A2(KEYINPUT118), .ZN(n373) );
  NAND2_X1 U428 ( .A1(G234), .A2(G237), .ZN(n496) );
  XOR2_X1 U429 ( .A(KEYINPUT89), .B(KEYINPUT14), .Z(n497) );
  NAND2_X1 U430 ( .A1(n349), .A2(n353), .ZN(n363) );
  XOR2_X1 U431 ( .A(KEYINPUT17), .B(KEYINPUT74), .Z(n489) );
  INV_X1 U432 ( .A(KEYINPUT84), .ZN(n420) );
  XNOR2_X1 U433 ( .A(G113), .B(G104), .ZN(n518) );
  XOR2_X1 U434 ( .A(KEYINPUT68), .B(G131), .Z(n512) );
  NOR2_X1 U435 ( .A1(n572), .A2(n564), .ZN(n609) );
  AND2_X1 U436 ( .A1(n550), .A2(n539), .ZN(n483) );
  NOR2_X1 U437 ( .A1(n402), .A2(n582), .ZN(n584) );
  INV_X1 U438 ( .A(KEYINPUT72), .ZN(n583) );
  XNOR2_X1 U439 ( .A(n470), .B(n469), .ZN(n678) );
  XNOR2_X1 U440 ( .A(n727), .B(n382), .ZN(n635) );
  XNOR2_X1 U441 ( .A(n480), .B(n383), .ZN(n382) );
  INV_X1 U442 ( .A(n492), .ZN(n383) );
  INV_X1 U443 ( .A(n663), .ZN(n617) );
  XNOR2_X1 U444 ( .A(n428), .B(n492), .ZN(n714) );
  XNOR2_X1 U445 ( .A(n494), .B(n526), .ZN(n428) );
  XNOR2_X1 U446 ( .A(n493), .B(n518), .ZN(n494) );
  XOR2_X1 U447 ( .A(G110), .B(KEYINPUT16), .Z(n493) );
  XNOR2_X1 U448 ( .A(G104), .B(G107), .ZN(n447) );
  XNOR2_X1 U449 ( .A(n446), .B(n445), .ZN(n449) );
  INV_X1 U450 ( .A(KEYINPUT92), .ZN(n445) );
  INV_X1 U451 ( .A(n700), .ZN(n374) );
  NAND2_X2 U452 ( .A1(n391), .A2(n388), .ZN(n542) );
  AND2_X1 U453 ( .A1(n393), .A2(n392), .ZN(n391) );
  NAND2_X1 U454 ( .A1(n390), .A2(n389), .ZN(n388) );
  NAND2_X1 U455 ( .A1(n674), .A2(n574), .ZN(n402) );
  BUF_X1 U456 ( .A(n678), .Z(n379) );
  NAND2_X1 U457 ( .A1(n422), .A2(G472), .ZN(n637) );
  XNOR2_X1 U458 ( .A(n380), .B(n529), .ZN(n532) );
  XNOR2_X1 U459 ( .A(n407), .B(n406), .ZN(n737) );
  XNOR2_X1 U460 ( .A(n599), .B(KEYINPUT109), .ZN(n406) );
  NAND2_X1 U461 ( .A1(n616), .A2(n598), .ZN(n407) );
  XNOR2_X1 U462 ( .A(n423), .B(n438), .ZN(n739) );
  XNOR2_X1 U463 ( .A(n439), .B(KEYINPUT35), .ZN(n438) );
  INV_X1 U464 ( .A(KEYINPUT83), .ZN(n439) );
  XNOR2_X1 U465 ( .A(n385), .B(n551), .ZN(n657) );
  XNOR2_X1 U466 ( .A(n430), .B(n429), .ZN(n707) );
  XNOR2_X1 U467 ( .A(n706), .B(n705), .ZN(n429) );
  INV_X1 U468 ( .A(KEYINPUT56), .ZN(n433) );
  NAND2_X1 U469 ( .A1(n436), .A2(n435), .ZN(n434) );
  INV_X1 U470 ( .A(n713), .ZN(n435) );
  INV_X1 U471 ( .A(KEYINPUT53), .ZN(n410) );
  NAND2_X1 U472 ( .A1(n370), .A2(KEYINPUT118), .ZN(n369) );
  AND2_X1 U473 ( .A1(n358), .A2(n360), .ZN(n349) );
  AND2_X1 U474 ( .A1(n729), .A2(KEYINPUT2), .ZN(n350) );
  AND2_X1 U475 ( .A1(n495), .A2(G210), .ZN(n351) );
  OR2_X1 U476 ( .A1(n557), .A2(KEYINPUT44), .ZN(n352) );
  INV_X1 U477 ( .A(G902), .ZN(n453) );
  AND2_X1 U478 ( .A1(n366), .A2(n364), .ZN(n353) );
  XNOR2_X1 U479 ( .A(KEYINPUT79), .B(KEYINPUT2), .ZN(n354) );
  NOR2_X1 U480 ( .A1(n355), .A2(n402), .ZN(n425) );
  NOR2_X1 U481 ( .A1(n355), .A2(n667), .ZN(n535) );
  NOR2_X1 U482 ( .A1(n355), .A2(n683), .ZN(n385) );
  NOR2_X1 U483 ( .A1(n693), .A2(n355), .ZN(n506) );
  XNOR2_X2 U484 ( .A(n505), .B(KEYINPUT0), .ZN(n355) );
  NAND2_X1 U485 ( .A1(n356), .A2(KEYINPUT104), .ZN(n365) );
  NAND2_X1 U486 ( .A1(n357), .A2(n358), .ZN(n356) );
  AND2_X1 U487 ( .A1(n359), .A2(n367), .ZN(n358) );
  NAND2_X1 U488 ( .A1(n657), .A2(KEYINPUT99), .ZN(n359) );
  INV_X1 U489 ( .A(n644), .ZN(n362) );
  NAND2_X1 U490 ( .A1(n365), .A2(n363), .ZN(n409) );
  NAND2_X1 U491 ( .A1(n721), .A2(n729), .ZN(n368) );
  NAND2_X1 U492 ( .A1(n721), .A2(n350), .ZN(n697) );
  AND2_X1 U493 ( .A1(n368), .A2(n354), .ZN(n405) );
  NAND2_X1 U494 ( .A1(n371), .A2(n369), .ZN(n377) );
  INV_X1 U495 ( .A(n699), .ZN(n370) );
  NAND2_X1 U496 ( .A1(n699), .A2(n376), .ZN(n375) );
  AND2_X1 U497 ( .A1(n700), .A2(n411), .ZN(n376) );
  XNOR2_X1 U498 ( .A(n377), .B(n410), .ZN(G75) );
  XNOR2_X1 U499 ( .A(n378), .B(n455), .ZN(n461) );
  XNOR2_X1 U500 ( .A(n456), .B(n454), .ZN(n378) );
  NAND2_X2 U501 ( .A1(n400), .A2(n622), .ZN(n633) );
  NOR2_X1 U502 ( .A1(n739), .A2(n648), .ZN(n547) );
  XNOR2_X1 U503 ( .A(n384), .B(n420), .ZN(n419) );
  NAND2_X1 U504 ( .A1(n555), .A2(n556), .ZN(n384) );
  XNOR2_X1 U505 ( .A(n486), .B(n487), .ZN(n491) );
  AND2_X2 U506 ( .A1(n386), .A2(n571), .ZN(n644) );
  XNOR2_X1 U507 ( .A(n425), .B(KEYINPUT96), .ZN(n386) );
  NAND2_X1 U508 ( .A1(n390), .A2(n387), .ZN(n574) );
  INV_X1 U509 ( .A(n394), .ZN(n387) );
  NAND2_X1 U510 ( .A1(n674), .A2(n542), .ZN(n474) );
  INV_X1 U511 ( .A(n397), .ZN(n390) );
  NAND2_X1 U512 ( .A1(n394), .A2(KEYINPUT1), .ZN(n392) );
  NAND2_X1 U513 ( .A1(n397), .A2(KEYINPUT1), .ZN(n393) );
  NAND2_X1 U514 ( .A1(G902), .A2(G469), .ZN(n398) );
  AND2_X4 U515 ( .A1(n697), .A2(n633), .ZN(n422) );
  NAND2_X1 U516 ( .A1(n401), .A2(n721), .ZN(n400) );
  NOR2_X1 U517 ( .A1(n403), .A2(G902), .ZN(n470) );
  XNOR2_X1 U518 ( .A(n711), .B(n403), .ZN(n712) );
  XNOR2_X1 U519 ( .A(n463), .B(n507), .ZN(n403) );
  XNOR2_X1 U520 ( .A(n405), .B(n404), .ZN(n698) );
  INV_X1 U521 ( .A(n641), .ZN(n408) );
  INV_X1 U522 ( .A(KEYINPUT118), .ZN(n411) );
  NAND2_X1 U523 ( .A1(n701), .A2(n619), .ZN(n412) );
  XNOR2_X1 U524 ( .A(n414), .B(n413), .ZN(n701) );
  XNOR2_X1 U525 ( .A(n491), .B(n415), .ZN(n414) );
  XNOR2_X1 U526 ( .A(n490), .B(KEYINPUT88), .ZN(n415) );
  XNOR2_X1 U527 ( .A(n417), .B(KEYINPUT48), .ZN(n416) );
  AND2_X2 U528 ( .A1(n416), .A2(n618), .ZN(n729) );
  XNOR2_X1 U529 ( .A(n584), .B(n583), .ZN(n585) );
  NAND2_X1 U530 ( .A1(n419), .A2(n352), .ZN(n418) );
  XNOR2_X2 U531 ( .A(n418), .B(KEYINPUT45), .ZN(n721) );
  XNOR2_X2 U532 ( .A(G128), .B(KEYINPUT76), .ZN(n421) );
  NAND2_X1 U533 ( .A1(n422), .A2(G210), .ZN(n437) );
  NAND2_X1 U534 ( .A1(n422), .A2(G478), .ZN(n708) );
  NAND2_X1 U535 ( .A1(n422), .A2(G217), .ZN(n711) );
  NAND2_X1 U536 ( .A1(n422), .A2(G469), .ZN(n430) );
  NAND2_X1 U537 ( .A1(n424), .A2(n587), .ZN(n423) );
  XNOR2_X1 U538 ( .A(n506), .B(KEYINPUT34), .ZN(n424) );
  INV_X1 U539 ( .A(n614), .ZN(n595) );
  XNOR2_X1 U540 ( .A(n434), .B(n433), .ZN(G51) );
  XNOR2_X1 U541 ( .A(n474), .B(n473), .ZN(n550) );
  XOR2_X1 U542 ( .A(G140), .B(G110), .Z(n440) );
  INV_X1 U543 ( .A(KEYINPUT12), .ZN(n514) );
  XNOR2_X1 U544 ( .A(n515), .B(n514), .ZN(n516) );
  XNOR2_X1 U545 ( .A(n479), .B(n478), .ZN(n480) );
  XNOR2_X1 U546 ( .A(n517), .B(n516), .ZN(n520) );
  INV_X1 U547 ( .A(KEYINPUT70), .ZN(n473) );
  NOR2_X1 U548 ( .A1(n738), .A2(n617), .ZN(n618) );
  XNOR2_X1 U549 ( .A(n567), .B(KEYINPUT112), .ZN(n568) );
  XNOR2_X1 U550 ( .A(n635), .B(n634), .ZN(n636) );
  XNOR2_X1 U551 ( .A(n627), .B(n626), .ZN(n628) );
  XNOR2_X1 U552 ( .A(n569), .B(n568), .ZN(n570) );
  XNOR2_X1 U553 ( .A(n637), .B(n636), .ZN(n638) );
  XNOR2_X1 U554 ( .A(n629), .B(n628), .ZN(n630) );
  XNOR2_X1 U555 ( .A(KEYINPUT60), .B(KEYINPUT66), .ZN(n631) );
  XNOR2_X1 U556 ( .A(n632), .B(n631), .ZN(G60) );
  XNOR2_X1 U557 ( .A(n484), .B(G137), .ZN(n442) );
  INV_X1 U558 ( .A(n512), .ZN(n441) );
  XNOR2_X1 U559 ( .A(n443), .B(n485), .ZN(n530) );
  XNOR2_X1 U560 ( .A(G101), .B(KEYINPUT73), .ZN(n451) );
  NAND2_X1 U561 ( .A1(G227), .A2(n457), .ZN(n446) );
  XNOR2_X1 U562 ( .A(n440), .B(n447), .ZN(n448) );
  XNOR2_X1 U563 ( .A(n451), .B(n450), .ZN(n452) );
  XOR2_X1 U564 ( .A(G137), .B(G110), .Z(n455) );
  XNOR2_X1 U565 ( .A(G128), .B(G119), .ZN(n454) );
  XOR2_X1 U566 ( .A(KEYINPUT24), .B(KEYINPUT23), .Z(n456) );
  NAND2_X1 U567 ( .A1(n457), .A2(G234), .ZN(n459) );
  XNOR2_X1 U568 ( .A(KEYINPUT81), .B(KEYINPUT8), .ZN(n458) );
  XNOR2_X1 U569 ( .A(n459), .B(n458), .ZN(n527) );
  NAND2_X1 U570 ( .A1(G221), .A2(n527), .ZN(n460) );
  XNOR2_X1 U571 ( .A(n461), .B(n460), .ZN(n463) );
  XNOR2_X1 U572 ( .A(G125), .B(G140), .ZN(n462) );
  XNOR2_X1 U573 ( .A(n462), .B(KEYINPUT10), .ZN(n726) );
  XNOR2_X1 U574 ( .A(G146), .B(n726), .ZN(n507) );
  XNOR2_X1 U575 ( .A(G902), .B(KEYINPUT15), .ZN(n619) );
  NAND2_X1 U576 ( .A1(n619), .A2(G234), .ZN(n465) );
  XNOR2_X1 U577 ( .A(n465), .B(n464), .ZN(n471) );
  NAND2_X1 U578 ( .A1(G217), .A2(n471), .ZN(n466) );
  XNOR2_X1 U579 ( .A(n467), .B(n466), .ZN(n468) );
  XNOR2_X1 U580 ( .A(KEYINPUT93), .B(n468), .ZN(n469) );
  NAND2_X1 U581 ( .A1(n471), .A2(G221), .ZN(n472) );
  XNOR2_X1 U582 ( .A(n472), .B(KEYINPUT21), .ZN(n677) );
  XNOR2_X1 U583 ( .A(G116), .B(KEYINPUT3), .ZN(n475) );
  XNOR2_X1 U584 ( .A(n477), .B(n476), .ZN(n479) );
  AND2_X1 U585 ( .A1(n513), .A2(G210), .ZN(n478) );
  XNOR2_X2 U586 ( .A(G472), .B(n481), .ZN(n580) );
  INV_X1 U587 ( .A(KEYINPUT6), .ZN(n482) );
  XNOR2_X1 U588 ( .A(n580), .B(n482), .ZN(n539) );
  XOR2_X1 U589 ( .A(n484), .B(KEYINPUT18), .Z(n487) );
  XNOR2_X1 U590 ( .A(n485), .B(G125), .ZN(n486) );
  NAND2_X1 U591 ( .A1(G224), .A2(n457), .ZN(n488) );
  XNOR2_X1 U592 ( .A(n489), .B(n488), .ZN(n490) );
  NAND2_X1 U593 ( .A1(G214), .A2(n495), .ZN(n664) );
  XNOR2_X1 U594 ( .A(n497), .B(n496), .ZN(n498) );
  XOR2_X1 U595 ( .A(KEYINPUT69), .B(n498), .Z(n500) );
  NAND2_X1 U596 ( .A1(n500), .A2(G952), .ZN(n692) );
  NOR2_X1 U597 ( .A1(G953), .A2(n692), .ZN(n499) );
  XOR2_X1 U598 ( .A(KEYINPUT90), .B(n499), .Z(n560) );
  NAND2_X1 U599 ( .A1(n500), .A2(G902), .ZN(n501) );
  XOR2_X1 U600 ( .A(KEYINPUT91), .B(n501), .Z(n558) );
  INV_X1 U601 ( .A(n558), .ZN(n502) );
  NOR2_X1 U602 ( .A1(G898), .A2(n457), .ZN(n716) );
  NAND2_X1 U603 ( .A1(n502), .A2(n716), .ZN(n503) );
  NAND2_X1 U604 ( .A1(n560), .A2(n503), .ZN(n504) );
  NAND2_X1 U605 ( .A1(n576), .A2(n504), .ZN(n505) );
  INV_X1 U606 ( .A(n507), .ZN(n511) );
  XOR2_X1 U607 ( .A(KEYINPUT102), .B(KEYINPUT11), .Z(n509) );
  XNOR2_X1 U608 ( .A(G122), .B(KEYINPUT101), .ZN(n508) );
  XNOR2_X1 U609 ( .A(n509), .B(n508), .ZN(n510) );
  XNOR2_X1 U610 ( .A(n511), .B(n510), .ZN(n522) );
  XOR2_X1 U611 ( .A(n512), .B(G143), .Z(n517) );
  NAND2_X1 U612 ( .A1(n513), .A2(G214), .ZN(n515) );
  XOR2_X1 U613 ( .A(n518), .B(KEYINPUT100), .Z(n519) );
  XNOR2_X1 U614 ( .A(n520), .B(n519), .ZN(n521) );
  XNOR2_X1 U615 ( .A(n522), .B(n521), .ZN(n627) );
  NOR2_X1 U616 ( .A1(G902), .A2(n627), .ZN(n525) );
  XNOR2_X1 U617 ( .A(KEYINPUT13), .B(KEYINPUT103), .ZN(n523) );
  XOR2_X1 U618 ( .A(n526), .B(KEYINPUT7), .Z(n529) );
  NAND2_X1 U619 ( .A1(G217), .A2(n527), .ZN(n528) );
  XNOR2_X1 U620 ( .A(G116), .B(n530), .ZN(n531) );
  XNOR2_X1 U621 ( .A(n532), .B(n531), .ZN(n709) );
  NOR2_X1 U622 ( .A1(G902), .A2(n709), .ZN(n533) );
  XNOR2_X1 U623 ( .A(G478), .B(n533), .ZN(n553) );
  NOR2_X1 U624 ( .A1(n552), .A2(n553), .ZN(n587) );
  INV_X1 U625 ( .A(n542), .ZN(n608) );
  XOR2_X1 U626 ( .A(KEYINPUT64), .B(KEYINPUT22), .Z(n537) );
  NAND2_X1 U627 ( .A1(n552), .A2(n553), .ZN(n667) );
  INV_X1 U628 ( .A(n677), .ZN(n534) );
  NAND2_X1 U629 ( .A1(n535), .A2(n534), .ZN(n536) );
  XNOR2_X1 U630 ( .A(n537), .B(n536), .ZN(n541) );
  NAND2_X1 U631 ( .A1(n608), .A2(n541), .ZN(n549) );
  INV_X1 U632 ( .A(n580), .ZN(n571) );
  NAND2_X1 U633 ( .A1(n379), .A2(n571), .ZN(n538) );
  NOR2_X1 U634 ( .A1(n549), .A2(n538), .ZN(n648) );
  INV_X1 U635 ( .A(n539), .ZN(n540) );
  NAND2_X1 U636 ( .A1(n541), .A2(n540), .ZN(n544) );
  NAND2_X1 U637 ( .A1(n379), .A2(n542), .ZN(n543) );
  NOR2_X1 U638 ( .A1(n544), .A2(n543), .ZN(n546) );
  XNOR2_X1 U639 ( .A(KEYINPUT75), .B(KEYINPUT32), .ZN(n545) );
  XNOR2_X1 U640 ( .A(n546), .B(n545), .ZN(n740) );
  NAND2_X1 U641 ( .A1(n547), .A2(n740), .ZN(n557) );
  NAND2_X1 U642 ( .A1(n557), .A2(KEYINPUT44), .ZN(n556) );
  OR2_X1 U643 ( .A1(n379), .A2(n539), .ZN(n548) );
  NOR2_X1 U644 ( .A1(n549), .A2(n548), .ZN(n641) );
  NAND2_X1 U645 ( .A1(n580), .A2(n550), .ZN(n683) );
  XOR2_X1 U646 ( .A(KEYINPUT98), .B(KEYINPUT31), .Z(n551) );
  INV_X1 U647 ( .A(n552), .ZN(n554) );
  NOR2_X1 U648 ( .A1(n554), .A2(n553), .ZN(n658) );
  NOR2_X1 U649 ( .A1(n598), .A2(n658), .ZN(n669) );
  NOR2_X1 U650 ( .A1(G900), .A2(n558), .ZN(n559) );
  NAND2_X1 U651 ( .A1(n559), .A2(G953), .ZN(n561) );
  NAND2_X1 U652 ( .A1(n561), .A2(n560), .ZN(n562) );
  XNOR2_X1 U653 ( .A(n562), .B(KEYINPUT77), .ZN(n582) );
  NOR2_X1 U654 ( .A1(n582), .A2(n677), .ZN(n563) );
  NAND2_X1 U655 ( .A1(n379), .A2(n563), .ZN(n572) );
  XOR2_X1 U656 ( .A(KEYINPUT105), .B(n598), .Z(n642) );
  NAND2_X1 U657 ( .A1(n539), .A2(n642), .ZN(n564) );
  INV_X1 U658 ( .A(n609), .ZN(n566) );
  NOR2_X1 U659 ( .A1(n566), .A2(n565), .ZN(n569) );
  XNOR2_X1 U660 ( .A(KEYINPUT36), .B(KEYINPUT85), .ZN(n567) );
  NOR2_X1 U661 ( .A1(n608), .A2(n570), .ZN(n661) );
  NOR2_X1 U662 ( .A1(n572), .A2(n571), .ZN(n573) );
  XNOR2_X1 U663 ( .A(KEYINPUT28), .B(n573), .ZN(n575) );
  NAND2_X1 U664 ( .A1(n575), .A2(n574), .ZN(n602) );
  INV_X1 U665 ( .A(n602), .ZN(n577) );
  NAND2_X1 U666 ( .A1(n577), .A2(n576), .ZN(n649) );
  OR2_X1 U667 ( .A1(n669), .A2(n649), .ZN(n578) );
  NOR2_X1 U668 ( .A1(KEYINPUT47), .A2(n578), .ZN(n579) );
  NAND2_X1 U669 ( .A1(n580), .A2(n664), .ZN(n581) );
  XNOR2_X1 U670 ( .A(KEYINPUT30), .B(n581), .ZN(n586) );
  NOR2_X1 U671 ( .A1(n586), .A2(n585), .ZN(n596) );
  NAND2_X1 U672 ( .A1(n596), .A2(n587), .ZN(n588) );
  NOR2_X1 U673 ( .A1(n595), .A2(n588), .ZN(n653) );
  NAND2_X1 U674 ( .A1(n669), .A2(KEYINPUT47), .ZN(n589) );
  XNOR2_X1 U675 ( .A(n589), .B(KEYINPUT80), .ZN(n591) );
  NAND2_X1 U676 ( .A1(n649), .A2(KEYINPUT47), .ZN(n590) );
  NAND2_X1 U677 ( .A1(n591), .A2(n590), .ZN(n592) );
  NOR2_X1 U678 ( .A1(n653), .A2(n592), .ZN(n593) );
  NAND2_X1 U679 ( .A1(n594), .A2(n593), .ZN(n607) );
  XOR2_X1 U680 ( .A(KEYINPUT40), .B(KEYINPUT108), .Z(n599) );
  XNOR2_X1 U681 ( .A(KEYINPUT38), .B(n595), .ZN(n665) );
  NAND2_X1 U682 ( .A1(n596), .A2(n665), .ZN(n597) );
  NAND2_X1 U683 ( .A1(n665), .A2(n664), .ZN(n668) );
  NOR2_X1 U684 ( .A1(n667), .A2(n668), .ZN(n601) );
  XNOR2_X1 U685 ( .A(KEYINPUT41), .B(KEYINPUT110), .ZN(n600) );
  XNOR2_X1 U686 ( .A(n601), .B(n600), .ZN(n694) );
  NOR2_X1 U687 ( .A1(n694), .A2(n602), .ZN(n604) );
  XNOR2_X1 U688 ( .A(KEYINPUT111), .B(KEYINPUT42), .ZN(n603) );
  XNOR2_X1 U689 ( .A(n604), .B(n603), .ZN(n742) );
  NAND2_X1 U690 ( .A1(n737), .A2(n742), .ZN(n605) );
  XNOR2_X1 U691 ( .A(n605), .B(KEYINPUT46), .ZN(n606) );
  INV_X1 U692 ( .A(n608), .ZN(n675) );
  NAND2_X1 U693 ( .A1(n609), .A2(n664), .ZN(n610) );
  NOR2_X1 U694 ( .A1(n675), .A2(n610), .ZN(n612) );
  XNOR2_X1 U695 ( .A(KEYINPUT106), .B(KEYINPUT43), .ZN(n611) );
  XNOR2_X1 U696 ( .A(n612), .B(n611), .ZN(n613) );
  NOR2_X1 U697 ( .A1(n614), .A2(n613), .ZN(n615) );
  XOR2_X1 U698 ( .A(KEYINPUT107), .B(n615), .Z(n738) );
  NAND2_X1 U699 ( .A1(n616), .A2(n658), .ZN(n663) );
  INV_X1 U700 ( .A(n619), .ZN(n620) );
  XNOR2_X1 U701 ( .A(n620), .B(KEYINPUT82), .ZN(n621) );
  NAND2_X1 U702 ( .A1(n621), .A2(KEYINPUT2), .ZN(n622) );
  AND2_X1 U703 ( .A1(n697), .A2(G475), .ZN(n623) );
  NAND2_X1 U704 ( .A1(n633), .A2(n623), .ZN(n629) );
  XOR2_X1 U705 ( .A(KEYINPUT65), .B(KEYINPUT120), .Z(n625) );
  XNOR2_X1 U706 ( .A(KEYINPUT119), .B(KEYINPUT59), .ZN(n624) );
  XNOR2_X1 U707 ( .A(n625), .B(n624), .ZN(n626) );
  NOR2_X1 U708 ( .A1(n713), .A2(n630), .ZN(n632) );
  XOR2_X1 U709 ( .A(KEYINPUT62), .B(KEYINPUT113), .Z(n634) );
  NOR2_X2 U710 ( .A1(n638), .A2(n713), .ZN(n640) );
  XNOR2_X1 U711 ( .A(KEYINPUT87), .B(KEYINPUT63), .ZN(n639) );
  XNOR2_X1 U712 ( .A(n640), .B(n639), .ZN(G57) );
  XOR2_X1 U713 ( .A(G101), .B(n641), .Z(G3) );
  NAND2_X1 U714 ( .A1(n644), .A2(n642), .ZN(n643) );
  XNOR2_X1 U715 ( .A(n643), .B(G104), .ZN(G6) );
  XOR2_X1 U716 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n646) );
  NAND2_X1 U717 ( .A1(n644), .A2(n658), .ZN(n645) );
  XNOR2_X1 U718 ( .A(n646), .B(n645), .ZN(n647) );
  XNOR2_X1 U719 ( .A(G107), .B(n647), .ZN(G9) );
  XOR2_X1 U720 ( .A(G110), .B(n648), .Z(G12) );
  XOR2_X1 U721 ( .A(KEYINPUT114), .B(KEYINPUT29), .Z(n651) );
  INV_X1 U722 ( .A(n649), .ZN(n654) );
  NAND2_X1 U723 ( .A1(n654), .A2(n658), .ZN(n650) );
  XNOR2_X1 U724 ( .A(n651), .B(n650), .ZN(n652) );
  XNOR2_X1 U725 ( .A(G128), .B(n652), .ZN(G30) );
  XOR2_X1 U726 ( .A(G143), .B(n653), .Z(G45) );
  NAND2_X1 U727 ( .A1(n654), .A2(n642), .ZN(n655) );
  XNOR2_X1 U728 ( .A(n655), .B(G146), .ZN(G48) );
  NAND2_X1 U729 ( .A1(n657), .A2(n642), .ZN(n656) );
  XNOR2_X1 U730 ( .A(n656), .B(G113), .ZN(G15) );
  XOR2_X1 U731 ( .A(G116), .B(KEYINPUT115), .Z(n660) );
  NAND2_X1 U732 ( .A1(n658), .A2(n657), .ZN(n659) );
  XNOR2_X1 U733 ( .A(n660), .B(n659), .ZN(G18) );
  XNOR2_X1 U734 ( .A(G125), .B(n661), .ZN(n662) );
  XNOR2_X1 U735 ( .A(n662), .B(KEYINPUT37), .ZN(G27) );
  XNOR2_X1 U736 ( .A(G134), .B(n663), .ZN(G36) );
  NOR2_X1 U737 ( .A1(n665), .A2(n664), .ZN(n666) );
  NOR2_X1 U738 ( .A1(n667), .A2(n666), .ZN(n671) );
  NOR2_X1 U739 ( .A1(n669), .A2(n668), .ZN(n670) );
  NOR2_X1 U740 ( .A1(n671), .A2(n670), .ZN(n672) );
  NOR2_X1 U741 ( .A1(n693), .A2(n672), .ZN(n689) );
  XNOR2_X1 U742 ( .A(KEYINPUT116), .B(KEYINPUT51), .ZN(n673) );
  XNOR2_X1 U743 ( .A(n673), .B(KEYINPUT117), .ZN(n686) );
  OR2_X1 U744 ( .A1(n675), .A2(n674), .ZN(n676) );
  XNOR2_X1 U745 ( .A(n676), .B(KEYINPUT50), .ZN(n682) );
  NAND2_X1 U746 ( .A1(n379), .A2(n677), .ZN(n679) );
  XNOR2_X1 U747 ( .A(KEYINPUT49), .B(n679), .ZN(n680) );
  NOR2_X1 U748 ( .A1(n580), .A2(n680), .ZN(n681) );
  NAND2_X1 U749 ( .A1(n682), .A2(n681), .ZN(n684) );
  NAND2_X1 U750 ( .A1(n684), .A2(n683), .ZN(n685) );
  XOR2_X1 U751 ( .A(n686), .B(n685), .Z(n687) );
  NOR2_X1 U752 ( .A1(n694), .A2(n687), .ZN(n688) );
  NOR2_X1 U753 ( .A1(n689), .A2(n688), .ZN(n690) );
  XNOR2_X1 U754 ( .A(n690), .B(KEYINPUT52), .ZN(n691) );
  NOR2_X1 U755 ( .A1(n692), .A2(n691), .ZN(n696) );
  NOR2_X1 U756 ( .A1(n694), .A2(n693), .ZN(n695) );
  NOR2_X1 U757 ( .A1(n696), .A2(n695), .ZN(n700) );
  NAND2_X1 U758 ( .A1(n698), .A2(n697), .ZN(n699) );
  XOR2_X1 U759 ( .A(KEYINPUT54), .B(KEYINPUT55), .Z(n703) );
  XNOR2_X1 U760 ( .A(n701), .B(KEYINPUT86), .ZN(n702) );
  XNOR2_X1 U761 ( .A(n703), .B(n702), .ZN(n704) );
  XOR2_X1 U762 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n705) );
  NOR2_X1 U763 ( .A1(n713), .A2(n707), .ZN(G54) );
  XNOR2_X1 U764 ( .A(n709), .B(n708), .ZN(n710) );
  NOR2_X1 U765 ( .A1(n713), .A2(n710), .ZN(G63) );
  NOR2_X1 U766 ( .A1(n713), .A2(n712), .ZN(G66) );
  XNOR2_X1 U767 ( .A(n714), .B(KEYINPUT122), .ZN(n715) );
  XNOR2_X1 U768 ( .A(n715), .B(KEYINPUT123), .ZN(n717) );
  NOR2_X1 U769 ( .A1(n717), .A2(n716), .ZN(n725) );
  XOR2_X1 U770 ( .A(KEYINPUT121), .B(KEYINPUT61), .Z(n719) );
  NAND2_X1 U771 ( .A1(G224), .A2(G953), .ZN(n718) );
  XNOR2_X1 U772 ( .A(n719), .B(n718), .ZN(n720) );
  NAND2_X1 U773 ( .A1(n720), .A2(G898), .ZN(n723) );
  NAND2_X1 U774 ( .A1(n721), .A2(n457), .ZN(n722) );
  NAND2_X1 U775 ( .A1(n723), .A2(n722), .ZN(n724) );
  XNOR2_X1 U776 ( .A(n725), .B(n724), .ZN(G69) );
  XOR2_X1 U777 ( .A(n727), .B(n726), .Z(n728) );
  XOR2_X1 U778 ( .A(KEYINPUT124), .B(n728), .Z(n731) );
  XOR2_X1 U779 ( .A(n731), .B(n729), .Z(n730) );
  NAND2_X1 U780 ( .A1(n730), .A2(n457), .ZN(n735) );
  XNOR2_X1 U781 ( .A(n731), .B(G227), .ZN(n732) );
  NOR2_X1 U782 ( .A1(n457), .A2(n732), .ZN(n733) );
  NAND2_X1 U783 ( .A1(G900), .A2(n733), .ZN(n734) );
  NAND2_X1 U784 ( .A1(n735), .A2(n734), .ZN(n736) );
  XNOR2_X1 U785 ( .A(KEYINPUT125), .B(n736), .ZN(G72) );
  XNOR2_X1 U786 ( .A(G131), .B(n737), .ZN(G33) );
  XOR2_X1 U787 ( .A(G140), .B(n738), .Z(G42) );
  XOR2_X1 U788 ( .A(n739), .B(G122), .Z(G24) );
  XNOR2_X1 U789 ( .A(G119), .B(n740), .ZN(n741) );
  XNOR2_X1 U790 ( .A(n741), .B(KEYINPUT126), .ZN(G21) );
  XOR2_X1 U791 ( .A(G137), .B(n742), .Z(n743) );
  XNOR2_X1 U792 ( .A(KEYINPUT127), .B(n743), .ZN(G39) );
endmodule

