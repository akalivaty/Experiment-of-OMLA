

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302,
         n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313,
         n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324,
         n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335,
         n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346,
         n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582;

  XNOR2_X1 U324 ( .A(n407), .B(n406), .ZN(n538) );
  NAND2_X1 U325 ( .A1(n482), .A2(n481), .ZN(n483) );
  XOR2_X1 U326 ( .A(n324), .B(n323), .Z(n521) );
  XNOR2_X1 U327 ( .A(n309), .B(n412), .ZN(n310) );
  XOR2_X1 U328 ( .A(KEYINPUT17), .B(KEYINPUT19), .Z(n292) );
  XOR2_X1 U329 ( .A(n318), .B(n388), .Z(n293) );
  OR2_X1 U330 ( .A1(n512), .A2(n510), .ZN(n451) );
  NOR2_X1 U331 ( .A1(n461), .A2(n452), .ZN(n453) );
  XNOR2_X1 U332 ( .A(n297), .B(n296), .ZN(n299) );
  XNOR2_X1 U333 ( .A(n299), .B(n298), .ZN(n301) );
  XNOR2_X1 U334 ( .A(KEYINPUT48), .B(KEYINPUT112), .ZN(n406) );
  NOR2_X1 U335 ( .A1(n512), .A2(n443), .ZN(n553) );
  XNOR2_X1 U336 ( .A(n483), .B(KEYINPUT37), .ZN(n506) );
  XNOR2_X1 U337 ( .A(G169GAT), .B(n314), .ZN(n416) );
  INV_X1 U338 ( .A(G190GAT), .ZN(n444) );
  XNOR2_X1 U339 ( .A(n311), .B(n310), .ZN(n547) );
  XNOR2_X1 U340 ( .A(KEYINPUT38), .B(n485), .ZN(n493) );
  XNOR2_X1 U341 ( .A(n445), .B(n444), .ZN(n446) );
  XNOR2_X1 U342 ( .A(n447), .B(n446), .ZN(G1351GAT) );
  XOR2_X1 U343 ( .A(KEYINPUT10), .B(KEYINPUT11), .Z(n295) );
  XNOR2_X1 U344 ( .A(KEYINPUT64), .B(KEYINPUT9), .ZN(n294) );
  XNOR2_X1 U345 ( .A(n295), .B(n294), .ZN(n297) );
  XOR2_X1 U346 ( .A(KEYINPUT75), .B(KEYINPUT76), .Z(n296) );
  XOR2_X1 U347 ( .A(G43GAT), .B(G134GAT), .Z(n315) );
  XOR2_X1 U348 ( .A(G50GAT), .B(G162GAT), .Z(n329) );
  XNOR2_X1 U349 ( .A(n315), .B(n329), .ZN(n298) );
  NAND2_X1 U350 ( .A1(G232GAT), .A2(G233GAT), .ZN(n300) );
  XNOR2_X1 U351 ( .A(n301), .B(n300), .ZN(n311) );
  XOR2_X1 U352 ( .A(G29GAT), .B(KEYINPUT7), .Z(n303) );
  XNOR2_X1 U353 ( .A(KEYINPUT68), .B(KEYINPUT8), .ZN(n302) );
  XNOR2_X1 U354 ( .A(n303), .B(n302), .ZN(n374) );
  XOR2_X1 U355 ( .A(KEYINPUT74), .B(KEYINPUT73), .Z(n305) );
  XNOR2_X1 U356 ( .A(G106GAT), .B(G85GAT), .ZN(n304) );
  XNOR2_X1 U357 ( .A(n305), .B(n304), .ZN(n306) );
  XOR2_X1 U358 ( .A(G99GAT), .B(n306), .Z(n358) );
  XNOR2_X1 U359 ( .A(n374), .B(n358), .ZN(n309) );
  XOR2_X1 U360 ( .A(G92GAT), .B(G218GAT), .Z(n308) );
  XNOR2_X1 U361 ( .A(G36GAT), .B(G190GAT), .ZN(n307) );
  XNOR2_X1 U362 ( .A(n308), .B(n307), .ZN(n412) );
  XNOR2_X1 U363 ( .A(KEYINPUT77), .B(n547), .ZN(n532) );
  XNOR2_X1 U364 ( .A(G113GAT), .B(KEYINPUT0), .ZN(n312) );
  XNOR2_X1 U365 ( .A(n312), .B(KEYINPUT81), .ZN(n434) );
  XOR2_X1 U366 ( .A(G120GAT), .B(G71GAT), .Z(n347) );
  XOR2_X1 U367 ( .A(n434), .B(n347), .Z(n317) );
  XNOR2_X1 U368 ( .A(KEYINPUT18), .B(G176GAT), .ZN(n313) );
  XNOR2_X1 U369 ( .A(n292), .B(n313), .ZN(n314) );
  XOR2_X1 U370 ( .A(n416), .B(n315), .Z(n316) );
  XNOR2_X1 U371 ( .A(n317), .B(n316), .ZN(n318) );
  XOR2_X1 U372 ( .A(G15GAT), .B(G127GAT), .Z(n388) );
  XNOR2_X1 U373 ( .A(G99GAT), .B(G190GAT), .ZN(n319) );
  XNOR2_X1 U374 ( .A(n293), .B(n319), .ZN(n324) );
  XOR2_X1 U375 ( .A(KEYINPUT20), .B(G183GAT), .Z(n321) );
  NAND2_X1 U376 ( .A1(G227GAT), .A2(G233GAT), .ZN(n320) );
  XNOR2_X1 U377 ( .A(n321), .B(n320), .ZN(n322) );
  XOR2_X1 U378 ( .A(KEYINPUT82), .B(n322), .Z(n323) );
  INV_X1 U379 ( .A(n521), .ZN(n512) );
  XOR2_X1 U380 ( .A(G204GAT), .B(KEYINPUT21), .Z(n326) );
  XNOR2_X1 U381 ( .A(G197GAT), .B(KEYINPUT86), .ZN(n325) );
  XNOR2_X1 U382 ( .A(n326), .B(n325), .ZN(n413) );
  XOR2_X1 U383 ( .A(G148GAT), .B(KEYINPUT2), .Z(n328) );
  XNOR2_X1 U384 ( .A(G141GAT), .B(KEYINPUT3), .ZN(n327) );
  XNOR2_X1 U385 ( .A(n328), .B(n327), .ZN(n426) );
  XOR2_X1 U386 ( .A(n426), .B(n329), .Z(n331) );
  XNOR2_X1 U387 ( .A(G218GAT), .B(G106GAT), .ZN(n330) );
  XNOR2_X1 U388 ( .A(n331), .B(n330), .ZN(n335) );
  XOR2_X1 U389 ( .A(KEYINPUT87), .B(KEYINPUT23), .Z(n333) );
  NAND2_X1 U390 ( .A1(G228GAT), .A2(G233GAT), .ZN(n332) );
  XNOR2_X1 U391 ( .A(n333), .B(n332), .ZN(n334) );
  XOR2_X1 U392 ( .A(n335), .B(n334), .Z(n340) );
  XOR2_X1 U393 ( .A(KEYINPUT85), .B(KEYINPUT22), .Z(n337) );
  XNOR2_X1 U394 ( .A(G211GAT), .B(KEYINPUT84), .ZN(n336) );
  XNOR2_X1 U395 ( .A(n337), .B(n336), .ZN(n338) );
  XNOR2_X1 U396 ( .A(n338), .B(KEYINPUT24), .ZN(n339) );
  XNOR2_X1 U397 ( .A(n340), .B(n339), .ZN(n341) );
  XNOR2_X1 U398 ( .A(n413), .B(n341), .ZN(n343) );
  XOR2_X1 U399 ( .A(G22GAT), .B(G155GAT), .Z(n342) );
  XOR2_X1 U400 ( .A(G78GAT), .B(n342), .Z(n393) );
  XOR2_X1 U401 ( .A(n343), .B(n393), .Z(n461) );
  XOR2_X1 U402 ( .A(KEYINPUT46), .B(KEYINPUT110), .Z(n380) );
  XOR2_X1 U403 ( .A(KEYINPUT33), .B(G148GAT), .Z(n345) );
  XNOR2_X1 U404 ( .A(G204GAT), .B(G78GAT), .ZN(n344) );
  XNOR2_X1 U405 ( .A(n345), .B(n344), .ZN(n346) );
  XOR2_X1 U406 ( .A(n346), .B(G92GAT), .Z(n349) );
  XNOR2_X1 U407 ( .A(G176GAT), .B(n347), .ZN(n348) );
  XNOR2_X1 U408 ( .A(n349), .B(n348), .ZN(n354) );
  XNOR2_X1 U409 ( .A(G57GAT), .B(KEYINPUT13), .ZN(n350) );
  XNOR2_X1 U410 ( .A(n350), .B(KEYINPUT70), .ZN(n389) );
  XOR2_X1 U411 ( .A(n389), .B(KEYINPUT71), .Z(n352) );
  NAND2_X1 U412 ( .A1(G230GAT), .A2(G233GAT), .ZN(n351) );
  XNOR2_X1 U413 ( .A(n352), .B(n351), .ZN(n353) );
  XOR2_X1 U414 ( .A(n354), .B(n353), .Z(n360) );
  XOR2_X1 U415 ( .A(KEYINPUT32), .B(KEYINPUT72), .Z(n356) );
  XNOR2_X1 U416 ( .A(G64GAT), .B(KEYINPUT31), .ZN(n355) );
  XNOR2_X1 U417 ( .A(n356), .B(n355), .ZN(n357) );
  XNOR2_X1 U418 ( .A(n358), .B(n357), .ZN(n359) );
  XNOR2_X1 U419 ( .A(n360), .B(n359), .ZN(n568) );
  XNOR2_X1 U420 ( .A(n568), .B(KEYINPUT41), .ZN(n524) );
  INV_X1 U421 ( .A(n524), .ZN(n552) );
  XOR2_X1 U422 ( .A(G1GAT), .B(G141GAT), .Z(n362) );
  XNOR2_X1 U423 ( .A(G197GAT), .B(G22GAT), .ZN(n361) );
  XNOR2_X1 U424 ( .A(n362), .B(n361), .ZN(n378) );
  XOR2_X1 U425 ( .A(KEYINPUT30), .B(KEYINPUT29), .Z(n364) );
  XNOR2_X1 U426 ( .A(KEYINPUT69), .B(KEYINPUT66), .ZN(n363) );
  XNOR2_X1 U427 ( .A(n364), .B(n363), .ZN(n372) );
  NAND2_X1 U428 ( .A1(G229GAT), .A2(G233GAT), .ZN(n370) );
  XOR2_X1 U429 ( .A(G113GAT), .B(G15GAT), .Z(n366) );
  XNOR2_X1 U430 ( .A(G169GAT), .B(G36GAT), .ZN(n365) );
  XNOR2_X1 U431 ( .A(n366), .B(n365), .ZN(n368) );
  XOR2_X1 U432 ( .A(G50GAT), .B(G43GAT), .Z(n367) );
  XNOR2_X1 U433 ( .A(n368), .B(n367), .ZN(n369) );
  XNOR2_X1 U434 ( .A(n370), .B(n369), .ZN(n371) );
  XNOR2_X1 U435 ( .A(n372), .B(n371), .ZN(n373) );
  XOR2_X1 U436 ( .A(n373), .B(KEYINPUT67), .Z(n376) );
  XNOR2_X1 U437 ( .A(n374), .B(G8GAT), .ZN(n375) );
  XNOR2_X1 U438 ( .A(n376), .B(n375), .ZN(n377) );
  XNOR2_X1 U439 ( .A(n378), .B(n377), .ZN(n522) );
  INV_X1 U440 ( .A(n522), .ZN(n564) );
  NAND2_X1 U441 ( .A1(n552), .A2(n564), .ZN(n379) );
  XNOR2_X1 U442 ( .A(n380), .B(n379), .ZN(n381) );
  NOR2_X1 U443 ( .A1(n547), .A2(n381), .ZN(n398) );
  XOR2_X1 U444 ( .A(KEYINPUT78), .B(G64GAT), .Z(n383) );
  XNOR2_X1 U445 ( .A(G183GAT), .B(G211GAT), .ZN(n382) );
  XNOR2_X1 U446 ( .A(n383), .B(n382), .ZN(n384) );
  XOR2_X1 U447 ( .A(G8GAT), .B(n384), .Z(n410) );
  XOR2_X1 U448 ( .A(KEYINPUT14), .B(KEYINPUT79), .Z(n386) );
  XNOR2_X1 U449 ( .A(G1GAT), .B(G71GAT), .ZN(n385) );
  XNOR2_X1 U450 ( .A(n386), .B(n385), .ZN(n387) );
  XNOR2_X1 U451 ( .A(n410), .B(n387), .ZN(n397) );
  XOR2_X1 U452 ( .A(n389), .B(n388), .Z(n391) );
  NAND2_X1 U453 ( .A1(G231GAT), .A2(G233GAT), .ZN(n390) );
  XNOR2_X1 U454 ( .A(n391), .B(n390), .ZN(n392) );
  XOR2_X1 U455 ( .A(n392), .B(KEYINPUT15), .Z(n395) );
  XNOR2_X1 U456 ( .A(n393), .B(KEYINPUT12), .ZN(n394) );
  XNOR2_X1 U457 ( .A(n395), .B(n394), .ZN(n396) );
  XOR2_X1 U458 ( .A(n397), .B(n396), .Z(n448) );
  XOR2_X1 U459 ( .A(n448), .B(KEYINPUT109), .Z(n559) );
  NAND2_X1 U460 ( .A1(n398), .A2(n559), .ZN(n399) );
  XNOR2_X1 U461 ( .A(n399), .B(KEYINPUT47), .ZN(n405) );
  XNOR2_X1 U462 ( .A(KEYINPUT36), .B(n532), .ZN(n580) );
  NOR2_X1 U463 ( .A1(n580), .A2(n448), .ZN(n401) );
  XOR2_X1 U464 ( .A(KEYINPUT45), .B(KEYINPUT111), .Z(n400) );
  XNOR2_X1 U465 ( .A(n401), .B(n400), .ZN(n402) );
  NAND2_X1 U466 ( .A1(n402), .A2(n522), .ZN(n403) );
  NOR2_X1 U467 ( .A1(n403), .A2(n568), .ZN(n404) );
  NOR2_X1 U468 ( .A1(n405), .A2(n404), .ZN(n407) );
  XOR2_X1 U469 ( .A(KEYINPUT92), .B(KEYINPUT93), .Z(n409) );
  NAND2_X1 U470 ( .A1(G226GAT), .A2(G233GAT), .ZN(n408) );
  XNOR2_X1 U471 ( .A(n409), .B(n408), .ZN(n411) );
  XOR2_X1 U472 ( .A(n411), .B(n410), .Z(n415) );
  XNOR2_X1 U473 ( .A(n413), .B(n412), .ZN(n414) );
  XNOR2_X1 U474 ( .A(n415), .B(n414), .ZN(n417) );
  XOR2_X1 U475 ( .A(n417), .B(n416), .Z(n510) );
  XOR2_X1 U476 ( .A(n510), .B(KEYINPUT119), .Z(n418) );
  NOR2_X1 U477 ( .A1(n538), .A2(n418), .ZN(n419) );
  XNOR2_X1 U478 ( .A(n419), .B(KEYINPUT54), .ZN(n441) );
  XOR2_X1 U479 ( .A(KEYINPUT88), .B(G155GAT), .Z(n421) );
  XNOR2_X1 U480 ( .A(G127GAT), .B(G120GAT), .ZN(n420) );
  XNOR2_X1 U481 ( .A(n421), .B(n420), .ZN(n425) );
  XOR2_X1 U482 ( .A(KEYINPUT6), .B(KEYINPUT90), .Z(n423) );
  XNOR2_X1 U483 ( .A(KEYINPUT5), .B(KEYINPUT4), .ZN(n422) );
  XNOR2_X1 U484 ( .A(n423), .B(n422), .ZN(n424) );
  XOR2_X1 U485 ( .A(n425), .B(n424), .Z(n431) );
  XOR2_X1 U486 ( .A(G85GAT), .B(n426), .Z(n428) );
  XNOR2_X1 U487 ( .A(G29GAT), .B(G162GAT), .ZN(n427) );
  XNOR2_X1 U488 ( .A(n428), .B(n427), .ZN(n429) );
  XNOR2_X1 U489 ( .A(G134GAT), .B(n429), .ZN(n430) );
  XNOR2_X1 U490 ( .A(n431), .B(n430), .ZN(n440) );
  XOR2_X1 U491 ( .A(G57GAT), .B(KEYINPUT89), .Z(n433) );
  XNOR2_X1 U492 ( .A(KEYINPUT91), .B(KEYINPUT1), .ZN(n432) );
  XNOR2_X1 U493 ( .A(n433), .B(n432), .ZN(n438) );
  XOR2_X1 U494 ( .A(n434), .B(G1GAT), .Z(n436) );
  NAND2_X1 U495 ( .A1(G225GAT), .A2(G233GAT), .ZN(n435) );
  XNOR2_X1 U496 ( .A(n436), .B(n435), .ZN(n437) );
  XOR2_X1 U497 ( .A(n438), .B(n437), .Z(n439) );
  XNOR2_X1 U498 ( .A(n440), .B(n439), .ZN(n507) );
  NAND2_X1 U499 ( .A1(n441), .A2(n507), .ZN(n562) );
  NOR2_X1 U500 ( .A1(n461), .A2(n562), .ZN(n442) );
  XNOR2_X1 U501 ( .A(n442), .B(KEYINPUT55), .ZN(n443) );
  INV_X1 U502 ( .A(n553), .ZN(n558) );
  NOR2_X1 U503 ( .A1(n532), .A2(n558), .ZN(n447) );
  XNOR2_X1 U504 ( .A(KEYINPUT58), .B(KEYINPUT122), .ZN(n445) );
  NOR2_X1 U505 ( .A1(n568), .A2(n522), .ZN(n484) );
  XOR2_X1 U506 ( .A(KEYINPUT80), .B(KEYINPUT16), .Z(n450) );
  INV_X1 U507 ( .A(n448), .ZN(n572) );
  NAND2_X1 U508 ( .A1(n572), .A2(n532), .ZN(n449) );
  XNOR2_X1 U509 ( .A(n450), .B(n449), .ZN(n467) );
  XNOR2_X1 U510 ( .A(KEYINPUT95), .B(n451), .ZN(n452) );
  XNOR2_X1 U511 ( .A(n453), .B(KEYINPUT25), .ZN(n456) );
  NAND2_X1 U512 ( .A1(n461), .A2(n512), .ZN(n454) );
  XOR2_X1 U513 ( .A(KEYINPUT26), .B(n454), .Z(n561) );
  XOR2_X1 U514 ( .A(n510), .B(KEYINPUT27), .Z(n459) );
  NAND2_X1 U515 ( .A1(n561), .A2(n459), .ZN(n455) );
  NAND2_X1 U516 ( .A1(n456), .A2(n455), .ZN(n457) );
  NAND2_X1 U517 ( .A1(n457), .A2(n507), .ZN(n458) );
  XNOR2_X1 U518 ( .A(n458), .B(KEYINPUT96), .ZN(n466) );
  XNOR2_X1 U519 ( .A(KEYINPUT83), .B(n521), .ZN(n464) );
  INV_X1 U520 ( .A(n459), .ZN(n460) );
  NOR2_X1 U521 ( .A1(n460), .A2(n507), .ZN(n536) );
  XNOR2_X1 U522 ( .A(KEYINPUT65), .B(KEYINPUT28), .ZN(n462) );
  XNOR2_X1 U523 ( .A(n462), .B(n461), .ZN(n516) );
  NAND2_X1 U524 ( .A1(n536), .A2(n516), .ZN(n519) );
  XOR2_X1 U525 ( .A(KEYINPUT94), .B(n519), .Z(n463) );
  NAND2_X1 U526 ( .A1(n464), .A2(n463), .ZN(n465) );
  NAND2_X1 U527 ( .A1(n466), .A2(n465), .ZN(n482) );
  AND2_X1 U528 ( .A1(n467), .A2(n482), .ZN(n496) );
  NAND2_X1 U529 ( .A1(n484), .A2(n496), .ZN(n468) );
  XOR2_X1 U530 ( .A(KEYINPUT97), .B(n468), .Z(n477) );
  NOR2_X1 U531 ( .A1(n507), .A2(n477), .ZN(n469) );
  XOR2_X1 U532 ( .A(G1GAT), .B(n469), .Z(n470) );
  XNOR2_X1 U533 ( .A(KEYINPUT34), .B(n470), .ZN(G1324GAT) );
  NOR2_X1 U534 ( .A1(n510), .A2(n477), .ZN(n471) );
  XOR2_X1 U535 ( .A(KEYINPUT98), .B(n471), .Z(n472) );
  XNOR2_X1 U536 ( .A(G8GAT), .B(n472), .ZN(G1325GAT) );
  NOR2_X1 U537 ( .A1(n477), .A2(n512), .ZN(n476) );
  XOR2_X1 U538 ( .A(KEYINPUT99), .B(KEYINPUT100), .Z(n474) );
  XNOR2_X1 U539 ( .A(G15GAT), .B(KEYINPUT35), .ZN(n473) );
  XNOR2_X1 U540 ( .A(n474), .B(n473), .ZN(n475) );
  XNOR2_X1 U541 ( .A(n476), .B(n475), .ZN(G1326GAT) );
  NOR2_X1 U542 ( .A1(n516), .A2(n477), .ZN(n478) );
  XOR2_X1 U543 ( .A(G22GAT), .B(n478), .Z(G1327GAT) );
  XOR2_X1 U544 ( .A(KEYINPUT103), .B(KEYINPUT102), .Z(n480) );
  XNOR2_X1 U545 ( .A(G29GAT), .B(KEYINPUT39), .ZN(n479) );
  XNOR2_X1 U546 ( .A(n480), .B(n479), .ZN(n487) );
  NOR2_X1 U547 ( .A1(n580), .A2(n572), .ZN(n481) );
  NAND2_X1 U548 ( .A1(n506), .A2(n484), .ZN(n485) );
  NOR2_X1 U549 ( .A1(n493), .A2(n507), .ZN(n486) );
  XOR2_X1 U550 ( .A(n487), .B(n486), .Z(n488) );
  XNOR2_X1 U551 ( .A(KEYINPUT101), .B(n488), .ZN(G1328GAT) );
  NOR2_X1 U552 ( .A1(n493), .A2(n510), .ZN(n489) );
  XOR2_X1 U553 ( .A(G36GAT), .B(n489), .Z(G1329GAT) );
  NOR2_X1 U554 ( .A1(n493), .A2(n512), .ZN(n491) );
  XNOR2_X1 U555 ( .A(KEYINPUT40), .B(KEYINPUT104), .ZN(n490) );
  XNOR2_X1 U556 ( .A(n491), .B(n490), .ZN(n492) );
  XOR2_X1 U557 ( .A(G43GAT), .B(n492), .Z(G1330GAT) );
  NOR2_X1 U558 ( .A1(n493), .A2(n516), .ZN(n495) );
  XNOR2_X1 U559 ( .A(G50GAT), .B(KEYINPUT105), .ZN(n494) );
  XNOR2_X1 U560 ( .A(n495), .B(n494), .ZN(G1331GAT) );
  NOR2_X1 U561 ( .A1(n564), .A2(n524), .ZN(n505) );
  NAND2_X1 U562 ( .A1(n496), .A2(n505), .ZN(n502) );
  NOR2_X1 U563 ( .A1(n507), .A2(n502), .ZN(n497) );
  XOR2_X1 U564 ( .A(G57GAT), .B(n497), .Z(n498) );
  XNOR2_X1 U565 ( .A(KEYINPUT42), .B(n498), .ZN(G1332GAT) );
  NOR2_X1 U566 ( .A1(n510), .A2(n502), .ZN(n499) );
  XOR2_X1 U567 ( .A(G64GAT), .B(n499), .Z(G1333GAT) );
  NOR2_X1 U568 ( .A1(n512), .A2(n502), .ZN(n500) );
  XOR2_X1 U569 ( .A(KEYINPUT106), .B(n500), .Z(n501) );
  XNOR2_X1 U570 ( .A(G71GAT), .B(n501), .ZN(G1334GAT) );
  NOR2_X1 U571 ( .A1(n516), .A2(n502), .ZN(n504) );
  XNOR2_X1 U572 ( .A(G78GAT), .B(KEYINPUT43), .ZN(n503) );
  XNOR2_X1 U573 ( .A(n504), .B(n503), .ZN(G1335GAT) );
  NAND2_X1 U574 ( .A1(n506), .A2(n505), .ZN(n515) );
  NOR2_X1 U575 ( .A1(n507), .A2(n515), .ZN(n509) );
  XNOR2_X1 U576 ( .A(G85GAT), .B(KEYINPUT107), .ZN(n508) );
  XNOR2_X1 U577 ( .A(n509), .B(n508), .ZN(G1336GAT) );
  NOR2_X1 U578 ( .A1(n510), .A2(n515), .ZN(n511) );
  XOR2_X1 U579 ( .A(G92GAT), .B(n511), .Z(G1337GAT) );
  NOR2_X1 U580 ( .A1(n512), .A2(n515), .ZN(n513) );
  XOR2_X1 U581 ( .A(KEYINPUT108), .B(n513), .Z(n514) );
  XNOR2_X1 U582 ( .A(G99GAT), .B(n514), .ZN(G1338GAT) );
  NOR2_X1 U583 ( .A1(n516), .A2(n515), .ZN(n517) );
  XOR2_X1 U584 ( .A(KEYINPUT44), .B(n517), .Z(n518) );
  XNOR2_X1 U585 ( .A(G106GAT), .B(n518), .ZN(G1339GAT) );
  NOR2_X1 U586 ( .A1(n538), .A2(n519), .ZN(n520) );
  NAND2_X1 U587 ( .A1(n521), .A2(n520), .ZN(n531) );
  NOR2_X1 U588 ( .A1(n522), .A2(n531), .ZN(n523) );
  XOR2_X1 U589 ( .A(G113GAT), .B(n523), .Z(G1340GAT) );
  NOR2_X1 U590 ( .A1(n524), .A2(n531), .ZN(n526) );
  XNOR2_X1 U591 ( .A(KEYINPUT113), .B(KEYINPUT49), .ZN(n525) );
  XNOR2_X1 U592 ( .A(n526), .B(n525), .ZN(n527) );
  XOR2_X1 U593 ( .A(G120GAT), .B(n527), .Z(G1341GAT) );
  NOR2_X1 U594 ( .A1(n559), .A2(n531), .ZN(n529) );
  XNOR2_X1 U595 ( .A(KEYINPUT50), .B(KEYINPUT114), .ZN(n528) );
  XNOR2_X1 U596 ( .A(n529), .B(n528), .ZN(n530) );
  XOR2_X1 U597 ( .A(G127GAT), .B(n530), .Z(G1342GAT) );
  NOR2_X1 U598 ( .A1(n532), .A2(n531), .ZN(n534) );
  XNOR2_X1 U599 ( .A(KEYINPUT115), .B(KEYINPUT51), .ZN(n533) );
  XNOR2_X1 U600 ( .A(n534), .B(n533), .ZN(n535) );
  XOR2_X1 U601 ( .A(G134GAT), .B(n535), .Z(G1343GAT) );
  NAND2_X1 U602 ( .A1(n536), .A2(n561), .ZN(n537) );
  NOR2_X1 U603 ( .A1(n538), .A2(n537), .ZN(n548) );
  NAND2_X1 U604 ( .A1(n548), .A2(n564), .ZN(n539) );
  XNOR2_X1 U605 ( .A(n539), .B(KEYINPUT116), .ZN(n540) );
  XNOR2_X1 U606 ( .A(G141GAT), .B(n540), .ZN(G1344GAT) );
  XOR2_X1 U607 ( .A(KEYINPUT52), .B(KEYINPUT117), .Z(n542) );
  NAND2_X1 U608 ( .A1(n548), .A2(n552), .ZN(n541) );
  XNOR2_X1 U609 ( .A(n542), .B(n541), .ZN(n544) );
  XOR2_X1 U610 ( .A(G148GAT), .B(KEYINPUT53), .Z(n543) );
  XNOR2_X1 U611 ( .A(n544), .B(n543), .ZN(G1345GAT) );
  NAND2_X1 U612 ( .A1(n548), .A2(n572), .ZN(n545) );
  XNOR2_X1 U613 ( .A(n545), .B(KEYINPUT118), .ZN(n546) );
  XNOR2_X1 U614 ( .A(G155GAT), .B(n546), .ZN(G1346GAT) );
  NAND2_X1 U615 ( .A1(n548), .A2(n547), .ZN(n549) );
  XNOR2_X1 U616 ( .A(n549), .B(G162GAT), .ZN(G1347GAT) );
  NAND2_X1 U617 ( .A1(n553), .A2(n564), .ZN(n550) );
  XNOR2_X1 U618 ( .A(n550), .B(KEYINPUT120), .ZN(n551) );
  XNOR2_X1 U619 ( .A(G169GAT), .B(n551), .ZN(G1348GAT) );
  XOR2_X1 U620 ( .A(KEYINPUT121), .B(KEYINPUT57), .Z(n555) );
  NAND2_X1 U621 ( .A1(n553), .A2(n552), .ZN(n554) );
  XNOR2_X1 U622 ( .A(n555), .B(n554), .ZN(n557) );
  XOR2_X1 U623 ( .A(G176GAT), .B(KEYINPUT56), .Z(n556) );
  XNOR2_X1 U624 ( .A(n557), .B(n556), .ZN(G1349GAT) );
  NOR2_X1 U625 ( .A1(n559), .A2(n558), .ZN(n560) );
  XOR2_X1 U626 ( .A(G183GAT), .B(n560), .Z(G1350GAT) );
  XOR2_X1 U627 ( .A(KEYINPUT60), .B(KEYINPUT59), .Z(n566) );
  INV_X1 U628 ( .A(n561), .ZN(n563) );
  NOR2_X1 U629 ( .A1(n563), .A2(n562), .ZN(n578) );
  NAND2_X1 U630 ( .A1(n578), .A2(n564), .ZN(n565) );
  XNOR2_X1 U631 ( .A(n566), .B(n565), .ZN(n567) );
  XNOR2_X1 U632 ( .A(G197GAT), .B(n567), .ZN(G1352GAT) );
  XOR2_X1 U633 ( .A(KEYINPUT123), .B(KEYINPUT61), .Z(n570) );
  NAND2_X1 U634 ( .A1(n578), .A2(n568), .ZN(n569) );
  XNOR2_X1 U635 ( .A(n570), .B(n569), .ZN(n571) );
  XOR2_X1 U636 ( .A(G204GAT), .B(n571), .Z(G1353GAT) );
  XOR2_X1 U637 ( .A(KEYINPUT124), .B(KEYINPUT125), .Z(n574) );
  NAND2_X1 U638 ( .A1(n578), .A2(n572), .ZN(n573) );
  XNOR2_X1 U639 ( .A(n574), .B(n573), .ZN(n575) );
  XNOR2_X1 U640 ( .A(G211GAT), .B(n575), .ZN(G1354GAT) );
  XOR2_X1 U641 ( .A(KEYINPUT126), .B(KEYINPUT62), .Z(n577) );
  XNOR2_X1 U642 ( .A(G218GAT), .B(KEYINPUT127), .ZN(n576) );
  XNOR2_X1 U643 ( .A(n577), .B(n576), .ZN(n582) );
  INV_X1 U644 ( .A(n578), .ZN(n579) );
  NOR2_X1 U645 ( .A1(n580), .A2(n579), .ZN(n581) );
  XOR2_X1 U646 ( .A(n582), .B(n581), .Z(G1355GAT) );
endmodule

