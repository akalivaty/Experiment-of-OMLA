//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 0 0 1 0 1 1 0 0 0 1 0 1 1 0 0 0 0 0 1 1 0 0 0 1 1 1 0 1 0 0 0 0 0 1 0 0 1 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 0 0 1 0 0 1 0 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:16:09 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n666, new_n667, new_n668, new_n669, new_n670, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n679, new_n680,
    new_n681, new_n682, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n726, new_n727, new_n728, new_n729, new_n730, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n738, new_n739, new_n740,
    new_n741, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n751, new_n752, new_n753, new_n754, new_n755, new_n757,
    new_n758, new_n759, new_n761, new_n762, new_n764, new_n765, new_n766,
    new_n767, new_n768, new_n769, new_n770, new_n771, new_n772, new_n773,
    new_n774, new_n775, new_n776, new_n777, new_n778, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n797, new_n798, new_n799, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n867, new_n868, new_n870, new_n871,
    new_n872, new_n873, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n933, new_n934, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n957, new_n958, new_n959, new_n961, new_n962,
    new_n963, new_n964, new_n965, new_n966, new_n967, new_n968, new_n969,
    new_n970, new_n971, new_n972, new_n973, new_n974, new_n975, new_n976,
    new_n977, new_n979, new_n980, new_n981, new_n982, new_n983, new_n984,
    new_n985, new_n987, new_n988, new_n989, new_n990, new_n991, new_n992,
    new_n993, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1009, new_n1010, new_n1011;
  XNOR2_X1  g000(.A(G113gat), .B(G141gat), .ZN(new_n202));
  XNOR2_X1  g001(.A(new_n202), .B(G197gat), .ZN(new_n203));
  XOR2_X1   g002(.A(KEYINPUT11), .B(G169gat), .Z(new_n204));
  XNOR2_X1  g003(.A(new_n203), .B(new_n204), .ZN(new_n205));
  XOR2_X1   g004(.A(new_n205), .B(KEYINPUT12), .Z(new_n206));
  INV_X1    g005(.A(new_n206), .ZN(new_n207));
  NAND2_X1  g006(.A1(G229gat), .A2(G233gat), .ZN(new_n208));
  XNOR2_X1  g007(.A(G15gat), .B(G22gat), .ZN(new_n209));
  NOR2_X1   g008(.A1(new_n209), .A2(G1gat), .ZN(new_n210));
  INV_X1    g009(.A(new_n210), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n211), .A2(KEYINPUT82), .ZN(new_n212));
  INV_X1    g011(.A(KEYINPUT82), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n210), .A2(new_n213), .ZN(new_n214));
  INV_X1    g013(.A(KEYINPUT16), .ZN(new_n215));
  OAI21_X1  g014(.A(new_n209), .B1(new_n215), .B2(G1gat), .ZN(new_n216));
  NAND3_X1  g015(.A1(new_n212), .A2(new_n214), .A3(new_n216), .ZN(new_n217));
  INV_X1    g016(.A(KEYINPUT83), .ZN(new_n218));
  INV_X1    g017(.A(G8gat), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n216), .A2(new_n219), .ZN(new_n220));
  OAI21_X1  g019(.A(new_n218), .B1(new_n220), .B2(new_n210), .ZN(new_n221));
  NAND4_X1  g020(.A1(new_n211), .A2(KEYINPUT83), .A3(new_n219), .A4(new_n216), .ZN(new_n222));
  AOI22_X1  g021(.A1(new_n217), .A2(G8gat), .B1(new_n221), .B2(new_n222), .ZN(new_n223));
  INV_X1    g022(.A(KEYINPUT17), .ZN(new_n224));
  XNOR2_X1  g023(.A(G43gat), .B(G50gat), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n225), .A2(KEYINPUT15), .ZN(new_n226));
  INV_X1    g025(.A(new_n226), .ZN(new_n227));
  XNOR2_X1  g026(.A(KEYINPUT79), .B(G29gat), .ZN(new_n228));
  XNOR2_X1  g027(.A(KEYINPUT80), .B(G36gat), .ZN(new_n229));
  NOR2_X1   g028(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  NOR2_X1   g029(.A1(G29gat), .A2(G36gat), .ZN(new_n231));
  XNOR2_X1  g030(.A(new_n231), .B(KEYINPUT14), .ZN(new_n232));
  OAI21_X1  g031(.A(new_n227), .B1(new_n230), .B2(new_n232), .ZN(new_n233));
  INV_X1    g032(.A(KEYINPUT81), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n230), .A2(new_n234), .ZN(new_n235));
  OAI21_X1  g034(.A(KEYINPUT81), .B1(new_n228), .B2(new_n229), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n235), .A2(new_n236), .ZN(new_n237));
  INV_X1    g036(.A(new_n232), .ZN(new_n238));
  OR2_X1    g037(.A1(new_n225), .A2(KEYINPUT15), .ZN(new_n239));
  NAND3_X1  g038(.A1(new_n238), .A2(new_n226), .A3(new_n239), .ZN(new_n240));
  OAI211_X1 g039(.A(new_n224), .B(new_n233), .C1(new_n237), .C2(new_n240), .ZN(new_n241));
  INV_X1    g040(.A(new_n241), .ZN(new_n242));
  NOR2_X1   g041(.A1(new_n227), .A2(new_n232), .ZN(new_n243));
  NAND4_X1  g042(.A1(new_n243), .A2(new_n239), .A3(new_n236), .A4(new_n235), .ZN(new_n244));
  AOI21_X1  g043(.A(new_n224), .B1(new_n244), .B2(new_n233), .ZN(new_n245));
  OAI21_X1  g044(.A(new_n223), .B1(new_n242), .B2(new_n245), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n221), .A2(new_n222), .ZN(new_n247));
  INV_X1    g046(.A(new_n214), .ZN(new_n248));
  OAI21_X1  g047(.A(new_n216), .B1(new_n210), .B2(new_n213), .ZN(new_n249));
  OAI21_X1  g048(.A(G8gat), .B1(new_n248), .B2(new_n249), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n247), .A2(new_n250), .ZN(new_n251));
  INV_X1    g050(.A(KEYINPUT84), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n244), .A2(new_n233), .ZN(new_n253));
  AND3_X1   g052(.A1(new_n251), .A2(new_n252), .A3(new_n253), .ZN(new_n254));
  AOI21_X1  g053(.A(new_n252), .B1(new_n251), .B2(new_n253), .ZN(new_n255));
  OAI211_X1 g054(.A(new_n208), .B(new_n246), .C1(new_n254), .C2(new_n255), .ZN(new_n256));
  NAND2_X1  g055(.A1(new_n256), .A2(KEYINPUT85), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n257), .A2(KEYINPUT18), .ZN(new_n258));
  INV_X1    g057(.A(KEYINPUT18), .ZN(new_n259));
  NAND3_X1  g058(.A1(new_n256), .A2(KEYINPUT85), .A3(new_n259), .ZN(new_n260));
  XOR2_X1   g059(.A(new_n208), .B(KEYINPUT13), .Z(new_n261));
  INV_X1    g060(.A(new_n261), .ZN(new_n262));
  INV_X1    g061(.A(new_n233), .ZN(new_n263));
  INV_X1    g062(.A(new_n237), .ZN(new_n264));
  INV_X1    g063(.A(new_n240), .ZN(new_n265));
  AOI21_X1  g064(.A(new_n263), .B1(new_n264), .B2(new_n265), .ZN(new_n266));
  OAI21_X1  g065(.A(KEYINPUT84), .B1(new_n223), .B2(new_n266), .ZN(new_n267));
  NAND3_X1  g066(.A1(new_n251), .A2(new_n252), .A3(new_n253), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n223), .A2(new_n266), .ZN(new_n270));
  AOI21_X1  g069(.A(new_n262), .B1(new_n269), .B2(new_n270), .ZN(new_n271));
  INV_X1    g070(.A(new_n271), .ZN(new_n272));
  AND4_X1   g071(.A1(new_n207), .A2(new_n258), .A3(new_n260), .A4(new_n272), .ZN(new_n273));
  AOI21_X1  g072(.A(new_n271), .B1(new_n257), .B2(KEYINPUT18), .ZN(new_n274));
  AOI21_X1  g073(.A(new_n207), .B1(new_n274), .B2(new_n260), .ZN(new_n275));
  NOR2_X1   g074(.A1(new_n273), .A2(new_n275), .ZN(new_n276));
  XNOR2_X1  g075(.A(G78gat), .B(G106gat), .ZN(new_n277));
  XNOR2_X1  g076(.A(KEYINPUT31), .B(G50gat), .ZN(new_n278));
  XOR2_X1   g077(.A(new_n277), .B(new_n278), .Z(new_n279));
  XNOR2_X1  g078(.A(new_n279), .B(KEYINPUT75), .ZN(new_n280));
  XNOR2_X1  g079(.A(KEYINPUT76), .B(G22gat), .ZN(new_n281));
  INV_X1    g080(.A(G141gat), .ZN(new_n282));
  INV_X1    g081(.A(G148gat), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  INV_X1    g083(.A(KEYINPUT2), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n285), .A2(KEYINPUT72), .ZN(new_n286));
  INV_X1    g085(.A(KEYINPUT72), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n287), .A2(KEYINPUT2), .ZN(new_n288));
  NAND2_X1  g087(.A1(G141gat), .A2(G148gat), .ZN(new_n289));
  NAND4_X1  g088(.A1(new_n284), .A2(new_n286), .A3(new_n288), .A4(new_n289), .ZN(new_n290));
  XOR2_X1   g089(.A(G155gat), .B(G162gat), .Z(new_n291));
  NAND2_X1  g090(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  XNOR2_X1  g091(.A(G155gat), .B(G162gat), .ZN(new_n293));
  INV_X1    g092(.A(G155gat), .ZN(new_n294));
  INV_X1    g093(.A(G162gat), .ZN(new_n295));
  OAI21_X1  g094(.A(KEYINPUT2), .B1(new_n294), .B2(new_n295), .ZN(new_n296));
  NAND4_X1  g095(.A1(new_n293), .A2(new_n284), .A3(new_n296), .A4(new_n289), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n292), .A2(new_n297), .ZN(new_n298));
  INV_X1    g097(.A(new_n298), .ZN(new_n299));
  XNOR2_X1  g098(.A(KEYINPUT73), .B(KEYINPUT3), .ZN(new_n300));
  NOR2_X1   g099(.A1(new_n299), .A2(new_n300), .ZN(new_n301));
  INV_X1    g100(.A(KEYINPUT22), .ZN(new_n302));
  AOI22_X1  g101(.A1(new_n302), .A2(KEYINPUT69), .B1(G211gat), .B2(G218gat), .ZN(new_n303));
  OAI21_X1  g102(.A(new_n303), .B1(KEYINPUT69), .B2(new_n302), .ZN(new_n304));
  XNOR2_X1  g103(.A(G197gat), .B(G204gat), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  XOR2_X1   g105(.A(G211gat), .B(G218gat), .Z(new_n307));
  NAND2_X1  g106(.A1(new_n306), .A2(new_n307), .ZN(new_n308));
  INV_X1    g107(.A(new_n307), .ZN(new_n309));
  NAND3_X1  g108(.A1(new_n309), .A2(new_n304), .A3(new_n305), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n308), .A2(new_n310), .ZN(new_n311));
  NOR2_X1   g110(.A1(new_n299), .A2(KEYINPUT29), .ZN(new_n312));
  AOI21_X1  g111(.A(new_n301), .B1(new_n311), .B2(new_n312), .ZN(new_n313));
  INV_X1    g112(.A(new_n311), .ZN(new_n314));
  NAND3_X1  g113(.A1(new_n292), .A2(new_n297), .A3(new_n300), .ZN(new_n315));
  INV_X1    g114(.A(KEYINPUT29), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n315), .A2(new_n316), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n314), .A2(new_n317), .ZN(new_n318));
  AOI22_X1  g117(.A1(new_n313), .A2(new_n318), .B1(G228gat), .B2(G233gat), .ZN(new_n319));
  INV_X1    g118(.A(new_n319), .ZN(new_n320));
  INV_X1    g119(.A(KEYINPUT70), .ZN(new_n321));
  NOR2_X1   g120(.A1(new_n311), .A2(new_n321), .ZN(new_n322));
  AOI21_X1  g121(.A(KEYINPUT70), .B1(new_n308), .B2(new_n310), .ZN(new_n323));
  OAI21_X1  g122(.A(new_n317), .B1(new_n322), .B2(new_n323), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n312), .A2(new_n311), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n298), .A2(KEYINPUT3), .ZN(new_n326));
  AND3_X1   g125(.A1(new_n326), .A2(G228gat), .A3(G233gat), .ZN(new_n327));
  NAND3_X1  g126(.A1(new_n324), .A2(new_n325), .A3(new_n327), .ZN(new_n328));
  AOI21_X1  g127(.A(new_n281), .B1(new_n320), .B2(new_n328), .ZN(new_n329));
  INV_X1    g128(.A(new_n328), .ZN(new_n330));
  INV_X1    g129(.A(new_n281), .ZN(new_n331));
  NOR3_X1   g130(.A1(new_n330), .A2(new_n319), .A3(new_n331), .ZN(new_n332));
  OAI21_X1  g131(.A(new_n280), .B1(new_n329), .B2(new_n332), .ZN(new_n333));
  OAI21_X1  g132(.A(G22gat), .B1(new_n330), .B2(new_n319), .ZN(new_n334));
  NAND3_X1  g133(.A1(new_n320), .A2(new_n281), .A3(new_n328), .ZN(new_n335));
  INV_X1    g134(.A(new_n279), .ZN(new_n336));
  NAND3_X1  g135(.A1(new_n334), .A2(new_n335), .A3(new_n336), .ZN(new_n337));
  AND2_X1   g136(.A1(new_n333), .A2(new_n337), .ZN(new_n338));
  XNOR2_X1  g137(.A(G8gat), .B(G36gat), .ZN(new_n339));
  XNOR2_X1  g138(.A(G64gat), .B(G92gat), .ZN(new_n340));
  XOR2_X1   g139(.A(new_n339), .B(new_n340), .Z(new_n341));
  INV_X1    g140(.A(new_n341), .ZN(new_n342));
  NAND2_X1  g141(.A1(G226gat), .A2(G233gat), .ZN(new_n343));
  INV_X1    g142(.A(new_n343), .ZN(new_n344));
  OR2_X1    g143(.A1(G169gat), .A2(G176gat), .ZN(new_n345));
  INV_X1    g144(.A(KEYINPUT26), .ZN(new_n346));
  NAND2_X1  g145(.A1(G169gat), .A2(G176gat), .ZN(new_n347));
  NAND3_X1  g146(.A1(new_n345), .A2(new_n346), .A3(new_n347), .ZN(new_n348));
  NAND2_X1  g147(.A1(G183gat), .A2(G190gat), .ZN(new_n349));
  NOR2_X1   g148(.A1(G169gat), .A2(G176gat), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n350), .A2(KEYINPUT26), .ZN(new_n351));
  NAND3_X1  g150(.A1(new_n348), .A2(new_n349), .A3(new_n351), .ZN(new_n352));
  XNOR2_X1  g151(.A(KEYINPUT27), .B(G183gat), .ZN(new_n353));
  INV_X1    g152(.A(G190gat), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  INV_X1    g154(.A(KEYINPUT28), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n355), .A2(new_n356), .ZN(new_n357));
  NAND3_X1  g156(.A1(new_n353), .A2(KEYINPUT28), .A3(new_n354), .ZN(new_n358));
  AOI21_X1  g157(.A(new_n352), .B1(new_n357), .B2(new_n358), .ZN(new_n359));
  INV_X1    g158(.A(new_n359), .ZN(new_n360));
  INV_X1    g159(.A(KEYINPUT23), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n345), .A2(new_n361), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n350), .A2(KEYINPUT23), .ZN(new_n363));
  NAND3_X1  g162(.A1(new_n362), .A2(new_n363), .A3(new_n347), .ZN(new_n364));
  NOR2_X1   g163(.A1(G183gat), .A2(G190gat), .ZN(new_n365));
  AND2_X1   g164(.A1(KEYINPUT24), .A2(G183gat), .ZN(new_n366));
  AOI21_X1  g165(.A(new_n365), .B1(new_n366), .B2(G190gat), .ZN(new_n367));
  AOI21_X1  g166(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n368));
  INV_X1    g167(.A(KEYINPUT65), .ZN(new_n369));
  NOR2_X1   g168(.A1(new_n368), .A2(new_n369), .ZN(new_n370));
  INV_X1    g169(.A(KEYINPUT24), .ZN(new_n371));
  AND3_X1   g170(.A1(new_n349), .A2(new_n369), .A3(new_n371), .ZN(new_n372));
  OAI21_X1  g171(.A(new_n367), .B1(new_n370), .B2(new_n372), .ZN(new_n373));
  AOI21_X1  g172(.A(new_n364), .B1(new_n373), .B2(KEYINPUT66), .ZN(new_n374));
  INV_X1    g173(.A(KEYINPUT66), .ZN(new_n375));
  OAI211_X1 g174(.A(new_n375), .B(new_n367), .C1(new_n370), .C2(new_n372), .ZN(new_n376));
  AOI21_X1  g175(.A(KEYINPUT25), .B1(new_n374), .B2(new_n376), .ZN(new_n377));
  NAND3_X1  g176(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n378));
  OAI21_X1  g177(.A(new_n378), .B1(G183gat), .B2(G190gat), .ZN(new_n379));
  NOR2_X1   g178(.A1(new_n379), .A2(new_n368), .ZN(new_n380));
  INV_X1    g179(.A(KEYINPUT25), .ZN(new_n381));
  NOR3_X1   g180(.A1(new_n364), .A2(new_n380), .A3(new_n381), .ZN(new_n382));
  OAI21_X1  g181(.A(new_n360), .B1(new_n377), .B2(new_n382), .ZN(new_n383));
  AOI21_X1  g182(.A(new_n344), .B1(new_n383), .B2(new_n316), .ZN(new_n384));
  AND3_X1   g183(.A1(new_n362), .A2(new_n363), .A3(new_n347), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n349), .A2(new_n371), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n386), .A2(KEYINPUT65), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n368), .A2(new_n369), .ZN(new_n388));
  AOI21_X1  g187(.A(new_n379), .B1(new_n387), .B2(new_n388), .ZN(new_n389));
  OAI21_X1  g188(.A(new_n385), .B1(new_n389), .B2(new_n375), .ZN(new_n390));
  INV_X1    g189(.A(new_n376), .ZN(new_n391));
  OAI21_X1  g190(.A(new_n381), .B1(new_n390), .B2(new_n391), .ZN(new_n392));
  INV_X1    g191(.A(new_n382), .ZN(new_n393));
  AOI21_X1  g192(.A(new_n359), .B1(new_n392), .B2(new_n393), .ZN(new_n394));
  XOR2_X1   g193(.A(new_n343), .B(KEYINPUT71), .Z(new_n395));
  INV_X1    g194(.A(new_n395), .ZN(new_n396));
  NOR2_X1   g195(.A1(new_n394), .A2(new_n396), .ZN(new_n397));
  NOR3_X1   g196(.A1(new_n384), .A2(new_n397), .A3(new_n314), .ZN(new_n398));
  NOR2_X1   g197(.A1(new_n322), .A2(new_n323), .ZN(new_n399));
  OAI21_X1  g198(.A(new_n396), .B1(new_n394), .B2(KEYINPUT29), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n383), .A2(new_n344), .ZN(new_n401));
  AOI21_X1  g200(.A(new_n399), .B1(new_n400), .B2(new_n401), .ZN(new_n402));
  OAI21_X1  g201(.A(new_n342), .B1(new_n398), .B2(new_n402), .ZN(new_n403));
  INV_X1    g202(.A(new_n399), .ZN(new_n404));
  AOI21_X1  g203(.A(new_n395), .B1(new_n383), .B2(new_n316), .ZN(new_n405));
  NOR2_X1   g204(.A1(new_n394), .A2(new_n343), .ZN(new_n406));
  OAI21_X1  g205(.A(new_n404), .B1(new_n405), .B2(new_n406), .ZN(new_n407));
  OAI21_X1  g206(.A(new_n343), .B1(new_n394), .B2(KEYINPUT29), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n383), .A2(new_n395), .ZN(new_n409));
  NAND3_X1  g208(.A1(new_n408), .A2(new_n311), .A3(new_n409), .ZN(new_n410));
  NAND3_X1  g209(.A1(new_n407), .A2(new_n410), .A3(new_n341), .ZN(new_n411));
  NAND3_X1  g210(.A1(new_n403), .A2(KEYINPUT30), .A3(new_n411), .ZN(new_n412));
  INV_X1    g211(.A(KEYINPUT30), .ZN(new_n413));
  NAND4_X1  g212(.A1(new_n407), .A2(new_n410), .A3(new_n413), .A4(new_n341), .ZN(new_n414));
  AND2_X1   g213(.A1(new_n412), .A2(new_n414), .ZN(new_n415));
  INV_X1    g214(.A(G113gat), .ZN(new_n416));
  INV_X1    g215(.A(G120gat), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  INV_X1    g217(.A(KEYINPUT1), .ZN(new_n419));
  NAND2_X1  g218(.A1(G113gat), .A2(G120gat), .ZN(new_n420));
  NAND3_X1  g219(.A1(new_n418), .A2(new_n419), .A3(new_n420), .ZN(new_n421));
  INV_X1    g220(.A(G127gat), .ZN(new_n422));
  INV_X1    g221(.A(G134gat), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  XNOR2_X1  g223(.A(KEYINPUT67), .B(G134gat), .ZN(new_n425));
  OAI211_X1 g224(.A(new_n421), .B(new_n424), .C1(new_n422), .C2(new_n425), .ZN(new_n426));
  AND2_X1   g225(.A1(KEYINPUT68), .A2(G120gat), .ZN(new_n427));
  NOR2_X1   g226(.A1(KEYINPUT68), .A2(G120gat), .ZN(new_n428));
  OAI21_X1  g227(.A(G113gat), .B1(new_n427), .B2(new_n428), .ZN(new_n429));
  OAI21_X1  g228(.A(new_n419), .B1(G113gat), .B2(G120gat), .ZN(new_n430));
  INV_X1    g229(.A(new_n430), .ZN(new_n431));
  NAND2_X1  g230(.A1(G127gat), .A2(G134gat), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n424), .A2(new_n432), .ZN(new_n433));
  NAND3_X1  g232(.A1(new_n429), .A2(new_n431), .A3(new_n433), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n426), .A2(new_n434), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n435), .A2(new_n298), .ZN(new_n436));
  NAND4_X1  g235(.A1(new_n426), .A2(new_n292), .A3(new_n297), .A4(new_n434), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n436), .A2(new_n437), .ZN(new_n438));
  NAND2_X1  g237(.A1(G225gat), .A2(G233gat), .ZN(new_n439));
  INV_X1    g238(.A(new_n439), .ZN(new_n440));
  OAI21_X1  g239(.A(KEYINPUT39), .B1(new_n438), .B2(new_n440), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n441), .A2(KEYINPUT77), .ZN(new_n442));
  INV_X1    g241(.A(KEYINPUT77), .ZN(new_n443));
  OAI211_X1 g242(.A(new_n443), .B(KEYINPUT39), .C1(new_n438), .C2(new_n440), .ZN(new_n444));
  XNOR2_X1  g243(.A(new_n437), .B(KEYINPUT4), .ZN(new_n445));
  NAND3_X1  g244(.A1(new_n326), .A2(new_n315), .A3(new_n435), .ZN(new_n446));
  AND2_X1   g245(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  OAI211_X1 g246(.A(new_n442), .B(new_n444), .C1(new_n447), .C2(new_n439), .ZN(new_n448));
  XOR2_X1   g247(.A(G1gat), .B(G29gat), .Z(new_n449));
  XNOR2_X1  g248(.A(new_n449), .B(KEYINPUT0), .ZN(new_n450));
  XNOR2_X1  g249(.A(G57gat), .B(G85gat), .ZN(new_n451));
  XNOR2_X1  g250(.A(new_n450), .B(new_n451), .ZN(new_n452));
  INV_X1    g251(.A(new_n452), .ZN(new_n453));
  AOI21_X1  g252(.A(new_n439), .B1(new_n445), .B2(new_n446), .ZN(new_n454));
  INV_X1    g253(.A(KEYINPUT39), .ZN(new_n455));
  AOI21_X1  g254(.A(new_n453), .B1(new_n454), .B2(new_n455), .ZN(new_n456));
  AND3_X1   g255(.A1(new_n448), .A2(KEYINPUT40), .A3(new_n456), .ZN(new_n457));
  AOI21_X1  g256(.A(KEYINPUT40), .B1(new_n448), .B2(new_n456), .ZN(new_n458));
  INV_X1    g257(.A(KEYINPUT74), .ZN(new_n459));
  INV_X1    g258(.A(new_n424), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n423), .A2(KEYINPUT67), .ZN(new_n461));
  INV_X1    g260(.A(KEYINPUT67), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n462), .A2(G134gat), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n461), .A2(new_n463), .ZN(new_n464));
  AOI21_X1  g263(.A(new_n460), .B1(new_n464), .B2(G127gat), .ZN(new_n465));
  AOI21_X1  g264(.A(new_n430), .B1(new_n424), .B2(new_n432), .ZN(new_n466));
  AOI22_X1  g265(.A1(new_n465), .A2(new_n421), .B1(new_n466), .B2(new_n429), .ZN(new_n467));
  NAND3_X1  g266(.A1(new_n299), .A2(new_n467), .A3(KEYINPUT4), .ZN(new_n468));
  INV_X1    g267(.A(KEYINPUT4), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n437), .A2(new_n469), .ZN(new_n470));
  NAND4_X1  g269(.A1(new_n446), .A2(new_n468), .A3(new_n439), .A4(new_n470), .ZN(new_n471));
  OAI21_X1  g270(.A(new_n459), .B1(new_n471), .B2(KEYINPUT5), .ZN(new_n472));
  INV_X1    g271(.A(KEYINPUT5), .ZN(new_n473));
  AOI21_X1  g272(.A(new_n473), .B1(new_n438), .B2(new_n440), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n474), .A2(new_n471), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n472), .A2(new_n475), .ZN(new_n476));
  NAND3_X1  g275(.A1(new_n474), .A2(new_n471), .A3(new_n459), .ZN(new_n477));
  AOI21_X1  g276(.A(new_n452), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  NOR3_X1   g277(.A1(new_n457), .A2(new_n458), .A3(new_n478), .ZN(new_n479));
  AOI21_X1  g278(.A(new_n338), .B1(new_n415), .B2(new_n479), .ZN(new_n480));
  NAND4_X1  g279(.A1(new_n445), .A2(new_n473), .A3(new_n439), .A4(new_n446), .ZN(new_n481));
  AOI22_X1  g280(.A1(new_n481), .A2(new_n459), .B1(new_n471), .B2(new_n474), .ZN(new_n482));
  INV_X1    g281(.A(new_n477), .ZN(new_n483));
  OAI21_X1  g282(.A(new_n453), .B1(new_n482), .B2(new_n483), .ZN(new_n484));
  INV_X1    g283(.A(KEYINPUT6), .ZN(new_n485));
  NAND3_X1  g284(.A1(new_n476), .A2(new_n452), .A3(new_n477), .ZN(new_n486));
  NAND4_X1  g285(.A1(new_n484), .A2(KEYINPUT78), .A3(new_n485), .A4(new_n486), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n478), .A2(KEYINPUT6), .ZN(new_n488));
  AND2_X1   g287(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  INV_X1    g288(.A(new_n411), .ZN(new_n490));
  INV_X1    g289(.A(KEYINPUT37), .ZN(new_n491));
  NOR2_X1   g290(.A1(new_n341), .A2(new_n491), .ZN(new_n492));
  INV_X1    g291(.A(new_n492), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n403), .A2(new_n493), .ZN(new_n494));
  OAI21_X1  g293(.A(new_n314), .B1(new_n384), .B2(new_n397), .ZN(new_n495));
  NAND3_X1  g294(.A1(new_n400), .A2(new_n401), .A3(new_n399), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  AOI21_X1  g296(.A(KEYINPUT38), .B1(new_n497), .B2(KEYINPUT37), .ZN(new_n498));
  AOI21_X1  g297(.A(new_n490), .B1(new_n494), .B2(new_n498), .ZN(new_n499));
  NAND3_X1  g298(.A1(new_n484), .A2(new_n485), .A3(new_n486), .ZN(new_n500));
  INV_X1    g299(.A(KEYINPUT78), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n407), .A2(new_n410), .ZN(new_n503));
  AOI21_X1  g302(.A(new_n492), .B1(new_n503), .B2(new_n342), .ZN(new_n504));
  AOI21_X1  g303(.A(new_n491), .B1(new_n407), .B2(new_n410), .ZN(new_n505));
  OAI21_X1  g304(.A(KEYINPUT38), .B1(new_n504), .B2(new_n505), .ZN(new_n506));
  NAND4_X1  g305(.A1(new_n489), .A2(new_n499), .A3(new_n502), .A4(new_n506), .ZN(new_n507));
  INV_X1    g306(.A(KEYINPUT36), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n373), .A2(KEYINPUT66), .ZN(new_n509));
  NAND3_X1  g308(.A1(new_n509), .A2(new_n376), .A3(new_n385), .ZN(new_n510));
  AOI21_X1  g309(.A(new_n382), .B1(new_n510), .B2(new_n381), .ZN(new_n511));
  OAI21_X1  g310(.A(new_n467), .B1(new_n511), .B2(new_n359), .ZN(new_n512));
  NAND2_X1  g311(.A1(G227gat), .A2(G233gat), .ZN(new_n513));
  XNOR2_X1  g312(.A(new_n513), .B(KEYINPUT64), .ZN(new_n514));
  OAI211_X1 g313(.A(new_n360), .B(new_n435), .C1(new_n377), .C2(new_n382), .ZN(new_n515));
  NAND3_X1  g314(.A1(new_n512), .A2(new_n514), .A3(new_n515), .ZN(new_n516));
  INV_X1    g315(.A(KEYINPUT33), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  XOR2_X1   g317(.A(G15gat), .B(G43gat), .Z(new_n519));
  XNOR2_X1  g318(.A(G71gat), .B(G99gat), .ZN(new_n520));
  XNOR2_X1  g319(.A(new_n519), .B(new_n520), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n518), .A2(new_n521), .ZN(new_n522));
  AND2_X1   g321(.A1(new_n512), .A2(new_n515), .ZN(new_n523));
  OAI21_X1  g322(.A(KEYINPUT34), .B1(new_n523), .B2(new_n514), .ZN(new_n524));
  AOI21_X1  g323(.A(new_n514), .B1(new_n512), .B2(new_n515), .ZN(new_n525));
  INV_X1    g324(.A(KEYINPUT34), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  NAND3_X1  g326(.A1(new_n522), .A2(new_n524), .A3(new_n527), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n516), .A2(KEYINPUT32), .ZN(new_n529));
  INV_X1    g328(.A(new_n529), .ZN(new_n530));
  INV_X1    g329(.A(new_n521), .ZN(new_n531));
  AOI21_X1  g330(.A(new_n531), .B1(new_n516), .B2(new_n517), .ZN(new_n532));
  NOR2_X1   g331(.A1(new_n525), .A2(new_n526), .ZN(new_n533));
  AOI211_X1 g332(.A(KEYINPUT34), .B(new_n514), .C1(new_n512), .C2(new_n515), .ZN(new_n534));
  OAI21_X1  g333(.A(new_n532), .B1(new_n533), .B2(new_n534), .ZN(new_n535));
  AND3_X1   g334(.A1(new_n528), .A2(new_n530), .A3(new_n535), .ZN(new_n536));
  AOI21_X1  g335(.A(new_n530), .B1(new_n528), .B2(new_n535), .ZN(new_n537));
  OAI21_X1  g336(.A(new_n508), .B1(new_n536), .B2(new_n537), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n528), .A2(new_n535), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n539), .A2(new_n529), .ZN(new_n540));
  NAND3_X1  g339(.A1(new_n528), .A2(new_n530), .A3(new_n535), .ZN(new_n541));
  NAND3_X1  g340(.A1(new_n540), .A2(KEYINPUT36), .A3(new_n541), .ZN(new_n542));
  AOI22_X1  g341(.A1(new_n480), .A2(new_n507), .B1(new_n538), .B2(new_n542), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n333), .A2(new_n337), .ZN(new_n544));
  NAND2_X1  g343(.A1(new_n412), .A2(new_n414), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n500), .A2(new_n488), .ZN(new_n546));
  AOI21_X1  g345(.A(new_n544), .B1(new_n545), .B2(new_n546), .ZN(new_n547));
  INV_X1    g346(.A(new_n547), .ZN(new_n548));
  NAND2_X1  g347(.A1(new_n543), .A2(new_n548), .ZN(new_n549));
  AND4_X1   g348(.A1(new_n545), .A2(new_n540), .A3(new_n544), .A4(new_n541), .ZN(new_n550));
  AOI21_X1  g349(.A(KEYINPUT35), .B1(new_n489), .B2(new_n502), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  AOI22_X1  g351(.A1(new_n412), .A2(new_n414), .B1(new_n500), .B2(new_n488), .ZN(new_n553));
  NAND4_X1  g352(.A1(new_n553), .A2(new_n544), .A3(new_n540), .A4(new_n541), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n554), .A2(KEYINPUT35), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n552), .A2(new_n555), .ZN(new_n556));
  AOI21_X1  g355(.A(new_n276), .B1(new_n549), .B2(new_n556), .ZN(new_n557));
  INV_X1    g356(.A(KEYINPUT96), .ZN(new_n558));
  XOR2_X1   g357(.A(G71gat), .B(G78gat), .Z(new_n559));
  NAND2_X1  g358(.A1(G71gat), .A2(G78gat), .ZN(new_n560));
  INV_X1    g359(.A(KEYINPUT9), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  INV_X1    g361(.A(G57gat), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n563), .A2(G64gat), .ZN(new_n564));
  INV_X1    g363(.A(G64gat), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n565), .A2(G57gat), .ZN(new_n566));
  AND2_X1   g365(.A1(new_n564), .A2(new_n566), .ZN(new_n567));
  INV_X1    g366(.A(KEYINPUT86), .ZN(new_n568));
  OAI21_X1  g367(.A(new_n562), .B1(new_n567), .B2(new_n568), .ZN(new_n569));
  AND3_X1   g368(.A1(new_n564), .A2(new_n566), .A3(new_n568), .ZN(new_n570));
  OAI21_X1  g369(.A(new_n559), .B1(new_n569), .B2(new_n570), .ZN(new_n571));
  OAI21_X1  g370(.A(KEYINPUT87), .B1(new_n563), .B2(G64gat), .ZN(new_n572));
  INV_X1    g371(.A(KEYINPUT87), .ZN(new_n573));
  NAND3_X1  g372(.A1(new_n573), .A2(new_n565), .A3(G57gat), .ZN(new_n574));
  NAND3_X1  g373(.A1(new_n572), .A2(new_n574), .A3(new_n564), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n575), .A2(KEYINPUT88), .ZN(new_n576));
  INV_X1    g375(.A(new_n559), .ZN(new_n577));
  INV_X1    g376(.A(KEYINPUT88), .ZN(new_n578));
  NAND4_X1  g377(.A1(new_n572), .A2(new_n574), .A3(new_n578), .A4(new_n564), .ZN(new_n579));
  NAND4_X1  g378(.A1(new_n576), .A2(new_n577), .A3(new_n562), .A4(new_n579), .ZN(new_n580));
  AOI21_X1  g379(.A(KEYINPUT21), .B1(new_n571), .B2(new_n580), .ZN(new_n581));
  NAND2_X1  g380(.A1(G231gat), .A2(G233gat), .ZN(new_n582));
  XNOR2_X1  g381(.A(new_n581), .B(new_n582), .ZN(new_n583));
  XNOR2_X1  g382(.A(new_n583), .B(G127gat), .ZN(new_n584));
  NAND2_X1  g383(.A1(new_n571), .A2(new_n580), .ZN(new_n585));
  NAND2_X1  g384(.A1(new_n585), .A2(KEYINPUT89), .ZN(new_n586));
  INV_X1    g385(.A(KEYINPUT89), .ZN(new_n587));
  NAND3_X1  g386(.A1(new_n571), .A2(new_n587), .A3(new_n580), .ZN(new_n588));
  NAND3_X1  g387(.A1(new_n586), .A2(KEYINPUT21), .A3(new_n588), .ZN(new_n589));
  NAND2_X1  g388(.A1(new_n589), .A2(new_n223), .ZN(new_n590));
  XNOR2_X1  g389(.A(new_n584), .B(new_n590), .ZN(new_n591));
  XNOR2_X1  g390(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n592));
  XNOR2_X1  g391(.A(new_n592), .B(new_n294), .ZN(new_n593));
  XNOR2_X1  g392(.A(G183gat), .B(G211gat), .ZN(new_n594));
  XOR2_X1   g393(.A(new_n593), .B(new_n594), .Z(new_n595));
  OR2_X1    g394(.A1(new_n591), .A2(new_n595), .ZN(new_n596));
  NAND2_X1  g395(.A1(new_n591), .A2(new_n595), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  XNOR2_X1  g397(.A(G190gat), .B(G218gat), .ZN(new_n599));
  XNOR2_X1  g398(.A(new_n599), .B(KEYINPUT93), .ZN(new_n600));
  INV_X1    g399(.A(new_n600), .ZN(new_n601));
  NAND3_X1  g400(.A1(KEYINPUT90), .A2(G85gat), .A3(G92gat), .ZN(new_n602));
  XNOR2_X1  g401(.A(new_n602), .B(KEYINPUT7), .ZN(new_n603));
  NAND2_X1  g402(.A1(G99gat), .A2(G106gat), .ZN(new_n604));
  INV_X1    g403(.A(G85gat), .ZN(new_n605));
  INV_X1    g404(.A(G92gat), .ZN(new_n606));
  AOI22_X1  g405(.A1(KEYINPUT8), .A2(new_n604), .B1(new_n605), .B2(new_n606), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n603), .A2(new_n607), .ZN(new_n608));
  XNOR2_X1  g407(.A(G99gat), .B(G106gat), .ZN(new_n609));
  INV_X1    g408(.A(new_n609), .ZN(new_n610));
  NAND2_X1  g409(.A1(new_n608), .A2(new_n610), .ZN(new_n611));
  NAND3_X1  g410(.A1(new_n603), .A2(new_n609), .A3(new_n607), .ZN(new_n612));
  NAND3_X1  g411(.A1(new_n611), .A2(KEYINPUT91), .A3(new_n612), .ZN(new_n613));
  AOI21_X1  g412(.A(new_n609), .B1(new_n603), .B2(new_n607), .ZN(new_n614));
  INV_X1    g413(.A(KEYINPUT91), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n613), .A2(new_n616), .ZN(new_n617));
  NAND2_X1  g416(.A1(G232gat), .A2(G233gat), .ZN(new_n618));
  INV_X1    g417(.A(new_n618), .ZN(new_n619));
  AOI22_X1  g418(.A1(new_n617), .A2(new_n253), .B1(KEYINPUT41), .B2(new_n619), .ZN(new_n620));
  INV_X1    g419(.A(KEYINPUT92), .ZN(new_n621));
  XNOR2_X1  g420(.A(new_n620), .B(new_n621), .ZN(new_n622));
  OAI211_X1 g421(.A(new_n616), .B(new_n613), .C1(new_n242), .C2(new_n245), .ZN(new_n623));
  AOI21_X1  g422(.A(new_n601), .B1(new_n622), .B2(new_n623), .ZN(new_n624));
  INV_X1    g423(.A(new_n624), .ZN(new_n625));
  NAND3_X1  g424(.A1(new_n622), .A2(new_n601), .A3(new_n623), .ZN(new_n626));
  NAND2_X1  g425(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  NOR2_X1   g426(.A1(new_n619), .A2(KEYINPUT41), .ZN(new_n628));
  XNOR2_X1  g427(.A(new_n628), .B(G134gat), .ZN(new_n629));
  XNOR2_X1  g428(.A(new_n629), .B(new_n295), .ZN(new_n630));
  INV_X1    g429(.A(KEYINPUT94), .ZN(new_n631));
  OAI21_X1  g430(.A(new_n630), .B1(new_n624), .B2(new_n631), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n627), .A2(new_n632), .ZN(new_n633));
  NAND4_X1  g432(.A1(new_n625), .A2(new_n631), .A3(new_n626), .A4(new_n630), .ZN(new_n634));
  NAND2_X1  g433(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n598), .A2(new_n635), .ZN(new_n636));
  NAND2_X1  g435(.A1(G230gat), .A2(G233gat), .ZN(new_n637));
  INV_X1    g436(.A(new_n637), .ZN(new_n638));
  NAND2_X1  g437(.A1(new_n611), .A2(new_n612), .ZN(new_n639));
  OAI21_X1  g438(.A(KEYINPUT95), .B1(new_n585), .B2(new_n639), .ZN(new_n640));
  NAND3_X1  g439(.A1(new_n585), .A2(new_n613), .A3(new_n616), .ZN(new_n641));
  AND3_X1   g440(.A1(new_n603), .A2(new_n609), .A3(new_n607), .ZN(new_n642));
  NOR2_X1   g441(.A1(new_n642), .A2(new_n614), .ZN(new_n643));
  INV_X1    g442(.A(KEYINPUT95), .ZN(new_n644));
  NAND4_X1  g443(.A1(new_n643), .A2(new_n644), .A3(new_n571), .A4(new_n580), .ZN(new_n645));
  INV_X1    g444(.A(KEYINPUT10), .ZN(new_n646));
  NAND4_X1  g445(.A1(new_n640), .A2(new_n641), .A3(new_n645), .A4(new_n646), .ZN(new_n647));
  NAND4_X1  g446(.A1(new_n586), .A2(new_n617), .A3(KEYINPUT10), .A4(new_n588), .ZN(new_n648));
  AOI21_X1  g447(.A(new_n638), .B1(new_n647), .B2(new_n648), .ZN(new_n649));
  NAND3_X1  g448(.A1(new_n640), .A2(new_n641), .A3(new_n645), .ZN(new_n650));
  AOI21_X1  g449(.A(new_n649), .B1(new_n638), .B2(new_n650), .ZN(new_n651));
  XNOR2_X1  g450(.A(G120gat), .B(G148gat), .ZN(new_n652));
  XNOR2_X1  g451(.A(G176gat), .B(G204gat), .ZN(new_n653));
  XOR2_X1   g452(.A(new_n652), .B(new_n653), .Z(new_n654));
  OR2_X1    g453(.A1(new_n651), .A2(new_n654), .ZN(new_n655));
  NAND2_X1  g454(.A1(new_n651), .A2(new_n654), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  NOR2_X1   g456(.A1(new_n636), .A2(new_n657), .ZN(new_n658));
  NAND3_X1  g457(.A1(new_n557), .A2(new_n558), .A3(new_n658), .ZN(new_n659));
  INV_X1    g458(.A(new_n659), .ZN(new_n660));
  AOI21_X1  g459(.A(new_n558), .B1(new_n557), .B2(new_n658), .ZN(new_n661));
  NOR2_X1   g460(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  NOR2_X1   g461(.A1(new_n662), .A2(new_n546), .ZN(new_n663));
  XNOR2_X1  g462(.A(KEYINPUT97), .B(G1gat), .ZN(new_n664));
  XNOR2_X1  g463(.A(new_n663), .B(new_n664), .ZN(G1324gat));
  OR2_X1    g464(.A1(new_n660), .A2(new_n661), .ZN(new_n666));
  AOI21_X1  g465(.A(new_n219), .B1(new_n666), .B2(new_n415), .ZN(new_n667));
  XNOR2_X1  g466(.A(KEYINPUT16), .B(G8gat), .ZN(new_n668));
  NOR3_X1   g467(.A1(new_n662), .A2(new_n545), .A3(new_n668), .ZN(new_n669));
  OAI21_X1  g468(.A(KEYINPUT42), .B1(new_n667), .B2(new_n669), .ZN(new_n670));
  OAI21_X1  g469(.A(new_n670), .B1(KEYINPUT42), .B2(new_n669), .ZN(G1325gat));
  INV_X1    g470(.A(G15gat), .ZN(new_n672));
  NOR2_X1   g471(.A1(new_n536), .A2(new_n537), .ZN(new_n673));
  NAND3_X1  g472(.A1(new_n666), .A2(new_n672), .A3(new_n673), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n538), .A2(new_n542), .ZN(new_n675));
  OAI21_X1  g474(.A(G15gat), .B1(new_n662), .B2(new_n675), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n674), .A2(new_n676), .ZN(new_n677));
  XOR2_X1   g476(.A(new_n677), .B(KEYINPUT98), .Z(G1326gat));
  OR3_X1    g477(.A1(new_n662), .A2(KEYINPUT99), .A3(new_n544), .ZN(new_n679));
  OAI21_X1  g478(.A(KEYINPUT99), .B1(new_n662), .B2(new_n544), .ZN(new_n680));
  NAND2_X1  g479(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  XNOR2_X1  g480(.A(KEYINPUT43), .B(G22gat), .ZN(new_n682));
  XNOR2_X1  g481(.A(new_n681), .B(new_n682), .ZN(G1327gat));
  NOR3_X1   g482(.A1(new_n598), .A2(new_n635), .A3(new_n657), .ZN(new_n684));
  NAND2_X1  g483(.A1(new_n557), .A2(new_n684), .ZN(new_n685));
  XOR2_X1   g484(.A(KEYINPUT79), .B(G29gat), .Z(new_n686));
  NOR3_X1   g485(.A1(new_n685), .A2(new_n546), .A3(new_n686), .ZN(new_n687));
  XOR2_X1   g486(.A(new_n687), .B(KEYINPUT45), .Z(new_n688));
  INV_X1    g487(.A(KEYINPUT44), .ZN(new_n689));
  INV_X1    g488(.A(KEYINPUT101), .ZN(new_n690));
  NOR2_X1   g489(.A1(new_n547), .A2(new_n690), .ZN(new_n691));
  NOR3_X1   g490(.A1(new_n553), .A2(KEYINPUT101), .A3(new_n544), .ZN(new_n692));
  NOR2_X1   g491(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  AOI22_X1  g492(.A1(new_n693), .A2(new_n543), .B1(new_n552), .B2(new_n555), .ZN(new_n694));
  OAI21_X1  g493(.A(new_n689), .B1(new_n694), .B2(new_n635), .ZN(new_n695));
  NOR2_X1   g494(.A1(new_n635), .A2(new_n689), .ZN(new_n696));
  NAND3_X1  g495(.A1(new_n479), .A2(new_n412), .A3(new_n414), .ZN(new_n697));
  NOR3_X1   g496(.A1(new_n405), .A2(new_n406), .A3(new_n404), .ZN(new_n698));
  AOI21_X1  g497(.A(new_n311), .B1(new_n408), .B2(new_n409), .ZN(new_n699));
  OAI21_X1  g498(.A(KEYINPUT37), .B1(new_n698), .B2(new_n699), .ZN(new_n700));
  INV_X1    g499(.A(KEYINPUT38), .ZN(new_n701));
  AOI21_X1  g500(.A(new_n341), .B1(new_n407), .B2(new_n410), .ZN(new_n702));
  OAI211_X1 g501(.A(new_n700), .B(new_n701), .C1(new_n702), .C2(new_n492), .ZN(new_n703));
  AOI21_X1  g502(.A(new_n505), .B1(new_n403), .B2(new_n493), .ZN(new_n704));
  OAI211_X1 g503(.A(new_n703), .B(new_n411), .C1(new_n704), .C2(new_n701), .ZN(new_n705));
  NAND3_X1  g504(.A1(new_n502), .A2(new_n488), .A3(new_n487), .ZN(new_n706));
  OAI211_X1 g505(.A(new_n544), .B(new_n697), .C1(new_n705), .C2(new_n706), .ZN(new_n707));
  AND3_X1   g506(.A1(new_n707), .A2(new_n548), .A3(new_n675), .ZN(new_n708));
  AOI22_X1  g507(.A1(new_n550), .A2(new_n551), .B1(new_n554), .B2(KEYINPUT35), .ZN(new_n709));
  OAI21_X1  g508(.A(new_n696), .B1(new_n708), .B2(new_n709), .ZN(new_n710));
  AND2_X1   g509(.A1(new_n695), .A2(new_n710), .ZN(new_n711));
  INV_X1    g510(.A(new_n546), .ZN(new_n712));
  INV_X1    g511(.A(new_n598), .ZN(new_n713));
  NAND2_X1  g512(.A1(new_n274), .A2(new_n260), .ZN(new_n714));
  NAND2_X1  g513(.A1(new_n714), .A2(new_n206), .ZN(new_n715));
  NAND3_X1  g514(.A1(new_n274), .A2(new_n207), .A3(new_n260), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  INV_X1    g516(.A(new_n657), .ZN(new_n718));
  NAND3_X1  g517(.A1(new_n713), .A2(new_n717), .A3(new_n718), .ZN(new_n719));
  XNOR2_X1  g518(.A(new_n719), .B(KEYINPUT100), .ZN(new_n720));
  NAND3_X1  g519(.A1(new_n711), .A2(new_n712), .A3(new_n720), .ZN(new_n721));
  INV_X1    g520(.A(KEYINPUT102), .ZN(new_n722));
  AND2_X1   g521(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  OAI21_X1  g522(.A(new_n686), .B1(new_n721), .B2(new_n722), .ZN(new_n724));
  OAI21_X1  g523(.A(new_n688), .B1(new_n723), .B2(new_n724), .ZN(G1328gat));
  XOR2_X1   g524(.A(KEYINPUT80), .B(G36gat), .Z(new_n726));
  NOR3_X1   g525(.A1(new_n685), .A2(new_n545), .A3(new_n726), .ZN(new_n727));
  XNOR2_X1  g526(.A(new_n727), .B(KEYINPUT46), .ZN(new_n728));
  NAND2_X1  g527(.A1(new_n711), .A2(new_n720), .ZN(new_n729));
  OAI21_X1  g528(.A(new_n726), .B1(new_n729), .B2(new_n545), .ZN(new_n730));
  NAND2_X1  g529(.A1(new_n728), .A2(new_n730), .ZN(G1329gat));
  INV_X1    g530(.A(new_n675), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n732), .A2(G43gat), .ZN(new_n733));
  INV_X1    g532(.A(new_n673), .ZN(new_n734));
  NOR2_X1   g533(.A1(new_n685), .A2(new_n734), .ZN(new_n735));
  OAI22_X1  g534(.A1(new_n729), .A2(new_n733), .B1(G43gat), .B2(new_n735), .ZN(new_n736));
  XNOR2_X1  g535(.A(new_n736), .B(KEYINPUT47), .ZN(G1330gat));
  OAI21_X1  g536(.A(G50gat), .B1(new_n729), .B2(new_n544), .ZN(new_n738));
  NOR2_X1   g537(.A1(new_n544), .A2(G50gat), .ZN(new_n739));
  XOR2_X1   g538(.A(new_n739), .B(KEYINPUT103), .Z(new_n740));
  OAI21_X1  g539(.A(new_n738), .B1(new_n685), .B2(new_n740), .ZN(new_n741));
  XOR2_X1   g540(.A(new_n741), .B(KEYINPUT48), .Z(G1331gat));
  NAND2_X1  g541(.A1(new_n547), .A2(new_n690), .ZN(new_n743));
  OAI21_X1  g542(.A(KEYINPUT101), .B1(new_n553), .B2(new_n544), .ZN(new_n744));
  NAND4_X1  g543(.A1(new_n707), .A2(new_n675), .A3(new_n743), .A4(new_n744), .ZN(new_n745));
  NAND2_X1  g544(.A1(new_n556), .A2(new_n745), .ZN(new_n746));
  NOR3_X1   g545(.A1(new_n636), .A2(new_n717), .A3(new_n718), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  NOR2_X1   g547(.A1(new_n748), .A2(new_n546), .ZN(new_n749));
  XNOR2_X1  g548(.A(new_n749), .B(new_n563), .ZN(G1332gat));
  INV_X1    g549(.A(new_n748), .ZN(new_n751));
  AOI21_X1  g550(.A(new_n545), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n752));
  XNOR2_X1  g551(.A(new_n752), .B(KEYINPUT104), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n751), .A2(new_n753), .ZN(new_n754));
  NOR2_X1   g553(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n755));
  XOR2_X1   g554(.A(new_n754), .B(new_n755), .Z(G1333gat));
  NOR3_X1   g555(.A1(new_n748), .A2(G71gat), .A3(new_n734), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n751), .A2(new_n732), .ZN(new_n758));
  AOI21_X1  g557(.A(new_n757), .B1(G71gat), .B2(new_n758), .ZN(new_n759));
  XNOR2_X1  g558(.A(new_n759), .B(KEYINPUT50), .ZN(G1334gat));
  NOR2_X1   g559(.A1(new_n748), .A2(new_n544), .ZN(new_n761));
  XNOR2_X1  g560(.A(KEYINPUT105), .B(G78gat), .ZN(new_n762));
  XNOR2_X1  g561(.A(new_n761), .B(new_n762), .ZN(G1335gat));
  INV_X1    g562(.A(new_n635), .ZN(new_n764));
  NOR2_X1   g563(.A1(new_n598), .A2(new_n717), .ZN(new_n765));
  NAND3_X1  g564(.A1(new_n746), .A2(new_n764), .A3(new_n765), .ZN(new_n766));
  INV_X1    g565(.A(KEYINPUT51), .ZN(new_n767));
  XNOR2_X1  g566(.A(new_n766), .B(new_n767), .ZN(new_n768));
  NAND2_X1  g567(.A1(new_n768), .A2(new_n657), .ZN(new_n769));
  NOR3_X1   g568(.A1(new_n769), .A2(G85gat), .A3(new_n546), .ZN(new_n770));
  NOR3_X1   g569(.A1(new_n598), .A2(new_n717), .A3(new_n718), .ZN(new_n771));
  AOI21_X1  g570(.A(new_n635), .B1(new_n556), .B2(new_n745), .ZN(new_n772));
  OAI211_X1 g571(.A(new_n710), .B(new_n771), .C1(new_n772), .C2(KEYINPUT44), .ZN(new_n773));
  INV_X1    g572(.A(KEYINPUT106), .ZN(new_n774));
  NAND2_X1  g573(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  NAND4_X1  g574(.A1(new_n695), .A2(KEYINPUT106), .A3(new_n710), .A4(new_n771), .ZN(new_n776));
  AND2_X1   g575(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  AOI21_X1  g576(.A(new_n605), .B1(new_n777), .B2(new_n712), .ZN(new_n778));
  OR2_X1    g577(.A1(new_n770), .A2(new_n778), .ZN(G1336gat));
  NOR2_X1   g578(.A1(new_n545), .A2(G92gat), .ZN(new_n780));
  NOR2_X1   g579(.A1(new_n766), .A2(new_n767), .ZN(new_n781));
  AOI21_X1  g580(.A(KEYINPUT51), .B1(new_n772), .B2(new_n765), .ZN(new_n782));
  OAI211_X1 g581(.A(new_n657), .B(new_n780), .C1(new_n781), .C2(new_n782), .ZN(new_n783));
  INV_X1    g582(.A(KEYINPUT52), .ZN(new_n784));
  OAI21_X1  g583(.A(G92gat), .B1(new_n773), .B2(new_n545), .ZN(new_n785));
  NAND3_X1  g584(.A1(new_n783), .A2(new_n784), .A3(new_n785), .ZN(new_n786));
  NAND3_X1  g585(.A1(new_n775), .A2(new_n415), .A3(new_n776), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n787), .A2(G92gat), .ZN(new_n788));
  INV_X1    g587(.A(KEYINPUT107), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n783), .A2(new_n789), .ZN(new_n790));
  NAND4_X1  g589(.A1(new_n768), .A2(KEYINPUT107), .A3(new_n657), .A4(new_n780), .ZN(new_n791));
  NAND3_X1  g590(.A1(new_n788), .A2(new_n790), .A3(new_n791), .ZN(new_n792));
  INV_X1    g591(.A(KEYINPUT108), .ZN(new_n793));
  AND3_X1   g592(.A1(new_n792), .A2(new_n793), .A3(KEYINPUT52), .ZN(new_n794));
  AOI21_X1  g593(.A(new_n793), .B1(new_n792), .B2(KEYINPUT52), .ZN(new_n795));
  OAI21_X1  g594(.A(new_n786), .B1(new_n794), .B2(new_n795), .ZN(G1337gat));
  NOR3_X1   g595(.A1(new_n769), .A2(G99gat), .A3(new_n734), .ZN(new_n797));
  INV_X1    g596(.A(G99gat), .ZN(new_n798));
  AOI21_X1  g597(.A(new_n798), .B1(new_n777), .B2(new_n732), .ZN(new_n799));
  OR2_X1    g598(.A1(new_n797), .A2(new_n799), .ZN(G1338gat));
  NOR3_X1   g599(.A1(new_n769), .A2(G106gat), .A3(new_n544), .ZN(new_n801));
  NOR2_X1   g600(.A1(new_n801), .A2(KEYINPUT53), .ZN(new_n802));
  OAI21_X1  g601(.A(G106gat), .B1(new_n773), .B2(new_n544), .ZN(new_n803));
  NAND2_X1  g602(.A1(new_n802), .A2(new_n803), .ZN(new_n804));
  INV_X1    g603(.A(G106gat), .ZN(new_n805));
  AOI21_X1  g604(.A(new_n805), .B1(new_n777), .B2(new_n338), .ZN(new_n806));
  OAI21_X1  g605(.A(KEYINPUT53), .B1(new_n801), .B2(new_n806), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n804), .A2(new_n807), .ZN(G1339gat));
  NAND3_X1  g607(.A1(new_n647), .A2(new_n638), .A3(new_n648), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n809), .A2(KEYINPUT109), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n647), .A2(new_n648), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n811), .A2(new_n637), .ZN(new_n812));
  INV_X1    g611(.A(KEYINPUT109), .ZN(new_n813));
  NAND4_X1  g612(.A1(new_n647), .A2(new_n813), .A3(new_n648), .A4(new_n638), .ZN(new_n814));
  NAND4_X1  g613(.A1(new_n810), .A2(new_n812), .A3(KEYINPUT54), .A4(new_n814), .ZN(new_n815));
  INV_X1    g614(.A(KEYINPUT54), .ZN(new_n816));
  AOI21_X1  g615(.A(new_n654), .B1(new_n649), .B2(new_n816), .ZN(new_n817));
  NAND4_X1  g616(.A1(new_n815), .A2(KEYINPUT110), .A3(KEYINPUT55), .A4(new_n817), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n818), .A2(new_n656), .ZN(new_n819));
  AND2_X1   g618(.A1(new_n817), .A2(KEYINPUT55), .ZN(new_n820));
  AOI21_X1  g619(.A(KEYINPUT110), .B1(new_n820), .B2(new_n815), .ZN(new_n821));
  NOR2_X1   g620(.A1(new_n819), .A2(new_n821), .ZN(new_n822));
  AOI21_X1  g621(.A(KEYINPUT55), .B1(new_n815), .B2(new_n817), .ZN(new_n823));
  INV_X1    g622(.A(KEYINPUT111), .ZN(new_n824));
  NOR2_X1   g623(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  AOI211_X1 g624(.A(KEYINPUT111), .B(KEYINPUT55), .C1(new_n815), .C2(new_n817), .ZN(new_n826));
  OAI211_X1 g625(.A(new_n822), .B(new_n717), .C1(new_n825), .C2(new_n826), .ZN(new_n827));
  AND3_X1   g626(.A1(new_n269), .A2(new_n270), .A3(new_n262), .ZN(new_n828));
  AOI21_X1  g627(.A(new_n208), .B1(new_n269), .B2(new_n246), .ZN(new_n829));
  OAI21_X1  g628(.A(new_n205), .B1(new_n828), .B2(new_n829), .ZN(new_n830));
  NAND3_X1  g629(.A1(new_n657), .A2(new_n716), .A3(new_n830), .ZN(new_n831));
  AOI21_X1  g630(.A(new_n764), .B1(new_n827), .B2(new_n831), .ZN(new_n832));
  NOR2_X1   g631(.A1(new_n825), .A2(new_n826), .ZN(new_n833));
  INV_X1    g632(.A(KEYINPUT110), .ZN(new_n834));
  INV_X1    g633(.A(new_n815), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n817), .A2(KEYINPUT55), .ZN(new_n836));
  OAI21_X1  g635(.A(new_n834), .B1(new_n835), .B2(new_n836), .ZN(new_n837));
  NAND3_X1  g636(.A1(new_n837), .A2(new_n656), .A3(new_n818), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n716), .A2(new_n830), .ZN(new_n839));
  NOR4_X1   g638(.A1(new_n833), .A2(new_n635), .A3(new_n838), .A4(new_n839), .ZN(new_n840));
  OAI21_X1  g639(.A(new_n713), .B1(new_n832), .B2(new_n840), .ZN(new_n841));
  NOR3_X1   g640(.A1(new_n636), .A2(new_n717), .A3(new_n657), .ZN(new_n842));
  INV_X1    g641(.A(new_n842), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n841), .A2(new_n843), .ZN(new_n844));
  NOR2_X1   g643(.A1(new_n415), .A2(new_n546), .ZN(new_n845));
  NAND4_X1  g644(.A1(new_n844), .A2(new_n544), .A3(new_n673), .A4(new_n845), .ZN(new_n846));
  OAI21_X1  g645(.A(G113gat), .B1(new_n846), .B2(new_n276), .ZN(new_n847));
  NOR3_X1   g646(.A1(new_n833), .A2(new_n838), .A3(new_n276), .ZN(new_n848));
  INV_X1    g647(.A(new_n831), .ZN(new_n849));
  OAI21_X1  g648(.A(new_n635), .B1(new_n848), .B2(new_n849), .ZN(new_n850));
  NOR2_X1   g649(.A1(new_n833), .A2(new_n838), .ZN(new_n851));
  INV_X1    g650(.A(new_n839), .ZN(new_n852));
  NAND3_X1  g651(.A1(new_n851), .A2(new_n764), .A3(new_n852), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n850), .A2(new_n853), .ZN(new_n854));
  AOI21_X1  g653(.A(new_n842), .B1(new_n854), .B2(new_n713), .ZN(new_n855));
  NOR2_X1   g654(.A1(new_n855), .A2(new_n546), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n856), .A2(new_n550), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n717), .A2(new_n416), .ZN(new_n858));
  OAI21_X1  g657(.A(new_n847), .B1(new_n857), .B2(new_n858), .ZN(new_n859));
  XNOR2_X1  g658(.A(new_n859), .B(KEYINPUT112), .ZN(G1340gat));
  NOR4_X1   g659(.A1(new_n857), .A2(new_n428), .A3(new_n427), .A4(new_n718), .ZN(new_n861));
  NOR2_X1   g660(.A1(new_n846), .A2(new_n718), .ZN(new_n862));
  NOR2_X1   g661(.A1(new_n862), .A2(new_n417), .ZN(new_n863));
  OR3_X1    g662(.A1(new_n861), .A2(KEYINPUT113), .A3(new_n863), .ZN(new_n864));
  OAI21_X1  g663(.A(KEYINPUT113), .B1(new_n861), .B2(new_n863), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n864), .A2(new_n865), .ZN(G1341gat));
  OAI21_X1  g665(.A(G127gat), .B1(new_n846), .B2(new_n713), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n598), .A2(new_n422), .ZN(new_n868));
  OAI21_X1  g667(.A(new_n867), .B1(new_n857), .B2(new_n868), .ZN(G1342gat));
  NOR3_X1   g668(.A1(new_n635), .A2(new_n464), .A3(new_n415), .ZN(new_n870));
  NAND4_X1  g669(.A1(new_n856), .A2(new_n544), .A3(new_n673), .A4(new_n870), .ZN(new_n871));
  XOR2_X1   g670(.A(new_n871), .B(KEYINPUT56), .Z(new_n872));
  OAI21_X1  g671(.A(G134gat), .B1(new_n846), .B2(new_n635), .ZN(new_n873));
  NAND2_X1  g672(.A1(new_n872), .A2(new_n873), .ZN(G1343gat));
  INV_X1    g673(.A(new_n845), .ZN(new_n875));
  NOR2_X1   g674(.A1(new_n732), .A2(new_n875), .ZN(new_n876));
  INV_X1    g675(.A(KEYINPUT57), .ZN(new_n877));
  NOR2_X1   g676(.A1(new_n544), .A2(new_n877), .ZN(new_n878));
  INV_X1    g677(.A(new_n878), .ZN(new_n879));
  AND2_X1   g678(.A1(new_n815), .A2(new_n817), .ZN(new_n880));
  OAI22_X1  g679(.A1(new_n273), .A2(new_n275), .B1(KEYINPUT55), .B2(new_n880), .ZN(new_n881));
  OAI21_X1  g680(.A(new_n831), .B1(new_n881), .B2(new_n838), .ZN(new_n882));
  NAND2_X1  g681(.A1(new_n882), .A2(new_n635), .ZN(new_n883));
  NAND2_X1  g682(.A1(new_n853), .A2(new_n883), .ZN(new_n884));
  NAND2_X1  g683(.A1(new_n884), .A2(new_n713), .ZN(new_n885));
  AOI21_X1  g684(.A(new_n842), .B1(new_n885), .B2(KEYINPUT115), .ZN(new_n886));
  AOI21_X1  g685(.A(new_n598), .B1(new_n853), .B2(new_n883), .ZN(new_n887));
  INV_X1    g686(.A(KEYINPUT115), .ZN(new_n888));
  NAND2_X1  g687(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  AOI21_X1  g688(.A(new_n879), .B1(new_n886), .B2(new_n889), .ZN(new_n890));
  AOI21_X1  g689(.A(new_n544), .B1(new_n841), .B2(new_n843), .ZN(new_n891));
  XNOR2_X1  g690(.A(KEYINPUT114), .B(KEYINPUT57), .ZN(new_n892));
  INV_X1    g691(.A(new_n892), .ZN(new_n893));
  NOR2_X1   g692(.A1(new_n891), .A2(new_n893), .ZN(new_n894));
  OAI21_X1  g693(.A(new_n876), .B1(new_n890), .B2(new_n894), .ZN(new_n895));
  OAI21_X1  g694(.A(G141gat), .B1(new_n895), .B2(new_n276), .ZN(new_n896));
  NAND2_X1  g695(.A1(new_n675), .A2(new_n338), .ZN(new_n897));
  NOR2_X1   g696(.A1(new_n897), .A2(new_n415), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n717), .A2(new_n282), .ZN(new_n899));
  XNOR2_X1  g698(.A(new_n899), .B(KEYINPUT117), .ZN(new_n900));
  NAND3_X1  g699(.A1(new_n856), .A2(new_n898), .A3(new_n900), .ZN(new_n901));
  NAND2_X1  g700(.A1(new_n896), .A2(new_n901), .ZN(new_n902));
  INV_X1    g701(.A(KEYINPUT116), .ZN(new_n903));
  NAND2_X1  g702(.A1(new_n901), .A2(new_n903), .ZN(new_n904));
  NAND2_X1  g703(.A1(new_n904), .A2(KEYINPUT58), .ZN(new_n905));
  INV_X1    g704(.A(new_n905), .ZN(new_n906));
  NAND2_X1  g705(.A1(new_n902), .A2(new_n906), .ZN(new_n907));
  NAND3_X1  g706(.A1(new_n896), .A2(new_n901), .A3(new_n905), .ZN(new_n908));
  NAND2_X1  g707(.A1(new_n907), .A2(new_n908), .ZN(G1344gat));
  AND2_X1   g708(.A1(new_n856), .A2(new_n898), .ZN(new_n910));
  NAND3_X1  g709(.A1(new_n910), .A2(new_n283), .A3(new_n657), .ZN(new_n911));
  NAND2_X1  g710(.A1(new_n876), .A2(new_n657), .ZN(new_n912));
  NAND2_X1  g711(.A1(new_n891), .A2(new_n893), .ZN(new_n913));
  OAI21_X1  g712(.A(new_n338), .B1(new_n887), .B2(new_n842), .ZN(new_n914));
  NAND2_X1  g713(.A1(new_n914), .A2(new_n877), .ZN(new_n915));
  AOI21_X1  g714(.A(new_n912), .B1(new_n913), .B2(new_n915), .ZN(new_n916));
  OAI211_X1 g715(.A(KEYINPUT118), .B(KEYINPUT59), .C1(new_n916), .C2(new_n283), .ZN(new_n917));
  INV_X1    g716(.A(new_n917), .ZN(new_n918));
  AOI22_X1  g717(.A1(new_n891), .A2(new_n893), .B1(new_n914), .B2(new_n877), .ZN(new_n919));
  OAI21_X1  g718(.A(G148gat), .B1(new_n919), .B2(new_n912), .ZN(new_n920));
  AOI21_X1  g719(.A(KEYINPUT118), .B1(new_n920), .B2(KEYINPUT59), .ZN(new_n921));
  NOR2_X1   g720(.A1(new_n918), .A2(new_n921), .ZN(new_n922));
  NOR2_X1   g721(.A1(new_n895), .A2(new_n718), .ZN(new_n923));
  NOR3_X1   g722(.A1(new_n923), .A2(KEYINPUT59), .A3(new_n283), .ZN(new_n924));
  OAI21_X1  g723(.A(new_n911), .B1(new_n922), .B2(new_n924), .ZN(G1345gat));
  OAI21_X1  g724(.A(G155gat), .B1(new_n895), .B2(new_n713), .ZN(new_n926));
  NAND3_X1  g725(.A1(new_n910), .A2(new_n294), .A3(new_n598), .ZN(new_n927));
  NAND2_X1  g726(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  INV_X1    g727(.A(KEYINPUT119), .ZN(new_n929));
  NAND2_X1  g728(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  NAND3_X1  g729(.A1(new_n926), .A2(KEYINPUT119), .A3(new_n927), .ZN(new_n931));
  NAND2_X1  g730(.A1(new_n930), .A2(new_n931), .ZN(G1346gat));
  OAI21_X1  g731(.A(G162gat), .B1(new_n895), .B2(new_n635), .ZN(new_n933));
  NAND3_X1  g732(.A1(new_n910), .A2(new_n295), .A3(new_n764), .ZN(new_n934));
  NAND2_X1  g733(.A1(new_n933), .A2(new_n934), .ZN(G1347gat));
  NOR2_X1   g734(.A1(new_n712), .A2(new_n545), .ZN(new_n936));
  INV_X1    g735(.A(new_n936), .ZN(new_n937));
  NOR2_X1   g736(.A1(new_n937), .A2(new_n734), .ZN(new_n938));
  NAND3_X1  g737(.A1(new_n844), .A2(new_n544), .A3(new_n938), .ZN(new_n939));
  OAI21_X1  g738(.A(G169gat), .B1(new_n939), .B2(new_n276), .ZN(new_n940));
  INV_X1    g739(.A(KEYINPUT122), .ZN(new_n941));
  NAND2_X1  g740(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  NOR3_X1   g741(.A1(new_n734), .A2(new_n545), .A3(new_n338), .ZN(new_n943));
  AOI21_X1  g742(.A(KEYINPUT120), .B1(new_n844), .B2(new_n546), .ZN(new_n944));
  INV_X1    g743(.A(KEYINPUT120), .ZN(new_n945));
  AOI211_X1 g744(.A(new_n945), .B(new_n712), .C1(new_n841), .C2(new_n843), .ZN(new_n946));
  OAI21_X1  g745(.A(new_n943), .B1(new_n944), .B2(new_n946), .ZN(new_n947));
  NAND2_X1  g746(.A1(new_n947), .A2(KEYINPUT121), .ZN(new_n948));
  INV_X1    g747(.A(KEYINPUT121), .ZN(new_n949));
  OAI211_X1 g748(.A(new_n949), .B(new_n943), .C1(new_n944), .C2(new_n946), .ZN(new_n950));
  NAND2_X1  g749(.A1(new_n948), .A2(new_n950), .ZN(new_n951));
  NOR2_X1   g750(.A1(new_n276), .A2(G169gat), .ZN(new_n952));
  AOI21_X1  g751(.A(new_n942), .B1(new_n951), .B2(new_n952), .ZN(new_n953));
  INV_X1    g752(.A(new_n952), .ZN(new_n954));
  AOI211_X1 g753(.A(new_n941), .B(new_n954), .C1(new_n948), .C2(new_n950), .ZN(new_n955));
  NOR2_X1   g754(.A1(new_n953), .A2(new_n955), .ZN(G1348gat));
  INV_X1    g755(.A(G176gat), .ZN(new_n957));
  NAND3_X1  g756(.A1(new_n951), .A2(new_n957), .A3(new_n657), .ZN(new_n958));
  OAI21_X1  g757(.A(G176gat), .B1(new_n939), .B2(new_n718), .ZN(new_n959));
  NAND2_X1  g758(.A1(new_n958), .A2(new_n959), .ZN(G1349gat));
  NOR2_X1   g759(.A1(KEYINPUT124), .A2(KEYINPUT60), .ZN(new_n961));
  INV_X1    g760(.A(new_n961), .ZN(new_n962));
  AND2_X1   g761(.A1(new_n598), .A2(new_n353), .ZN(new_n963));
  OAI211_X1 g762(.A(new_n943), .B(new_n963), .C1(new_n944), .C2(new_n946), .ZN(new_n964));
  NAND2_X1  g763(.A1(new_n964), .A2(KEYINPUT123), .ZN(new_n965));
  OAI21_X1  g764(.A(new_n945), .B1(new_n855), .B2(new_n712), .ZN(new_n966));
  NAND3_X1  g765(.A1(new_n844), .A2(KEYINPUT120), .A3(new_n546), .ZN(new_n967));
  NAND2_X1  g766(.A1(new_n966), .A2(new_n967), .ZN(new_n968));
  INV_X1    g767(.A(KEYINPUT123), .ZN(new_n969));
  NAND4_X1  g768(.A1(new_n968), .A2(new_n969), .A3(new_n943), .A4(new_n963), .ZN(new_n970));
  NAND2_X1  g769(.A1(new_n965), .A2(new_n970), .ZN(new_n971));
  OAI21_X1  g770(.A(G183gat), .B1(new_n939), .B2(new_n713), .ZN(new_n972));
  NAND2_X1  g771(.A1(KEYINPUT124), .A2(KEYINPUT60), .ZN(new_n973));
  NAND2_X1  g772(.A1(new_n972), .A2(new_n973), .ZN(new_n974));
  INV_X1    g773(.A(new_n974), .ZN(new_n975));
  AOI21_X1  g774(.A(new_n962), .B1(new_n971), .B2(new_n975), .ZN(new_n976));
  AOI211_X1 g775(.A(new_n961), .B(new_n974), .C1(new_n965), .C2(new_n970), .ZN(new_n977));
  NOR2_X1   g776(.A1(new_n976), .A2(new_n977), .ZN(G1350gat));
  OAI21_X1  g777(.A(G190gat), .B1(new_n939), .B2(new_n635), .ZN(new_n979));
  XNOR2_X1  g778(.A(new_n979), .B(KEYINPUT61), .ZN(new_n980));
  INV_X1    g779(.A(KEYINPUT125), .ZN(new_n981));
  NOR2_X1   g780(.A1(new_n635), .A2(G190gat), .ZN(new_n982));
  AOI21_X1  g781(.A(new_n981), .B1(new_n951), .B2(new_n982), .ZN(new_n983));
  INV_X1    g782(.A(new_n982), .ZN(new_n984));
  AOI211_X1 g783(.A(KEYINPUT125), .B(new_n984), .C1(new_n948), .C2(new_n950), .ZN(new_n985));
  OAI21_X1  g784(.A(new_n980), .B1(new_n983), .B2(new_n985), .ZN(G1351gat));
  NOR2_X1   g785(.A1(new_n732), .A2(new_n937), .ZN(new_n987));
  OR2_X1    g786(.A1(new_n987), .A2(KEYINPUT126), .ZN(new_n988));
  NAND2_X1  g787(.A1(new_n987), .A2(KEYINPUT126), .ZN(new_n989));
  AOI21_X1  g788(.A(new_n919), .B1(new_n988), .B2(new_n989), .ZN(new_n990));
  AND3_X1   g789(.A1(new_n990), .A2(G197gat), .A3(new_n717), .ZN(new_n991));
  AOI211_X1 g790(.A(new_n545), .B(new_n897), .C1(new_n966), .C2(new_n967), .ZN(new_n992));
  AOI21_X1  g791(.A(G197gat), .B1(new_n992), .B2(new_n717), .ZN(new_n993));
  NOR2_X1   g792(.A1(new_n991), .A2(new_n993), .ZN(G1352gat));
  XOR2_X1   g793(.A(KEYINPUT127), .B(G204gat), .Z(new_n995));
  NOR2_X1   g794(.A1(new_n718), .A2(new_n995), .ZN(new_n996));
  NAND2_X1  g795(.A1(new_n992), .A2(new_n996), .ZN(new_n997));
  OR2_X1    g796(.A1(new_n997), .A2(KEYINPUT62), .ZN(new_n998));
  INV_X1    g797(.A(new_n990), .ZN(new_n999));
  OAI21_X1  g798(.A(new_n995), .B1(new_n999), .B2(new_n718), .ZN(new_n1000));
  NAND2_X1  g799(.A1(new_n997), .A2(KEYINPUT62), .ZN(new_n1001));
  NAND3_X1  g800(.A1(new_n998), .A2(new_n1000), .A3(new_n1001), .ZN(G1353gat));
  INV_X1    g801(.A(G211gat), .ZN(new_n1003));
  NAND3_X1  g802(.A1(new_n992), .A2(new_n1003), .A3(new_n598), .ZN(new_n1004));
  NAND2_X1  g803(.A1(new_n990), .A2(new_n598), .ZN(new_n1005));
  AND3_X1   g804(.A1(new_n1005), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n1006));
  AOI21_X1  g805(.A(KEYINPUT63), .B1(new_n1005), .B2(G211gat), .ZN(new_n1007));
  OAI21_X1  g806(.A(new_n1004), .B1(new_n1006), .B2(new_n1007), .ZN(G1354gat));
  OAI21_X1  g807(.A(G218gat), .B1(new_n999), .B2(new_n635), .ZN(new_n1009));
  INV_X1    g808(.A(G218gat), .ZN(new_n1010));
  NAND3_X1  g809(.A1(new_n992), .A2(new_n1010), .A3(new_n764), .ZN(new_n1011));
  NAND2_X1  g810(.A1(new_n1009), .A2(new_n1011), .ZN(G1355gat));
endmodule


