//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 0 0 1 0 0 0 1 0 1 1 1 0 0 1 0 1 1 0 1 1 1 0 0 1 0 0 1 1 1 1 1 1 1 1 1 0 0 1 0 1 0 1 0 0 1 0 0 1 0 1 0 0 0 1 1 1 1 0 0 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:15:58 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n684, new_n685, new_n686,
    new_n688, new_n689, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n707, new_n708, new_n709, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n742,
    new_n743, new_n744, new_n746, new_n747, new_n748, new_n749, new_n750,
    new_n751, new_n752, new_n754, new_n756, new_n757, new_n758, new_n759,
    new_n760, new_n761, new_n762, new_n763, new_n764, new_n765, new_n766,
    new_n767, new_n768, new_n769, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n780, new_n781, new_n782,
    new_n783, new_n784, new_n785, new_n786, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n842, new_n843, new_n845, new_n846, new_n847, new_n848, new_n850,
    new_n851, new_n852, new_n853, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n907, new_n908, new_n910,
    new_n911, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n932, new_n933, new_n934,
    new_n936, new_n937, new_n938, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n957, new_n958, new_n959,
    new_n960, new_n961, new_n962, new_n963, new_n964, new_n966, new_n967,
    new_n968;
  XOR2_X1   g000(.A(G141gat), .B(G148gat), .Z(new_n202));
  INV_X1    g001(.A(G155gat), .ZN(new_n203));
  INV_X1    g002(.A(G162gat), .ZN(new_n204));
  NAND2_X1  g003(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  NAND2_X1  g004(.A1(G155gat), .A2(G162gat), .ZN(new_n206));
  NAND2_X1  g005(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  NAND2_X1  g006(.A1(new_n206), .A2(KEYINPUT2), .ZN(new_n208));
  NAND3_X1  g007(.A1(new_n202), .A2(new_n207), .A3(new_n208), .ZN(new_n209));
  XNOR2_X1  g008(.A(G141gat), .B(G148gat), .ZN(new_n210));
  OAI211_X1 g009(.A(new_n206), .B(new_n205), .C1(new_n210), .C2(KEYINPUT2), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n209), .A2(new_n211), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n212), .A2(KEYINPUT3), .ZN(new_n213));
  NOR2_X1   g012(.A1(G127gat), .A2(G134gat), .ZN(new_n214));
  INV_X1    g013(.A(G127gat), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n215), .A2(KEYINPUT70), .ZN(new_n216));
  INV_X1    g015(.A(KEYINPUT70), .ZN(new_n217));
  NAND2_X1  g016(.A1(new_n217), .A2(G127gat), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n216), .A2(new_n218), .ZN(new_n219));
  AOI21_X1  g018(.A(new_n214), .B1(new_n219), .B2(G134gat), .ZN(new_n220));
  INV_X1    g019(.A(KEYINPUT1), .ZN(new_n221));
  OAI21_X1  g020(.A(new_n221), .B1(G113gat), .B2(G120gat), .ZN(new_n222));
  INV_X1    g021(.A(new_n222), .ZN(new_n223));
  NAND2_X1  g022(.A1(G113gat), .A2(G120gat), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n220), .A2(new_n225), .ZN(new_n226));
  INV_X1    g025(.A(new_n214), .ZN(new_n227));
  NAND2_X1  g026(.A1(G127gat), .A2(G134gat), .ZN(new_n228));
  AOI21_X1  g027(.A(new_n222), .B1(new_n227), .B2(new_n228), .ZN(new_n229));
  INV_X1    g028(.A(G120gat), .ZN(new_n230));
  AND2_X1   g029(.A1(new_n230), .A2(KEYINPUT71), .ZN(new_n231));
  NOR2_X1   g030(.A1(new_n230), .A2(KEYINPUT71), .ZN(new_n232));
  OAI21_X1  g031(.A(G113gat), .B1(new_n231), .B2(new_n232), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n229), .A2(new_n233), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n226), .A2(new_n234), .ZN(new_n235));
  INV_X1    g034(.A(KEYINPUT3), .ZN(new_n236));
  NAND3_X1  g035(.A1(new_n209), .A2(new_n211), .A3(new_n236), .ZN(new_n237));
  NAND3_X1  g036(.A1(new_n213), .A2(new_n235), .A3(new_n237), .ZN(new_n238));
  NAND2_X1  g037(.A1(G225gat), .A2(G233gat), .ZN(new_n239));
  XNOR2_X1  g038(.A(new_n239), .B(KEYINPUT77), .ZN(new_n240));
  INV_X1    g039(.A(new_n240), .ZN(new_n241));
  AND2_X1   g040(.A1(new_n238), .A2(new_n241), .ZN(new_n242));
  INV_X1    g041(.A(KEYINPUT5), .ZN(new_n243));
  INV_X1    g042(.A(KEYINPUT78), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n212), .A2(new_n244), .ZN(new_n245));
  AOI22_X1  g044(.A1(new_n220), .A2(new_n225), .B1(new_n229), .B2(new_n233), .ZN(new_n246));
  NAND3_X1  g045(.A1(new_n209), .A2(new_n211), .A3(KEYINPUT78), .ZN(new_n247));
  NAND3_X1  g046(.A1(new_n245), .A2(new_n246), .A3(new_n247), .ZN(new_n248));
  INV_X1    g047(.A(KEYINPUT4), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n248), .A2(new_n249), .ZN(new_n250));
  OAI21_X1  g049(.A(KEYINPUT79), .B1(new_n235), .B2(new_n212), .ZN(new_n251));
  INV_X1    g050(.A(KEYINPUT79), .ZN(new_n252));
  NAND4_X1  g051(.A1(new_n246), .A2(new_n252), .A3(new_n211), .A4(new_n209), .ZN(new_n253));
  NAND3_X1  g052(.A1(new_n251), .A2(new_n253), .A3(KEYINPUT4), .ZN(new_n254));
  NAND4_X1  g053(.A1(new_n242), .A2(new_n243), .A3(new_n250), .A4(new_n254), .ZN(new_n255));
  AOI22_X1  g054(.A1(new_n251), .A2(new_n253), .B1(new_n212), .B2(new_n235), .ZN(new_n256));
  OAI21_X1  g055(.A(KEYINPUT5), .B1(new_n256), .B2(new_n241), .ZN(new_n257));
  OAI211_X1 g056(.A(new_n241), .B(new_n238), .C1(new_n248), .C2(new_n249), .ZN(new_n258));
  AOI21_X1  g057(.A(KEYINPUT4), .B1(new_n251), .B2(new_n253), .ZN(new_n259));
  NOR2_X1   g058(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  OAI21_X1  g059(.A(new_n255), .B1(new_n257), .B2(new_n260), .ZN(new_n261));
  XOR2_X1   g060(.A(G1gat), .B(G29gat), .Z(new_n262));
  XNOR2_X1  g061(.A(KEYINPUT80), .B(KEYINPUT0), .ZN(new_n263));
  XNOR2_X1  g062(.A(new_n262), .B(new_n263), .ZN(new_n264));
  XNOR2_X1  g063(.A(G57gat), .B(G85gat), .ZN(new_n265));
  XOR2_X1   g064(.A(new_n264), .B(new_n265), .Z(new_n266));
  INV_X1    g065(.A(new_n266), .ZN(new_n267));
  XOR2_X1   g066(.A(KEYINPUT81), .B(KEYINPUT6), .Z(new_n268));
  INV_X1    g067(.A(new_n268), .ZN(new_n269));
  NAND3_X1  g068(.A1(new_n261), .A2(new_n267), .A3(new_n269), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n270), .A2(KEYINPUT82), .ZN(new_n271));
  INV_X1    g070(.A(KEYINPUT82), .ZN(new_n272));
  NAND4_X1  g071(.A1(new_n261), .A2(new_n272), .A3(new_n267), .A4(new_n269), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n271), .A2(new_n273), .ZN(new_n274));
  AOI21_X1  g073(.A(new_n269), .B1(new_n261), .B2(new_n267), .ZN(new_n275));
  OAI21_X1  g074(.A(new_n275), .B1(new_n267), .B2(new_n261), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n274), .A2(new_n276), .ZN(new_n277));
  INV_X1    g076(.A(new_n277), .ZN(new_n278));
  XNOR2_X1  g077(.A(G8gat), .B(G36gat), .ZN(new_n279));
  XNOR2_X1  g078(.A(G64gat), .B(G92gat), .ZN(new_n280));
  XOR2_X1   g079(.A(new_n279), .B(new_n280), .Z(new_n281));
  XNOR2_X1  g080(.A(G197gat), .B(G204gat), .ZN(new_n282));
  INV_X1    g081(.A(KEYINPUT22), .ZN(new_n283));
  INV_X1    g082(.A(G211gat), .ZN(new_n284));
  INV_X1    g083(.A(G218gat), .ZN(new_n285));
  OAI21_X1  g084(.A(new_n283), .B1(new_n284), .B2(new_n285), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n282), .A2(new_n286), .ZN(new_n287));
  XNOR2_X1  g086(.A(G211gat), .B(G218gat), .ZN(new_n288));
  INV_X1    g087(.A(new_n288), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n287), .A2(new_n289), .ZN(new_n290));
  NAND3_X1  g089(.A1(new_n288), .A2(new_n282), .A3(new_n286), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  INV_X1    g091(.A(new_n292), .ZN(new_n293));
  INV_X1    g092(.A(KEYINPUT25), .ZN(new_n294));
  INV_X1    g093(.A(KEYINPUT65), .ZN(new_n295));
  NAND2_X1  g094(.A1(G169gat), .A2(G176gat), .ZN(new_n296));
  NAND2_X1  g095(.A1(new_n296), .A2(KEYINPUT23), .ZN(new_n297));
  INV_X1    g096(.A(G169gat), .ZN(new_n298));
  INV_X1    g097(.A(G176gat), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n298), .A2(new_n299), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n297), .A2(new_n300), .ZN(new_n301));
  INV_X1    g100(.A(KEYINPUT64), .ZN(new_n302));
  AND4_X1   g101(.A1(new_n302), .A2(new_n298), .A3(new_n299), .A4(KEYINPUT23), .ZN(new_n303));
  NOR2_X1   g102(.A1(G169gat), .A2(G176gat), .ZN(new_n304));
  AOI21_X1  g103(.A(new_n302), .B1(new_n304), .B2(KEYINPUT23), .ZN(new_n305));
  OAI211_X1 g104(.A(new_n295), .B(new_n301), .C1(new_n303), .C2(new_n305), .ZN(new_n306));
  OAI21_X1  g105(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n307));
  INV_X1    g106(.A(G183gat), .ZN(new_n308));
  INV_X1    g107(.A(G190gat), .ZN(new_n309));
  OAI21_X1  g108(.A(new_n307), .B1(new_n308), .B2(new_n309), .ZN(new_n310));
  NAND3_X1  g109(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n306), .A2(new_n312), .ZN(new_n313));
  NAND3_X1  g112(.A1(new_n298), .A2(new_n299), .A3(KEYINPUT23), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n314), .A2(KEYINPUT64), .ZN(new_n315));
  NAND3_X1  g114(.A1(new_n304), .A2(new_n302), .A3(KEYINPUT23), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n315), .A2(new_n316), .ZN(new_n317));
  AOI21_X1  g116(.A(new_n295), .B1(new_n317), .B2(new_n301), .ZN(new_n318));
  OAI21_X1  g117(.A(new_n294), .B1(new_n313), .B2(new_n318), .ZN(new_n319));
  XOR2_X1   g118(.A(new_n311), .B(KEYINPUT66), .Z(new_n320));
  NAND2_X1  g119(.A1(new_n320), .A2(new_n310), .ZN(new_n321));
  NAND4_X1  g120(.A1(new_n321), .A2(KEYINPUT25), .A3(new_n301), .A4(new_n314), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n319), .A2(new_n322), .ZN(new_n323));
  INV_X1    g122(.A(G226gat), .ZN(new_n324));
  INV_X1    g123(.A(G233gat), .ZN(new_n325));
  NOR2_X1   g124(.A1(new_n324), .A2(new_n325), .ZN(new_n326));
  INV_X1    g125(.A(new_n326), .ZN(new_n327));
  INV_X1    g126(.A(KEYINPUT68), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n308), .A2(KEYINPUT27), .ZN(new_n329));
  INV_X1    g128(.A(KEYINPUT27), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n330), .A2(G183gat), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n329), .A2(new_n331), .ZN(new_n332));
  NOR3_X1   g131(.A1(new_n332), .A2(KEYINPUT28), .A3(G190gat), .ZN(new_n333));
  INV_X1    g132(.A(new_n333), .ZN(new_n334));
  AND3_X1   g133(.A1(new_n329), .A2(new_n331), .A3(KEYINPUT67), .ZN(new_n335));
  AOI21_X1  g134(.A(KEYINPUT67), .B1(new_n329), .B2(new_n331), .ZN(new_n336));
  NOR3_X1   g135(.A1(new_n335), .A2(new_n336), .A3(G190gat), .ZN(new_n337));
  INV_X1    g136(.A(KEYINPUT28), .ZN(new_n338));
  OAI211_X1 g137(.A(new_n328), .B(new_n334), .C1(new_n337), .C2(new_n338), .ZN(new_n339));
  INV_X1    g138(.A(KEYINPUT69), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n304), .A2(new_n340), .ZN(new_n341));
  OR2_X1    g140(.A1(new_n341), .A2(KEYINPUT26), .ZN(new_n342));
  AOI22_X1  g141(.A1(new_n341), .A2(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n343));
  AOI22_X1  g142(.A1(new_n342), .A2(new_n343), .B1(G183gat), .B2(G190gat), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n339), .A2(new_n344), .ZN(new_n345));
  INV_X1    g144(.A(KEYINPUT67), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n332), .A2(new_n346), .ZN(new_n347));
  XNOR2_X1  g146(.A(KEYINPUT27), .B(G183gat), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n348), .A2(KEYINPUT67), .ZN(new_n349));
  NAND3_X1  g148(.A1(new_n347), .A2(new_n349), .A3(new_n309), .ZN(new_n350));
  AOI21_X1  g149(.A(new_n333), .B1(new_n350), .B2(KEYINPUT28), .ZN(new_n351));
  NOR2_X1   g150(.A1(new_n351), .A2(new_n328), .ZN(new_n352));
  OAI211_X1 g151(.A(new_n323), .B(new_n327), .C1(new_n345), .C2(new_n352), .ZN(new_n353));
  OR2_X1    g152(.A1(new_n351), .A2(new_n328), .ZN(new_n354));
  INV_X1    g153(.A(new_n344), .ZN(new_n355));
  AOI21_X1  g154(.A(new_n355), .B1(new_n351), .B2(new_n328), .ZN(new_n356));
  AOI22_X1  g155(.A1(new_n354), .A2(new_n356), .B1(new_n319), .B2(new_n322), .ZN(new_n357));
  NOR2_X1   g156(.A1(new_n326), .A2(KEYINPUT29), .ZN(new_n358));
  OAI211_X1 g157(.A(new_n293), .B(new_n353), .C1(new_n357), .C2(new_n358), .ZN(new_n359));
  INV_X1    g158(.A(new_n359), .ZN(new_n360));
  AND3_X1   g159(.A1(new_n290), .A2(KEYINPUT75), .A3(new_n291), .ZN(new_n361));
  AOI21_X1  g160(.A(KEYINPUT75), .B1(new_n290), .B2(new_n291), .ZN(new_n362));
  NOR2_X1   g161(.A1(new_n361), .A2(new_n362), .ZN(new_n363));
  INV_X1    g162(.A(new_n363), .ZN(new_n364));
  OAI21_X1  g163(.A(new_n323), .B1(new_n345), .B2(new_n352), .ZN(new_n365));
  INV_X1    g164(.A(new_n358), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n365), .A2(new_n366), .ZN(new_n367));
  AOI21_X1  g166(.A(new_n364), .B1(new_n367), .B2(new_n353), .ZN(new_n368));
  OAI21_X1  g167(.A(new_n281), .B1(new_n360), .B2(new_n368), .ZN(new_n369));
  INV_X1    g168(.A(KEYINPUT37), .ZN(new_n370));
  OAI21_X1  g169(.A(new_n370), .B1(new_n360), .B2(new_n368), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n371), .A2(KEYINPUT86), .ZN(new_n372));
  INV_X1    g171(.A(KEYINPUT86), .ZN(new_n373));
  OAI211_X1 g172(.A(new_n373), .B(new_n370), .C1(new_n360), .C2(new_n368), .ZN(new_n374));
  NAND2_X1  g173(.A1(new_n372), .A2(new_n374), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n367), .A2(new_n353), .ZN(new_n376));
  AOI21_X1  g175(.A(new_n370), .B1(new_n376), .B2(new_n292), .ZN(new_n377));
  NAND3_X1  g176(.A1(new_n367), .A2(new_n353), .A3(new_n364), .ZN(new_n378));
  AOI21_X1  g177(.A(new_n281), .B1(new_n377), .B2(new_n378), .ZN(new_n379));
  AOI21_X1  g178(.A(KEYINPUT38), .B1(new_n375), .B2(new_n379), .ZN(new_n380));
  INV_X1    g179(.A(new_n368), .ZN(new_n381));
  NAND3_X1  g180(.A1(new_n381), .A2(KEYINPUT37), .A3(new_n359), .ZN(new_n382));
  INV_X1    g181(.A(new_n281), .ZN(new_n383));
  NAND3_X1  g182(.A1(new_n382), .A2(KEYINPUT38), .A3(new_n383), .ZN(new_n384));
  AOI21_X1  g183(.A(new_n384), .B1(new_n372), .B2(new_n374), .ZN(new_n385));
  OAI211_X1 g184(.A(new_n278), .B(new_n369), .C1(new_n380), .C2(new_n385), .ZN(new_n386));
  AND2_X1   g185(.A1(G228gat), .A2(G233gat), .ZN(new_n387));
  AOI21_X1  g186(.A(KEYINPUT29), .B1(new_n290), .B2(new_n291), .ZN(new_n388));
  OAI21_X1  g187(.A(new_n212), .B1(new_n388), .B2(KEYINPUT3), .ZN(new_n389));
  INV_X1    g188(.A(KEYINPUT29), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n237), .A2(new_n390), .ZN(new_n391));
  INV_X1    g190(.A(new_n391), .ZN(new_n392));
  OAI211_X1 g191(.A(new_n387), .B(new_n389), .C1(new_n363), .C2(new_n392), .ZN(new_n393));
  OR2_X1    g192(.A1(new_n388), .A2(KEYINPUT3), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n245), .A2(new_n247), .ZN(new_n395));
  AOI22_X1  g194(.A1(new_n394), .A2(new_n395), .B1(new_n293), .B2(new_n391), .ZN(new_n396));
  OAI21_X1  g195(.A(new_n393), .B1(new_n396), .B2(new_n387), .ZN(new_n397));
  XNOR2_X1  g196(.A(new_n397), .B(G22gat), .ZN(new_n398));
  INV_X1    g197(.A(KEYINPUT84), .ZN(new_n399));
  XNOR2_X1  g198(.A(G78gat), .B(G106gat), .ZN(new_n400));
  INV_X1    g199(.A(G50gat), .ZN(new_n401));
  XNOR2_X1  g200(.A(new_n400), .B(new_n401), .ZN(new_n402));
  XOR2_X1   g201(.A(KEYINPUT83), .B(KEYINPUT31), .Z(new_n403));
  XNOR2_X1  g202(.A(new_n402), .B(new_n403), .ZN(new_n404));
  INV_X1    g203(.A(new_n404), .ZN(new_n405));
  NOR3_X1   g204(.A1(new_n398), .A2(new_n399), .A3(new_n405), .ZN(new_n406));
  INV_X1    g205(.A(new_n406), .ZN(new_n407));
  INV_X1    g206(.A(G22gat), .ZN(new_n408));
  XNOR2_X1  g207(.A(new_n397), .B(new_n408), .ZN(new_n409));
  AOI21_X1  g208(.A(new_n404), .B1(new_n409), .B2(KEYINPUT84), .ZN(new_n410));
  INV_X1    g209(.A(new_n410), .ZN(new_n411));
  NOR2_X1   g210(.A1(new_n409), .A2(KEYINPUT84), .ZN(new_n412));
  OAI21_X1  g211(.A(new_n407), .B1(new_n411), .B2(new_n412), .ZN(new_n413));
  NAND3_X1  g212(.A1(new_n254), .A2(new_n250), .A3(new_n238), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n414), .A2(new_n240), .ZN(new_n415));
  INV_X1    g214(.A(KEYINPUT39), .ZN(new_n416));
  AOI21_X1  g215(.A(new_n416), .B1(new_n256), .B2(new_n241), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n415), .A2(new_n417), .ZN(new_n418));
  NAND3_X1  g217(.A1(new_n414), .A2(new_n416), .A3(new_n240), .ZN(new_n419));
  AND3_X1   g218(.A1(new_n419), .A2(KEYINPUT85), .A3(new_n266), .ZN(new_n420));
  AOI21_X1  g219(.A(KEYINPUT85), .B1(new_n419), .B2(new_n266), .ZN(new_n421));
  OAI21_X1  g220(.A(new_n418), .B1(new_n420), .B2(new_n421), .ZN(new_n422));
  INV_X1    g221(.A(KEYINPUT40), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n261), .A2(new_n267), .ZN(new_n425));
  OAI211_X1 g224(.A(KEYINPUT40), .B(new_n418), .C1(new_n420), .C2(new_n421), .ZN(new_n426));
  AND3_X1   g225(.A1(new_n424), .A2(new_n425), .A3(new_n426), .ZN(new_n427));
  OAI211_X1 g226(.A(KEYINPUT30), .B(new_n281), .C1(new_n360), .C2(new_n368), .ZN(new_n428));
  NAND3_X1  g227(.A1(new_n381), .A2(new_n359), .A3(new_n383), .ZN(new_n429));
  NAND2_X1  g228(.A1(new_n428), .A2(new_n429), .ZN(new_n430));
  INV_X1    g229(.A(new_n430), .ZN(new_n431));
  INV_X1    g230(.A(KEYINPUT76), .ZN(new_n432));
  INV_X1    g231(.A(KEYINPUT30), .ZN(new_n433));
  AND3_X1   g232(.A1(new_n369), .A2(new_n432), .A3(new_n433), .ZN(new_n434));
  AOI21_X1  g233(.A(new_n432), .B1(new_n369), .B2(new_n433), .ZN(new_n435));
  OAI21_X1  g234(.A(new_n431), .B1(new_n434), .B2(new_n435), .ZN(new_n436));
  AOI21_X1  g235(.A(new_n413), .B1(new_n427), .B2(new_n436), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n386), .A2(new_n437), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n365), .A2(new_n246), .ZN(new_n439));
  OAI211_X1 g238(.A(new_n323), .B(new_n235), .C1(new_n345), .C2(new_n352), .ZN(new_n440));
  INV_X1    g239(.A(G227gat), .ZN(new_n441));
  NOR2_X1   g240(.A1(new_n441), .A2(new_n325), .ZN(new_n442));
  NAND3_X1  g241(.A1(new_n439), .A2(new_n440), .A3(new_n442), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n443), .A2(KEYINPUT32), .ZN(new_n444));
  INV_X1    g243(.A(KEYINPUT33), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n443), .A2(new_n445), .ZN(new_n446));
  XOR2_X1   g245(.A(G15gat), .B(G43gat), .Z(new_n447));
  XNOR2_X1  g246(.A(G71gat), .B(G99gat), .ZN(new_n448));
  XNOR2_X1  g247(.A(new_n447), .B(new_n448), .ZN(new_n449));
  NAND3_X1  g248(.A1(new_n444), .A2(new_n446), .A3(new_n449), .ZN(new_n450));
  INV_X1    g249(.A(new_n449), .ZN(new_n451));
  OAI211_X1 g250(.A(new_n443), .B(KEYINPUT32), .C1(new_n445), .C2(new_n451), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n450), .A2(new_n452), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n439), .A2(new_n440), .ZN(new_n454));
  OAI21_X1  g253(.A(new_n454), .B1(new_n441), .B2(new_n325), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n455), .A2(KEYINPUT34), .ZN(new_n456));
  INV_X1    g255(.A(KEYINPUT34), .ZN(new_n457));
  OAI211_X1 g256(.A(new_n454), .B(new_n457), .C1(new_n441), .C2(new_n325), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n456), .A2(new_n458), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n453), .A2(new_n459), .ZN(new_n460));
  NAND4_X1  g259(.A1(new_n450), .A2(new_n456), .A3(new_n458), .A4(new_n452), .ZN(new_n461));
  NAND3_X1  g260(.A1(new_n460), .A2(KEYINPUT74), .A3(new_n461), .ZN(new_n462));
  INV_X1    g261(.A(KEYINPUT74), .ZN(new_n463));
  NAND3_X1  g262(.A1(new_n453), .A2(new_n459), .A3(new_n463), .ZN(new_n464));
  XNOR2_X1  g263(.A(KEYINPUT73), .B(KEYINPUT36), .ZN(new_n465));
  NAND3_X1  g264(.A1(new_n462), .A2(new_n464), .A3(new_n465), .ZN(new_n466));
  INV_X1    g265(.A(KEYINPUT72), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n460), .A2(new_n467), .ZN(new_n468));
  NAND3_X1  g267(.A1(new_n453), .A2(new_n459), .A3(KEYINPUT72), .ZN(new_n469));
  NAND4_X1  g268(.A1(new_n468), .A2(KEYINPUT36), .A3(new_n469), .A4(new_n461), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n369), .A2(new_n433), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n471), .A2(KEYINPUT76), .ZN(new_n472));
  NAND3_X1  g271(.A1(new_n369), .A2(new_n432), .A3(new_n433), .ZN(new_n473));
  AOI21_X1  g272(.A(new_n430), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n474), .A2(new_n277), .ZN(new_n475));
  AOI22_X1  g274(.A1(new_n466), .A2(new_n470), .B1(new_n475), .B2(new_n413), .ZN(new_n476));
  NOR2_X1   g275(.A1(new_n278), .A2(new_n436), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n462), .A2(new_n464), .ZN(new_n478));
  INV_X1    g277(.A(KEYINPUT35), .ZN(new_n479));
  INV_X1    g278(.A(new_n412), .ZN(new_n480));
  AOI21_X1  g279(.A(new_n406), .B1(new_n480), .B2(new_n410), .ZN(new_n481));
  NAND4_X1  g280(.A1(new_n477), .A2(new_n478), .A3(new_n479), .A4(new_n481), .ZN(new_n482));
  NAND4_X1  g281(.A1(new_n468), .A2(new_n481), .A3(new_n469), .A4(new_n461), .ZN(new_n483));
  OAI21_X1  g282(.A(KEYINPUT35), .B1(new_n483), .B2(new_n475), .ZN(new_n484));
  AOI22_X1  g283(.A1(new_n438), .A2(new_n476), .B1(new_n482), .B2(new_n484), .ZN(new_n485));
  XNOR2_X1  g284(.A(G113gat), .B(G141gat), .ZN(new_n486));
  XNOR2_X1  g285(.A(new_n486), .B(G197gat), .ZN(new_n487));
  XOR2_X1   g286(.A(KEYINPUT11), .B(G169gat), .Z(new_n488));
  XNOR2_X1  g287(.A(new_n487), .B(new_n488), .ZN(new_n489));
  XOR2_X1   g288(.A(new_n489), .B(KEYINPUT12), .Z(new_n490));
  NAND2_X1  g289(.A1(G229gat), .A2(G233gat), .ZN(new_n491));
  XOR2_X1   g290(.A(new_n491), .B(KEYINPUT13), .Z(new_n492));
  XNOR2_X1  g291(.A(G15gat), .B(G22gat), .ZN(new_n493));
  INV_X1    g292(.A(G1gat), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n494), .A2(KEYINPUT16), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n493), .A2(new_n495), .ZN(new_n496));
  INV_X1    g295(.A(new_n496), .ZN(new_n497));
  INV_X1    g296(.A(KEYINPUT88), .ZN(new_n498));
  OAI21_X1  g297(.A(new_n498), .B1(new_n493), .B2(G1gat), .ZN(new_n499));
  OAI21_X1  g298(.A(G8gat), .B1(new_n497), .B2(new_n499), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n408), .A2(G15gat), .ZN(new_n501));
  INV_X1    g300(.A(G15gat), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n502), .A2(G22gat), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n501), .A2(new_n503), .ZN(new_n504));
  AOI21_X1  g303(.A(KEYINPUT88), .B1(new_n504), .B2(new_n494), .ZN(new_n505));
  INV_X1    g304(.A(G8gat), .ZN(new_n506));
  NAND3_X1  g305(.A1(new_n505), .A2(new_n506), .A3(new_n496), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n500), .A2(new_n507), .ZN(new_n508));
  INV_X1    g307(.A(G29gat), .ZN(new_n509));
  INV_X1    g308(.A(G36gat), .ZN(new_n510));
  NAND3_X1  g309(.A1(new_n509), .A2(new_n510), .A3(KEYINPUT14), .ZN(new_n511));
  INV_X1    g310(.A(KEYINPUT14), .ZN(new_n512));
  OAI21_X1  g311(.A(new_n512), .B1(G29gat), .B2(G36gat), .ZN(new_n513));
  AND2_X1   g312(.A1(new_n511), .A2(new_n513), .ZN(new_n514));
  INV_X1    g313(.A(KEYINPUT15), .ZN(new_n515));
  INV_X1    g314(.A(G43gat), .ZN(new_n516));
  NOR2_X1   g315(.A1(new_n516), .A2(G50gat), .ZN(new_n517));
  NOR2_X1   g316(.A1(new_n401), .A2(G43gat), .ZN(new_n518));
  OAI21_X1  g317(.A(new_n515), .B1(new_n517), .B2(new_n518), .ZN(new_n519));
  NAND2_X1  g318(.A1(G29gat), .A2(G36gat), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n520), .A2(KEYINPUT87), .ZN(new_n521));
  INV_X1    g320(.A(KEYINPUT87), .ZN(new_n522));
  NAND3_X1  g321(.A1(new_n522), .A2(G29gat), .A3(G36gat), .ZN(new_n523));
  AND2_X1   g322(.A1(new_n521), .A2(new_n523), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n401), .A2(G43gat), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n516), .A2(G50gat), .ZN(new_n526));
  NAND3_X1  g325(.A1(new_n525), .A2(new_n526), .A3(KEYINPUT15), .ZN(new_n527));
  NAND4_X1  g326(.A1(new_n514), .A2(new_n519), .A3(new_n524), .A4(new_n527), .ZN(new_n528));
  NAND3_X1  g327(.A1(new_n511), .A2(new_n513), .A3(new_n520), .ZN(new_n529));
  NOR2_X1   g328(.A1(new_n517), .A2(new_n518), .ZN(new_n530));
  NAND3_X1  g329(.A1(new_n529), .A2(new_n530), .A3(KEYINPUT15), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n528), .A2(new_n531), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n508), .A2(new_n532), .ZN(new_n533));
  INV_X1    g332(.A(new_n533), .ZN(new_n534));
  NOR2_X1   g333(.A1(new_n508), .A2(new_n532), .ZN(new_n535));
  OAI21_X1  g334(.A(new_n492), .B1(new_n534), .B2(new_n535), .ZN(new_n536));
  INV_X1    g335(.A(new_n491), .ZN(new_n537));
  INV_X1    g336(.A(KEYINPUT89), .ZN(new_n538));
  AOI21_X1  g337(.A(new_n538), .B1(new_n508), .B2(new_n532), .ZN(new_n539));
  INV_X1    g338(.A(KEYINPUT17), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n519), .A2(new_n527), .ZN(new_n541));
  NAND4_X1  g340(.A1(new_n511), .A2(new_n521), .A3(new_n513), .A4(new_n523), .ZN(new_n542));
  OAI211_X1 g341(.A(new_n531), .B(new_n540), .C1(new_n541), .C2(new_n542), .ZN(new_n543));
  INV_X1    g342(.A(new_n543), .ZN(new_n544));
  AOI21_X1  g343(.A(new_n540), .B1(new_n528), .B2(new_n531), .ZN(new_n545));
  NOR2_X1   g344(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  OAI21_X1  g345(.A(new_n539), .B1(new_n546), .B2(new_n508), .ZN(new_n547));
  AND2_X1   g346(.A1(new_n500), .A2(new_n507), .ZN(new_n548));
  OAI211_X1 g347(.A(new_n548), .B(new_n538), .C1(new_n544), .C2(new_n545), .ZN(new_n549));
  AOI21_X1  g348(.A(new_n537), .B1(new_n547), .B2(new_n549), .ZN(new_n550));
  OAI21_X1  g349(.A(new_n536), .B1(new_n550), .B2(KEYINPUT18), .ZN(new_n551));
  INV_X1    g350(.A(KEYINPUT18), .ZN(new_n552));
  AOI211_X1 g351(.A(new_n552), .B(new_n537), .C1(new_n547), .C2(new_n549), .ZN(new_n553));
  OAI21_X1  g352(.A(new_n490), .B1(new_n551), .B2(new_n553), .ZN(new_n554));
  INV_X1    g353(.A(KEYINPUT90), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n533), .A2(KEYINPUT89), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n532), .A2(KEYINPUT17), .ZN(new_n557));
  AOI21_X1  g356(.A(new_n508), .B1(new_n557), .B2(new_n543), .ZN(new_n558));
  OAI21_X1  g357(.A(new_n549), .B1(new_n556), .B2(new_n558), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n559), .A2(new_n491), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n560), .A2(new_n552), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n550), .A2(KEYINPUT18), .ZN(new_n562));
  INV_X1    g361(.A(new_n490), .ZN(new_n563));
  NAND4_X1  g362(.A1(new_n561), .A2(new_n562), .A3(new_n563), .A4(new_n536), .ZN(new_n564));
  NAND3_X1  g363(.A1(new_n554), .A2(new_n555), .A3(new_n564), .ZN(new_n565));
  OAI211_X1 g364(.A(KEYINPUT90), .B(new_n490), .C1(new_n551), .C2(new_n553), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  INV_X1    g366(.A(KEYINPUT99), .ZN(new_n568));
  NAND2_X1  g367(.A1(G230gat), .A2(G233gat), .ZN(new_n569));
  INV_X1    g368(.A(new_n569), .ZN(new_n570));
  INV_X1    g369(.A(KEYINPUT91), .ZN(new_n571));
  INV_X1    g370(.A(KEYINPUT9), .ZN(new_n572));
  INV_X1    g371(.A(G57gat), .ZN(new_n573));
  NAND2_X1  g372(.A1(new_n573), .A2(G64gat), .ZN(new_n574));
  INV_X1    g373(.A(G64gat), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n575), .A2(G57gat), .ZN(new_n576));
  AOI21_X1  g375(.A(new_n572), .B1(new_n574), .B2(new_n576), .ZN(new_n577));
  OR2_X1    g376(.A1(G71gat), .A2(G78gat), .ZN(new_n578));
  NAND2_X1  g377(.A1(G71gat), .A2(G78gat), .ZN(new_n579));
  NAND2_X1  g378(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  OAI21_X1  g379(.A(new_n571), .B1(new_n577), .B2(new_n580), .ZN(new_n581));
  INV_X1    g380(.A(new_n579), .ZN(new_n582));
  NOR2_X1   g381(.A1(G71gat), .A2(G78gat), .ZN(new_n583));
  NOR2_X1   g382(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  XNOR2_X1  g383(.A(G57gat), .B(G64gat), .ZN(new_n585));
  OAI211_X1 g384(.A(new_n584), .B(KEYINPUT91), .C1(new_n585), .C2(new_n572), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n581), .A2(new_n586), .ZN(new_n587));
  INV_X1    g386(.A(KEYINPUT92), .ZN(new_n588));
  OAI21_X1  g387(.A(new_n588), .B1(new_n575), .B2(G57gat), .ZN(new_n589));
  INV_X1    g388(.A(KEYINPUT93), .ZN(new_n590));
  OAI21_X1  g389(.A(new_n590), .B1(new_n573), .B2(G64gat), .ZN(new_n591));
  NAND3_X1  g390(.A1(new_n573), .A2(KEYINPUT92), .A3(G64gat), .ZN(new_n592));
  NAND3_X1  g391(.A1(new_n575), .A2(KEYINPUT93), .A3(G57gat), .ZN(new_n593));
  NAND4_X1  g392(.A1(new_n589), .A2(new_n591), .A3(new_n592), .A4(new_n593), .ZN(new_n594));
  INV_X1    g393(.A(KEYINPUT94), .ZN(new_n595));
  OAI21_X1  g394(.A(new_n579), .B1(new_n578), .B2(new_n572), .ZN(new_n596));
  AND3_X1   g395(.A1(new_n594), .A2(new_n595), .A3(new_n596), .ZN(new_n597));
  AOI21_X1  g396(.A(new_n595), .B1(new_n594), .B2(new_n596), .ZN(new_n598));
  OAI21_X1  g397(.A(new_n587), .B1(new_n597), .B2(new_n598), .ZN(new_n599));
  NAND2_X1  g398(.A1(G85gat), .A2(G92gat), .ZN(new_n600));
  NAND2_X1  g399(.A1(new_n600), .A2(KEYINPUT7), .ZN(new_n601));
  INV_X1    g400(.A(KEYINPUT7), .ZN(new_n602));
  NAND3_X1  g401(.A1(new_n602), .A2(G85gat), .A3(G92gat), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n601), .A2(new_n603), .ZN(new_n604));
  XNOR2_X1  g403(.A(G99gat), .B(G106gat), .ZN(new_n605));
  NAND2_X1  g404(.A1(G99gat), .A2(G106gat), .ZN(new_n606));
  INV_X1    g405(.A(G85gat), .ZN(new_n607));
  INV_X1    g406(.A(G92gat), .ZN(new_n608));
  AOI22_X1  g407(.A1(KEYINPUT8), .A2(new_n606), .B1(new_n607), .B2(new_n608), .ZN(new_n609));
  AND3_X1   g408(.A1(new_n604), .A2(new_n605), .A3(new_n609), .ZN(new_n610));
  AOI21_X1  g409(.A(new_n605), .B1(new_n604), .B2(new_n609), .ZN(new_n611));
  NOR2_X1   g410(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  INV_X1    g411(.A(new_n612), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n599), .A2(new_n613), .ZN(new_n614));
  INV_X1    g413(.A(KEYINPUT10), .ZN(new_n615));
  OAI211_X1 g414(.A(new_n612), .B(new_n587), .C1(new_n598), .C2(new_n597), .ZN(new_n616));
  NAND3_X1  g415(.A1(new_n614), .A2(new_n615), .A3(new_n616), .ZN(new_n617));
  INV_X1    g416(.A(new_n611), .ZN(new_n618));
  NAND3_X1  g417(.A1(new_n604), .A2(new_n609), .A3(new_n605), .ZN(new_n619));
  NAND3_X1  g418(.A1(new_n618), .A2(KEYINPUT97), .A3(new_n619), .ZN(new_n620));
  INV_X1    g419(.A(KEYINPUT97), .ZN(new_n621));
  OAI21_X1  g420(.A(new_n621), .B1(new_n610), .B2(new_n611), .ZN(new_n622));
  NAND2_X1  g421(.A1(new_n620), .A2(new_n622), .ZN(new_n623));
  OR2_X1    g422(.A1(new_n597), .A2(new_n598), .ZN(new_n624));
  NAND4_X1  g423(.A1(new_n623), .A2(new_n624), .A3(KEYINPUT10), .A4(new_n587), .ZN(new_n625));
  AOI21_X1  g424(.A(new_n570), .B1(new_n617), .B2(new_n625), .ZN(new_n626));
  AOI21_X1  g425(.A(new_n569), .B1(new_n614), .B2(new_n616), .ZN(new_n627));
  NOR2_X1   g426(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  XNOR2_X1  g427(.A(G120gat), .B(G148gat), .ZN(new_n629));
  XNOR2_X1  g428(.A(G176gat), .B(G204gat), .ZN(new_n630));
  XOR2_X1   g429(.A(new_n629), .B(new_n630), .Z(new_n631));
  AOI21_X1  g430(.A(new_n568), .B1(new_n628), .B2(new_n631), .ZN(new_n632));
  INV_X1    g431(.A(new_n631), .ZN(new_n633));
  NOR4_X1   g432(.A1(new_n626), .A2(KEYINPUT99), .A3(new_n627), .A4(new_n633), .ZN(new_n634));
  OAI22_X1  g433(.A1(new_n632), .A2(new_n634), .B1(new_n628), .B2(new_n631), .ZN(new_n635));
  INV_X1    g434(.A(KEYINPUT21), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n599), .A2(new_n636), .ZN(new_n637));
  NAND2_X1  g436(.A1(G231gat), .A2(G233gat), .ZN(new_n638));
  XNOR2_X1  g437(.A(new_n637), .B(new_n638), .ZN(new_n639));
  XOR2_X1   g438(.A(G127gat), .B(G155gat), .Z(new_n640));
  XNOR2_X1  g439(.A(new_n640), .B(KEYINPUT20), .ZN(new_n641));
  XNOR2_X1  g440(.A(new_n639), .B(new_n641), .ZN(new_n642));
  XNOR2_X1  g441(.A(G183gat), .B(G211gat), .ZN(new_n643));
  OR2_X1    g442(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n642), .A2(new_n643), .ZN(new_n645));
  NAND2_X1  g444(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  OAI21_X1  g445(.A(new_n548), .B1(new_n599), .B2(new_n636), .ZN(new_n647));
  XOR2_X1   g446(.A(KEYINPUT95), .B(KEYINPUT19), .Z(new_n648));
  XNOR2_X1  g447(.A(new_n647), .B(new_n648), .ZN(new_n649));
  INV_X1    g448(.A(new_n649), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n646), .A2(new_n650), .ZN(new_n651));
  NAND3_X1  g450(.A1(new_n644), .A2(new_n649), .A3(new_n645), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  OR2_X1    g452(.A1(new_n546), .A2(new_n623), .ZN(new_n654));
  NAND3_X1  g453(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n655));
  XNOR2_X1  g454(.A(G190gat), .B(G218gat), .ZN(new_n656));
  INV_X1    g455(.A(new_n656), .ZN(new_n657));
  OAI21_X1  g456(.A(new_n655), .B1(new_n657), .B2(KEYINPUT98), .ZN(new_n658));
  AOI21_X1  g457(.A(new_n658), .B1(new_n623), .B2(new_n532), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n654), .A2(new_n659), .ZN(new_n660));
  NAND3_X1  g459(.A1(new_n660), .A2(KEYINPUT98), .A3(new_n657), .ZN(new_n661));
  NAND2_X1  g460(.A1(new_n657), .A2(KEYINPUT98), .ZN(new_n662));
  NAND3_X1  g461(.A1(new_n654), .A2(new_n662), .A3(new_n659), .ZN(new_n663));
  NAND2_X1  g462(.A1(new_n661), .A2(new_n663), .ZN(new_n664));
  AOI21_X1  g463(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n665));
  XOR2_X1   g464(.A(new_n665), .B(KEYINPUT96), .Z(new_n666));
  XNOR2_X1  g465(.A(G134gat), .B(G162gat), .ZN(new_n667));
  XNOR2_X1  g466(.A(new_n666), .B(new_n667), .ZN(new_n668));
  INV_X1    g467(.A(new_n668), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n664), .A2(new_n669), .ZN(new_n670));
  NAND3_X1  g469(.A1(new_n661), .A2(new_n668), .A3(new_n663), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  INV_X1    g471(.A(new_n672), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n653), .A2(new_n673), .ZN(new_n674));
  NOR4_X1   g473(.A1(new_n485), .A2(new_n567), .A3(new_n635), .A4(new_n674), .ZN(new_n675));
  NAND2_X1  g474(.A1(new_n675), .A2(new_n278), .ZN(new_n676));
  XNOR2_X1  g475(.A(new_n676), .B(G1gat), .ZN(G1324gat));
  XNOR2_X1  g476(.A(KEYINPUT100), .B(KEYINPUT16), .ZN(new_n678));
  XNOR2_X1  g477(.A(new_n678), .B(new_n506), .ZN(new_n679));
  AND3_X1   g478(.A1(new_n675), .A2(new_n436), .A3(new_n679), .ZN(new_n680));
  AOI21_X1  g479(.A(new_n506), .B1(new_n675), .B2(new_n436), .ZN(new_n681));
  OAI21_X1  g480(.A(KEYINPUT42), .B1(new_n680), .B2(new_n681), .ZN(new_n682));
  OAI21_X1  g481(.A(new_n682), .B1(KEYINPUT42), .B2(new_n680), .ZN(G1325gat));
  NAND3_X1  g482(.A1(new_n675), .A2(new_n502), .A3(new_n478), .ZN(new_n684));
  AND2_X1   g483(.A1(new_n466), .A2(new_n470), .ZN(new_n685));
  AND2_X1   g484(.A1(new_n675), .A2(new_n685), .ZN(new_n686));
  OAI21_X1  g485(.A(new_n684), .B1(new_n686), .B2(new_n502), .ZN(G1326gat));
  NAND2_X1  g486(.A1(new_n675), .A2(new_n413), .ZN(new_n688));
  XNOR2_X1  g487(.A(KEYINPUT43), .B(G22gat), .ZN(new_n689));
  XNOR2_X1  g488(.A(new_n688), .B(new_n689), .ZN(G1327gat));
  NAND2_X1  g489(.A1(new_n476), .A2(new_n438), .ZN(new_n691));
  NAND2_X1  g490(.A1(new_n482), .A2(new_n484), .ZN(new_n692));
  AOI21_X1  g491(.A(new_n673), .B1(new_n691), .B2(new_n692), .ZN(new_n693));
  NOR3_X1   g492(.A1(new_n653), .A2(new_n567), .A3(new_n635), .ZN(new_n694));
  AND2_X1   g493(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  NAND3_X1  g494(.A1(new_n695), .A2(new_n509), .A3(new_n278), .ZN(new_n696));
  XNOR2_X1  g495(.A(new_n696), .B(KEYINPUT45), .ZN(new_n697));
  INV_X1    g496(.A(KEYINPUT44), .ZN(new_n698));
  OAI21_X1  g497(.A(new_n698), .B1(new_n485), .B2(new_n673), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n691), .A2(new_n692), .ZN(new_n700));
  NAND3_X1  g499(.A1(new_n700), .A2(KEYINPUT44), .A3(new_n672), .ZN(new_n701));
  AND2_X1   g500(.A1(new_n699), .A2(new_n701), .ZN(new_n702));
  XOR2_X1   g501(.A(new_n694), .B(KEYINPUT101), .Z(new_n703));
  NAND2_X1  g502(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  OAI21_X1  g503(.A(G29gat), .B1(new_n704), .B2(new_n277), .ZN(new_n705));
  NAND2_X1  g504(.A1(new_n697), .A2(new_n705), .ZN(G1328gat));
  NAND3_X1  g505(.A1(new_n695), .A2(new_n510), .A3(new_n436), .ZN(new_n707));
  XOR2_X1   g506(.A(new_n707), .B(KEYINPUT46), .Z(new_n708));
  OAI21_X1  g507(.A(G36gat), .B1(new_n704), .B2(new_n474), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n708), .A2(new_n709), .ZN(G1329gat));
  NAND4_X1  g509(.A1(new_n699), .A2(new_n701), .A3(new_n685), .A4(new_n703), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n711), .A2(G43gat), .ZN(new_n712));
  NAND3_X1  g511(.A1(new_n695), .A2(new_n516), .A3(new_n478), .ZN(new_n713));
  NAND2_X1  g512(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  AOI21_X1  g513(.A(KEYINPUT47), .B1(new_n713), .B2(KEYINPUT102), .ZN(new_n715));
  XNOR2_X1  g514(.A(new_n714), .B(new_n715), .ZN(G1330gat));
  NAND4_X1  g515(.A1(new_n699), .A2(new_n701), .A3(new_n413), .A4(new_n703), .ZN(new_n717));
  NAND2_X1  g516(.A1(new_n717), .A2(G50gat), .ZN(new_n718));
  INV_X1    g517(.A(KEYINPUT103), .ZN(new_n719));
  AOI21_X1  g518(.A(KEYINPUT48), .B1(new_n718), .B2(new_n719), .ZN(new_n720));
  NAND3_X1  g519(.A1(new_n695), .A2(new_n401), .A3(new_n413), .ZN(new_n721));
  NAND2_X1  g520(.A1(new_n718), .A2(new_n721), .ZN(new_n722));
  XNOR2_X1  g521(.A(new_n720), .B(new_n722), .ZN(G1331gat));
  INV_X1    g522(.A(new_n567), .ZN(new_n724));
  NOR2_X1   g523(.A1(new_n628), .A2(new_n631), .ZN(new_n725));
  NAND2_X1  g524(.A1(new_n617), .A2(new_n625), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n726), .A2(new_n569), .ZN(new_n727));
  INV_X1    g526(.A(new_n627), .ZN(new_n728));
  NAND3_X1  g527(.A1(new_n727), .A2(new_n728), .A3(new_n631), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n729), .A2(KEYINPUT99), .ZN(new_n730));
  NAND3_X1  g529(.A1(new_n628), .A2(new_n568), .A3(new_n631), .ZN(new_n731));
  AOI21_X1  g530(.A(new_n725), .B1(new_n730), .B2(new_n731), .ZN(new_n732));
  NOR3_X1   g531(.A1(new_n674), .A2(new_n724), .A3(new_n732), .ZN(new_n733));
  NAND2_X1  g532(.A1(new_n700), .A2(new_n733), .ZN(new_n734));
  INV_X1    g533(.A(KEYINPUT104), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  NAND3_X1  g535(.A1(new_n700), .A2(KEYINPUT104), .A3(new_n733), .ZN(new_n737));
  AND2_X1   g536(.A1(new_n736), .A2(new_n737), .ZN(new_n738));
  NAND2_X1  g537(.A1(new_n738), .A2(new_n278), .ZN(new_n739));
  XNOR2_X1  g538(.A(KEYINPUT105), .B(G57gat), .ZN(new_n740));
  XNOR2_X1  g539(.A(new_n739), .B(new_n740), .ZN(G1332gat));
  NAND2_X1  g540(.A1(new_n738), .A2(new_n436), .ZN(new_n742));
  OAI21_X1  g541(.A(new_n742), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n743));
  XOR2_X1   g542(.A(KEYINPUT49), .B(G64gat), .Z(new_n744));
  OAI21_X1  g543(.A(new_n743), .B1(new_n742), .B2(new_n744), .ZN(G1333gat));
  INV_X1    g544(.A(G71gat), .ZN(new_n746));
  NAND3_X1  g545(.A1(new_n738), .A2(new_n746), .A3(new_n478), .ZN(new_n747));
  NAND3_X1  g546(.A1(new_n736), .A2(new_n685), .A3(new_n737), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n748), .A2(G71gat), .ZN(new_n749));
  XNOR2_X1  g548(.A(KEYINPUT106), .B(KEYINPUT50), .ZN(new_n750));
  AND3_X1   g549(.A1(new_n747), .A2(new_n749), .A3(new_n750), .ZN(new_n751));
  AOI21_X1  g550(.A(new_n750), .B1(new_n747), .B2(new_n749), .ZN(new_n752));
  NOR2_X1   g551(.A1(new_n751), .A2(new_n752), .ZN(G1334gat));
  NAND2_X1  g552(.A1(new_n738), .A2(new_n413), .ZN(new_n754));
  XNOR2_X1  g553(.A(new_n754), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g554(.A1(new_n653), .A2(new_n724), .ZN(new_n756));
  INV_X1    g555(.A(new_n756), .ZN(new_n757));
  NOR2_X1   g556(.A1(new_n757), .A2(new_n732), .ZN(new_n758));
  NAND3_X1  g557(.A1(new_n702), .A2(new_n278), .A3(new_n758), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n759), .A2(G85gat), .ZN(new_n760));
  NAND2_X1  g559(.A1(new_n693), .A2(new_n756), .ZN(new_n761));
  INV_X1    g560(.A(KEYINPUT51), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  OR2_X1    g562(.A1(new_n763), .A2(KEYINPUT107), .ZN(new_n764));
  NOR4_X1   g563(.A1(new_n485), .A2(new_n762), .A3(new_n673), .A4(new_n757), .ZN(new_n765));
  INV_X1    g564(.A(new_n765), .ZN(new_n766));
  NAND3_X1  g565(.A1(new_n766), .A2(KEYINPUT107), .A3(new_n763), .ZN(new_n767));
  NAND3_X1  g566(.A1(new_n764), .A2(new_n767), .A3(new_n635), .ZN(new_n768));
  NAND2_X1  g567(.A1(new_n278), .A2(new_n607), .ZN(new_n769));
  OAI21_X1  g568(.A(new_n760), .B1(new_n768), .B2(new_n769), .ZN(G1336gat));
  NOR3_X1   g569(.A1(new_n474), .A2(G92gat), .A3(new_n732), .ZN(new_n771));
  AND3_X1   g570(.A1(new_n764), .A2(new_n767), .A3(new_n771), .ZN(new_n772));
  NAND4_X1  g571(.A1(new_n699), .A2(new_n701), .A3(new_n436), .A4(new_n758), .ZN(new_n773));
  NAND2_X1  g572(.A1(new_n773), .A2(G92gat), .ZN(new_n774));
  INV_X1    g573(.A(KEYINPUT52), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n766), .A2(new_n763), .ZN(new_n777));
  AOI22_X1  g576(.A1(new_n777), .A2(new_n771), .B1(new_n773), .B2(G92gat), .ZN(new_n778));
  OAI22_X1  g577(.A1(new_n772), .A2(new_n776), .B1(new_n775), .B2(new_n778), .ZN(G1337gat));
  NAND3_X1  g578(.A1(new_n702), .A2(new_n685), .A3(new_n758), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n780), .A2(KEYINPUT108), .ZN(new_n781));
  XOR2_X1   g580(.A(KEYINPUT109), .B(G99gat), .Z(new_n782));
  NAND2_X1  g581(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  NOR2_X1   g582(.A1(new_n780), .A2(KEYINPUT108), .ZN(new_n784));
  INV_X1    g583(.A(new_n478), .ZN(new_n785));
  OR2_X1    g584(.A1(new_n785), .A2(new_n782), .ZN(new_n786));
  OAI22_X1  g585(.A1(new_n783), .A2(new_n784), .B1(new_n768), .B2(new_n786), .ZN(G1338gat));
  NOR3_X1   g586(.A1(new_n481), .A2(G106gat), .A3(new_n732), .ZN(new_n788));
  NAND3_X1  g587(.A1(new_n764), .A2(new_n767), .A3(new_n788), .ZN(new_n789));
  NAND4_X1  g588(.A1(new_n699), .A2(new_n701), .A3(new_n413), .A4(new_n758), .ZN(new_n790));
  AOI21_X1  g589(.A(KEYINPUT53), .B1(new_n790), .B2(G106gat), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n789), .A2(new_n791), .ZN(new_n792));
  INV_X1    g591(.A(KEYINPUT110), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n790), .A2(G106gat), .ZN(new_n794));
  AOI21_X1  g593(.A(KEYINPUT51), .B1(new_n693), .B2(new_n756), .ZN(new_n795));
  OAI21_X1  g594(.A(new_n788), .B1(new_n765), .B2(new_n795), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n794), .A2(new_n796), .ZN(new_n797));
  AOI21_X1  g596(.A(new_n793), .B1(new_n797), .B2(KEYINPUT53), .ZN(new_n798));
  INV_X1    g597(.A(KEYINPUT53), .ZN(new_n799));
  AOI211_X1 g598(.A(KEYINPUT110), .B(new_n799), .C1(new_n794), .C2(new_n796), .ZN(new_n800));
  OAI21_X1  g599(.A(new_n792), .B1(new_n798), .B2(new_n800), .ZN(G1339gat));
  INV_X1    g600(.A(G113gat), .ZN(new_n802));
  NAND4_X1  g601(.A1(new_n653), .A2(new_n567), .A3(new_n732), .A4(new_n673), .ZN(new_n803));
  NAND2_X1  g602(.A1(new_n730), .A2(new_n731), .ZN(new_n804));
  INV_X1    g603(.A(KEYINPUT55), .ZN(new_n805));
  INV_X1    g604(.A(KEYINPUT54), .ZN(new_n806));
  AOI211_X1 g605(.A(new_n805), .B(new_n631), .C1(new_n626), .C2(new_n806), .ZN(new_n807));
  NAND3_X1  g606(.A1(new_n617), .A2(new_n570), .A3(new_n625), .ZN(new_n808));
  AND4_X1   g607(.A1(KEYINPUT111), .A2(new_n727), .A3(KEYINPUT54), .A4(new_n808), .ZN(new_n809));
  AOI21_X1  g608(.A(new_n806), .B1(new_n726), .B2(new_n569), .ZN(new_n810));
  AOI21_X1  g609(.A(KEYINPUT111), .B1(new_n810), .B2(new_n808), .ZN(new_n811));
  OAI21_X1  g610(.A(new_n807), .B1(new_n809), .B2(new_n811), .ZN(new_n812));
  OAI21_X1  g611(.A(new_n633), .B1(new_n727), .B2(KEYINPUT54), .ZN(new_n813));
  NAND3_X1  g612(.A1(new_n727), .A2(KEYINPUT54), .A3(new_n808), .ZN(new_n814));
  INV_X1    g613(.A(KEYINPUT111), .ZN(new_n815));
  NAND2_X1  g614(.A1(new_n814), .A2(new_n815), .ZN(new_n816));
  NAND3_X1  g615(.A1(new_n810), .A2(KEYINPUT111), .A3(new_n808), .ZN(new_n817));
  AOI21_X1  g616(.A(new_n813), .B1(new_n816), .B2(new_n817), .ZN(new_n818));
  OAI211_X1 g617(.A(new_n804), .B(new_n812), .C1(new_n818), .C2(KEYINPUT55), .ZN(new_n819));
  OR3_X1    g618(.A1(new_n534), .A2(new_n535), .A3(new_n492), .ZN(new_n820));
  OAI21_X1  g619(.A(new_n820), .B1(new_n559), .B2(new_n491), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n821), .A2(new_n489), .ZN(new_n822));
  NAND3_X1  g621(.A1(new_n672), .A2(new_n564), .A3(new_n822), .ZN(new_n823));
  NOR2_X1   g622(.A1(new_n819), .A2(new_n823), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n564), .A2(new_n822), .ZN(new_n825));
  OAI22_X1  g624(.A1(new_n819), .A2(new_n567), .B1(new_n732), .B2(new_n825), .ZN(new_n826));
  AOI21_X1  g625(.A(new_n824), .B1(new_n826), .B2(new_n673), .ZN(new_n827));
  OAI21_X1  g626(.A(new_n803), .B1(new_n827), .B2(new_n653), .ZN(new_n828));
  AND2_X1   g627(.A1(new_n828), .A2(new_n481), .ZN(new_n829));
  NOR2_X1   g628(.A1(new_n436), .A2(new_n277), .ZN(new_n830));
  INV_X1    g629(.A(new_n830), .ZN(new_n831));
  NOR2_X1   g630(.A1(new_n831), .A2(new_n785), .ZN(new_n832));
  AND2_X1   g631(.A1(new_n829), .A2(new_n832), .ZN(new_n833));
  AOI21_X1  g632(.A(new_n802), .B1(new_n833), .B2(new_n724), .ZN(new_n834));
  XNOR2_X1  g633(.A(new_n834), .B(KEYINPUT112), .ZN(new_n835));
  AND2_X1   g634(.A1(new_n828), .A2(new_n278), .ZN(new_n836));
  NOR2_X1   g635(.A1(new_n483), .A2(new_n436), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n724), .A2(new_n802), .ZN(new_n839));
  XNOR2_X1  g638(.A(new_n839), .B(KEYINPUT113), .ZN(new_n840));
  OAI21_X1  g639(.A(new_n835), .B1(new_n838), .B2(new_n840), .ZN(G1340gat));
  NOR4_X1   g640(.A1(new_n838), .A2(new_n231), .A3(new_n232), .A4(new_n732), .ZN(new_n842));
  AOI21_X1  g641(.A(new_n230), .B1(new_n833), .B2(new_n635), .ZN(new_n843));
  OR2_X1    g642(.A1(new_n842), .A2(new_n843), .ZN(G1341gat));
  INV_X1    g643(.A(new_n833), .ZN(new_n845));
  INV_X1    g644(.A(new_n653), .ZN(new_n846));
  OAI21_X1  g645(.A(new_n219), .B1(new_n845), .B2(new_n846), .ZN(new_n847));
  OR3_X1    g646(.A1(new_n838), .A2(new_n219), .A3(new_n846), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n847), .A2(new_n848), .ZN(G1342gat));
  OR3_X1    g648(.A1(new_n838), .A2(G134gat), .A3(new_n673), .ZN(new_n850));
  OR2_X1    g649(.A1(new_n850), .A2(KEYINPUT56), .ZN(new_n851));
  OAI21_X1  g650(.A(G134gat), .B1(new_n845), .B2(new_n673), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n850), .A2(KEYINPUT56), .ZN(new_n853));
  NAND3_X1  g652(.A1(new_n851), .A2(new_n852), .A3(new_n853), .ZN(G1343gat));
  NOR3_X1   g653(.A1(new_n685), .A2(new_n481), .A3(new_n436), .ZN(new_n855));
  NOR2_X1   g654(.A1(new_n567), .A2(G141gat), .ZN(new_n856));
  XNOR2_X1  g655(.A(new_n856), .B(KEYINPUT115), .ZN(new_n857));
  NAND3_X1  g656(.A1(new_n836), .A2(new_n855), .A3(new_n857), .ZN(new_n858));
  NAND2_X1  g657(.A1(new_n858), .A2(KEYINPUT116), .ZN(new_n859));
  INV_X1    g658(.A(KEYINPUT58), .ZN(new_n860));
  INV_X1    g659(.A(KEYINPUT116), .ZN(new_n861));
  NAND4_X1  g660(.A1(new_n836), .A2(new_n861), .A3(new_n855), .A4(new_n857), .ZN(new_n862));
  AND3_X1   g661(.A1(new_n859), .A2(new_n860), .A3(new_n862), .ZN(new_n863));
  NOR2_X1   g662(.A1(new_n819), .A2(new_n567), .ZN(new_n864));
  OAI21_X1  g663(.A(KEYINPUT114), .B1(new_n732), .B2(new_n825), .ZN(new_n865));
  INV_X1    g664(.A(KEYINPUT114), .ZN(new_n866));
  NAND4_X1  g665(.A1(new_n635), .A2(new_n866), .A3(new_n564), .A4(new_n822), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n865), .A2(new_n867), .ZN(new_n868));
  OAI21_X1  g667(.A(new_n673), .B1(new_n864), .B2(new_n868), .ZN(new_n869));
  INV_X1    g668(.A(new_n824), .ZN(new_n870));
  AOI21_X1  g669(.A(new_n653), .B1(new_n869), .B2(new_n870), .ZN(new_n871));
  INV_X1    g670(.A(new_n803), .ZN(new_n872));
  NOR2_X1   g671(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  OAI21_X1  g672(.A(KEYINPUT57), .B1(new_n873), .B2(new_n481), .ZN(new_n874));
  INV_X1    g673(.A(KEYINPUT57), .ZN(new_n875));
  NAND3_X1  g674(.A1(new_n828), .A2(new_n875), .A3(new_n413), .ZN(new_n876));
  NOR2_X1   g675(.A1(new_n685), .A2(new_n831), .ZN(new_n877));
  NAND3_X1  g676(.A1(new_n874), .A2(new_n876), .A3(new_n877), .ZN(new_n878));
  OAI21_X1  g677(.A(G141gat), .B1(new_n878), .B2(new_n567), .ZN(new_n879));
  AND3_X1   g678(.A1(new_n863), .A2(KEYINPUT117), .A3(new_n879), .ZN(new_n880));
  AOI21_X1  g679(.A(KEYINPUT117), .B1(new_n863), .B2(new_n879), .ZN(new_n881));
  AND2_X1   g680(.A1(new_n879), .A2(new_n858), .ZN(new_n882));
  OAI22_X1  g681(.A1(new_n880), .A2(new_n881), .B1(new_n860), .B2(new_n882), .ZN(G1344gat));
  OAI21_X1  g682(.A(KEYINPUT118), .B1(new_n871), .B2(new_n872), .ZN(new_n884));
  INV_X1    g683(.A(KEYINPUT118), .ZN(new_n885));
  OAI211_X1 g684(.A(new_n865), .B(new_n867), .C1(new_n819), .C2(new_n567), .ZN(new_n886));
  AOI21_X1  g685(.A(new_n824), .B1(new_n886), .B2(new_n673), .ZN(new_n887));
  OAI211_X1 g686(.A(new_n885), .B(new_n803), .C1(new_n887), .C2(new_n653), .ZN(new_n888));
  NOR2_X1   g687(.A1(new_n481), .A2(KEYINPUT57), .ZN(new_n889));
  NAND3_X1  g688(.A1(new_n884), .A2(new_n888), .A3(new_n889), .ZN(new_n890));
  NAND2_X1  g689(.A1(new_n828), .A2(new_n413), .ZN(new_n891));
  NAND2_X1  g690(.A1(new_n891), .A2(KEYINPUT57), .ZN(new_n892));
  AND2_X1   g691(.A1(new_n890), .A2(new_n892), .ZN(new_n893));
  NOR3_X1   g692(.A1(new_n685), .A2(new_n732), .A3(new_n831), .ZN(new_n894));
  AOI21_X1  g693(.A(KEYINPUT119), .B1(new_n893), .B2(new_n894), .ZN(new_n895));
  NAND4_X1  g694(.A1(new_n890), .A2(KEYINPUT119), .A3(new_n892), .A4(new_n894), .ZN(new_n896));
  NAND2_X1  g695(.A1(new_n896), .A2(G148gat), .ZN(new_n897));
  OAI21_X1  g696(.A(KEYINPUT59), .B1(new_n895), .B2(new_n897), .ZN(new_n898));
  INV_X1    g697(.A(G148gat), .ZN(new_n899));
  NOR2_X1   g698(.A1(new_n899), .A2(KEYINPUT59), .ZN(new_n900));
  OAI21_X1  g699(.A(new_n900), .B1(new_n878), .B2(new_n732), .ZN(new_n901));
  NAND2_X1  g700(.A1(new_n898), .A2(new_n901), .ZN(new_n902));
  NAND2_X1  g701(.A1(new_n836), .A2(new_n855), .ZN(new_n903));
  INV_X1    g702(.A(new_n903), .ZN(new_n904));
  NAND3_X1  g703(.A1(new_n904), .A2(new_n899), .A3(new_n635), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n902), .A2(new_n905), .ZN(G1345gat));
  OAI21_X1  g705(.A(G155gat), .B1(new_n878), .B2(new_n846), .ZN(new_n907));
  NAND3_X1  g706(.A1(new_n904), .A2(new_n203), .A3(new_n653), .ZN(new_n908));
  NAND2_X1  g707(.A1(new_n907), .A2(new_n908), .ZN(G1346gat));
  NOR3_X1   g708(.A1(new_n878), .A2(new_n204), .A3(new_n673), .ZN(new_n910));
  AOI21_X1  g709(.A(G162gat), .B1(new_n904), .B2(new_n672), .ZN(new_n911));
  NOR2_X1   g710(.A1(new_n910), .A2(new_n911), .ZN(G1347gat));
  NAND2_X1  g711(.A1(new_n436), .A2(new_n277), .ZN(new_n913));
  NOR2_X1   g712(.A1(new_n785), .A2(new_n913), .ZN(new_n914));
  NAND2_X1  g713(.A1(new_n829), .A2(new_n914), .ZN(new_n915));
  NOR3_X1   g714(.A1(new_n915), .A2(new_n298), .A3(new_n567), .ZN(new_n916));
  AND2_X1   g715(.A1(new_n828), .A2(new_n277), .ZN(new_n917));
  NOR2_X1   g716(.A1(new_n483), .A2(new_n474), .ZN(new_n918));
  XNOR2_X1  g717(.A(new_n918), .B(KEYINPUT120), .ZN(new_n919));
  NAND2_X1  g718(.A1(new_n917), .A2(new_n919), .ZN(new_n920));
  NAND2_X1  g719(.A1(new_n920), .A2(KEYINPUT121), .ZN(new_n921));
  INV_X1    g720(.A(KEYINPUT121), .ZN(new_n922));
  NAND3_X1  g721(.A1(new_n917), .A2(new_n922), .A3(new_n919), .ZN(new_n923));
  NAND3_X1  g722(.A1(new_n921), .A2(new_n724), .A3(new_n923), .ZN(new_n924));
  AOI21_X1  g723(.A(new_n916), .B1(new_n924), .B2(new_n298), .ZN(G1348gat));
  NOR3_X1   g724(.A1(new_n915), .A2(new_n299), .A3(new_n732), .ZN(new_n926));
  XOR2_X1   g725(.A(new_n926), .B(KEYINPUT123), .Z(new_n927));
  NAND3_X1  g726(.A1(new_n921), .A2(new_n635), .A3(new_n923), .ZN(new_n928));
  AND3_X1   g727(.A1(new_n928), .A2(KEYINPUT122), .A3(new_n299), .ZN(new_n929));
  AOI21_X1  g728(.A(KEYINPUT122), .B1(new_n928), .B2(new_n299), .ZN(new_n930));
  NOR3_X1   g729(.A1(new_n927), .A2(new_n929), .A3(new_n930), .ZN(G1349gat));
  OAI21_X1  g730(.A(G183gat), .B1(new_n915), .B2(new_n846), .ZN(new_n932));
  NAND3_X1  g731(.A1(new_n653), .A2(new_n347), .A3(new_n349), .ZN(new_n933));
  OAI21_X1  g732(.A(new_n932), .B1(new_n920), .B2(new_n933), .ZN(new_n934));
  XNOR2_X1  g733(.A(new_n934), .B(KEYINPUT60), .ZN(G1350gat));
  OAI21_X1  g734(.A(G190gat), .B1(new_n915), .B2(new_n673), .ZN(new_n936));
  XNOR2_X1  g735(.A(new_n936), .B(KEYINPUT61), .ZN(new_n937));
  NAND4_X1  g736(.A1(new_n921), .A2(new_n309), .A3(new_n672), .A4(new_n923), .ZN(new_n938));
  NAND2_X1  g737(.A1(new_n937), .A2(new_n938), .ZN(G1351gat));
  INV_X1    g738(.A(G197gat), .ZN(new_n940));
  NOR2_X1   g739(.A1(new_n685), .A2(new_n913), .ZN(new_n941));
  AND2_X1   g740(.A1(new_n893), .A2(new_n941), .ZN(new_n942));
  AOI21_X1  g741(.A(new_n940), .B1(new_n942), .B2(new_n724), .ZN(new_n943));
  NOR3_X1   g742(.A1(new_n685), .A2(new_n481), .A3(new_n474), .ZN(new_n944));
  AND2_X1   g743(.A1(new_n917), .A2(new_n944), .ZN(new_n945));
  NAND3_X1  g744(.A1(new_n945), .A2(new_n940), .A3(new_n724), .ZN(new_n946));
  XNOR2_X1  g745(.A(new_n946), .B(KEYINPUT124), .ZN(new_n947));
  OR2_X1    g746(.A1(new_n943), .A2(new_n947), .ZN(G1352gat));
  NOR2_X1   g747(.A1(new_n732), .A2(G204gat), .ZN(new_n949));
  NAND3_X1  g748(.A1(new_n917), .A2(new_n944), .A3(new_n949), .ZN(new_n950));
  INV_X1    g749(.A(KEYINPUT62), .ZN(new_n951));
  XNOR2_X1  g750(.A(new_n950), .B(new_n951), .ZN(new_n952));
  NAND4_X1  g751(.A1(new_n890), .A2(new_n635), .A3(new_n892), .A4(new_n941), .ZN(new_n953));
  NAND2_X1  g752(.A1(new_n953), .A2(G204gat), .ZN(new_n954));
  NAND2_X1  g753(.A1(new_n952), .A2(new_n954), .ZN(new_n955));
  XNOR2_X1  g754(.A(new_n955), .B(KEYINPUT125), .ZN(G1353gat));
  NAND3_X1  g755(.A1(new_n945), .A2(new_n284), .A3(new_n653), .ZN(new_n957));
  NAND4_X1  g756(.A1(new_n890), .A2(new_n653), .A3(new_n892), .A4(new_n941), .ZN(new_n958));
  AND3_X1   g757(.A1(new_n958), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n959));
  AOI21_X1  g758(.A(KEYINPUT63), .B1(new_n958), .B2(G211gat), .ZN(new_n960));
  OAI21_X1  g759(.A(new_n957), .B1(new_n959), .B2(new_n960), .ZN(new_n961));
  INV_X1    g760(.A(KEYINPUT126), .ZN(new_n962));
  NAND2_X1  g761(.A1(new_n961), .A2(new_n962), .ZN(new_n963));
  OAI211_X1 g762(.A(KEYINPUT126), .B(new_n957), .C1(new_n959), .C2(new_n960), .ZN(new_n964));
  NAND2_X1  g763(.A1(new_n963), .A2(new_n964), .ZN(G1354gat));
  AOI21_X1  g764(.A(G218gat), .B1(new_n945), .B2(new_n672), .ZN(new_n966));
  NAND2_X1  g765(.A1(new_n672), .A2(G218gat), .ZN(new_n967));
  XNOR2_X1  g766(.A(new_n967), .B(KEYINPUT127), .ZN(new_n968));
  AOI21_X1  g767(.A(new_n966), .B1(new_n942), .B2(new_n968), .ZN(G1355gat));
endmodule


