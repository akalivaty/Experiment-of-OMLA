

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n514, n515, n516, n517,
         n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583,
         n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594,
         n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605,
         n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616,
         n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627,
         n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638,
         n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649,
         n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660,
         n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671,
         n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682,
         n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693,
         n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704,
         n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715,
         n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726,
         n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737,
         n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748,
         n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759,
         n760, n761, n762, n763, n764, n765, n766, n767, n768, n769, n770,
         n771, n772, n773, n774, n775, n776, n777, n778, n779, n780, n781,
         n782, n783, n784, n785, n786, n787, n788, n789, n790, n791, n792,
         n793, n794, n795, n796, n797, n798, n799, n800, n801, n802, n803,
         n804, n805, n806, n807, n808, n809, n810, n811, n812, n813, n814,
         n815, n816, n817, n818, n819, n820, n821, n822, n823, n824, n825,
         n826, n827, n828, n829, n830, n831, n832, n833, n834, n835, n836,
         n837, n838, n839, n840, n841, n842, n843, n844, n845, n846, n847,
         n848, n849, n850, n851, n852, n853, n854, n855, n856, n857, n858,
         n859, n860, n861, n862, n863, n864, n865, n866, n867, n868, n869,
         n870, n871, n872, n873, n874, n875, n876, n877, n878, n879, n880,
         n881, n882, n883, n884, n885, n886, n887, n888, n889, n890, n891,
         n892, n893, n894, n895, n896, n897, n898, n899, n900, n901, n902,
         n903, n904, n905, n906, n907, n908, n909, n910, n911, n912, n913,
         n914, n915, n916, n917, n918, n919, n920, n921, n922, n923, n924,
         n925, n926, n927, n928, n929, n930, n931, n932, n933, n934, n935,
         n936, n937, n938, n939, n940, n941, n942, n943, n944, n945, n946,
         n947, n948, n949, n950, n951, n952, n953, n954, n955, n956, n957,
         n958, n959, n960, n961, n962, n963, n964, n965, n966, n967, n968,
         n969, n970, n971, n972, n973, n974, n975, n976, n977, n978, n979,
         n980, n981, n982, n983, n984, n985, n986, n987, n988, n989, n990,
         n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001,
         n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011,
         n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  AND2_X1 U549 ( .A1(n735), .A2(n734), .ZN(n737) );
  XNOR2_X1 U550 ( .A(n531), .B(n530), .ZN(n635) );
  XOR2_X1 U551 ( .A(n539), .B(KEYINPUT64), .Z(n514) );
  OR2_X1 U552 ( .A1(n763), .A2(n762), .ZN(n515) );
  INV_X1 U553 ( .A(KEYINPUT28), .ZN(n703) );
  XNOR2_X1 U554 ( .A(KEYINPUT32), .B(KEYINPUT102), .ZN(n736) );
  INV_X1 U555 ( .A(n970), .ZN(n743) );
  NOR2_X2 U556 ( .A1(n767), .A2(n681), .ZN(n708) );
  AND2_X1 U557 ( .A1(n744), .A2(n743), .ZN(n745) );
  NAND2_X1 U558 ( .A1(n764), .A2(n515), .ZN(n765) );
  NOR2_X1 U559 ( .A1(n572), .A2(n571), .ZN(n573) );
  AND2_X1 U560 ( .A1(n520), .A2(G2105), .ZN(n884) );
  NOR2_X2 U561 ( .A1(G2105), .A2(n520), .ZN(n888) );
  NOR2_X1 U562 ( .A1(G651), .A2(n618), .ZN(n643) );
  NOR2_X1 U563 ( .A1(G2105), .A2(G2104), .ZN(n516) );
  XOR2_X1 U564 ( .A(KEYINPUT17), .B(n516), .Z(n517) );
  XNOR2_X1 U565 ( .A(n517), .B(KEYINPUT66), .ZN(n889) );
  NAND2_X1 U566 ( .A1(n889), .A2(G138), .ZN(n523) );
  INV_X1 U567 ( .A(G2104), .ZN(n520) );
  NAND2_X1 U568 ( .A1(G126), .A2(n884), .ZN(n519) );
  AND2_X1 U569 ( .A1(G2105), .A2(G2104), .ZN(n885) );
  NAND2_X1 U570 ( .A1(G114), .A2(n885), .ZN(n518) );
  AND2_X1 U571 ( .A1(n519), .A2(n518), .ZN(n522) );
  NAND2_X1 U572 ( .A1(G102), .A2(n888), .ZN(n521) );
  AND2_X1 U573 ( .A1(n522), .A2(n521), .ZN(n678) );
  AND2_X1 U574 ( .A1(n523), .A2(n678), .ZN(G164) );
  AND2_X1 U575 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U576 ( .A(G57), .ZN(G237) );
  INV_X1 U577 ( .A(G132), .ZN(G219) );
  NOR2_X1 U578 ( .A1(G651), .A2(G543), .ZN(n636) );
  NAND2_X1 U579 ( .A1(n636), .A2(G89), .ZN(n524) );
  XNOR2_X1 U580 ( .A(n524), .B(KEYINPUT4), .ZN(n526) );
  XOR2_X1 U581 ( .A(KEYINPUT0), .B(G543), .Z(n618) );
  INV_X1 U582 ( .A(G651), .ZN(n529) );
  NOR2_X1 U583 ( .A1(n618), .A2(n529), .ZN(n639) );
  NAND2_X1 U584 ( .A1(G76), .A2(n639), .ZN(n525) );
  NAND2_X1 U585 ( .A1(n526), .A2(n525), .ZN(n527) );
  XNOR2_X1 U586 ( .A(n527), .B(KEYINPUT5), .ZN(n536) );
  NAND2_X1 U587 ( .A1(n643), .A2(G51), .ZN(n528) );
  XNOR2_X1 U588 ( .A(n528), .B(KEYINPUT76), .ZN(n533) );
  NOR2_X1 U589 ( .A1(G543), .A2(n529), .ZN(n531) );
  XNOR2_X1 U590 ( .A(KEYINPUT67), .B(KEYINPUT1), .ZN(n530) );
  NAND2_X1 U591 ( .A1(G63), .A2(n635), .ZN(n532) );
  NAND2_X1 U592 ( .A1(n533), .A2(n532), .ZN(n534) );
  XOR2_X1 U593 ( .A(KEYINPUT6), .B(n534), .Z(n535) );
  NAND2_X1 U594 ( .A1(n536), .A2(n535), .ZN(n537) );
  XNOR2_X1 U595 ( .A(n537), .B(KEYINPUT7), .ZN(G168) );
  XOR2_X1 U596 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U597 ( .A1(G101), .A2(n888), .ZN(n538) );
  XNOR2_X1 U598 ( .A(n538), .B(KEYINPUT23), .ZN(n540) );
  NAND2_X1 U599 ( .A1(G125), .A2(n884), .ZN(n539) );
  NOR2_X1 U600 ( .A1(n540), .A2(n514), .ZN(n542) );
  NAND2_X1 U601 ( .A1(G137), .A2(n889), .ZN(n541) );
  NAND2_X1 U602 ( .A1(n542), .A2(n541), .ZN(n675) );
  NAND2_X1 U603 ( .A1(G113), .A2(n885), .ZN(n543) );
  XNOR2_X1 U604 ( .A(KEYINPUT65), .B(n543), .ZN(n673) );
  NOR2_X1 U605 ( .A1(n675), .A2(n673), .ZN(G160) );
  NAND2_X1 U606 ( .A1(G7), .A2(G661), .ZN(n544) );
  XOR2_X1 U607 ( .A(n544), .B(KEYINPUT10), .Z(n915) );
  NAND2_X1 U608 ( .A1(n915), .A2(G567), .ZN(n545) );
  XOR2_X1 U609 ( .A(KEYINPUT11), .B(n545), .Z(G234) );
  NAND2_X1 U610 ( .A1(G56), .A2(n635), .ZN(n546) );
  XOR2_X1 U611 ( .A(KEYINPUT14), .B(n546), .Z(n552) );
  NAND2_X1 U612 ( .A1(n636), .A2(G81), .ZN(n547) );
  XNOR2_X1 U613 ( .A(n547), .B(KEYINPUT12), .ZN(n549) );
  NAND2_X1 U614 ( .A1(G68), .A2(n639), .ZN(n548) );
  NAND2_X1 U615 ( .A1(n549), .A2(n548), .ZN(n550) );
  XOR2_X1 U616 ( .A(KEYINPUT13), .B(n550), .Z(n551) );
  NOR2_X1 U617 ( .A1(n552), .A2(n551), .ZN(n554) );
  NAND2_X1 U618 ( .A1(n643), .A2(G43), .ZN(n553) );
  NAND2_X1 U619 ( .A1(n554), .A2(n553), .ZN(n975) );
  INV_X1 U620 ( .A(G860), .ZN(n587) );
  OR2_X1 U621 ( .A1(n975), .A2(n587), .ZN(G153) );
  NAND2_X1 U622 ( .A1(G64), .A2(n635), .ZN(n556) );
  NAND2_X1 U623 ( .A1(G52), .A2(n643), .ZN(n555) );
  NAND2_X1 U624 ( .A1(n556), .A2(n555), .ZN(n557) );
  XNOR2_X1 U625 ( .A(KEYINPUT68), .B(n557), .ZN(n563) );
  NAND2_X1 U626 ( .A1(n639), .A2(G77), .ZN(n558) );
  XOR2_X1 U627 ( .A(KEYINPUT69), .B(n558), .Z(n560) );
  NAND2_X1 U628 ( .A1(n636), .A2(G90), .ZN(n559) );
  NAND2_X1 U629 ( .A1(n560), .A2(n559), .ZN(n561) );
  XOR2_X1 U630 ( .A(KEYINPUT9), .B(n561), .Z(n562) );
  NOR2_X1 U631 ( .A1(n563), .A2(n562), .ZN(n564) );
  XOR2_X1 U632 ( .A(KEYINPUT70), .B(n564), .Z(G301) );
  NAND2_X1 U633 ( .A1(G301), .A2(G868), .ZN(n576) );
  NAND2_X1 U634 ( .A1(G66), .A2(n635), .ZN(n566) );
  NAND2_X1 U635 ( .A1(G92), .A2(n636), .ZN(n565) );
  NAND2_X1 U636 ( .A1(n566), .A2(n565), .ZN(n567) );
  XNOR2_X1 U637 ( .A(n567), .B(KEYINPUT73), .ZN(n569) );
  NAND2_X1 U638 ( .A1(G79), .A2(n639), .ZN(n568) );
  NAND2_X1 U639 ( .A1(n569), .A2(n568), .ZN(n572) );
  NAND2_X1 U640 ( .A1(n643), .A2(G54), .ZN(n570) );
  XOR2_X1 U641 ( .A(KEYINPUT74), .B(n570), .Z(n571) );
  XNOR2_X1 U642 ( .A(n573), .B(KEYINPUT15), .ZN(n574) );
  XNOR2_X2 U643 ( .A(n574), .B(KEYINPUT75), .ZN(n980) );
  OR2_X1 U644 ( .A1(n980), .A2(G868), .ZN(n575) );
  NAND2_X1 U645 ( .A1(n576), .A2(n575), .ZN(G284) );
  NAND2_X1 U646 ( .A1(G65), .A2(n635), .ZN(n578) );
  NAND2_X1 U647 ( .A1(G53), .A2(n643), .ZN(n577) );
  NAND2_X1 U648 ( .A1(n578), .A2(n577), .ZN(n582) );
  NAND2_X1 U649 ( .A1(G91), .A2(n636), .ZN(n580) );
  NAND2_X1 U650 ( .A1(G78), .A2(n639), .ZN(n579) );
  NAND2_X1 U651 ( .A1(n580), .A2(n579), .ZN(n581) );
  NOR2_X1 U652 ( .A1(n582), .A2(n581), .ZN(n968) );
  XNOR2_X1 U653 ( .A(n968), .B(KEYINPUT71), .ZN(G299) );
  INV_X1 U654 ( .A(G868), .ZN(n590) );
  NOR2_X1 U655 ( .A1(G286), .A2(n590), .ZN(n583) );
  XOR2_X1 U656 ( .A(KEYINPUT77), .B(n583), .Z(n586) );
  NOR2_X1 U657 ( .A1(G868), .A2(G299), .ZN(n584) );
  XNOR2_X1 U658 ( .A(KEYINPUT78), .B(n584), .ZN(n585) );
  NOR2_X1 U659 ( .A1(n586), .A2(n585), .ZN(G297) );
  NAND2_X1 U660 ( .A1(n587), .A2(G559), .ZN(n588) );
  NAND2_X1 U661 ( .A1(n588), .A2(n980), .ZN(n589) );
  XNOR2_X1 U662 ( .A(n589), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U663 ( .A1(G559), .A2(n590), .ZN(n591) );
  NAND2_X1 U664 ( .A1(n980), .A2(n591), .ZN(n592) );
  XNOR2_X1 U665 ( .A(n592), .B(KEYINPUT79), .ZN(n594) );
  NOR2_X1 U666 ( .A1(n975), .A2(G868), .ZN(n593) );
  NOR2_X1 U667 ( .A1(n594), .A2(n593), .ZN(G282) );
  XOR2_X1 U668 ( .A(KEYINPUT80), .B(KEYINPUT18), .Z(n596) );
  NAND2_X1 U669 ( .A1(G123), .A2(n884), .ZN(n595) );
  XNOR2_X1 U670 ( .A(n596), .B(n595), .ZN(n603) );
  NAND2_X1 U671 ( .A1(G99), .A2(n888), .ZN(n598) );
  NAND2_X1 U672 ( .A1(G111), .A2(n885), .ZN(n597) );
  NAND2_X1 U673 ( .A1(n598), .A2(n597), .ZN(n599) );
  XNOR2_X1 U674 ( .A(n599), .B(KEYINPUT81), .ZN(n601) );
  NAND2_X1 U675 ( .A1(G135), .A2(n889), .ZN(n600) );
  NAND2_X1 U676 ( .A1(n601), .A2(n600), .ZN(n602) );
  NOR2_X1 U677 ( .A1(n603), .A2(n602), .ZN(n921) );
  XNOR2_X1 U678 ( .A(G2096), .B(n921), .ZN(n604) );
  INV_X1 U679 ( .A(G2100), .ZN(n842) );
  NAND2_X1 U680 ( .A1(n604), .A2(n842), .ZN(G156) );
  NAND2_X1 U681 ( .A1(G80), .A2(n639), .ZN(n605) );
  XNOR2_X1 U682 ( .A(n605), .B(KEYINPUT82), .ZN(n607) );
  NAND2_X1 U683 ( .A1(n635), .A2(G67), .ZN(n606) );
  NAND2_X1 U684 ( .A1(n607), .A2(n606), .ZN(n611) );
  NAND2_X1 U685 ( .A1(G93), .A2(n636), .ZN(n609) );
  NAND2_X1 U686 ( .A1(G55), .A2(n643), .ZN(n608) );
  NAND2_X1 U687 ( .A1(n609), .A2(n608), .ZN(n610) );
  NOR2_X1 U688 ( .A1(n611), .A2(n610), .ZN(n652) );
  NAND2_X1 U689 ( .A1(G559), .A2(n980), .ZN(n612) );
  XNOR2_X1 U690 ( .A(n612), .B(n975), .ZN(n655) );
  NOR2_X1 U691 ( .A1(G860), .A2(n655), .ZN(n613) );
  XOR2_X1 U692 ( .A(KEYINPUT83), .B(n613), .Z(n614) );
  XNOR2_X1 U693 ( .A(n652), .B(n614), .ZN(G145) );
  NAND2_X1 U694 ( .A1(G49), .A2(n643), .ZN(n616) );
  NAND2_X1 U695 ( .A1(G74), .A2(G651), .ZN(n615) );
  NAND2_X1 U696 ( .A1(n616), .A2(n615), .ZN(n617) );
  NOR2_X1 U697 ( .A1(n635), .A2(n617), .ZN(n620) );
  NAND2_X1 U698 ( .A1(n618), .A2(G87), .ZN(n619) );
  NAND2_X1 U699 ( .A1(n620), .A2(n619), .ZN(G288) );
  NAND2_X1 U700 ( .A1(n635), .A2(G62), .ZN(n627) );
  NAND2_X1 U701 ( .A1(G88), .A2(n636), .ZN(n622) );
  NAND2_X1 U702 ( .A1(G75), .A2(n639), .ZN(n621) );
  NAND2_X1 U703 ( .A1(n622), .A2(n621), .ZN(n625) );
  NAND2_X1 U704 ( .A1(n643), .A2(G50), .ZN(n623) );
  XOR2_X1 U705 ( .A(KEYINPUT84), .B(n623), .Z(n624) );
  NOR2_X1 U706 ( .A1(n625), .A2(n624), .ZN(n626) );
  NAND2_X1 U707 ( .A1(n627), .A2(n626), .ZN(n628) );
  XNOR2_X1 U708 ( .A(KEYINPUT85), .B(n628), .ZN(G166) );
  INV_X1 U709 ( .A(G166), .ZN(G303) );
  AND2_X1 U710 ( .A1(n635), .A2(G60), .ZN(n632) );
  NAND2_X1 U711 ( .A1(G85), .A2(n636), .ZN(n630) );
  NAND2_X1 U712 ( .A1(G72), .A2(n639), .ZN(n629) );
  NAND2_X1 U713 ( .A1(n630), .A2(n629), .ZN(n631) );
  NOR2_X1 U714 ( .A1(n632), .A2(n631), .ZN(n634) );
  NAND2_X1 U715 ( .A1(n643), .A2(G47), .ZN(n633) );
  NAND2_X1 U716 ( .A1(n634), .A2(n633), .ZN(G290) );
  NAND2_X1 U717 ( .A1(G61), .A2(n635), .ZN(n638) );
  NAND2_X1 U718 ( .A1(G86), .A2(n636), .ZN(n637) );
  NAND2_X1 U719 ( .A1(n638), .A2(n637), .ZN(n642) );
  NAND2_X1 U720 ( .A1(n639), .A2(G73), .ZN(n640) );
  XOR2_X1 U721 ( .A(KEYINPUT2), .B(n640), .Z(n641) );
  NOR2_X1 U722 ( .A1(n642), .A2(n641), .ZN(n645) );
  NAND2_X1 U723 ( .A1(n643), .A2(G48), .ZN(n644) );
  NAND2_X1 U724 ( .A1(n645), .A2(n644), .ZN(G305) );
  NOR2_X1 U725 ( .A1(G868), .A2(n652), .ZN(n646) );
  XOR2_X1 U726 ( .A(n646), .B(KEYINPUT88), .Z(n658) );
  XNOR2_X1 U727 ( .A(KEYINPUT19), .B(KEYINPUT86), .ZN(n648) );
  XNOR2_X1 U728 ( .A(G288), .B(KEYINPUT87), .ZN(n647) );
  XNOR2_X1 U729 ( .A(n648), .B(n647), .ZN(n651) );
  XOR2_X1 U730 ( .A(G303), .B(G290), .Z(n649) );
  XNOR2_X1 U731 ( .A(n649), .B(G305), .ZN(n650) );
  XNOR2_X1 U732 ( .A(n651), .B(n650), .ZN(n654) );
  XNOR2_X1 U733 ( .A(G299), .B(n652), .ZN(n653) );
  XNOR2_X1 U734 ( .A(n654), .B(n653), .ZN(n903) );
  XNOR2_X1 U735 ( .A(n903), .B(n655), .ZN(n656) );
  NAND2_X1 U736 ( .A1(G868), .A2(n656), .ZN(n657) );
  NAND2_X1 U737 ( .A1(n658), .A2(n657), .ZN(G295) );
  NAND2_X1 U738 ( .A1(G2078), .A2(G2084), .ZN(n659) );
  XOR2_X1 U739 ( .A(KEYINPUT20), .B(n659), .Z(n660) );
  NAND2_X1 U740 ( .A1(G2090), .A2(n660), .ZN(n661) );
  XNOR2_X1 U741 ( .A(KEYINPUT21), .B(n661), .ZN(n662) );
  NAND2_X1 U742 ( .A1(n662), .A2(G2072), .ZN(n663) );
  XOR2_X1 U743 ( .A(KEYINPUT89), .B(n663), .Z(G158) );
  XNOR2_X1 U744 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  XOR2_X1 U745 ( .A(KEYINPUT72), .B(G82), .Z(G220) );
  NOR2_X1 U746 ( .A1(G220), .A2(G219), .ZN(n664) );
  XOR2_X1 U747 ( .A(KEYINPUT22), .B(n664), .Z(n665) );
  NOR2_X1 U748 ( .A1(G218), .A2(n665), .ZN(n666) );
  NAND2_X1 U749 ( .A1(G96), .A2(n666), .ZN(n824) );
  NAND2_X1 U750 ( .A1(n824), .A2(G2106), .ZN(n670) );
  NAND2_X1 U751 ( .A1(G108), .A2(G120), .ZN(n667) );
  NOR2_X1 U752 ( .A1(G237), .A2(n667), .ZN(n668) );
  NAND2_X1 U753 ( .A1(G69), .A2(n668), .ZN(n825) );
  NAND2_X1 U754 ( .A1(n825), .A2(G567), .ZN(n669) );
  NAND2_X1 U755 ( .A1(n670), .A2(n669), .ZN(n857) );
  NAND2_X1 U756 ( .A1(G661), .A2(G483), .ZN(n671) );
  NOR2_X1 U757 ( .A1(n857), .A2(n671), .ZN(n823) );
  NAND2_X1 U758 ( .A1(n823), .A2(G36), .ZN(G176) );
  XNOR2_X1 U759 ( .A(G1981), .B(G305), .ZN(n986) );
  INV_X1 U760 ( .A(G40), .ZN(n672) );
  OR2_X1 U761 ( .A1(n673), .A2(n672), .ZN(n674) );
  OR2_X1 U762 ( .A1(n675), .A2(n674), .ZN(n767) );
  INV_X1 U763 ( .A(G1384), .ZN(n676) );
  AND2_X1 U764 ( .A1(G138), .A2(n676), .ZN(n677) );
  NAND2_X1 U765 ( .A1(n889), .A2(n677), .ZN(n680) );
  OR2_X1 U766 ( .A1(G1384), .A2(n678), .ZN(n679) );
  NAND2_X1 U767 ( .A1(n680), .A2(n679), .ZN(n768) );
  INV_X1 U768 ( .A(n768), .ZN(n681) );
  INV_X1 U769 ( .A(n708), .ZN(n728) );
  NOR2_X1 U770 ( .A1(G2084), .A2(n728), .ZN(n713) );
  NAND2_X1 U771 ( .A1(n713), .A2(G8), .ZN(n725) );
  NAND2_X1 U772 ( .A1(G8), .A2(n728), .ZN(n763) );
  NOR2_X1 U773 ( .A1(G1966), .A2(n763), .ZN(n723) );
  NAND2_X1 U774 ( .A1(n708), .A2(G1996), .ZN(n682) );
  XNOR2_X1 U775 ( .A(n682), .B(KEYINPUT26), .ZN(n684) );
  NAND2_X1 U776 ( .A1(n728), .A2(G1341), .ZN(n683) );
  NAND2_X1 U777 ( .A1(n684), .A2(n683), .ZN(n685) );
  NOR2_X1 U778 ( .A1(n975), .A2(n685), .ZN(n687) );
  NOR2_X1 U779 ( .A1(n687), .A2(n980), .ZN(n686) );
  XNOR2_X1 U780 ( .A(n686), .B(KEYINPUT101), .ZN(n694) );
  NAND2_X1 U781 ( .A1(n687), .A2(n980), .ZN(n692) );
  AND2_X1 U782 ( .A1(n708), .A2(G2067), .ZN(n688) );
  XOR2_X1 U783 ( .A(n688), .B(KEYINPUT100), .Z(n690) );
  NAND2_X1 U784 ( .A1(n728), .A2(G1348), .ZN(n689) );
  NAND2_X1 U785 ( .A1(n690), .A2(n689), .ZN(n691) );
  NAND2_X1 U786 ( .A1(n692), .A2(n691), .ZN(n693) );
  NAND2_X1 U787 ( .A1(n694), .A2(n693), .ZN(n701) );
  NAND2_X1 U788 ( .A1(n708), .A2(G2072), .ZN(n696) );
  INV_X1 U789 ( .A(KEYINPUT99), .ZN(n695) );
  XNOR2_X1 U790 ( .A(n696), .B(n695), .ZN(n697) );
  XNOR2_X1 U791 ( .A(n697), .B(KEYINPUT27), .ZN(n699) );
  INV_X1 U792 ( .A(G1956), .ZN(n947) );
  NOR2_X1 U793 ( .A1(n708), .A2(n947), .ZN(n698) );
  NOR2_X1 U794 ( .A1(n699), .A2(n698), .ZN(n702) );
  NAND2_X1 U795 ( .A1(n968), .A2(n702), .ZN(n700) );
  NAND2_X1 U796 ( .A1(n701), .A2(n700), .ZN(n706) );
  NOR2_X1 U797 ( .A1(n968), .A2(n702), .ZN(n704) );
  XNOR2_X1 U798 ( .A(n704), .B(n703), .ZN(n705) );
  NAND2_X1 U799 ( .A1(n706), .A2(n705), .ZN(n707) );
  XNOR2_X1 U800 ( .A(n707), .B(KEYINPUT29), .ZN(n712) );
  XOR2_X1 U801 ( .A(G2078), .B(KEYINPUT25), .Z(n1001) );
  NOR2_X1 U802 ( .A1(n1001), .A2(n728), .ZN(n710) );
  XNOR2_X1 U803 ( .A(G1961), .B(KEYINPUT98), .ZN(n952) );
  NOR2_X1 U804 ( .A1(n708), .A2(n952), .ZN(n709) );
  NOR2_X1 U805 ( .A1(n710), .A2(n709), .ZN(n717) );
  NOR2_X1 U806 ( .A1(G301), .A2(n717), .ZN(n711) );
  NOR2_X1 U807 ( .A1(n712), .A2(n711), .ZN(n722) );
  NOR2_X1 U808 ( .A1(n723), .A2(n713), .ZN(n714) );
  NAND2_X1 U809 ( .A1(G8), .A2(n714), .ZN(n715) );
  XNOR2_X1 U810 ( .A(KEYINPUT30), .B(n715), .ZN(n716) );
  NOR2_X1 U811 ( .A1(G168), .A2(n716), .ZN(n719) );
  AND2_X1 U812 ( .A1(n717), .A2(G301), .ZN(n718) );
  NOR2_X1 U813 ( .A1(n719), .A2(n718), .ZN(n720) );
  XNOR2_X1 U814 ( .A(n720), .B(KEYINPUT31), .ZN(n721) );
  NOR2_X1 U815 ( .A1(n722), .A2(n721), .ZN(n726) );
  NOR2_X1 U816 ( .A1(n723), .A2(n726), .ZN(n724) );
  NAND2_X1 U817 ( .A1(n725), .A2(n724), .ZN(n739) );
  INV_X1 U818 ( .A(n726), .ZN(n727) );
  NAND2_X1 U819 ( .A1(n727), .A2(G286), .ZN(n735) );
  INV_X1 U820 ( .A(G8), .ZN(n733) );
  NOR2_X1 U821 ( .A1(G1971), .A2(n763), .ZN(n730) );
  NOR2_X1 U822 ( .A1(G2090), .A2(n728), .ZN(n729) );
  NOR2_X1 U823 ( .A1(n730), .A2(n729), .ZN(n731) );
  NAND2_X1 U824 ( .A1(n731), .A2(G303), .ZN(n732) );
  OR2_X1 U825 ( .A1(n733), .A2(n732), .ZN(n734) );
  XNOR2_X1 U826 ( .A(n737), .B(n736), .ZN(n738) );
  NAND2_X1 U827 ( .A1(n739), .A2(n738), .ZN(n759) );
  NOR2_X1 U828 ( .A1(G1971), .A2(G303), .ZN(n740) );
  XNOR2_X1 U829 ( .A(n740), .B(KEYINPUT103), .ZN(n742) );
  INV_X1 U830 ( .A(KEYINPUT33), .ZN(n741) );
  AND2_X1 U831 ( .A1(n742), .A2(n741), .ZN(n744) );
  NOR2_X1 U832 ( .A1(G1976), .A2(G288), .ZN(n970) );
  NAND2_X1 U833 ( .A1(n759), .A2(n745), .ZN(n754) );
  INV_X1 U834 ( .A(n763), .ZN(n746) );
  NAND2_X1 U835 ( .A1(G1976), .A2(G288), .ZN(n971) );
  AND2_X1 U836 ( .A1(n746), .A2(n971), .ZN(n747) );
  NOR2_X1 U837 ( .A1(KEYINPUT33), .A2(n747), .ZN(n752) );
  NAND2_X1 U838 ( .A1(KEYINPUT33), .A2(n970), .ZN(n748) );
  XNOR2_X1 U839 ( .A(KEYINPUT104), .B(n748), .ZN(n749) );
  NOR2_X1 U840 ( .A1(n763), .A2(n749), .ZN(n750) );
  XOR2_X1 U841 ( .A(KEYINPUT105), .B(n750), .Z(n751) );
  NOR2_X1 U842 ( .A1(n752), .A2(n751), .ZN(n753) );
  AND2_X1 U843 ( .A1(n754), .A2(n753), .ZN(n755) );
  XOR2_X1 U844 ( .A(KEYINPUT106), .B(n755), .Z(n756) );
  NOR2_X1 U845 ( .A1(n986), .A2(n756), .ZN(n766) );
  NOR2_X1 U846 ( .A1(G2090), .A2(G303), .ZN(n757) );
  NAND2_X1 U847 ( .A1(G8), .A2(n757), .ZN(n758) );
  NAND2_X1 U848 ( .A1(n759), .A2(n758), .ZN(n760) );
  NAND2_X1 U849 ( .A1(n760), .A2(n763), .ZN(n764) );
  NOR2_X1 U850 ( .A1(G1981), .A2(G305), .ZN(n761) );
  XOR2_X1 U851 ( .A(n761), .B(KEYINPUT24), .Z(n762) );
  OR2_X1 U852 ( .A1(n766), .A2(n765), .ZN(n780) );
  NOR2_X1 U853 ( .A1(n768), .A2(n767), .ZN(n815) );
  NAND2_X1 U854 ( .A1(G128), .A2(n884), .ZN(n770) );
  NAND2_X1 U855 ( .A1(G116), .A2(n885), .ZN(n769) );
  NAND2_X1 U856 ( .A1(n770), .A2(n769), .ZN(n771) );
  XNOR2_X1 U857 ( .A(KEYINPUT35), .B(n771), .ZN(n777) );
  NAND2_X1 U858 ( .A1(G104), .A2(n888), .ZN(n773) );
  NAND2_X1 U859 ( .A1(G140), .A2(n889), .ZN(n772) );
  NAND2_X1 U860 ( .A1(n773), .A2(n772), .ZN(n775) );
  XOR2_X1 U861 ( .A(KEYINPUT34), .B(KEYINPUT90), .Z(n774) );
  XNOR2_X1 U862 ( .A(n775), .B(n774), .ZN(n776) );
  NAND2_X1 U863 ( .A1(n777), .A2(n776), .ZN(n778) );
  XNOR2_X1 U864 ( .A(KEYINPUT36), .B(n778), .ZN(n881) );
  XOR2_X1 U865 ( .A(KEYINPUT37), .B(G2067), .Z(n812) );
  NAND2_X1 U866 ( .A1(n881), .A2(n812), .ZN(n779) );
  XNOR2_X1 U867 ( .A(n779), .B(KEYINPUT91), .ZN(n938) );
  NAND2_X1 U868 ( .A1(n815), .A2(n938), .ZN(n810) );
  AND2_X1 U869 ( .A1(n780), .A2(n810), .ZN(n804) );
  NAND2_X1 U870 ( .A1(n888), .A2(G95), .ZN(n781) );
  XOR2_X1 U871 ( .A(KEYINPUT93), .B(n781), .Z(n783) );
  NAND2_X1 U872 ( .A1(G131), .A2(n889), .ZN(n782) );
  NAND2_X1 U873 ( .A1(n783), .A2(n782), .ZN(n784) );
  XNOR2_X1 U874 ( .A(KEYINPUT94), .B(n784), .ZN(n787) );
  NAND2_X1 U875 ( .A1(n885), .A2(G107), .ZN(n785) );
  XOR2_X1 U876 ( .A(KEYINPUT92), .B(n785), .Z(n786) );
  NOR2_X1 U877 ( .A1(n787), .A2(n786), .ZN(n789) );
  NAND2_X1 U878 ( .A1(n884), .A2(G119), .ZN(n788) );
  AND2_X1 U879 ( .A1(n789), .A2(n788), .ZN(n880) );
  XNOR2_X1 U880 ( .A(KEYINPUT95), .B(G1991), .ZN(n992) );
  NOR2_X1 U881 ( .A1(n880), .A2(n992), .ZN(n799) );
  NAND2_X1 U882 ( .A1(G129), .A2(n884), .ZN(n791) );
  NAND2_X1 U883 ( .A1(G117), .A2(n885), .ZN(n790) );
  NAND2_X1 U884 ( .A1(n791), .A2(n790), .ZN(n792) );
  XNOR2_X1 U885 ( .A(KEYINPUT96), .B(n792), .ZN(n795) );
  NAND2_X1 U886 ( .A1(n888), .A2(G105), .ZN(n793) );
  XOR2_X1 U887 ( .A(KEYINPUT38), .B(n793), .Z(n794) );
  NOR2_X1 U888 ( .A1(n795), .A2(n794), .ZN(n797) );
  NAND2_X1 U889 ( .A1(G141), .A2(n889), .ZN(n796) );
  NAND2_X1 U890 ( .A1(n797), .A2(n796), .ZN(n866) );
  AND2_X1 U891 ( .A1(n866), .A2(G1996), .ZN(n798) );
  NOR2_X1 U892 ( .A1(n799), .A2(n798), .ZN(n927) );
  INV_X1 U893 ( .A(n815), .ZN(n800) );
  NOR2_X1 U894 ( .A1(n927), .A2(n800), .ZN(n807) );
  XOR2_X1 U895 ( .A(KEYINPUT97), .B(n807), .Z(n802) );
  XNOR2_X1 U896 ( .A(G1986), .B(G290), .ZN(n974) );
  AND2_X1 U897 ( .A1(n974), .A2(n815), .ZN(n801) );
  NOR2_X1 U898 ( .A1(n802), .A2(n801), .ZN(n803) );
  NAND2_X1 U899 ( .A1(n804), .A2(n803), .ZN(n818) );
  NOR2_X1 U900 ( .A1(G1996), .A2(n866), .ZN(n917) );
  AND2_X1 U901 ( .A1(n992), .A2(n880), .ZN(n925) );
  NOR2_X1 U902 ( .A1(G1986), .A2(G290), .ZN(n805) );
  NOR2_X1 U903 ( .A1(n925), .A2(n805), .ZN(n806) );
  NOR2_X1 U904 ( .A1(n807), .A2(n806), .ZN(n808) );
  NOR2_X1 U905 ( .A1(n917), .A2(n808), .ZN(n809) );
  XNOR2_X1 U906 ( .A(n809), .B(KEYINPUT39), .ZN(n811) );
  NAND2_X1 U907 ( .A1(n811), .A2(n810), .ZN(n814) );
  NOR2_X1 U908 ( .A1(n881), .A2(n812), .ZN(n813) );
  XNOR2_X1 U909 ( .A(n813), .B(KEYINPUT107), .ZN(n935) );
  NAND2_X1 U910 ( .A1(n814), .A2(n935), .ZN(n816) );
  NAND2_X1 U911 ( .A1(n816), .A2(n815), .ZN(n817) );
  NAND2_X1 U912 ( .A1(n818), .A2(n817), .ZN(n819) );
  XNOR2_X1 U913 ( .A(KEYINPUT40), .B(n819), .ZN(G329) );
  NAND2_X1 U914 ( .A1(n915), .A2(G2106), .ZN(n820) );
  XOR2_X1 U915 ( .A(KEYINPUT111), .B(n820), .Z(G217) );
  AND2_X1 U916 ( .A1(G15), .A2(G2), .ZN(n821) );
  NAND2_X1 U917 ( .A1(G661), .A2(n821), .ZN(G259) );
  NAND2_X1 U918 ( .A1(G3), .A2(G1), .ZN(n822) );
  NAND2_X1 U919 ( .A1(n823), .A2(n822), .ZN(G188) );
  XOR2_X1 U920 ( .A(G120), .B(KEYINPUT112), .Z(G236) );
  NOR2_X1 U921 ( .A1(n825), .A2(n824), .ZN(G325) );
  XNOR2_X1 U922 ( .A(KEYINPUT113), .B(G325), .ZN(G261) );
  INV_X1 U924 ( .A(G108), .ZN(G238) );
  INV_X1 U925 ( .A(G96), .ZN(G221) );
  XNOR2_X1 U926 ( .A(KEYINPUT108), .B(G2454), .ZN(n834) );
  XNOR2_X1 U927 ( .A(G2430), .B(G2435), .ZN(n832) );
  XOR2_X1 U928 ( .A(G2451), .B(G2427), .Z(n827) );
  XNOR2_X1 U929 ( .A(G2438), .B(G2446), .ZN(n826) );
  XNOR2_X1 U930 ( .A(n827), .B(n826), .ZN(n828) );
  XOR2_X1 U931 ( .A(n828), .B(G2443), .Z(n830) );
  XNOR2_X1 U932 ( .A(G1348), .B(G1341), .ZN(n829) );
  XNOR2_X1 U933 ( .A(n830), .B(n829), .ZN(n831) );
  XNOR2_X1 U934 ( .A(n832), .B(n831), .ZN(n833) );
  XNOR2_X1 U935 ( .A(n834), .B(n833), .ZN(n835) );
  NAND2_X1 U936 ( .A1(n835), .A2(G14), .ZN(n836) );
  XOR2_X1 U937 ( .A(KEYINPUT109), .B(n836), .Z(n910) );
  XOR2_X1 U938 ( .A(KEYINPUT110), .B(n910), .Z(G401) );
  XOR2_X1 U939 ( .A(G2096), .B(KEYINPUT43), .Z(n838) );
  XNOR2_X1 U940 ( .A(G2090), .B(G2678), .ZN(n837) );
  XNOR2_X1 U941 ( .A(n838), .B(n837), .ZN(n839) );
  XOR2_X1 U942 ( .A(n839), .B(KEYINPUT42), .Z(n841) );
  XNOR2_X1 U943 ( .A(G2067), .B(G2072), .ZN(n840) );
  XNOR2_X1 U944 ( .A(n841), .B(n840), .ZN(n846) );
  XNOR2_X1 U945 ( .A(KEYINPUT114), .B(n842), .ZN(n844) );
  XNOR2_X1 U946 ( .A(G2078), .B(G2084), .ZN(n843) );
  XNOR2_X1 U947 ( .A(n844), .B(n843), .ZN(n845) );
  XNOR2_X1 U948 ( .A(n846), .B(n845), .ZN(G227) );
  XOR2_X1 U949 ( .A(G1981), .B(G1966), .Z(n848) );
  XOR2_X1 U950 ( .A(G1986), .B(n947), .Z(n847) );
  XNOR2_X1 U951 ( .A(n848), .B(n847), .ZN(n852) );
  XOR2_X1 U952 ( .A(G1961), .B(G1971), .Z(n850) );
  XNOR2_X1 U953 ( .A(G1996), .B(G1991), .ZN(n849) );
  XNOR2_X1 U954 ( .A(n850), .B(n849), .ZN(n851) );
  XOR2_X1 U955 ( .A(n852), .B(n851), .Z(n854) );
  XNOR2_X1 U956 ( .A(KEYINPUT41), .B(G2474), .ZN(n853) );
  XNOR2_X1 U957 ( .A(n854), .B(n853), .ZN(n856) );
  XOR2_X1 U958 ( .A(G1976), .B(KEYINPUT115), .Z(n855) );
  XNOR2_X1 U959 ( .A(n856), .B(n855), .ZN(G229) );
  INV_X1 U960 ( .A(n857), .ZN(G319) );
  NAND2_X1 U961 ( .A1(G124), .A2(n884), .ZN(n858) );
  XNOR2_X1 U962 ( .A(n858), .B(KEYINPUT116), .ZN(n859) );
  XNOR2_X1 U963 ( .A(n859), .B(KEYINPUT44), .ZN(n861) );
  NAND2_X1 U964 ( .A1(G100), .A2(n888), .ZN(n860) );
  NAND2_X1 U965 ( .A1(n861), .A2(n860), .ZN(n865) );
  NAND2_X1 U966 ( .A1(n885), .A2(G112), .ZN(n863) );
  NAND2_X1 U967 ( .A1(G136), .A2(n889), .ZN(n862) );
  NAND2_X1 U968 ( .A1(n863), .A2(n862), .ZN(n864) );
  NOR2_X1 U969 ( .A1(n865), .A2(n864), .ZN(G162) );
  XOR2_X1 U970 ( .A(n921), .B(G162), .Z(n868) );
  XOR2_X1 U971 ( .A(G160), .B(n866), .Z(n867) );
  XNOR2_X1 U972 ( .A(n868), .B(n867), .ZN(n879) );
  NAND2_X1 U973 ( .A1(G103), .A2(n888), .ZN(n870) );
  NAND2_X1 U974 ( .A1(G139), .A2(n889), .ZN(n869) );
  NAND2_X1 U975 ( .A1(n870), .A2(n869), .ZN(n877) );
  NAND2_X1 U976 ( .A1(n885), .A2(G115), .ZN(n871) );
  XNOR2_X1 U977 ( .A(KEYINPUT119), .B(n871), .ZN(n874) );
  NAND2_X1 U978 ( .A1(n884), .A2(G127), .ZN(n872) );
  XOR2_X1 U979 ( .A(KEYINPUT118), .B(n872), .Z(n873) );
  NOR2_X1 U980 ( .A1(n874), .A2(n873), .ZN(n875) );
  XNOR2_X1 U981 ( .A(n875), .B(KEYINPUT47), .ZN(n876) );
  NOR2_X1 U982 ( .A1(n877), .A2(n876), .ZN(n878) );
  XOR2_X1 U983 ( .A(KEYINPUT120), .B(n878), .Z(n929) );
  XOR2_X1 U984 ( .A(n879), .B(n929), .Z(n883) );
  XNOR2_X1 U985 ( .A(n881), .B(n880), .ZN(n882) );
  XNOR2_X1 U986 ( .A(n883), .B(n882), .ZN(n901) );
  XOR2_X1 U987 ( .A(KEYINPUT121), .B(KEYINPUT46), .Z(n898) );
  NAND2_X1 U988 ( .A1(G130), .A2(n884), .ZN(n887) );
  NAND2_X1 U989 ( .A1(G118), .A2(n885), .ZN(n886) );
  NAND2_X1 U990 ( .A1(n887), .A2(n886), .ZN(n895) );
  NAND2_X1 U991 ( .A1(G106), .A2(n888), .ZN(n891) );
  NAND2_X1 U992 ( .A1(G142), .A2(n889), .ZN(n890) );
  NAND2_X1 U993 ( .A1(n891), .A2(n890), .ZN(n892) );
  XNOR2_X1 U994 ( .A(KEYINPUT45), .B(n892), .ZN(n893) );
  XNOR2_X1 U995 ( .A(KEYINPUT117), .B(n893), .ZN(n894) );
  NOR2_X1 U996 ( .A1(n895), .A2(n894), .ZN(n896) );
  XNOR2_X1 U997 ( .A(KEYINPUT48), .B(n896), .ZN(n897) );
  XNOR2_X1 U998 ( .A(n898), .B(n897), .ZN(n899) );
  XNOR2_X1 U999 ( .A(G164), .B(n899), .ZN(n900) );
  XNOR2_X1 U1000 ( .A(n901), .B(n900), .ZN(n902) );
  NOR2_X1 U1001 ( .A1(G37), .A2(n902), .ZN(G395) );
  INV_X1 U1002 ( .A(G301), .ZN(G171) );
  XNOR2_X1 U1003 ( .A(n975), .B(n903), .ZN(n905) );
  XOR2_X1 U1004 ( .A(G171), .B(n980), .Z(n904) );
  XNOR2_X1 U1005 ( .A(n905), .B(n904), .ZN(n906) );
  XNOR2_X1 U1006 ( .A(n906), .B(G286), .ZN(n907) );
  NOR2_X1 U1007 ( .A1(G37), .A2(n907), .ZN(G397) );
  NOR2_X1 U1008 ( .A1(G227), .A2(G229), .ZN(n909) );
  XNOR2_X1 U1009 ( .A(KEYINPUT122), .B(KEYINPUT49), .ZN(n908) );
  XNOR2_X1 U1010 ( .A(n909), .B(n908), .ZN(n912) );
  NAND2_X1 U1011 ( .A1(G319), .A2(n910), .ZN(n911) );
  NOR2_X1 U1012 ( .A1(n912), .A2(n911), .ZN(n914) );
  NOR2_X1 U1013 ( .A1(G395), .A2(G397), .ZN(n913) );
  NAND2_X1 U1014 ( .A1(n914), .A2(n913), .ZN(G225) );
  INV_X1 U1015 ( .A(G225), .ZN(G308) );
  INV_X1 U1016 ( .A(G69), .ZN(G235) );
  INV_X1 U1017 ( .A(n915), .ZN(G223) );
  XOR2_X1 U1018 ( .A(G2090), .B(G162), .Z(n916) );
  NOR2_X1 U1019 ( .A1(n917), .A2(n916), .ZN(n918) );
  XOR2_X1 U1020 ( .A(KEYINPUT51), .B(n918), .Z(n923) );
  XNOR2_X1 U1021 ( .A(G160), .B(G2084), .ZN(n919) );
  XNOR2_X1 U1022 ( .A(n919), .B(KEYINPUT123), .ZN(n920) );
  NOR2_X1 U1023 ( .A1(n921), .A2(n920), .ZN(n922) );
  NAND2_X1 U1024 ( .A1(n923), .A2(n922), .ZN(n924) );
  NOR2_X1 U1025 ( .A1(n925), .A2(n924), .ZN(n926) );
  NAND2_X1 U1026 ( .A1(n927), .A2(n926), .ZN(n934) );
  XOR2_X1 U1027 ( .A(G164), .B(G2078), .Z(n928) );
  XNOR2_X1 U1028 ( .A(KEYINPUT124), .B(n928), .ZN(n931) );
  XNOR2_X1 U1029 ( .A(n929), .B(G2072), .ZN(n930) );
  NOR2_X1 U1030 ( .A1(n931), .A2(n930), .ZN(n932) );
  XOR2_X1 U1031 ( .A(KEYINPUT50), .B(n932), .Z(n933) );
  NOR2_X1 U1032 ( .A1(n934), .A2(n933), .ZN(n936) );
  NAND2_X1 U1033 ( .A1(n936), .A2(n935), .ZN(n937) );
  NOR2_X1 U1034 ( .A1(n938), .A2(n937), .ZN(n939) );
  XNOR2_X1 U1035 ( .A(KEYINPUT52), .B(n939), .ZN(n940) );
  INV_X1 U1036 ( .A(KEYINPUT55), .ZN(n1011) );
  NAND2_X1 U1037 ( .A1(n940), .A2(n1011), .ZN(n941) );
  NAND2_X1 U1038 ( .A1(n941), .A2(G29), .ZN(n1019) );
  XNOR2_X1 U1039 ( .A(G1348), .B(KEYINPUT59), .ZN(n942) );
  XNOR2_X1 U1040 ( .A(n942), .B(G4), .ZN(n946) );
  XNOR2_X1 U1041 ( .A(G1341), .B(G19), .ZN(n944) );
  XNOR2_X1 U1042 ( .A(G6), .B(G1981), .ZN(n943) );
  NOR2_X1 U1043 ( .A1(n944), .A2(n943), .ZN(n945) );
  NAND2_X1 U1044 ( .A1(n946), .A2(n945), .ZN(n950) );
  XNOR2_X1 U1045 ( .A(G20), .B(n947), .ZN(n948) );
  XNOR2_X1 U1046 ( .A(KEYINPUT127), .B(n948), .ZN(n949) );
  NOR2_X1 U1047 ( .A1(n950), .A2(n949), .ZN(n951) );
  XNOR2_X1 U1048 ( .A(KEYINPUT60), .B(n951), .ZN(n956) );
  XNOR2_X1 U1049 ( .A(n952), .B(G5), .ZN(n954) );
  XNOR2_X1 U1050 ( .A(G21), .B(G1966), .ZN(n953) );
  NOR2_X1 U1051 ( .A1(n954), .A2(n953), .ZN(n955) );
  NAND2_X1 U1052 ( .A1(n956), .A2(n955), .ZN(n963) );
  XNOR2_X1 U1053 ( .A(G1971), .B(G22), .ZN(n958) );
  XNOR2_X1 U1054 ( .A(G23), .B(G1976), .ZN(n957) );
  NOR2_X1 U1055 ( .A1(n958), .A2(n957), .ZN(n960) );
  XOR2_X1 U1056 ( .A(G1986), .B(G24), .Z(n959) );
  NAND2_X1 U1057 ( .A1(n960), .A2(n959), .ZN(n961) );
  XNOR2_X1 U1058 ( .A(KEYINPUT58), .B(n961), .ZN(n962) );
  NOR2_X1 U1059 ( .A1(n963), .A2(n962), .ZN(n964) );
  XNOR2_X1 U1060 ( .A(KEYINPUT61), .B(n964), .ZN(n965) );
  INV_X1 U1061 ( .A(G16), .ZN(n967) );
  NAND2_X1 U1062 ( .A1(n965), .A2(n967), .ZN(n966) );
  NAND2_X1 U1063 ( .A1(n966), .A2(G11), .ZN(n1017) );
  XOR2_X1 U1064 ( .A(KEYINPUT56), .B(n967), .Z(n991) );
  XOR2_X1 U1065 ( .A(n968), .B(G1956), .Z(n969) );
  NOR2_X1 U1066 ( .A1(n970), .A2(n969), .ZN(n972) );
  NAND2_X1 U1067 ( .A1(n972), .A2(n971), .ZN(n973) );
  NOR2_X1 U1068 ( .A1(n974), .A2(n973), .ZN(n979) );
  XOR2_X1 U1069 ( .A(G166), .B(G1971), .Z(n977) );
  XNOR2_X1 U1070 ( .A(n975), .B(G1341), .ZN(n976) );
  NOR2_X1 U1071 ( .A1(n977), .A2(n976), .ZN(n978) );
  NAND2_X1 U1072 ( .A1(n979), .A2(n978), .ZN(n984) );
  XNOR2_X1 U1073 ( .A(G1348), .B(n980), .ZN(n982) );
  XOR2_X1 U1074 ( .A(G301), .B(G1961), .Z(n981) );
  NAND2_X1 U1075 ( .A1(n982), .A2(n981), .ZN(n983) );
  NOR2_X1 U1076 ( .A1(n984), .A2(n983), .ZN(n989) );
  XOR2_X1 U1077 ( .A(G1966), .B(G168), .Z(n985) );
  NOR2_X1 U1078 ( .A1(n986), .A2(n985), .ZN(n987) );
  XOR2_X1 U1079 ( .A(KEYINPUT57), .B(n987), .Z(n988) );
  NAND2_X1 U1080 ( .A1(n989), .A2(n988), .ZN(n990) );
  NAND2_X1 U1081 ( .A1(n991), .A2(n990), .ZN(n1015) );
  XNOR2_X1 U1082 ( .A(G2090), .B(G35), .ZN(n1006) );
  XNOR2_X1 U1083 ( .A(G25), .B(n992), .ZN(n1000) );
  XNOR2_X1 U1084 ( .A(G1996), .B(G32), .ZN(n994) );
  XNOR2_X1 U1085 ( .A(G33), .B(G2072), .ZN(n993) );
  NOR2_X1 U1086 ( .A1(n994), .A2(n993), .ZN(n995) );
  NAND2_X1 U1087 ( .A1(G28), .A2(n995), .ZN(n998) );
  XOR2_X1 U1088 ( .A(KEYINPUT125), .B(G2067), .Z(n996) );
  XNOR2_X1 U1089 ( .A(G26), .B(n996), .ZN(n997) );
  NOR2_X1 U1090 ( .A1(n998), .A2(n997), .ZN(n999) );
  NAND2_X1 U1091 ( .A1(n1000), .A2(n999), .ZN(n1003) );
  XNOR2_X1 U1092 ( .A(G27), .B(n1001), .ZN(n1002) );
  NOR2_X1 U1093 ( .A1(n1003), .A2(n1002), .ZN(n1004) );
  XNOR2_X1 U1094 ( .A(KEYINPUT53), .B(n1004), .ZN(n1005) );
  NOR2_X1 U1095 ( .A1(n1006), .A2(n1005), .ZN(n1009) );
  XOR2_X1 U1096 ( .A(G2084), .B(G34), .Z(n1007) );
  XNOR2_X1 U1097 ( .A(KEYINPUT54), .B(n1007), .ZN(n1008) );
  NAND2_X1 U1098 ( .A1(n1009), .A2(n1008), .ZN(n1010) );
  XOR2_X1 U1099 ( .A(n1011), .B(n1010), .Z(n1012) );
  NOR2_X1 U1100 ( .A1(n1012), .A2(G29), .ZN(n1013) );
  XOR2_X1 U1101 ( .A(KEYINPUT126), .B(n1013), .Z(n1014) );
  NAND2_X1 U1102 ( .A1(n1015), .A2(n1014), .ZN(n1016) );
  NOR2_X1 U1103 ( .A1(n1017), .A2(n1016), .ZN(n1018) );
  NAND2_X1 U1104 ( .A1(n1019), .A2(n1018), .ZN(n1020) );
  XNOR2_X1 U1105 ( .A(KEYINPUT62), .B(n1020), .ZN(G150) );
  INV_X1 U1106 ( .A(G150), .ZN(G311) );
endmodule

