//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 0 1 0 0 1 0 0 0 1 1 1 1 0 0 0 0 1 0 0 0 0 0 1 1 1 1 0 1 0 1 0 0 0 0 1 0 1 1 0 1 1 1 0 1 0 1 0 0 0 1 0 1 1 1 1 0 0 1 1 1 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:28:02 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n723, new_n724,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n737, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n752, new_n753, new_n754, new_n755, new_n756,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n770, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n781, new_n782, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n805, new_n806, new_n807, new_n808, new_n809, new_n810,
    new_n811, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n909, new_n910,
    new_n911, new_n912, new_n913, new_n914, new_n915, new_n916, new_n917,
    new_n918, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n930, new_n931, new_n932, new_n934,
    new_n935, new_n936, new_n937, new_n938, new_n939, new_n940, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n951, new_n952, new_n953, new_n954, new_n955, new_n956,
    new_n957, new_n958, new_n959, new_n960, new_n961, new_n963, new_n964,
    new_n965, new_n966, new_n967, new_n968, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008;
  XNOR2_X1  g000(.A(KEYINPUT76), .B(G217), .ZN(new_n187));
  INV_X1    g001(.A(new_n187), .ZN(new_n188));
  INV_X1    g002(.A(G902), .ZN(new_n189));
  AOI21_X1  g003(.A(new_n188), .B1(G234), .B2(new_n189), .ZN(new_n190));
  INV_X1    g004(.A(new_n190), .ZN(new_n191));
  INV_X1    g005(.A(KEYINPUT25), .ZN(new_n192));
  OR2_X1    g006(.A1(KEYINPUT68), .A2(G119), .ZN(new_n193));
  NAND2_X1  g007(.A1(KEYINPUT68), .A2(G119), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n193), .A2(new_n194), .ZN(new_n195));
  INV_X1    g009(.A(KEYINPUT23), .ZN(new_n196));
  OAI21_X1  g010(.A(new_n195), .B1(new_n196), .B2(G128), .ZN(new_n197));
  INV_X1    g011(.A(G128), .ZN(new_n198));
  NAND3_X1  g012(.A1(new_n198), .A2(KEYINPUT23), .A3(G119), .ZN(new_n199));
  OAI211_X1 g013(.A(new_n197), .B(new_n199), .C1(KEYINPUT23), .C2(new_n198), .ZN(new_n200));
  INV_X1    g014(.A(G119), .ZN(new_n201));
  NOR2_X1   g015(.A1(new_n201), .A2(G128), .ZN(new_n202));
  AOI21_X1  g016(.A(new_n202), .B1(new_n195), .B2(G128), .ZN(new_n203));
  XOR2_X1   g017(.A(KEYINPUT24), .B(G110), .Z(new_n204));
  OAI22_X1  g018(.A1(new_n200), .A2(G110), .B1(new_n203), .B2(new_n204), .ZN(new_n205));
  XNOR2_X1  g019(.A(G125), .B(G140), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n206), .A2(KEYINPUT16), .ZN(new_n207));
  INV_X1    g021(.A(G140), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n208), .A2(G125), .ZN(new_n209));
  OR2_X1    g023(.A1(new_n209), .A2(KEYINPUT16), .ZN(new_n210));
  NAND3_X1  g024(.A1(new_n207), .A2(G146), .A3(new_n210), .ZN(new_n211));
  INV_X1    g025(.A(G125), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n212), .A2(G140), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n209), .A2(new_n213), .ZN(new_n214));
  INV_X1    g028(.A(KEYINPUT77), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n214), .A2(new_n215), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n206), .A2(KEYINPUT77), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  INV_X1    g032(.A(G146), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n219), .A2(KEYINPUT65), .ZN(new_n220));
  INV_X1    g034(.A(KEYINPUT65), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n221), .A2(G146), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n220), .A2(new_n222), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n218), .A2(new_n223), .ZN(new_n224));
  NAND3_X1  g038(.A1(new_n205), .A2(new_n211), .A3(new_n224), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n200), .A2(G110), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n207), .A2(new_n210), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n227), .A2(new_n219), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n228), .A2(new_n211), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n203), .A2(new_n204), .ZN(new_n230));
  NAND3_X1  g044(.A1(new_n226), .A2(new_n229), .A3(new_n230), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n225), .A2(new_n231), .ZN(new_n232));
  INV_X1    g046(.A(G953), .ZN(new_n233));
  NAND3_X1  g047(.A1(new_n233), .A2(G221), .A3(G234), .ZN(new_n234));
  XNOR2_X1  g048(.A(new_n234), .B(KEYINPUT22), .ZN(new_n235));
  XNOR2_X1  g049(.A(new_n235), .B(G137), .ZN(new_n236));
  XNOR2_X1  g050(.A(new_n236), .B(KEYINPUT78), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n232), .A2(new_n237), .ZN(new_n238));
  NAND3_X1  g052(.A1(new_n225), .A2(new_n236), .A3(new_n231), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n238), .A2(new_n239), .ZN(new_n240));
  OAI21_X1  g054(.A(new_n192), .B1(new_n240), .B2(G902), .ZN(new_n241));
  NAND4_X1  g055(.A1(new_n238), .A2(KEYINPUT25), .A3(new_n189), .A4(new_n239), .ZN(new_n242));
  AOI21_X1  g056(.A(new_n191), .B1(new_n241), .B2(new_n242), .ZN(new_n243));
  INV_X1    g057(.A(new_n243), .ZN(new_n244));
  NOR2_X1   g058(.A1(new_n190), .A2(G902), .ZN(new_n245));
  NAND3_X1  g059(.A1(new_n238), .A2(new_n239), .A3(new_n245), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n244), .A2(new_n246), .ZN(new_n247));
  XNOR2_X1  g061(.A(KEYINPUT2), .B(G113), .ZN(new_n248));
  INV_X1    g062(.A(G116), .ZN(new_n249));
  AOI21_X1  g063(.A(new_n249), .B1(new_n193), .B2(new_n194), .ZN(new_n250));
  NOR2_X1   g064(.A1(new_n201), .A2(G116), .ZN(new_n251));
  OAI21_X1  g065(.A(new_n248), .B1(new_n250), .B2(new_n251), .ZN(new_n252));
  XOR2_X1   g066(.A(KEYINPUT2), .B(G113), .Z(new_n253));
  AND2_X1   g067(.A1(KEYINPUT68), .A2(G119), .ZN(new_n254));
  NOR2_X1   g068(.A1(KEYINPUT68), .A2(G119), .ZN(new_n255));
  OAI21_X1  g069(.A(G116), .B1(new_n254), .B2(new_n255), .ZN(new_n256));
  INV_X1    g070(.A(new_n251), .ZN(new_n257));
  NAND3_X1  g071(.A1(new_n253), .A2(new_n256), .A3(new_n257), .ZN(new_n258));
  AND3_X1   g072(.A1(new_n252), .A2(KEYINPUT69), .A3(new_n258), .ZN(new_n259));
  AOI21_X1  g073(.A(KEYINPUT69), .B1(new_n252), .B2(new_n258), .ZN(new_n260));
  NOR2_X1   g074(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  INV_X1    g075(.A(KEYINPUT66), .ZN(new_n262));
  INV_X1    g076(.A(G134), .ZN(new_n263));
  OAI21_X1  g077(.A(new_n262), .B1(new_n263), .B2(G137), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n264), .A2(KEYINPUT11), .ZN(new_n265));
  INV_X1    g079(.A(G131), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n263), .A2(G137), .ZN(new_n267));
  INV_X1    g081(.A(KEYINPUT11), .ZN(new_n268));
  OAI211_X1 g082(.A(new_n262), .B(new_n268), .C1(new_n263), .C2(G137), .ZN(new_n269));
  NAND4_X1  g083(.A1(new_n265), .A2(new_n266), .A3(new_n267), .A4(new_n269), .ZN(new_n270));
  INV_X1    g084(.A(KEYINPUT67), .ZN(new_n271));
  OAI21_X1  g085(.A(new_n271), .B1(new_n263), .B2(G137), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n272), .A2(new_n267), .ZN(new_n273));
  NOR3_X1   g087(.A1(new_n271), .A2(new_n263), .A3(G137), .ZN(new_n274));
  OAI21_X1  g088(.A(G131), .B1(new_n273), .B2(new_n274), .ZN(new_n275));
  XNOR2_X1  g089(.A(KEYINPUT65), .B(G146), .ZN(new_n276));
  INV_X1    g090(.A(G143), .ZN(new_n277));
  OAI21_X1  g091(.A(KEYINPUT1), .B1(new_n276), .B2(new_n277), .ZN(new_n278));
  NOR2_X1   g092(.A1(new_n277), .A2(G146), .ZN(new_n279));
  INV_X1    g093(.A(new_n279), .ZN(new_n280));
  NAND3_X1  g094(.A1(new_n220), .A2(new_n222), .A3(new_n277), .ZN(new_n281));
  AOI22_X1  g095(.A1(new_n278), .A2(G128), .B1(new_n280), .B2(new_n281), .ZN(new_n282));
  AOI21_X1  g096(.A(new_n277), .B1(new_n220), .B2(new_n222), .ZN(new_n283));
  NOR2_X1   g097(.A1(new_n219), .A2(G143), .ZN(new_n284));
  NOR4_X1   g098(.A1(new_n283), .A2(KEYINPUT1), .A3(new_n198), .A4(new_n284), .ZN(new_n285));
  OAI211_X1 g099(.A(new_n270), .B(new_n275), .C1(new_n282), .C2(new_n285), .ZN(new_n286));
  NAND3_X1  g100(.A1(new_n265), .A2(new_n267), .A3(new_n269), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n287), .A2(G131), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n288), .A2(new_n270), .ZN(new_n289));
  NOR2_X1   g103(.A1(KEYINPUT0), .A2(G128), .ZN(new_n290));
  AOI21_X1  g104(.A(new_n290), .B1(new_n281), .B2(new_n280), .ZN(new_n291));
  NAND2_X1  g105(.A1(KEYINPUT0), .A2(G128), .ZN(new_n292));
  XNOR2_X1  g106(.A(new_n292), .B(KEYINPUT64), .ZN(new_n293));
  AOI21_X1  g107(.A(new_n284), .B1(new_n223), .B2(G143), .ZN(new_n294));
  INV_X1    g108(.A(new_n292), .ZN(new_n295));
  AOI22_X1  g109(.A1(new_n291), .A2(new_n293), .B1(new_n294), .B2(new_n295), .ZN(new_n296));
  INV_X1    g110(.A(KEYINPUT70), .ZN(new_n297));
  AND3_X1   g111(.A1(new_n289), .A2(new_n296), .A3(new_n297), .ZN(new_n298));
  AOI21_X1  g112(.A(new_n297), .B1(new_n289), .B2(new_n296), .ZN(new_n299));
  OAI211_X1 g113(.A(new_n261), .B(new_n286), .C1(new_n298), .C2(new_n299), .ZN(new_n300));
  INV_X1    g114(.A(G101), .ZN(new_n301));
  NOR2_X1   g115(.A1(KEYINPUT71), .A2(G237), .ZN(new_n302));
  INV_X1    g116(.A(new_n302), .ZN(new_n303));
  NAND2_X1  g117(.A1(KEYINPUT71), .A2(G237), .ZN(new_n304));
  AOI21_X1  g118(.A(G953), .B1(new_n303), .B2(new_n304), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n305), .A2(G210), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n306), .A2(KEYINPUT27), .ZN(new_n307));
  INV_X1    g121(.A(KEYINPUT26), .ZN(new_n308));
  INV_X1    g122(.A(KEYINPUT27), .ZN(new_n309));
  NAND3_X1  g123(.A1(new_n305), .A2(new_n309), .A3(G210), .ZN(new_n310));
  NAND3_X1  g124(.A1(new_n307), .A2(new_n308), .A3(new_n310), .ZN(new_n311));
  INV_X1    g125(.A(new_n311), .ZN(new_n312));
  AOI21_X1  g126(.A(new_n308), .B1(new_n307), .B2(new_n310), .ZN(new_n313));
  OAI21_X1  g127(.A(new_n301), .B1(new_n312), .B2(new_n313), .ZN(new_n314));
  INV_X1    g128(.A(new_n313), .ZN(new_n315));
  NAND3_X1  g129(.A1(new_n315), .A2(G101), .A3(new_n311), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n314), .A2(new_n316), .ZN(new_n317));
  INV_X1    g131(.A(new_n317), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n289), .A2(new_n296), .ZN(new_n319));
  INV_X1    g133(.A(KEYINPUT30), .ZN(new_n320));
  AND3_X1   g134(.A1(new_n286), .A2(new_n319), .A3(new_n320), .ZN(new_n321));
  OAI21_X1  g135(.A(new_n286), .B1(new_n298), .B2(new_n299), .ZN(new_n322));
  AOI21_X1  g136(.A(new_n321), .B1(new_n322), .B2(KEYINPUT30), .ZN(new_n323));
  OAI211_X1 g137(.A(new_n300), .B(new_n318), .C1(new_n323), .C2(new_n261), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n324), .A2(KEYINPUT31), .ZN(new_n325));
  OR2_X1    g139(.A1(new_n259), .A2(new_n260), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n319), .A2(KEYINPUT70), .ZN(new_n327));
  NAND3_X1  g141(.A1(new_n289), .A2(new_n296), .A3(new_n297), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n327), .A2(new_n328), .ZN(new_n329));
  AOI21_X1  g143(.A(new_n320), .B1(new_n329), .B2(new_n286), .ZN(new_n330));
  OAI21_X1  g144(.A(new_n326), .B1(new_n330), .B2(new_n321), .ZN(new_n331));
  INV_X1    g145(.A(KEYINPUT31), .ZN(new_n332));
  NAND4_X1  g146(.A1(new_n331), .A2(new_n332), .A3(new_n300), .A4(new_n318), .ZN(new_n333));
  INV_X1    g147(.A(KEYINPUT28), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n286), .A2(new_n319), .ZN(new_n335));
  OAI21_X1  g149(.A(new_n334), .B1(new_n335), .B2(new_n326), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n336), .A2(KEYINPUT73), .ZN(new_n337));
  INV_X1    g151(.A(KEYINPUT73), .ZN(new_n338));
  OAI211_X1 g152(.A(new_n338), .B(new_n334), .C1(new_n335), .C2(new_n326), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n337), .A2(new_n339), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n335), .A2(new_n326), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n341), .A2(KEYINPUT72), .ZN(new_n342));
  INV_X1    g156(.A(KEYINPUT72), .ZN(new_n343));
  NAND3_X1  g157(.A1(new_n335), .A2(new_n326), .A3(new_n343), .ZN(new_n344));
  NAND3_X1  g158(.A1(new_n342), .A2(new_n300), .A3(new_n344), .ZN(new_n345));
  AOI21_X1  g159(.A(new_n340), .B1(KEYINPUT28), .B2(new_n345), .ZN(new_n346));
  OAI211_X1 g160(.A(new_n325), .B(new_n333), .C1(new_n346), .C2(new_n318), .ZN(new_n347));
  NOR2_X1   g161(.A1(G472), .A2(G902), .ZN(new_n348));
  AND3_X1   g162(.A1(new_n347), .A2(KEYINPUT32), .A3(new_n348), .ZN(new_n349));
  AOI21_X1  g163(.A(KEYINPUT32), .B1(new_n347), .B2(new_n348), .ZN(new_n350));
  NOR2_X1   g164(.A1(new_n349), .A2(new_n350), .ZN(new_n351));
  INV_X1    g165(.A(KEYINPUT74), .ZN(new_n352));
  INV_X1    g166(.A(new_n300), .ZN(new_n353));
  INV_X1    g167(.A(new_n321), .ZN(new_n354));
  INV_X1    g168(.A(new_n270), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n278), .A2(G128), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n281), .A2(new_n280), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  NOR2_X1   g172(.A1(new_n221), .A2(G146), .ZN(new_n359));
  NOR2_X1   g173(.A1(new_n219), .A2(KEYINPUT65), .ZN(new_n360));
  OAI21_X1  g174(.A(G143), .B1(new_n359), .B2(new_n360), .ZN(new_n361));
  INV_X1    g175(.A(KEYINPUT1), .ZN(new_n362));
  INV_X1    g176(.A(new_n284), .ZN(new_n363));
  NAND4_X1  g177(.A1(new_n361), .A2(new_n362), .A3(G128), .A4(new_n363), .ZN(new_n364));
  AOI21_X1  g178(.A(new_n355), .B1(new_n358), .B2(new_n364), .ZN(new_n365));
  AOI22_X1  g179(.A1(new_n327), .A2(new_n328), .B1(new_n275), .B2(new_n365), .ZN(new_n366));
  OAI21_X1  g180(.A(new_n354), .B1(new_n366), .B2(new_n320), .ZN(new_n367));
  AOI21_X1  g181(.A(new_n353), .B1(new_n367), .B2(new_n326), .ZN(new_n368));
  OAI21_X1  g182(.A(new_n352), .B1(new_n368), .B2(new_n318), .ZN(new_n369));
  INV_X1    g183(.A(KEYINPUT29), .ZN(new_n370));
  OAI21_X1  g184(.A(new_n300), .B1(new_n323), .B2(new_n261), .ZN(new_n371));
  NAND3_X1  g185(.A1(new_n371), .A2(KEYINPUT74), .A3(new_n317), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n345), .A2(KEYINPUT28), .ZN(new_n373));
  AND2_X1   g187(.A1(new_n337), .A2(new_n339), .ZN(new_n374));
  NAND3_X1  g188(.A1(new_n373), .A2(new_n374), .A3(new_n318), .ZN(new_n375));
  NAND4_X1  g189(.A1(new_n369), .A2(new_n370), .A3(new_n372), .A4(new_n375), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n322), .A2(new_n326), .ZN(new_n377));
  NAND3_X1  g191(.A1(new_n377), .A2(KEYINPUT75), .A3(new_n300), .ZN(new_n378));
  INV_X1    g192(.A(KEYINPUT75), .ZN(new_n379));
  NAND3_X1  g193(.A1(new_n322), .A2(new_n379), .A3(new_n326), .ZN(new_n380));
  NAND3_X1  g194(.A1(new_n378), .A2(KEYINPUT28), .A3(new_n380), .ZN(new_n381));
  NAND4_X1  g195(.A1(new_n381), .A2(KEYINPUT29), .A3(new_n374), .A4(new_n318), .ZN(new_n382));
  NAND3_X1  g196(.A1(new_n376), .A2(new_n382), .A3(new_n189), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n383), .A2(G472), .ZN(new_n384));
  AOI21_X1  g198(.A(new_n247), .B1(new_n351), .B2(new_n384), .ZN(new_n385));
  NOR2_X1   g199(.A1(G475), .A2(G902), .ZN(new_n386));
  XNOR2_X1  g200(.A(G113), .B(G122), .ZN(new_n387));
  INV_X1    g201(.A(G104), .ZN(new_n388));
  XNOR2_X1  g202(.A(new_n387), .B(new_n388), .ZN(new_n389));
  AND2_X1   g203(.A1(KEYINPUT71), .A2(G237), .ZN(new_n390));
  OAI211_X1 g204(.A(G214), .B(new_n233), .C1(new_n390), .C2(new_n302), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n391), .A2(new_n277), .ZN(new_n392));
  XNOR2_X1  g206(.A(KEYINPUT71), .B(G237), .ZN(new_n393));
  NAND4_X1  g207(.A1(new_n393), .A2(G143), .A3(G214), .A4(new_n233), .ZN(new_n394));
  NAND3_X1  g208(.A1(new_n392), .A2(new_n394), .A3(new_n266), .ZN(new_n395));
  INV_X1    g209(.A(KEYINPUT88), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n395), .A2(new_n396), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n392), .A2(new_n394), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n398), .A2(G131), .ZN(new_n399));
  NAND4_X1  g213(.A1(new_n392), .A2(new_n394), .A3(KEYINPUT88), .A4(new_n266), .ZN(new_n400));
  NAND3_X1  g214(.A1(new_n397), .A2(new_n399), .A3(new_n400), .ZN(new_n401));
  INV_X1    g215(.A(KEYINPUT89), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n401), .A2(new_n402), .ZN(new_n403));
  AOI21_X1  g217(.A(KEYINPUT19), .B1(new_n216), .B2(new_n217), .ZN(new_n404));
  XNOR2_X1  g218(.A(new_n206), .B(KEYINPUT87), .ZN(new_n405));
  AOI21_X1  g219(.A(new_n404), .B1(KEYINPUT19), .B2(new_n405), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n406), .A2(new_n223), .ZN(new_n407));
  NAND4_X1  g221(.A1(new_n397), .A2(new_n399), .A3(KEYINPUT89), .A4(new_n400), .ZN(new_n408));
  NAND4_X1  g222(.A1(new_n403), .A2(new_n211), .A3(new_n407), .A4(new_n408), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n405), .A2(G146), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n410), .A2(new_n224), .ZN(new_n411));
  INV_X1    g225(.A(KEYINPUT18), .ZN(new_n412));
  NOR2_X1   g226(.A1(new_n412), .A2(new_n266), .ZN(new_n413));
  OAI221_X1 g227(.A(new_n411), .B1(new_n398), .B2(new_n413), .C1(new_n412), .C2(new_n399), .ZN(new_n414));
  AOI21_X1  g228(.A(new_n389), .B1(new_n409), .B2(new_n414), .ZN(new_n415));
  INV_X1    g229(.A(KEYINPUT17), .ZN(new_n416));
  NAND4_X1  g230(.A1(new_n397), .A2(new_n399), .A3(new_n416), .A4(new_n400), .ZN(new_n417));
  INV_X1    g231(.A(new_n229), .ZN(new_n418));
  INV_X1    g232(.A(KEYINPUT90), .ZN(new_n419));
  AOI21_X1  g233(.A(new_n266), .B1(new_n392), .B2(new_n394), .ZN(new_n420));
  AOI21_X1  g234(.A(new_n419), .B1(new_n420), .B2(KEYINPUT17), .ZN(new_n421));
  AND3_X1   g235(.A1(new_n420), .A2(new_n419), .A3(KEYINPUT17), .ZN(new_n422));
  OAI211_X1 g236(.A(new_n417), .B(new_n418), .C1(new_n421), .C2(new_n422), .ZN(new_n423));
  AND3_X1   g237(.A1(new_n423), .A2(new_n389), .A3(new_n414), .ZN(new_n424));
  OAI21_X1  g238(.A(new_n386), .B1(new_n415), .B2(new_n424), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n425), .A2(KEYINPUT20), .ZN(new_n426));
  INV_X1    g240(.A(KEYINPUT20), .ZN(new_n427));
  OAI211_X1 g241(.A(new_n427), .B(new_n386), .C1(new_n415), .C2(new_n424), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n426), .A2(new_n428), .ZN(new_n429));
  INV_X1    g243(.A(G475), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n423), .A2(new_n414), .ZN(new_n431));
  INV_X1    g245(.A(new_n389), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n431), .A2(new_n432), .ZN(new_n433));
  NAND3_X1  g247(.A1(new_n423), .A2(new_n389), .A3(new_n414), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n433), .A2(new_n434), .ZN(new_n435));
  AOI21_X1  g249(.A(new_n430), .B1(new_n435), .B2(new_n189), .ZN(new_n436));
  INV_X1    g250(.A(new_n436), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n429), .A2(new_n437), .ZN(new_n438));
  INV_X1    g252(.A(KEYINPUT94), .ZN(new_n439));
  AOI21_X1  g253(.A(KEYINPUT13), .B1(new_n277), .B2(G128), .ZN(new_n440));
  NOR2_X1   g254(.A1(new_n277), .A2(G128), .ZN(new_n441));
  OAI21_X1  g255(.A(KEYINPUT91), .B1(new_n440), .B2(new_n441), .ZN(new_n442));
  NAND3_X1  g256(.A1(new_n277), .A2(KEYINPUT13), .A3(G128), .ZN(new_n443));
  INV_X1    g257(.A(KEYINPUT13), .ZN(new_n444));
  OAI21_X1  g258(.A(new_n444), .B1(new_n198), .B2(G143), .ZN(new_n445));
  INV_X1    g259(.A(KEYINPUT91), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n198), .A2(G143), .ZN(new_n447));
  NAND3_X1  g261(.A1(new_n445), .A2(new_n446), .A3(new_n447), .ZN(new_n448));
  NAND3_X1  g262(.A1(new_n442), .A2(new_n443), .A3(new_n448), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n449), .A2(G134), .ZN(new_n450));
  INV_X1    g264(.A(G122), .ZN(new_n451));
  NOR2_X1   g265(.A1(new_n451), .A2(G116), .ZN(new_n452));
  NOR2_X1   g266(.A1(new_n249), .A2(G122), .ZN(new_n453));
  OR3_X1    g267(.A1(new_n452), .A2(new_n453), .A3(G107), .ZN(new_n454));
  OAI21_X1  g268(.A(G107), .B1(new_n452), .B2(new_n453), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n277), .A2(G128), .ZN(new_n457));
  NAND3_X1  g271(.A1(new_n457), .A2(new_n447), .A3(new_n263), .ZN(new_n458));
  INV_X1    g272(.A(KEYINPUT92), .ZN(new_n459));
  XNOR2_X1  g273(.A(new_n458), .B(new_n459), .ZN(new_n460));
  NAND3_X1  g274(.A1(new_n450), .A2(new_n456), .A3(new_n460), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n457), .A2(new_n447), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n462), .A2(G134), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n463), .A2(new_n458), .ZN(new_n464));
  INV_X1    g278(.A(new_n453), .ZN(new_n465));
  INV_X1    g279(.A(KEYINPUT14), .ZN(new_n466));
  NAND3_X1  g280(.A1(new_n466), .A2(new_n249), .A3(G122), .ZN(new_n467));
  INV_X1    g281(.A(KEYINPUT93), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  OAI21_X1  g283(.A(KEYINPUT14), .B1(new_n451), .B2(G116), .ZN(new_n470));
  NAND4_X1  g284(.A1(new_n466), .A2(new_n249), .A3(KEYINPUT93), .A4(G122), .ZN(new_n471));
  AND4_X1   g285(.A1(new_n465), .A2(new_n469), .A3(new_n470), .A4(new_n471), .ZN(new_n472));
  INV_X1    g286(.A(G107), .ZN(new_n473));
  OAI211_X1 g287(.A(new_n464), .B(new_n454), .C1(new_n472), .C2(new_n473), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n461), .A2(new_n474), .ZN(new_n475));
  XOR2_X1   g289(.A(KEYINPUT9), .B(G234), .Z(new_n476));
  AND3_X1   g290(.A1(new_n476), .A2(new_n233), .A3(new_n187), .ZN(new_n477));
  INV_X1    g291(.A(new_n477), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n475), .A2(new_n478), .ZN(new_n479));
  NAND3_X1  g293(.A1(new_n461), .A2(new_n474), .A3(new_n477), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  AOI21_X1  g295(.A(new_n439), .B1(new_n481), .B2(new_n189), .ZN(new_n482));
  AND3_X1   g296(.A1(new_n461), .A2(new_n474), .A3(new_n477), .ZN(new_n483));
  AOI21_X1  g297(.A(new_n477), .B1(new_n461), .B2(new_n474), .ZN(new_n484));
  OAI211_X1 g298(.A(new_n439), .B(new_n189), .C1(new_n483), .C2(new_n484), .ZN(new_n485));
  INV_X1    g299(.A(new_n485), .ZN(new_n486));
  INV_X1    g300(.A(G478), .ZN(new_n487));
  OAI22_X1  g301(.A1(new_n482), .A2(new_n486), .B1(KEYINPUT15), .B2(new_n487), .ZN(new_n488));
  INV_X1    g302(.A(KEYINPUT95), .ZN(new_n489));
  NOR2_X1   g303(.A1(new_n487), .A2(KEYINPUT15), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n485), .A2(new_n490), .ZN(new_n491));
  NAND3_X1  g305(.A1(new_n488), .A2(new_n489), .A3(new_n491), .ZN(new_n492));
  OAI21_X1  g306(.A(new_n189), .B1(new_n483), .B2(new_n484), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n493), .A2(KEYINPUT94), .ZN(new_n494));
  AOI21_X1  g308(.A(new_n490), .B1(new_n494), .B2(new_n485), .ZN(new_n495));
  INV_X1    g309(.A(new_n491), .ZN(new_n496));
  OAI21_X1  g310(.A(KEYINPUT95), .B1(new_n495), .B2(new_n496), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n492), .A2(new_n497), .ZN(new_n498));
  NOR2_X1   g312(.A1(new_n438), .A2(new_n498), .ZN(new_n499));
  INV_X1    g313(.A(KEYINPUT10), .ZN(new_n500));
  NOR3_X1   g314(.A1(new_n283), .A2(new_n198), .A3(new_n284), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n361), .A2(new_n363), .ZN(new_n502));
  OAI21_X1  g316(.A(G128), .B1(new_n279), .B2(new_n362), .ZN(new_n503));
  AOI22_X1  g317(.A1(new_n501), .A2(new_n362), .B1(new_n502), .B2(new_n503), .ZN(new_n504));
  OAI21_X1  g318(.A(KEYINPUT80), .B1(new_n388), .B2(G107), .ZN(new_n505));
  OAI21_X1  g319(.A(KEYINPUT81), .B1(new_n473), .B2(G104), .ZN(new_n506));
  INV_X1    g320(.A(KEYINPUT80), .ZN(new_n507));
  NAND3_X1  g321(.A1(new_n507), .A2(new_n473), .A3(G104), .ZN(new_n508));
  INV_X1    g322(.A(KEYINPUT81), .ZN(new_n509));
  NAND3_X1  g323(.A1(new_n509), .A2(new_n388), .A3(G107), .ZN(new_n510));
  NAND4_X1  g324(.A1(new_n505), .A2(new_n506), .A3(new_n508), .A4(new_n510), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n511), .A2(G101), .ZN(new_n512));
  NOR2_X1   g326(.A1(new_n388), .A2(G107), .ZN(new_n513));
  AND2_X1   g327(.A1(KEYINPUT79), .A2(KEYINPUT3), .ZN(new_n514));
  NOR2_X1   g328(.A1(KEYINPUT79), .A2(KEYINPUT3), .ZN(new_n515));
  OAI21_X1  g329(.A(new_n513), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  OAI22_X1  g330(.A1(new_n388), .A2(G107), .B1(KEYINPUT79), .B2(KEYINPUT3), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n388), .A2(G107), .ZN(new_n518));
  NAND4_X1  g332(.A1(new_n516), .A2(new_n517), .A3(new_n301), .A4(new_n518), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n512), .A2(new_n519), .ZN(new_n520));
  OAI21_X1  g334(.A(new_n500), .B1(new_n504), .B2(new_n520), .ZN(new_n521));
  NAND3_X1  g335(.A1(new_n516), .A2(new_n518), .A3(new_n517), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n522), .A2(G101), .ZN(new_n523));
  NAND3_X1  g337(.A1(new_n523), .A2(KEYINPUT4), .A3(new_n519), .ZN(new_n524));
  INV_X1    g338(.A(KEYINPUT4), .ZN(new_n525));
  NAND3_X1  g339(.A1(new_n522), .A2(new_n525), .A3(G101), .ZN(new_n526));
  NAND3_X1  g340(.A1(new_n524), .A2(new_n296), .A3(new_n526), .ZN(new_n527));
  AOI21_X1  g341(.A(new_n198), .B1(new_n361), .B2(KEYINPUT1), .ZN(new_n528));
  INV_X1    g342(.A(new_n357), .ZN(new_n529));
  OAI21_X1  g343(.A(new_n364), .B1(new_n528), .B2(new_n529), .ZN(new_n530));
  AND2_X1   g344(.A1(new_n512), .A2(new_n519), .ZN(new_n531));
  NAND3_X1  g345(.A1(new_n530), .A2(new_n531), .A3(KEYINPUT10), .ZN(new_n532));
  INV_X1    g346(.A(new_n289), .ZN(new_n533));
  NAND4_X1  g347(.A1(new_n521), .A2(new_n527), .A3(new_n532), .A4(new_n533), .ZN(new_n534));
  NAND3_X1  g348(.A1(new_n358), .A2(new_n520), .A3(new_n364), .ZN(new_n535));
  OAI21_X1  g349(.A(new_n535), .B1(new_n520), .B2(new_n504), .ZN(new_n536));
  AND3_X1   g350(.A1(new_n536), .A2(KEYINPUT12), .A3(new_n289), .ZN(new_n537));
  AOI21_X1  g351(.A(KEYINPUT12), .B1(new_n536), .B2(new_n289), .ZN(new_n538));
  OAI21_X1  g352(.A(new_n534), .B1(new_n537), .B2(new_n538), .ZN(new_n539));
  XNOR2_X1  g353(.A(G110), .B(G140), .ZN(new_n540));
  INV_X1    g354(.A(G227), .ZN(new_n541));
  NOR2_X1   g355(.A1(new_n541), .A2(G953), .ZN(new_n542));
  XOR2_X1   g356(.A(new_n540), .B(new_n542), .Z(new_n543));
  INV_X1    g357(.A(new_n543), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n539), .A2(new_n544), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n534), .A2(new_n543), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n546), .A2(KEYINPUT82), .ZN(new_n547));
  NAND3_X1  g361(.A1(new_n521), .A2(new_n527), .A3(new_n532), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n548), .A2(new_n289), .ZN(new_n549));
  INV_X1    g363(.A(KEYINPUT82), .ZN(new_n550));
  NAND3_X1  g364(.A1(new_n534), .A2(new_n550), .A3(new_n543), .ZN(new_n551));
  NAND3_X1  g365(.A1(new_n547), .A2(new_n549), .A3(new_n551), .ZN(new_n552));
  NAND3_X1  g366(.A1(new_n545), .A2(new_n552), .A3(G469), .ZN(new_n553));
  INV_X1    g367(.A(G469), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n536), .A2(new_n289), .ZN(new_n555));
  INV_X1    g369(.A(KEYINPUT12), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  NAND3_X1  g371(.A1(new_n536), .A2(KEYINPUT12), .A3(new_n289), .ZN(new_n558));
  AOI21_X1  g372(.A(new_n546), .B1(new_n557), .B2(new_n558), .ZN(new_n559));
  AOI21_X1  g373(.A(new_n543), .B1(new_n549), .B2(new_n534), .ZN(new_n560));
  OAI211_X1 g374(.A(new_n554), .B(new_n189), .C1(new_n559), .C2(new_n560), .ZN(new_n561));
  NAND2_X1  g375(.A1(G469), .A2(G902), .ZN(new_n562));
  NAND3_X1  g376(.A1(new_n553), .A2(new_n561), .A3(new_n562), .ZN(new_n563));
  INV_X1    g377(.A(KEYINPUT83), .ZN(new_n564));
  INV_X1    g378(.A(G221), .ZN(new_n565));
  AOI21_X1  g379(.A(new_n565), .B1(new_n476), .B2(new_n189), .ZN(new_n566));
  INV_X1    g380(.A(new_n566), .ZN(new_n567));
  AND3_X1   g381(.A1(new_n563), .A2(new_n564), .A3(new_n567), .ZN(new_n568));
  AOI21_X1  g382(.A(new_n564), .B1(new_n563), .B2(new_n567), .ZN(new_n569));
  OAI21_X1  g383(.A(new_n499), .B1(new_n568), .B2(new_n569), .ZN(new_n570));
  NAND2_X1  g384(.A1(G234), .A2(G237), .ZN(new_n571));
  NAND3_X1  g385(.A1(new_n571), .A2(G952), .A3(new_n233), .ZN(new_n572));
  XOR2_X1   g386(.A(KEYINPUT21), .B(G898), .Z(new_n573));
  NAND3_X1  g387(.A1(new_n571), .A2(G902), .A3(G953), .ZN(new_n574));
  OAI21_X1  g388(.A(new_n572), .B1(new_n573), .B2(new_n574), .ZN(new_n575));
  INV_X1    g389(.A(new_n575), .ZN(new_n576));
  XOR2_X1   g390(.A(G110), .B(G122), .Z(new_n577));
  INV_X1    g391(.A(new_n577), .ZN(new_n578));
  OAI211_X1 g392(.A(new_n524), .B(new_n526), .C1(new_n259), .C2(new_n260), .ZN(new_n579));
  OR3_X1    g393(.A1(new_n256), .A2(KEYINPUT85), .A3(KEYINPUT5), .ZN(new_n580));
  OAI21_X1  g394(.A(KEYINPUT85), .B1(new_n256), .B2(KEYINPUT5), .ZN(new_n581));
  NAND3_X1  g395(.A1(new_n256), .A2(KEYINPUT5), .A3(new_n257), .ZN(new_n582));
  NAND4_X1  g396(.A1(new_n580), .A2(new_n581), .A3(G113), .A4(new_n582), .ZN(new_n583));
  NAND3_X1  g397(.A1(new_n583), .A2(new_n258), .A3(new_n531), .ZN(new_n584));
  AOI211_X1 g398(.A(KEYINPUT86), .B(new_n578), .C1(new_n579), .C2(new_n584), .ZN(new_n585));
  NAND3_X1  g399(.A1(new_n579), .A2(new_n584), .A3(new_n578), .ZN(new_n586));
  INV_X1    g400(.A(new_n586), .ZN(new_n587));
  OAI21_X1  g401(.A(KEYINPUT6), .B1(new_n585), .B2(new_n587), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n579), .A2(new_n584), .ZN(new_n589));
  INV_X1    g403(.A(KEYINPUT86), .ZN(new_n590));
  NAND3_X1  g404(.A1(new_n589), .A2(new_n590), .A3(new_n577), .ZN(new_n591));
  INV_X1    g405(.A(KEYINPUT6), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n588), .A2(new_n593), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n530), .A2(new_n212), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n296), .A2(G125), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  INV_X1    g411(.A(G224), .ZN(new_n598));
  NOR2_X1   g412(.A1(new_n598), .A2(G953), .ZN(new_n599));
  XOR2_X1   g413(.A(new_n597), .B(new_n599), .Z(new_n600));
  AOI21_X1  g414(.A(G902), .B1(new_n594), .B2(new_n600), .ZN(new_n601));
  OAI21_X1  g415(.A(G210), .B1(G237), .B2(G902), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n583), .A2(new_n258), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n603), .A2(new_n520), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n604), .A2(new_n584), .ZN(new_n605));
  XOR2_X1   g419(.A(new_n577), .B(KEYINPUT8), .Z(new_n606));
  NAND2_X1  g420(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  INV_X1    g421(.A(KEYINPUT7), .ZN(new_n608));
  OAI211_X1 g422(.A(new_n595), .B(new_n596), .C1(new_n608), .C2(new_n599), .ZN(new_n609));
  OAI211_X1 g423(.A(new_n597), .B(KEYINPUT7), .C1(new_n598), .C2(G953), .ZN(new_n610));
  NAND4_X1  g424(.A1(new_n607), .A2(new_n609), .A3(new_n586), .A4(new_n610), .ZN(new_n611));
  NAND3_X1  g425(.A1(new_n601), .A2(new_n602), .A3(new_n611), .ZN(new_n612));
  AOI21_X1  g426(.A(new_n592), .B1(new_n591), .B2(new_n586), .ZN(new_n613));
  NOR2_X1   g427(.A1(new_n585), .A2(KEYINPUT6), .ZN(new_n614));
  OAI21_X1  g428(.A(new_n600), .B1(new_n613), .B2(new_n614), .ZN(new_n615));
  NAND3_X1  g429(.A1(new_n615), .A2(new_n189), .A3(new_n611), .ZN(new_n616));
  INV_X1    g430(.A(new_n602), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  AOI21_X1  g432(.A(new_n576), .B1(new_n612), .B2(new_n618), .ZN(new_n619));
  OAI21_X1  g433(.A(G214), .B1(G237), .B2(G902), .ZN(new_n620));
  XOR2_X1   g434(.A(new_n620), .B(KEYINPUT84), .Z(new_n621));
  NAND2_X1  g435(.A1(new_n619), .A2(new_n621), .ZN(new_n622));
  NOR2_X1   g436(.A1(new_n570), .A2(new_n622), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n385), .A2(new_n623), .ZN(new_n624));
  XNOR2_X1  g438(.A(new_n624), .B(G101), .ZN(G3));
  NAND2_X1  g439(.A1(new_n563), .A2(new_n567), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n626), .A2(KEYINPUT83), .ZN(new_n627));
  NAND3_X1  g441(.A1(new_n563), .A2(new_n564), .A3(new_n567), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n347), .A2(new_n189), .ZN(new_n630));
  AOI22_X1  g444(.A1(new_n630), .A2(G472), .B1(new_n348), .B2(new_n347), .ZN(new_n631));
  INV_X1    g445(.A(new_n247), .ZN(new_n632));
  AND3_X1   g446(.A1(new_n629), .A2(new_n631), .A3(new_n632), .ZN(new_n633));
  AOI21_X1  g447(.A(new_n602), .B1(new_n601), .B2(new_n611), .ZN(new_n634));
  AND4_X1   g448(.A1(new_n189), .A2(new_n615), .A3(new_n602), .A4(new_n611), .ZN(new_n635));
  OAI211_X1 g449(.A(new_n620), .B(new_n575), .C1(new_n634), .C2(new_n635), .ZN(new_n636));
  AOI21_X1  g450(.A(G478), .B1(new_n481), .B2(new_n189), .ZN(new_n637));
  NOR2_X1   g451(.A1(new_n483), .A2(new_n484), .ZN(new_n638));
  INV_X1    g452(.A(KEYINPUT96), .ZN(new_n639));
  OAI21_X1  g453(.A(KEYINPUT33), .B1(new_n484), .B2(new_n639), .ZN(new_n640));
  OR2_X1    g454(.A1(new_n638), .A2(new_n640), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n638), .A2(new_n640), .ZN(new_n642));
  AOI21_X1  g456(.A(G902), .B1(new_n641), .B2(new_n642), .ZN(new_n643));
  AOI21_X1  g457(.A(new_n637), .B1(new_n643), .B2(G478), .ZN(new_n644));
  INV_X1    g458(.A(new_n644), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n438), .A2(new_n645), .ZN(new_n646));
  NOR2_X1   g460(.A1(new_n636), .A2(new_n646), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n633), .A2(new_n647), .ZN(new_n648));
  XOR2_X1   g462(.A(KEYINPUT34), .B(G104), .Z(new_n649));
  XNOR2_X1  g463(.A(new_n648), .B(new_n649), .ZN(G6));
  AOI21_X1  g464(.A(new_n436), .B1(new_n492), .B2(new_n497), .ZN(new_n651));
  NAND3_X1  g465(.A1(new_n426), .A2(KEYINPUT97), .A3(new_n428), .ZN(new_n652));
  INV_X1    g466(.A(new_n652), .ZN(new_n653));
  AOI21_X1  g467(.A(KEYINPUT97), .B1(new_n426), .B2(new_n428), .ZN(new_n654));
  OAI21_X1  g468(.A(new_n651), .B1(new_n653), .B2(new_n654), .ZN(new_n655));
  NOR2_X1   g469(.A1(new_n636), .A2(new_n655), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n633), .A2(new_n656), .ZN(new_n657));
  XOR2_X1   g471(.A(KEYINPUT35), .B(G107), .Z(new_n658));
  XNOR2_X1  g472(.A(new_n657), .B(new_n658), .ZN(G9));
  NAND2_X1  g473(.A1(new_n630), .A2(G472), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n347), .A2(new_n348), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  XOR2_X1   g476(.A(new_n236), .B(KEYINPUT78), .Z(new_n663));
  INV_X1    g477(.A(KEYINPUT36), .ZN(new_n664));
  NAND2_X1  g478(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  OR2_X1    g479(.A1(new_n665), .A2(new_n232), .ZN(new_n666));
  NAND2_X1  g480(.A1(new_n665), .A2(new_n232), .ZN(new_n667));
  AND3_X1   g481(.A1(new_n666), .A2(new_n245), .A3(new_n667), .ZN(new_n668));
  INV_X1    g482(.A(new_n668), .ZN(new_n669));
  AOI21_X1  g483(.A(KEYINPUT98), .B1(new_n669), .B2(new_n244), .ZN(new_n670));
  INV_X1    g484(.A(KEYINPUT98), .ZN(new_n671));
  NOR3_X1   g485(.A1(new_n668), .A2(new_n243), .A3(new_n671), .ZN(new_n672));
  NOR2_X1   g486(.A1(new_n670), .A2(new_n672), .ZN(new_n673));
  NOR2_X1   g487(.A1(new_n662), .A2(new_n673), .ZN(new_n674));
  NAND2_X1  g488(.A1(new_n623), .A2(new_n674), .ZN(new_n675));
  XOR2_X1   g489(.A(new_n675), .B(KEYINPUT37), .Z(new_n676));
  XNOR2_X1  g490(.A(new_n676), .B(G110), .ZN(G12));
  AOI21_X1  g491(.A(new_n673), .B1(new_n351), .B2(new_n384), .ZN(new_n678));
  AOI21_X1  g492(.A(new_n489), .B1(new_n488), .B2(new_n491), .ZN(new_n679));
  NOR3_X1   g493(.A1(new_n495), .A2(new_n496), .A3(KEYINPUT95), .ZN(new_n680));
  OAI21_X1  g494(.A(new_n437), .B1(new_n679), .B2(new_n680), .ZN(new_n681));
  INV_X1    g495(.A(new_n654), .ZN(new_n682));
  AOI21_X1  g496(.A(new_n681), .B1(new_n682), .B2(new_n652), .ZN(new_n683));
  INV_X1    g497(.A(KEYINPUT100), .ZN(new_n684));
  INV_X1    g498(.A(new_n620), .ZN(new_n685));
  AOI21_X1  g499(.A(new_n685), .B1(new_n612), .B2(new_n618), .ZN(new_n686));
  INV_X1    g500(.A(new_n572), .ZN(new_n687));
  INV_X1    g501(.A(new_n574), .ZN(new_n688));
  XNOR2_X1  g502(.A(KEYINPUT99), .B(G900), .ZN(new_n689));
  AOI21_X1  g503(.A(new_n687), .B1(new_n688), .B2(new_n689), .ZN(new_n690));
  INV_X1    g504(.A(new_n690), .ZN(new_n691));
  NAND4_X1  g505(.A1(new_n683), .A2(new_n684), .A3(new_n686), .A4(new_n691), .ZN(new_n692));
  OAI211_X1 g506(.A(new_n651), .B(new_n691), .C1(new_n653), .C2(new_n654), .ZN(new_n693));
  OAI21_X1  g507(.A(new_n620), .B1(new_n634), .B2(new_n635), .ZN(new_n694));
  OAI21_X1  g508(.A(KEYINPUT100), .B1(new_n693), .B2(new_n694), .ZN(new_n695));
  NAND4_X1  g509(.A1(new_n678), .A2(new_n629), .A3(new_n692), .A4(new_n695), .ZN(new_n696));
  XNOR2_X1  g510(.A(new_n696), .B(G128), .ZN(G30));
  NAND2_X1  g511(.A1(new_n612), .A2(new_n618), .ZN(new_n698));
  INV_X1    g512(.A(KEYINPUT101), .ZN(new_n699));
  XNOR2_X1  g513(.A(new_n698), .B(new_n699), .ZN(new_n700));
  XNOR2_X1  g514(.A(new_n700), .B(KEYINPUT38), .ZN(new_n701));
  XNOR2_X1  g515(.A(new_n690), .B(KEYINPUT39), .ZN(new_n702));
  AOI21_X1  g516(.A(new_n702), .B1(new_n627), .B2(new_n628), .ZN(new_n703));
  INV_X1    g517(.A(KEYINPUT40), .ZN(new_n704));
  NAND2_X1  g518(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  INV_X1    g519(.A(new_n498), .ZN(new_n706));
  AOI21_X1  g520(.A(new_n436), .B1(new_n426), .B2(new_n428), .ZN(new_n707));
  NOR2_X1   g521(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  NAND3_X1  g522(.A1(new_n701), .A2(new_n705), .A3(new_n708), .ZN(new_n709));
  INV_X1    g523(.A(new_n709), .ZN(new_n710));
  AND2_X1   g524(.A1(new_n378), .A2(new_n380), .ZN(new_n711));
  OAI21_X1  g525(.A(new_n189), .B1(new_n711), .B2(new_n318), .ZN(new_n712));
  NAND2_X1  g526(.A1(new_n371), .A2(new_n318), .ZN(new_n713));
  INV_X1    g527(.A(new_n713), .ZN(new_n714));
  OAI21_X1  g528(.A(G472), .B1(new_n712), .B2(new_n714), .ZN(new_n715));
  NAND2_X1  g529(.A1(new_n351), .A2(new_n715), .ZN(new_n716));
  XOR2_X1   g530(.A(new_n716), .B(KEYINPUT102), .Z(new_n717));
  NAND2_X1  g531(.A1(new_n669), .A2(new_n244), .ZN(new_n718));
  NOR2_X1   g532(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  OR2_X1    g533(.A1(new_n703), .A2(new_n704), .ZN(new_n720));
  NAND4_X1  g534(.A1(new_n710), .A2(new_n719), .A3(new_n620), .A4(new_n720), .ZN(new_n721));
  XNOR2_X1  g535(.A(new_n721), .B(G143), .ZN(G45));
  NOR2_X1   g536(.A1(new_n646), .A2(new_n690), .ZN(new_n723));
  NAND4_X1  g537(.A1(new_n678), .A2(new_n629), .A3(new_n686), .A4(new_n723), .ZN(new_n724));
  XNOR2_X1  g538(.A(new_n724), .B(G146), .ZN(G48));
  INV_X1    g539(.A(KEYINPUT32), .ZN(new_n726));
  NAND2_X1  g540(.A1(new_n661), .A2(new_n726), .ZN(new_n727));
  NAND3_X1  g541(.A1(new_n347), .A2(KEYINPUT32), .A3(new_n348), .ZN(new_n728));
  NAND3_X1  g542(.A1(new_n384), .A2(new_n727), .A3(new_n728), .ZN(new_n729));
  OAI21_X1  g543(.A(new_n189), .B1(new_n559), .B2(new_n560), .ZN(new_n730));
  NAND2_X1  g544(.A1(new_n730), .A2(G469), .ZN(new_n731));
  NAND2_X1  g545(.A1(new_n731), .A2(new_n561), .ZN(new_n732));
  NOR2_X1   g546(.A1(new_n732), .A2(new_n566), .ZN(new_n733));
  NAND4_X1  g547(.A1(new_n729), .A2(new_n647), .A3(new_n632), .A4(new_n733), .ZN(new_n734));
  XNOR2_X1  g548(.A(KEYINPUT41), .B(G113), .ZN(new_n735));
  XNOR2_X1  g549(.A(new_n734), .B(new_n735), .ZN(G15));
  NAND4_X1  g550(.A1(new_n729), .A2(new_n656), .A3(new_n632), .A4(new_n733), .ZN(new_n737));
  XNOR2_X1  g551(.A(new_n737), .B(G116), .ZN(G18));
  OR2_X1    g552(.A1(new_n670), .A2(new_n672), .ZN(new_n739));
  AND2_X1   g553(.A1(new_n383), .A2(G472), .ZN(new_n740));
  NAND2_X1  g554(.A1(new_n727), .A2(new_n728), .ZN(new_n741));
  OAI211_X1 g555(.A(new_n499), .B(new_n739), .C1(new_n740), .C2(new_n741), .ZN(new_n742));
  NAND2_X1  g556(.A1(new_n686), .A2(new_n733), .ZN(new_n743));
  INV_X1    g557(.A(new_n743), .ZN(new_n744));
  NAND2_X1  g558(.A1(new_n744), .A2(new_n575), .ZN(new_n745));
  OAI21_X1  g559(.A(KEYINPUT103), .B1(new_n742), .B2(new_n745), .ZN(new_n746));
  NOR2_X1   g560(.A1(new_n743), .A2(new_n576), .ZN(new_n747));
  INV_X1    g561(.A(KEYINPUT103), .ZN(new_n748));
  NAND4_X1  g562(.A1(new_n678), .A2(new_n747), .A3(new_n748), .A4(new_n499), .ZN(new_n749));
  NAND2_X1  g563(.A1(new_n746), .A2(new_n749), .ZN(new_n750));
  XNOR2_X1  g564(.A(new_n750), .B(G119), .ZN(G21));
  INV_X1    g565(.A(G472), .ZN(new_n752));
  AOI21_X1  g566(.A(new_n752), .B1(new_n347), .B2(new_n189), .ZN(new_n753));
  NAND2_X1  g567(.A1(new_n381), .A2(new_n374), .ZN(new_n754));
  NAND2_X1  g568(.A1(new_n754), .A2(new_n317), .ZN(new_n755));
  NAND3_X1  g569(.A1(new_n755), .A2(KEYINPUT104), .A3(new_n325), .ZN(new_n756));
  INV_X1    g570(.A(KEYINPUT104), .ZN(new_n757));
  AOI21_X1  g571(.A(new_n318), .B1(new_n381), .B2(new_n374), .ZN(new_n758));
  AOI21_X1  g572(.A(new_n332), .B1(new_n368), .B2(new_n318), .ZN(new_n759));
  OAI21_X1  g573(.A(new_n757), .B1(new_n758), .B2(new_n759), .ZN(new_n760));
  NAND3_X1  g574(.A1(new_n756), .A2(new_n333), .A3(new_n760), .ZN(new_n761));
  AOI21_X1  g575(.A(new_n753), .B1(new_n761), .B2(new_n348), .ZN(new_n762));
  AND2_X1   g576(.A1(new_n762), .A2(new_n632), .ZN(new_n763));
  OAI21_X1  g577(.A(KEYINPUT105), .B1(new_n706), .B2(new_n707), .ZN(new_n764));
  INV_X1    g578(.A(KEYINPUT105), .ZN(new_n765));
  NAND3_X1  g579(.A1(new_n438), .A2(new_n765), .A3(new_n498), .ZN(new_n766));
  AND3_X1   g580(.A1(new_n764), .A2(new_n686), .A3(new_n766), .ZN(new_n767));
  NAND4_X1  g581(.A1(new_n763), .A2(new_n575), .A3(new_n733), .A4(new_n767), .ZN(new_n768));
  XNOR2_X1  g582(.A(new_n768), .B(G122), .ZN(G24));
  NAND4_X1  g583(.A1(new_n744), .A2(new_n762), .A3(new_n718), .A4(new_n723), .ZN(new_n770));
  XNOR2_X1  g584(.A(new_n770), .B(G125), .ZN(G27));
  INV_X1    g585(.A(KEYINPUT42), .ZN(new_n772));
  NAND3_X1  g586(.A1(new_n612), .A2(new_n618), .A3(new_n620), .ZN(new_n773));
  NOR2_X1   g587(.A1(new_n773), .A2(new_n626), .ZN(new_n774));
  OAI211_X1 g588(.A(new_n632), .B(new_n774), .C1(new_n740), .C2(new_n741), .ZN(new_n775));
  INV_X1    g589(.A(new_n723), .ZN(new_n776));
  OAI21_X1  g590(.A(new_n772), .B1(new_n775), .B2(new_n776), .ZN(new_n777));
  NAND4_X1  g591(.A1(new_n385), .A2(KEYINPUT42), .A3(new_n723), .A4(new_n774), .ZN(new_n778));
  NAND2_X1  g592(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  XNOR2_X1  g593(.A(new_n779), .B(G131), .ZN(G33));
  INV_X1    g594(.A(new_n693), .ZN(new_n781));
  NAND4_X1  g595(.A1(new_n729), .A2(new_n632), .A3(new_n781), .A4(new_n774), .ZN(new_n782));
  XNOR2_X1  g596(.A(new_n782), .B(G134), .ZN(G36));
  INV_X1    g597(.A(KEYINPUT107), .ZN(new_n784));
  AOI21_X1  g598(.A(KEYINPUT43), .B1(new_n707), .B2(new_n784), .ZN(new_n785));
  NAND2_X1  g599(.A1(new_n707), .A2(new_n645), .ZN(new_n786));
  XNOR2_X1  g600(.A(new_n785), .B(new_n786), .ZN(new_n787));
  NAND3_X1  g601(.A1(new_n787), .A2(new_n662), .A3(new_n718), .ZN(new_n788));
  XNOR2_X1  g602(.A(new_n788), .B(KEYINPUT44), .ZN(new_n789));
  INV_X1    g603(.A(new_n773), .ZN(new_n790));
  NAND2_X1  g604(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  XNOR2_X1  g605(.A(new_n791), .B(KEYINPUT108), .ZN(new_n792));
  NAND2_X1  g606(.A1(new_n545), .A2(new_n552), .ZN(new_n793));
  XNOR2_X1  g607(.A(new_n793), .B(KEYINPUT45), .ZN(new_n794));
  NAND2_X1  g608(.A1(new_n794), .A2(G469), .ZN(new_n795));
  NAND3_X1  g609(.A1(new_n795), .A2(KEYINPUT46), .A3(new_n562), .ZN(new_n796));
  INV_X1    g610(.A(KEYINPUT46), .ZN(new_n797));
  OAI211_X1 g611(.A(new_n797), .B(G469), .C1(new_n794), .C2(G902), .ZN(new_n798));
  NAND3_X1  g612(.A1(new_n796), .A2(new_n561), .A3(new_n798), .ZN(new_n799));
  NAND2_X1  g613(.A1(new_n799), .A2(new_n567), .ZN(new_n800));
  OR2_X1    g614(.A1(new_n800), .A2(new_n702), .ZN(new_n801));
  XOR2_X1   g615(.A(new_n801), .B(KEYINPUT106), .Z(new_n802));
  NAND2_X1  g616(.A1(new_n792), .A2(new_n802), .ZN(new_n803));
  XNOR2_X1  g617(.A(new_n803), .B(G137), .ZN(G39));
  AND2_X1   g618(.A1(new_n800), .A2(KEYINPUT109), .ZN(new_n805));
  NOR2_X1   g619(.A1(new_n800), .A2(KEYINPUT109), .ZN(new_n806));
  INV_X1    g620(.A(KEYINPUT47), .ZN(new_n807));
  OR3_X1    g621(.A1(new_n805), .A2(new_n806), .A3(new_n807), .ZN(new_n808));
  OAI21_X1  g622(.A(new_n807), .B1(new_n805), .B2(new_n806), .ZN(new_n809));
  AOI21_X1  g623(.A(new_n729), .B1(new_n808), .B2(new_n809), .ZN(new_n810));
  NAND4_X1  g624(.A1(new_n810), .A2(new_n247), .A3(new_n723), .A4(new_n790), .ZN(new_n811));
  XNOR2_X1  g625(.A(new_n811), .B(G140), .ZN(G42));
  INV_X1    g626(.A(new_n701), .ZN(new_n813));
  AND2_X1   g627(.A1(new_n763), .A2(new_n733), .ZN(new_n814));
  AND2_X1   g628(.A1(new_n787), .A2(new_n687), .ZN(new_n815));
  NAND4_X1  g629(.A1(new_n813), .A2(new_n685), .A3(new_n814), .A4(new_n815), .ZN(new_n816));
  XOR2_X1   g630(.A(new_n816), .B(KEYINPUT50), .Z(new_n817));
  NOR3_X1   g631(.A1(new_n773), .A2(new_n566), .A3(new_n732), .ZN(new_n818));
  AND4_X1   g632(.A1(new_n632), .A2(new_n717), .A3(new_n687), .A4(new_n818), .ZN(new_n819));
  NAND3_X1  g633(.A1(new_n819), .A2(new_n707), .A3(new_n644), .ZN(new_n820));
  NAND2_X1  g634(.A1(new_n815), .A2(new_n818), .ZN(new_n821));
  XNOR2_X1  g635(.A(new_n821), .B(KEYINPUT116), .ZN(new_n822));
  AND2_X1   g636(.A1(new_n762), .A2(new_n718), .ZN(new_n823));
  NAND2_X1  g637(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  AND2_X1   g638(.A1(new_n824), .A2(KEYINPUT117), .ZN(new_n825));
  NOR2_X1   g639(.A1(new_n824), .A2(KEYINPUT117), .ZN(new_n826));
  OAI211_X1 g640(.A(new_n817), .B(new_n820), .C1(new_n825), .C2(new_n826), .ZN(new_n827));
  INV_X1    g641(.A(new_n827), .ZN(new_n828));
  XNOR2_X1  g642(.A(new_n732), .B(KEYINPUT110), .ZN(new_n829));
  NAND2_X1  g643(.A1(new_n829), .A2(new_n566), .ZN(new_n830));
  NAND3_X1  g644(.A1(new_n808), .A2(new_n809), .A3(new_n830), .ZN(new_n831));
  AND3_X1   g645(.A1(new_n815), .A2(new_n763), .A3(new_n790), .ZN(new_n832));
  NAND2_X1  g646(.A1(new_n831), .A2(new_n832), .ZN(new_n833));
  NAND3_X1  g647(.A1(new_n828), .A2(KEYINPUT51), .A3(new_n833), .ZN(new_n834));
  NAND2_X1  g648(.A1(new_n233), .A2(G952), .ZN(new_n835));
  AOI21_X1  g649(.A(new_n644), .B1(new_n429), .B2(new_n437), .ZN(new_n836));
  AOI21_X1  g650(.A(new_n835), .B1(new_n819), .B2(new_n836), .ZN(new_n837));
  AND2_X1   g651(.A1(new_n822), .A2(new_n385), .ZN(new_n838));
  OAI21_X1  g652(.A(new_n837), .B1(new_n838), .B2(KEYINPUT48), .ZN(new_n839));
  AOI21_X1  g653(.A(new_n839), .B1(KEYINPUT48), .B2(new_n838), .ZN(new_n840));
  AND2_X1   g654(.A1(new_n834), .A2(new_n840), .ZN(new_n841));
  NAND3_X1  g655(.A1(new_n814), .A2(new_n686), .A3(new_n815), .ZN(new_n842));
  AND3_X1   g656(.A1(new_n729), .A2(new_n629), .A3(new_n739), .ZN(new_n843));
  NAND2_X1  g657(.A1(new_n488), .A2(new_n491), .ZN(new_n844));
  NOR2_X1   g658(.A1(new_n844), .A2(new_n690), .ZN(new_n845));
  OAI211_X1 g659(.A(new_n437), .B(new_n845), .C1(new_n653), .C2(new_n654), .ZN(new_n846));
  INV_X1    g660(.A(KEYINPUT112), .ZN(new_n847));
  OR2_X1    g661(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  NAND2_X1  g662(.A1(new_n846), .A2(new_n847), .ZN(new_n849));
  NAND4_X1  g663(.A1(new_n843), .A2(new_n848), .A3(new_n790), .A4(new_n849), .ZN(new_n850));
  NAND4_X1  g664(.A1(new_n762), .A2(new_n718), .A3(new_n723), .A4(new_n774), .ZN(new_n851));
  NAND2_X1  g665(.A1(new_n782), .A2(new_n851), .ZN(new_n852));
  INV_X1    g666(.A(new_n852), .ZN(new_n853));
  NAND3_X1  g667(.A1(new_n779), .A2(new_n850), .A3(new_n853), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n734), .A2(new_n737), .ZN(new_n855));
  INV_X1    g669(.A(new_n855), .ZN(new_n856));
  NAND2_X1  g670(.A1(new_n750), .A2(new_n856), .ZN(new_n857));
  NAND4_X1  g671(.A1(new_n698), .A2(new_n836), .A3(new_n621), .A4(new_n575), .ZN(new_n858));
  INV_X1    g672(.A(KEYINPUT111), .ZN(new_n859));
  NAND2_X1  g673(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  NAND4_X1  g674(.A1(new_n619), .A2(KEYINPUT111), .A3(new_n621), .A4(new_n836), .ZN(new_n861));
  NAND2_X1  g675(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  AOI22_X1  g676(.A1(new_n862), .A2(new_n633), .B1(new_n385), .B2(new_n623), .ZN(new_n863));
  NAND2_X1  g677(.A1(new_n707), .A2(new_n844), .ZN(new_n864));
  NOR2_X1   g678(.A1(new_n622), .A2(new_n864), .ZN(new_n865));
  AOI22_X1  g679(.A1(new_n633), .A2(new_n865), .B1(new_n623), .B2(new_n674), .ZN(new_n866));
  NAND3_X1  g680(.A1(new_n863), .A2(new_n768), .A3(new_n866), .ZN(new_n867));
  NOR3_X1   g681(.A1(new_n854), .A2(new_n857), .A3(new_n867), .ZN(new_n868));
  INV_X1    g682(.A(new_n626), .ZN(new_n869));
  NOR2_X1   g683(.A1(new_n718), .A2(new_n690), .ZN(new_n870));
  NAND4_X1  g684(.A1(new_n716), .A2(new_n767), .A3(new_n869), .A4(new_n870), .ZN(new_n871));
  NAND4_X1  g685(.A1(new_n696), .A2(new_n724), .A3(new_n770), .A4(new_n871), .ZN(new_n872));
  INV_X1    g686(.A(KEYINPUT52), .ZN(new_n873));
  XNOR2_X1  g687(.A(new_n872), .B(new_n873), .ZN(new_n874));
  XOR2_X1   g688(.A(KEYINPUT114), .B(KEYINPUT53), .Z(new_n875));
  NAND3_X1  g689(.A1(new_n868), .A2(new_n874), .A3(new_n875), .ZN(new_n876));
  INV_X1    g690(.A(KEYINPUT114), .ZN(new_n877));
  NAND2_X1  g691(.A1(new_n877), .A2(KEYINPUT53), .ZN(new_n878));
  AND3_X1   g692(.A1(new_n863), .A2(new_n768), .A3(new_n866), .ZN(new_n879));
  AOI21_X1  g693(.A(new_n855), .B1(new_n749), .B2(new_n746), .ZN(new_n880));
  AOI21_X1  g694(.A(new_n852), .B1(new_n777), .B2(new_n778), .ZN(new_n881));
  NAND4_X1  g695(.A1(new_n879), .A2(new_n880), .A3(new_n850), .A4(new_n881), .ZN(new_n882));
  AND2_X1   g696(.A1(new_n692), .A2(new_n695), .ZN(new_n883));
  NAND2_X1  g697(.A1(new_n761), .A2(new_n348), .ZN(new_n884));
  AND4_X1   g698(.A1(new_n660), .A2(new_n884), .A3(new_n718), .A4(new_n723), .ZN(new_n885));
  AOI22_X1  g699(.A1(new_n843), .A2(new_n883), .B1(new_n885), .B2(new_n744), .ZN(new_n886));
  NAND4_X1  g700(.A1(new_n886), .A2(new_n873), .A3(new_n724), .A4(new_n871), .ZN(new_n887));
  NAND2_X1  g701(.A1(new_n872), .A2(KEYINPUT52), .ZN(new_n888));
  NAND2_X1  g702(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  OAI21_X1  g703(.A(new_n878), .B1(new_n882), .B2(new_n889), .ZN(new_n890));
  NAND2_X1  g704(.A1(new_n876), .A2(new_n890), .ZN(new_n891));
  NOR2_X1   g705(.A1(new_n891), .A2(KEYINPUT54), .ZN(new_n892));
  AOI21_X1  g706(.A(KEYINPUT53), .B1(new_n874), .B2(KEYINPUT113), .ZN(new_n893));
  NAND2_X1  g707(.A1(new_n868), .A2(new_n874), .ZN(new_n894));
  XNOR2_X1  g708(.A(new_n893), .B(new_n894), .ZN(new_n895));
  AOI21_X1  g709(.A(new_n892), .B1(new_n895), .B2(KEYINPUT54), .ZN(new_n896));
  INV_X1    g710(.A(KEYINPUT51), .ZN(new_n897));
  XNOR2_X1  g711(.A(new_n830), .B(KEYINPUT115), .ZN(new_n898));
  NAND3_X1  g712(.A1(new_n808), .A2(new_n809), .A3(new_n898), .ZN(new_n899));
  AND2_X1   g713(.A1(new_n899), .A2(new_n832), .ZN(new_n900));
  OAI21_X1  g714(.A(new_n897), .B1(new_n827), .B2(new_n900), .ZN(new_n901));
  NAND4_X1  g715(.A1(new_n841), .A2(new_n842), .A3(new_n896), .A4(new_n901), .ZN(new_n902));
  OAI21_X1  g716(.A(new_n902), .B1(G952), .B2(G953), .ZN(new_n903));
  XNOR2_X1  g717(.A(new_n829), .B(KEYINPUT49), .ZN(new_n904));
  AND4_X1   g718(.A1(new_n632), .A2(new_n904), .A3(new_n621), .A4(new_n567), .ZN(new_n905));
  INV_X1    g719(.A(new_n786), .ZN(new_n906));
  NAND3_X1  g720(.A1(new_n905), .A2(new_n717), .A3(new_n906), .ZN(new_n907));
  OAI21_X1  g721(.A(new_n903), .B1(new_n701), .B2(new_n907), .ZN(G75));
  INV_X1    g722(.A(new_n891), .ZN(new_n909));
  NOR2_X1   g723(.A1(new_n909), .A2(new_n189), .ZN(new_n910));
  NAND2_X1  g724(.A1(new_n910), .A2(G210), .ZN(new_n911));
  XOR2_X1   g725(.A(new_n594), .B(new_n600), .Z(new_n912));
  XNOR2_X1  g726(.A(new_n912), .B(KEYINPUT55), .ZN(new_n913));
  XOR2_X1   g727(.A(KEYINPUT118), .B(KEYINPUT56), .Z(new_n914));
  AND3_X1   g728(.A1(new_n911), .A2(new_n913), .A3(new_n914), .ZN(new_n915));
  INV_X1    g729(.A(KEYINPUT56), .ZN(new_n916));
  AOI21_X1  g730(.A(new_n913), .B1(new_n911), .B2(new_n916), .ZN(new_n917));
  NOR2_X1   g731(.A1(new_n233), .A2(G952), .ZN(new_n918));
  NOR3_X1   g732(.A1(new_n915), .A2(new_n917), .A3(new_n918), .ZN(G51));
  AND2_X1   g733(.A1(new_n891), .A2(KEYINPUT54), .ZN(new_n920));
  OR2_X1    g734(.A1(new_n920), .A2(new_n892), .ZN(new_n921));
  XOR2_X1   g735(.A(new_n562), .B(KEYINPUT57), .Z(new_n922));
  NAND2_X1  g736(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  INV_X1    g737(.A(KEYINPUT119), .ZN(new_n924));
  NAND2_X1  g738(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  NAND3_X1  g739(.A1(new_n921), .A2(KEYINPUT119), .A3(new_n922), .ZN(new_n926));
  OAI211_X1 g740(.A(new_n925), .B(new_n926), .C1(new_n560), .C2(new_n559), .ZN(new_n927));
  NAND3_X1  g741(.A1(new_n910), .A2(G469), .A3(new_n794), .ZN(new_n928));
  AOI21_X1  g742(.A(new_n918), .B1(new_n927), .B2(new_n928), .ZN(G54));
  NAND3_X1  g743(.A1(new_n910), .A2(KEYINPUT58), .A3(G475), .ZN(new_n930));
  NOR2_X1   g744(.A1(new_n415), .A2(new_n424), .ZN(new_n931));
  XNOR2_X1  g745(.A(new_n930), .B(new_n931), .ZN(new_n932));
  NOR2_X1   g746(.A1(new_n932), .A2(new_n918), .ZN(G60));
  NOR2_X1   g747(.A1(new_n920), .A2(new_n892), .ZN(new_n934));
  NAND2_X1  g748(.A1(G478), .A2(G902), .ZN(new_n935));
  XOR2_X1   g749(.A(new_n935), .B(KEYINPUT59), .Z(new_n936));
  NAND2_X1  g750(.A1(new_n641), .A2(new_n642), .ZN(new_n937));
  XOR2_X1   g751(.A(new_n937), .B(KEYINPUT120), .Z(new_n938));
  NOR3_X1   g752(.A1(new_n934), .A2(new_n936), .A3(new_n938), .ZN(new_n939));
  OR2_X1    g753(.A1(new_n896), .A2(new_n936), .ZN(new_n940));
  AOI211_X1 g754(.A(new_n918), .B(new_n939), .C1(new_n938), .C2(new_n940), .ZN(G63));
  INV_X1    g755(.A(KEYINPUT122), .ZN(new_n942));
  NAND2_X1  g756(.A1(G217), .A2(G902), .ZN(new_n943));
  XOR2_X1   g757(.A(new_n943), .B(KEYINPUT121), .Z(new_n944));
  XOR2_X1   g758(.A(new_n944), .B(KEYINPUT60), .Z(new_n945));
  AOI21_X1  g759(.A(new_n942), .B1(new_n891), .B2(new_n945), .ZN(new_n946));
  INV_X1    g760(.A(new_n945), .ZN(new_n947));
  AOI211_X1 g761(.A(KEYINPUT122), .B(new_n947), .C1(new_n876), .C2(new_n890), .ZN(new_n948));
  NOR2_X1   g762(.A1(new_n946), .A2(new_n948), .ZN(new_n949));
  AOI21_X1  g763(.A(new_n918), .B1(new_n949), .B2(new_n240), .ZN(new_n950));
  AND2_X1   g764(.A1(new_n666), .A2(new_n667), .ZN(new_n951));
  OAI21_X1  g765(.A(new_n951), .B1(new_n946), .B2(new_n948), .ZN(new_n952));
  NAND3_X1  g766(.A1(new_n950), .A2(KEYINPUT61), .A3(new_n952), .ZN(new_n953));
  INV_X1    g767(.A(KEYINPUT123), .ZN(new_n954));
  NAND2_X1  g768(.A1(new_n952), .A2(new_n954), .ZN(new_n955));
  OAI211_X1 g769(.A(KEYINPUT123), .B(new_n951), .C1(new_n946), .C2(new_n948), .ZN(new_n956));
  NAND3_X1  g770(.A1(new_n950), .A2(new_n955), .A3(new_n956), .ZN(new_n957));
  INV_X1    g771(.A(KEYINPUT124), .ZN(new_n958));
  INV_X1    g772(.A(KEYINPUT61), .ZN(new_n959));
  AND3_X1   g773(.A1(new_n957), .A2(new_n958), .A3(new_n959), .ZN(new_n960));
  AOI21_X1  g774(.A(new_n958), .B1(new_n957), .B2(new_n959), .ZN(new_n961));
  OAI21_X1  g775(.A(new_n953), .B1(new_n960), .B2(new_n961), .ZN(G66));
  NOR2_X1   g776(.A1(new_n857), .A2(new_n867), .ZN(new_n963));
  NOR2_X1   g777(.A1(new_n963), .A2(G953), .ZN(new_n964));
  AOI21_X1  g778(.A(new_n233), .B1(new_n573), .B2(G224), .ZN(new_n965));
  OAI21_X1  g779(.A(KEYINPUT125), .B1(new_n964), .B2(new_n965), .ZN(new_n966));
  OAI21_X1  g780(.A(new_n966), .B1(KEYINPUT125), .B2(new_n965), .ZN(new_n967));
  OAI211_X1 g781(.A(new_n588), .B(new_n593), .C1(G898), .C2(new_n233), .ZN(new_n968));
  XNOR2_X1  g782(.A(new_n967), .B(new_n968), .ZN(G69));
  AND2_X1   g783(.A1(new_n886), .A2(new_n724), .ZN(new_n970));
  AND2_X1   g784(.A1(new_n811), .A2(new_n970), .ZN(new_n971));
  AND2_X1   g785(.A1(new_n385), .A2(new_n767), .ZN(new_n972));
  OAI21_X1  g786(.A(new_n802), .B1(new_n792), .B2(new_n972), .ZN(new_n973));
  AND2_X1   g787(.A1(new_n779), .A2(new_n782), .ZN(new_n974));
  NAND4_X1  g788(.A1(new_n971), .A2(new_n233), .A3(new_n973), .A4(new_n974), .ZN(new_n975));
  INV_X1    g789(.A(G900), .ZN(new_n976));
  NOR2_X1   g790(.A1(new_n976), .A2(new_n233), .ZN(new_n977));
  INV_X1    g791(.A(new_n977), .ZN(new_n978));
  NAND2_X1  g792(.A1(new_n975), .A2(new_n978), .ZN(new_n979));
  NAND2_X1  g793(.A1(new_n721), .A2(new_n970), .ZN(new_n980));
  INV_X1    g794(.A(KEYINPUT62), .ZN(new_n981));
  XNOR2_X1  g795(.A(new_n980), .B(new_n981), .ZN(new_n982));
  AND2_X1   g796(.A1(new_n982), .A2(new_n811), .ZN(new_n983));
  NAND2_X1  g797(.A1(new_n646), .A2(new_n864), .ZN(new_n984));
  NAND4_X1  g798(.A1(new_n385), .A2(new_n703), .A3(new_n790), .A4(new_n984), .ZN(new_n985));
  AND2_X1   g799(.A1(new_n803), .A2(new_n985), .ZN(new_n986));
  AOI21_X1  g800(.A(G953), .B1(new_n983), .B2(new_n986), .ZN(new_n987));
  XNOR2_X1  g801(.A(new_n323), .B(new_n406), .ZN(new_n988));
  NOR2_X1   g802(.A1(new_n988), .A2(KEYINPUT126), .ZN(new_n989));
  OAI21_X1  g803(.A(new_n979), .B1(new_n987), .B2(new_n989), .ZN(new_n990));
  OAI21_X1  g804(.A(new_n988), .B1(new_n987), .B2(KEYINPUT126), .ZN(new_n991));
  NAND2_X1  g805(.A1(new_n990), .A2(new_n991), .ZN(new_n992));
  OAI21_X1  g806(.A(G953), .B1(new_n541), .B2(new_n976), .ZN(new_n993));
  XOR2_X1   g807(.A(new_n993), .B(KEYINPUT127), .Z(new_n994));
  INV_X1    g808(.A(new_n994), .ZN(new_n995));
  NAND2_X1  g809(.A1(new_n992), .A2(new_n995), .ZN(new_n996));
  NAND3_X1  g810(.A1(new_n991), .A2(new_n990), .A3(new_n994), .ZN(new_n997));
  NAND2_X1  g811(.A1(new_n996), .A2(new_n997), .ZN(G72));
  NAND3_X1  g812(.A1(new_n983), .A2(new_n963), .A3(new_n986), .ZN(new_n999));
  NAND2_X1  g813(.A1(G472), .A2(G902), .ZN(new_n1000));
  XOR2_X1   g814(.A(new_n1000), .B(KEYINPUT63), .Z(new_n1001));
  NAND2_X1  g815(.A1(new_n999), .A2(new_n1001), .ZN(new_n1002));
  AOI21_X1  g816(.A(new_n918), .B1(new_n1002), .B2(new_n714), .ZN(new_n1003));
  AND4_X1   g817(.A1(new_n963), .A2(new_n971), .A3(new_n973), .A4(new_n974), .ZN(new_n1004));
  INV_X1    g818(.A(new_n1001), .ZN(new_n1005));
  OAI211_X1 g819(.A(new_n317), .B(new_n368), .C1(new_n1004), .C2(new_n1005), .ZN(new_n1006));
  NAND3_X1  g820(.A1(new_n369), .A2(new_n324), .A3(new_n372), .ZN(new_n1007));
  NAND3_X1  g821(.A1(new_n895), .A2(new_n1001), .A3(new_n1007), .ZN(new_n1008));
  AND3_X1   g822(.A1(new_n1003), .A2(new_n1006), .A3(new_n1008), .ZN(G57));
endmodule


