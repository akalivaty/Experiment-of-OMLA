

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n513, n514, n515, n516,
         n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527,
         n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538,
         n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549,
         n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560,
         n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571,
         n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582,
         n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593,
         n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604,
         n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615,
         n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626,
         n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637,
         n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648,
         n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659,
         n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670,
         n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681,
         n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692,
         n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703,
         n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714,
         n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725,
         n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736,
         n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747,
         n748, n749, n750, n751, n752, n753, n754, n755, n756, n757, n758,
         n759, n760, n761, n762, n763, n764, n765, n766, n767, n768, n769,
         n770, n771, n772, n773, n774, n775, n776, n777, n778, n779, n780,
         n781, n782, n783, n784, n785, n786, n787, n788, n789, n790, n791,
         n792, n793, n794, n795, n796, n797, n798, n799, n800, n801, n802,
         n803, n804, n805, n806, n807, n808, n809, n810, n811, n812, n813,
         n814, n815, n816, n817, n818, n819, n820, n821, n822, n823, n824,
         n825, n826, n827, n828, n829, n830, n831, n832, n833, n834, n835,
         n836, n837, n838, n839, n840, n841, n842, n843, n844, n845, n846,
         n847, n848, n849, n850, n851, n852, n853, n854, n855, n856, n857,
         n858, n859, n860, n861, n862, n863, n864, n865, n866, n867, n868,
         n869, n870, n871, n872, n873, n874, n875, n876, n877, n878, n879,
         n880, n881, n882, n883, n884, n885, n886, n887, n888, n889, n890,
         n891, n892, n893, n894, n895, n896, n897, n898, n899, n900, n901,
         n902, n903, n904, n905, n906, n907, n908, n909, n910, n911, n912,
         n913, n914, n915, n916, n917, n918, n919, n920, n921, n922, n923,
         n924, n925, n926, n927, n928, n929, n930, n931, n932, n933, n934,
         n935, n936, n937, n938, n939, n940, n941, n942, n943, n944, n945,
         n946, n947, n948, n949, n950, n951, n952, n953, n954, n955, n956,
         n957, n958, n959, n960, n961, n962, n963, n964, n965, n966, n967,
         n968, n969, n970, n971, n972, n973, n974, n975, n976, n977, n978,
         n979, n980, n981, n982, n983, n984, n985, n986, n987, n988, n989,
         n990, n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000,
         n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  XNOR2_X1 U550 ( .A(n524), .B(KEYINPUT66), .ZN(n882) );
  XOR2_X1 U551 ( .A(KEYINPUT76), .B(n597), .Z(n513) );
  OR2_X1 U552 ( .A1(n694), .A2(n683), .ZN(n514) );
  NAND2_X1 U553 ( .A1(n698), .A2(n697), .ZN(n515) );
  OR2_X1 U554 ( .A1(n686), .A2(n685), .ZN(n516) );
  NOR2_X1 U555 ( .A1(n912), .A2(n618), .ZN(n620) );
  NAND2_X1 U556 ( .A1(n673), .A2(n672), .ZN(n689) );
  NAND2_X1 U557 ( .A1(n680), .A2(n614), .ZN(n656) );
  NAND2_X1 U558 ( .A1(n684), .A2(n514), .ZN(n685) );
  NOR2_X2 U559 ( .A1(G2105), .A2(n522), .ZN(n881) );
  XOR2_X1 U560 ( .A(KEYINPUT77), .B(n602), .Z(n906) );
  NOR2_X1 U561 ( .A1(G651), .A2(n571), .ZN(n788) );
  XOR2_X1 U562 ( .A(KEYINPUT23), .B(KEYINPUT64), .Z(n518) );
  INV_X1 U563 ( .A(G2104), .ZN(n522) );
  NAND2_X1 U564 ( .A1(G101), .A2(n881), .ZN(n517) );
  XNOR2_X1 U565 ( .A(n518), .B(n517), .ZN(n521) );
  AND2_X1 U566 ( .A1(G2104), .A2(G2105), .ZN(n877) );
  NAND2_X1 U567 ( .A1(G113), .A2(n877), .ZN(n519) );
  XOR2_X1 U568 ( .A(KEYINPUT65), .B(n519), .Z(n520) );
  NAND2_X1 U569 ( .A1(n521), .A2(n520), .ZN(n528) );
  AND2_X1 U570 ( .A1(n522), .A2(G2105), .ZN(n876) );
  NAND2_X1 U571 ( .A1(G125), .A2(n876), .ZN(n526) );
  NOR2_X1 U572 ( .A1(G2104), .A2(G2105), .ZN(n523) );
  XOR2_X1 U573 ( .A(n523), .B(KEYINPUT17), .Z(n524) );
  NAND2_X1 U574 ( .A1(G137), .A2(n882), .ZN(n525) );
  NAND2_X1 U575 ( .A1(n526), .A2(n525), .ZN(n527) );
  NOR2_X1 U576 ( .A1(n528), .A2(n527), .ZN(G160) );
  NAND2_X1 U577 ( .A1(G138), .A2(n882), .ZN(n531) );
  NAND2_X1 U578 ( .A1(G126), .A2(n876), .ZN(n529) );
  XOR2_X1 U579 ( .A(KEYINPUT93), .B(n529), .Z(n530) );
  NAND2_X1 U580 ( .A1(n531), .A2(n530), .ZN(n535) );
  NAND2_X1 U581 ( .A1(G114), .A2(n877), .ZN(n533) );
  NAND2_X1 U582 ( .A1(G102), .A2(n881), .ZN(n532) );
  NAND2_X1 U583 ( .A1(n533), .A2(n532), .ZN(n534) );
  NOR2_X1 U584 ( .A1(n535), .A2(n534), .ZN(G164) );
  XOR2_X1 U585 ( .A(KEYINPUT0), .B(G543), .Z(n571) );
  INV_X1 U586 ( .A(G651), .ZN(n536) );
  NOR2_X2 U587 ( .A1(n571), .A2(n536), .ZN(n784) );
  NAND2_X1 U588 ( .A1(G78), .A2(n784), .ZN(n539) );
  NOR2_X1 U589 ( .A1(G543), .A2(n536), .ZN(n537) );
  XOR2_X1 U590 ( .A(KEYINPUT1), .B(n537), .Z(n787) );
  NAND2_X1 U591 ( .A1(G65), .A2(n787), .ZN(n538) );
  NAND2_X1 U592 ( .A1(n539), .A2(n538), .ZN(n542) );
  NOR2_X1 U593 ( .A1(G651), .A2(G543), .ZN(n783) );
  NAND2_X1 U594 ( .A1(n783), .A2(G91), .ZN(n540) );
  XOR2_X1 U595 ( .A(KEYINPUT68), .B(n540), .Z(n541) );
  NOR2_X1 U596 ( .A1(n542), .A2(n541), .ZN(n544) );
  NAND2_X1 U597 ( .A1(n788), .A2(G53), .ZN(n543) );
  NAND2_X1 U598 ( .A1(n544), .A2(n543), .ZN(G299) );
  NAND2_X1 U599 ( .A1(G64), .A2(n787), .ZN(n546) );
  NAND2_X1 U600 ( .A1(G52), .A2(n788), .ZN(n545) );
  NAND2_X1 U601 ( .A1(n546), .A2(n545), .ZN(n551) );
  NAND2_X1 U602 ( .A1(G90), .A2(n783), .ZN(n548) );
  NAND2_X1 U603 ( .A1(G77), .A2(n784), .ZN(n547) );
  NAND2_X1 U604 ( .A1(n548), .A2(n547), .ZN(n549) );
  XOR2_X1 U605 ( .A(KEYINPUT9), .B(n549), .Z(n550) );
  NOR2_X1 U606 ( .A1(n551), .A2(n550), .ZN(G171) );
  NAND2_X1 U607 ( .A1(n783), .A2(G89), .ZN(n552) );
  XOR2_X1 U608 ( .A(KEYINPUT4), .B(n552), .Z(n555) );
  NAND2_X1 U609 ( .A1(n784), .A2(G76), .ZN(n553) );
  XOR2_X1 U610 ( .A(KEYINPUT78), .B(n553), .Z(n554) );
  NOR2_X1 U611 ( .A1(n555), .A2(n554), .ZN(n556) );
  XNOR2_X1 U612 ( .A(KEYINPUT5), .B(n556), .ZN(n557) );
  XNOR2_X1 U613 ( .A(n557), .B(KEYINPUT79), .ZN(n562) );
  NAND2_X1 U614 ( .A1(G63), .A2(n787), .ZN(n559) );
  NAND2_X1 U615 ( .A1(G51), .A2(n788), .ZN(n558) );
  NAND2_X1 U616 ( .A1(n559), .A2(n558), .ZN(n560) );
  XOR2_X1 U617 ( .A(KEYINPUT6), .B(n560), .Z(n561) );
  NAND2_X1 U618 ( .A1(n562), .A2(n561), .ZN(n563) );
  XNOR2_X1 U619 ( .A(KEYINPUT7), .B(n563), .ZN(G168) );
  XOR2_X1 U620 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U621 ( .A1(G75), .A2(n784), .ZN(n565) );
  NAND2_X1 U622 ( .A1(G62), .A2(n787), .ZN(n564) );
  NAND2_X1 U623 ( .A1(n565), .A2(n564), .ZN(n568) );
  NAND2_X1 U624 ( .A1(n783), .A2(G88), .ZN(n566) );
  XOR2_X1 U625 ( .A(KEYINPUT88), .B(n566), .Z(n567) );
  NOR2_X1 U626 ( .A1(n568), .A2(n567), .ZN(n570) );
  NAND2_X1 U627 ( .A1(n788), .A2(G50), .ZN(n569) );
  NAND2_X1 U628 ( .A1(n570), .A2(n569), .ZN(G303) );
  NAND2_X1 U629 ( .A1(G74), .A2(G651), .ZN(n576) );
  NAND2_X1 U630 ( .A1(G49), .A2(n788), .ZN(n573) );
  NAND2_X1 U631 ( .A1(G87), .A2(n571), .ZN(n572) );
  NAND2_X1 U632 ( .A1(n573), .A2(n572), .ZN(n574) );
  NOR2_X1 U633 ( .A1(n787), .A2(n574), .ZN(n575) );
  NAND2_X1 U634 ( .A1(n576), .A2(n575), .ZN(n577) );
  XNOR2_X1 U635 ( .A(n577), .B(KEYINPUT84), .ZN(G288) );
  NAND2_X1 U636 ( .A1(G86), .A2(n783), .ZN(n579) );
  NAND2_X1 U637 ( .A1(G61), .A2(n787), .ZN(n578) );
  NAND2_X1 U638 ( .A1(n579), .A2(n578), .ZN(n580) );
  XOR2_X1 U639 ( .A(KEYINPUT85), .B(n580), .Z(n585) );
  XOR2_X1 U640 ( .A(KEYINPUT2), .B(KEYINPUT87), .Z(n582) );
  NAND2_X1 U641 ( .A1(G73), .A2(n784), .ZN(n581) );
  XNOR2_X1 U642 ( .A(n582), .B(n581), .ZN(n583) );
  XOR2_X1 U643 ( .A(KEYINPUT86), .B(n583), .Z(n584) );
  NOR2_X1 U644 ( .A1(n585), .A2(n584), .ZN(n587) );
  NAND2_X1 U645 ( .A1(n788), .A2(G48), .ZN(n586) );
  NAND2_X1 U646 ( .A1(n587), .A2(n586), .ZN(G305) );
  NAND2_X1 U647 ( .A1(G85), .A2(n783), .ZN(n589) );
  NAND2_X1 U648 ( .A1(G72), .A2(n784), .ZN(n588) );
  NAND2_X1 U649 ( .A1(n589), .A2(n588), .ZN(n590) );
  XNOR2_X1 U650 ( .A(KEYINPUT67), .B(n590), .ZN(n594) );
  NAND2_X1 U651 ( .A1(G60), .A2(n787), .ZN(n592) );
  NAND2_X1 U652 ( .A1(G47), .A2(n788), .ZN(n591) );
  AND2_X1 U653 ( .A1(n592), .A2(n591), .ZN(n593) );
  NAND2_X1 U654 ( .A1(n594), .A2(n593), .ZN(G290) );
  NAND2_X1 U655 ( .A1(G54), .A2(n788), .ZN(n600) );
  NAND2_X1 U656 ( .A1(G92), .A2(n783), .ZN(n596) );
  NAND2_X1 U657 ( .A1(G66), .A2(n787), .ZN(n595) );
  NAND2_X1 U658 ( .A1(n596), .A2(n595), .ZN(n598) );
  NAND2_X1 U659 ( .A1(n784), .A2(G79), .ZN(n597) );
  NOR2_X1 U660 ( .A1(n598), .A2(n513), .ZN(n599) );
  NAND2_X1 U661 ( .A1(n600), .A2(n599), .ZN(n601) );
  XNOR2_X1 U662 ( .A(n601), .B(KEYINPUT15), .ZN(n602) );
  XNOR2_X1 U663 ( .A(KEYINPUT74), .B(KEYINPUT75), .ZN(n608) );
  NAND2_X1 U664 ( .A1(n783), .A2(G81), .ZN(n603) );
  XNOR2_X1 U665 ( .A(n603), .B(KEYINPUT12), .ZN(n605) );
  NAND2_X1 U666 ( .A1(G68), .A2(n784), .ZN(n604) );
  NAND2_X1 U667 ( .A1(n605), .A2(n604), .ZN(n606) );
  XNOR2_X1 U668 ( .A(n606), .B(KEYINPUT13), .ZN(n607) );
  XNOR2_X1 U669 ( .A(n608), .B(n607), .ZN(n611) );
  NAND2_X1 U670 ( .A1(n787), .A2(G56), .ZN(n609) );
  XOR2_X1 U671 ( .A(KEYINPUT14), .B(n609), .Z(n610) );
  NOR2_X1 U672 ( .A1(n611), .A2(n610), .ZN(n613) );
  NAND2_X1 U673 ( .A1(n788), .A2(G43), .ZN(n612) );
  NAND2_X1 U674 ( .A1(n613), .A2(n612), .ZN(n912) );
  NOR2_X1 U675 ( .A1(G164), .A2(G1384), .ZN(n680) );
  NAND2_X1 U676 ( .A1(G160), .A2(G40), .ZN(n679) );
  INV_X1 U677 ( .A(n679), .ZN(n614) );
  INV_X1 U678 ( .A(G1996), .ZN(n959) );
  NOR2_X1 U679 ( .A1(n656), .A2(n959), .ZN(n615) );
  XOR2_X1 U680 ( .A(n615), .B(KEYINPUT26), .Z(n617) );
  NAND2_X1 U681 ( .A1(n656), .A2(G1341), .ZN(n616) );
  NAND2_X1 U682 ( .A1(n617), .A2(n616), .ZN(n618) );
  NOR2_X1 U683 ( .A1(n906), .A2(n620), .ZN(n619) );
  XNOR2_X1 U684 ( .A(KEYINPUT101), .B(n619), .ZN(n627) );
  NAND2_X1 U685 ( .A1(n906), .A2(n620), .ZN(n624) );
  NAND2_X1 U686 ( .A1(n656), .A2(G1348), .ZN(n622) );
  XOR2_X1 U687 ( .A(n656), .B(KEYINPUT98), .Z(n642) );
  NAND2_X1 U688 ( .A1(G2067), .A2(n642), .ZN(n621) );
  NAND2_X1 U689 ( .A1(n622), .A2(n621), .ZN(n623) );
  NAND2_X1 U690 ( .A1(n624), .A2(n623), .ZN(n625) );
  XNOR2_X1 U691 ( .A(n625), .B(KEYINPUT100), .ZN(n626) );
  NAND2_X1 U692 ( .A1(n627), .A2(n626), .ZN(n633) );
  INV_X1 U693 ( .A(G299), .ZN(n909) );
  NAND2_X1 U694 ( .A1(G2072), .A2(n642), .ZN(n628) );
  XNOR2_X1 U695 ( .A(n628), .B(KEYINPUT27), .ZN(n631) );
  INV_X1 U696 ( .A(G1956), .ZN(n629) );
  NOR2_X1 U697 ( .A1(n642), .A2(n629), .ZN(n630) );
  NOR2_X1 U698 ( .A1(n631), .A2(n630), .ZN(n634) );
  NAND2_X1 U699 ( .A1(n909), .A2(n634), .ZN(n632) );
  NAND2_X1 U700 ( .A1(n633), .A2(n632), .ZN(n638) );
  NOR2_X1 U701 ( .A1(n909), .A2(n634), .ZN(n636) );
  XNOR2_X1 U702 ( .A(KEYINPUT28), .B(KEYINPUT99), .ZN(n635) );
  XNOR2_X1 U703 ( .A(n636), .B(n635), .ZN(n637) );
  NAND2_X1 U704 ( .A1(n638), .A2(n637), .ZN(n641) );
  XNOR2_X1 U705 ( .A(KEYINPUT102), .B(KEYINPUT103), .ZN(n639) );
  XNOR2_X1 U706 ( .A(n639), .B(KEYINPUT29), .ZN(n640) );
  XNOR2_X1 U707 ( .A(n641), .B(n640), .ZN(n646) );
  XNOR2_X1 U708 ( .A(KEYINPUT25), .B(G2078), .ZN(n965) );
  NAND2_X1 U709 ( .A1(n642), .A2(n965), .ZN(n644) );
  INV_X1 U710 ( .A(G1961), .ZN(n929) );
  NAND2_X1 U711 ( .A1(n929), .A2(n656), .ZN(n643) );
  NAND2_X1 U712 ( .A1(n644), .A2(n643), .ZN(n650) );
  NAND2_X1 U713 ( .A1(n650), .A2(G171), .ZN(n645) );
  NAND2_X1 U714 ( .A1(n646), .A2(n645), .ZN(n655) );
  NAND2_X1 U715 ( .A1(G8), .A2(n656), .ZN(n694) );
  NOR2_X1 U716 ( .A1(G1966), .A2(n694), .ZN(n669) );
  NOR2_X1 U717 ( .A1(G2084), .A2(n656), .ZN(n666) );
  NOR2_X1 U718 ( .A1(n669), .A2(n666), .ZN(n647) );
  NAND2_X1 U719 ( .A1(G8), .A2(n647), .ZN(n648) );
  XNOR2_X1 U720 ( .A(KEYINPUT30), .B(n648), .ZN(n649) );
  NOR2_X1 U721 ( .A1(G168), .A2(n649), .ZN(n652) );
  NOR2_X1 U722 ( .A1(G171), .A2(n650), .ZN(n651) );
  NOR2_X1 U723 ( .A1(n652), .A2(n651), .ZN(n653) );
  XOR2_X1 U724 ( .A(KEYINPUT31), .B(n653), .Z(n654) );
  NAND2_X1 U725 ( .A1(n655), .A2(n654), .ZN(n667) );
  NAND2_X1 U726 ( .A1(n667), .A2(G286), .ZN(n664) );
  INV_X1 U727 ( .A(G8), .ZN(n662) );
  NOR2_X1 U728 ( .A1(G1971), .A2(n694), .ZN(n658) );
  NOR2_X1 U729 ( .A1(G2090), .A2(n656), .ZN(n657) );
  NOR2_X1 U730 ( .A1(n658), .A2(n657), .ZN(n659) );
  XNOR2_X1 U731 ( .A(n659), .B(KEYINPUT104), .ZN(n660) );
  NAND2_X1 U732 ( .A1(n660), .A2(G303), .ZN(n661) );
  OR2_X1 U733 ( .A1(n662), .A2(n661), .ZN(n663) );
  AND2_X1 U734 ( .A1(n664), .A2(n663), .ZN(n665) );
  XNOR2_X1 U735 ( .A(KEYINPUT32), .B(n665), .ZN(n673) );
  NAND2_X1 U736 ( .A1(G8), .A2(n666), .ZN(n671) );
  INV_X1 U737 ( .A(n667), .ZN(n668) );
  NOR2_X1 U738 ( .A1(n669), .A2(n668), .ZN(n670) );
  NAND2_X1 U739 ( .A1(n671), .A2(n670), .ZN(n672) );
  NOR2_X1 U740 ( .A1(G1976), .A2(G288), .ZN(n682) );
  NOR2_X1 U741 ( .A1(G1971), .A2(G303), .ZN(n674) );
  NOR2_X1 U742 ( .A1(n682), .A2(n674), .ZN(n904) );
  NAND2_X1 U743 ( .A1(n689), .A2(n904), .ZN(n676) );
  NAND2_X1 U744 ( .A1(G288), .A2(G1976), .ZN(n675) );
  XOR2_X1 U745 ( .A(KEYINPUT105), .B(n675), .Z(n915) );
  NAND2_X1 U746 ( .A1(n676), .A2(n915), .ZN(n677) );
  NOR2_X1 U747 ( .A1(n677), .A2(n694), .ZN(n678) );
  NOR2_X1 U748 ( .A1(n678), .A2(KEYINPUT33), .ZN(n686) );
  XOR2_X1 U749 ( .A(G1981), .B(G305), .Z(n917) );
  NOR2_X1 U750 ( .A1(n680), .A2(n679), .ZN(n742) );
  XNOR2_X1 U751 ( .A(G1986), .B(G290), .ZN(n908) );
  NAND2_X1 U752 ( .A1(n742), .A2(n908), .ZN(n681) );
  XNOR2_X1 U753 ( .A(KEYINPUT94), .B(n681), .ZN(n698) );
  AND2_X1 U754 ( .A1(n917), .A2(n698), .ZN(n684) );
  NAND2_X1 U755 ( .A1(n682), .A2(KEYINPUT33), .ZN(n683) );
  NOR2_X1 U756 ( .A1(G2090), .A2(G303), .ZN(n687) );
  NAND2_X1 U757 ( .A1(G8), .A2(n687), .ZN(n688) );
  XNOR2_X1 U758 ( .A(n688), .B(KEYINPUT106), .ZN(n690) );
  NAND2_X1 U759 ( .A1(n690), .A2(n689), .ZN(n691) );
  NAND2_X1 U760 ( .A1(n691), .A2(n694), .ZN(n696) );
  NOR2_X1 U761 ( .A1(G1981), .A2(G305), .ZN(n692) );
  XOR2_X1 U762 ( .A(n692), .B(KEYINPUT24), .Z(n693) );
  OR2_X1 U763 ( .A1(n694), .A2(n693), .ZN(n695) );
  NAND2_X1 U764 ( .A1(n696), .A2(n695), .ZN(n697) );
  NAND2_X1 U765 ( .A1(n516), .A2(n515), .ZN(n728) );
  NAND2_X1 U766 ( .A1(G119), .A2(n876), .ZN(n700) );
  NAND2_X1 U767 ( .A1(G107), .A2(n877), .ZN(n699) );
  NAND2_X1 U768 ( .A1(n700), .A2(n699), .ZN(n701) );
  XNOR2_X1 U769 ( .A(KEYINPUT97), .B(n701), .ZN(n705) );
  NAND2_X1 U770 ( .A1(n882), .A2(G131), .ZN(n703) );
  NAND2_X1 U771 ( .A1(n881), .A2(G95), .ZN(n702) );
  AND2_X1 U772 ( .A1(n703), .A2(n702), .ZN(n704) );
  NAND2_X1 U773 ( .A1(n705), .A2(n704), .ZN(n871) );
  NAND2_X1 U774 ( .A1(G1991), .A2(n871), .ZN(n714) );
  NAND2_X1 U775 ( .A1(G129), .A2(n876), .ZN(n707) );
  NAND2_X1 U776 ( .A1(G141), .A2(n882), .ZN(n706) );
  NAND2_X1 U777 ( .A1(n707), .A2(n706), .ZN(n710) );
  NAND2_X1 U778 ( .A1(n881), .A2(G105), .ZN(n708) );
  XOR2_X1 U779 ( .A(KEYINPUT38), .B(n708), .Z(n709) );
  NOR2_X1 U780 ( .A1(n710), .A2(n709), .ZN(n712) );
  NAND2_X1 U781 ( .A1(n877), .A2(G117), .ZN(n711) );
  NAND2_X1 U782 ( .A1(n712), .A2(n711), .ZN(n869) );
  NAND2_X1 U783 ( .A1(G1996), .A2(n869), .ZN(n713) );
  NAND2_X1 U784 ( .A1(n714), .A2(n713), .ZN(n978) );
  NAND2_X1 U785 ( .A1(n978), .A2(n742), .ZN(n726) );
  XOR2_X1 U786 ( .A(G2067), .B(KEYINPUT37), .Z(n740) );
  NAND2_X1 U787 ( .A1(G128), .A2(n876), .ZN(n716) );
  NAND2_X1 U788 ( .A1(G116), .A2(n877), .ZN(n715) );
  NAND2_X1 U789 ( .A1(n716), .A2(n715), .ZN(n717) );
  XOR2_X1 U790 ( .A(KEYINPUT35), .B(n717), .Z(n724) );
  NAND2_X1 U791 ( .A1(G104), .A2(n881), .ZN(n720) );
  NAND2_X1 U792 ( .A1(G140), .A2(n882), .ZN(n718) );
  XOR2_X1 U793 ( .A(KEYINPUT95), .B(n718), .Z(n719) );
  NAND2_X1 U794 ( .A1(n720), .A2(n719), .ZN(n721) );
  XNOR2_X1 U795 ( .A(n721), .B(KEYINPUT34), .ZN(n722) );
  XNOR2_X1 U796 ( .A(n722), .B(KEYINPUT96), .ZN(n723) );
  NOR2_X1 U797 ( .A1(n724), .A2(n723), .ZN(n725) );
  XOR2_X1 U798 ( .A(KEYINPUT36), .B(n725), .Z(n889) );
  AND2_X1 U799 ( .A1(n740), .A2(n889), .ZN(n979) );
  NAND2_X1 U800 ( .A1(n979), .A2(n742), .ZN(n729) );
  AND2_X1 U801 ( .A1(n726), .A2(n729), .ZN(n727) );
  NAND2_X1 U802 ( .A1(n728), .A2(n727), .ZN(n739) );
  INV_X1 U803 ( .A(n729), .ZN(n737) );
  NOR2_X1 U804 ( .A1(G1996), .A2(n869), .ZN(n988) );
  NOR2_X1 U805 ( .A1(G1986), .A2(G290), .ZN(n730) );
  NOR2_X1 U806 ( .A1(G1991), .A2(n871), .ZN(n983) );
  NOR2_X1 U807 ( .A1(n730), .A2(n983), .ZN(n731) );
  XOR2_X1 U808 ( .A(KEYINPUT107), .B(n731), .Z(n732) );
  NOR2_X1 U809 ( .A1(n978), .A2(n732), .ZN(n733) );
  NOR2_X1 U810 ( .A1(n988), .A2(n733), .ZN(n734) );
  XNOR2_X1 U811 ( .A(KEYINPUT39), .B(n734), .ZN(n735) );
  NAND2_X1 U812 ( .A1(n735), .A2(n742), .ZN(n736) );
  OR2_X1 U813 ( .A1(n737), .A2(n736), .ZN(n738) );
  AND2_X1 U814 ( .A1(n739), .A2(n738), .ZN(n744) );
  NOR2_X1 U815 ( .A1(n889), .A2(n740), .ZN(n741) );
  XNOR2_X1 U816 ( .A(n741), .B(KEYINPUT108), .ZN(n997) );
  NAND2_X1 U817 ( .A1(n997), .A2(n742), .ZN(n743) );
  NAND2_X1 U818 ( .A1(n744), .A2(n743), .ZN(n745) );
  XNOR2_X1 U819 ( .A(n745), .B(KEYINPUT40), .ZN(G329) );
  XOR2_X1 U820 ( .A(G2435), .B(G2454), .Z(n747) );
  XNOR2_X1 U821 ( .A(G2430), .B(G2438), .ZN(n746) );
  XNOR2_X1 U822 ( .A(n747), .B(n746), .ZN(n754) );
  XOR2_X1 U823 ( .A(G2446), .B(KEYINPUT109), .Z(n749) );
  XNOR2_X1 U824 ( .A(G2451), .B(G2443), .ZN(n748) );
  XNOR2_X1 U825 ( .A(n749), .B(n748), .ZN(n750) );
  XOR2_X1 U826 ( .A(n750), .B(G2427), .Z(n752) );
  XNOR2_X1 U827 ( .A(G1341), .B(G1348), .ZN(n751) );
  XNOR2_X1 U828 ( .A(n752), .B(n751), .ZN(n753) );
  XNOR2_X1 U829 ( .A(n754), .B(n753), .ZN(n755) );
  AND2_X1 U830 ( .A1(n755), .A2(G14), .ZN(G401) );
  AND2_X1 U831 ( .A1(G452), .A2(G94), .ZN(G173) );
  XOR2_X1 U832 ( .A(KEYINPUT73), .B(KEYINPUT10), .Z(n757) );
  NAND2_X1 U833 ( .A1(G7), .A2(G661), .ZN(n756) );
  XNOR2_X1 U834 ( .A(n757), .B(n756), .ZN(n758) );
  XNOR2_X1 U835 ( .A(KEYINPUT72), .B(n758), .ZN(G223) );
  INV_X1 U836 ( .A(G223), .ZN(n822) );
  NAND2_X1 U837 ( .A1(n822), .A2(G567), .ZN(n759) );
  XOR2_X1 U838 ( .A(KEYINPUT11), .B(n759), .Z(G234) );
  INV_X1 U839 ( .A(G860), .ZN(n782) );
  OR2_X1 U840 ( .A1(n912), .A2(n782), .ZN(G153) );
  INV_X1 U841 ( .A(G171), .ZN(G301) );
  NAND2_X1 U842 ( .A1(G868), .A2(G301), .ZN(n761) );
  OR2_X1 U843 ( .A1(n906), .A2(G868), .ZN(n760) );
  NAND2_X1 U844 ( .A1(n761), .A2(n760), .ZN(G284) );
  INV_X1 U845 ( .A(G868), .ZN(n802) );
  NOR2_X1 U846 ( .A1(G286), .A2(n802), .ZN(n763) );
  NOR2_X1 U847 ( .A1(G868), .A2(G299), .ZN(n762) );
  NOR2_X1 U848 ( .A1(n763), .A2(n762), .ZN(G297) );
  NAND2_X1 U849 ( .A1(n782), .A2(G559), .ZN(n764) );
  NAND2_X1 U850 ( .A1(n764), .A2(n906), .ZN(n765) );
  XNOR2_X1 U851 ( .A(n765), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U852 ( .A1(G868), .A2(n912), .ZN(n768) );
  NAND2_X1 U853 ( .A1(G868), .A2(n906), .ZN(n766) );
  NOR2_X1 U854 ( .A1(G559), .A2(n766), .ZN(n767) );
  NOR2_X1 U855 ( .A1(n768), .A2(n767), .ZN(n769) );
  XNOR2_X1 U856 ( .A(KEYINPUT80), .B(n769), .ZN(G282) );
  NAND2_X1 U857 ( .A1(G123), .A2(n876), .ZN(n770) );
  XNOR2_X1 U858 ( .A(n770), .B(KEYINPUT18), .ZN(n777) );
  NAND2_X1 U859 ( .A1(n881), .A2(G99), .ZN(n772) );
  NAND2_X1 U860 ( .A1(G135), .A2(n882), .ZN(n771) );
  NAND2_X1 U861 ( .A1(n772), .A2(n771), .ZN(n775) );
  NAND2_X1 U862 ( .A1(G111), .A2(n877), .ZN(n773) );
  XNOR2_X1 U863 ( .A(KEYINPUT81), .B(n773), .ZN(n774) );
  NOR2_X1 U864 ( .A1(n775), .A2(n774), .ZN(n776) );
  NAND2_X1 U865 ( .A1(n777), .A2(n776), .ZN(n980) );
  XNOR2_X1 U866 ( .A(G2096), .B(n980), .ZN(n778) );
  NOR2_X1 U867 ( .A1(G2100), .A2(n778), .ZN(n779) );
  XOR2_X1 U868 ( .A(KEYINPUT82), .B(n779), .Z(G156) );
  XNOR2_X1 U869 ( .A(n912), .B(KEYINPUT83), .ZN(n781) );
  NAND2_X1 U870 ( .A1(n906), .A2(G559), .ZN(n780) );
  XNOR2_X1 U871 ( .A(n781), .B(n780), .ZN(n799) );
  NAND2_X1 U872 ( .A1(n782), .A2(n799), .ZN(n793) );
  NAND2_X1 U873 ( .A1(G93), .A2(n783), .ZN(n786) );
  NAND2_X1 U874 ( .A1(G80), .A2(n784), .ZN(n785) );
  NAND2_X1 U875 ( .A1(n786), .A2(n785), .ZN(n792) );
  NAND2_X1 U876 ( .A1(G67), .A2(n787), .ZN(n790) );
  NAND2_X1 U877 ( .A1(G55), .A2(n788), .ZN(n789) );
  NAND2_X1 U878 ( .A1(n790), .A2(n789), .ZN(n791) );
  NOR2_X1 U879 ( .A1(n792), .A2(n791), .ZN(n801) );
  XOR2_X1 U880 ( .A(n793), .B(n801), .Z(G145) );
  XNOR2_X1 U881 ( .A(n801), .B(G303), .ZN(n794) );
  XNOR2_X1 U882 ( .A(n794), .B(G305), .ZN(n795) );
  XOR2_X1 U883 ( .A(n795), .B(KEYINPUT19), .Z(n797) );
  XNOR2_X1 U884 ( .A(n909), .B(G288), .ZN(n796) );
  XNOR2_X1 U885 ( .A(n797), .B(n796), .ZN(n798) );
  XNOR2_X1 U886 ( .A(n798), .B(G290), .ZN(n895) );
  XOR2_X1 U887 ( .A(n895), .B(n799), .Z(n800) );
  NOR2_X1 U888 ( .A1(n802), .A2(n800), .ZN(n804) );
  AND2_X1 U889 ( .A1(n802), .A2(n801), .ZN(n803) );
  NOR2_X1 U890 ( .A1(n804), .A2(n803), .ZN(G295) );
  NAND2_X1 U891 ( .A1(G2078), .A2(G2084), .ZN(n805) );
  XOR2_X1 U892 ( .A(KEYINPUT20), .B(n805), .Z(n806) );
  NAND2_X1 U893 ( .A1(G2090), .A2(n806), .ZN(n807) );
  XNOR2_X1 U894 ( .A(KEYINPUT21), .B(n807), .ZN(n808) );
  NAND2_X1 U895 ( .A1(n808), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U896 ( .A(KEYINPUT69), .B(G57), .ZN(G237) );
  XOR2_X1 U897 ( .A(KEYINPUT70), .B(G132), .Z(G219) );
  XNOR2_X1 U898 ( .A(KEYINPUT71), .B(G82), .ZN(G220) );
  XNOR2_X1 U899 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NAND2_X1 U900 ( .A1(G120), .A2(G108), .ZN(n809) );
  NOR2_X1 U901 ( .A1(G237), .A2(n809), .ZN(n810) );
  NAND2_X1 U902 ( .A1(G69), .A2(n810), .ZN(n828) );
  NAND2_X1 U903 ( .A1(G567), .A2(n828), .ZN(n818) );
  NOR2_X1 U904 ( .A1(G219), .A2(G220), .ZN(n812) );
  XNOR2_X1 U905 ( .A(KEYINPUT22), .B(KEYINPUT89), .ZN(n811) );
  XNOR2_X1 U906 ( .A(n812), .B(n811), .ZN(n813) );
  NOR2_X1 U907 ( .A1(n813), .A2(G218), .ZN(n814) );
  NAND2_X1 U908 ( .A1(G96), .A2(n814), .ZN(n815) );
  XNOR2_X1 U909 ( .A(KEYINPUT90), .B(n815), .ZN(n829) );
  NAND2_X1 U910 ( .A1(n829), .A2(G2106), .ZN(n816) );
  XOR2_X1 U911 ( .A(KEYINPUT91), .B(n816), .Z(n817) );
  NAND2_X1 U912 ( .A1(n818), .A2(n817), .ZN(n819) );
  XOR2_X1 U913 ( .A(KEYINPUT92), .B(n819), .Z(G319) );
  INV_X1 U914 ( .A(G319), .ZN(n821) );
  NAND2_X1 U915 ( .A1(G661), .A2(G483), .ZN(n820) );
  NOR2_X1 U916 ( .A1(n821), .A2(n820), .ZN(n827) );
  NAND2_X1 U917 ( .A1(n827), .A2(G36), .ZN(G176) );
  NAND2_X1 U918 ( .A1(G2106), .A2(n822), .ZN(G217) );
  INV_X1 U919 ( .A(G661), .ZN(n824) );
  NAND2_X1 U920 ( .A1(G2), .A2(G15), .ZN(n823) );
  NOR2_X1 U921 ( .A1(n824), .A2(n823), .ZN(n825) );
  XOR2_X1 U922 ( .A(KEYINPUT110), .B(n825), .Z(G259) );
  NAND2_X1 U923 ( .A1(G3), .A2(G1), .ZN(n826) );
  NAND2_X1 U924 ( .A1(n827), .A2(n826), .ZN(G188) );
  XNOR2_X1 U925 ( .A(G108), .B(KEYINPUT119), .ZN(G238) );
  INV_X1 U927 ( .A(G120), .ZN(G236) );
  INV_X1 U928 ( .A(G96), .ZN(G221) );
  INV_X1 U929 ( .A(G69), .ZN(G235) );
  NOR2_X1 U930 ( .A1(n829), .A2(n828), .ZN(G325) );
  INV_X1 U931 ( .A(G325), .ZN(G261) );
  XOR2_X1 U932 ( .A(G2100), .B(G2096), .Z(n831) );
  XNOR2_X1 U933 ( .A(KEYINPUT42), .B(G2678), .ZN(n830) );
  XNOR2_X1 U934 ( .A(n831), .B(n830), .ZN(n835) );
  XOR2_X1 U935 ( .A(KEYINPUT43), .B(G2090), .Z(n833) );
  XNOR2_X1 U936 ( .A(G2067), .B(G2072), .ZN(n832) );
  XNOR2_X1 U937 ( .A(n833), .B(n832), .ZN(n834) );
  XOR2_X1 U938 ( .A(n835), .B(n834), .Z(n837) );
  XNOR2_X1 U939 ( .A(G2078), .B(G2084), .ZN(n836) );
  XNOR2_X1 U940 ( .A(n837), .B(n836), .ZN(G227) );
  XOR2_X1 U941 ( .A(KEYINPUT112), .B(G1961), .Z(n839) );
  XNOR2_X1 U942 ( .A(G1996), .B(G1991), .ZN(n838) );
  XNOR2_X1 U943 ( .A(n839), .B(n838), .ZN(n840) );
  XOR2_X1 U944 ( .A(n840), .B(KEYINPUT41), .Z(n842) );
  XNOR2_X1 U945 ( .A(G1966), .B(G1981), .ZN(n841) );
  XNOR2_X1 U946 ( .A(n842), .B(n841), .ZN(n846) );
  XOR2_X1 U947 ( .A(G1976), .B(G1971), .Z(n844) );
  XNOR2_X1 U948 ( .A(G1986), .B(G1956), .ZN(n843) );
  XNOR2_X1 U949 ( .A(n844), .B(n843), .ZN(n845) );
  XOR2_X1 U950 ( .A(n846), .B(n845), .Z(n848) );
  XNOR2_X1 U951 ( .A(KEYINPUT111), .B(G2474), .ZN(n847) );
  XNOR2_X1 U952 ( .A(n848), .B(n847), .ZN(G229) );
  NAND2_X1 U953 ( .A1(G124), .A2(n876), .ZN(n849) );
  XOR2_X1 U954 ( .A(KEYINPUT44), .B(n849), .Z(n850) );
  XNOR2_X1 U955 ( .A(n850), .B(KEYINPUT113), .ZN(n852) );
  NAND2_X1 U956 ( .A1(G136), .A2(n882), .ZN(n851) );
  NAND2_X1 U957 ( .A1(n852), .A2(n851), .ZN(n853) );
  XOR2_X1 U958 ( .A(KEYINPUT114), .B(n853), .Z(n855) );
  NAND2_X1 U959 ( .A1(n881), .A2(G100), .ZN(n854) );
  NAND2_X1 U960 ( .A1(n855), .A2(n854), .ZN(n858) );
  NAND2_X1 U961 ( .A1(G112), .A2(n877), .ZN(n856) );
  XNOR2_X1 U962 ( .A(KEYINPUT115), .B(n856), .ZN(n857) );
  NOR2_X1 U963 ( .A1(n858), .A2(n857), .ZN(G162) );
  XOR2_X1 U964 ( .A(KEYINPUT48), .B(KEYINPUT46), .Z(n868) );
  NAND2_X1 U965 ( .A1(G130), .A2(n876), .ZN(n860) );
  NAND2_X1 U966 ( .A1(G118), .A2(n877), .ZN(n859) );
  NAND2_X1 U967 ( .A1(n860), .A2(n859), .ZN(n865) );
  NAND2_X1 U968 ( .A1(n881), .A2(G106), .ZN(n862) );
  NAND2_X1 U969 ( .A1(G142), .A2(n882), .ZN(n861) );
  NAND2_X1 U970 ( .A1(n862), .A2(n861), .ZN(n863) );
  XOR2_X1 U971 ( .A(KEYINPUT45), .B(n863), .Z(n864) );
  NOR2_X1 U972 ( .A1(n865), .A2(n864), .ZN(n866) );
  XNOR2_X1 U973 ( .A(G164), .B(n866), .ZN(n867) );
  XNOR2_X1 U974 ( .A(n868), .B(n867), .ZN(n870) );
  XNOR2_X1 U975 ( .A(n870), .B(n869), .ZN(n872) );
  XNOR2_X1 U976 ( .A(n872), .B(n871), .ZN(n873) );
  XNOR2_X1 U977 ( .A(n980), .B(n873), .ZN(n875) );
  XNOR2_X1 U978 ( .A(G160), .B(G162), .ZN(n874) );
  XNOR2_X1 U979 ( .A(n875), .B(n874), .ZN(n891) );
  NAND2_X1 U980 ( .A1(G127), .A2(n876), .ZN(n879) );
  NAND2_X1 U981 ( .A1(G115), .A2(n877), .ZN(n878) );
  NAND2_X1 U982 ( .A1(n879), .A2(n878), .ZN(n880) );
  XNOR2_X1 U983 ( .A(n880), .B(KEYINPUT47), .ZN(n887) );
  NAND2_X1 U984 ( .A1(n881), .A2(G103), .ZN(n884) );
  NAND2_X1 U985 ( .A1(G139), .A2(n882), .ZN(n883) );
  NAND2_X1 U986 ( .A1(n884), .A2(n883), .ZN(n885) );
  XOR2_X1 U987 ( .A(KEYINPUT116), .B(n885), .Z(n886) );
  NAND2_X1 U988 ( .A1(n887), .A2(n886), .ZN(n888) );
  XNOR2_X1 U989 ( .A(n888), .B(KEYINPUT117), .ZN(n992) );
  XOR2_X1 U990 ( .A(n992), .B(n889), .Z(n890) );
  XNOR2_X1 U991 ( .A(n891), .B(n890), .ZN(n892) );
  NOR2_X1 U992 ( .A1(G37), .A2(n892), .ZN(G395) );
  XNOR2_X1 U993 ( .A(n912), .B(KEYINPUT118), .ZN(n894) );
  XNOR2_X1 U994 ( .A(G171), .B(n906), .ZN(n893) );
  XNOR2_X1 U995 ( .A(n894), .B(n893), .ZN(n897) );
  XOR2_X1 U996 ( .A(G286), .B(n895), .Z(n896) );
  XNOR2_X1 U997 ( .A(n897), .B(n896), .ZN(n898) );
  NOR2_X1 U998 ( .A1(G37), .A2(n898), .ZN(G397) );
  NOR2_X1 U999 ( .A1(G227), .A2(G229), .ZN(n899) );
  XNOR2_X1 U1000 ( .A(KEYINPUT49), .B(n899), .ZN(n900) );
  NOR2_X1 U1001 ( .A1(G401), .A2(n900), .ZN(n901) );
  AND2_X1 U1002 ( .A1(n901), .A2(G319), .ZN(n903) );
  NOR2_X1 U1003 ( .A1(G395), .A2(G397), .ZN(n902) );
  NAND2_X1 U1004 ( .A1(n903), .A2(n902), .ZN(G225) );
  INV_X1 U1005 ( .A(G225), .ZN(G308) );
  INV_X1 U1006 ( .A(G303), .ZN(G166) );
  XNOR2_X1 U1007 ( .A(KEYINPUT56), .B(G16), .ZN(n928) );
  XNOR2_X1 U1008 ( .A(G171), .B(G1961), .ZN(n905) );
  NAND2_X1 U1009 ( .A1(n905), .A2(n904), .ZN(n925) );
  XOR2_X1 U1010 ( .A(n906), .B(G1348), .Z(n907) );
  NOR2_X1 U1011 ( .A1(n908), .A2(n907), .ZN(n923) );
  XNOR2_X1 U1012 ( .A(n909), .B(G1956), .ZN(n911) );
  NAND2_X1 U1013 ( .A1(G1971), .A2(G303), .ZN(n910) );
  NAND2_X1 U1014 ( .A1(n911), .A2(n910), .ZN(n914) );
  XNOR2_X1 U1015 ( .A(G1341), .B(n912), .ZN(n913) );
  NOR2_X1 U1016 ( .A1(n914), .A2(n913), .ZN(n916) );
  NAND2_X1 U1017 ( .A1(n916), .A2(n915), .ZN(n921) );
  XNOR2_X1 U1018 ( .A(G1966), .B(G168), .ZN(n918) );
  NAND2_X1 U1019 ( .A1(n918), .A2(n917), .ZN(n919) );
  XOR2_X1 U1020 ( .A(KEYINPUT57), .B(n919), .Z(n920) );
  NOR2_X1 U1021 ( .A1(n921), .A2(n920), .ZN(n922) );
  NAND2_X1 U1022 ( .A1(n923), .A2(n922), .ZN(n924) );
  NOR2_X1 U1023 ( .A1(n925), .A2(n924), .ZN(n926) );
  XNOR2_X1 U1024 ( .A(KEYINPUT125), .B(n926), .ZN(n927) );
  NAND2_X1 U1025 ( .A1(n928), .A2(n927), .ZN(n1007) );
  XNOR2_X1 U1026 ( .A(G5), .B(n929), .ZN(n938) );
  XNOR2_X1 U1027 ( .A(G1966), .B(G21), .ZN(n936) );
  XNOR2_X1 U1028 ( .A(G1986), .B(G24), .ZN(n931) );
  XNOR2_X1 U1029 ( .A(G1971), .B(G22), .ZN(n930) );
  NOR2_X1 U1030 ( .A1(n931), .A2(n930), .ZN(n933) );
  XOR2_X1 U1031 ( .A(G1976), .B(G23), .Z(n932) );
  NAND2_X1 U1032 ( .A1(n933), .A2(n932), .ZN(n934) );
  XNOR2_X1 U1033 ( .A(KEYINPUT58), .B(n934), .ZN(n935) );
  NOR2_X1 U1034 ( .A1(n936), .A2(n935), .ZN(n937) );
  NAND2_X1 U1035 ( .A1(n938), .A2(n937), .ZN(n950) );
  XOR2_X1 U1036 ( .A(G1348), .B(KEYINPUT59), .Z(n939) );
  XNOR2_X1 U1037 ( .A(G4), .B(n939), .ZN(n947) );
  XOR2_X1 U1038 ( .A(G1981), .B(G6), .Z(n942) );
  XOR2_X1 U1039 ( .A(KEYINPUT126), .B(G20), .Z(n940) );
  XNOR2_X1 U1040 ( .A(n940), .B(G1956), .ZN(n941) );
  NAND2_X1 U1041 ( .A1(n942), .A2(n941), .ZN(n944) );
  XNOR2_X1 U1042 ( .A(G19), .B(G1341), .ZN(n943) );
  NOR2_X1 U1043 ( .A1(n944), .A2(n943), .ZN(n945) );
  XNOR2_X1 U1044 ( .A(n945), .B(KEYINPUT127), .ZN(n946) );
  NOR2_X1 U1045 ( .A1(n947), .A2(n946), .ZN(n948) );
  XOR2_X1 U1046 ( .A(KEYINPUT60), .B(n948), .Z(n949) );
  NOR2_X1 U1047 ( .A1(n950), .A2(n949), .ZN(n951) );
  XNOR2_X1 U1048 ( .A(KEYINPUT61), .B(n951), .ZN(n953) );
  INV_X1 U1049 ( .A(G16), .ZN(n952) );
  NAND2_X1 U1050 ( .A1(n953), .A2(n952), .ZN(n954) );
  NAND2_X1 U1051 ( .A1(n954), .A2(G11), .ZN(n1005) );
  XNOR2_X1 U1052 ( .A(KEYINPUT121), .B(G2072), .ZN(n955) );
  XNOR2_X1 U1053 ( .A(n955), .B(G33), .ZN(n964) );
  XNOR2_X1 U1054 ( .A(G2067), .B(G26), .ZN(n957) );
  XNOR2_X1 U1055 ( .A(G1991), .B(G25), .ZN(n956) );
  NOR2_X1 U1056 ( .A1(n957), .A2(n956), .ZN(n958) );
  NAND2_X1 U1057 ( .A1(G28), .A2(n958), .ZN(n962) );
  XOR2_X1 U1058 ( .A(KEYINPUT122), .B(n959), .Z(n960) );
  XNOR2_X1 U1059 ( .A(G32), .B(n960), .ZN(n961) );
  NOR2_X1 U1060 ( .A1(n962), .A2(n961), .ZN(n963) );
  NAND2_X1 U1061 ( .A1(n964), .A2(n963), .ZN(n967) );
  XOR2_X1 U1062 ( .A(G27), .B(n965), .Z(n966) );
  NOR2_X1 U1063 ( .A1(n967), .A2(n966), .ZN(n968) );
  XOR2_X1 U1064 ( .A(KEYINPUT53), .B(n968), .Z(n972) );
  XNOR2_X1 U1065 ( .A(KEYINPUT54), .B(G34), .ZN(n969) );
  XNOR2_X1 U1066 ( .A(n969), .B(KEYINPUT123), .ZN(n970) );
  XNOR2_X1 U1067 ( .A(G2084), .B(n970), .ZN(n971) );
  NAND2_X1 U1068 ( .A1(n972), .A2(n971), .ZN(n974) );
  XNOR2_X1 U1069 ( .A(G35), .B(G2090), .ZN(n973) );
  NOR2_X1 U1070 ( .A1(n974), .A2(n973), .ZN(n975) );
  XNOR2_X1 U1071 ( .A(KEYINPUT124), .B(n975), .ZN(n976) );
  NOR2_X1 U1072 ( .A1(G29), .A2(n976), .ZN(n977) );
  XNOR2_X1 U1073 ( .A(n977), .B(KEYINPUT55), .ZN(n1003) );
  NOR2_X1 U1074 ( .A1(n979), .A2(n978), .ZN(n986) );
  XNOR2_X1 U1075 ( .A(G160), .B(G2084), .ZN(n981) );
  NAND2_X1 U1076 ( .A1(n981), .A2(n980), .ZN(n982) );
  NOR2_X1 U1077 ( .A1(n983), .A2(n982), .ZN(n984) );
  XNOR2_X1 U1078 ( .A(n984), .B(KEYINPUT120), .ZN(n985) );
  NAND2_X1 U1079 ( .A1(n986), .A2(n985), .ZN(n991) );
  XOR2_X1 U1080 ( .A(G2090), .B(G162), .Z(n987) );
  NOR2_X1 U1081 ( .A1(n988), .A2(n987), .ZN(n989) );
  XNOR2_X1 U1082 ( .A(n989), .B(KEYINPUT51), .ZN(n990) );
  NOR2_X1 U1083 ( .A1(n991), .A2(n990), .ZN(n999) );
  XOR2_X1 U1084 ( .A(G2072), .B(n992), .Z(n994) );
  XOR2_X1 U1085 ( .A(G164), .B(G2078), .Z(n993) );
  NOR2_X1 U1086 ( .A1(n994), .A2(n993), .ZN(n995) );
  XOR2_X1 U1087 ( .A(KEYINPUT50), .B(n995), .Z(n996) );
  NOR2_X1 U1088 ( .A1(n997), .A2(n996), .ZN(n998) );
  NAND2_X1 U1089 ( .A1(n999), .A2(n998), .ZN(n1000) );
  XNOR2_X1 U1090 ( .A(KEYINPUT52), .B(n1000), .ZN(n1001) );
  NAND2_X1 U1091 ( .A1(G29), .A2(n1001), .ZN(n1002) );
  NAND2_X1 U1092 ( .A1(n1003), .A2(n1002), .ZN(n1004) );
  NOR2_X1 U1093 ( .A1(n1005), .A2(n1004), .ZN(n1006) );
  NAND2_X1 U1094 ( .A1(n1007), .A2(n1006), .ZN(n1008) );
  XOR2_X1 U1095 ( .A(KEYINPUT62), .B(n1008), .Z(G311) );
  INV_X1 U1096 ( .A(G311), .ZN(G150) );
endmodule

