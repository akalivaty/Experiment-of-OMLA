//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 1 1 1 0 0 0 1 1 0 1 1 1 1 1 1 1 0 1 1 0 1 0 1 1 1 1 0 0 0 1 1 1 0 0 0 0 0 0 1 0 0 0 0 0 1 0 0 0 0 1 0 0 1 1 0 0 1 0 0 1 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:22:12 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n698, new_n699, new_n700, new_n701, new_n702, new_n703,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n716, new_n717, new_n719, new_n720,
    new_n721, new_n723, new_n724, new_n725, new_n726, new_n727, new_n728,
    new_n729, new_n730, new_n731, new_n733, new_n734, new_n735, new_n736,
    new_n737, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n762, new_n763, new_n764, new_n765, new_n766,
    new_n767, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n797, new_n798, new_n799, new_n800, new_n801, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n917,
    new_n918, new_n919, new_n920, new_n921, new_n922, new_n923, new_n924,
    new_n925, new_n926, new_n927, new_n928, new_n929, new_n930, new_n931,
    new_n932, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n948, new_n949, new_n950, new_n951, new_n953, new_n954, new_n955,
    new_n956, new_n957, new_n958, new_n959, new_n960, new_n961, new_n962,
    new_n963, new_n964, new_n965, new_n966, new_n967, new_n968, new_n970,
    new_n971, new_n972, new_n973, new_n974, new_n975, new_n976, new_n977,
    new_n978, new_n979, new_n980, new_n981, new_n982, new_n984, new_n985,
    new_n986, new_n987, new_n988, new_n989, new_n990, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1019,
    new_n1020, new_n1021, new_n1022, new_n1023, new_n1024, new_n1025,
    new_n1026, new_n1027, new_n1028, new_n1029;
  XNOR2_X1  g000(.A(G119), .B(G128), .ZN(new_n187));
  XNOR2_X1  g001(.A(new_n187), .B(KEYINPUT76), .ZN(new_n188));
  XOR2_X1   g002(.A(KEYINPUT24), .B(G110), .Z(new_n189));
  INV_X1    g003(.A(G128), .ZN(new_n190));
  INV_X1    g004(.A(KEYINPUT77), .ZN(new_n191));
  OAI211_X1 g005(.A(G119), .B(new_n190), .C1(new_n191), .C2(KEYINPUT23), .ZN(new_n192));
  INV_X1    g006(.A(KEYINPUT23), .ZN(new_n193));
  INV_X1    g007(.A(G119), .ZN(new_n194));
  AOI21_X1  g008(.A(new_n193), .B1(new_n194), .B2(G128), .ZN(new_n195));
  OAI21_X1  g009(.A(KEYINPUT77), .B1(new_n194), .B2(G128), .ZN(new_n196));
  OAI21_X1  g010(.A(new_n192), .B1(new_n195), .B2(new_n196), .ZN(new_n197));
  AOI22_X1  g011(.A1(new_n188), .A2(new_n189), .B1(G110), .B2(new_n197), .ZN(new_n198));
  INV_X1    g012(.A(KEYINPUT79), .ZN(new_n199));
  INV_X1    g013(.A(G125), .ZN(new_n200));
  AOI21_X1  g014(.A(new_n199), .B1(new_n200), .B2(G140), .ZN(new_n201));
  XNOR2_X1  g015(.A(KEYINPUT78), .B(G140), .ZN(new_n202));
  OAI21_X1  g016(.A(new_n201), .B1(new_n202), .B2(new_n200), .ZN(new_n203));
  INV_X1    g017(.A(G140), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n204), .A2(KEYINPUT78), .ZN(new_n205));
  INV_X1    g019(.A(KEYINPUT78), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n206), .A2(G140), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n205), .A2(new_n207), .ZN(new_n208));
  NAND3_X1  g022(.A1(new_n208), .A2(new_n199), .A3(G125), .ZN(new_n209));
  NAND3_X1  g023(.A1(new_n203), .A2(new_n209), .A3(KEYINPUT16), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n204), .A2(G125), .ZN(new_n211));
  INV_X1    g025(.A(KEYINPUT16), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n210), .A2(new_n213), .ZN(new_n214));
  NOR2_X1   g028(.A1(new_n214), .A2(G146), .ZN(new_n215));
  INV_X1    g029(.A(G146), .ZN(new_n216));
  AOI21_X1  g030(.A(new_n216), .B1(new_n210), .B2(new_n213), .ZN(new_n217));
  OAI21_X1  g031(.A(new_n198), .B1(new_n215), .B2(new_n217), .ZN(new_n218));
  INV_X1    g032(.A(new_n217), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n200), .A2(G140), .ZN(new_n220));
  NAND3_X1  g034(.A1(new_n211), .A2(new_n220), .A3(new_n216), .ZN(new_n221));
  XOR2_X1   g035(.A(new_n221), .B(KEYINPUT80), .Z(new_n222));
  INV_X1    g036(.A(new_n222), .ZN(new_n223));
  OAI22_X1  g037(.A1(new_n188), .A2(new_n189), .B1(G110), .B2(new_n197), .ZN(new_n224));
  NAND3_X1  g038(.A1(new_n219), .A2(new_n223), .A3(new_n224), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n218), .A2(new_n225), .ZN(new_n226));
  XNOR2_X1  g040(.A(KEYINPUT22), .B(G137), .ZN(new_n227));
  INV_X1    g041(.A(G221), .ZN(new_n228));
  INV_X1    g042(.A(G234), .ZN(new_n229));
  NOR3_X1   g043(.A1(new_n228), .A2(new_n229), .A3(G953), .ZN(new_n230));
  XOR2_X1   g044(.A(new_n227), .B(new_n230), .Z(new_n231));
  INV_X1    g045(.A(new_n231), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n226), .A2(new_n232), .ZN(new_n233));
  NAND3_X1  g047(.A1(new_n218), .A2(new_n225), .A3(new_n231), .ZN(new_n234));
  INV_X1    g048(.A(KEYINPUT81), .ZN(new_n235));
  INV_X1    g049(.A(KEYINPUT25), .ZN(new_n236));
  AOI21_X1  g050(.A(G902), .B1(new_n235), .B2(new_n236), .ZN(new_n237));
  NAND3_X1  g051(.A1(new_n233), .A2(new_n234), .A3(new_n237), .ZN(new_n238));
  NOR2_X1   g052(.A1(new_n235), .A2(new_n236), .ZN(new_n239));
  OR2_X1    g053(.A1(new_n238), .A2(new_n239), .ZN(new_n240));
  OAI21_X1  g054(.A(G217), .B1(new_n229), .B2(G902), .ZN(new_n241));
  AOI21_X1  g055(.A(new_n241), .B1(new_n238), .B2(new_n239), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n240), .A2(new_n242), .ZN(new_n243));
  AND2_X1   g057(.A1(new_n233), .A2(new_n234), .ZN(new_n244));
  AOI21_X1  g058(.A(G902), .B1(new_n229), .B2(G217), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n244), .A2(new_n245), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n243), .A2(new_n246), .ZN(new_n247));
  INV_X1    g061(.A(G472), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n216), .A2(G143), .ZN(new_n249));
  INV_X1    g063(.A(KEYINPUT64), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  NAND2_X1  g065(.A1(KEYINPUT0), .A2(G128), .ZN(new_n252));
  INV_X1    g066(.A(new_n252), .ZN(new_n253));
  NAND3_X1  g067(.A1(new_n216), .A2(KEYINPUT64), .A3(G143), .ZN(new_n254));
  INV_X1    g068(.A(G143), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n255), .A2(G146), .ZN(new_n256));
  NAND4_X1  g070(.A1(new_n251), .A2(new_n253), .A3(new_n254), .A4(new_n256), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n249), .A2(new_n256), .ZN(new_n258));
  OR2_X1    g072(.A1(KEYINPUT0), .A2(G128), .ZN(new_n259));
  NAND3_X1  g073(.A1(new_n258), .A2(new_n252), .A3(new_n259), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n257), .A2(new_n260), .ZN(new_n261));
  INV_X1    g075(.A(new_n261), .ZN(new_n262));
  INV_X1    g076(.A(KEYINPUT11), .ZN(new_n263));
  INV_X1    g077(.A(G134), .ZN(new_n264));
  OAI21_X1  g078(.A(new_n263), .B1(new_n264), .B2(G137), .ZN(new_n265));
  INV_X1    g079(.A(G137), .ZN(new_n266));
  NAND3_X1  g080(.A1(new_n266), .A2(KEYINPUT11), .A3(G134), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n264), .A2(G137), .ZN(new_n268));
  NAND3_X1  g082(.A1(new_n265), .A2(new_n267), .A3(new_n268), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n269), .A2(G131), .ZN(new_n270));
  INV_X1    g084(.A(G131), .ZN(new_n271));
  NAND4_X1  g085(.A1(new_n265), .A2(new_n267), .A3(new_n271), .A4(new_n268), .ZN(new_n272));
  AND3_X1   g086(.A1(new_n270), .A2(KEYINPUT69), .A3(new_n272), .ZN(new_n273));
  AOI21_X1  g087(.A(KEYINPUT69), .B1(new_n270), .B2(new_n272), .ZN(new_n274));
  OAI21_X1  g088(.A(new_n262), .B1(new_n273), .B2(new_n274), .ZN(new_n275));
  NOR2_X1   g089(.A1(new_n190), .A2(KEYINPUT1), .ZN(new_n276));
  NAND4_X1  g090(.A1(new_n251), .A2(new_n254), .A3(new_n256), .A4(new_n276), .ZN(new_n277));
  AOI21_X1  g091(.A(new_n190), .B1(new_n249), .B2(KEYINPUT1), .ZN(new_n278));
  XNOR2_X1  g092(.A(G143), .B(G146), .ZN(new_n279));
  NOR3_X1   g093(.A1(new_n278), .A2(new_n279), .A3(KEYINPUT66), .ZN(new_n280));
  INV_X1    g094(.A(KEYINPUT66), .ZN(new_n281));
  OAI21_X1  g095(.A(KEYINPUT1), .B1(new_n255), .B2(G146), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n282), .A2(G128), .ZN(new_n283));
  AOI21_X1  g097(.A(new_n281), .B1(new_n283), .B2(new_n258), .ZN(new_n284));
  OAI21_X1  g098(.A(new_n277), .B1(new_n280), .B2(new_n284), .ZN(new_n285));
  XNOR2_X1  g099(.A(G134), .B(G137), .ZN(new_n286));
  OAI21_X1  g100(.A(KEYINPUT65), .B1(new_n286), .B2(new_n271), .ZN(new_n287));
  INV_X1    g101(.A(KEYINPUT65), .ZN(new_n288));
  NOR2_X1   g102(.A1(new_n264), .A2(G137), .ZN(new_n289));
  NOR2_X1   g103(.A1(new_n266), .A2(G134), .ZN(new_n290));
  OAI211_X1 g104(.A(new_n288), .B(G131), .C1(new_n289), .C2(new_n290), .ZN(new_n291));
  NAND3_X1  g105(.A1(new_n287), .A2(new_n272), .A3(new_n291), .ZN(new_n292));
  INV_X1    g106(.A(new_n292), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n285), .A2(new_n293), .ZN(new_n294));
  INV_X1    g108(.A(KEYINPUT67), .ZN(new_n295));
  INV_X1    g109(.A(G116), .ZN(new_n296));
  OAI21_X1  g110(.A(new_n295), .B1(new_n296), .B2(G119), .ZN(new_n297));
  NAND3_X1  g111(.A1(new_n194), .A2(KEYINPUT67), .A3(G116), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n296), .A2(G119), .ZN(new_n299));
  NAND3_X1  g113(.A1(new_n297), .A2(new_n298), .A3(new_n299), .ZN(new_n300));
  INV_X1    g114(.A(G113), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n301), .A2(KEYINPUT2), .ZN(new_n302));
  INV_X1    g116(.A(KEYINPUT2), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n303), .A2(G113), .ZN(new_n304));
  AND2_X1   g118(.A1(new_n302), .A2(new_n304), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n300), .A2(new_n305), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n302), .A2(new_n304), .ZN(new_n307));
  NAND4_X1  g121(.A1(new_n307), .A2(new_n297), .A3(new_n298), .A4(new_n299), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n306), .A2(new_n308), .ZN(new_n309));
  INV_X1    g123(.A(KEYINPUT68), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  NAND3_X1  g125(.A1(new_n306), .A2(new_n308), .A3(KEYINPUT68), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  NAND3_X1  g127(.A1(new_n275), .A2(new_n294), .A3(new_n313), .ZN(new_n314));
  INV_X1    g128(.A(new_n314), .ZN(new_n315));
  AOI21_X1  g129(.A(new_n313), .B1(new_n275), .B2(new_n294), .ZN(new_n316));
  OAI21_X1  g130(.A(KEYINPUT28), .B1(new_n315), .B2(new_n316), .ZN(new_n317));
  INV_X1    g131(.A(KEYINPUT28), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n314), .A2(new_n318), .ZN(new_n319));
  NOR2_X1   g133(.A1(G237), .A2(G953), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n320), .A2(G210), .ZN(new_n321));
  XNOR2_X1  g135(.A(new_n321), .B(KEYINPUT27), .ZN(new_n322));
  XNOR2_X1  g136(.A(KEYINPUT26), .B(G101), .ZN(new_n323));
  XNOR2_X1  g137(.A(new_n322), .B(new_n323), .ZN(new_n324));
  INV_X1    g138(.A(new_n324), .ZN(new_n325));
  INV_X1    g139(.A(KEYINPUT29), .ZN(new_n326));
  NOR2_X1   g140(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  NAND3_X1  g141(.A1(new_n317), .A2(new_n319), .A3(new_n327), .ZN(new_n328));
  INV_X1    g142(.A(G902), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n328), .A2(new_n329), .ZN(new_n330));
  AND3_X1   g144(.A1(new_n306), .A2(new_n308), .A3(KEYINPUT68), .ZN(new_n331));
  AOI21_X1  g145(.A(KEYINPUT68), .B1(new_n306), .B2(new_n308), .ZN(new_n332));
  NOR2_X1   g146(.A1(new_n331), .A2(new_n332), .ZN(new_n333));
  OAI21_X1  g147(.A(KEYINPUT66), .B1(new_n278), .B2(new_n279), .ZN(new_n334));
  NAND3_X1  g148(.A1(new_n283), .A2(new_n281), .A3(new_n258), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  AOI21_X1  g150(.A(new_n292), .B1(new_n336), .B2(new_n277), .ZN(new_n337));
  AOI21_X1  g151(.A(new_n261), .B1(new_n272), .B2(new_n270), .ZN(new_n338));
  OAI21_X1  g152(.A(new_n333), .B1(new_n337), .B2(new_n338), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n314), .A2(new_n339), .ZN(new_n340));
  XOR2_X1   g154(.A(KEYINPUT71), .B(KEYINPUT28), .Z(new_n341));
  NAND2_X1  g155(.A1(new_n340), .A2(new_n341), .ZN(new_n342));
  XNOR2_X1  g156(.A(new_n324), .B(KEYINPUT70), .ZN(new_n343));
  INV_X1    g157(.A(new_n343), .ZN(new_n344));
  NAND3_X1  g158(.A1(new_n342), .A2(new_n344), .A3(new_n319), .ZN(new_n345));
  NAND3_X1  g159(.A1(new_n275), .A2(KEYINPUT30), .A3(new_n294), .ZN(new_n346));
  INV_X1    g160(.A(KEYINPUT30), .ZN(new_n347));
  OAI21_X1  g161(.A(new_n347), .B1(new_n337), .B2(new_n338), .ZN(new_n348));
  NAND3_X1  g162(.A1(new_n346), .A2(new_n333), .A3(new_n348), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n349), .A2(new_n314), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n350), .A2(new_n325), .ZN(new_n351));
  NAND3_X1  g165(.A1(new_n345), .A2(new_n351), .A3(new_n326), .ZN(new_n352));
  INV_X1    g166(.A(KEYINPUT75), .ZN(new_n353));
  AOI21_X1  g167(.A(new_n330), .B1(new_n352), .B2(new_n353), .ZN(new_n354));
  NAND4_X1  g168(.A1(new_n345), .A2(new_n351), .A3(KEYINPUT75), .A4(new_n326), .ZN(new_n355));
  AOI21_X1  g169(.A(new_n248), .B1(new_n354), .B2(new_n355), .ZN(new_n356));
  NAND3_X1  g170(.A1(new_n349), .A2(new_n314), .A3(new_n324), .ZN(new_n357));
  INV_X1    g171(.A(KEYINPUT31), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n357), .A2(new_n358), .ZN(new_n359));
  NAND4_X1  g173(.A1(new_n349), .A2(KEYINPUT31), .A3(new_n314), .A4(new_n324), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n359), .A2(new_n360), .ZN(new_n361));
  INV_X1    g175(.A(KEYINPUT72), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n342), .A2(new_n319), .ZN(new_n363));
  AOI21_X1  g177(.A(new_n362), .B1(new_n363), .B2(new_n343), .ZN(new_n364));
  INV_X1    g178(.A(new_n341), .ZN(new_n365));
  AOI21_X1  g179(.A(new_n365), .B1(new_n314), .B2(new_n339), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n270), .A2(new_n272), .ZN(new_n367));
  INV_X1    g181(.A(KEYINPUT69), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  NAND3_X1  g183(.A1(new_n270), .A2(KEYINPUT69), .A3(new_n272), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n369), .A2(new_n370), .ZN(new_n371));
  AOI21_X1  g185(.A(new_n337), .B1(new_n371), .B2(new_n262), .ZN(new_n372));
  AOI21_X1  g186(.A(KEYINPUT28), .B1(new_n372), .B2(new_n313), .ZN(new_n373));
  OAI211_X1 g187(.A(new_n362), .B(new_n343), .C1(new_n366), .C2(new_n373), .ZN(new_n374));
  INV_X1    g188(.A(new_n374), .ZN(new_n375));
  OAI21_X1  g189(.A(new_n361), .B1(new_n364), .B2(new_n375), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n376), .A2(KEYINPUT73), .ZN(new_n377));
  AOI22_X1  g191(.A1(new_n340), .A2(new_n341), .B1(new_n318), .B2(new_n314), .ZN(new_n378));
  OAI21_X1  g192(.A(KEYINPUT72), .B1(new_n378), .B2(new_n344), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n379), .A2(new_n374), .ZN(new_n380));
  INV_X1    g194(.A(KEYINPUT73), .ZN(new_n381));
  NAND3_X1  g195(.A1(new_n380), .A2(new_n381), .A3(new_n361), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n377), .A2(new_n382), .ZN(new_n383));
  NOR2_X1   g197(.A1(G472), .A2(G902), .ZN(new_n384));
  AND2_X1   g198(.A1(new_n384), .A2(KEYINPUT32), .ZN(new_n385));
  AOI21_X1  g199(.A(new_n356), .B1(new_n383), .B2(new_n385), .ZN(new_n386));
  AOI221_X4 g200(.A(KEYINPUT73), .B1(new_n359), .B2(new_n360), .C1(new_n379), .C2(new_n374), .ZN(new_n387));
  AOI21_X1  g201(.A(new_n381), .B1(new_n380), .B2(new_n361), .ZN(new_n388));
  OAI21_X1  g202(.A(new_n384), .B1(new_n387), .B2(new_n388), .ZN(new_n389));
  XOR2_X1   g203(.A(KEYINPUT74), .B(KEYINPUT32), .Z(new_n390));
  INV_X1    g204(.A(new_n390), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n389), .A2(new_n391), .ZN(new_n392));
  AOI21_X1  g206(.A(new_n247), .B1(new_n386), .B2(new_n392), .ZN(new_n393));
  INV_X1    g207(.A(KEYINPUT92), .ZN(new_n394));
  XNOR2_X1  g208(.A(KEYINPUT9), .B(G234), .ZN(new_n395));
  INV_X1    g209(.A(new_n395), .ZN(new_n396));
  AOI21_X1  g210(.A(new_n228), .B1(new_n396), .B2(new_n329), .ZN(new_n397));
  INV_X1    g211(.A(G469), .ZN(new_n398));
  NOR2_X1   g212(.A1(new_n398), .A2(new_n329), .ZN(new_n399));
  INV_X1    g213(.A(KEYINPUT10), .ZN(new_n400));
  NAND3_X1  g214(.A1(new_n251), .A2(new_n254), .A3(new_n256), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n401), .A2(new_n283), .ZN(new_n402));
  AND2_X1   g216(.A1(new_n402), .A2(new_n277), .ZN(new_n403));
  INV_X1    g217(.A(G104), .ZN(new_n404));
  NOR2_X1   g218(.A1(new_n404), .A2(G107), .ZN(new_n405));
  INV_X1    g219(.A(G107), .ZN(new_n406));
  NOR2_X1   g220(.A1(new_n406), .A2(G104), .ZN(new_n407));
  OAI21_X1  g221(.A(G101), .B1(new_n405), .B2(new_n407), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n408), .A2(KEYINPUT82), .ZN(new_n409));
  OAI21_X1  g223(.A(KEYINPUT3), .B1(new_n404), .B2(G107), .ZN(new_n410));
  INV_X1    g224(.A(KEYINPUT3), .ZN(new_n411));
  NAND3_X1  g225(.A1(new_n411), .A2(new_n406), .A3(G104), .ZN(new_n412));
  INV_X1    g226(.A(G101), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n404), .A2(G107), .ZN(new_n414));
  NAND4_X1  g228(.A1(new_n410), .A2(new_n412), .A3(new_n413), .A4(new_n414), .ZN(new_n415));
  INV_X1    g229(.A(KEYINPUT82), .ZN(new_n416));
  OAI211_X1 g230(.A(new_n416), .B(G101), .C1(new_n405), .C2(new_n407), .ZN(new_n417));
  NAND3_X1  g231(.A1(new_n409), .A2(new_n415), .A3(new_n417), .ZN(new_n418));
  OAI21_X1  g232(.A(new_n400), .B1(new_n403), .B2(new_n418), .ZN(new_n419));
  AND3_X1   g233(.A1(new_n409), .A2(new_n415), .A3(new_n417), .ZN(new_n420));
  NAND3_X1  g234(.A1(new_n420), .A2(new_n285), .A3(KEYINPUT10), .ZN(new_n421));
  NAND3_X1  g235(.A1(new_n410), .A2(new_n412), .A3(new_n414), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n422), .A2(G101), .ZN(new_n423));
  NAND3_X1  g237(.A1(new_n423), .A2(KEYINPUT4), .A3(new_n415), .ZN(new_n424));
  INV_X1    g238(.A(KEYINPUT4), .ZN(new_n425));
  NAND3_X1  g239(.A1(new_n422), .A2(new_n425), .A3(G101), .ZN(new_n426));
  NAND3_X1  g240(.A1(new_n262), .A2(new_n424), .A3(new_n426), .ZN(new_n427));
  NAND3_X1  g241(.A1(new_n419), .A2(new_n421), .A3(new_n427), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n428), .A2(new_n371), .ZN(new_n429));
  INV_X1    g243(.A(new_n371), .ZN(new_n430));
  NAND4_X1  g244(.A1(new_n430), .A2(new_n419), .A3(new_n427), .A4(new_n421), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n429), .A2(new_n431), .ZN(new_n432));
  XNOR2_X1  g246(.A(G110), .B(G140), .ZN(new_n433));
  INV_X1    g247(.A(G953), .ZN(new_n434));
  AND2_X1   g248(.A1(new_n434), .A2(G227), .ZN(new_n435));
  XNOR2_X1  g249(.A(new_n433), .B(new_n435), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n432), .A2(new_n436), .ZN(new_n437));
  INV_X1    g251(.A(new_n436), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n402), .A2(new_n277), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n420), .A2(new_n439), .ZN(new_n440));
  NAND3_X1  g254(.A1(new_n418), .A2(new_n277), .A3(new_n336), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n440), .A2(new_n441), .ZN(new_n442));
  AOI21_X1  g256(.A(KEYINPUT12), .B1(new_n442), .B2(new_n371), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n367), .A2(KEYINPUT12), .ZN(new_n444));
  AOI21_X1  g258(.A(new_n444), .B1(new_n440), .B2(new_n441), .ZN(new_n445));
  OAI211_X1 g259(.A(new_n431), .B(new_n438), .C1(new_n443), .C2(new_n445), .ZN(new_n446));
  AOI21_X1  g260(.A(G902), .B1(new_n437), .B2(new_n446), .ZN(new_n447));
  AOI21_X1  g261(.A(new_n399), .B1(new_n447), .B2(new_n398), .ZN(new_n448));
  NOR2_X1   g262(.A1(new_n443), .A2(new_n445), .ZN(new_n449));
  INV_X1    g263(.A(new_n431), .ZN(new_n450));
  OAI21_X1  g264(.A(new_n436), .B1(new_n449), .B2(new_n450), .ZN(new_n451));
  NAND3_X1  g265(.A1(new_n429), .A2(new_n431), .A3(new_n438), .ZN(new_n452));
  NAND3_X1  g266(.A1(new_n451), .A2(G469), .A3(new_n452), .ZN(new_n453));
  AOI21_X1  g267(.A(new_n397), .B1(new_n448), .B2(new_n453), .ZN(new_n454));
  OAI21_X1  g268(.A(G214), .B1(G237), .B2(G902), .ZN(new_n455));
  INV_X1    g269(.A(new_n455), .ZN(new_n456));
  OAI21_X1  g270(.A(G210), .B1(G237), .B2(G902), .ZN(new_n457));
  NOR2_X1   g271(.A1(new_n296), .A2(G119), .ZN(new_n458));
  INV_X1    g272(.A(KEYINPUT5), .ZN(new_n459));
  AOI21_X1  g273(.A(new_n301), .B1(new_n458), .B2(new_n459), .ZN(new_n460));
  OAI21_X1  g274(.A(new_n460), .B1(new_n300), .B2(new_n459), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n461), .A2(new_n308), .ZN(new_n462));
  NOR2_X1   g276(.A1(new_n462), .A2(new_n418), .ZN(new_n463));
  AND2_X1   g277(.A1(new_n424), .A2(new_n426), .ZN(new_n464));
  AOI21_X1  g278(.A(new_n463), .B1(new_n333), .B2(new_n464), .ZN(new_n465));
  XNOR2_X1  g279(.A(G110), .B(G122), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n424), .A2(new_n426), .ZN(new_n468));
  OAI22_X1  g282(.A1(new_n313), .A2(new_n468), .B1(new_n418), .B2(new_n462), .ZN(new_n469));
  INV_X1    g283(.A(new_n466), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  NAND3_X1  g285(.A1(new_n467), .A2(new_n471), .A3(KEYINPUT6), .ZN(new_n472));
  OR3_X1    g286(.A1(new_n465), .A2(KEYINPUT6), .A3(new_n466), .ZN(new_n473));
  INV_X1    g287(.A(KEYINPUT83), .ZN(new_n474));
  OAI21_X1  g288(.A(new_n474), .B1(new_n262), .B2(new_n200), .ZN(new_n475));
  NAND3_X1  g289(.A1(new_n261), .A2(KEYINPUT83), .A3(G125), .ZN(new_n476));
  NAND3_X1  g290(.A1(new_n336), .A2(new_n200), .A3(new_n277), .ZN(new_n477));
  NAND3_X1  g291(.A1(new_n475), .A2(new_n476), .A3(new_n477), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n434), .A2(G224), .ZN(new_n479));
  XNOR2_X1  g293(.A(new_n479), .B(KEYINPUT84), .ZN(new_n480));
  INV_X1    g294(.A(new_n480), .ZN(new_n481));
  XNOR2_X1  g295(.A(new_n478), .B(new_n481), .ZN(new_n482));
  NAND3_X1  g296(.A1(new_n472), .A2(new_n473), .A3(new_n482), .ZN(new_n483));
  AND3_X1   g297(.A1(new_n475), .A2(new_n476), .A3(new_n477), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n480), .A2(KEYINPUT7), .ZN(new_n485));
  INV_X1    g299(.A(new_n485), .ZN(new_n486));
  AOI22_X1  g300(.A1(new_n484), .A2(new_n486), .B1(new_n465), .B2(new_n466), .ZN(new_n487));
  XNOR2_X1  g301(.A(new_n462), .B(new_n418), .ZN(new_n488));
  XNOR2_X1  g302(.A(new_n466), .B(KEYINPUT8), .ZN(new_n489));
  AOI22_X1  g303(.A1(new_n478), .A2(new_n485), .B1(new_n488), .B2(new_n489), .ZN(new_n490));
  AOI21_X1  g304(.A(G902), .B1(new_n487), .B2(new_n490), .ZN(new_n491));
  AOI21_X1  g305(.A(new_n457), .B1(new_n483), .B2(new_n491), .ZN(new_n492));
  INV_X1    g306(.A(new_n492), .ZN(new_n493));
  NAND3_X1  g307(.A1(new_n483), .A2(new_n491), .A3(new_n457), .ZN(new_n494));
  AOI21_X1  g308(.A(new_n456), .B1(new_n493), .B2(new_n494), .ZN(new_n495));
  OR2_X1    g309(.A1(KEYINPUT91), .A2(G952), .ZN(new_n496));
  NAND2_X1  g310(.A1(KEYINPUT91), .A2(G952), .ZN(new_n497));
  AOI21_X1  g311(.A(G953), .B1(new_n496), .B2(new_n497), .ZN(new_n498));
  INV_X1    g312(.A(G237), .ZN(new_n499));
  OAI21_X1  g313(.A(new_n498), .B1(new_n229), .B2(new_n499), .ZN(new_n500));
  INV_X1    g314(.A(new_n500), .ZN(new_n501));
  XNOR2_X1  g315(.A(KEYINPUT21), .B(G898), .ZN(new_n502));
  AOI211_X1 g316(.A(new_n329), .B(new_n434), .C1(G234), .C2(G237), .ZN(new_n503));
  AOI21_X1  g317(.A(new_n501), .B1(new_n502), .B2(new_n503), .ZN(new_n504));
  INV_X1    g318(.A(new_n504), .ZN(new_n505));
  NAND3_X1  g319(.A1(new_n454), .A2(new_n495), .A3(new_n505), .ZN(new_n506));
  INV_X1    g320(.A(KEYINPUT20), .ZN(new_n507));
  NOR2_X1   g321(.A1(G475), .A2(G902), .ZN(new_n508));
  XNOR2_X1  g322(.A(G113), .B(G122), .ZN(new_n509));
  XNOR2_X1  g323(.A(new_n509), .B(new_n404), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n320), .A2(G214), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n511), .A2(new_n255), .ZN(new_n512));
  NAND3_X1  g326(.A1(new_n320), .A2(G143), .A3(G214), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  NAND2_X1  g328(.A1(KEYINPUT18), .A2(G131), .ZN(new_n515));
  INV_X1    g329(.A(new_n515), .ZN(new_n516));
  XNOR2_X1  g330(.A(new_n514), .B(new_n516), .ZN(new_n517));
  INV_X1    g331(.A(new_n517), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n220), .A2(KEYINPUT79), .ZN(new_n519));
  AOI21_X1  g333(.A(new_n519), .B1(new_n208), .B2(G125), .ZN(new_n520));
  AOI211_X1 g334(.A(KEYINPUT79), .B(new_n200), .C1(new_n205), .C2(new_n207), .ZN(new_n521));
  OAI21_X1  g335(.A(KEYINPUT85), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  INV_X1    g336(.A(KEYINPUT85), .ZN(new_n523));
  NAND3_X1  g337(.A1(new_n203), .A2(new_n209), .A3(new_n523), .ZN(new_n524));
  AOI21_X1  g338(.A(new_n216), .B1(new_n522), .B2(new_n524), .ZN(new_n525));
  NOR3_X1   g339(.A1(new_n525), .A2(KEYINPUT86), .A3(new_n222), .ZN(new_n526));
  INV_X1    g340(.A(KEYINPUT86), .ZN(new_n527));
  AND3_X1   g341(.A1(new_n203), .A2(new_n209), .A3(new_n523), .ZN(new_n528));
  AOI21_X1  g342(.A(new_n523), .B1(new_n203), .B2(new_n209), .ZN(new_n529));
  OAI21_X1  g343(.A(G146), .B1(new_n528), .B2(new_n529), .ZN(new_n530));
  AOI21_X1  g344(.A(new_n527), .B1(new_n530), .B2(new_n223), .ZN(new_n531));
  OAI21_X1  g345(.A(new_n518), .B1(new_n526), .B2(new_n531), .ZN(new_n532));
  INV_X1    g346(.A(KEYINPUT19), .ZN(new_n533));
  NAND3_X1  g347(.A1(new_n211), .A2(new_n220), .A3(new_n533), .ZN(new_n534));
  INV_X1    g348(.A(new_n534), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n522), .A2(new_n524), .ZN(new_n536));
  AOI21_X1  g350(.A(new_n535), .B1(new_n536), .B2(KEYINPUT19), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n537), .A2(new_n216), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n514), .A2(G131), .ZN(new_n539));
  NAND3_X1  g353(.A1(new_n512), .A2(new_n271), .A3(new_n513), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  NAND3_X1  g355(.A1(new_n538), .A2(new_n219), .A3(new_n541), .ZN(new_n542));
  AOI21_X1  g356(.A(new_n510), .B1(new_n532), .B2(new_n542), .ZN(new_n543));
  OAI21_X1  g357(.A(KEYINPUT86), .B1(new_n525), .B2(new_n222), .ZN(new_n544));
  NAND3_X1  g358(.A1(new_n530), .A2(new_n527), .A3(new_n223), .ZN(new_n545));
  AOI21_X1  g359(.A(new_n517), .B1(new_n544), .B2(new_n545), .ZN(new_n546));
  INV_X1    g360(.A(new_n510), .ZN(new_n547));
  NAND3_X1  g361(.A1(new_n514), .A2(KEYINPUT17), .A3(G131), .ZN(new_n548));
  OAI21_X1  g362(.A(new_n548), .B1(new_n541), .B2(KEYINPUT17), .ZN(new_n549));
  NOR3_X1   g363(.A1(new_n549), .A2(new_n215), .A3(new_n217), .ZN(new_n550));
  NOR3_X1   g364(.A1(new_n546), .A2(new_n547), .A3(new_n550), .ZN(new_n551));
  OAI211_X1 g365(.A(new_n507), .B(new_n508), .C1(new_n543), .C2(new_n551), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n552), .A2(KEYINPUT87), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n219), .A2(new_n541), .ZN(new_n554));
  AOI21_X1  g368(.A(new_n554), .B1(new_n216), .B2(new_n537), .ZN(new_n555));
  OAI21_X1  g369(.A(new_n547), .B1(new_n555), .B2(new_n546), .ZN(new_n556));
  INV_X1    g370(.A(new_n550), .ZN(new_n557));
  NAND3_X1  g371(.A1(new_n532), .A2(new_n557), .A3(new_n510), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n556), .A2(new_n558), .ZN(new_n559));
  INV_X1    g373(.A(KEYINPUT87), .ZN(new_n560));
  NAND4_X1  g374(.A1(new_n559), .A2(new_n560), .A3(new_n507), .A4(new_n508), .ZN(new_n561));
  OAI21_X1  g375(.A(new_n508), .B1(new_n543), .B2(new_n551), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n562), .A2(KEYINPUT20), .ZN(new_n563));
  NAND3_X1  g377(.A1(new_n553), .A2(new_n561), .A3(new_n563), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n255), .A2(G128), .ZN(new_n565));
  INV_X1    g379(.A(KEYINPUT13), .ZN(new_n566));
  XNOR2_X1  g380(.A(new_n565), .B(new_n566), .ZN(new_n567));
  OAI21_X1  g381(.A(KEYINPUT88), .B1(new_n255), .B2(G128), .ZN(new_n568));
  INV_X1    g382(.A(KEYINPUT88), .ZN(new_n569));
  NAND3_X1  g383(.A1(new_n569), .A2(new_n190), .A3(G143), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n568), .A2(new_n570), .ZN(new_n571));
  INV_X1    g385(.A(new_n571), .ZN(new_n572));
  OAI21_X1  g386(.A(G134), .B1(new_n567), .B2(new_n572), .ZN(new_n573));
  INV_X1    g387(.A(G122), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n574), .A2(G116), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n296), .A2(G122), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  XNOR2_X1  g391(.A(new_n577), .B(G107), .ZN(new_n578));
  AND2_X1   g392(.A1(new_n573), .A2(new_n578), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n571), .A2(new_n565), .ZN(new_n580));
  INV_X1    g394(.A(KEYINPUT89), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  NAND3_X1  g396(.A1(new_n571), .A2(KEYINPUT89), .A3(new_n565), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n584), .A2(new_n264), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n579), .A2(new_n585), .ZN(new_n586));
  INV_X1    g400(.A(new_n586), .ZN(new_n587));
  AOI21_X1  g401(.A(new_n406), .B1(new_n575), .B2(KEYINPUT14), .ZN(new_n588));
  XOR2_X1   g402(.A(new_n588), .B(new_n577), .Z(new_n589));
  INV_X1    g403(.A(new_n589), .ZN(new_n590));
  NAND3_X1  g404(.A1(new_n582), .A2(G134), .A3(new_n583), .ZN(new_n591));
  AOI21_X1  g405(.A(new_n590), .B1(new_n585), .B2(new_n591), .ZN(new_n592));
  NOR2_X1   g406(.A1(new_n587), .A2(new_n592), .ZN(new_n593));
  NAND3_X1  g407(.A1(new_n396), .A2(G217), .A3(new_n434), .ZN(new_n594));
  INV_X1    g408(.A(new_n594), .ZN(new_n595));
  AOI21_X1  g409(.A(KEYINPUT90), .B1(new_n593), .B2(new_n595), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n585), .A2(new_n591), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n597), .A2(new_n589), .ZN(new_n598));
  NAND4_X1  g412(.A1(new_n598), .A2(KEYINPUT90), .A3(new_n586), .A4(new_n595), .ZN(new_n599));
  OAI21_X1  g413(.A(new_n594), .B1(new_n587), .B2(new_n592), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  OAI21_X1  g415(.A(new_n329), .B1(new_n596), .B2(new_n601), .ZN(new_n602));
  INV_X1    g416(.A(G478), .ZN(new_n603));
  NOR2_X1   g417(.A1(new_n603), .A2(KEYINPUT15), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n602), .A2(new_n604), .ZN(new_n605));
  NAND3_X1  g419(.A1(new_n598), .A2(new_n586), .A3(new_n595), .ZN(new_n606));
  INV_X1    g420(.A(KEYINPUT90), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  NAND3_X1  g422(.A1(new_n608), .A2(new_n600), .A3(new_n599), .ZN(new_n609));
  OAI211_X1 g423(.A(new_n609), .B(new_n329), .C1(KEYINPUT15), .C2(new_n603), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n605), .A2(new_n610), .ZN(new_n611));
  INV_X1    g425(.A(new_n611), .ZN(new_n612));
  OAI21_X1  g426(.A(new_n547), .B1(new_n546), .B2(new_n550), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n558), .A2(new_n613), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n614), .A2(new_n329), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n615), .A2(G475), .ZN(new_n616));
  NAND3_X1  g430(.A1(new_n564), .A2(new_n612), .A3(new_n616), .ZN(new_n617));
  OAI21_X1  g431(.A(new_n394), .B1(new_n506), .B2(new_n617), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n564), .A2(new_n616), .ZN(new_n619));
  INV_X1    g433(.A(new_n619), .ZN(new_n620));
  INV_X1    g434(.A(new_n494), .ZN(new_n621));
  OAI211_X1 g435(.A(new_n505), .B(new_n455), .C1(new_n621), .C2(new_n492), .ZN(new_n622));
  INV_X1    g436(.A(new_n446), .ZN(new_n623));
  AOI21_X1  g437(.A(new_n438), .B1(new_n429), .B2(new_n431), .ZN(new_n624));
  OAI211_X1 g438(.A(new_n398), .B(new_n329), .C1(new_n623), .C2(new_n624), .ZN(new_n625));
  INV_X1    g439(.A(new_n399), .ZN(new_n626));
  NAND3_X1  g440(.A1(new_n625), .A2(new_n453), .A3(new_n626), .ZN(new_n627));
  INV_X1    g441(.A(new_n397), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  NOR2_X1   g443(.A1(new_n622), .A2(new_n629), .ZN(new_n630));
  NAND4_X1  g444(.A1(new_n620), .A2(KEYINPUT92), .A3(new_n630), .A4(new_n612), .ZN(new_n631));
  NAND3_X1  g445(.A1(new_n393), .A2(new_n618), .A3(new_n631), .ZN(new_n632));
  XNOR2_X1  g446(.A(new_n632), .B(G101), .ZN(G3));
  INV_X1    g447(.A(new_n384), .ZN(new_n634));
  AOI21_X1  g448(.A(new_n634), .B1(new_n377), .B2(new_n382), .ZN(new_n635));
  OAI21_X1  g449(.A(new_n329), .B1(new_n387), .B2(new_n388), .ZN(new_n636));
  AOI21_X1  g450(.A(new_n635), .B1(G472), .B2(new_n636), .ZN(new_n637));
  AND3_X1   g451(.A1(new_n600), .A2(new_n606), .A3(KEYINPUT33), .ZN(new_n638));
  INV_X1    g452(.A(KEYINPUT33), .ZN(new_n639));
  AOI21_X1  g453(.A(new_n638), .B1(new_n609), .B2(new_n639), .ZN(new_n640));
  NOR2_X1   g454(.A1(new_n603), .A2(G902), .ZN(new_n641));
  XNOR2_X1  g455(.A(KEYINPUT93), .B(G478), .ZN(new_n642));
  AOI22_X1  g456(.A1(new_n640), .A2(new_n641), .B1(new_n602), .B2(new_n642), .ZN(new_n643));
  AOI21_X1  g457(.A(new_n643), .B1(new_n564), .B2(new_n616), .ZN(new_n644));
  NOR3_X1   g458(.A1(new_n622), .A2(new_n629), .A3(new_n247), .ZN(new_n645));
  NAND3_X1  g459(.A1(new_n637), .A2(new_n644), .A3(new_n645), .ZN(new_n646));
  XOR2_X1   g460(.A(KEYINPUT34), .B(G104), .Z(new_n647));
  XNOR2_X1  g461(.A(new_n646), .B(new_n647), .ZN(G6));
  INV_X1    g462(.A(KEYINPUT94), .ZN(new_n649));
  NAND3_X1  g463(.A1(new_n615), .A2(new_n649), .A3(G475), .ZN(new_n650));
  AOI21_X1  g464(.A(G902), .B1(new_n558), .B2(new_n613), .ZN(new_n651));
  INV_X1    g465(.A(G475), .ZN(new_n652));
  OAI21_X1  g466(.A(KEYINPUT94), .B1(new_n651), .B2(new_n652), .ZN(new_n653));
  NAND2_X1  g467(.A1(new_n650), .A2(new_n653), .ZN(new_n654));
  INV_X1    g468(.A(new_n654), .ZN(new_n655));
  AOI22_X1  g469(.A1(new_n563), .A2(new_n552), .B1(new_n605), .B2(new_n610), .ZN(new_n656));
  AND4_X1   g470(.A1(new_n637), .A2(new_n645), .A3(new_n655), .A4(new_n656), .ZN(new_n657));
  XNOR2_X1  g471(.A(KEYINPUT35), .B(G107), .ZN(new_n658));
  XNOR2_X1  g472(.A(new_n657), .B(new_n658), .ZN(G9));
  NOR2_X1   g473(.A1(new_n232), .A2(KEYINPUT36), .ZN(new_n660));
  XNOR2_X1  g474(.A(new_n226), .B(new_n660), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n661), .A2(new_n245), .ZN(new_n662));
  NAND2_X1  g476(.A1(new_n243), .A2(new_n662), .ZN(new_n663));
  NAND4_X1  g477(.A1(new_n631), .A2(new_n618), .A3(new_n637), .A4(new_n663), .ZN(new_n664));
  XOR2_X1   g478(.A(KEYINPUT37), .B(G110), .Z(new_n665));
  XNOR2_X1  g479(.A(new_n665), .B(KEYINPUT95), .ZN(new_n666));
  XNOR2_X1  g480(.A(new_n664), .B(new_n666), .ZN(G12));
  INV_X1    g481(.A(new_n663), .ZN(new_n668));
  AOI21_X1  g482(.A(new_n668), .B1(new_n386), .B2(new_n392), .ZN(new_n669));
  INV_X1    g483(.A(new_n552), .ZN(new_n670));
  AOI21_X1  g484(.A(new_n507), .B1(new_n559), .B2(new_n508), .ZN(new_n671));
  OAI21_X1  g485(.A(new_n611), .B1(new_n670), .B2(new_n671), .ZN(new_n672));
  INV_X1    g486(.A(G900), .ZN(new_n673));
  AOI21_X1  g487(.A(new_n501), .B1(new_n673), .B2(new_n503), .ZN(new_n674));
  NOR3_X1   g488(.A1(new_n672), .A2(new_n654), .A3(new_n674), .ZN(new_n675));
  INV_X1    g489(.A(KEYINPUT96), .ZN(new_n676));
  NAND3_X1  g490(.A1(new_n675), .A2(new_n676), .A3(new_n495), .ZN(new_n677));
  INV_X1    g491(.A(new_n674), .ZN(new_n678));
  NAND4_X1  g492(.A1(new_n655), .A2(new_n495), .A3(new_n656), .A4(new_n678), .ZN(new_n679));
  NAND2_X1  g493(.A1(new_n679), .A2(KEYINPUT96), .ZN(new_n680));
  NAND4_X1  g494(.A1(new_n669), .A2(new_n454), .A3(new_n677), .A4(new_n680), .ZN(new_n681));
  XNOR2_X1  g495(.A(new_n681), .B(G128), .ZN(G30));
  OAI21_X1  g496(.A(new_n343), .B1(new_n315), .B2(new_n316), .ZN(new_n683));
  NAND2_X1  g497(.A1(new_n357), .A2(new_n683), .ZN(new_n684));
  AOI21_X1  g498(.A(new_n248), .B1(new_n684), .B2(new_n329), .ZN(new_n685));
  AOI21_X1  g499(.A(new_n685), .B1(new_n383), .B2(new_n385), .ZN(new_n686));
  NAND2_X1  g500(.A1(new_n686), .A2(new_n392), .ZN(new_n687));
  NAND2_X1  g501(.A1(new_n687), .A2(new_n668), .ZN(new_n688));
  XOR2_X1   g502(.A(new_n674), .B(KEYINPUT39), .Z(new_n689));
  NAND2_X1  g503(.A1(new_n454), .A2(new_n689), .ZN(new_n690));
  XNOR2_X1  g504(.A(new_n690), .B(KEYINPUT40), .ZN(new_n691));
  NAND2_X1  g505(.A1(new_n493), .A2(new_n494), .ZN(new_n692));
  XNOR2_X1  g506(.A(new_n692), .B(KEYINPUT38), .ZN(new_n693));
  NAND3_X1  g507(.A1(new_n693), .A2(new_n611), .A3(new_n455), .ZN(new_n694));
  NOR4_X1   g508(.A1(new_n688), .A2(new_n691), .A3(new_n694), .A4(new_n620), .ZN(new_n695));
  XOR2_X1   g509(.A(KEYINPUT97), .B(G143), .Z(new_n696));
  XNOR2_X1  g510(.A(new_n695), .B(new_n696), .ZN(G45));
  NAND3_X1  g511(.A1(new_n644), .A2(new_n495), .A3(new_n678), .ZN(new_n698));
  INV_X1    g512(.A(KEYINPUT98), .ZN(new_n699));
  NAND2_X1  g513(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  AOI211_X1 g514(.A(new_n674), .B(new_n643), .C1(new_n564), .C2(new_n616), .ZN(new_n701));
  NAND3_X1  g515(.A1(new_n701), .A2(KEYINPUT98), .A3(new_n495), .ZN(new_n702));
  NAND4_X1  g516(.A1(new_n700), .A2(new_n669), .A3(new_n702), .A4(new_n454), .ZN(new_n703));
  XNOR2_X1  g517(.A(new_n703), .B(G146), .ZN(G48));
  AOI211_X1 g518(.A(new_n643), .B(new_n622), .C1(new_n616), .C2(new_n564), .ZN(new_n705));
  OAI21_X1  g519(.A(new_n385), .B1(new_n387), .B2(new_n388), .ZN(new_n706));
  INV_X1    g520(.A(new_n356), .ZN(new_n707));
  OAI211_X1 g521(.A(new_n706), .B(new_n707), .C1(new_n635), .C2(new_n390), .ZN(new_n708));
  AND2_X1   g522(.A1(new_n243), .A2(new_n246), .ZN(new_n709));
  NOR2_X1   g523(.A1(new_n447), .A2(new_n398), .ZN(new_n710));
  INV_X1    g524(.A(new_n625), .ZN(new_n711));
  NOR3_X1   g525(.A1(new_n710), .A2(new_n711), .A3(new_n397), .ZN(new_n712));
  NAND4_X1  g526(.A1(new_n705), .A2(new_n708), .A3(new_n709), .A4(new_n712), .ZN(new_n713));
  XNOR2_X1  g527(.A(KEYINPUT41), .B(G113), .ZN(new_n714));
  XNOR2_X1  g528(.A(new_n713), .B(new_n714), .ZN(G15));
  NOR3_X1   g529(.A1(new_n672), .A2(new_n622), .A3(new_n654), .ZN(new_n716));
  NAND4_X1  g530(.A1(new_n708), .A2(new_n709), .A3(new_n712), .A4(new_n716), .ZN(new_n717));
  XNOR2_X1  g531(.A(new_n717), .B(G116), .ZN(G18));
  NAND3_X1  g532(.A1(new_n712), .A2(new_n505), .A3(new_n495), .ZN(new_n719));
  NOR2_X1   g533(.A1(new_n719), .A2(new_n617), .ZN(new_n720));
  NAND2_X1  g534(.A1(new_n669), .A2(new_n720), .ZN(new_n721));
  XNOR2_X1  g535(.A(new_n721), .B(G119), .ZN(G21));
  NAND2_X1  g536(.A1(new_n712), .A2(new_n505), .ZN(new_n723));
  NAND2_X1  g537(.A1(new_n495), .A2(new_n611), .ZN(new_n724));
  NOR3_X1   g538(.A1(new_n620), .A2(new_n723), .A3(new_n724), .ZN(new_n725));
  NAND2_X1  g539(.A1(new_n317), .A2(new_n319), .ZN(new_n726));
  AOI21_X1  g540(.A(new_n344), .B1(new_n726), .B2(KEYINPUT99), .ZN(new_n727));
  OAI21_X1  g541(.A(new_n727), .B1(KEYINPUT99), .B2(new_n726), .ZN(new_n728));
  AOI21_X1  g542(.A(new_n634), .B1(new_n728), .B2(new_n361), .ZN(new_n729));
  AOI211_X1 g543(.A(new_n247), .B(new_n729), .C1(new_n636), .C2(G472), .ZN(new_n730));
  NAND2_X1  g544(.A1(new_n725), .A2(new_n730), .ZN(new_n731));
  XNOR2_X1  g545(.A(new_n731), .B(G122), .ZN(G24));
  NAND2_X1  g546(.A1(new_n636), .A2(G472), .ZN(new_n733));
  INV_X1    g547(.A(new_n729), .ZN(new_n734));
  NAND3_X1  g548(.A1(new_n733), .A2(new_n663), .A3(new_n734), .ZN(new_n735));
  NAND4_X1  g549(.A1(new_n644), .A2(new_n495), .A3(new_n678), .A4(new_n712), .ZN(new_n736));
  NOR2_X1   g550(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  XNOR2_X1  g551(.A(new_n737), .B(new_n200), .ZN(G27));
  INV_X1    g552(.A(KEYINPUT100), .ZN(new_n739));
  NAND4_X1  g553(.A1(new_n451), .A2(new_n739), .A3(new_n452), .A4(G469), .ZN(new_n740));
  NAND3_X1  g554(.A1(new_n625), .A2(new_n740), .A3(new_n626), .ZN(new_n741));
  AND2_X1   g555(.A1(new_n453), .A2(KEYINPUT100), .ZN(new_n742));
  OAI21_X1  g556(.A(new_n628), .B1(new_n741), .B2(new_n742), .ZN(new_n743));
  NAND3_X1  g557(.A1(new_n493), .A2(new_n455), .A3(new_n494), .ZN(new_n744));
  NOR3_X1   g558(.A1(new_n743), .A2(new_n247), .A3(new_n744), .ZN(new_n745));
  NAND3_X1  g559(.A1(new_n708), .A2(new_n701), .A3(new_n745), .ZN(new_n746));
  NAND2_X1  g560(.A1(new_n746), .A2(KEYINPUT101), .ZN(new_n747));
  INV_X1    g561(.A(KEYINPUT42), .ZN(new_n748));
  INV_X1    g562(.A(KEYINPUT101), .ZN(new_n749));
  NAND4_X1  g563(.A1(new_n708), .A2(new_n749), .A3(new_n745), .A4(new_n701), .ZN(new_n750));
  NAND3_X1  g564(.A1(new_n747), .A2(new_n748), .A3(new_n750), .ZN(new_n751));
  NOR2_X1   g565(.A1(new_n743), .A2(new_n744), .ZN(new_n752));
  NAND3_X1  g566(.A1(new_n701), .A2(KEYINPUT42), .A3(new_n752), .ZN(new_n753));
  INV_X1    g567(.A(new_n753), .ZN(new_n754));
  OAI211_X1 g568(.A(new_n706), .B(new_n707), .C1(new_n635), .C2(KEYINPUT32), .ZN(new_n755));
  INV_X1    g569(.A(KEYINPUT102), .ZN(new_n756));
  AND3_X1   g570(.A1(new_n755), .A2(new_n756), .A3(new_n709), .ZN(new_n757));
  AOI21_X1  g571(.A(new_n756), .B1(new_n755), .B2(new_n709), .ZN(new_n758));
  OAI21_X1  g572(.A(new_n754), .B1(new_n757), .B2(new_n758), .ZN(new_n759));
  NAND2_X1  g573(.A1(new_n751), .A2(new_n759), .ZN(new_n760));
  XNOR2_X1  g574(.A(new_n760), .B(G131), .ZN(G33));
  NAND2_X1  g575(.A1(new_n453), .A2(KEYINPUT100), .ZN(new_n762));
  NAND3_X1  g576(.A1(new_n448), .A2(new_n762), .A3(new_n740), .ZN(new_n763));
  NOR3_X1   g577(.A1(new_n621), .A2(new_n492), .A3(new_n456), .ZN(new_n764));
  NAND4_X1  g578(.A1(new_n709), .A2(new_n763), .A3(new_n764), .A4(new_n628), .ZN(new_n765));
  AOI21_X1  g579(.A(new_n765), .B1(new_n386), .B2(new_n392), .ZN(new_n766));
  NAND2_X1  g580(.A1(new_n766), .A2(new_n675), .ZN(new_n767));
  XNOR2_X1  g581(.A(new_n767), .B(G134), .ZN(G36));
  XNOR2_X1  g582(.A(new_n619), .B(KEYINPUT105), .ZN(new_n769));
  INV_X1    g583(.A(new_n643), .ZN(new_n770));
  NAND3_X1  g584(.A1(new_n769), .A2(KEYINPUT43), .A3(new_n770), .ZN(new_n771));
  INV_X1    g585(.A(KEYINPUT43), .ZN(new_n772));
  XNOR2_X1  g586(.A(new_n643), .B(KEYINPUT104), .ZN(new_n773));
  OAI21_X1  g587(.A(new_n772), .B1(new_n773), .B2(new_n619), .ZN(new_n774));
  NAND2_X1  g588(.A1(new_n771), .A2(new_n774), .ZN(new_n775));
  INV_X1    g589(.A(new_n637), .ZN(new_n776));
  NAND3_X1  g590(.A1(new_n775), .A2(new_n776), .A3(new_n663), .ZN(new_n777));
  INV_X1    g591(.A(KEYINPUT44), .ZN(new_n778));
  OR2_X1    g592(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  NAND2_X1  g593(.A1(new_n777), .A2(new_n778), .ZN(new_n780));
  INV_X1    g594(.A(KEYINPUT46), .ZN(new_n781));
  NAND2_X1  g595(.A1(new_n451), .A2(new_n452), .ZN(new_n782));
  INV_X1    g596(.A(KEYINPUT45), .ZN(new_n783));
  NAND2_X1  g597(.A1(new_n782), .A2(new_n783), .ZN(new_n784));
  NAND3_X1  g598(.A1(new_n451), .A2(KEYINPUT45), .A3(new_n452), .ZN(new_n785));
  NAND3_X1  g599(.A1(new_n784), .A2(G469), .A3(new_n785), .ZN(new_n786));
  INV_X1    g600(.A(new_n786), .ZN(new_n787));
  OAI21_X1  g601(.A(new_n781), .B1(new_n787), .B2(new_n399), .ZN(new_n788));
  NAND3_X1  g602(.A1(new_n786), .A2(KEYINPUT46), .A3(new_n626), .ZN(new_n789));
  NAND3_X1  g603(.A1(new_n788), .A2(new_n625), .A3(new_n789), .ZN(new_n790));
  NAND3_X1  g604(.A1(new_n790), .A2(new_n628), .A3(new_n689), .ZN(new_n791));
  XNOR2_X1  g605(.A(new_n791), .B(KEYINPUT103), .ZN(new_n792));
  XNOR2_X1  g606(.A(new_n744), .B(KEYINPUT106), .ZN(new_n793));
  NAND4_X1  g607(.A1(new_n779), .A2(new_n780), .A3(new_n792), .A4(new_n793), .ZN(new_n794));
  XOR2_X1   g608(.A(KEYINPUT107), .B(G137), .Z(new_n795));
  XNOR2_X1  g609(.A(new_n794), .B(new_n795), .ZN(G39));
  NAND2_X1  g610(.A1(new_n790), .A2(new_n628), .ZN(new_n797));
  XNOR2_X1  g611(.A(new_n797), .B(KEYINPUT47), .ZN(new_n798));
  INV_X1    g612(.A(new_n708), .ZN(new_n799));
  NAND4_X1  g613(.A1(new_n799), .A2(new_n247), .A3(new_n701), .A4(new_n764), .ZN(new_n800));
  NOR2_X1   g614(.A1(new_n798), .A2(new_n800), .ZN(new_n801));
  XNOR2_X1  g615(.A(new_n801), .B(new_n204), .ZN(G42));
  NOR2_X1   g616(.A1(new_n710), .A2(new_n711), .ZN(new_n803));
  INV_X1    g617(.A(new_n803), .ZN(new_n804));
  AOI21_X1  g618(.A(new_n643), .B1(new_n804), .B2(KEYINPUT49), .ZN(new_n805));
  OAI21_X1  g619(.A(new_n805), .B1(KEYINPUT49), .B2(new_n804), .ZN(new_n806));
  NAND3_X1  g620(.A1(new_n709), .A2(new_n455), .A3(new_n628), .ZN(new_n807));
  NOR3_X1   g621(.A1(new_n806), .A2(new_n693), .A3(new_n807), .ZN(new_n808));
  INV_X1    g622(.A(new_n687), .ZN(new_n809));
  NAND3_X1  g623(.A1(new_n808), .A2(new_n809), .A3(new_n769), .ZN(new_n810));
  XOR2_X1   g624(.A(new_n810), .B(KEYINPUT108), .Z(new_n811));
  INV_X1    g625(.A(KEYINPUT51), .ZN(new_n812));
  AOI21_X1  g626(.A(new_n500), .B1(new_n771), .B2(new_n774), .ZN(new_n813));
  AND2_X1   g627(.A1(new_n813), .A2(new_n730), .ZN(new_n814));
  AND2_X1   g628(.A1(new_n814), .A2(new_n793), .ZN(new_n815));
  OR2_X1    g629(.A1(new_n815), .A2(KEYINPUT111), .ZN(new_n816));
  NAND2_X1  g630(.A1(new_n815), .A2(KEYINPUT111), .ZN(new_n817));
  OAI21_X1  g631(.A(new_n798), .B1(new_n628), .B2(new_n804), .ZN(new_n818));
  AND3_X1   g632(.A1(new_n816), .A2(new_n817), .A3(new_n818), .ZN(new_n819));
  INV_X1    g633(.A(new_n712), .ZN(new_n820));
  NOR3_X1   g634(.A1(new_n693), .A2(new_n455), .A3(new_n820), .ZN(new_n821));
  NAND2_X1  g635(.A1(new_n814), .A2(new_n821), .ZN(new_n822));
  XOR2_X1   g636(.A(KEYINPUT112), .B(KEYINPUT50), .Z(new_n823));
  NAND2_X1  g637(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  AND3_X1   g638(.A1(new_n813), .A2(new_n712), .A3(new_n764), .ZN(new_n825));
  AOI21_X1  g639(.A(new_n729), .B1(new_n636), .B2(G472), .ZN(new_n826));
  NAND3_X1  g640(.A1(new_n825), .A2(new_n663), .A3(new_n826), .ZN(new_n827));
  NOR4_X1   g641(.A1(new_n820), .A2(new_n247), .A3(new_n500), .A4(new_n744), .ZN(new_n828));
  NAND4_X1  g642(.A1(new_n809), .A2(new_n620), .A3(new_n643), .A4(new_n828), .ZN(new_n829));
  AND3_X1   g643(.A1(new_n824), .A2(new_n827), .A3(new_n829), .ZN(new_n830));
  NOR2_X1   g644(.A1(KEYINPUT112), .A2(KEYINPUT50), .ZN(new_n831));
  NAND3_X1  g645(.A1(new_n814), .A2(new_n831), .A3(new_n821), .ZN(new_n832));
  NAND2_X1  g646(.A1(new_n830), .A2(new_n832), .ZN(new_n833));
  OAI21_X1  g647(.A(new_n812), .B1(new_n819), .B2(new_n833), .ZN(new_n834));
  INV_X1    g648(.A(KEYINPUT113), .ZN(new_n835));
  NAND2_X1  g649(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  OAI211_X1 g650(.A(KEYINPUT113), .B(new_n812), .C1(new_n819), .C2(new_n833), .ZN(new_n837));
  AND2_X1   g651(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  INV_X1    g652(.A(KEYINPUT54), .ZN(new_n839));
  INV_X1    g653(.A(new_n737), .ZN(new_n840));
  NOR4_X1   g654(.A1(new_n620), .A2(new_n724), .A3(new_n743), .A4(new_n674), .ZN(new_n841));
  NAND3_X1  g655(.A1(new_n841), .A2(new_n668), .A3(new_n687), .ZN(new_n842));
  NAND4_X1  g656(.A1(new_n703), .A2(new_n840), .A3(new_n681), .A4(new_n842), .ZN(new_n843));
  NAND2_X1  g657(.A1(new_n843), .A2(KEYINPUT52), .ZN(new_n844));
  AND2_X1   g658(.A1(new_n677), .A2(new_n680), .ZN(new_n845));
  AOI211_X1 g659(.A(new_n629), .B(new_n668), .C1(new_n386), .C2(new_n392), .ZN(new_n846));
  AOI21_X1  g660(.A(new_n737), .B1(new_n845), .B2(new_n846), .ZN(new_n847));
  INV_X1    g661(.A(KEYINPUT52), .ZN(new_n848));
  NAND4_X1  g662(.A1(new_n847), .A2(new_n848), .A3(new_n703), .A4(new_n842), .ZN(new_n849));
  NAND2_X1  g663(.A1(new_n844), .A2(new_n849), .ZN(new_n850));
  INV_X1    g664(.A(new_n850), .ZN(new_n851));
  OAI211_X1 g665(.A(new_n612), .B(new_n678), .C1(new_n670), .C2(new_n671), .ZN(new_n852));
  NOR3_X1   g666(.A1(new_n852), .A2(new_n654), .A3(new_n744), .ZN(new_n853));
  NAND4_X1  g667(.A1(new_n853), .A2(new_n708), .A3(new_n454), .A4(new_n663), .ZN(new_n854));
  NAND4_X1  g668(.A1(new_n826), .A2(new_n701), .A3(new_n663), .A4(new_n752), .ZN(new_n855));
  NAND3_X1  g669(.A1(new_n854), .A2(new_n767), .A3(new_n855), .ZN(new_n856));
  AOI21_X1  g670(.A(new_n856), .B1(new_n751), .B2(new_n759), .ZN(new_n857));
  NAND4_X1  g671(.A1(new_n632), .A2(new_n664), .A3(new_n713), .A4(new_n717), .ZN(new_n858));
  NAND2_X1  g672(.A1(new_n619), .A2(new_n643), .ZN(new_n859));
  NAND4_X1  g673(.A1(new_n637), .A2(new_n617), .A3(new_n645), .A4(new_n859), .ZN(new_n860));
  NAND3_X1  g674(.A1(new_n721), .A2(new_n731), .A3(new_n860), .ZN(new_n861));
  NOR2_X1   g675(.A1(new_n858), .A2(new_n861), .ZN(new_n862));
  INV_X1    g676(.A(KEYINPUT109), .ZN(new_n863));
  AND3_X1   g677(.A1(new_n857), .A2(new_n862), .A3(new_n863), .ZN(new_n864));
  AOI21_X1  g678(.A(new_n863), .B1(new_n857), .B2(new_n862), .ZN(new_n865));
  OAI21_X1  g679(.A(new_n851), .B1(new_n864), .B2(new_n865), .ZN(new_n866));
  INV_X1    g680(.A(KEYINPUT53), .ZN(new_n867));
  NAND2_X1  g681(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  OAI21_X1  g682(.A(new_n867), .B1(new_n847), .B2(new_n848), .ZN(new_n869));
  OAI211_X1 g683(.A(new_n851), .B(new_n869), .C1(new_n864), .C2(new_n865), .ZN(new_n870));
  AOI21_X1  g684(.A(new_n839), .B1(new_n868), .B2(new_n870), .ZN(new_n871));
  NAND2_X1  g685(.A1(new_n840), .A2(new_n681), .ZN(new_n872));
  AOI21_X1  g686(.A(new_n867), .B1(new_n872), .B2(KEYINPUT52), .ZN(new_n873));
  NAND3_X1  g687(.A1(new_n844), .A2(new_n849), .A3(new_n873), .ZN(new_n874));
  NAND2_X1  g688(.A1(new_n857), .A2(new_n862), .ZN(new_n875));
  NOR2_X1   g689(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  AOI211_X1 g690(.A(KEYINPUT54), .B(new_n876), .C1(new_n866), .C2(new_n867), .ZN(new_n877));
  OAI21_X1  g691(.A(KEYINPUT110), .B1(new_n871), .B2(new_n877), .ZN(new_n878));
  AND3_X1   g692(.A1(new_n854), .A2(new_n767), .A3(new_n855), .ZN(new_n879));
  NAND2_X1  g693(.A1(new_n750), .A2(new_n748), .ZN(new_n880));
  AOI21_X1  g694(.A(new_n749), .B1(new_n766), .B2(new_n701), .ZN(new_n881));
  NOR2_X1   g695(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  NAND2_X1  g696(.A1(new_n755), .A2(new_n709), .ZN(new_n883));
  NAND2_X1  g697(.A1(new_n883), .A2(KEYINPUT102), .ZN(new_n884));
  NAND3_X1  g698(.A1(new_n755), .A2(new_n756), .A3(new_n709), .ZN(new_n885));
  AOI21_X1  g699(.A(new_n753), .B1(new_n884), .B2(new_n885), .ZN(new_n886));
  OAI21_X1  g700(.A(new_n879), .B1(new_n882), .B2(new_n886), .ZN(new_n887));
  AND2_X1   g701(.A1(new_n713), .A2(new_n717), .ZN(new_n888));
  NAND3_X1  g702(.A1(new_n733), .A2(new_n389), .A3(new_n663), .ZN(new_n889));
  INV_X1    g703(.A(new_n889), .ZN(new_n890));
  OAI211_X1 g704(.A(new_n618), .B(new_n631), .C1(new_n890), .C2(new_n393), .ZN(new_n891));
  AOI22_X1  g705(.A1(new_n669), .A2(new_n720), .B1(new_n725), .B2(new_n730), .ZN(new_n892));
  NAND4_X1  g706(.A1(new_n888), .A2(new_n891), .A3(new_n860), .A4(new_n892), .ZN(new_n893));
  OAI21_X1  g707(.A(KEYINPUT109), .B1(new_n887), .B2(new_n893), .ZN(new_n894));
  NAND3_X1  g708(.A1(new_n857), .A2(new_n862), .A3(new_n863), .ZN(new_n895));
  AOI21_X1  g709(.A(new_n850), .B1(new_n894), .B2(new_n895), .ZN(new_n896));
  OAI21_X1  g710(.A(new_n870), .B1(new_n896), .B2(KEYINPUT53), .ZN(new_n897));
  NAND2_X1  g711(.A1(new_n897), .A2(KEYINPUT54), .ZN(new_n898));
  INV_X1    g712(.A(KEYINPUT110), .ZN(new_n899));
  OR2_X1    g713(.A1(new_n874), .A2(new_n875), .ZN(new_n900));
  OAI211_X1 g714(.A(new_n839), .B(new_n900), .C1(new_n896), .C2(KEYINPUT53), .ZN(new_n901));
  NAND3_X1  g715(.A1(new_n898), .A2(new_n899), .A3(new_n901), .ZN(new_n902));
  NAND2_X1  g716(.A1(new_n878), .A2(new_n902), .ZN(new_n903));
  NAND3_X1  g717(.A1(new_n816), .A2(new_n817), .A3(new_n818), .ZN(new_n904));
  NAND4_X1  g718(.A1(new_n904), .A2(KEYINPUT51), .A3(new_n832), .A4(new_n830), .ZN(new_n905));
  NAND2_X1  g719(.A1(new_n884), .A2(new_n885), .ZN(new_n906));
  NAND2_X1  g720(.A1(new_n825), .A2(new_n906), .ZN(new_n907));
  XNOR2_X1  g721(.A(new_n907), .B(KEYINPUT48), .ZN(new_n908));
  NAND3_X1  g722(.A1(new_n814), .A2(new_n495), .A3(new_n712), .ZN(new_n909));
  NAND3_X1  g723(.A1(new_n809), .A2(new_n644), .A3(new_n828), .ZN(new_n910));
  AND3_X1   g724(.A1(new_n909), .A2(new_n498), .A3(new_n910), .ZN(new_n911));
  NAND3_X1  g725(.A1(new_n905), .A2(new_n908), .A3(new_n911), .ZN(new_n912));
  NOR3_X1   g726(.A1(new_n838), .A2(new_n903), .A3(new_n912), .ZN(new_n913));
  NOR2_X1   g727(.A1(G952), .A2(G953), .ZN(new_n914));
  XOR2_X1   g728(.A(new_n914), .B(KEYINPUT114), .Z(new_n915));
  OAI21_X1  g729(.A(new_n811), .B1(new_n913), .B2(new_n915), .ZN(G75));
  NOR2_X1   g730(.A1(new_n434), .A2(G952), .ZN(new_n917));
  OAI21_X1  g731(.A(new_n900), .B1(new_n896), .B2(KEYINPUT53), .ZN(new_n918));
  INV_X1    g732(.A(new_n918), .ZN(new_n919));
  NOR2_X1   g733(.A1(new_n919), .A2(new_n329), .ZN(new_n920));
  NAND2_X1  g734(.A1(new_n920), .A2(G210), .ZN(new_n921));
  INV_X1    g735(.A(KEYINPUT56), .ZN(new_n922));
  NAND2_X1  g736(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  NAND2_X1  g737(.A1(new_n472), .A2(new_n473), .ZN(new_n924));
  XOR2_X1   g738(.A(new_n924), .B(new_n482), .Z(new_n925));
  XNOR2_X1  g739(.A(new_n925), .B(KEYINPUT55), .ZN(new_n926));
  AOI21_X1  g740(.A(new_n917), .B1(new_n923), .B2(new_n926), .ZN(new_n927));
  INV_X1    g741(.A(KEYINPUT115), .ZN(new_n928));
  NAND2_X1  g742(.A1(new_n921), .A2(new_n928), .ZN(new_n929));
  NAND3_X1  g743(.A1(new_n920), .A2(KEYINPUT115), .A3(G210), .ZN(new_n930));
  NOR2_X1   g744(.A1(new_n926), .A2(KEYINPUT56), .ZN(new_n931));
  NAND3_X1  g745(.A1(new_n929), .A2(new_n930), .A3(new_n931), .ZN(new_n932));
  AND2_X1   g746(.A1(new_n927), .A2(new_n932), .ZN(G51));
  NAND2_X1  g747(.A1(new_n918), .A2(KEYINPUT54), .ZN(new_n934));
  INV_X1    g748(.A(KEYINPUT116), .ZN(new_n935));
  NAND3_X1  g749(.A1(new_n934), .A2(new_n935), .A3(new_n901), .ZN(new_n936));
  NAND3_X1  g750(.A1(new_n918), .A2(KEYINPUT116), .A3(KEYINPUT54), .ZN(new_n937));
  XNOR2_X1  g751(.A(new_n399), .B(KEYINPUT57), .ZN(new_n938));
  NAND3_X1  g752(.A1(new_n936), .A2(new_n937), .A3(new_n938), .ZN(new_n939));
  INV_X1    g753(.A(KEYINPUT117), .ZN(new_n940));
  NAND2_X1  g754(.A1(new_n437), .A2(new_n446), .ZN(new_n941));
  NAND3_X1  g755(.A1(new_n939), .A2(new_n940), .A3(new_n941), .ZN(new_n942));
  NAND2_X1  g756(.A1(new_n920), .A2(new_n787), .ZN(new_n943));
  AND2_X1   g757(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  NAND2_X1  g758(.A1(new_n939), .A2(new_n941), .ZN(new_n945));
  NAND2_X1  g759(.A1(new_n945), .A2(KEYINPUT117), .ZN(new_n946));
  AOI21_X1  g760(.A(new_n917), .B1(new_n944), .B2(new_n946), .ZN(G54));
  NAND3_X1  g761(.A1(new_n920), .A2(KEYINPUT58), .A3(G475), .ZN(new_n948));
  INV_X1    g762(.A(new_n559), .ZN(new_n949));
  AND2_X1   g763(.A1(new_n948), .A2(new_n949), .ZN(new_n950));
  NOR2_X1   g764(.A1(new_n948), .A2(new_n949), .ZN(new_n951));
  NOR3_X1   g765(.A1(new_n950), .A2(new_n951), .A3(new_n917), .ZN(G60));
  XOR2_X1   g766(.A(KEYINPUT118), .B(KEYINPUT59), .Z(new_n953));
  NOR2_X1   g767(.A1(new_n603), .A2(new_n329), .ZN(new_n954));
  XNOR2_X1  g768(.A(new_n953), .B(new_n954), .ZN(new_n955));
  NOR3_X1   g769(.A1(new_n871), .A2(new_n877), .A3(KEYINPUT110), .ZN(new_n956));
  AOI21_X1  g770(.A(new_n899), .B1(new_n898), .B2(new_n901), .ZN(new_n957));
  OAI21_X1  g771(.A(new_n955), .B1(new_n956), .B2(new_n957), .ZN(new_n958));
  INV_X1    g772(.A(new_n640), .ZN(new_n959));
  NAND2_X1  g773(.A1(new_n958), .A2(new_n959), .ZN(new_n960));
  NAND4_X1  g774(.A1(new_n936), .A2(new_n640), .A3(new_n937), .A4(new_n955), .ZN(new_n961));
  INV_X1    g775(.A(new_n917), .ZN(new_n962));
  AND2_X1   g776(.A1(new_n961), .A2(new_n962), .ZN(new_n963));
  NAND3_X1  g777(.A1(new_n960), .A2(new_n963), .A3(KEYINPUT119), .ZN(new_n964));
  INV_X1    g778(.A(KEYINPUT119), .ZN(new_n965));
  AOI21_X1  g779(.A(new_n640), .B1(new_n903), .B2(new_n955), .ZN(new_n966));
  NAND2_X1  g780(.A1(new_n961), .A2(new_n962), .ZN(new_n967));
  OAI21_X1  g781(.A(new_n965), .B1(new_n966), .B2(new_n967), .ZN(new_n968));
  NAND2_X1  g782(.A1(new_n964), .A2(new_n968), .ZN(G63));
  NAND2_X1  g783(.A1(G217), .A2(G902), .ZN(new_n970));
  XNOR2_X1  g784(.A(new_n970), .B(KEYINPUT60), .ZN(new_n971));
  NOR2_X1   g785(.A1(new_n919), .A2(new_n971), .ZN(new_n972));
  NAND2_X1  g786(.A1(new_n972), .A2(new_n661), .ZN(new_n973));
  OR2_X1    g787(.A1(new_n973), .A2(KEYINPUT120), .ZN(new_n974));
  OAI21_X1  g788(.A(new_n962), .B1(new_n972), .B2(new_n244), .ZN(new_n975));
  INV_X1    g789(.A(KEYINPUT121), .ZN(new_n976));
  NAND2_X1  g790(.A1(new_n975), .A2(new_n976), .ZN(new_n977));
  OAI221_X1 g791(.A(new_n962), .B1(KEYINPUT121), .B2(KEYINPUT61), .C1(new_n972), .C2(new_n244), .ZN(new_n978));
  NAND2_X1  g792(.A1(new_n973), .A2(KEYINPUT120), .ZN(new_n979));
  NAND4_X1  g793(.A1(new_n974), .A2(new_n977), .A3(new_n978), .A4(new_n979), .ZN(new_n980));
  INV_X1    g794(.A(new_n973), .ZN(new_n981));
  OAI21_X1  g795(.A(KEYINPUT61), .B1(new_n978), .B2(new_n981), .ZN(new_n982));
  AND2_X1   g796(.A1(new_n980), .A2(new_n982), .ZN(G66));
  INV_X1    g797(.A(G224), .ZN(new_n984));
  OAI21_X1  g798(.A(G953), .B1(new_n502), .B2(new_n984), .ZN(new_n985));
  XOR2_X1   g799(.A(new_n985), .B(KEYINPUT123), .Z(new_n986));
  XNOR2_X1  g800(.A(new_n862), .B(KEYINPUT122), .ZN(new_n987));
  OAI21_X1  g801(.A(new_n986), .B1(new_n987), .B2(G953), .ZN(new_n988));
  XOR2_X1   g802(.A(new_n988), .B(KEYINPUT124), .Z(new_n989));
  OAI21_X1  g803(.A(new_n924), .B1(G898), .B2(new_n434), .ZN(new_n990));
  XNOR2_X1  g804(.A(new_n989), .B(new_n990), .ZN(G69));
  NAND2_X1  g805(.A1(new_n346), .A2(new_n348), .ZN(new_n992));
  XOR2_X1   g806(.A(new_n992), .B(new_n537), .Z(new_n993));
  AND2_X1   g807(.A1(new_n847), .A2(new_n703), .ZN(new_n994));
  INV_X1    g808(.A(KEYINPUT125), .ZN(new_n995));
  XNOR2_X1  g809(.A(new_n994), .B(new_n995), .ZN(new_n996));
  OR3_X1    g810(.A1(new_n996), .A2(KEYINPUT62), .A3(new_n695), .ZN(new_n997));
  OAI21_X1  g811(.A(KEYINPUT62), .B1(new_n996), .B2(new_n695), .ZN(new_n998));
  INV_X1    g812(.A(new_n801), .ZN(new_n999));
  NOR2_X1   g813(.A1(new_n690), .A2(new_n744), .ZN(new_n1000));
  NAND4_X1  g814(.A1(new_n393), .A2(new_n617), .A3(new_n859), .A4(new_n1000), .ZN(new_n1001));
  AND3_X1   g815(.A1(new_n794), .A2(new_n999), .A3(new_n1001), .ZN(new_n1002));
  NAND3_X1  g816(.A1(new_n997), .A2(new_n998), .A3(new_n1002), .ZN(new_n1003));
  AOI21_X1  g817(.A(new_n993), .B1(new_n1003), .B2(new_n434), .ZN(new_n1004));
  INV_X1    g818(.A(new_n993), .ZN(new_n1005));
  NOR2_X1   g819(.A1(new_n673), .A2(new_n434), .ZN(new_n1006));
  NOR2_X1   g820(.A1(new_n620), .A2(new_n724), .ZN(new_n1007));
  NAND3_X1  g821(.A1(new_n792), .A2(new_n1007), .A3(new_n906), .ZN(new_n1008));
  AND4_X1   g822(.A1(new_n760), .A2(new_n999), .A3(new_n767), .A4(new_n1008), .ZN(new_n1009));
  NAND2_X1  g823(.A1(new_n1009), .A2(new_n794), .ZN(new_n1010));
  NOR2_X1   g824(.A1(new_n1010), .A2(new_n996), .ZN(new_n1011));
  AOI211_X1 g825(.A(new_n1005), .B(new_n1006), .C1(new_n1011), .C2(new_n434), .ZN(new_n1012));
  AOI21_X1  g826(.A(new_n434), .B1(G227), .B2(G900), .ZN(new_n1013));
  INV_X1    g827(.A(KEYINPUT126), .ZN(new_n1014));
  AND2_X1   g828(.A1(new_n1013), .A2(new_n1014), .ZN(new_n1015));
  NOR3_X1   g829(.A1(new_n1004), .A2(new_n1012), .A3(new_n1015), .ZN(new_n1016));
  NOR2_X1   g830(.A1(new_n1013), .A2(new_n1014), .ZN(new_n1017));
  XNOR2_X1  g831(.A(new_n1016), .B(new_n1017), .ZN(G72));
  NAND2_X1  g832(.A1(G472), .A2(G902), .ZN(new_n1019));
  XOR2_X1   g833(.A(new_n1019), .B(KEYINPUT63), .Z(new_n1020));
  INV_X1    g834(.A(new_n1020), .ZN(new_n1021));
  AOI21_X1  g835(.A(new_n1021), .B1(new_n1011), .B2(new_n987), .ZN(new_n1022));
  XOR2_X1   g836(.A(new_n350), .B(KEYINPUT127), .Z(new_n1023));
  INV_X1    g837(.A(new_n1023), .ZN(new_n1024));
  NAND2_X1  g838(.A1(new_n1024), .A2(new_n325), .ZN(new_n1025));
  OAI21_X1  g839(.A(new_n962), .B1(new_n1022), .B2(new_n1025), .ZN(new_n1026));
  NAND4_X1  g840(.A1(new_n997), .A2(new_n987), .A3(new_n998), .A4(new_n1002), .ZN(new_n1027));
  AOI211_X1 g841(.A(new_n325), .B(new_n1024), .C1(new_n1027), .C2(new_n1020), .ZN(new_n1028));
  AOI21_X1  g842(.A(new_n1021), .B1(new_n351), .B2(new_n357), .ZN(new_n1029));
  AOI211_X1 g843(.A(new_n1026), .B(new_n1028), .C1(new_n897), .C2(new_n1029), .ZN(G57));
endmodule


