

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304,
         n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315,
         n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326,
         n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, n337,
         n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, n348,
         n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359,
         n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370,
         n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381,
         n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392,
         n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403,
         n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414,
         n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425,
         n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436,
         n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447,
         n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458,
         n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469,
         n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480,
         n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491,
         n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502,
         n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513,
         n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591;

  AND2_X1 U326 ( .A1(n387), .A2(n473), .ZN(n388) );
  XNOR2_X1 U327 ( .A(n378), .B(n377), .ZN(n379) );
  XOR2_X1 U328 ( .A(G176GAT), .B(KEYINPUT82), .Z(n294) );
  XOR2_X1 U329 ( .A(n435), .B(n371), .Z(n295) );
  INV_X1 U330 ( .A(KEYINPUT98), .ZN(n385) );
  INV_X1 U331 ( .A(KEYINPUT48), .ZN(n467) );
  XNOR2_X1 U332 ( .A(n467), .B(KEYINPUT64), .ZN(n468) );
  XOR2_X1 U333 ( .A(KEYINPUT75), .B(G162GAT), .Z(n318) );
  XNOR2_X1 U334 ( .A(n469), .B(n468), .ZN(n530) );
  INV_X1 U335 ( .A(KEYINPUT85), .ZN(n375) );
  XNOR2_X1 U336 ( .A(n376), .B(n375), .ZN(n377) );
  NAND2_X1 U337 ( .A1(n415), .A2(n414), .ZN(n481) );
  NOR2_X1 U338 ( .A1(n589), .A2(n417), .ZN(n418) );
  XOR2_X1 U339 ( .A(KEYINPUT36), .B(n561), .Z(n589) );
  XOR2_X1 U340 ( .A(n334), .B(n333), .Z(n561) );
  XNOR2_X1 U341 ( .A(n382), .B(n381), .ZN(n521) );
  XNOR2_X1 U342 ( .A(KEYINPUT38), .B(n451), .ZN(n501) );
  XNOR2_X1 U343 ( .A(G190GAT), .B(KEYINPUT58), .ZN(n476) );
  INV_X1 U344 ( .A(G50GAT), .ZN(n452) );
  XNOR2_X1 U345 ( .A(n477), .B(n476), .ZN(G1351GAT) );
  XNOR2_X1 U346 ( .A(n453), .B(n452), .ZN(G1331GAT) );
  XNOR2_X1 U347 ( .A(KEYINPUT28), .B(KEYINPUT66), .ZN(n315) );
  XOR2_X1 U348 ( .A(G211GAT), .B(KEYINPUT21), .Z(n297) );
  XNOR2_X1 U349 ( .A(G197GAT), .B(G218GAT), .ZN(n296) );
  XNOR2_X1 U350 ( .A(n297), .B(n296), .ZN(n358) );
  XOR2_X1 U351 ( .A(n358), .B(G204GAT), .Z(n299) );
  NAND2_X1 U352 ( .A1(G228GAT), .A2(G233GAT), .ZN(n298) );
  XNOR2_X1 U353 ( .A(n299), .B(n298), .ZN(n314) );
  XOR2_X1 U354 ( .A(G78GAT), .B(G148GAT), .Z(n301) );
  XNOR2_X1 U355 ( .A(G106GAT), .B(KEYINPUT72), .ZN(n300) );
  XNOR2_X1 U356 ( .A(n301), .B(n300), .ZN(n440) );
  XOR2_X1 U357 ( .A(n440), .B(KEYINPUT89), .Z(n303) );
  XNOR2_X1 U358 ( .A(n318), .B(KEYINPUT22), .ZN(n302) );
  XNOR2_X1 U359 ( .A(n303), .B(n302), .ZN(n307) );
  XOR2_X1 U360 ( .A(KEYINPUT86), .B(KEYINPUT24), .Z(n305) );
  XNOR2_X1 U361 ( .A(KEYINPUT23), .B(KEYINPUT87), .ZN(n304) );
  XNOR2_X1 U362 ( .A(n305), .B(n304), .ZN(n306) );
  XOR2_X1 U363 ( .A(n307), .B(n306), .Z(n312) );
  XNOR2_X1 U364 ( .A(G50GAT), .B(G22GAT), .ZN(n308) );
  XNOR2_X1 U365 ( .A(n308), .B(G141GAT), .ZN(n423) );
  XOR2_X1 U366 ( .A(G155GAT), .B(KEYINPUT3), .Z(n310) );
  XNOR2_X1 U367 ( .A(KEYINPUT2), .B(KEYINPUT88), .ZN(n309) );
  XNOR2_X1 U368 ( .A(n310), .B(n309), .ZN(n406) );
  XNOR2_X1 U369 ( .A(n423), .B(n406), .ZN(n311) );
  XNOR2_X1 U370 ( .A(n312), .B(n311), .ZN(n313) );
  XNOR2_X1 U371 ( .A(n314), .B(n313), .ZN(n473) );
  XNOR2_X1 U372 ( .A(n315), .B(n473), .ZN(n534) );
  INV_X1 U373 ( .A(KEYINPUT104), .ZN(n450) );
  XOR2_X1 U374 ( .A(KEYINPUT77), .B(KEYINPUT11), .Z(n317) );
  XNOR2_X1 U375 ( .A(G190GAT), .B(KEYINPUT10), .ZN(n316) );
  XNOR2_X1 U376 ( .A(n317), .B(n316), .ZN(n334) );
  XOR2_X1 U377 ( .A(n318), .B(G92GAT), .Z(n320) );
  NAND2_X1 U378 ( .A1(G232GAT), .A2(G233GAT), .ZN(n319) );
  XOR2_X1 U379 ( .A(n320), .B(n319), .Z(n327) );
  XOR2_X1 U380 ( .A(KEYINPUT76), .B(KEYINPUT9), .Z(n322) );
  XNOR2_X1 U381 ( .A(G106GAT), .B(KEYINPUT78), .ZN(n321) );
  XNOR2_X1 U382 ( .A(n322), .B(n321), .ZN(n323) );
  XOR2_X1 U383 ( .A(G99GAT), .B(G85GAT), .Z(n434) );
  XNOR2_X1 U384 ( .A(n323), .B(n434), .ZN(n325) );
  XOR2_X1 U385 ( .A(G134GAT), .B(G218GAT), .Z(n324) );
  XNOR2_X1 U386 ( .A(n325), .B(n324), .ZN(n326) );
  XNOR2_X1 U387 ( .A(n327), .B(n326), .ZN(n332) );
  XOR2_X1 U388 ( .A(KEYINPUT8), .B(G43GAT), .Z(n329) );
  XNOR2_X1 U389 ( .A(G36GAT), .B(G29GAT), .ZN(n328) );
  XNOR2_X1 U390 ( .A(n329), .B(n328), .ZN(n330) );
  XOR2_X1 U391 ( .A(KEYINPUT7), .B(n330), .Z(n431) );
  XNOR2_X1 U392 ( .A(n431), .B(G50GAT), .ZN(n331) );
  XNOR2_X1 U393 ( .A(n332), .B(n331), .ZN(n333) );
  XOR2_X1 U394 ( .A(G211GAT), .B(G155GAT), .Z(n336) );
  XNOR2_X1 U395 ( .A(G183GAT), .B(G71GAT), .ZN(n335) );
  XNOR2_X1 U396 ( .A(n336), .B(n335), .ZN(n337) );
  XOR2_X1 U397 ( .A(G57GAT), .B(KEYINPUT13), .Z(n444) );
  XOR2_X1 U398 ( .A(n337), .B(n444), .Z(n339) );
  XNOR2_X1 U399 ( .A(G22GAT), .B(G78GAT), .ZN(n338) );
  XNOR2_X1 U400 ( .A(n339), .B(n338), .ZN(n344) );
  XNOR2_X1 U401 ( .A(G15GAT), .B(G1GAT), .ZN(n340) );
  XNOR2_X1 U402 ( .A(n340), .B(KEYINPUT69), .ZN(n419) );
  XOR2_X1 U403 ( .A(n419), .B(KEYINPUT79), .Z(n342) );
  NAND2_X1 U404 ( .A1(G231GAT), .A2(G233GAT), .ZN(n341) );
  XNOR2_X1 U405 ( .A(n342), .B(n341), .ZN(n343) );
  XOR2_X1 U406 ( .A(n344), .B(n343), .Z(n352) );
  XOR2_X1 U407 ( .A(KEYINPUT80), .B(KEYINPUT14), .Z(n346) );
  XNOR2_X1 U408 ( .A(G127GAT), .B(KEYINPUT15), .ZN(n345) );
  XNOR2_X1 U409 ( .A(n346), .B(n345), .ZN(n350) );
  XOR2_X1 U410 ( .A(G64GAT), .B(KEYINPUT12), .Z(n348) );
  XNOR2_X1 U411 ( .A(G8GAT), .B(KEYINPUT81), .ZN(n347) );
  XNOR2_X1 U412 ( .A(n348), .B(n347), .ZN(n349) );
  XNOR2_X1 U413 ( .A(n350), .B(n349), .ZN(n351) );
  XNOR2_X1 U414 ( .A(n352), .B(n351), .ZN(n540) );
  XOR2_X1 U415 ( .A(KEYINPUT17), .B(G190GAT), .Z(n354) );
  XNOR2_X1 U416 ( .A(KEYINPUT18), .B(G183GAT), .ZN(n353) );
  XNOR2_X1 U417 ( .A(n354), .B(n353), .ZN(n355) );
  XOR2_X1 U418 ( .A(KEYINPUT19), .B(n355), .Z(n382) );
  XOR2_X1 U419 ( .A(G64GAT), .B(G92GAT), .Z(n357) );
  XNOR2_X1 U420 ( .A(G176GAT), .B(G204GAT), .ZN(n356) );
  XNOR2_X1 U421 ( .A(n357), .B(n356), .ZN(n439) );
  XNOR2_X1 U422 ( .A(n358), .B(n439), .ZN(n365) );
  XOR2_X1 U423 ( .A(G169GAT), .B(G8GAT), .Z(n420) );
  XOR2_X1 U424 ( .A(KEYINPUT94), .B(KEYINPUT93), .Z(n360) );
  XNOR2_X1 U425 ( .A(G36GAT), .B(KEYINPUT79), .ZN(n359) );
  XNOR2_X1 U426 ( .A(n360), .B(n359), .ZN(n361) );
  XOR2_X1 U427 ( .A(n420), .B(n361), .Z(n363) );
  NAND2_X1 U428 ( .A1(G226GAT), .A2(G233GAT), .ZN(n362) );
  XNOR2_X1 U429 ( .A(n363), .B(n362), .ZN(n364) );
  XNOR2_X1 U430 ( .A(n365), .B(n364), .ZN(n366) );
  XNOR2_X1 U431 ( .A(n382), .B(n366), .ZN(n496) );
  XOR2_X1 U432 ( .A(KEYINPUT27), .B(KEYINPUT95), .Z(n367) );
  XNOR2_X1 U433 ( .A(n496), .B(n367), .ZN(n529) );
  XOR2_X1 U434 ( .A(KEYINPUT83), .B(KEYINPUT84), .Z(n369) );
  XNOR2_X1 U435 ( .A(G169GAT), .B(G15GAT), .ZN(n368) );
  XNOR2_X1 U436 ( .A(n369), .B(n368), .ZN(n380) );
  XOR2_X1 U437 ( .A(G120GAT), .B(G71GAT), .Z(n435) );
  XNOR2_X1 U438 ( .A(G43GAT), .B(G99GAT), .ZN(n370) );
  XNOR2_X1 U439 ( .A(n294), .B(n370), .ZN(n371) );
  NAND2_X1 U440 ( .A1(G227GAT), .A2(G233GAT), .ZN(n372) );
  XNOR2_X1 U441 ( .A(n295), .B(n372), .ZN(n378) );
  XOR2_X1 U442 ( .A(G127GAT), .B(KEYINPUT0), .Z(n374) );
  XNOR2_X1 U443 ( .A(G113GAT), .B(G134GAT), .ZN(n373) );
  XNOR2_X1 U444 ( .A(n374), .B(n373), .ZN(n407) );
  XNOR2_X1 U445 ( .A(n407), .B(KEYINPUT20), .ZN(n376) );
  XOR2_X1 U446 ( .A(n380), .B(n379), .Z(n381) );
  NOR2_X1 U447 ( .A1(n521), .A2(n473), .ZN(n383) );
  XOR2_X1 U448 ( .A(KEYINPUT26), .B(n383), .Z(n547) );
  NOR2_X1 U449 ( .A1(n529), .A2(n547), .ZN(n384) );
  XNOR2_X1 U450 ( .A(n384), .B(KEYINPUT97), .ZN(n390) );
  INV_X1 U451 ( .A(n521), .ZN(n536) );
  NOR2_X1 U452 ( .A1(n536), .A2(n496), .ZN(n386) );
  XNOR2_X1 U453 ( .A(n386), .B(n385), .ZN(n387) );
  XNOR2_X1 U454 ( .A(KEYINPUT25), .B(n388), .ZN(n389) );
  NAND2_X1 U455 ( .A1(n390), .A2(n389), .ZN(n410) );
  XOR2_X1 U456 ( .A(G85GAT), .B(G162GAT), .Z(n392) );
  XNOR2_X1 U457 ( .A(G29GAT), .B(G141GAT), .ZN(n391) );
  XNOR2_X1 U458 ( .A(n392), .B(n391), .ZN(n396) );
  XOR2_X1 U459 ( .A(G57GAT), .B(G148GAT), .Z(n394) );
  XNOR2_X1 U460 ( .A(G1GAT), .B(G120GAT), .ZN(n393) );
  XNOR2_X1 U461 ( .A(n394), .B(n393), .ZN(n395) );
  XOR2_X1 U462 ( .A(n396), .B(n395), .Z(n401) );
  XOR2_X1 U463 ( .A(KEYINPUT4), .B(KEYINPUT5), .Z(n398) );
  NAND2_X1 U464 ( .A1(G225GAT), .A2(G233GAT), .ZN(n397) );
  XNOR2_X1 U465 ( .A(n398), .B(n397), .ZN(n399) );
  XNOR2_X1 U466 ( .A(KEYINPUT90), .B(n399), .ZN(n400) );
  XNOR2_X1 U467 ( .A(n401), .B(n400), .ZN(n405) );
  XOR2_X1 U468 ( .A(KEYINPUT91), .B(KEYINPUT92), .Z(n403) );
  XNOR2_X1 U469 ( .A(KEYINPUT6), .B(KEYINPUT1), .ZN(n402) );
  XNOR2_X1 U470 ( .A(n403), .B(n402), .ZN(n404) );
  XOR2_X1 U471 ( .A(n405), .B(n404), .Z(n409) );
  XNOR2_X1 U472 ( .A(n407), .B(n406), .ZN(n408) );
  XNOR2_X1 U473 ( .A(n409), .B(n408), .ZN(n493) );
  NAND2_X1 U474 ( .A1(n410), .A2(n493), .ZN(n415) );
  INV_X1 U475 ( .A(n493), .ZN(n532) );
  NAND2_X1 U476 ( .A1(n536), .A2(n534), .ZN(n411) );
  NOR2_X1 U477 ( .A1(n529), .A2(n411), .ZN(n412) );
  NAND2_X1 U478 ( .A1(n532), .A2(n412), .ZN(n413) );
  XNOR2_X1 U479 ( .A(n413), .B(KEYINPUT96), .ZN(n414) );
  NAND2_X1 U480 ( .A1(n540), .A2(n481), .ZN(n416) );
  XOR2_X1 U481 ( .A(KEYINPUT103), .B(n416), .Z(n417) );
  XNOR2_X1 U482 ( .A(KEYINPUT37), .B(n418), .ZN(n515) );
  XOR2_X1 U483 ( .A(n420), .B(n419), .Z(n422) );
  XNOR2_X1 U484 ( .A(G197GAT), .B(G113GAT), .ZN(n421) );
  XNOR2_X1 U485 ( .A(n422), .B(n421), .ZN(n427) );
  XOR2_X1 U486 ( .A(n423), .B(KEYINPUT70), .Z(n425) );
  NAND2_X1 U487 ( .A1(G229GAT), .A2(G233GAT), .ZN(n424) );
  XNOR2_X1 U488 ( .A(n425), .B(n424), .ZN(n426) );
  XOR2_X1 U489 ( .A(n427), .B(n426), .Z(n433) );
  XOR2_X1 U490 ( .A(KEYINPUT68), .B(KEYINPUT29), .Z(n429) );
  XNOR2_X1 U491 ( .A(KEYINPUT67), .B(KEYINPUT30), .ZN(n428) );
  XNOR2_X1 U492 ( .A(n429), .B(n428), .ZN(n430) );
  XNOR2_X1 U493 ( .A(n431), .B(n430), .ZN(n432) );
  XNOR2_X1 U494 ( .A(n433), .B(n432), .ZN(n577) );
  XOR2_X1 U495 ( .A(KEYINPUT71), .B(n577), .Z(n564) );
  XNOR2_X1 U496 ( .A(n435), .B(n434), .ZN(n448) );
  XOR2_X1 U497 ( .A(KEYINPUT31), .B(KEYINPUT33), .Z(n437) );
  NAND2_X1 U498 ( .A1(G230GAT), .A2(G233GAT), .ZN(n436) );
  XNOR2_X1 U499 ( .A(n437), .B(n436), .ZN(n438) );
  XOR2_X1 U500 ( .A(n438), .B(KEYINPUT73), .Z(n442) );
  XNOR2_X1 U501 ( .A(n440), .B(n439), .ZN(n441) );
  XNOR2_X1 U502 ( .A(n442), .B(n441), .ZN(n443) );
  XOR2_X1 U503 ( .A(n443), .B(KEYINPUT32), .Z(n446) );
  XNOR2_X1 U504 ( .A(n444), .B(KEYINPUT74), .ZN(n445) );
  XNOR2_X1 U505 ( .A(n446), .B(n445), .ZN(n447) );
  XNOR2_X1 U506 ( .A(n448), .B(n447), .ZN(n581) );
  NAND2_X1 U507 ( .A1(n564), .A2(n581), .ZN(n484) );
  NOR2_X1 U508 ( .A1(n515), .A2(n484), .ZN(n449) );
  XNOR2_X1 U509 ( .A(n450), .B(n449), .ZN(n451) );
  NOR2_X1 U510 ( .A1(n534), .A2(n501), .ZN(n453) );
  NOR2_X1 U511 ( .A1(n540), .A2(n589), .ZN(n454) );
  XNOR2_X1 U512 ( .A(n454), .B(KEYINPUT45), .ZN(n457) );
  INV_X1 U513 ( .A(n581), .ZN(n455) );
  NOR2_X1 U514 ( .A1(n564), .A2(n455), .ZN(n456) );
  AND2_X1 U515 ( .A1(n457), .A2(n456), .ZN(n458) );
  XNOR2_X1 U516 ( .A(n458), .B(KEYINPUT117), .ZN(n466) );
  XNOR2_X1 U517 ( .A(n581), .B(KEYINPUT41), .ZN(n555) );
  NAND2_X1 U518 ( .A1(n555), .A2(n577), .ZN(n460) );
  XOR2_X1 U519 ( .A(KEYINPUT115), .B(KEYINPUT46), .Z(n459) );
  XNOR2_X1 U520 ( .A(n460), .B(n459), .ZN(n461) );
  NAND2_X1 U521 ( .A1(n461), .A2(n540), .ZN(n462) );
  NOR2_X1 U522 ( .A1(n561), .A2(n462), .ZN(n464) );
  XNOR2_X1 U523 ( .A(KEYINPUT116), .B(KEYINPUT47), .ZN(n463) );
  XNOR2_X1 U524 ( .A(n464), .B(n463), .ZN(n465) );
  NAND2_X1 U525 ( .A1(n466), .A2(n465), .ZN(n469) );
  NOR2_X1 U526 ( .A1(n530), .A2(n496), .ZN(n470) );
  XNOR2_X1 U527 ( .A(n470), .B(KEYINPUT54), .ZN(n471) );
  NAND2_X1 U528 ( .A1(n471), .A2(n493), .ZN(n472) );
  XNOR2_X1 U529 ( .A(n472), .B(KEYINPUT65), .ZN(n575) );
  NAND2_X1 U530 ( .A1(n575), .A2(n473), .ZN(n474) );
  XNOR2_X1 U531 ( .A(n474), .B(KEYINPUT55), .ZN(n475) );
  AND2_X1 U532 ( .A1(n475), .A2(n521), .ZN(n573) );
  NAND2_X1 U533 ( .A1(n573), .A2(n561), .ZN(n477) );
  XNOR2_X1 U534 ( .A(G1GAT), .B(KEYINPUT100), .ZN(n478) );
  XNOR2_X1 U535 ( .A(n478), .B(KEYINPUT101), .ZN(n479) );
  XOR2_X1 U536 ( .A(KEYINPUT34), .B(n479), .Z(n486) );
  NOR2_X1 U537 ( .A1(n561), .A2(n540), .ZN(n480) );
  XNOR2_X1 U538 ( .A(n480), .B(KEYINPUT16), .ZN(n482) );
  NAND2_X1 U539 ( .A1(n482), .A2(n481), .ZN(n483) );
  XOR2_X1 U540 ( .A(KEYINPUT99), .B(n483), .Z(n504) );
  NOR2_X1 U541 ( .A1(n484), .A2(n504), .ZN(n491) );
  NAND2_X1 U542 ( .A1(n491), .A2(n532), .ZN(n485) );
  XNOR2_X1 U543 ( .A(n486), .B(n485), .ZN(G1324GAT) );
  INV_X1 U544 ( .A(n496), .ZN(n518) );
  NAND2_X1 U545 ( .A1(n491), .A2(n518), .ZN(n487) );
  XNOR2_X1 U546 ( .A(n487), .B(G8GAT), .ZN(G1325GAT) );
  XOR2_X1 U547 ( .A(KEYINPUT35), .B(KEYINPUT102), .Z(n489) );
  NAND2_X1 U548 ( .A1(n491), .A2(n521), .ZN(n488) );
  XNOR2_X1 U549 ( .A(n489), .B(n488), .ZN(n490) );
  XNOR2_X1 U550 ( .A(G15GAT), .B(n490), .ZN(G1326GAT) );
  INV_X1 U551 ( .A(n534), .ZN(n524) );
  NAND2_X1 U552 ( .A1(n491), .A2(n524), .ZN(n492) );
  XNOR2_X1 U553 ( .A(n492), .B(G22GAT), .ZN(G1327GAT) );
  NOR2_X1 U554 ( .A1(n493), .A2(n501), .ZN(n495) );
  XNOR2_X1 U555 ( .A(G29GAT), .B(KEYINPUT39), .ZN(n494) );
  XNOR2_X1 U556 ( .A(n495), .B(n494), .ZN(G1328GAT) );
  NOR2_X1 U557 ( .A1(n496), .A2(n501), .ZN(n498) );
  XNOR2_X1 U558 ( .A(G36GAT), .B(KEYINPUT105), .ZN(n497) );
  XNOR2_X1 U559 ( .A(n498), .B(n497), .ZN(G1329GAT) );
  XOR2_X1 U560 ( .A(KEYINPUT107), .B(KEYINPUT40), .Z(n500) );
  XNOR2_X1 U561 ( .A(G43GAT), .B(KEYINPUT106), .ZN(n499) );
  XNOR2_X1 U562 ( .A(n500), .B(n499), .ZN(n503) );
  NOR2_X1 U563 ( .A1(n536), .A2(n501), .ZN(n502) );
  XOR2_X1 U564 ( .A(n503), .B(n502), .Z(G1330GAT) );
  XOR2_X1 U565 ( .A(KEYINPUT42), .B(KEYINPUT110), .Z(n507) );
  XNOR2_X1 U566 ( .A(KEYINPUT108), .B(n555), .ZN(n570) );
  INV_X1 U567 ( .A(n577), .ZN(n549) );
  NAND2_X1 U568 ( .A1(n570), .A2(n549), .ZN(n514) );
  NOR2_X1 U569 ( .A1(n514), .A2(n504), .ZN(n505) );
  XOR2_X1 U570 ( .A(KEYINPUT109), .B(n505), .Z(n511) );
  NAND2_X1 U571 ( .A1(n511), .A2(n532), .ZN(n506) );
  XNOR2_X1 U572 ( .A(n507), .B(n506), .ZN(n508) );
  XOR2_X1 U573 ( .A(G57GAT), .B(n508), .Z(G1332GAT) );
  NAND2_X1 U574 ( .A1(n511), .A2(n518), .ZN(n509) );
  XNOR2_X1 U575 ( .A(n509), .B(G64GAT), .ZN(G1333GAT) );
  NAND2_X1 U576 ( .A1(n521), .A2(n511), .ZN(n510) );
  XNOR2_X1 U577 ( .A(n510), .B(G71GAT), .ZN(G1334GAT) );
  XOR2_X1 U578 ( .A(G78GAT), .B(KEYINPUT43), .Z(n513) );
  NAND2_X1 U579 ( .A1(n511), .A2(n524), .ZN(n512) );
  XNOR2_X1 U580 ( .A(n513), .B(n512), .ZN(G1335GAT) );
  XOR2_X1 U581 ( .A(G85GAT), .B(KEYINPUT111), .Z(n517) );
  NOR2_X1 U582 ( .A1(n515), .A2(n514), .ZN(n525) );
  NAND2_X1 U583 ( .A1(n525), .A2(n532), .ZN(n516) );
  XNOR2_X1 U584 ( .A(n517), .B(n516), .ZN(G1336GAT) );
  XNOR2_X1 U585 ( .A(G92GAT), .B(KEYINPUT112), .ZN(n520) );
  NAND2_X1 U586 ( .A1(n518), .A2(n525), .ZN(n519) );
  XNOR2_X1 U587 ( .A(n520), .B(n519), .ZN(G1337GAT) );
  XOR2_X1 U588 ( .A(G99GAT), .B(KEYINPUT113), .Z(n523) );
  NAND2_X1 U589 ( .A1(n525), .A2(n521), .ZN(n522) );
  XNOR2_X1 U590 ( .A(n523), .B(n522), .ZN(G1338GAT) );
  XOR2_X1 U591 ( .A(KEYINPUT44), .B(KEYINPUT114), .Z(n527) );
  NAND2_X1 U592 ( .A1(n525), .A2(n524), .ZN(n526) );
  XNOR2_X1 U593 ( .A(n527), .B(n526), .ZN(n528) );
  XOR2_X1 U594 ( .A(G106GAT), .B(n528), .Z(G1339GAT) );
  NOR2_X1 U595 ( .A1(n530), .A2(n529), .ZN(n531) );
  NAND2_X1 U596 ( .A1(n532), .A2(n531), .ZN(n533) );
  XOR2_X1 U597 ( .A(KEYINPUT118), .B(n533), .Z(n548) );
  NAND2_X1 U598 ( .A1(n534), .A2(n548), .ZN(n535) );
  NOR2_X1 U599 ( .A1(n536), .A2(n535), .ZN(n543) );
  NAND2_X1 U600 ( .A1(n543), .A2(n564), .ZN(n537) );
  XNOR2_X1 U601 ( .A(n537), .B(G113GAT), .ZN(G1340GAT) );
  XOR2_X1 U602 ( .A(G120GAT), .B(KEYINPUT49), .Z(n539) );
  NAND2_X1 U603 ( .A1(n543), .A2(n570), .ZN(n538) );
  XNOR2_X1 U604 ( .A(n539), .B(n538), .ZN(G1341GAT) );
  INV_X1 U605 ( .A(n540), .ZN(n584) );
  NAND2_X1 U606 ( .A1(n584), .A2(n543), .ZN(n541) );
  XNOR2_X1 U607 ( .A(n541), .B(KEYINPUT50), .ZN(n542) );
  XNOR2_X1 U608 ( .A(G127GAT), .B(n542), .ZN(G1342GAT) );
  XOR2_X1 U609 ( .A(KEYINPUT119), .B(KEYINPUT51), .Z(n545) );
  NAND2_X1 U610 ( .A1(n543), .A2(n561), .ZN(n544) );
  XNOR2_X1 U611 ( .A(n545), .B(n544), .ZN(n546) );
  XOR2_X1 U612 ( .A(G134GAT), .B(n546), .Z(G1343GAT) );
  INV_X1 U613 ( .A(n547), .ZN(n576) );
  NAND2_X1 U614 ( .A1(n576), .A2(n548), .ZN(n554) );
  NOR2_X1 U615 ( .A1(n549), .A2(n554), .ZN(n550) );
  XOR2_X1 U616 ( .A(G141GAT), .B(n550), .Z(n551) );
  XNOR2_X1 U617 ( .A(KEYINPUT120), .B(n551), .ZN(G1344GAT) );
  XOR2_X1 U618 ( .A(KEYINPUT123), .B(KEYINPUT53), .Z(n553) );
  XNOR2_X1 U619 ( .A(KEYINPUT121), .B(KEYINPUT122), .ZN(n552) );
  XNOR2_X1 U620 ( .A(n553), .B(n552), .ZN(n559) );
  XOR2_X1 U621 ( .A(G148GAT), .B(KEYINPUT52), .Z(n557) );
  INV_X1 U622 ( .A(n554), .ZN(n562) );
  NAND2_X1 U623 ( .A1(n562), .A2(n555), .ZN(n556) );
  XNOR2_X1 U624 ( .A(n557), .B(n556), .ZN(n558) );
  XOR2_X1 U625 ( .A(n559), .B(n558), .Z(G1345GAT) );
  NAND2_X1 U626 ( .A1(n584), .A2(n562), .ZN(n560) );
  XNOR2_X1 U627 ( .A(n560), .B(G155GAT), .ZN(G1346GAT) );
  NAND2_X1 U628 ( .A1(n562), .A2(n561), .ZN(n563) );
  XNOR2_X1 U629 ( .A(n563), .B(G162GAT), .ZN(G1347GAT) );
  NAND2_X1 U630 ( .A1(n573), .A2(n564), .ZN(n565) );
  XNOR2_X1 U631 ( .A(n565), .B(KEYINPUT124), .ZN(n566) );
  XNOR2_X1 U632 ( .A(G169GAT), .B(n566), .ZN(G1348GAT) );
  XOR2_X1 U633 ( .A(KEYINPUT57), .B(KEYINPUT126), .Z(n568) );
  XNOR2_X1 U634 ( .A(G176GAT), .B(KEYINPUT125), .ZN(n567) );
  XNOR2_X1 U635 ( .A(n568), .B(n567), .ZN(n569) );
  XOR2_X1 U636 ( .A(KEYINPUT56), .B(n569), .Z(n572) );
  NAND2_X1 U637 ( .A1(n570), .A2(n573), .ZN(n571) );
  XNOR2_X1 U638 ( .A(n572), .B(n571), .ZN(G1349GAT) );
  NAND2_X1 U639 ( .A1(n584), .A2(n573), .ZN(n574) );
  XNOR2_X1 U640 ( .A(n574), .B(G183GAT), .ZN(G1350GAT) );
  XOR2_X1 U641 ( .A(KEYINPUT60), .B(KEYINPUT59), .Z(n579) );
  NAND2_X1 U642 ( .A1(n576), .A2(n575), .ZN(n588) );
  INV_X1 U643 ( .A(n588), .ZN(n585) );
  NAND2_X1 U644 ( .A1(n585), .A2(n577), .ZN(n578) );
  XNOR2_X1 U645 ( .A(n579), .B(n578), .ZN(n580) );
  XNOR2_X1 U646 ( .A(G197GAT), .B(n580), .ZN(G1352GAT) );
  XOR2_X1 U647 ( .A(G204GAT), .B(KEYINPUT61), .Z(n583) );
  OR2_X1 U648 ( .A1(n588), .A2(n581), .ZN(n582) );
  XNOR2_X1 U649 ( .A(n583), .B(n582), .ZN(G1353GAT) );
  XOR2_X1 U650 ( .A(G211GAT), .B(KEYINPUT127), .Z(n587) );
  NAND2_X1 U651 ( .A1(n585), .A2(n584), .ZN(n586) );
  XNOR2_X1 U652 ( .A(n587), .B(n586), .ZN(G1354GAT) );
  NOR2_X1 U653 ( .A1(n589), .A2(n588), .ZN(n590) );
  XOR2_X1 U654 ( .A(KEYINPUT62), .B(n590), .Z(n591) );
  XNOR2_X1 U655 ( .A(G218GAT), .B(n591), .ZN(G1355GAT) );
endmodule

