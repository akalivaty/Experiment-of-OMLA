//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 1 1 0 0 1 0 0 1 0 1 1 1 0 0 0 0 0 0 0 0 1 1 0 0 1 0 0 0 1 0 1 0 0 0 0 0 1 0 1 1 0 0 1 1 1 1 1 0 1 0 1 0 0 1 1 1 1 1 0 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:20:15 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n696, new_n697, new_n698, new_n699,
    new_n700, new_n701, new_n703, new_n704, new_n705, new_n706, new_n707,
    new_n708, new_n710, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n743, new_n744, new_n745,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n762,
    new_n763, new_n764, new_n765, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n773, new_n774, new_n775, new_n777, new_n779, new_n780,
    new_n781, new_n782, new_n783, new_n784, new_n785, new_n786, new_n787,
    new_n788, new_n789, new_n790, new_n791, new_n792, new_n793, new_n794,
    new_n795, new_n796, new_n797, new_n798, new_n799, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n812, new_n813, new_n814, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n863, new_n864, new_n865, new_n867, new_n868, new_n870, new_n871,
    new_n872, new_n873, new_n874, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n915, new_n916, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n930, new_n931, new_n932, new_n934,
    new_n935, new_n936, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n952, new_n953, new_n954, new_n955, new_n956, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n970, new_n971, new_n972, new_n973,
    new_n974, new_n975, new_n976, new_n977, new_n978, new_n980, new_n981;
  INV_X1    g000(.A(G22gat), .ZN(new_n202));
  INV_X1    g001(.A(KEYINPUT81), .ZN(new_n203));
  XNOR2_X1  g002(.A(G197gat), .B(G204gat), .ZN(new_n204));
  NAND2_X1  g003(.A1(G211gat), .A2(G218gat), .ZN(new_n205));
  INV_X1    g004(.A(KEYINPUT22), .ZN(new_n206));
  NAND2_X1  g005(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  NAND2_X1  g006(.A1(new_n204), .A2(new_n207), .ZN(new_n208));
  XNOR2_X1  g007(.A(G211gat), .B(G218gat), .ZN(new_n209));
  INV_X1    g008(.A(new_n209), .ZN(new_n210));
  NAND2_X1  g009(.A1(new_n208), .A2(new_n210), .ZN(new_n211));
  NAND3_X1  g010(.A1(new_n209), .A2(new_n204), .A3(new_n207), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  INV_X1    g012(.A(KEYINPUT29), .ZN(new_n214));
  AOI21_X1  g013(.A(KEYINPUT3), .B1(new_n213), .B2(new_n214), .ZN(new_n215));
  INV_X1    g014(.A(G148gat), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n216), .A2(KEYINPUT74), .ZN(new_n217));
  INV_X1    g016(.A(KEYINPUT74), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n218), .A2(G148gat), .ZN(new_n219));
  NAND3_X1  g018(.A1(new_n217), .A2(new_n219), .A3(G141gat), .ZN(new_n220));
  INV_X1    g019(.A(G141gat), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n221), .A2(G148gat), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n222), .A2(KEYINPUT75), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n220), .A2(new_n223), .ZN(new_n224));
  XNOR2_X1  g023(.A(KEYINPUT74), .B(G148gat), .ZN(new_n225));
  NAND3_X1  g024(.A1(new_n225), .A2(KEYINPUT75), .A3(G141gat), .ZN(new_n226));
  NAND2_X1  g025(.A1(G155gat), .A2(G162gat), .ZN(new_n227));
  NOR2_X1   g026(.A1(G155gat), .A2(G162gat), .ZN(new_n228));
  INV_X1    g027(.A(KEYINPUT2), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  AOI22_X1  g029(.A1(new_n224), .A2(new_n226), .B1(new_n227), .B2(new_n230), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n216), .A2(G141gat), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n222), .A2(new_n232), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n233), .A2(new_n229), .ZN(new_n234));
  INV_X1    g033(.A(new_n228), .ZN(new_n235));
  AND3_X1   g034(.A1(new_n234), .A2(new_n227), .A3(new_n235), .ZN(new_n236));
  NOR2_X1   g035(.A1(new_n231), .A2(new_n236), .ZN(new_n237));
  OAI21_X1  g036(.A(new_n203), .B1(new_n215), .B2(new_n237), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n230), .A2(new_n227), .ZN(new_n239));
  AOI22_X1  g038(.A1(new_n225), .A2(G141gat), .B1(KEYINPUT75), .B2(new_n222), .ZN(new_n240));
  AND4_X1   g039(.A1(KEYINPUT75), .A2(new_n217), .A3(new_n219), .A4(G141gat), .ZN(new_n241));
  OAI21_X1  g040(.A(new_n239), .B1(new_n240), .B2(new_n241), .ZN(new_n242));
  NAND3_X1  g041(.A1(new_n234), .A2(new_n227), .A3(new_n235), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n242), .A2(new_n243), .ZN(new_n244));
  AOI21_X1  g043(.A(KEYINPUT29), .B1(new_n211), .B2(new_n212), .ZN(new_n245));
  OAI211_X1 g044(.A(new_n244), .B(KEYINPUT81), .C1(KEYINPUT3), .C2(new_n245), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n238), .A2(new_n246), .ZN(new_n247));
  INV_X1    g046(.A(KEYINPUT3), .ZN(new_n248));
  NAND3_X1  g047(.A1(new_n242), .A2(new_n248), .A3(new_n243), .ZN(new_n249));
  AOI21_X1  g048(.A(new_n213), .B1(new_n249), .B2(new_n214), .ZN(new_n250));
  INV_X1    g049(.A(new_n250), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n247), .A2(new_n251), .ZN(new_n252));
  NAND2_X1  g051(.A1(G228gat), .A2(G233gat), .ZN(new_n253));
  XOR2_X1   g052(.A(new_n253), .B(KEYINPUT80), .Z(new_n254));
  NAND2_X1  g053(.A1(new_n252), .A2(new_n254), .ZN(new_n255));
  NOR2_X1   g054(.A1(new_n215), .A2(new_n237), .ZN(new_n256));
  NOR3_X1   g055(.A1(new_n250), .A2(new_n256), .A3(new_n253), .ZN(new_n257));
  INV_X1    g056(.A(new_n257), .ZN(new_n258));
  AOI21_X1  g057(.A(new_n202), .B1(new_n255), .B2(new_n258), .ZN(new_n259));
  INV_X1    g058(.A(new_n254), .ZN(new_n260));
  AOI21_X1  g059(.A(new_n260), .B1(new_n247), .B2(new_n251), .ZN(new_n261));
  NOR3_X1   g060(.A1(new_n261), .A2(G22gat), .A3(new_n257), .ZN(new_n262));
  OAI21_X1  g061(.A(KEYINPUT82), .B1(new_n259), .B2(new_n262), .ZN(new_n263));
  XNOR2_X1  g062(.A(G78gat), .B(G106gat), .ZN(new_n264));
  INV_X1    g063(.A(G50gat), .ZN(new_n265));
  XNOR2_X1  g064(.A(new_n264), .B(new_n265), .ZN(new_n266));
  XOR2_X1   g065(.A(KEYINPUT79), .B(KEYINPUT31), .Z(new_n267));
  XNOR2_X1  g066(.A(new_n266), .B(new_n267), .ZN(new_n268));
  INV_X1    g067(.A(new_n268), .ZN(new_n269));
  NAND3_X1  g068(.A1(new_n255), .A2(new_n202), .A3(new_n258), .ZN(new_n270));
  INV_X1    g069(.A(KEYINPUT82), .ZN(new_n271));
  OAI21_X1  g070(.A(G22gat), .B1(new_n261), .B2(new_n257), .ZN(new_n272));
  NAND3_X1  g071(.A1(new_n270), .A2(new_n271), .A3(new_n272), .ZN(new_n273));
  NAND3_X1  g072(.A1(new_n263), .A2(new_n269), .A3(new_n273), .ZN(new_n274));
  NAND4_X1  g073(.A1(new_n270), .A2(new_n272), .A3(new_n271), .A4(new_n268), .ZN(new_n275));
  AND2_X1   g074(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  INV_X1    g075(.A(KEYINPUT25), .ZN(new_n277));
  OR2_X1    g076(.A1(G183gat), .A2(G190gat), .ZN(new_n278));
  NAND3_X1  g077(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n279));
  AOI21_X1  g078(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n280));
  INV_X1    g079(.A(KEYINPUT65), .ZN(new_n281));
  OAI211_X1 g080(.A(new_n278), .B(new_n279), .C1(new_n280), .C2(new_n281), .ZN(new_n282));
  NAND2_X1  g081(.A1(G183gat), .A2(G190gat), .ZN(new_n283));
  INV_X1    g082(.A(KEYINPUT24), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  NOR2_X1   g084(.A1(new_n285), .A2(KEYINPUT65), .ZN(new_n286));
  NOR2_X1   g085(.A1(new_n282), .A2(new_n286), .ZN(new_n287));
  NAND2_X1  g086(.A1(G169gat), .A2(G176gat), .ZN(new_n288));
  NOR2_X1   g087(.A1(G169gat), .A2(G176gat), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n289), .A2(KEYINPUT23), .ZN(new_n290));
  XNOR2_X1  g089(.A(KEYINPUT66), .B(KEYINPUT23), .ZN(new_n291));
  OAI211_X1 g090(.A(new_n288), .B(new_n290), .C1(new_n291), .C2(new_n289), .ZN(new_n292));
  OAI21_X1  g091(.A(new_n277), .B1(new_n287), .B2(new_n292), .ZN(new_n293));
  NAND2_X1  g092(.A1(new_n285), .A2(KEYINPUT68), .ZN(new_n294));
  INV_X1    g093(.A(KEYINPUT68), .ZN(new_n295));
  NAND2_X1  g094(.A1(new_n280), .A2(new_n295), .ZN(new_n296));
  NAND4_X1  g095(.A1(new_n294), .A2(new_n278), .A3(new_n279), .A4(new_n296), .ZN(new_n297));
  OR2_X1    g096(.A1(new_n291), .A2(new_n289), .ZN(new_n298));
  INV_X1    g097(.A(KEYINPUT67), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n289), .A2(new_n299), .ZN(new_n300));
  OAI21_X1  g099(.A(KEYINPUT67), .B1(G169gat), .B2(G176gat), .ZN(new_n301));
  NAND3_X1  g100(.A1(new_n300), .A2(KEYINPUT23), .A3(new_n301), .ZN(new_n302));
  AOI21_X1  g101(.A(new_n277), .B1(G169gat), .B2(G176gat), .ZN(new_n303));
  NAND4_X1  g102(.A1(new_n297), .A2(new_n298), .A3(new_n302), .A4(new_n303), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n293), .A2(new_n304), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n305), .A2(KEYINPUT69), .ZN(new_n306));
  INV_X1    g105(.A(KEYINPUT69), .ZN(new_n307));
  NAND3_X1  g106(.A1(new_n293), .A2(new_n304), .A3(new_n307), .ZN(new_n308));
  XNOR2_X1  g107(.A(KEYINPUT27), .B(G183gat), .ZN(new_n309));
  INV_X1    g108(.A(G190gat), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  INV_X1    g110(.A(KEYINPUT28), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  NAND3_X1  g112(.A1(new_n309), .A2(KEYINPUT28), .A3(new_n310), .ZN(new_n314));
  AOI22_X1  g113(.A1(new_n313), .A2(new_n314), .B1(G183gat), .B2(G190gat), .ZN(new_n315));
  INV_X1    g114(.A(KEYINPUT26), .ZN(new_n316));
  NAND3_X1  g115(.A1(new_n300), .A2(new_n316), .A3(new_n301), .ZN(new_n317));
  INV_X1    g116(.A(KEYINPUT70), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n317), .A2(new_n318), .ZN(new_n319));
  NAND4_X1  g118(.A1(new_n300), .A2(KEYINPUT70), .A3(new_n316), .A4(new_n301), .ZN(new_n320));
  OAI21_X1  g119(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n321));
  NAND4_X1  g120(.A1(new_n319), .A2(new_n288), .A3(new_n320), .A4(new_n321), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n315), .A2(new_n322), .ZN(new_n323));
  NAND3_X1  g122(.A1(new_n306), .A2(new_n308), .A3(new_n323), .ZN(new_n324));
  AND2_X1   g123(.A1(G226gat), .A2(G233gat), .ZN(new_n325));
  NOR2_X1   g124(.A1(new_n325), .A2(KEYINPUT29), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n324), .A2(new_n326), .ZN(new_n327));
  INV_X1    g126(.A(new_n213), .ZN(new_n328));
  AOI22_X1  g127(.A1(new_n322), .A2(new_n315), .B1(new_n293), .B2(new_n304), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n329), .A2(new_n325), .ZN(new_n330));
  NAND3_X1  g129(.A1(new_n327), .A2(new_n328), .A3(new_n330), .ZN(new_n331));
  NAND4_X1  g130(.A1(new_n306), .A2(new_n308), .A3(new_n323), .A4(new_n325), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n323), .A2(new_n305), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n333), .A2(new_n326), .ZN(new_n334));
  NAND2_X1  g133(.A1(new_n332), .A2(new_n334), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n335), .A2(new_n213), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n331), .A2(new_n336), .ZN(new_n337));
  XNOR2_X1  g136(.A(G8gat), .B(G36gat), .ZN(new_n338));
  XNOR2_X1  g137(.A(G64gat), .B(G92gat), .ZN(new_n339));
  XNOR2_X1  g138(.A(new_n338), .B(new_n339), .ZN(new_n340));
  NOR3_X1   g139(.A1(new_n337), .A2(KEYINPUT30), .A3(new_n340), .ZN(new_n341));
  INV_X1    g140(.A(KEYINPUT73), .ZN(new_n342));
  AOI221_X4 g141(.A(new_n213), .B1(new_n325), .B2(new_n329), .C1(new_n324), .C2(new_n326), .ZN(new_n343));
  AOI21_X1  g142(.A(new_n328), .B1(new_n332), .B2(new_n334), .ZN(new_n344));
  OAI21_X1  g143(.A(new_n342), .B1(new_n343), .B2(new_n344), .ZN(new_n345));
  NAND3_X1  g144(.A1(new_n331), .A2(new_n336), .A3(KEYINPUT73), .ZN(new_n346));
  NAND3_X1  g145(.A1(new_n345), .A2(new_n340), .A3(new_n346), .ZN(new_n347));
  INV_X1    g146(.A(KEYINPUT30), .ZN(new_n348));
  AOI22_X1  g147(.A1(new_n324), .A2(new_n326), .B1(new_n325), .B2(new_n329), .ZN(new_n349));
  AOI21_X1  g148(.A(new_n344), .B1(new_n328), .B2(new_n349), .ZN(new_n350));
  INV_X1    g149(.A(new_n340), .ZN(new_n351));
  AOI21_X1  g150(.A(new_n348), .B1(new_n350), .B2(new_n351), .ZN(new_n352));
  AOI21_X1  g151(.A(new_n341), .B1(new_n347), .B2(new_n352), .ZN(new_n353));
  XNOR2_X1  g152(.A(G1gat), .B(G29gat), .ZN(new_n354));
  XNOR2_X1  g153(.A(new_n354), .B(KEYINPUT0), .ZN(new_n355));
  XNOR2_X1  g154(.A(new_n355), .B(KEYINPUT76), .ZN(new_n356));
  XOR2_X1   g155(.A(G57gat), .B(G85gat), .Z(new_n357));
  XNOR2_X1  g156(.A(new_n356), .B(new_n357), .ZN(new_n358));
  OAI21_X1  g157(.A(KEYINPUT3), .B1(new_n231), .B2(new_n236), .ZN(new_n359));
  XOR2_X1   g158(.A(G113gat), .B(G120gat), .Z(new_n360));
  INV_X1    g159(.A(KEYINPUT1), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  XNOR2_X1  g161(.A(G127gat), .B(G134gat), .ZN(new_n363));
  INV_X1    g162(.A(new_n363), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n362), .A2(new_n364), .ZN(new_n365));
  NAND3_X1  g164(.A1(new_n360), .A2(new_n361), .A3(new_n363), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n365), .A2(new_n366), .ZN(new_n367));
  NAND3_X1  g166(.A1(new_n359), .A2(new_n249), .A3(new_n367), .ZN(new_n368));
  INV_X1    g167(.A(KEYINPUT4), .ZN(new_n369));
  OAI21_X1  g168(.A(new_n369), .B1(new_n244), .B2(new_n367), .ZN(new_n370));
  AND2_X1   g169(.A1(new_n365), .A2(new_n366), .ZN(new_n371));
  NAND3_X1  g170(.A1(new_n237), .A2(new_n371), .A3(KEYINPUT4), .ZN(new_n372));
  NAND3_X1  g171(.A1(new_n368), .A2(new_n370), .A3(new_n372), .ZN(new_n373));
  INV_X1    g172(.A(KEYINPUT39), .ZN(new_n374));
  NAND2_X1  g173(.A1(G225gat), .A2(G233gat), .ZN(new_n375));
  INV_X1    g174(.A(new_n375), .ZN(new_n376));
  NAND3_X1  g175(.A1(new_n373), .A2(new_n374), .A3(new_n376), .ZN(new_n377));
  NOR2_X1   g176(.A1(new_n237), .A2(new_n371), .ZN(new_n378));
  NOR2_X1   g177(.A1(new_n244), .A2(new_n367), .ZN(new_n379));
  OR2_X1    g178(.A1(new_n378), .A2(new_n379), .ZN(new_n380));
  OAI21_X1  g179(.A(KEYINPUT39), .B1(new_n380), .B2(new_n376), .ZN(new_n381));
  AND2_X1   g180(.A1(new_n373), .A2(new_n376), .ZN(new_n382));
  OAI211_X1 g181(.A(new_n358), .B(new_n377), .C1(new_n381), .C2(new_n382), .ZN(new_n383));
  NOR2_X1   g182(.A1(KEYINPUT83), .A2(KEYINPUT40), .ZN(new_n384));
  NAND4_X1  g183(.A1(new_n368), .A2(new_n370), .A3(new_n372), .A4(new_n375), .ZN(new_n385));
  INV_X1    g184(.A(KEYINPUT5), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n385), .A2(new_n386), .ZN(new_n387));
  INV_X1    g186(.A(new_n387), .ZN(new_n388));
  OAI21_X1  g187(.A(new_n376), .B1(new_n378), .B2(new_n379), .ZN(new_n389));
  AOI21_X1  g188(.A(new_n386), .B1(new_n385), .B2(new_n389), .ZN(new_n390));
  NOR2_X1   g189(.A1(new_n388), .A2(new_n390), .ZN(new_n391));
  INV_X1    g190(.A(new_n358), .ZN(new_n392));
  AOI22_X1  g191(.A1(new_n383), .A2(new_n384), .B1(new_n391), .B2(new_n392), .ZN(new_n393));
  OR2_X1    g192(.A1(new_n383), .A2(new_n384), .ZN(new_n394));
  NAND3_X1  g193(.A1(new_n353), .A2(new_n393), .A3(new_n394), .ZN(new_n395));
  INV_X1    g194(.A(KEYINPUT6), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n385), .A2(new_n389), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n397), .A2(KEYINPUT5), .ZN(new_n398));
  NAND3_X1  g197(.A1(new_n398), .A2(new_n392), .A3(new_n387), .ZN(new_n399));
  INV_X1    g198(.A(KEYINPUT77), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n398), .A2(new_n387), .ZN(new_n401));
  AOI21_X1  g200(.A(new_n400), .B1(new_n401), .B2(new_n358), .ZN(new_n402));
  OAI211_X1 g201(.A(new_n400), .B(new_n358), .C1(new_n388), .C2(new_n390), .ZN(new_n403));
  INV_X1    g202(.A(new_n403), .ZN(new_n404));
  OAI211_X1 g203(.A(new_n396), .B(new_n399), .C1(new_n402), .C2(new_n404), .ZN(new_n405));
  NAND4_X1  g204(.A1(new_n398), .A2(KEYINPUT6), .A3(new_n392), .A4(new_n387), .ZN(new_n406));
  INV_X1    g205(.A(KEYINPUT84), .ZN(new_n407));
  XNOR2_X1  g206(.A(new_n406), .B(new_n407), .ZN(new_n408));
  INV_X1    g207(.A(KEYINPUT37), .ZN(new_n409));
  AOI21_X1  g208(.A(new_n351), .B1(new_n350), .B2(new_n409), .ZN(new_n410));
  AOI21_X1  g209(.A(new_n409), .B1(new_n349), .B2(new_n213), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n335), .A2(new_n328), .ZN(new_n412));
  AOI21_X1  g211(.A(KEYINPUT38), .B1(new_n411), .B2(new_n412), .ZN(new_n413));
  AOI22_X1  g212(.A1(new_n410), .A2(new_n413), .B1(new_n351), .B2(new_n350), .ZN(new_n414));
  NAND3_X1  g213(.A1(new_n405), .A2(new_n408), .A3(new_n414), .ZN(new_n415));
  INV_X1    g214(.A(KEYINPUT38), .ZN(new_n416));
  NAND3_X1  g215(.A1(new_n345), .A2(KEYINPUT37), .A3(new_n346), .ZN(new_n417));
  AOI21_X1  g216(.A(new_n416), .B1(new_n417), .B2(new_n410), .ZN(new_n418));
  OAI211_X1 g217(.A(new_n276), .B(new_n395), .C1(new_n415), .C2(new_n418), .ZN(new_n419));
  INV_X1    g218(.A(KEYINPUT36), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n308), .A2(new_n323), .ZN(new_n421));
  AOI21_X1  g220(.A(new_n307), .B1(new_n293), .B2(new_n304), .ZN(new_n422));
  OAI21_X1  g221(.A(new_n371), .B1(new_n421), .B2(new_n422), .ZN(new_n423));
  NAND4_X1  g222(.A1(new_n306), .A2(new_n367), .A3(new_n308), .A4(new_n323), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n423), .A2(new_n424), .ZN(new_n425));
  NAND2_X1  g224(.A1(G227gat), .A2(G233gat), .ZN(new_n426));
  XNOR2_X1  g225(.A(new_n426), .B(KEYINPUT64), .ZN(new_n427));
  INV_X1    g226(.A(new_n427), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n425), .A2(new_n428), .ZN(new_n429));
  INV_X1    g228(.A(KEYINPUT71), .ZN(new_n430));
  NAND3_X1  g229(.A1(new_n429), .A2(new_n430), .A3(KEYINPUT34), .ZN(new_n431));
  AOI21_X1  g230(.A(new_n427), .B1(new_n423), .B2(new_n424), .ZN(new_n432));
  INV_X1    g231(.A(KEYINPUT34), .ZN(new_n433));
  OAI21_X1  g232(.A(KEYINPUT71), .B1(new_n432), .B2(new_n433), .ZN(new_n434));
  AND3_X1   g233(.A1(new_n432), .A2(KEYINPUT72), .A3(new_n433), .ZN(new_n435));
  AOI21_X1  g234(.A(KEYINPUT72), .B1(new_n432), .B2(new_n433), .ZN(new_n436));
  OAI211_X1 g235(.A(new_n431), .B(new_n434), .C1(new_n435), .C2(new_n436), .ZN(new_n437));
  NAND3_X1  g236(.A1(new_n423), .A2(new_n427), .A3(new_n424), .ZN(new_n438));
  INV_X1    g237(.A(KEYINPUT33), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n438), .A2(new_n439), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n438), .A2(KEYINPUT32), .ZN(new_n441));
  XOR2_X1   g240(.A(G15gat), .B(G43gat), .Z(new_n442));
  XNOR2_X1  g241(.A(G71gat), .B(G99gat), .ZN(new_n443));
  XNOR2_X1  g242(.A(new_n442), .B(new_n443), .ZN(new_n444));
  NAND3_X1  g243(.A1(new_n440), .A2(new_n441), .A3(new_n444), .ZN(new_n445));
  INV_X1    g244(.A(new_n444), .ZN(new_n446));
  OAI211_X1 g245(.A(new_n438), .B(KEYINPUT32), .C1(new_n439), .C2(new_n446), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n445), .A2(new_n447), .ZN(new_n448));
  AND2_X1   g247(.A1(new_n437), .A2(new_n448), .ZN(new_n449));
  NOR2_X1   g248(.A1(new_n437), .A2(new_n448), .ZN(new_n450));
  OAI21_X1  g249(.A(new_n420), .B1(new_n449), .B2(new_n450), .ZN(new_n451));
  AND2_X1   g250(.A1(new_n431), .A2(new_n434), .ZN(new_n452));
  INV_X1    g251(.A(KEYINPUT72), .ZN(new_n453));
  OAI21_X1  g252(.A(new_n453), .B1(new_n429), .B2(KEYINPUT34), .ZN(new_n454));
  NAND3_X1  g253(.A1(new_n432), .A2(KEYINPUT72), .A3(new_n433), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  NAND4_X1  g255(.A1(new_n452), .A2(new_n456), .A3(new_n447), .A4(new_n445), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n437), .A2(new_n448), .ZN(new_n458));
  NAND3_X1  g257(.A1(new_n457), .A2(new_n458), .A3(KEYINPUT36), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n451), .A2(new_n459), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n274), .A2(new_n275), .ZN(new_n461));
  INV_X1    g260(.A(new_n406), .ZN(new_n462));
  OAI21_X1  g261(.A(KEYINPUT77), .B1(new_n391), .B2(new_n392), .ZN(new_n463));
  AOI21_X1  g262(.A(KEYINPUT6), .B1(new_n463), .B2(new_n403), .ZN(new_n464));
  INV_X1    g263(.A(KEYINPUT78), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n399), .A2(new_n465), .ZN(new_n466));
  NAND3_X1  g265(.A1(new_n391), .A2(KEYINPUT78), .A3(new_n392), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  AOI21_X1  g267(.A(new_n462), .B1(new_n464), .B2(new_n468), .ZN(new_n469));
  OAI21_X1  g268(.A(new_n461), .B1(new_n469), .B2(new_n353), .ZN(new_n470));
  AND3_X1   g269(.A1(new_n419), .A2(new_n460), .A3(new_n470), .ZN(new_n471));
  INV_X1    g270(.A(new_n471), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n405), .A2(new_n408), .ZN(new_n473));
  XNOR2_X1  g272(.A(KEYINPUT86), .B(KEYINPUT35), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n347), .A2(new_n352), .ZN(new_n475));
  INV_X1    g274(.A(new_n341), .ZN(new_n476));
  AOI21_X1  g275(.A(new_n474), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  AND2_X1   g276(.A1(new_n473), .A2(new_n477), .ZN(new_n478));
  AOI21_X1  g277(.A(KEYINPUT85), .B1(new_n457), .B2(new_n458), .ZN(new_n479));
  INV_X1    g278(.A(new_n479), .ZN(new_n480));
  NAND3_X1  g279(.A1(new_n457), .A2(new_n458), .A3(KEYINPUT85), .ZN(new_n481));
  NAND4_X1  g280(.A1(new_n478), .A2(new_n276), .A3(new_n480), .A4(new_n481), .ZN(new_n482));
  NOR2_X1   g281(.A1(new_n449), .A2(new_n450), .ZN(new_n483));
  OAI21_X1  g282(.A(new_n396), .B1(new_n402), .B2(new_n404), .ZN(new_n484));
  AND2_X1   g283(.A1(new_n466), .A2(new_n467), .ZN(new_n485));
  OAI21_X1  g284(.A(new_n406), .B1(new_n484), .B2(new_n485), .ZN(new_n486));
  INV_X1    g285(.A(new_n353), .ZN(new_n487));
  NAND4_X1  g286(.A1(new_n483), .A2(new_n486), .A3(new_n276), .A4(new_n487), .ZN(new_n488));
  NAND2_X1  g287(.A1(new_n488), .A2(KEYINPUT35), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n482), .A2(new_n489), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n472), .A2(new_n490), .ZN(new_n491));
  XNOR2_X1  g290(.A(G127gat), .B(G155gat), .ZN(new_n492));
  XOR2_X1   g291(.A(new_n492), .B(KEYINPUT94), .Z(new_n493));
  AND2_X1   g292(.A1(G71gat), .A2(G78gat), .ZN(new_n494));
  NOR2_X1   g293(.A1(G71gat), .A2(G78gat), .ZN(new_n495));
  NOR2_X1   g294(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  NAND2_X1  g295(.A1(G57gat), .A2(G64gat), .ZN(new_n497));
  INV_X1    g296(.A(new_n497), .ZN(new_n498));
  NOR2_X1   g297(.A1(G57gat), .A2(G64gat), .ZN(new_n499));
  NOR3_X1   g298(.A1(new_n498), .A2(new_n499), .A3(KEYINPUT91), .ZN(new_n500));
  INV_X1    g299(.A(KEYINPUT91), .ZN(new_n501));
  INV_X1    g300(.A(G57gat), .ZN(new_n502));
  INV_X1    g301(.A(G64gat), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  AOI21_X1  g303(.A(new_n501), .B1(new_n504), .B2(new_n497), .ZN(new_n505));
  OAI21_X1  g304(.A(KEYINPUT9), .B1(new_n500), .B2(new_n505), .ZN(new_n506));
  INV_X1    g305(.A(KEYINPUT92), .ZN(new_n507));
  AOI21_X1  g306(.A(new_n494), .B1(KEYINPUT9), .B2(new_n495), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n504), .A2(new_n497), .ZN(new_n509));
  OAI21_X1  g308(.A(new_n507), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  NAND2_X1  g309(.A1(G71gat), .A2(G78gat), .ZN(new_n511));
  INV_X1    g310(.A(G71gat), .ZN(new_n512));
  INV_X1    g311(.A(G78gat), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  INV_X1    g313(.A(KEYINPUT9), .ZN(new_n515));
  OAI21_X1  g314(.A(new_n511), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  NOR2_X1   g315(.A1(new_n498), .A2(new_n499), .ZN(new_n517));
  NAND3_X1  g316(.A1(new_n516), .A2(KEYINPUT92), .A3(new_n517), .ZN(new_n518));
  AOI22_X1  g317(.A1(new_n496), .A2(new_n506), .B1(new_n510), .B2(new_n518), .ZN(new_n519));
  XOR2_X1   g318(.A(KEYINPUT93), .B(KEYINPUT21), .Z(new_n520));
  NOR2_X1   g319(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  NAND2_X1  g320(.A1(G231gat), .A2(G233gat), .ZN(new_n522));
  INV_X1    g321(.A(new_n522), .ZN(new_n523));
  XNOR2_X1  g322(.A(new_n521), .B(new_n523), .ZN(new_n524));
  XOR2_X1   g323(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n525));
  NAND2_X1  g324(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  XNOR2_X1  g325(.A(new_n521), .B(new_n522), .ZN(new_n527));
  INV_X1    g326(.A(new_n525), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  AOI21_X1  g328(.A(new_n493), .B1(new_n526), .B2(new_n529), .ZN(new_n530));
  INV_X1    g329(.A(new_n530), .ZN(new_n531));
  INV_X1    g330(.A(KEYINPUT89), .ZN(new_n532));
  XNOR2_X1  g331(.A(G15gat), .B(G22gat), .ZN(new_n533));
  OR2_X1    g332(.A1(new_n533), .A2(G1gat), .ZN(new_n534));
  INV_X1    g333(.A(KEYINPUT16), .ZN(new_n535));
  OAI21_X1  g334(.A(new_n533), .B1(new_n535), .B2(G1gat), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n534), .A2(new_n536), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n534), .A2(KEYINPUT88), .ZN(new_n538));
  INV_X1    g337(.A(G8gat), .ZN(new_n539));
  NAND3_X1  g338(.A1(new_n537), .A2(new_n538), .A3(new_n539), .ZN(new_n540));
  OAI211_X1 g339(.A(new_n534), .B(new_n536), .C1(KEYINPUT88), .C2(G8gat), .ZN(new_n541));
  AOI21_X1  g340(.A(new_n532), .B1(new_n540), .B2(new_n541), .ZN(new_n542));
  INV_X1    g341(.A(new_n542), .ZN(new_n543));
  NAND3_X1  g342(.A1(new_n540), .A2(new_n532), .A3(new_n541), .ZN(new_n544));
  NAND2_X1  g343(.A1(new_n519), .A2(KEYINPUT21), .ZN(new_n545));
  NAND3_X1  g344(.A1(new_n543), .A2(new_n544), .A3(new_n545), .ZN(new_n546));
  XNOR2_X1  g345(.A(new_n546), .B(KEYINPUT95), .ZN(new_n547));
  NAND3_X1  g346(.A1(new_n526), .A2(new_n529), .A3(new_n493), .ZN(new_n548));
  NAND3_X1  g347(.A1(new_n531), .A2(new_n547), .A3(new_n548), .ZN(new_n549));
  INV_X1    g348(.A(new_n547), .ZN(new_n550));
  INV_X1    g349(.A(new_n548), .ZN(new_n551));
  OAI21_X1  g350(.A(new_n550), .B1(new_n551), .B2(new_n530), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n549), .A2(new_n552), .ZN(new_n553));
  XOR2_X1   g352(.A(G183gat), .B(G211gat), .Z(new_n554));
  NAND2_X1  g353(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  INV_X1    g354(.A(new_n554), .ZN(new_n556));
  NAND3_X1  g355(.A1(new_n549), .A2(new_n552), .A3(new_n556), .ZN(new_n557));
  NAND2_X1  g356(.A1(G232gat), .A2(G233gat), .ZN(new_n558));
  INV_X1    g357(.A(KEYINPUT41), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  XNOR2_X1  g359(.A(new_n560), .B(KEYINPUT96), .ZN(new_n561));
  XNOR2_X1  g360(.A(new_n561), .B(KEYINPUT97), .ZN(new_n562));
  XNOR2_X1  g361(.A(G134gat), .B(G162gat), .ZN(new_n563));
  XNOR2_X1  g362(.A(new_n562), .B(new_n563), .ZN(new_n564));
  NAND2_X1  g363(.A1(G99gat), .A2(G106gat), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n565), .A2(KEYINPUT8), .ZN(new_n566));
  NAND2_X1  g365(.A1(G85gat), .A2(G92gat), .ZN(new_n567));
  INV_X1    g366(.A(KEYINPUT7), .ZN(new_n568));
  NAND2_X1  g367(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  OR2_X1    g368(.A1(G85gat), .A2(G92gat), .ZN(new_n570));
  NAND3_X1  g369(.A1(KEYINPUT7), .A2(G85gat), .A3(G92gat), .ZN(new_n571));
  NAND4_X1  g370(.A1(new_n566), .A2(new_n569), .A3(new_n570), .A4(new_n571), .ZN(new_n572));
  XNOR2_X1  g371(.A(G99gat), .B(G106gat), .ZN(new_n573));
  INV_X1    g372(.A(new_n573), .ZN(new_n574));
  XNOR2_X1  g373(.A(new_n572), .B(new_n574), .ZN(new_n575));
  INV_X1    g374(.A(KEYINPUT14), .ZN(new_n576));
  INV_X1    g375(.A(G29gat), .ZN(new_n577));
  INV_X1    g376(.A(G36gat), .ZN(new_n578));
  NAND3_X1  g377(.A1(new_n576), .A2(new_n577), .A3(new_n578), .ZN(new_n579));
  OAI21_X1  g378(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n580));
  NAND2_X1  g379(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  NAND2_X1  g380(.A1(G29gat), .A2(G36gat), .ZN(new_n582));
  NAND2_X1  g381(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  INV_X1    g382(.A(KEYINPUT15), .ZN(new_n584));
  NAND2_X1  g383(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  XOR2_X1   g384(.A(G43gat), .B(G50gat), .Z(new_n586));
  INV_X1    g385(.A(new_n586), .ZN(new_n587));
  AOI22_X1  g386(.A1(new_n579), .A2(new_n580), .B1(G29gat), .B2(G36gat), .ZN(new_n588));
  NAND2_X1  g387(.A1(new_n588), .A2(KEYINPUT15), .ZN(new_n589));
  NAND3_X1  g388(.A1(new_n585), .A2(new_n587), .A3(new_n589), .ZN(new_n590));
  NAND3_X1  g389(.A1(new_n588), .A2(KEYINPUT15), .A3(new_n586), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  AOI21_X1  g391(.A(KEYINPUT17), .B1(new_n592), .B2(KEYINPUT87), .ZN(new_n593));
  INV_X1    g392(.A(KEYINPUT87), .ZN(new_n594));
  INV_X1    g393(.A(KEYINPUT17), .ZN(new_n595));
  AOI211_X1 g394(.A(new_n594), .B(new_n595), .C1(new_n590), .C2(new_n591), .ZN(new_n596));
  OAI21_X1  g395(.A(new_n575), .B1(new_n593), .B2(new_n596), .ZN(new_n597));
  NOR2_X1   g396(.A1(new_n558), .A2(new_n559), .ZN(new_n598));
  XNOR2_X1  g397(.A(new_n572), .B(new_n573), .ZN(new_n599));
  AOI21_X1  g398(.A(new_n598), .B1(new_n592), .B2(new_n599), .ZN(new_n600));
  XNOR2_X1  g399(.A(G190gat), .B(G218gat), .ZN(new_n601));
  INV_X1    g400(.A(new_n601), .ZN(new_n602));
  NAND3_X1  g401(.A1(new_n597), .A2(new_n600), .A3(new_n602), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n603), .A2(KEYINPUT98), .ZN(new_n604));
  NAND2_X1  g403(.A1(new_n597), .A2(new_n600), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n605), .A2(new_n601), .ZN(new_n606));
  AND2_X1   g405(.A1(new_n604), .A2(new_n606), .ZN(new_n607));
  OR2_X1    g406(.A1(new_n603), .A2(KEYINPUT98), .ZN(new_n608));
  AOI21_X1  g407(.A(new_n564), .B1(new_n607), .B2(new_n608), .ZN(new_n609));
  NAND3_X1  g408(.A1(new_n606), .A2(new_n564), .A3(new_n603), .ZN(new_n610));
  NAND2_X1  g409(.A1(new_n610), .A2(KEYINPUT99), .ZN(new_n611));
  INV_X1    g410(.A(KEYINPUT99), .ZN(new_n612));
  NAND4_X1  g411(.A1(new_n606), .A2(new_n612), .A3(new_n564), .A4(new_n603), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n611), .A2(new_n613), .ZN(new_n614));
  NOR2_X1   g413(.A1(new_n609), .A2(new_n614), .ZN(new_n615));
  NAND3_X1  g414(.A1(new_n555), .A2(new_n557), .A3(new_n615), .ZN(new_n616));
  OAI21_X1  g415(.A(KEYINPUT100), .B1(new_n519), .B2(new_n599), .ZN(new_n617));
  INV_X1    g416(.A(KEYINPUT10), .ZN(new_n618));
  NOR3_X1   g417(.A1(new_n508), .A2(new_n507), .A3(new_n509), .ZN(new_n619));
  AOI21_X1  g418(.A(KEYINPUT92), .B1(new_n516), .B2(new_n517), .ZN(new_n620));
  OAI21_X1  g419(.A(KEYINPUT91), .B1(new_n498), .B2(new_n499), .ZN(new_n621));
  NAND3_X1  g420(.A1(new_n504), .A2(new_n501), .A3(new_n497), .ZN(new_n622));
  AOI21_X1  g421(.A(new_n515), .B1(new_n621), .B2(new_n622), .ZN(new_n623));
  INV_X1    g422(.A(new_n496), .ZN(new_n624));
  OAI22_X1  g423(.A1(new_n619), .A2(new_n620), .B1(new_n623), .B2(new_n624), .ZN(new_n625));
  INV_X1    g424(.A(KEYINPUT100), .ZN(new_n626));
  NAND3_X1  g425(.A1(new_n625), .A2(new_n575), .A3(new_n626), .ZN(new_n627));
  INV_X1    g426(.A(KEYINPUT101), .ZN(new_n628));
  OAI21_X1  g427(.A(new_n628), .B1(new_n572), .B2(new_n574), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n572), .A2(new_n574), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  NAND2_X1  g430(.A1(new_n506), .A2(new_n496), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n510), .A2(new_n518), .ZN(new_n633));
  NAND3_X1  g432(.A1(new_n572), .A2(new_n628), .A3(new_n574), .ZN(new_n634));
  NAND4_X1  g433(.A1(new_n631), .A2(new_n632), .A3(new_n633), .A4(new_n634), .ZN(new_n635));
  NAND4_X1  g434(.A1(new_n617), .A2(new_n618), .A3(new_n627), .A4(new_n635), .ZN(new_n636));
  NAND3_X1  g435(.A1(new_n519), .A2(KEYINPUT10), .A3(new_n599), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  NAND2_X1  g437(.A1(G230gat), .A2(G233gat), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  NAND3_X1  g439(.A1(new_n617), .A2(new_n627), .A3(new_n635), .ZN(new_n641));
  INV_X1    g440(.A(new_n639), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  INV_X1    g442(.A(KEYINPUT102), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  NAND3_X1  g444(.A1(new_n641), .A2(KEYINPUT102), .A3(new_n642), .ZN(new_n646));
  XOR2_X1   g445(.A(G120gat), .B(G148gat), .Z(new_n647));
  XNOR2_X1  g446(.A(new_n647), .B(KEYINPUT103), .ZN(new_n648));
  XOR2_X1   g447(.A(G176gat), .B(G204gat), .Z(new_n649));
  XNOR2_X1  g448(.A(new_n648), .B(new_n649), .ZN(new_n650));
  NAND4_X1  g449(.A1(new_n640), .A2(new_n645), .A3(new_n646), .A4(new_n650), .ZN(new_n651));
  AND2_X1   g450(.A1(new_n645), .A2(new_n646), .ZN(new_n652));
  XOR2_X1   g451(.A(new_n639), .B(KEYINPUT104), .Z(new_n653));
  AOI21_X1  g452(.A(new_n653), .B1(new_n636), .B2(new_n637), .ZN(new_n654));
  INV_X1    g453(.A(new_n654), .ZN(new_n655));
  AND2_X1   g454(.A1(new_n652), .A2(new_n655), .ZN(new_n656));
  OAI21_X1  g455(.A(new_n651), .B1(new_n656), .B2(new_n650), .ZN(new_n657));
  OAI21_X1  g456(.A(KEYINPUT105), .B1(new_n616), .B2(new_n657), .ZN(new_n658));
  AND3_X1   g457(.A1(new_n549), .A2(new_n552), .A3(new_n556), .ZN(new_n659));
  AOI21_X1  g458(.A(new_n556), .B1(new_n549), .B2(new_n552), .ZN(new_n660));
  NOR2_X1   g459(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  INV_X1    g460(.A(KEYINPUT105), .ZN(new_n662));
  INV_X1    g461(.A(new_n657), .ZN(new_n663));
  NAND4_X1  g462(.A1(new_n661), .A2(new_n662), .A3(new_n615), .A4(new_n663), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n540), .A2(new_n541), .ZN(new_n665));
  OAI21_X1  g464(.A(new_n665), .B1(new_n593), .B2(new_n596), .ZN(new_n666));
  INV_X1    g465(.A(new_n544), .ZN(new_n667));
  OAI21_X1  g466(.A(new_n592), .B1(new_n667), .B2(new_n542), .ZN(new_n668));
  NAND2_X1  g467(.A1(G229gat), .A2(G233gat), .ZN(new_n669));
  NAND3_X1  g468(.A1(new_n666), .A2(new_n668), .A3(new_n669), .ZN(new_n670));
  INV_X1    g469(.A(KEYINPUT90), .ZN(new_n671));
  NOR2_X1   g470(.A1(new_n671), .A2(KEYINPUT18), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n670), .A2(new_n672), .ZN(new_n673));
  INV_X1    g472(.A(new_n672), .ZN(new_n674));
  NAND4_X1  g473(.A1(new_n666), .A2(new_n668), .A3(new_n669), .A4(new_n674), .ZN(new_n675));
  INV_X1    g474(.A(new_n592), .ZN(new_n676));
  NAND3_X1  g475(.A1(new_n543), .A2(new_n676), .A3(new_n544), .ZN(new_n677));
  NAND2_X1  g476(.A1(new_n668), .A2(new_n677), .ZN(new_n678));
  XOR2_X1   g477(.A(new_n669), .B(KEYINPUT13), .Z(new_n679));
  NAND2_X1  g478(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  NAND3_X1  g479(.A1(new_n673), .A2(new_n675), .A3(new_n680), .ZN(new_n681));
  XNOR2_X1  g480(.A(G113gat), .B(G141gat), .ZN(new_n682));
  XNOR2_X1  g481(.A(new_n682), .B(KEYINPUT11), .ZN(new_n683));
  INV_X1    g482(.A(G169gat), .ZN(new_n684));
  XNOR2_X1  g483(.A(new_n683), .B(new_n684), .ZN(new_n685));
  XNOR2_X1  g484(.A(new_n685), .B(G197gat), .ZN(new_n686));
  XNOR2_X1  g485(.A(new_n686), .B(KEYINPUT12), .ZN(new_n687));
  INV_X1    g486(.A(new_n687), .ZN(new_n688));
  NAND2_X1  g487(.A1(new_n681), .A2(new_n688), .ZN(new_n689));
  NAND4_X1  g488(.A1(new_n687), .A2(new_n673), .A3(new_n675), .A4(new_n680), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  AND3_X1   g490(.A1(new_n658), .A2(new_n664), .A3(new_n691), .ZN(new_n692));
  AND2_X1   g491(.A1(new_n491), .A2(new_n692), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n693), .A2(new_n469), .ZN(new_n694));
  XNOR2_X1  g493(.A(new_n694), .B(G1gat), .ZN(G1324gat));
  XOR2_X1   g494(.A(KEYINPUT16), .B(G8gat), .Z(new_n696));
  NAND4_X1  g495(.A1(new_n491), .A2(new_n353), .A3(new_n692), .A4(new_n696), .ZN(new_n697));
  OR2_X1    g496(.A1(new_n697), .A2(KEYINPUT42), .ZN(new_n698));
  AOI21_X1  g497(.A(new_n539), .B1(new_n693), .B2(new_n353), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n697), .A2(KEYINPUT42), .ZN(new_n700));
  OAI21_X1  g499(.A(new_n698), .B1(new_n699), .B2(new_n700), .ZN(new_n701));
  XNOR2_X1  g500(.A(new_n701), .B(KEYINPUT106), .ZN(G1325gat));
  INV_X1    g501(.A(G15gat), .ZN(new_n703));
  AND3_X1   g502(.A1(new_n457), .A2(KEYINPUT85), .A3(new_n458), .ZN(new_n704));
  NOR2_X1   g503(.A1(new_n704), .A2(new_n479), .ZN(new_n705));
  NAND3_X1  g504(.A1(new_n693), .A2(new_n703), .A3(new_n705), .ZN(new_n706));
  INV_X1    g505(.A(new_n460), .ZN(new_n707));
  AND2_X1   g506(.A1(new_n693), .A2(new_n707), .ZN(new_n708));
  OAI21_X1  g507(.A(new_n706), .B1(new_n708), .B2(new_n703), .ZN(G1326gat));
  NAND2_X1  g508(.A1(new_n693), .A2(new_n461), .ZN(new_n710));
  OR2_X1    g509(.A1(new_n710), .A2(KEYINPUT107), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n710), .A2(KEYINPUT107), .ZN(new_n712));
  XOR2_X1   g511(.A(KEYINPUT43), .B(G22gat), .Z(new_n713));
  AND3_X1   g512(.A1(new_n711), .A2(new_n712), .A3(new_n713), .ZN(new_n714));
  AOI21_X1  g513(.A(new_n713), .B1(new_n711), .B2(new_n712), .ZN(new_n715));
  NOR2_X1   g514(.A1(new_n714), .A2(new_n715), .ZN(G1327gat));
  AOI21_X1  g515(.A(new_n615), .B1(new_n472), .B2(new_n490), .ZN(new_n717));
  INV_X1    g516(.A(new_n691), .ZN(new_n718));
  NOR3_X1   g517(.A1(new_n661), .A2(new_n718), .A3(new_n657), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n717), .A2(new_n719), .ZN(new_n720));
  NOR3_X1   g519(.A1(new_n720), .A2(G29gat), .A3(new_n486), .ZN(new_n721));
  XOR2_X1   g520(.A(new_n721), .B(KEYINPUT45), .Z(new_n722));
  INV_X1    g521(.A(KEYINPUT108), .ZN(new_n723));
  NAND2_X1  g522(.A1(new_n463), .A2(new_n403), .ZN(new_n724));
  NAND3_X1  g523(.A1(new_n724), .A2(new_n468), .A3(new_n396), .ZN(new_n725));
  AOI21_X1  g524(.A(new_n353), .B1(new_n725), .B2(new_n406), .ZN(new_n726));
  OAI21_X1  g525(.A(new_n723), .B1(new_n726), .B2(new_n276), .ZN(new_n727));
  OAI211_X1 g526(.A(KEYINPUT108), .B(new_n461), .C1(new_n469), .C2(new_n353), .ZN(new_n728));
  NAND4_X1  g527(.A1(new_n727), .A2(new_n419), .A3(new_n460), .A4(new_n728), .ZN(new_n729));
  AOI21_X1  g528(.A(new_n615), .B1(new_n490), .B2(new_n729), .ZN(new_n730));
  OR2_X1    g529(.A1(new_n730), .A2(KEYINPUT44), .ZN(new_n731));
  INV_X1    g530(.A(new_n614), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n607), .A2(new_n608), .ZN(new_n733));
  INV_X1    g532(.A(new_n564), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n732), .A2(new_n735), .ZN(new_n736));
  NOR3_X1   g535(.A1(new_n704), .A2(new_n479), .A3(new_n461), .ZN(new_n737));
  AOI22_X1  g536(.A1(new_n737), .A2(new_n478), .B1(new_n488), .B2(KEYINPUT35), .ZN(new_n738));
  OAI211_X1 g537(.A(KEYINPUT44), .B(new_n736), .C1(new_n738), .C2(new_n471), .ZN(new_n739));
  NAND3_X1  g538(.A1(new_n731), .A2(new_n719), .A3(new_n739), .ZN(new_n740));
  OAI21_X1  g539(.A(G29gat), .B1(new_n740), .B2(new_n486), .ZN(new_n741));
  NAND2_X1  g540(.A1(new_n722), .A2(new_n741), .ZN(G1328gat));
  NOR3_X1   g541(.A1(new_n720), .A2(G36gat), .A3(new_n487), .ZN(new_n743));
  XNOR2_X1  g542(.A(new_n743), .B(KEYINPUT46), .ZN(new_n744));
  OAI21_X1  g543(.A(G36gat), .B1(new_n740), .B2(new_n487), .ZN(new_n745));
  NAND2_X1  g544(.A1(new_n744), .A2(new_n745), .ZN(G1329gat));
  INV_X1    g545(.A(G43gat), .ZN(new_n747));
  INV_X1    g546(.A(new_n705), .ZN(new_n748));
  OAI21_X1  g547(.A(new_n747), .B1(new_n720), .B2(new_n748), .ZN(new_n749));
  NAND2_X1  g548(.A1(new_n707), .A2(G43gat), .ZN(new_n750));
  OAI21_X1  g549(.A(new_n749), .B1(new_n740), .B2(new_n750), .ZN(new_n751));
  XOR2_X1   g550(.A(KEYINPUT109), .B(KEYINPUT47), .Z(new_n752));
  XOR2_X1   g551(.A(new_n751), .B(new_n752), .Z(G1330gat));
  NOR2_X1   g552(.A1(new_n276), .A2(new_n265), .ZN(new_n754));
  NAND4_X1  g553(.A1(new_n731), .A2(new_n719), .A3(new_n739), .A4(new_n754), .ZN(new_n755));
  OAI21_X1  g554(.A(new_n265), .B1(new_n720), .B2(new_n276), .ZN(new_n756));
  INV_X1    g555(.A(KEYINPUT110), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n757), .A2(KEYINPUT48), .ZN(new_n758));
  NAND3_X1  g557(.A1(new_n755), .A2(new_n756), .A3(new_n758), .ZN(new_n759));
  NOR2_X1   g558(.A1(new_n757), .A2(KEYINPUT48), .ZN(new_n760));
  XOR2_X1   g559(.A(new_n759), .B(new_n760), .Z(G1331gat));
  NAND2_X1  g560(.A1(new_n490), .A2(new_n729), .ZN(new_n762));
  NOR3_X1   g561(.A1(new_n616), .A2(new_n691), .A3(new_n663), .ZN(new_n763));
  NAND2_X1  g562(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  NOR2_X1   g563(.A1(new_n764), .A2(new_n486), .ZN(new_n765));
  XNOR2_X1  g564(.A(new_n765), .B(new_n502), .ZN(G1332gat));
  INV_X1    g565(.A(new_n764), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n767), .A2(new_n353), .ZN(new_n768));
  NOR2_X1   g567(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n769));
  AND2_X1   g568(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n770));
  NOR3_X1   g569(.A1(new_n768), .A2(new_n769), .A3(new_n770), .ZN(new_n771));
  AOI21_X1  g570(.A(new_n771), .B1(new_n769), .B2(new_n768), .ZN(G1333gat));
  OAI21_X1  g571(.A(new_n512), .B1(new_n764), .B2(new_n748), .ZN(new_n773));
  NAND2_X1  g572(.A1(new_n707), .A2(G71gat), .ZN(new_n774));
  OAI21_X1  g573(.A(new_n773), .B1(new_n764), .B2(new_n774), .ZN(new_n775));
  XNOR2_X1  g574(.A(new_n775), .B(KEYINPUT50), .ZN(G1334gat));
  NOR2_X1   g575(.A1(new_n764), .A2(new_n276), .ZN(new_n777));
  XNOR2_X1  g576(.A(new_n777), .B(new_n513), .ZN(G1335gat));
  INV_X1    g577(.A(KEYINPUT113), .ZN(new_n779));
  NOR2_X1   g578(.A1(new_n661), .A2(new_n691), .ZN(new_n780));
  NAND3_X1  g579(.A1(new_n762), .A2(new_n736), .A3(new_n780), .ZN(new_n781));
  INV_X1    g580(.A(KEYINPUT51), .ZN(new_n782));
  NAND3_X1  g581(.A1(new_n781), .A2(KEYINPUT112), .A3(new_n782), .ZN(new_n783));
  NAND3_X1  g582(.A1(new_n730), .A2(KEYINPUT51), .A3(new_n780), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  AOI21_X1  g584(.A(KEYINPUT51), .B1(new_n730), .B2(new_n780), .ZN(new_n786));
  NOR2_X1   g585(.A1(new_n786), .A2(KEYINPUT112), .ZN(new_n787));
  OAI21_X1  g586(.A(new_n779), .B1(new_n785), .B2(new_n787), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n781), .A2(new_n782), .ZN(new_n789));
  INV_X1    g588(.A(KEYINPUT112), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  NAND4_X1  g590(.A1(new_n791), .A2(KEYINPUT113), .A3(new_n783), .A4(new_n784), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n788), .A2(new_n792), .ZN(new_n793));
  NOR2_X1   g592(.A1(new_n486), .A2(G85gat), .ZN(new_n794));
  NAND3_X1  g593(.A1(new_n793), .A2(new_n657), .A3(new_n794), .ZN(new_n795));
  NOR3_X1   g594(.A1(new_n661), .A2(new_n691), .A3(new_n663), .ZN(new_n796));
  XNOR2_X1  g595(.A(new_n796), .B(KEYINPUT111), .ZN(new_n797));
  OAI211_X1 g596(.A(new_n739), .B(new_n797), .C1(new_n730), .C2(KEYINPUT44), .ZN(new_n798));
  OAI21_X1  g597(.A(G85gat), .B1(new_n798), .B2(new_n486), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n795), .A2(new_n799), .ZN(G1336gat));
  OAI21_X1  g599(.A(G92gat), .B1(new_n798), .B2(new_n487), .ZN(new_n801));
  XNOR2_X1  g600(.A(KEYINPUT115), .B(KEYINPUT52), .ZN(new_n802));
  NOR2_X1   g601(.A1(new_n785), .A2(new_n787), .ZN(new_n803));
  NOR3_X1   g602(.A1(new_n487), .A2(new_n663), .A3(G92gat), .ZN(new_n804));
  XOR2_X1   g603(.A(new_n804), .B(KEYINPUT114), .Z(new_n805));
  OAI211_X1 g604(.A(new_n801), .B(new_n802), .C1(new_n803), .C2(new_n805), .ZN(new_n806));
  INV_X1    g605(.A(new_n784), .ZN(new_n807));
  NOR2_X1   g606(.A1(new_n807), .A2(new_n786), .ZN(new_n808));
  OAI21_X1  g607(.A(new_n801), .B1(new_n808), .B2(new_n805), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n809), .A2(KEYINPUT52), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n806), .A2(new_n810), .ZN(G1337gat));
  NOR2_X1   g610(.A1(new_n748), .A2(G99gat), .ZN(new_n812));
  NAND3_X1  g611(.A1(new_n793), .A2(new_n657), .A3(new_n812), .ZN(new_n813));
  OAI21_X1  g612(.A(G99gat), .B1(new_n798), .B2(new_n460), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n813), .A2(new_n814), .ZN(G1338gat));
  INV_X1    g614(.A(KEYINPUT53), .ZN(new_n816));
  OAI21_X1  g615(.A(G106gat), .B1(new_n798), .B2(new_n276), .ZN(new_n817));
  NOR3_X1   g616(.A1(new_n276), .A2(G106gat), .A3(new_n663), .ZN(new_n818));
  INV_X1    g617(.A(new_n818), .ZN(new_n819));
  OAI211_X1 g618(.A(new_n816), .B(new_n817), .C1(new_n803), .C2(new_n819), .ZN(new_n820));
  INV_X1    g619(.A(KEYINPUT116), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n817), .A2(new_n821), .ZN(new_n822));
  OAI211_X1 g621(.A(KEYINPUT116), .B(G106gat), .C1(new_n798), .C2(new_n276), .ZN(new_n823));
  OAI21_X1  g622(.A(new_n818), .B1(new_n807), .B2(new_n786), .ZN(new_n824));
  AND3_X1   g623(.A1(new_n822), .A2(new_n823), .A3(new_n824), .ZN(new_n825));
  OAI21_X1  g624(.A(new_n820), .B1(new_n825), .B2(new_n816), .ZN(G1339gat));
  NOR2_X1   g625(.A1(new_n486), .A2(new_n353), .ZN(new_n827));
  INV_X1    g626(.A(new_n827), .ZN(new_n828));
  INV_X1    g627(.A(new_n661), .ZN(new_n829));
  NAND3_X1  g628(.A1(new_n636), .A2(new_n637), .A3(new_n653), .ZN(new_n830));
  NAND3_X1  g629(.A1(new_n640), .A2(KEYINPUT54), .A3(new_n830), .ZN(new_n831));
  INV_X1    g630(.A(KEYINPUT54), .ZN(new_n832));
  AOI21_X1  g631(.A(new_n650), .B1(new_n654), .B2(new_n832), .ZN(new_n833));
  NAND3_X1  g632(.A1(new_n831), .A2(KEYINPUT55), .A3(new_n833), .ZN(new_n834));
  NAND2_X1  g633(.A1(new_n834), .A2(new_n651), .ZN(new_n835));
  INV_X1    g634(.A(KEYINPUT117), .ZN(new_n836));
  NAND2_X1  g635(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  NAND3_X1  g636(.A1(new_n834), .A2(KEYINPUT117), .A3(new_n651), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n831), .A2(new_n833), .ZN(new_n839));
  INV_X1    g638(.A(KEYINPUT55), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n839), .A2(new_n840), .ZN(new_n841));
  NAND4_X1  g640(.A1(new_n837), .A2(new_n691), .A3(new_n838), .A4(new_n841), .ZN(new_n842));
  NOR2_X1   g641(.A1(new_n678), .A2(new_n679), .ZN(new_n843));
  AOI21_X1  g642(.A(new_n669), .B1(new_n666), .B2(new_n668), .ZN(new_n844));
  OAI21_X1  g643(.A(new_n686), .B1(new_n843), .B2(new_n844), .ZN(new_n845));
  AND2_X1   g644(.A1(new_n690), .A2(new_n845), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n657), .A2(new_n846), .ZN(new_n847));
  AOI21_X1  g646(.A(new_n736), .B1(new_n842), .B2(new_n847), .ZN(new_n848));
  NAND3_X1  g647(.A1(new_n837), .A2(new_n838), .A3(new_n841), .ZN(new_n849));
  OAI21_X1  g648(.A(new_n846), .B1(new_n609), .B2(new_n614), .ZN(new_n850));
  NOR2_X1   g649(.A1(new_n849), .A2(new_n850), .ZN(new_n851));
  OAI21_X1  g650(.A(new_n829), .B1(new_n848), .B2(new_n851), .ZN(new_n852));
  NAND4_X1  g651(.A1(new_n661), .A2(new_n718), .A3(new_n615), .A4(new_n663), .ZN(new_n853));
  AOI21_X1  g652(.A(new_n828), .B1(new_n852), .B2(new_n853), .ZN(new_n854));
  NOR3_X1   g653(.A1(new_n461), .A2(new_n449), .A3(new_n450), .ZN(new_n855));
  NAND2_X1  g654(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  XNOR2_X1  g655(.A(new_n856), .B(KEYINPUT118), .ZN(new_n857));
  INV_X1    g656(.A(G113gat), .ZN(new_n858));
  NAND3_X1  g657(.A1(new_n857), .A2(new_n858), .A3(new_n691), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n854), .A2(new_n737), .ZN(new_n860));
  OAI21_X1  g659(.A(G113gat), .B1(new_n860), .B2(new_n718), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n859), .A2(new_n861), .ZN(G1340gat));
  INV_X1    g661(.A(G120gat), .ZN(new_n863));
  NAND3_X1  g662(.A1(new_n857), .A2(new_n863), .A3(new_n657), .ZN(new_n864));
  OAI21_X1  g663(.A(G120gat), .B1(new_n860), .B2(new_n663), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n864), .A2(new_n865), .ZN(G1341gat));
  OAI21_X1  g665(.A(G127gat), .B1(new_n860), .B2(new_n829), .ZN(new_n867));
  OR2_X1    g666(.A1(new_n829), .A2(G127gat), .ZN(new_n868));
  OAI21_X1  g667(.A(new_n867), .B1(new_n856), .B2(new_n868), .ZN(G1342gat));
  NOR2_X1   g668(.A1(new_n615), .A2(G134gat), .ZN(new_n870));
  NAND3_X1  g669(.A1(new_n854), .A2(new_n855), .A3(new_n870), .ZN(new_n871));
  XOR2_X1   g670(.A(new_n871), .B(KEYINPUT119), .Z(new_n872));
  XNOR2_X1  g671(.A(new_n872), .B(KEYINPUT56), .ZN(new_n873));
  OAI21_X1  g672(.A(G134gat), .B1(new_n860), .B2(new_n615), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n873), .A2(new_n874), .ZN(G1343gat));
  NOR2_X1   g674(.A1(new_n707), .A2(new_n276), .ZN(new_n876));
  NAND2_X1  g675(.A1(new_n854), .A2(new_n876), .ZN(new_n877));
  OAI21_X1  g676(.A(new_n221), .B1(new_n877), .B2(new_n718), .ZN(new_n878));
  NOR2_X1   g677(.A1(new_n707), .A2(new_n828), .ZN(new_n879));
  INV_X1    g678(.A(KEYINPUT57), .ZN(new_n880));
  INV_X1    g679(.A(new_n851), .ZN(new_n881));
  NAND2_X1  g680(.A1(new_n691), .A2(new_n841), .ZN(new_n882));
  OAI21_X1  g681(.A(new_n847), .B1(new_n882), .B2(new_n835), .ZN(new_n883));
  NAND2_X1  g682(.A1(new_n883), .A2(new_n615), .ZN(new_n884));
  NAND2_X1  g683(.A1(new_n881), .A2(new_n884), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n885), .A2(new_n829), .ZN(new_n886));
  AOI211_X1 g685(.A(new_n880), .B(new_n276), .C1(new_n886), .C2(new_n853), .ZN(new_n887));
  AOI21_X1  g686(.A(new_n276), .B1(new_n852), .B2(new_n853), .ZN(new_n888));
  NOR2_X1   g687(.A1(new_n888), .A2(KEYINPUT57), .ZN(new_n889));
  OAI21_X1  g688(.A(new_n879), .B1(new_n887), .B2(new_n889), .ZN(new_n890));
  NAND2_X1  g689(.A1(new_n691), .A2(G141gat), .ZN(new_n891));
  OAI21_X1  g690(.A(new_n878), .B1(new_n890), .B2(new_n891), .ZN(new_n892));
  XOR2_X1   g691(.A(new_n892), .B(KEYINPUT58), .Z(G1344gat));
  NOR2_X1   g692(.A1(new_n225), .A2(KEYINPUT59), .ZN(new_n894));
  OAI211_X1 g693(.A(KEYINPUT120), .B(new_n894), .C1(new_n890), .C2(new_n663), .ZN(new_n895));
  OR2_X1    g694(.A1(new_n888), .A2(new_n880), .ZN(new_n896));
  AND3_X1   g695(.A1(new_n658), .A2(new_n664), .A3(new_n718), .ZN(new_n897));
  AOI21_X1  g696(.A(new_n661), .B1(new_n881), .B2(new_n884), .ZN(new_n898));
  OAI211_X1 g697(.A(new_n880), .B(new_n461), .C1(new_n897), .C2(new_n898), .ZN(new_n899));
  NAND3_X1  g698(.A1(new_n896), .A2(new_n657), .A3(new_n899), .ZN(new_n900));
  INV_X1    g699(.A(new_n900), .ZN(new_n901));
  AOI21_X1  g700(.A(new_n216), .B1(new_n901), .B2(new_n879), .ZN(new_n902));
  XOR2_X1   g701(.A(KEYINPUT121), .B(KEYINPUT59), .Z(new_n903));
  OAI21_X1  g702(.A(new_n895), .B1(new_n902), .B2(new_n903), .ZN(new_n904));
  OR2_X1    g703(.A1(new_n890), .A2(new_n663), .ZN(new_n905));
  AOI21_X1  g704(.A(KEYINPUT120), .B1(new_n905), .B2(new_n894), .ZN(new_n906));
  NAND2_X1  g705(.A1(new_n657), .A2(new_n225), .ZN(new_n907));
  OAI22_X1  g706(.A1(new_n904), .A2(new_n906), .B1(new_n877), .B2(new_n907), .ZN(G1345gat));
  NAND2_X1  g707(.A1(new_n661), .A2(G155gat), .ZN(new_n909));
  XNOR2_X1  g708(.A(new_n909), .B(KEYINPUT122), .ZN(new_n910));
  NOR2_X1   g709(.A1(new_n890), .A2(new_n910), .ZN(new_n911));
  INV_X1    g710(.A(G155gat), .ZN(new_n912));
  NAND3_X1  g711(.A1(new_n854), .A2(new_n661), .A3(new_n876), .ZN(new_n913));
  AOI21_X1  g712(.A(new_n911), .B1(new_n912), .B2(new_n913), .ZN(G1346gat));
  OAI21_X1  g713(.A(G162gat), .B1(new_n890), .B2(new_n615), .ZN(new_n915));
  OR2_X1    g714(.A1(new_n615), .A2(G162gat), .ZN(new_n916));
  OAI21_X1  g715(.A(new_n915), .B1(new_n877), .B2(new_n916), .ZN(G1347gat));
  NAND2_X1  g716(.A1(new_n852), .A2(new_n853), .ZN(new_n918));
  NOR2_X1   g717(.A1(new_n469), .A2(new_n487), .ZN(new_n919));
  AND2_X1   g718(.A1(new_n737), .A2(new_n919), .ZN(new_n920));
  NAND2_X1  g719(.A1(new_n918), .A2(new_n920), .ZN(new_n921));
  NOR3_X1   g720(.A1(new_n921), .A2(new_n684), .A3(new_n718), .ZN(new_n922));
  NAND2_X1  g721(.A1(new_n918), .A2(new_n486), .ZN(new_n923));
  INV_X1    g722(.A(KEYINPUT123), .ZN(new_n924));
  NAND2_X1  g723(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  NAND3_X1  g724(.A1(new_n918), .A2(KEYINPUT123), .A3(new_n486), .ZN(new_n926));
  AOI21_X1  g725(.A(new_n487), .B1(new_n925), .B2(new_n926), .ZN(new_n927));
  NAND3_X1  g726(.A1(new_n927), .A2(new_n855), .A3(new_n691), .ZN(new_n928));
  AOI21_X1  g727(.A(new_n922), .B1(new_n928), .B2(new_n684), .ZN(G1348gat));
  OAI21_X1  g728(.A(G176gat), .B1(new_n921), .B2(new_n663), .ZN(new_n930));
  NAND2_X1  g729(.A1(new_n927), .A2(new_n855), .ZN(new_n931));
  OR2_X1    g730(.A1(new_n663), .A2(G176gat), .ZN(new_n932));
  OAI21_X1  g731(.A(new_n930), .B1(new_n931), .B2(new_n932), .ZN(G1349gat));
  OAI21_X1  g732(.A(G183gat), .B1(new_n921), .B2(new_n829), .ZN(new_n934));
  NAND2_X1  g733(.A1(new_n661), .A2(new_n309), .ZN(new_n935));
  OAI21_X1  g734(.A(new_n934), .B1(new_n931), .B2(new_n935), .ZN(new_n936));
  XNOR2_X1  g735(.A(new_n936), .B(KEYINPUT60), .ZN(G1350gat));
  NAND3_X1  g736(.A1(new_n918), .A2(new_n736), .A3(new_n920), .ZN(new_n938));
  AND2_X1   g737(.A1(new_n938), .A2(G190gat), .ZN(new_n939));
  INV_X1    g738(.A(KEYINPUT61), .ZN(new_n940));
  NOR2_X1   g739(.A1(new_n939), .A2(new_n940), .ZN(new_n941));
  NAND2_X1  g740(.A1(new_n939), .A2(new_n940), .ZN(new_n942));
  AOI21_X1  g741(.A(new_n941), .B1(KEYINPUT124), .B2(new_n942), .ZN(new_n943));
  OAI21_X1  g742(.A(new_n943), .B1(KEYINPUT124), .B2(new_n942), .ZN(new_n944));
  NAND2_X1  g743(.A1(new_n736), .A2(new_n310), .ZN(new_n945));
  OAI21_X1  g744(.A(new_n944), .B1(new_n931), .B2(new_n945), .ZN(G1351gat));
  AOI21_X1  g745(.A(KEYINPUT123), .B1(new_n918), .B2(new_n486), .ZN(new_n947));
  AOI211_X1 g746(.A(new_n924), .B(new_n469), .C1(new_n852), .C2(new_n853), .ZN(new_n948));
  OAI211_X1 g747(.A(new_n353), .B(new_n876), .C1(new_n947), .C2(new_n948), .ZN(new_n949));
  NOR3_X1   g748(.A1(new_n949), .A2(G197gat), .A3(new_n718), .ZN(new_n950));
  OR2_X1    g749(.A1(new_n950), .A2(KEYINPUT125), .ZN(new_n951));
  NAND2_X1  g750(.A1(new_n950), .A2(KEYINPUT125), .ZN(new_n952));
  NAND2_X1  g751(.A1(new_n460), .A2(new_n919), .ZN(new_n953));
  INV_X1    g752(.A(new_n953), .ZN(new_n954));
  NAND3_X1  g753(.A1(new_n896), .A2(new_n899), .A3(new_n954), .ZN(new_n955));
  OAI21_X1  g754(.A(G197gat), .B1(new_n955), .B2(new_n718), .ZN(new_n956));
  NAND3_X1  g755(.A1(new_n951), .A2(new_n952), .A3(new_n956), .ZN(G1352gat));
  NOR2_X1   g756(.A1(new_n663), .A2(G204gat), .ZN(new_n958));
  NAND4_X1  g757(.A1(new_n927), .A2(KEYINPUT62), .A3(new_n876), .A4(new_n958), .ZN(new_n959));
  INV_X1    g758(.A(KEYINPUT62), .ZN(new_n960));
  INV_X1    g759(.A(new_n958), .ZN(new_n961));
  OAI21_X1  g760(.A(new_n960), .B1(new_n949), .B2(new_n961), .ZN(new_n962));
  NAND2_X1  g761(.A1(new_n959), .A2(new_n962), .ZN(new_n963));
  OAI21_X1  g762(.A(G204gat), .B1(new_n900), .B2(new_n953), .ZN(new_n964));
  NAND2_X1  g763(.A1(new_n963), .A2(new_n964), .ZN(new_n965));
  NAND2_X1  g764(.A1(new_n965), .A2(KEYINPUT126), .ZN(new_n966));
  INV_X1    g765(.A(KEYINPUT126), .ZN(new_n967));
  NAND3_X1  g766(.A1(new_n963), .A2(new_n967), .A3(new_n964), .ZN(new_n968));
  NAND2_X1  g767(.A1(new_n966), .A2(new_n968), .ZN(G1353gat));
  INV_X1    g768(.A(KEYINPUT127), .ZN(new_n970));
  NAND4_X1  g769(.A1(new_n896), .A2(new_n899), .A3(new_n661), .A4(new_n954), .ZN(new_n971));
  NAND2_X1  g770(.A1(new_n971), .A2(G211gat), .ZN(new_n972));
  INV_X1    g771(.A(KEYINPUT63), .ZN(new_n973));
  OAI21_X1  g772(.A(new_n970), .B1(new_n972), .B2(new_n973), .ZN(new_n974));
  NAND2_X1  g773(.A1(new_n972), .A2(new_n973), .ZN(new_n975));
  NAND2_X1  g774(.A1(new_n974), .A2(new_n975), .ZN(new_n976));
  NOR3_X1   g775(.A1(new_n972), .A2(new_n970), .A3(new_n973), .ZN(new_n977));
  OR2_X1    g776(.A1(new_n829), .A2(G211gat), .ZN(new_n978));
  OAI22_X1  g777(.A1(new_n976), .A2(new_n977), .B1(new_n949), .B2(new_n978), .ZN(G1354gat));
  OAI21_X1  g778(.A(G218gat), .B1(new_n955), .B2(new_n615), .ZN(new_n980));
  OR2_X1    g779(.A1(new_n615), .A2(G218gat), .ZN(new_n981));
  OAI21_X1  g780(.A(new_n980), .B1(new_n949), .B2(new_n981), .ZN(G1355gat));
endmodule


