

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n678, n679, n680, n681, n682, n683, n684, n685,
         n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696,
         n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707,
         n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718,
         n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729,
         n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740,
         n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751,
         n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762,
         n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773,
         n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784,
         n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, n795,
         n796, n797, n798, n799, n800, n801, n802, n803, n804, n805, n806,
         n807, n808, n809, n810, n811, n812, n813, n814, n815, n816, n817,
         n818, n819, n820, n821, n822, n823, n824, n825, n826, n827, n828,
         n829, n830, n831, n832, n833, n834, n835, n836, n837, n838, n839,
         n840, n841, n842, n843, n844, n845, n846, n847, n848, n849, n850,
         n851, n852, n853, n854, n855, n856, n857, n858, n859, n860, n861,
         n862, n863, n864, n865, n866, n867, n868, n869, n870, n871, n872,
         n873, n874, n875, n876, n877, n878, n879, n880, n881, n882, n883,
         n884, n885, n886, n887, n888, n889, n890, n891, n892, n893, n894,
         n895, n896, n897, n898, n899, n900, n901, n902, n903, n904, n905,
         n906, n907, n908, n909, n910, n911, n912, n913, n914, n915, n916,
         n917, n918, n919, n920, n921, n922, n923, n924, n925, n926, n927,
         n928, n929, n930, n931, n932, n933, n934, n935, n936, n937, n938,
         n939, n940, n941, n942, n943, n944, n945, n946, n947, n948, n949,
         n950, n951, n952, n953, n954, n955, n956, n957, n958, n959, n960,
         n961, n962, n963, n964, n965, n966, n967, n968, n969, n970, n971,
         n972, n973, n974, n975, n976, n977, n978, n979, n980, n981, n982,
         n983, n984, n985, n986, n987, n988, n989, n990, n991, n992, n993,
         n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NOR2_X2 U551 ( .A1(n774), .A2(n678), .ZN(n707) );
  NOR2_X1 U552 ( .A1(n757), .A2(n754), .ZN(n516) );
  AND2_X1 U553 ( .A1(n792), .A2(n807), .ZN(n517) );
  INV_X1 U554 ( .A(KEYINPUT95), .ZN(n683) );
  INV_X1 U555 ( .A(KEYINPUT97), .ZN(n714) );
  XNOR2_X1 U556 ( .A(n714), .B(KEYINPUT30), .ZN(n715) );
  XNOR2_X1 U557 ( .A(n716), .B(n715), .ZN(n717) );
  NOR2_X1 U558 ( .A1(n711), .A2(n710), .ZN(n712) );
  AND2_X1 U559 ( .A1(n736), .A2(n735), .ZN(n737) );
  NOR2_X1 U560 ( .A1(n524), .A2(G2105), .ZN(n602) );
  NOR2_X1 U561 ( .A1(G1384), .A2(G164), .ZN(n775) );
  NOR2_X1 U562 ( .A1(n566), .A2(n565), .ZN(n567) );
  AND2_X1 U563 ( .A1(n795), .A2(n794), .ZN(n796) );
  NOR2_X1 U564 ( .A1(G543), .A2(n543), .ZN(n544) );
  NOR2_X1 U565 ( .A1(G543), .A2(G651), .ZN(n642) );
  AND2_X1 U566 ( .A1(G2105), .A2(n524), .ZN(n871) );
  XNOR2_X1 U567 ( .A(n569), .B(KEYINPUT15), .ZN(n962) );
  NOR2_X1 U568 ( .A1(n618), .A2(G651), .ZN(n639) );
  NOR2_X1 U569 ( .A1(n528), .A2(n527), .ZN(G160) );
  XOR2_X1 U570 ( .A(G2104), .B(KEYINPUT64), .Z(n524) );
  NAND2_X1 U571 ( .A1(G101), .A2(n602), .ZN(n518) );
  XNOR2_X1 U572 ( .A(n518), .B(KEYINPUT23), .ZN(n519) );
  XNOR2_X1 U573 ( .A(n519), .B(KEYINPUT65), .ZN(n522) );
  AND2_X1 U574 ( .A1(G2105), .A2(G2104), .ZN(n870) );
  NAND2_X1 U575 ( .A1(G113), .A2(n870), .ZN(n520) );
  XNOR2_X1 U576 ( .A(n520), .B(KEYINPUT66), .ZN(n521) );
  NAND2_X1 U577 ( .A1(n522), .A2(n521), .ZN(n528) );
  NOR2_X1 U578 ( .A1(G2105), .A2(G2104), .ZN(n523) );
  XOR2_X1 U579 ( .A(KEYINPUT17), .B(n523), .Z(n531) );
  BUF_X1 U580 ( .A(n531), .Z(n875) );
  NAND2_X1 U581 ( .A1(G137), .A2(n875), .ZN(n526) );
  NAND2_X1 U582 ( .A1(G125), .A2(n871), .ZN(n525) );
  NAND2_X1 U583 ( .A1(n526), .A2(n525), .ZN(n527) );
  NAND2_X1 U584 ( .A1(G114), .A2(n870), .ZN(n530) );
  NAND2_X1 U585 ( .A1(G102), .A2(n602), .ZN(n529) );
  NAND2_X1 U586 ( .A1(n530), .A2(n529), .ZN(n535) );
  NAND2_X1 U587 ( .A1(G138), .A2(n531), .ZN(n533) );
  NAND2_X1 U588 ( .A1(G126), .A2(n871), .ZN(n532) );
  NAND2_X1 U589 ( .A1(n533), .A2(n532), .ZN(n534) );
  NOR2_X1 U590 ( .A1(n535), .A2(n534), .ZN(n536) );
  XNOR2_X1 U591 ( .A(n536), .B(KEYINPUT86), .ZN(G164) );
  AND2_X1 U592 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U593 ( .A(G132), .ZN(G219) );
  INV_X1 U594 ( .A(G82), .ZN(G220) );
  NAND2_X1 U595 ( .A1(G90), .A2(n642), .ZN(n539) );
  XOR2_X1 U596 ( .A(KEYINPUT0), .B(G543), .Z(n618) );
  XNOR2_X1 U597 ( .A(KEYINPUT67), .B(G651), .ZN(n543) );
  NOR2_X1 U598 ( .A1(n618), .A2(n543), .ZN(n537) );
  XNOR2_X1 U599 ( .A(KEYINPUT68), .B(n537), .ZN(n638) );
  NAND2_X1 U600 ( .A1(G77), .A2(n638), .ZN(n538) );
  NAND2_X1 U601 ( .A1(n539), .A2(n538), .ZN(n542) );
  XOR2_X1 U602 ( .A(KEYINPUT70), .B(KEYINPUT71), .Z(n540) );
  XNOR2_X1 U603 ( .A(KEYINPUT9), .B(n540), .ZN(n541) );
  XNOR2_X1 U604 ( .A(n542), .B(n541), .ZN(n548) );
  XOR2_X1 U605 ( .A(KEYINPUT1), .B(n544), .Z(n643) );
  NAND2_X1 U606 ( .A1(n643), .A2(G64), .ZN(n546) );
  NAND2_X1 U607 ( .A1(n639), .A2(G52), .ZN(n545) );
  AND2_X1 U608 ( .A1(n546), .A2(n545), .ZN(n547) );
  NAND2_X1 U609 ( .A1(n548), .A2(n547), .ZN(G301) );
  XOR2_X1 U610 ( .A(KEYINPUT10), .B(KEYINPUT75), .Z(n550) );
  NAND2_X1 U611 ( .A1(G7), .A2(G661), .ZN(n549) );
  XOR2_X1 U612 ( .A(n550), .B(n549), .Z(n907) );
  NAND2_X1 U613 ( .A1(n907), .A2(G567), .ZN(n551) );
  XOR2_X1 U614 ( .A(KEYINPUT11), .B(n551), .Z(G234) );
  NAND2_X1 U615 ( .A1(n643), .A2(G56), .ZN(n552) );
  XOR2_X1 U616 ( .A(KEYINPUT14), .B(n552), .Z(n559) );
  NAND2_X1 U617 ( .A1(n642), .A2(G81), .ZN(n553) );
  XOR2_X1 U618 ( .A(KEYINPUT12), .B(n553), .Z(n556) );
  NAND2_X1 U619 ( .A1(n638), .A2(G68), .ZN(n554) );
  XOR2_X1 U620 ( .A(KEYINPUT76), .B(n554), .Z(n555) );
  NOR2_X1 U621 ( .A1(n556), .A2(n555), .ZN(n557) );
  XNOR2_X1 U622 ( .A(n557), .B(KEYINPUT13), .ZN(n558) );
  NOR2_X1 U623 ( .A1(n559), .A2(n558), .ZN(n561) );
  NAND2_X1 U624 ( .A1(n639), .A2(G43), .ZN(n560) );
  NAND2_X1 U625 ( .A1(n561), .A2(n560), .ZN(n978) );
  INV_X1 U626 ( .A(G860), .ZN(n609) );
  OR2_X1 U627 ( .A1(n978), .A2(n609), .ZN(G153) );
  NAND2_X1 U628 ( .A1(G868), .A2(G301), .ZN(n571) );
  NAND2_X1 U629 ( .A1(G54), .A2(n639), .ZN(n568) );
  NAND2_X1 U630 ( .A1(G92), .A2(n642), .ZN(n563) );
  NAND2_X1 U631 ( .A1(G79), .A2(n638), .ZN(n562) );
  NAND2_X1 U632 ( .A1(n563), .A2(n562), .ZN(n566) );
  NAND2_X1 U633 ( .A1(G66), .A2(n643), .ZN(n564) );
  XNOR2_X1 U634 ( .A(KEYINPUT77), .B(n564), .ZN(n565) );
  NAND2_X1 U635 ( .A1(n568), .A2(n567), .ZN(n569) );
  OR2_X1 U636 ( .A1(n962), .A2(G868), .ZN(n570) );
  NAND2_X1 U637 ( .A1(n571), .A2(n570), .ZN(G284) );
  NAND2_X1 U638 ( .A1(n639), .A2(G51), .ZN(n573) );
  NAND2_X1 U639 ( .A1(G63), .A2(n643), .ZN(n572) );
  NAND2_X1 U640 ( .A1(n573), .A2(n572), .ZN(n574) );
  XNOR2_X1 U641 ( .A(KEYINPUT6), .B(n574), .ZN(n581) );
  NAND2_X1 U642 ( .A1(n642), .A2(G89), .ZN(n575) );
  XNOR2_X1 U643 ( .A(n575), .B(KEYINPUT4), .ZN(n577) );
  NAND2_X1 U644 ( .A1(G76), .A2(n638), .ZN(n576) );
  NAND2_X1 U645 ( .A1(n577), .A2(n576), .ZN(n578) );
  XOR2_X1 U646 ( .A(KEYINPUT78), .B(n578), .Z(n579) );
  XNOR2_X1 U647 ( .A(KEYINPUT5), .B(n579), .ZN(n580) );
  NOR2_X1 U648 ( .A1(n581), .A2(n580), .ZN(n583) );
  XNOR2_X1 U649 ( .A(KEYINPUT79), .B(KEYINPUT7), .ZN(n582) );
  XNOR2_X1 U650 ( .A(n583), .B(n582), .ZN(G168) );
  XOR2_X1 U651 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U652 ( .A1(n639), .A2(G53), .ZN(n585) );
  NAND2_X1 U653 ( .A1(G65), .A2(n643), .ZN(n584) );
  NAND2_X1 U654 ( .A1(n585), .A2(n584), .ZN(n586) );
  XOR2_X1 U655 ( .A(KEYINPUT72), .B(n586), .Z(n590) );
  NAND2_X1 U656 ( .A1(n642), .A2(G91), .ZN(n588) );
  NAND2_X1 U657 ( .A1(G78), .A2(n638), .ZN(n587) );
  AND2_X1 U658 ( .A1(n588), .A2(n587), .ZN(n589) );
  NAND2_X1 U659 ( .A1(n590), .A2(n589), .ZN(n969) );
  XOR2_X1 U660 ( .A(KEYINPUT73), .B(n969), .Z(G299) );
  NAND2_X1 U661 ( .A1(G286), .A2(G868), .ZN(n592) );
  INV_X1 U662 ( .A(G868), .ZN(n659) );
  NAND2_X1 U663 ( .A1(n659), .A2(G299), .ZN(n591) );
  NAND2_X1 U664 ( .A1(n592), .A2(n591), .ZN(G297) );
  NAND2_X1 U665 ( .A1(n609), .A2(G559), .ZN(n593) );
  NAND2_X1 U666 ( .A1(n593), .A2(n962), .ZN(n594) );
  XNOR2_X1 U667 ( .A(n594), .B(KEYINPUT16), .ZN(n595) );
  XNOR2_X1 U668 ( .A(KEYINPUT80), .B(n595), .ZN(G148) );
  NOR2_X1 U669 ( .A1(G868), .A2(n978), .ZN(n598) );
  NAND2_X1 U670 ( .A1(G868), .A2(n962), .ZN(n596) );
  NOR2_X1 U671 ( .A1(G559), .A2(n596), .ZN(n597) );
  NOR2_X1 U672 ( .A1(n598), .A2(n597), .ZN(G282) );
  NAND2_X1 U673 ( .A1(G111), .A2(n870), .ZN(n600) );
  NAND2_X1 U674 ( .A1(G135), .A2(n875), .ZN(n599) );
  NAND2_X1 U675 ( .A1(n600), .A2(n599), .ZN(n606) );
  NAND2_X1 U676 ( .A1(n871), .A2(G123), .ZN(n601) );
  XNOR2_X1 U677 ( .A(n601), .B(KEYINPUT18), .ZN(n604) );
  BUF_X1 U678 ( .A(n602), .Z(n877) );
  NAND2_X1 U679 ( .A1(G99), .A2(n877), .ZN(n603) );
  NAND2_X1 U680 ( .A1(n604), .A2(n603), .ZN(n605) );
  NOR2_X1 U681 ( .A1(n606), .A2(n605), .ZN(n908) );
  XNOR2_X1 U682 ( .A(n908), .B(G2096), .ZN(n607) );
  INV_X1 U683 ( .A(G2100), .ZN(n819) );
  NAND2_X1 U684 ( .A1(n607), .A2(n819), .ZN(G156) );
  NAND2_X1 U685 ( .A1(G559), .A2(n962), .ZN(n608) );
  XOR2_X1 U686 ( .A(n978), .B(n608), .Z(n655) );
  NAND2_X1 U687 ( .A1(n609), .A2(n655), .ZN(n617) );
  NAND2_X1 U688 ( .A1(n638), .A2(G80), .ZN(n611) );
  NAND2_X1 U689 ( .A1(G67), .A2(n643), .ZN(n610) );
  NAND2_X1 U690 ( .A1(n611), .A2(n610), .ZN(n614) );
  NAND2_X1 U691 ( .A1(G55), .A2(n639), .ZN(n612) );
  XNOR2_X1 U692 ( .A(KEYINPUT81), .B(n612), .ZN(n613) );
  NOR2_X1 U693 ( .A1(n614), .A2(n613), .ZN(n616) );
  NAND2_X1 U694 ( .A1(n642), .A2(G93), .ZN(n615) );
  NAND2_X1 U695 ( .A1(n616), .A2(n615), .ZN(n658) );
  XNOR2_X1 U696 ( .A(n617), .B(n658), .ZN(G145) );
  NAND2_X1 U697 ( .A1(G74), .A2(G651), .ZN(n620) );
  NAND2_X1 U698 ( .A1(G87), .A2(n618), .ZN(n619) );
  NAND2_X1 U699 ( .A1(n620), .A2(n619), .ZN(n621) );
  NOR2_X1 U700 ( .A1(n643), .A2(n621), .ZN(n623) );
  NAND2_X1 U701 ( .A1(n639), .A2(G49), .ZN(n622) );
  NAND2_X1 U702 ( .A1(n623), .A2(n622), .ZN(G288) );
  NAND2_X1 U703 ( .A1(n638), .A2(G75), .ZN(n625) );
  NAND2_X1 U704 ( .A1(G62), .A2(n643), .ZN(n624) );
  NAND2_X1 U705 ( .A1(n625), .A2(n624), .ZN(n629) );
  NAND2_X1 U706 ( .A1(G88), .A2(n642), .ZN(n627) );
  NAND2_X1 U707 ( .A1(G50), .A2(n639), .ZN(n626) );
  NAND2_X1 U708 ( .A1(n627), .A2(n626), .ZN(n628) );
  NOR2_X1 U709 ( .A1(n629), .A2(n628), .ZN(G166) );
  INV_X1 U710 ( .A(G166), .ZN(G303) );
  NAND2_X1 U711 ( .A1(G73), .A2(n638), .ZN(n630) );
  XNOR2_X1 U712 ( .A(n630), .B(KEYINPUT2), .ZN(n637) );
  NAND2_X1 U713 ( .A1(n642), .A2(G86), .ZN(n632) );
  NAND2_X1 U714 ( .A1(G61), .A2(n643), .ZN(n631) );
  NAND2_X1 U715 ( .A1(n632), .A2(n631), .ZN(n635) );
  NAND2_X1 U716 ( .A1(n639), .A2(G48), .ZN(n633) );
  XOR2_X1 U717 ( .A(KEYINPUT82), .B(n633), .Z(n634) );
  NOR2_X1 U718 ( .A1(n635), .A2(n634), .ZN(n636) );
  NAND2_X1 U719 ( .A1(n637), .A2(n636), .ZN(G305) );
  NAND2_X1 U720 ( .A1(G72), .A2(n638), .ZN(n641) );
  NAND2_X1 U721 ( .A1(G47), .A2(n639), .ZN(n640) );
  NAND2_X1 U722 ( .A1(n641), .A2(n640), .ZN(n647) );
  NAND2_X1 U723 ( .A1(n642), .A2(G85), .ZN(n645) );
  NAND2_X1 U724 ( .A1(G60), .A2(n643), .ZN(n644) );
  NAND2_X1 U725 ( .A1(n645), .A2(n644), .ZN(n646) );
  NOR2_X1 U726 ( .A1(n647), .A2(n646), .ZN(n648) );
  XNOR2_X1 U727 ( .A(n648), .B(KEYINPUT69), .ZN(G290) );
  XNOR2_X1 U728 ( .A(KEYINPUT83), .B(KEYINPUT19), .ZN(n650) );
  XOR2_X1 U729 ( .A(G288), .B(G303), .Z(n649) );
  XNOR2_X1 U730 ( .A(n650), .B(n649), .ZN(n651) );
  XNOR2_X1 U731 ( .A(n651), .B(G305), .ZN(n652) );
  XNOR2_X1 U732 ( .A(n652), .B(n658), .ZN(n653) );
  XNOR2_X1 U733 ( .A(n653), .B(G290), .ZN(n654) );
  XNOR2_X1 U734 ( .A(n654), .B(G299), .ZN(n888) );
  XNOR2_X1 U735 ( .A(n888), .B(n655), .ZN(n656) );
  NAND2_X1 U736 ( .A1(n656), .A2(G868), .ZN(n657) );
  XNOR2_X1 U737 ( .A(n657), .B(KEYINPUT84), .ZN(n661) );
  NAND2_X1 U738 ( .A1(n659), .A2(n658), .ZN(n660) );
  NAND2_X1 U739 ( .A1(n661), .A2(n660), .ZN(G295) );
  NAND2_X1 U740 ( .A1(G2084), .A2(G2078), .ZN(n662) );
  XOR2_X1 U741 ( .A(KEYINPUT20), .B(n662), .Z(n663) );
  NAND2_X1 U742 ( .A1(G2090), .A2(n663), .ZN(n664) );
  XNOR2_X1 U743 ( .A(KEYINPUT21), .B(n664), .ZN(n665) );
  NAND2_X1 U744 ( .A1(n665), .A2(G2072), .ZN(G158) );
  XOR2_X1 U745 ( .A(KEYINPUT74), .B(G57), .Z(G237) );
  XOR2_X1 U746 ( .A(KEYINPUT85), .B(G44), .Z(n666) );
  XNOR2_X1 U747 ( .A(KEYINPUT3), .B(n666), .ZN(G218) );
  NAND2_X1 U748 ( .A1(G108), .A2(G120), .ZN(n667) );
  NOR2_X1 U749 ( .A1(G237), .A2(n667), .ZN(n668) );
  NAND2_X1 U750 ( .A1(G69), .A2(n668), .ZN(n816) );
  NAND2_X1 U751 ( .A1(n816), .A2(G567), .ZN(n673) );
  NOR2_X1 U752 ( .A1(G220), .A2(G219), .ZN(n669) );
  XOR2_X1 U753 ( .A(KEYINPUT22), .B(n669), .Z(n670) );
  NOR2_X1 U754 ( .A1(G218), .A2(n670), .ZN(n671) );
  NAND2_X1 U755 ( .A1(G96), .A2(n671), .ZN(n817) );
  NAND2_X1 U756 ( .A1(n817), .A2(G2106), .ZN(n672) );
  NAND2_X1 U757 ( .A1(n673), .A2(n672), .ZN(n818) );
  NAND2_X1 U758 ( .A1(G661), .A2(G483), .ZN(n674) );
  NOR2_X1 U759 ( .A1(n818), .A2(n674), .ZN(n813) );
  NAND2_X1 U760 ( .A1(n813), .A2(G36), .ZN(G176) );
  NOR2_X1 U761 ( .A1(G2090), .A2(G303), .ZN(n675) );
  NAND2_X1 U762 ( .A1(G8), .A2(n675), .ZN(n676) );
  XNOR2_X1 U763 ( .A(n676), .B(KEYINPUT102), .ZN(n743) );
  NAND2_X1 U764 ( .A1(G160), .A2(G40), .ZN(n774) );
  INV_X1 U765 ( .A(n775), .ZN(n678) );
  XOR2_X2 U766 ( .A(KEYINPUT92), .B(n707), .Z(n706) );
  INV_X1 U767 ( .A(G2072), .ZN(n923) );
  NOR2_X1 U768 ( .A1(n706), .A2(n923), .ZN(n680) );
  XOR2_X1 U769 ( .A(KEYINPUT27), .B(KEYINPUT93), .Z(n679) );
  XNOR2_X1 U770 ( .A(n680), .B(n679), .ZN(n700) );
  NAND2_X1 U771 ( .A1(n706), .A2(G1956), .ZN(n699) );
  INV_X1 U772 ( .A(n969), .ZN(n681) );
  AND2_X1 U773 ( .A1(n699), .A2(n681), .ZN(n682) );
  NAND2_X1 U774 ( .A1(n700), .A2(n682), .ZN(n684) );
  XNOR2_X1 U775 ( .A(n684), .B(n683), .ZN(n698) );
  INV_X1 U776 ( .A(n707), .ZN(n725) );
  NAND2_X1 U777 ( .A1(G1348), .A2(n725), .ZN(n685) );
  XOR2_X1 U778 ( .A(KEYINPUT94), .B(n685), .Z(n687) );
  INV_X1 U779 ( .A(G2067), .ZN(n822) );
  NOR2_X1 U780 ( .A1(n706), .A2(n822), .ZN(n686) );
  NOR2_X1 U781 ( .A1(n687), .A2(n686), .ZN(n688) );
  OR2_X1 U782 ( .A1(n962), .A2(n688), .ZN(n696) );
  NAND2_X1 U783 ( .A1(n962), .A2(n688), .ZN(n694) );
  AND2_X1 U784 ( .A1(n707), .A2(G1996), .ZN(n689) );
  XOR2_X1 U785 ( .A(n689), .B(KEYINPUT26), .Z(n691) );
  NAND2_X1 U786 ( .A1(n725), .A2(G1341), .ZN(n690) );
  NAND2_X1 U787 ( .A1(n691), .A2(n690), .ZN(n692) );
  OR2_X1 U788 ( .A1(n978), .A2(n692), .ZN(n693) );
  NAND2_X1 U789 ( .A1(n694), .A2(n693), .ZN(n695) );
  NAND2_X1 U790 ( .A1(n696), .A2(n695), .ZN(n697) );
  NAND2_X1 U791 ( .A1(n698), .A2(n697), .ZN(n704) );
  NAND2_X1 U792 ( .A1(n700), .A2(n699), .ZN(n701) );
  NAND2_X1 U793 ( .A1(n969), .A2(n701), .ZN(n702) );
  XNOR2_X1 U794 ( .A(n702), .B(KEYINPUT28), .ZN(n703) );
  NAND2_X1 U795 ( .A1(n704), .A2(n703), .ZN(n705) );
  XNOR2_X1 U796 ( .A(n705), .B(KEYINPUT29), .ZN(n711) );
  XOR2_X1 U797 ( .A(KEYINPUT25), .B(G2078), .Z(n941) );
  NOR2_X1 U798 ( .A1(n941), .A2(n706), .ZN(n709) );
  NOR2_X1 U799 ( .A1(n707), .A2(G1961), .ZN(n708) );
  NOR2_X1 U800 ( .A1(n709), .A2(n708), .ZN(n718) );
  NOR2_X1 U801 ( .A1(G301), .A2(n718), .ZN(n710) );
  XOR2_X1 U802 ( .A(KEYINPUT96), .B(n712), .Z(n723) );
  NOR2_X1 U803 ( .A1(G2084), .A2(n725), .ZN(n738) );
  NAND2_X1 U804 ( .A1(G8), .A2(n725), .ZN(n757) );
  NOR2_X1 U805 ( .A1(G1966), .A2(n757), .ZN(n734) );
  NOR2_X1 U806 ( .A1(n738), .A2(n734), .ZN(n713) );
  NAND2_X1 U807 ( .A1(G8), .A2(n713), .ZN(n716) );
  NOR2_X1 U808 ( .A1(G168), .A2(n717), .ZN(n720) );
  AND2_X1 U809 ( .A1(G301), .A2(n718), .ZN(n719) );
  NOR2_X1 U810 ( .A1(n720), .A2(n719), .ZN(n721) );
  XOR2_X1 U811 ( .A(KEYINPUT31), .B(n721), .Z(n722) );
  NAND2_X1 U812 ( .A1(n723), .A2(n722), .ZN(n735) );
  NAND2_X1 U813 ( .A1(n735), .A2(G286), .ZN(n731) );
  NOR2_X1 U814 ( .A1(G1971), .A2(n757), .ZN(n724) );
  XNOR2_X1 U815 ( .A(KEYINPUT99), .B(n724), .ZN(n729) );
  NOR2_X1 U816 ( .A1(G2090), .A2(n725), .ZN(n726) );
  XNOR2_X1 U817 ( .A(KEYINPUT100), .B(n726), .ZN(n727) );
  NOR2_X1 U818 ( .A1(G166), .A2(n727), .ZN(n728) );
  NAND2_X1 U819 ( .A1(n729), .A2(n728), .ZN(n730) );
  NAND2_X1 U820 ( .A1(n731), .A2(n730), .ZN(n732) );
  NAND2_X1 U821 ( .A1(n732), .A2(G8), .ZN(n733) );
  XNOR2_X1 U822 ( .A(n733), .B(KEYINPUT32), .ZN(n742) );
  INV_X1 U823 ( .A(n734), .ZN(n736) );
  XNOR2_X1 U824 ( .A(n737), .B(KEYINPUT98), .ZN(n740) );
  NAND2_X1 U825 ( .A1(n738), .A2(G8), .ZN(n739) );
  NAND2_X1 U826 ( .A1(n740), .A2(n739), .ZN(n741) );
  NAND2_X1 U827 ( .A1(n742), .A2(n741), .ZN(n753) );
  NAND2_X1 U828 ( .A1(n743), .A2(n753), .ZN(n744) );
  NAND2_X1 U829 ( .A1(n744), .A2(n757), .ZN(n745) );
  XNOR2_X1 U830 ( .A(n745), .B(KEYINPUT103), .ZN(n750) );
  NOR2_X1 U831 ( .A1(G1981), .A2(G305), .ZN(n746) );
  XNOR2_X1 U832 ( .A(n746), .B(KEYINPUT24), .ZN(n747) );
  XNOR2_X1 U833 ( .A(n747), .B(KEYINPUT91), .ZN(n748) );
  NOR2_X1 U834 ( .A1(n757), .A2(n748), .ZN(n749) );
  NOR2_X1 U835 ( .A1(n750), .A2(n749), .ZN(n764) );
  NOR2_X1 U836 ( .A1(G1971), .A2(G303), .ZN(n751) );
  NOR2_X1 U837 ( .A1(G1976), .A2(G288), .ZN(n966) );
  NOR2_X1 U838 ( .A1(n751), .A2(n966), .ZN(n752) );
  NAND2_X1 U839 ( .A1(n753), .A2(n752), .ZN(n755) );
  NAND2_X1 U840 ( .A1(G1976), .A2(G288), .ZN(n967) );
  INV_X1 U841 ( .A(n967), .ZN(n754) );
  AND2_X1 U842 ( .A1(n755), .A2(n516), .ZN(n756) );
  NOR2_X1 U843 ( .A1(KEYINPUT33), .A2(n756), .ZN(n760) );
  NAND2_X1 U844 ( .A1(n966), .A2(KEYINPUT33), .ZN(n758) );
  NOR2_X1 U845 ( .A1(n758), .A2(n757), .ZN(n759) );
  NOR2_X1 U846 ( .A1(n760), .A2(n759), .ZN(n762) );
  XNOR2_X1 U847 ( .A(KEYINPUT101), .B(G1981), .ZN(n761) );
  XNOR2_X1 U848 ( .A(n761), .B(G305), .ZN(n959) );
  NAND2_X1 U849 ( .A1(n762), .A2(n959), .ZN(n763) );
  NAND2_X1 U850 ( .A1(n764), .A2(n763), .ZN(n797) );
  XOR2_X1 U851 ( .A(n822), .B(KEYINPUT37), .Z(n805) );
  NAND2_X1 U852 ( .A1(G140), .A2(n875), .ZN(n766) );
  NAND2_X1 U853 ( .A1(G104), .A2(n877), .ZN(n765) );
  NAND2_X1 U854 ( .A1(n766), .A2(n765), .ZN(n767) );
  XNOR2_X1 U855 ( .A(KEYINPUT34), .B(n767), .ZN(n772) );
  NAND2_X1 U856 ( .A1(G116), .A2(n870), .ZN(n769) );
  NAND2_X1 U857 ( .A1(G128), .A2(n871), .ZN(n768) );
  NAND2_X1 U858 ( .A1(n769), .A2(n768), .ZN(n770) );
  XOR2_X1 U859 ( .A(KEYINPUT35), .B(n770), .Z(n771) );
  NOR2_X1 U860 ( .A1(n772), .A2(n771), .ZN(n773) );
  XNOR2_X1 U861 ( .A(KEYINPUT36), .B(n773), .ZN(n847) );
  NOR2_X1 U862 ( .A1(n805), .A2(n847), .ZN(n928) );
  NOR2_X1 U863 ( .A1(n775), .A2(n774), .ZN(n807) );
  NAND2_X1 U864 ( .A1(n928), .A2(n807), .ZN(n776) );
  XOR2_X1 U865 ( .A(n776), .B(KEYINPUT88), .Z(n802) );
  XOR2_X1 U866 ( .A(KEYINPUT90), .B(KEYINPUT38), .Z(n778) );
  NAND2_X1 U867 ( .A1(G105), .A2(n877), .ZN(n777) );
  XNOR2_X1 U868 ( .A(n778), .B(n777), .ZN(n783) );
  NAND2_X1 U869 ( .A1(G117), .A2(n870), .ZN(n780) );
  NAND2_X1 U870 ( .A1(G129), .A2(n871), .ZN(n779) );
  NAND2_X1 U871 ( .A1(n780), .A2(n779), .ZN(n781) );
  XOR2_X1 U872 ( .A(KEYINPUT89), .B(n781), .Z(n782) );
  NOR2_X1 U873 ( .A1(n783), .A2(n782), .ZN(n785) );
  NAND2_X1 U874 ( .A1(n875), .A2(G141), .ZN(n784) );
  NAND2_X1 U875 ( .A1(n785), .A2(n784), .ZN(n867) );
  AND2_X1 U876 ( .A1(n867), .A2(G1996), .ZN(n915) );
  NAND2_X1 U877 ( .A1(G107), .A2(n870), .ZN(n787) );
  NAND2_X1 U878 ( .A1(G131), .A2(n875), .ZN(n786) );
  NAND2_X1 U879 ( .A1(n787), .A2(n786), .ZN(n791) );
  NAND2_X1 U880 ( .A1(G119), .A2(n871), .ZN(n789) );
  NAND2_X1 U881 ( .A1(G95), .A2(n877), .ZN(n788) );
  NAND2_X1 U882 ( .A1(n789), .A2(n788), .ZN(n790) );
  OR2_X1 U883 ( .A1(n791), .A2(n790), .ZN(n866) );
  AND2_X1 U884 ( .A1(n866), .A2(G1991), .ZN(n909) );
  OR2_X1 U885 ( .A1(n915), .A2(n909), .ZN(n792) );
  NOR2_X1 U886 ( .A1(n802), .A2(n517), .ZN(n795) );
  XOR2_X1 U887 ( .A(G1986), .B(KEYINPUT87), .Z(n793) );
  XNOR2_X1 U888 ( .A(G290), .B(n793), .ZN(n975) );
  NAND2_X1 U889 ( .A1(n975), .A2(n807), .ZN(n794) );
  NAND2_X1 U890 ( .A1(n797), .A2(n796), .ZN(n810) );
  NOR2_X1 U891 ( .A1(G1996), .A2(n867), .ZN(n918) );
  NOR2_X1 U892 ( .A1(G1986), .A2(G290), .ZN(n798) );
  NOR2_X1 U893 ( .A1(G1991), .A2(n866), .ZN(n911) );
  NOR2_X1 U894 ( .A1(n798), .A2(n911), .ZN(n799) );
  NOR2_X1 U895 ( .A1(n517), .A2(n799), .ZN(n800) );
  NOR2_X1 U896 ( .A1(n918), .A2(n800), .ZN(n801) );
  XNOR2_X1 U897 ( .A(KEYINPUT39), .B(n801), .ZN(n804) );
  INV_X1 U898 ( .A(n802), .ZN(n803) );
  NAND2_X1 U899 ( .A1(n804), .A2(n803), .ZN(n806) );
  NAND2_X1 U900 ( .A1(n805), .A2(n847), .ZN(n927) );
  NAND2_X1 U901 ( .A1(n806), .A2(n927), .ZN(n808) );
  NAND2_X1 U902 ( .A1(n808), .A2(n807), .ZN(n809) );
  NAND2_X1 U903 ( .A1(n810), .A2(n809), .ZN(n811) );
  XNOR2_X1 U904 ( .A(KEYINPUT40), .B(n811), .ZN(G329) );
  NAND2_X1 U905 ( .A1(G2106), .A2(n907), .ZN(G217) );
  AND2_X1 U906 ( .A1(G15), .A2(G2), .ZN(n812) );
  NAND2_X1 U907 ( .A1(G661), .A2(n812), .ZN(G259) );
  NAND2_X1 U908 ( .A1(G1), .A2(G3), .ZN(n814) );
  NAND2_X1 U909 ( .A1(n814), .A2(n813), .ZN(n815) );
  XNOR2_X1 U910 ( .A(n815), .B(KEYINPUT104), .ZN(G188) );
  XNOR2_X1 U911 ( .A(G96), .B(KEYINPUT105), .ZN(G221) );
  NOR2_X1 U912 ( .A1(n817), .A2(n816), .ZN(G325) );
  XOR2_X1 U913 ( .A(KEYINPUT106), .B(G325), .Z(G261) );
  INV_X1 U915 ( .A(G120), .ZN(G236) );
  INV_X1 U916 ( .A(G108), .ZN(G238) );
  INV_X1 U917 ( .A(G69), .ZN(G235) );
  INV_X1 U918 ( .A(G301), .ZN(G171) );
  INV_X1 U919 ( .A(n818), .ZN(G319) );
  XNOR2_X1 U920 ( .A(n819), .B(G2096), .ZN(n821) );
  XNOR2_X1 U921 ( .A(KEYINPUT42), .B(G2678), .ZN(n820) );
  XNOR2_X1 U922 ( .A(n821), .B(n820), .ZN(n826) );
  XOR2_X1 U923 ( .A(KEYINPUT43), .B(G2090), .Z(n824) );
  XOR2_X1 U924 ( .A(n822), .B(G2072), .Z(n823) );
  XNOR2_X1 U925 ( .A(n824), .B(n823), .ZN(n825) );
  XOR2_X1 U926 ( .A(n826), .B(n825), .Z(n828) );
  XNOR2_X1 U927 ( .A(G2084), .B(G2078), .ZN(n827) );
  XNOR2_X1 U928 ( .A(n828), .B(n827), .ZN(G227) );
  XOR2_X1 U929 ( .A(G1956), .B(G1961), .Z(n830) );
  XNOR2_X1 U930 ( .A(G1991), .B(G1986), .ZN(n829) );
  XNOR2_X1 U931 ( .A(n830), .B(n829), .ZN(n834) );
  XOR2_X1 U932 ( .A(G1966), .B(G1971), .Z(n832) );
  XNOR2_X1 U933 ( .A(G1981), .B(G1976), .ZN(n831) );
  XNOR2_X1 U934 ( .A(n832), .B(n831), .ZN(n833) );
  XOR2_X1 U935 ( .A(n834), .B(n833), .Z(n836) );
  XNOR2_X1 U936 ( .A(G2474), .B(KEYINPUT107), .ZN(n835) );
  XNOR2_X1 U937 ( .A(n836), .B(n835), .ZN(n837) );
  XNOR2_X1 U938 ( .A(KEYINPUT41), .B(n837), .ZN(n838) );
  XOR2_X1 U939 ( .A(n838), .B(G1996), .Z(G229) );
  NAND2_X1 U940 ( .A1(G112), .A2(n870), .ZN(n840) );
  NAND2_X1 U941 ( .A1(G136), .A2(n875), .ZN(n839) );
  NAND2_X1 U942 ( .A1(n840), .A2(n839), .ZN(n846) );
  NAND2_X1 U943 ( .A1(G100), .A2(n877), .ZN(n841) );
  XNOR2_X1 U944 ( .A(n841), .B(KEYINPUT108), .ZN(n844) );
  NAND2_X1 U945 ( .A1(G124), .A2(n871), .ZN(n842) );
  XNOR2_X1 U946 ( .A(n842), .B(KEYINPUT44), .ZN(n843) );
  NAND2_X1 U947 ( .A1(n844), .A2(n843), .ZN(n845) );
  NOR2_X1 U948 ( .A1(n846), .A2(n845), .ZN(G162) );
  XNOR2_X1 U949 ( .A(G162), .B(G164), .ZN(n848) );
  XNOR2_X1 U950 ( .A(n848), .B(n847), .ZN(n859) );
  NAND2_X1 U951 ( .A1(G118), .A2(n870), .ZN(n849) );
  XNOR2_X1 U952 ( .A(n849), .B(KEYINPUT110), .ZN(n852) );
  NAND2_X1 U953 ( .A1(G130), .A2(n871), .ZN(n850) );
  XOR2_X1 U954 ( .A(KEYINPUT109), .B(n850), .Z(n851) );
  NAND2_X1 U955 ( .A1(n852), .A2(n851), .ZN(n857) );
  NAND2_X1 U956 ( .A1(G142), .A2(n875), .ZN(n854) );
  NAND2_X1 U957 ( .A1(G106), .A2(n877), .ZN(n853) );
  NAND2_X1 U958 ( .A1(n854), .A2(n853), .ZN(n855) );
  XOR2_X1 U959 ( .A(KEYINPUT45), .B(n855), .Z(n856) );
  NOR2_X1 U960 ( .A1(n857), .A2(n856), .ZN(n858) );
  XOR2_X1 U961 ( .A(n859), .B(n858), .Z(n861) );
  XNOR2_X1 U962 ( .A(G160), .B(n908), .ZN(n860) );
  XNOR2_X1 U963 ( .A(n861), .B(n860), .ZN(n865) );
  XOR2_X1 U964 ( .A(KEYINPUT114), .B(KEYINPUT48), .Z(n863) );
  XNOR2_X1 U965 ( .A(KEYINPUT46), .B(KEYINPUT115), .ZN(n862) );
  XNOR2_X1 U966 ( .A(n863), .B(n862), .ZN(n864) );
  XOR2_X1 U967 ( .A(n865), .B(n864), .Z(n869) );
  XNOR2_X1 U968 ( .A(n867), .B(n866), .ZN(n868) );
  XNOR2_X1 U969 ( .A(n869), .B(n868), .ZN(n884) );
  NAND2_X1 U970 ( .A1(G115), .A2(n870), .ZN(n873) );
  NAND2_X1 U971 ( .A1(G127), .A2(n871), .ZN(n872) );
  NAND2_X1 U972 ( .A1(n873), .A2(n872), .ZN(n874) );
  XNOR2_X1 U973 ( .A(KEYINPUT47), .B(n874), .ZN(n882) );
  NAND2_X1 U974 ( .A1(G139), .A2(n875), .ZN(n876) );
  XOR2_X1 U975 ( .A(KEYINPUT112), .B(n876), .Z(n880) );
  NAND2_X1 U976 ( .A1(G103), .A2(n877), .ZN(n878) );
  XNOR2_X1 U977 ( .A(KEYINPUT111), .B(n878), .ZN(n879) );
  NOR2_X1 U978 ( .A1(n880), .A2(n879), .ZN(n881) );
  NAND2_X1 U979 ( .A1(n882), .A2(n881), .ZN(n883) );
  XNOR2_X1 U980 ( .A(KEYINPUT113), .B(n883), .ZN(n922) );
  XNOR2_X1 U981 ( .A(n884), .B(n922), .ZN(n885) );
  NOR2_X1 U982 ( .A1(G37), .A2(n885), .ZN(G395) );
  XNOR2_X1 U983 ( .A(n978), .B(KEYINPUT116), .ZN(n887) );
  XOR2_X1 U984 ( .A(G301), .B(n962), .Z(n886) );
  XNOR2_X1 U985 ( .A(n887), .B(n886), .ZN(n890) );
  XNOR2_X1 U986 ( .A(n888), .B(G286), .ZN(n889) );
  XNOR2_X1 U987 ( .A(n890), .B(n889), .ZN(n891) );
  NOR2_X1 U988 ( .A1(G37), .A2(n891), .ZN(G397) );
  XOR2_X1 U989 ( .A(G2451), .B(G2430), .Z(n893) );
  XNOR2_X1 U990 ( .A(G2438), .B(G2443), .ZN(n892) );
  XNOR2_X1 U991 ( .A(n893), .B(n892), .ZN(n899) );
  XOR2_X1 U992 ( .A(G2435), .B(G2454), .Z(n895) );
  XNOR2_X1 U993 ( .A(G1348), .B(G1341), .ZN(n894) );
  XNOR2_X1 U994 ( .A(n895), .B(n894), .ZN(n897) );
  XOR2_X1 U995 ( .A(G2446), .B(G2427), .Z(n896) );
  XNOR2_X1 U996 ( .A(n897), .B(n896), .ZN(n898) );
  XOR2_X1 U997 ( .A(n899), .B(n898), .Z(n900) );
  NAND2_X1 U998 ( .A1(G14), .A2(n900), .ZN(n906) );
  NAND2_X1 U999 ( .A1(G319), .A2(n906), .ZN(n903) );
  NOR2_X1 U1000 ( .A1(G227), .A2(G229), .ZN(n901) );
  XNOR2_X1 U1001 ( .A(KEYINPUT49), .B(n901), .ZN(n902) );
  NOR2_X1 U1002 ( .A1(n903), .A2(n902), .ZN(n905) );
  NOR2_X1 U1003 ( .A1(G395), .A2(G397), .ZN(n904) );
  NAND2_X1 U1004 ( .A1(n905), .A2(n904), .ZN(G225) );
  INV_X1 U1005 ( .A(G225), .ZN(G308) );
  INV_X1 U1006 ( .A(n906), .ZN(G401) );
  INV_X1 U1007 ( .A(n907), .ZN(G223) );
  XNOR2_X1 U1008 ( .A(KEYINPUT127), .B(KEYINPUT62), .ZN(n1019) );
  INV_X1 U1009 ( .A(KEYINPUT55), .ZN(n957) );
  NOR2_X1 U1010 ( .A1(n909), .A2(n908), .ZN(n913) );
  XOR2_X1 U1011 ( .A(G160), .B(G2084), .Z(n910) );
  NOR2_X1 U1012 ( .A1(n911), .A2(n910), .ZN(n912) );
  NAND2_X1 U1013 ( .A1(n913), .A2(n912), .ZN(n914) );
  NOR2_X1 U1014 ( .A1(n915), .A2(n914), .ZN(n921) );
  XNOR2_X1 U1015 ( .A(G2090), .B(G162), .ZN(n916) );
  XNOR2_X1 U1016 ( .A(n916), .B(KEYINPUT117), .ZN(n917) );
  NOR2_X1 U1017 ( .A1(n918), .A2(n917), .ZN(n919) );
  XOR2_X1 U1018 ( .A(KEYINPUT51), .B(n919), .Z(n920) );
  NAND2_X1 U1019 ( .A1(n921), .A2(n920), .ZN(n933) );
  XNOR2_X1 U1020 ( .A(n923), .B(n922), .ZN(n925) );
  XOR2_X1 U1021 ( .A(G164), .B(G2078), .Z(n924) );
  NOR2_X1 U1022 ( .A1(n925), .A2(n924), .ZN(n926) );
  XNOR2_X1 U1023 ( .A(KEYINPUT50), .B(n926), .ZN(n931) );
  INV_X1 U1024 ( .A(n927), .ZN(n929) );
  NOR2_X1 U1025 ( .A1(n929), .A2(n928), .ZN(n930) );
  NAND2_X1 U1026 ( .A1(n931), .A2(n930), .ZN(n932) );
  NOR2_X1 U1027 ( .A1(n933), .A2(n932), .ZN(n934) );
  XNOR2_X1 U1028 ( .A(KEYINPUT52), .B(n934), .ZN(n935) );
  NAND2_X1 U1029 ( .A1(n957), .A2(n935), .ZN(n936) );
  NAND2_X1 U1030 ( .A1(n936), .A2(G29), .ZN(n1017) );
  XOR2_X1 U1031 ( .A(G2072), .B(G33), .Z(n938) );
  XOR2_X1 U1032 ( .A(G1996), .B(G32), .Z(n937) );
  NAND2_X1 U1033 ( .A1(n938), .A2(n937), .ZN(n948) );
  XNOR2_X1 U1034 ( .A(G25), .B(G1991), .ZN(n939) );
  XNOR2_X1 U1035 ( .A(n939), .B(KEYINPUT119), .ZN(n946) );
  XOR2_X1 U1036 ( .A(G26), .B(G2067), .Z(n940) );
  NAND2_X1 U1037 ( .A1(n940), .A2(G28), .ZN(n944) );
  XNOR2_X1 U1038 ( .A(G27), .B(n941), .ZN(n942) );
  XNOR2_X1 U1039 ( .A(KEYINPUT120), .B(n942), .ZN(n943) );
  NOR2_X1 U1040 ( .A1(n944), .A2(n943), .ZN(n945) );
  NAND2_X1 U1041 ( .A1(n946), .A2(n945), .ZN(n947) );
  NOR2_X1 U1042 ( .A1(n948), .A2(n947), .ZN(n949) );
  XOR2_X1 U1043 ( .A(KEYINPUT53), .B(n949), .Z(n952) );
  XOR2_X1 U1044 ( .A(KEYINPUT54), .B(G34), .Z(n950) );
  XNOR2_X1 U1045 ( .A(G2084), .B(n950), .ZN(n951) );
  NAND2_X1 U1046 ( .A1(n952), .A2(n951), .ZN(n955) );
  XNOR2_X1 U1047 ( .A(KEYINPUT118), .B(G2090), .ZN(n953) );
  XNOR2_X1 U1048 ( .A(G35), .B(n953), .ZN(n954) );
  NOR2_X1 U1049 ( .A1(n955), .A2(n954), .ZN(n956) );
  XNOR2_X1 U1050 ( .A(n957), .B(n956), .ZN(n958) );
  NOR2_X1 U1051 ( .A1(G29), .A2(n958), .ZN(n1013) );
  INV_X1 U1052 ( .A(G16), .ZN(n1009) );
  XOR2_X1 U1053 ( .A(n1009), .B(KEYINPUT56), .Z(n984) );
  XNOR2_X1 U1054 ( .A(G1966), .B(G168), .ZN(n960) );
  NAND2_X1 U1055 ( .A1(n960), .A2(n959), .ZN(n961) );
  XNOR2_X1 U1056 ( .A(n961), .B(KEYINPUT57), .ZN(n982) );
  XNOR2_X1 U1057 ( .A(n962), .B(G1348), .ZN(n964) );
  XOR2_X1 U1058 ( .A(G301), .B(G1961), .Z(n963) );
  NAND2_X1 U1059 ( .A1(n964), .A2(n963), .ZN(n965) );
  XNOR2_X1 U1060 ( .A(KEYINPUT121), .B(n965), .ZN(n977) );
  XOR2_X1 U1061 ( .A(G1971), .B(G303), .Z(n973) );
  XOR2_X1 U1062 ( .A(n966), .B(KEYINPUT122), .Z(n968) );
  NAND2_X1 U1063 ( .A1(n968), .A2(n967), .ZN(n971) );
  XNOR2_X1 U1064 ( .A(G1956), .B(n969), .ZN(n970) );
  NOR2_X1 U1065 ( .A1(n971), .A2(n970), .ZN(n972) );
  NAND2_X1 U1066 ( .A1(n973), .A2(n972), .ZN(n974) );
  NOR2_X1 U1067 ( .A1(n975), .A2(n974), .ZN(n976) );
  NAND2_X1 U1068 ( .A1(n977), .A2(n976), .ZN(n980) );
  XNOR2_X1 U1069 ( .A(G1341), .B(n978), .ZN(n979) );
  NOR2_X1 U1070 ( .A1(n980), .A2(n979), .ZN(n981) );
  NAND2_X1 U1071 ( .A1(n982), .A2(n981), .ZN(n983) );
  NAND2_X1 U1072 ( .A1(n984), .A2(n983), .ZN(n1011) );
  XOR2_X1 U1073 ( .A(G1961), .B(G5), .Z(n998) );
  XOR2_X1 U1074 ( .A(G1348), .B(KEYINPUT59), .Z(n985) );
  XNOR2_X1 U1075 ( .A(G4), .B(n985), .ZN(n987) );
  XNOR2_X1 U1076 ( .A(G6), .B(G1981), .ZN(n986) );
  NOR2_X1 U1077 ( .A1(n987), .A2(n986), .ZN(n991) );
  XNOR2_X1 U1078 ( .A(G1341), .B(G19), .ZN(n989) );
  XNOR2_X1 U1079 ( .A(G20), .B(G1956), .ZN(n988) );
  NOR2_X1 U1080 ( .A1(n989), .A2(n988), .ZN(n990) );
  NAND2_X1 U1081 ( .A1(n991), .A2(n990), .ZN(n992) );
  XNOR2_X1 U1082 ( .A(n992), .B(KEYINPUT123), .ZN(n993) );
  XOR2_X1 U1083 ( .A(KEYINPUT60), .B(n993), .Z(n995) );
  XNOR2_X1 U1084 ( .A(G1966), .B(G21), .ZN(n994) );
  NOR2_X1 U1085 ( .A1(n995), .A2(n994), .ZN(n996) );
  XNOR2_X1 U1086 ( .A(KEYINPUT124), .B(n996), .ZN(n997) );
  NAND2_X1 U1087 ( .A1(n998), .A2(n997), .ZN(n1006) );
  XOR2_X1 U1088 ( .A(G1986), .B(G24), .Z(n1002) );
  XNOR2_X1 U1089 ( .A(G1976), .B(G23), .ZN(n1000) );
  XNOR2_X1 U1090 ( .A(G1971), .B(G22), .ZN(n999) );
  NOR2_X1 U1091 ( .A1(n1000), .A2(n999), .ZN(n1001) );
  NAND2_X1 U1092 ( .A1(n1002), .A2(n1001), .ZN(n1003) );
  XOR2_X1 U1093 ( .A(KEYINPUT125), .B(n1003), .Z(n1004) );
  XNOR2_X1 U1094 ( .A(KEYINPUT58), .B(n1004), .ZN(n1005) );
  NOR2_X1 U1095 ( .A1(n1006), .A2(n1005), .ZN(n1007) );
  XNOR2_X1 U1096 ( .A(KEYINPUT61), .B(n1007), .ZN(n1008) );
  NAND2_X1 U1097 ( .A1(n1009), .A2(n1008), .ZN(n1010) );
  NAND2_X1 U1098 ( .A1(n1011), .A2(n1010), .ZN(n1012) );
  NOR2_X1 U1099 ( .A1(n1013), .A2(n1012), .ZN(n1014) );
  NAND2_X1 U1100 ( .A1(G11), .A2(n1014), .ZN(n1015) );
  XOR2_X1 U1101 ( .A(KEYINPUT126), .B(n1015), .Z(n1016) );
  NAND2_X1 U1102 ( .A1(n1017), .A2(n1016), .ZN(n1018) );
  XOR2_X1 U1103 ( .A(n1019), .B(n1018), .Z(G150) );
  INV_X1 U1104 ( .A(G150), .ZN(G311) );
endmodule

