

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601,
         n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612,
         n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623,
         n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634,
         n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645,
         n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656,
         n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667,
         n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678,
         n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689,
         n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700,
         n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711,
         n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722,
         n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733,
         n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744,
         n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, n755,
         n756, n757, n758, n759, n760, n761, n762, n763, n764, n765, n766,
         n767, n768, n769, n770, n771, n772, n773, n774, n775, n776, n777,
         n778, n779, n780, n781, n782, n783, n784, n785, n786, n787, n788,
         n789, n790, n791, n792, n793, n794, n795, n796, n797, n798, n799,
         n800, n801, n802, n803, n804, n805, n806, n807, n808, n809, n810,
         n811, n812, n813, n814, n815, n816, n817, n818, n819, n820, n821,
         n822, n823, n824, n825, n826, n827, n828, n829, n830, n831, n832,
         n833, n834, n835, n836, n837, n838, n839, n840, n841, n842, n843,
         n844, n845, n846, n847, n848, n849, n850, n851, n852, n853, n854,
         n855, n856, n857, n858, n859, n860, n861, n862, n863, n864, n865,
         n866, n867, n868, n869, n870, n871, n872, n873, n874, n875, n876,
         n877, n878, n879, n880, n881, n882, n883, n884, n885, n886, n887,
         n888, n889, n890, n891, n892, n893, n894, n895, n896, n897, n898,
         n899, n900, n901, n902, n903, n904, n905, n906, n907, n908, n909,
         n910, n911, n912, n913, n914, n915, n916, n917, n918, n919, n920,
         n921, n922, n923, n924, n925, n926, n927, n928, n929, n930, n931,
         n932, n933, n934, n935, n936, n937, n938, n939, n940, n941, n942,
         n943, n944, n945, n946, n947, n948, n949, n950, n951, n952, n953,
         n954, n955, n956, n957, n958, n959, n960, n961, n962, n963, n964,
         n965, n966, n967, n968, n969, n970, n971, n972, n973, n974, n975,
         n976, n977, n978, n979, n980, n981, n982, n983, n984, n985, n986,
         n987, n988, n989, n990, n991, n992, n993, n994, n995, n996, n997,
         n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007,
         n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017,
         n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027,
         n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NAND2_X2 U555 ( .A1(n675), .A2(n753), .ZN(n726) );
  OR2_X1 U556 ( .A1(n809), .A2(n808), .ZN(n810) );
  AND2_X1 U557 ( .A1(n558), .A2(n557), .ZN(n559) );
  INV_X1 U558 ( .A(n726), .ZN(n680) );
  BUF_X1 U559 ( .A(n680), .Z(n701) );
  INV_X1 U560 ( .A(KEYINPUT31), .ZN(n714) );
  XNOR2_X1 U561 ( .A(n714), .B(KEYINPUT94), .ZN(n715) );
  XNOR2_X1 U562 ( .A(n716), .B(n715), .ZN(n717) );
  NAND2_X1 U563 ( .A1(G160), .A2(G40), .ZN(n752) );
  NAND2_X1 U564 ( .A1(G8), .A2(n726), .ZN(n795) );
  NOR2_X1 U565 ( .A1(G651), .A2(n619), .ZN(n643) );
  NOR2_X1 U566 ( .A1(n531), .A2(n530), .ZN(G160) );
  XNOR2_X1 U567 ( .A(G2104), .B(KEYINPUT65), .ZN(n526) );
  NOR2_X1 U568 ( .A1(G2105), .A2(n526), .ZN(n885) );
  NAND2_X1 U569 ( .A1(G101), .A2(n885), .ZN(n521) );
  XOR2_X1 U570 ( .A(KEYINPUT23), .B(n521), .Z(n525) );
  NOR2_X1 U571 ( .A1(G2104), .A2(G2105), .ZN(n522) );
  XOR2_X2 U572 ( .A(KEYINPUT17), .B(n522), .Z(n882) );
  NAND2_X1 U573 ( .A1(n882), .A2(G137), .ZN(n523) );
  XOR2_X1 U574 ( .A(KEYINPUT67), .B(n523), .Z(n524) );
  NAND2_X1 U575 ( .A1(n525), .A2(n524), .ZN(n531) );
  AND2_X2 U576 ( .A1(n526), .A2(G2105), .ZN(n877) );
  NAND2_X1 U577 ( .A1(G125), .A2(n877), .ZN(n529) );
  NAND2_X1 U578 ( .A1(G2105), .A2(G2104), .ZN(n527) );
  XOR2_X2 U579 ( .A(KEYINPUT66), .B(n527), .Z(n878) );
  NAND2_X1 U580 ( .A1(G113), .A2(n878), .ZN(n528) );
  NAND2_X1 U581 ( .A1(n529), .A2(n528), .ZN(n530) );
  AND2_X1 U582 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U583 ( .A(G651), .ZN(n536) );
  NOR2_X1 U584 ( .A1(G543), .A2(n536), .ZN(n532) );
  XOR2_X1 U585 ( .A(KEYINPUT1), .B(n532), .Z(n644) );
  NAND2_X1 U586 ( .A1(n644), .A2(G65), .ZN(n535) );
  NOR2_X1 U587 ( .A1(G651), .A2(G543), .ZN(n533) );
  XNOR2_X1 U588 ( .A(n533), .B(KEYINPUT64), .ZN(n639) );
  NAND2_X1 U589 ( .A1(G91), .A2(n639), .ZN(n534) );
  NAND2_X1 U590 ( .A1(n535), .A2(n534), .ZN(n540) );
  XOR2_X1 U591 ( .A(G543), .B(KEYINPUT0), .Z(n619) );
  NAND2_X1 U592 ( .A1(G53), .A2(n643), .ZN(n538) );
  NOR2_X1 U593 ( .A1(n619), .A2(n536), .ZN(n638) );
  NAND2_X1 U594 ( .A1(G78), .A2(n638), .ZN(n537) );
  NAND2_X1 U595 ( .A1(n538), .A2(n537), .ZN(n539) );
  NOR2_X1 U596 ( .A1(n540), .A2(n539), .ZN(n694) );
  INV_X1 U597 ( .A(n694), .ZN(G299) );
  INV_X1 U598 ( .A(G57), .ZN(G237) );
  INV_X1 U599 ( .A(G132), .ZN(G219) );
  NAND2_X1 U600 ( .A1(G89), .A2(n639), .ZN(n541) );
  XNOR2_X1 U601 ( .A(n541), .B(KEYINPUT4), .ZN(n543) );
  NAND2_X1 U602 ( .A1(G76), .A2(n638), .ZN(n542) );
  NAND2_X1 U603 ( .A1(n543), .A2(n542), .ZN(n544) );
  XNOR2_X1 U604 ( .A(n544), .B(KEYINPUT5), .ZN(n549) );
  NAND2_X1 U605 ( .A1(G51), .A2(n643), .ZN(n546) );
  NAND2_X1 U606 ( .A1(G63), .A2(n644), .ZN(n545) );
  NAND2_X1 U607 ( .A1(n546), .A2(n545), .ZN(n547) );
  XOR2_X1 U608 ( .A(KEYINPUT6), .B(n547), .Z(n548) );
  NAND2_X1 U609 ( .A1(n549), .A2(n548), .ZN(n550) );
  XNOR2_X1 U610 ( .A(n550), .B(KEYINPUT7), .ZN(G168) );
  XOR2_X1 U611 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U612 ( .A1(n877), .A2(G126), .ZN(n551) );
  XNOR2_X1 U613 ( .A(n551), .B(KEYINPUT80), .ZN(n553) );
  NAND2_X1 U614 ( .A1(G114), .A2(n878), .ZN(n552) );
  NAND2_X1 U615 ( .A1(n553), .A2(n552), .ZN(n554) );
  XNOR2_X1 U616 ( .A(n554), .B(KEYINPUT81), .ZN(n558) );
  NAND2_X1 U617 ( .A1(G138), .A2(n882), .ZN(n556) );
  NAND2_X1 U618 ( .A1(G102), .A2(n885), .ZN(n555) );
  AND2_X1 U619 ( .A1(n556), .A2(n555), .ZN(n557) );
  XNOR2_X1 U620 ( .A(KEYINPUT82), .B(n559), .ZN(G164) );
  NAND2_X1 U621 ( .A1(G7), .A2(G661), .ZN(n560) );
  XNOR2_X1 U622 ( .A(n560), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U623 ( .A(G223), .ZN(n829) );
  NAND2_X1 U624 ( .A1(n829), .A2(G567), .ZN(n561) );
  XOR2_X1 U625 ( .A(KEYINPUT11), .B(n561), .Z(G234) );
  NAND2_X1 U626 ( .A1(G56), .A2(n644), .ZN(n562) );
  XOR2_X1 U627 ( .A(KEYINPUT14), .B(n562), .Z(n568) );
  NAND2_X1 U628 ( .A1(G81), .A2(n639), .ZN(n563) );
  XNOR2_X1 U629 ( .A(n563), .B(KEYINPUT12), .ZN(n565) );
  NAND2_X1 U630 ( .A1(G68), .A2(n638), .ZN(n564) );
  NAND2_X1 U631 ( .A1(n565), .A2(n564), .ZN(n566) );
  XOR2_X1 U632 ( .A(KEYINPUT13), .B(n566), .Z(n567) );
  NOR2_X1 U633 ( .A1(n568), .A2(n567), .ZN(n570) );
  NAND2_X1 U634 ( .A1(n643), .A2(G43), .ZN(n569) );
  NAND2_X1 U635 ( .A1(n570), .A2(n569), .ZN(n989) );
  INV_X1 U636 ( .A(G860), .ZN(n607) );
  OR2_X1 U637 ( .A1(n989), .A2(n607), .ZN(G153) );
  NAND2_X1 U638 ( .A1(G64), .A2(n644), .ZN(n571) );
  XNOR2_X1 U639 ( .A(n571), .B(KEYINPUT69), .ZN(n576) );
  NAND2_X1 U640 ( .A1(n638), .A2(G77), .ZN(n573) );
  NAND2_X1 U641 ( .A1(G90), .A2(n639), .ZN(n572) );
  NAND2_X1 U642 ( .A1(n573), .A2(n572), .ZN(n574) );
  XOR2_X1 U643 ( .A(KEYINPUT9), .B(n574), .Z(n575) );
  NOR2_X1 U644 ( .A1(n576), .A2(n575), .ZN(n578) );
  NAND2_X1 U645 ( .A1(n643), .A2(G52), .ZN(n577) );
  NAND2_X1 U646 ( .A1(n578), .A2(n577), .ZN(G301) );
  NAND2_X1 U647 ( .A1(G868), .A2(G301), .ZN(n587) );
  NAND2_X1 U648 ( .A1(n644), .A2(G66), .ZN(n580) );
  NAND2_X1 U649 ( .A1(G92), .A2(n639), .ZN(n579) );
  NAND2_X1 U650 ( .A1(n580), .A2(n579), .ZN(n584) );
  NAND2_X1 U651 ( .A1(G54), .A2(n643), .ZN(n582) );
  NAND2_X1 U652 ( .A1(G79), .A2(n638), .ZN(n581) );
  NAND2_X1 U653 ( .A1(n582), .A2(n581), .ZN(n583) );
  NOR2_X1 U654 ( .A1(n584), .A2(n583), .ZN(n585) );
  XOR2_X1 U655 ( .A(KEYINPUT15), .B(n585), .Z(n899) );
  INV_X1 U656 ( .A(n899), .ZN(n975) );
  INV_X1 U657 ( .A(G868), .ZN(n588) );
  NAND2_X1 U658 ( .A1(n975), .A2(n588), .ZN(n586) );
  NAND2_X1 U659 ( .A1(n587), .A2(n586), .ZN(G284) );
  NOR2_X1 U660 ( .A1(G286), .A2(n588), .ZN(n590) );
  NOR2_X1 U661 ( .A1(G868), .A2(G299), .ZN(n589) );
  NOR2_X1 U662 ( .A1(n590), .A2(n589), .ZN(G297) );
  NAND2_X1 U663 ( .A1(n607), .A2(G559), .ZN(n591) );
  NAND2_X1 U664 ( .A1(n591), .A2(n899), .ZN(n592) );
  XNOR2_X1 U665 ( .A(n592), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U666 ( .A1(G868), .A2(n989), .ZN(n595) );
  NAND2_X1 U667 ( .A1(G868), .A2(n899), .ZN(n593) );
  NOR2_X1 U668 ( .A1(G559), .A2(n593), .ZN(n594) );
  NOR2_X1 U669 ( .A1(n595), .A2(n594), .ZN(G282) );
  NAND2_X1 U670 ( .A1(G123), .A2(n877), .ZN(n596) );
  XNOR2_X1 U671 ( .A(n596), .B(KEYINPUT18), .ZN(n599) );
  NAND2_X1 U672 ( .A1(n878), .A2(G111), .ZN(n597) );
  XOR2_X1 U673 ( .A(KEYINPUT71), .B(n597), .Z(n598) );
  NAND2_X1 U674 ( .A1(n599), .A2(n598), .ZN(n603) );
  NAND2_X1 U675 ( .A1(G135), .A2(n882), .ZN(n601) );
  NAND2_X1 U676 ( .A1(G99), .A2(n885), .ZN(n600) );
  NAND2_X1 U677 ( .A1(n601), .A2(n600), .ZN(n602) );
  NOR2_X1 U678 ( .A1(n603), .A2(n602), .ZN(n930) );
  XNOR2_X1 U679 ( .A(G2096), .B(n930), .ZN(n605) );
  INV_X1 U680 ( .A(G2100), .ZN(n604) );
  NAND2_X1 U681 ( .A1(n605), .A2(n604), .ZN(G156) );
  NAND2_X1 U682 ( .A1(G559), .A2(n899), .ZN(n606) );
  XOR2_X1 U683 ( .A(n989), .B(n606), .Z(n657) );
  NAND2_X1 U684 ( .A1(n607), .A2(n657), .ZN(n615) );
  NAND2_X1 U685 ( .A1(n638), .A2(G80), .ZN(n609) );
  NAND2_X1 U686 ( .A1(G93), .A2(n639), .ZN(n608) );
  NAND2_X1 U687 ( .A1(n609), .A2(n608), .ZN(n614) );
  NAND2_X1 U688 ( .A1(n643), .A2(G55), .ZN(n610) );
  XNOR2_X1 U689 ( .A(n610), .B(KEYINPUT72), .ZN(n612) );
  NAND2_X1 U690 ( .A1(G67), .A2(n644), .ZN(n611) );
  NAND2_X1 U691 ( .A1(n612), .A2(n611), .ZN(n613) );
  NOR2_X1 U692 ( .A1(n614), .A2(n613), .ZN(n659) );
  XOR2_X1 U693 ( .A(n615), .B(n659), .Z(G145) );
  NAND2_X1 U694 ( .A1(G49), .A2(n643), .ZN(n617) );
  NAND2_X1 U695 ( .A1(G74), .A2(G651), .ZN(n616) );
  NAND2_X1 U696 ( .A1(n617), .A2(n616), .ZN(n618) );
  NOR2_X1 U697 ( .A1(n644), .A2(n618), .ZN(n622) );
  NAND2_X1 U698 ( .A1(G87), .A2(n619), .ZN(n620) );
  XOR2_X1 U699 ( .A(KEYINPUT73), .B(n620), .Z(n621) );
  NAND2_X1 U700 ( .A1(n622), .A2(n621), .ZN(G288) );
  NAND2_X1 U701 ( .A1(n644), .A2(G61), .ZN(n623) );
  XNOR2_X1 U702 ( .A(n623), .B(KEYINPUT74), .ZN(n630) );
  NAND2_X1 U703 ( .A1(n643), .A2(G48), .ZN(n625) );
  NAND2_X1 U704 ( .A1(G86), .A2(n639), .ZN(n624) );
  NAND2_X1 U705 ( .A1(n625), .A2(n624), .ZN(n628) );
  NAND2_X1 U706 ( .A1(G73), .A2(n638), .ZN(n626) );
  XOR2_X1 U707 ( .A(KEYINPUT2), .B(n626), .Z(n627) );
  NOR2_X1 U708 ( .A1(n628), .A2(n627), .ZN(n629) );
  NAND2_X1 U709 ( .A1(n630), .A2(n629), .ZN(G305) );
  NAND2_X1 U710 ( .A1(n644), .A2(G62), .ZN(n632) );
  NAND2_X1 U711 ( .A1(G88), .A2(n639), .ZN(n631) );
  NAND2_X1 U712 ( .A1(n632), .A2(n631), .ZN(n636) );
  NAND2_X1 U713 ( .A1(G50), .A2(n643), .ZN(n634) );
  NAND2_X1 U714 ( .A1(G75), .A2(n638), .ZN(n633) );
  NAND2_X1 U715 ( .A1(n634), .A2(n633), .ZN(n635) );
  NOR2_X1 U716 ( .A1(n636), .A2(n635), .ZN(n637) );
  XOR2_X1 U717 ( .A(KEYINPUT75), .B(n637), .Z(G166) );
  NAND2_X1 U718 ( .A1(n638), .A2(G72), .ZN(n641) );
  NAND2_X1 U719 ( .A1(G85), .A2(n639), .ZN(n640) );
  NAND2_X1 U720 ( .A1(n641), .A2(n640), .ZN(n642) );
  XOR2_X1 U721 ( .A(KEYINPUT68), .B(n642), .Z(n648) );
  NAND2_X1 U722 ( .A1(n643), .A2(G47), .ZN(n646) );
  NAND2_X1 U723 ( .A1(G60), .A2(n644), .ZN(n645) );
  AND2_X1 U724 ( .A1(n646), .A2(n645), .ZN(n647) );
  NAND2_X1 U725 ( .A1(n648), .A2(n647), .ZN(G290) );
  XNOR2_X1 U726 ( .A(n694), .B(n659), .ZN(n655) );
  XNOR2_X1 U727 ( .A(KEYINPUT77), .B(KEYINPUT78), .ZN(n650) );
  XNOR2_X1 U728 ( .A(G288), .B(KEYINPUT19), .ZN(n649) );
  XNOR2_X1 U729 ( .A(n650), .B(n649), .ZN(n651) );
  XNOR2_X1 U730 ( .A(KEYINPUT76), .B(n651), .ZN(n653) );
  XNOR2_X1 U731 ( .A(G305), .B(G166), .ZN(n652) );
  XNOR2_X1 U732 ( .A(n653), .B(n652), .ZN(n654) );
  XNOR2_X1 U733 ( .A(n655), .B(n654), .ZN(n656) );
  XNOR2_X1 U734 ( .A(n656), .B(G290), .ZN(n902) );
  XNOR2_X1 U735 ( .A(n657), .B(n902), .ZN(n658) );
  NAND2_X1 U736 ( .A1(n658), .A2(G868), .ZN(n661) );
  OR2_X1 U737 ( .A1(G868), .A2(n659), .ZN(n660) );
  NAND2_X1 U738 ( .A1(n661), .A2(n660), .ZN(G295) );
  NAND2_X1 U739 ( .A1(G2084), .A2(G2078), .ZN(n662) );
  XNOR2_X1 U740 ( .A(n662), .B(KEYINPUT20), .ZN(n663) );
  XNOR2_X1 U741 ( .A(n663), .B(KEYINPUT79), .ZN(n664) );
  NAND2_X1 U742 ( .A1(n664), .A2(G2090), .ZN(n665) );
  XNOR2_X1 U743 ( .A(KEYINPUT21), .B(n665), .ZN(n666) );
  NAND2_X1 U744 ( .A1(n666), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U745 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  XOR2_X1 U746 ( .A(KEYINPUT70), .B(G82), .Z(G220) );
  NOR2_X1 U747 ( .A1(G220), .A2(G219), .ZN(n667) );
  XOR2_X1 U748 ( .A(KEYINPUT22), .B(n667), .Z(n668) );
  NOR2_X1 U749 ( .A1(G218), .A2(n668), .ZN(n669) );
  NAND2_X1 U750 ( .A1(G96), .A2(n669), .ZN(n834) );
  NAND2_X1 U751 ( .A1(n834), .A2(G2106), .ZN(n673) );
  NAND2_X1 U752 ( .A1(G108), .A2(G120), .ZN(n670) );
  NOR2_X1 U753 ( .A1(G237), .A2(n670), .ZN(n671) );
  NAND2_X1 U754 ( .A1(G69), .A2(n671), .ZN(n835) );
  NAND2_X1 U755 ( .A1(n835), .A2(G567), .ZN(n672) );
  NAND2_X1 U756 ( .A1(n673), .A2(n672), .ZN(n836) );
  NAND2_X1 U757 ( .A1(G483), .A2(G661), .ZN(n674) );
  NOR2_X1 U758 ( .A1(n836), .A2(n674), .ZN(n832) );
  NAND2_X1 U759 ( .A1(n832), .A2(G36), .ZN(G176) );
  INV_X1 U760 ( .A(G166), .ZN(G303) );
  INV_X1 U761 ( .A(n752), .ZN(n675) );
  NOR2_X1 U762 ( .A1(G1384), .A2(G164), .ZN(n753) );
  NOR2_X1 U763 ( .A1(G1966), .A2(n795), .ZN(n720) );
  NAND2_X1 U764 ( .A1(n680), .A2(G2072), .ZN(n676) );
  XNOR2_X1 U765 ( .A(n676), .B(KEYINPUT27), .ZN(n678) );
  INV_X1 U766 ( .A(G1956), .ZN(n1012) );
  NOR2_X1 U767 ( .A1(n1012), .A2(n701), .ZN(n677) );
  NOR2_X1 U768 ( .A1(n678), .A2(n677), .ZN(n693) );
  NOR2_X1 U769 ( .A1(n694), .A2(n693), .ZN(n679) );
  XOR2_X1 U770 ( .A(n679), .B(KEYINPUT28), .Z(n698) );
  XNOR2_X1 U771 ( .A(G1996), .B(KEYINPUT90), .ZN(n955) );
  NAND2_X1 U772 ( .A1(n955), .A2(n680), .ZN(n681) );
  XNOR2_X1 U773 ( .A(n681), .B(KEYINPUT26), .ZN(n683) );
  NAND2_X1 U774 ( .A1(n726), .A2(G1341), .ZN(n682) );
  NAND2_X1 U775 ( .A1(n683), .A2(n682), .ZN(n684) );
  NOR2_X1 U776 ( .A1(n684), .A2(n989), .ZN(n690) );
  NAND2_X1 U777 ( .A1(n690), .A2(n899), .ZN(n689) );
  AND2_X1 U778 ( .A1(n701), .A2(G2067), .ZN(n685) );
  XNOR2_X1 U779 ( .A(n685), .B(KEYINPUT91), .ZN(n687) );
  NAND2_X1 U780 ( .A1(n726), .A2(G1348), .ZN(n686) );
  NAND2_X1 U781 ( .A1(n687), .A2(n686), .ZN(n688) );
  NAND2_X1 U782 ( .A1(n689), .A2(n688), .ZN(n692) );
  OR2_X1 U783 ( .A1(n899), .A2(n690), .ZN(n691) );
  NAND2_X1 U784 ( .A1(n692), .A2(n691), .ZN(n696) );
  NAND2_X1 U785 ( .A1(n694), .A2(n693), .ZN(n695) );
  NAND2_X1 U786 ( .A1(n696), .A2(n695), .ZN(n697) );
  NAND2_X1 U787 ( .A1(n698), .A2(n697), .ZN(n700) );
  XOR2_X1 U788 ( .A(KEYINPUT29), .B(KEYINPUT92), .Z(n699) );
  XNOR2_X1 U789 ( .A(n700), .B(n699), .ZN(n706) );
  NAND2_X1 U790 ( .A1(G1961), .A2(n726), .ZN(n703) );
  XOR2_X1 U791 ( .A(G2078), .B(KEYINPUT25), .Z(n956) );
  NAND2_X1 U792 ( .A1(n701), .A2(n956), .ZN(n702) );
  NAND2_X1 U793 ( .A1(n703), .A2(n702), .ZN(n707) );
  NOR2_X1 U794 ( .A1(G301), .A2(n707), .ZN(n704) );
  XNOR2_X1 U795 ( .A(n704), .B(KEYINPUT89), .ZN(n705) );
  NAND2_X1 U796 ( .A1(n706), .A2(n705), .ZN(n718) );
  NAND2_X1 U797 ( .A1(G301), .A2(n707), .ZN(n708) );
  XNOR2_X1 U798 ( .A(n708), .B(KEYINPUT93), .ZN(n713) );
  NOR2_X1 U799 ( .A1(G2084), .A2(n726), .ZN(n789) );
  NOR2_X1 U800 ( .A1(n789), .A2(n720), .ZN(n709) );
  NAND2_X1 U801 ( .A1(G8), .A2(n709), .ZN(n710) );
  XNOR2_X1 U802 ( .A(n710), .B(KEYINPUT30), .ZN(n711) );
  NOR2_X1 U803 ( .A1(n711), .A2(G168), .ZN(n712) );
  NOR2_X1 U804 ( .A1(n713), .A2(n712), .ZN(n716) );
  NAND2_X1 U805 ( .A1(n718), .A2(n717), .ZN(n724) );
  XNOR2_X1 U806 ( .A(KEYINPUT95), .B(n724), .ZN(n719) );
  NOR2_X1 U807 ( .A1(n720), .A2(n719), .ZN(n721) );
  XNOR2_X1 U808 ( .A(n721), .B(KEYINPUT96), .ZN(n791) );
  INV_X1 U809 ( .A(G1971), .ZN(n1004) );
  NAND2_X1 U810 ( .A1(G166), .A2(n1004), .ZN(n722) );
  AND2_X1 U811 ( .A1(n791), .A2(n722), .ZN(n738) );
  INV_X1 U812 ( .A(n722), .ZN(n736) );
  AND2_X1 U813 ( .A1(G286), .A2(G8), .ZN(n723) );
  NAND2_X1 U814 ( .A1(n724), .A2(n723), .ZN(n734) );
  INV_X1 U815 ( .A(G8), .ZN(n732) );
  NOR2_X1 U816 ( .A1(G1971), .A2(n795), .ZN(n725) );
  XNOR2_X1 U817 ( .A(KEYINPUT97), .B(n725), .ZN(n730) );
  NOR2_X1 U818 ( .A1(G2090), .A2(n726), .ZN(n727) );
  XNOR2_X1 U819 ( .A(KEYINPUT98), .B(n727), .ZN(n728) );
  NOR2_X1 U820 ( .A1(G166), .A2(n728), .ZN(n729) );
  NAND2_X1 U821 ( .A1(n730), .A2(n729), .ZN(n731) );
  OR2_X1 U822 ( .A1(n732), .A2(n731), .ZN(n733) );
  AND2_X1 U823 ( .A1(n734), .A2(n733), .ZN(n735) );
  XNOR2_X1 U824 ( .A(n735), .B(KEYINPUT32), .ZN(n796) );
  NOR2_X1 U825 ( .A1(n736), .A2(n796), .ZN(n737) );
  NOR2_X1 U826 ( .A1(n738), .A2(n737), .ZN(n739) );
  NOR2_X1 U827 ( .A1(G1976), .A2(G288), .ZN(n979) );
  NOR2_X1 U828 ( .A1(n739), .A2(n979), .ZN(n740) );
  NOR2_X1 U829 ( .A1(n795), .A2(n740), .ZN(n743) );
  NAND2_X1 U830 ( .A1(G1976), .A2(G288), .ZN(n980) );
  INV_X1 U831 ( .A(n980), .ZN(n741) );
  NOR2_X1 U832 ( .A1(n741), .A2(KEYINPUT99), .ZN(n742) );
  AND2_X1 U833 ( .A1(n743), .A2(n742), .ZN(n744) );
  NOR2_X1 U834 ( .A1(n744), .A2(KEYINPUT33), .ZN(n751) );
  INV_X1 U835 ( .A(KEYINPUT99), .ZN(n746) );
  NAND2_X1 U836 ( .A1(n979), .A2(KEYINPUT33), .ZN(n745) );
  NAND2_X1 U837 ( .A1(n746), .A2(n745), .ZN(n748) );
  NAND2_X1 U838 ( .A1(n979), .A2(KEYINPUT99), .ZN(n747) );
  NAND2_X1 U839 ( .A1(n748), .A2(n747), .ZN(n749) );
  NOR2_X1 U840 ( .A1(n795), .A2(n749), .ZN(n750) );
  NOR2_X1 U841 ( .A1(n751), .A2(n750), .ZN(n787) );
  XOR2_X1 U842 ( .A(G1981), .B(G305), .Z(n995) );
  NOR2_X1 U843 ( .A1(n753), .A2(n752), .ZN(n822) );
  XNOR2_X1 U844 ( .A(G2067), .B(KEYINPUT37), .ZN(n819) );
  XNOR2_X1 U845 ( .A(KEYINPUT85), .B(KEYINPUT36), .ZN(n765) );
  NAND2_X1 U846 ( .A1(G128), .A2(n877), .ZN(n755) );
  NAND2_X1 U847 ( .A1(G116), .A2(n878), .ZN(n754) );
  NAND2_X1 U848 ( .A1(n755), .A2(n754), .ZN(n756) );
  XNOR2_X1 U849 ( .A(KEYINPUT35), .B(n756), .ZN(n763) );
  XNOR2_X1 U850 ( .A(KEYINPUT34), .B(KEYINPUT84), .ZN(n761) );
  NAND2_X1 U851 ( .A1(n882), .A2(G140), .ZN(n759) );
  NAND2_X1 U852 ( .A1(n885), .A2(G104), .ZN(n757) );
  XOR2_X1 U853 ( .A(KEYINPUT83), .B(n757), .Z(n758) );
  NAND2_X1 U854 ( .A1(n759), .A2(n758), .ZN(n760) );
  XOR2_X1 U855 ( .A(n761), .B(n760), .Z(n762) );
  NAND2_X1 U856 ( .A1(n763), .A2(n762), .ZN(n764) );
  XNOR2_X1 U857 ( .A(n765), .B(n764), .ZN(n894) );
  NOR2_X1 U858 ( .A1(n819), .A2(n894), .ZN(n766) );
  XNOR2_X1 U859 ( .A(n766), .B(KEYINPUT86), .ZN(n946) );
  NAND2_X1 U860 ( .A1(n822), .A2(n946), .ZN(n817) );
  NAND2_X1 U861 ( .A1(G141), .A2(n882), .ZN(n768) );
  NAND2_X1 U862 ( .A1(G117), .A2(n878), .ZN(n767) );
  NAND2_X1 U863 ( .A1(n768), .A2(n767), .ZN(n771) );
  NAND2_X1 U864 ( .A1(n885), .A2(G105), .ZN(n769) );
  XOR2_X1 U865 ( .A(KEYINPUT38), .B(n769), .Z(n770) );
  NOR2_X1 U866 ( .A1(n771), .A2(n770), .ZN(n773) );
  NAND2_X1 U867 ( .A1(n877), .A2(G129), .ZN(n772) );
  NAND2_X1 U868 ( .A1(n773), .A2(n772), .ZN(n866) );
  NAND2_X1 U869 ( .A1(G1996), .A2(n866), .ZN(n781) );
  NAND2_X1 U870 ( .A1(G119), .A2(n877), .ZN(n775) );
  NAND2_X1 U871 ( .A1(G107), .A2(n878), .ZN(n774) );
  NAND2_X1 U872 ( .A1(n775), .A2(n774), .ZN(n779) );
  NAND2_X1 U873 ( .A1(G131), .A2(n882), .ZN(n777) );
  NAND2_X1 U874 ( .A1(G95), .A2(n885), .ZN(n776) );
  NAND2_X1 U875 ( .A1(n777), .A2(n776), .ZN(n778) );
  OR2_X1 U876 ( .A1(n779), .A2(n778), .ZN(n874) );
  NAND2_X1 U877 ( .A1(G1991), .A2(n874), .ZN(n780) );
  NAND2_X1 U878 ( .A1(n781), .A2(n780), .ZN(n934) );
  NAND2_X1 U879 ( .A1(n934), .A2(n822), .ZN(n782) );
  XNOR2_X1 U880 ( .A(n782), .B(KEYINPUT87), .ZN(n814) );
  INV_X1 U881 ( .A(n814), .ZN(n783) );
  NAND2_X1 U882 ( .A1(n817), .A2(n783), .ZN(n809) );
  INV_X1 U883 ( .A(n809), .ZN(n784) );
  AND2_X1 U884 ( .A1(n995), .A2(n784), .ZN(n785) );
  XNOR2_X1 U885 ( .A(G1986), .B(G290), .ZN(n991) );
  NAND2_X1 U886 ( .A1(n991), .A2(n822), .ZN(n788) );
  AND2_X1 U887 ( .A1(n785), .A2(n788), .ZN(n786) );
  NAND2_X1 U888 ( .A1(n787), .A2(n786), .ZN(n827) );
  INV_X1 U889 ( .A(n788), .ZN(n811) );
  NAND2_X1 U890 ( .A1(n789), .A2(G8), .ZN(n790) );
  NAND2_X1 U891 ( .A1(n791), .A2(n790), .ZN(n798) );
  NOR2_X1 U892 ( .A1(G1981), .A2(G305), .ZN(n792) );
  XOR2_X1 U893 ( .A(n792), .B(KEYINPUT24), .Z(n793) );
  NOR2_X1 U894 ( .A1(n795), .A2(n793), .ZN(n794) );
  XNOR2_X1 U895 ( .A(n794), .B(KEYINPUT88), .ZN(n801) );
  OR2_X1 U896 ( .A1(n801), .A2(n795), .ZN(n799) );
  AND2_X1 U897 ( .A1(n796), .A2(n799), .ZN(n797) );
  NAND2_X1 U898 ( .A1(n798), .A2(n797), .ZN(n807) );
  INV_X1 U899 ( .A(n799), .ZN(n805) );
  NOR2_X1 U900 ( .A1(G2090), .A2(G303), .ZN(n800) );
  NAND2_X1 U901 ( .A1(G8), .A2(n800), .ZN(n803) );
  INV_X1 U902 ( .A(n801), .ZN(n802) );
  AND2_X1 U903 ( .A1(n803), .A2(n802), .ZN(n804) );
  OR2_X1 U904 ( .A1(n805), .A2(n804), .ZN(n806) );
  AND2_X1 U905 ( .A1(n807), .A2(n806), .ZN(n808) );
  OR2_X1 U906 ( .A1(n811), .A2(n810), .ZN(n825) );
  NOR2_X1 U907 ( .A1(G1996), .A2(n866), .ZN(n926) );
  NOR2_X1 U908 ( .A1(G1986), .A2(G290), .ZN(n812) );
  NOR2_X1 U909 ( .A1(G1991), .A2(n874), .ZN(n931) );
  NOR2_X1 U910 ( .A1(n812), .A2(n931), .ZN(n813) );
  NOR2_X1 U911 ( .A1(n814), .A2(n813), .ZN(n815) );
  NOR2_X1 U912 ( .A1(n926), .A2(n815), .ZN(n816) );
  XNOR2_X1 U913 ( .A(n816), .B(KEYINPUT39), .ZN(n818) );
  NAND2_X1 U914 ( .A1(n818), .A2(n817), .ZN(n820) );
  NAND2_X1 U915 ( .A1(n894), .A2(n819), .ZN(n943) );
  NAND2_X1 U916 ( .A1(n820), .A2(n943), .ZN(n821) );
  NAND2_X1 U917 ( .A1(n822), .A2(n821), .ZN(n823) );
  XNOR2_X1 U918 ( .A(KEYINPUT100), .B(n823), .ZN(n824) );
  AND2_X1 U919 ( .A1(n825), .A2(n824), .ZN(n826) );
  NAND2_X1 U920 ( .A1(n827), .A2(n826), .ZN(n828) );
  XNOR2_X1 U921 ( .A(n828), .B(KEYINPUT40), .ZN(G329) );
  NAND2_X1 U922 ( .A1(G2106), .A2(n829), .ZN(G217) );
  AND2_X1 U923 ( .A1(G15), .A2(G2), .ZN(n830) );
  NAND2_X1 U924 ( .A1(G661), .A2(n830), .ZN(G259) );
  NAND2_X1 U925 ( .A1(G3), .A2(G1), .ZN(n831) );
  XNOR2_X1 U926 ( .A(KEYINPUT104), .B(n831), .ZN(n833) );
  NAND2_X1 U927 ( .A1(n833), .A2(n832), .ZN(G188) );
  XNOR2_X1 U928 ( .A(G120), .B(KEYINPUT105), .ZN(G236) );
  INV_X1 U930 ( .A(G108), .ZN(G238) );
  INV_X1 U931 ( .A(G96), .ZN(G221) );
  NOR2_X1 U932 ( .A1(n835), .A2(n834), .ZN(G325) );
  INV_X1 U933 ( .A(G325), .ZN(G261) );
  INV_X1 U934 ( .A(n836), .ZN(G319) );
  XOR2_X1 U935 ( .A(G1991), .B(G1996), .Z(n838) );
  XNOR2_X1 U936 ( .A(G1981), .B(G1966), .ZN(n837) );
  XNOR2_X1 U937 ( .A(n838), .B(n837), .ZN(n848) );
  XOR2_X1 U938 ( .A(KEYINPUT107), .B(KEYINPUT41), .Z(n840) );
  XNOR2_X1 U939 ( .A(G1956), .B(KEYINPUT108), .ZN(n839) );
  XNOR2_X1 U940 ( .A(n840), .B(n839), .ZN(n844) );
  XOR2_X1 U941 ( .A(G1986), .B(G1961), .Z(n842) );
  XNOR2_X1 U942 ( .A(G1976), .B(G1971), .ZN(n841) );
  XNOR2_X1 U943 ( .A(n842), .B(n841), .ZN(n843) );
  XOR2_X1 U944 ( .A(n844), .B(n843), .Z(n846) );
  XNOR2_X1 U945 ( .A(KEYINPUT109), .B(G2474), .ZN(n845) );
  XNOR2_X1 U946 ( .A(n846), .B(n845), .ZN(n847) );
  XOR2_X1 U947 ( .A(n848), .B(n847), .Z(G229) );
  XOR2_X1 U948 ( .A(G2096), .B(KEYINPUT43), .Z(n850) );
  XNOR2_X1 U949 ( .A(G2090), .B(KEYINPUT106), .ZN(n849) );
  XNOR2_X1 U950 ( .A(n850), .B(n849), .ZN(n851) );
  XOR2_X1 U951 ( .A(n851), .B(G2678), .Z(n853) );
  XNOR2_X1 U952 ( .A(G2067), .B(G2072), .ZN(n852) );
  XNOR2_X1 U953 ( .A(n853), .B(n852), .ZN(n857) );
  XOR2_X1 U954 ( .A(KEYINPUT42), .B(G2100), .Z(n855) );
  XNOR2_X1 U955 ( .A(G2084), .B(G2078), .ZN(n854) );
  XNOR2_X1 U956 ( .A(n855), .B(n854), .ZN(n856) );
  XNOR2_X1 U957 ( .A(n857), .B(n856), .ZN(G227) );
  NAND2_X1 U958 ( .A1(n877), .A2(G124), .ZN(n858) );
  XNOR2_X1 U959 ( .A(n858), .B(KEYINPUT44), .ZN(n860) );
  NAND2_X1 U960 ( .A1(G112), .A2(n878), .ZN(n859) );
  NAND2_X1 U961 ( .A1(n860), .A2(n859), .ZN(n864) );
  NAND2_X1 U962 ( .A1(G136), .A2(n882), .ZN(n862) );
  NAND2_X1 U963 ( .A1(G100), .A2(n885), .ZN(n861) );
  NAND2_X1 U964 ( .A1(n862), .A2(n861), .ZN(n863) );
  NOR2_X1 U965 ( .A1(n864), .A2(n863), .ZN(G162) );
  XOR2_X1 U966 ( .A(G160), .B(G162), .Z(n865) );
  XNOR2_X1 U967 ( .A(n866), .B(n865), .ZN(n893) );
  NAND2_X1 U968 ( .A1(G130), .A2(n877), .ZN(n868) );
  NAND2_X1 U969 ( .A1(G118), .A2(n878), .ZN(n867) );
  NAND2_X1 U970 ( .A1(n868), .A2(n867), .ZN(n873) );
  NAND2_X1 U971 ( .A1(G142), .A2(n882), .ZN(n870) );
  NAND2_X1 U972 ( .A1(G106), .A2(n885), .ZN(n869) );
  NAND2_X1 U973 ( .A1(n870), .A2(n869), .ZN(n871) );
  XOR2_X1 U974 ( .A(n871), .B(KEYINPUT45), .Z(n872) );
  NOR2_X1 U975 ( .A1(n873), .A2(n872), .ZN(n875) );
  XNOR2_X1 U976 ( .A(n875), .B(n874), .ZN(n876) );
  XOR2_X1 U977 ( .A(n876), .B(KEYINPUT48), .Z(n891) );
  NAND2_X1 U978 ( .A1(G127), .A2(n877), .ZN(n880) );
  NAND2_X1 U979 ( .A1(G115), .A2(n878), .ZN(n879) );
  NAND2_X1 U980 ( .A1(n880), .A2(n879), .ZN(n881) );
  XNOR2_X1 U981 ( .A(n881), .B(KEYINPUT47), .ZN(n884) );
  NAND2_X1 U982 ( .A1(G139), .A2(n882), .ZN(n883) );
  NAND2_X1 U983 ( .A1(n884), .A2(n883), .ZN(n888) );
  NAND2_X1 U984 ( .A1(n885), .A2(G103), .ZN(n886) );
  XOR2_X1 U985 ( .A(KEYINPUT110), .B(n886), .Z(n887) );
  NOR2_X1 U986 ( .A1(n888), .A2(n887), .ZN(n889) );
  XOR2_X1 U987 ( .A(KEYINPUT111), .B(n889), .Z(n937) );
  XNOR2_X1 U988 ( .A(n937), .B(KEYINPUT46), .ZN(n890) );
  XNOR2_X1 U989 ( .A(n891), .B(n890), .ZN(n892) );
  XNOR2_X1 U990 ( .A(n893), .B(n892), .ZN(n896) );
  XNOR2_X1 U991 ( .A(n894), .B(n930), .ZN(n895) );
  XNOR2_X1 U992 ( .A(n896), .B(n895), .ZN(n897) );
  XNOR2_X1 U993 ( .A(G164), .B(n897), .ZN(n898) );
  NOR2_X1 U994 ( .A1(G37), .A2(n898), .ZN(G395) );
  INV_X1 U995 ( .A(G301), .ZN(G171) );
  XOR2_X1 U996 ( .A(KEYINPUT112), .B(G286), .Z(n901) );
  XNOR2_X1 U997 ( .A(G171), .B(n899), .ZN(n900) );
  XNOR2_X1 U998 ( .A(n901), .B(n900), .ZN(n904) );
  XOR2_X1 U999 ( .A(n989), .B(n902), .Z(n903) );
  XNOR2_X1 U1000 ( .A(n904), .B(n903), .ZN(n905) );
  NOR2_X1 U1001 ( .A1(G37), .A2(n905), .ZN(n906) );
  XOR2_X1 U1002 ( .A(KEYINPUT113), .B(n906), .Z(G397) );
  XOR2_X1 U1003 ( .A(KEYINPUT103), .B(G2446), .Z(n908) );
  XNOR2_X1 U1004 ( .A(G2454), .B(G2451), .ZN(n907) );
  XNOR2_X1 U1005 ( .A(n908), .B(n907), .ZN(n909) );
  XOR2_X1 U1006 ( .A(n909), .B(G2430), .Z(n911) );
  XNOR2_X1 U1007 ( .A(G1341), .B(G1348), .ZN(n910) );
  XNOR2_X1 U1008 ( .A(n911), .B(n910), .ZN(n915) );
  XOR2_X1 U1009 ( .A(KEYINPUT101), .B(G2435), .Z(n913) );
  XNOR2_X1 U1010 ( .A(KEYINPUT102), .B(G2438), .ZN(n912) );
  XNOR2_X1 U1011 ( .A(n913), .B(n912), .ZN(n914) );
  XOR2_X1 U1012 ( .A(n915), .B(n914), .Z(n917) );
  XNOR2_X1 U1013 ( .A(G2443), .B(G2427), .ZN(n916) );
  XNOR2_X1 U1014 ( .A(n917), .B(n916), .ZN(n918) );
  NAND2_X1 U1015 ( .A1(n918), .A2(G14), .ZN(n924) );
  NAND2_X1 U1016 ( .A1(G319), .A2(n924), .ZN(n921) );
  NOR2_X1 U1017 ( .A1(G229), .A2(G227), .ZN(n919) );
  XNOR2_X1 U1018 ( .A(KEYINPUT49), .B(n919), .ZN(n920) );
  NOR2_X1 U1019 ( .A1(n921), .A2(n920), .ZN(n923) );
  NOR2_X1 U1020 ( .A1(G395), .A2(G397), .ZN(n922) );
  NAND2_X1 U1021 ( .A1(n923), .A2(n922), .ZN(G225) );
  INV_X1 U1022 ( .A(G225), .ZN(G308) );
  INV_X1 U1023 ( .A(G69), .ZN(G235) );
  INV_X1 U1024 ( .A(n924), .ZN(G401) );
  XOR2_X1 U1025 ( .A(G160), .B(G2084), .Z(n929) );
  XOR2_X1 U1026 ( .A(G2090), .B(G162), .Z(n925) );
  NOR2_X1 U1027 ( .A1(n926), .A2(n925), .ZN(n927) );
  XNOR2_X1 U1028 ( .A(KEYINPUT51), .B(n927), .ZN(n928) );
  NOR2_X1 U1029 ( .A1(n929), .A2(n928), .ZN(n936) );
  NOR2_X1 U1030 ( .A1(n931), .A2(n930), .ZN(n932) );
  XOR2_X1 U1031 ( .A(KEYINPUT114), .B(n932), .Z(n933) );
  NOR2_X1 U1032 ( .A1(n934), .A2(n933), .ZN(n935) );
  NAND2_X1 U1033 ( .A1(n936), .A2(n935), .ZN(n942) );
  XOR2_X1 U1034 ( .A(G2072), .B(n937), .Z(n939) );
  XOR2_X1 U1035 ( .A(G164), .B(G2078), .Z(n938) );
  NOR2_X1 U1036 ( .A1(n939), .A2(n938), .ZN(n940) );
  XOR2_X1 U1037 ( .A(KEYINPUT50), .B(n940), .Z(n941) );
  NOR2_X1 U1038 ( .A1(n942), .A2(n941), .ZN(n944) );
  NAND2_X1 U1039 ( .A1(n944), .A2(n943), .ZN(n945) );
  NOR2_X1 U1040 ( .A1(n946), .A2(n945), .ZN(n947) );
  XNOR2_X1 U1041 ( .A(KEYINPUT52), .B(n947), .ZN(n949) );
  INV_X1 U1042 ( .A(KEYINPUT55), .ZN(n948) );
  NAND2_X1 U1043 ( .A1(n949), .A2(n948), .ZN(n950) );
  NAND2_X1 U1044 ( .A1(n950), .A2(G29), .ZN(n1036) );
  XOR2_X1 U1045 ( .A(KEYINPUT116), .B(G34), .Z(n952) );
  XNOR2_X1 U1046 ( .A(G2084), .B(KEYINPUT54), .ZN(n951) );
  XNOR2_X1 U1047 ( .A(n952), .B(n951), .ZN(n969) );
  XNOR2_X1 U1048 ( .A(G2090), .B(G35), .ZN(n967) );
  XNOR2_X1 U1049 ( .A(G2067), .B(G26), .ZN(n954) );
  XNOR2_X1 U1050 ( .A(G2072), .B(G33), .ZN(n953) );
  NOR2_X1 U1051 ( .A1(n954), .A2(n953), .ZN(n960) );
  XNOR2_X1 U1052 ( .A(n955), .B(G32), .ZN(n958) );
  XNOR2_X1 U1053 ( .A(G27), .B(n956), .ZN(n957) );
  NOR2_X1 U1054 ( .A1(n958), .A2(n957), .ZN(n959) );
  NAND2_X1 U1055 ( .A1(n960), .A2(n959), .ZN(n964) );
  XOR2_X1 U1056 ( .A(G1991), .B(G25), .Z(n961) );
  NAND2_X1 U1057 ( .A1(n961), .A2(G28), .ZN(n962) );
  XOR2_X1 U1058 ( .A(KEYINPUT115), .B(n962), .Z(n963) );
  NOR2_X1 U1059 ( .A1(n964), .A2(n963), .ZN(n965) );
  XNOR2_X1 U1060 ( .A(KEYINPUT53), .B(n965), .ZN(n966) );
  NOR2_X1 U1061 ( .A1(n967), .A2(n966), .ZN(n968) );
  NAND2_X1 U1062 ( .A1(n969), .A2(n968), .ZN(n970) );
  XNOR2_X1 U1063 ( .A(KEYINPUT55), .B(n970), .ZN(n971) );
  NOR2_X1 U1064 ( .A1(G29), .A2(n971), .ZN(n972) );
  XNOR2_X1 U1065 ( .A(n972), .B(KEYINPUT117), .ZN(n973) );
  NAND2_X1 U1066 ( .A1(G11), .A2(n973), .ZN(n1034) );
  INV_X1 U1067 ( .A(G16), .ZN(n1030) );
  XOR2_X1 U1068 ( .A(KEYINPUT56), .B(KEYINPUT118), .Z(n974) );
  XNOR2_X1 U1069 ( .A(n1030), .B(n974), .ZN(n1003) );
  XNOR2_X1 U1070 ( .A(G301), .B(G1961), .ZN(n977) );
  XNOR2_X1 U1071 ( .A(n975), .B(G1348), .ZN(n976) );
  NOR2_X1 U1072 ( .A1(n977), .A2(n976), .ZN(n978) );
  XOR2_X1 U1073 ( .A(KEYINPUT120), .B(n978), .Z(n987) );
  XNOR2_X1 U1074 ( .A(KEYINPUT121), .B(n979), .ZN(n981) );
  NAND2_X1 U1075 ( .A1(n981), .A2(n980), .ZN(n982) );
  XNOR2_X1 U1076 ( .A(KEYINPUT122), .B(n982), .ZN(n984) );
  XNOR2_X1 U1077 ( .A(G166), .B(n1004), .ZN(n983) );
  NOR2_X1 U1078 ( .A1(n984), .A2(n983), .ZN(n985) );
  XNOR2_X1 U1079 ( .A(KEYINPUT123), .B(n985), .ZN(n986) );
  NOR2_X1 U1080 ( .A1(n987), .A2(n986), .ZN(n1001) );
  XOR2_X1 U1081 ( .A(G1341), .B(KEYINPUT124), .Z(n988) );
  XNOR2_X1 U1082 ( .A(n989), .B(n988), .ZN(n993) );
  XNOR2_X1 U1083 ( .A(G1956), .B(G299), .ZN(n990) );
  NOR2_X1 U1084 ( .A1(n991), .A2(n990), .ZN(n992) );
  NAND2_X1 U1085 ( .A1(n993), .A2(n992), .ZN(n999) );
  XOR2_X1 U1086 ( .A(G1966), .B(G168), .Z(n994) );
  XNOR2_X1 U1087 ( .A(KEYINPUT119), .B(n994), .ZN(n996) );
  NAND2_X1 U1088 ( .A1(n996), .A2(n995), .ZN(n997) );
  XOR2_X1 U1089 ( .A(KEYINPUT57), .B(n997), .Z(n998) );
  NOR2_X1 U1090 ( .A1(n999), .A2(n998), .ZN(n1000) );
  NAND2_X1 U1091 ( .A1(n1001), .A2(n1000), .ZN(n1002) );
  NAND2_X1 U1092 ( .A1(n1003), .A2(n1002), .ZN(n1032) );
  XOR2_X1 U1093 ( .A(G1961), .B(G5), .Z(n1011) );
  XOR2_X1 U1094 ( .A(G1976), .B(G23), .Z(n1006) );
  XNOR2_X1 U1095 ( .A(n1004), .B(G22), .ZN(n1005) );
  NAND2_X1 U1096 ( .A1(n1006), .A2(n1005), .ZN(n1008) );
  XNOR2_X1 U1097 ( .A(G24), .B(G1986), .ZN(n1007) );
  NOR2_X1 U1098 ( .A1(n1008), .A2(n1007), .ZN(n1009) );
  XNOR2_X1 U1099 ( .A(KEYINPUT58), .B(n1009), .ZN(n1010) );
  NAND2_X1 U1100 ( .A1(n1011), .A2(n1010), .ZN(n1027) );
  XOR2_X1 U1101 ( .A(G1966), .B(G21), .Z(n1024) );
  XOR2_X1 U1102 ( .A(G1341), .B(G19), .Z(n1014) );
  XNOR2_X1 U1103 ( .A(n1012), .B(G20), .ZN(n1013) );
  NAND2_X1 U1104 ( .A1(n1014), .A2(n1013), .ZN(n1016) );
  XNOR2_X1 U1105 ( .A(G6), .B(G1981), .ZN(n1015) );
  NOR2_X1 U1106 ( .A1(n1016), .A2(n1015), .ZN(n1020) );
  XOR2_X1 U1107 ( .A(G4), .B(KEYINPUT125), .Z(n1018) );
  XNOR2_X1 U1108 ( .A(G1348), .B(KEYINPUT59), .ZN(n1017) );
  XNOR2_X1 U1109 ( .A(n1018), .B(n1017), .ZN(n1019) );
  NAND2_X1 U1110 ( .A1(n1020), .A2(n1019), .ZN(n1021) );
  XOR2_X1 U1111 ( .A(KEYINPUT60), .B(n1021), .Z(n1022) );
  XNOR2_X1 U1112 ( .A(n1022), .B(KEYINPUT126), .ZN(n1023) );
  NAND2_X1 U1113 ( .A1(n1024), .A2(n1023), .ZN(n1025) );
  XOR2_X1 U1114 ( .A(KEYINPUT127), .B(n1025), .Z(n1026) );
  NOR2_X1 U1115 ( .A1(n1027), .A2(n1026), .ZN(n1028) );
  XNOR2_X1 U1116 ( .A(KEYINPUT61), .B(n1028), .ZN(n1029) );
  NAND2_X1 U1117 ( .A1(n1030), .A2(n1029), .ZN(n1031) );
  NAND2_X1 U1118 ( .A1(n1032), .A2(n1031), .ZN(n1033) );
  NOR2_X1 U1119 ( .A1(n1034), .A2(n1033), .ZN(n1035) );
  NAND2_X1 U1120 ( .A1(n1036), .A2(n1035), .ZN(n1037) );
  XOR2_X1 U1121 ( .A(KEYINPUT62), .B(n1037), .Z(G311) );
  INV_X1 U1122 ( .A(G311), .ZN(G150) );
endmodule

