

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n513, n514, n515, n516,
         n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527,
         n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538,
         n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549,
         n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560,
         n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571,
         n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582,
         n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593,
         n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604,
         n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615,
         n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626,
         n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637,
         n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648,
         n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659,
         n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670,
         n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681,
         n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692,
         n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703,
         n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714,
         n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725,
         n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736,
         n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747,
         n748, n749, n750, n751, n752, n753, n754, n755, n756, n757, n758,
         n759, n760, n761, n762, n763, n764, n765, n766, n767, n768, n769,
         n770, n771, n772, n773, n774, n775, n776, n777, n778, n779, n780,
         n781, n782, n783, n784, n785, n786, n787, n788, n789, n790, n791,
         n792, n793, n794, n795, n796, n797, n798, n799, n800, n801, n802,
         n803, n804, n805, n806, n807, n808, n809, n810, n811, n812, n813,
         n814, n815, n816, n817, n818, n819, n820, n821, n822, n823, n824,
         n825, n826, n827, n828, n829, n830, n831, n832, n833, n834, n835,
         n836, n837, n838, n839, n840, n841, n842, n843, n844, n845, n846,
         n847, n848, n849, n850, n851, n852, n853, n854, n855, n856, n857,
         n858, n859, n860, n861, n862, n863, n864, n865, n866, n867, n868,
         n869, n870, n871, n872, n873, n874, n875, n876, n877, n878, n879,
         n880, n881, n882, n883, n884, n885, n886, n887, n888, n889, n890,
         n891, n892, n893, n894, n895, n896, n897, n898, n899, n900, n901,
         n902, n903, n904, n905, n906, n907, n908, n909, n910, n911, n912,
         n913, n914, n915, n916, n917, n918, n919, n920, n921, n922, n923,
         n924, n925, n926, n927, n928, n929, n930, n931, n932, n933, n934,
         n935, n936, n937, n938, n939, n940, n941, n942, n943, n944, n945,
         n946, n947, n948, n949, n950, n951, n952, n953, n954, n955, n956,
         n957, n958, n959, n960, n961, n962, n963, n964, n965, n966, n967,
         n968, n969, n970, n971, n972, n973, n974, n975, n976, n977, n978,
         n979, n980, n981, n982, n983, n984, n985, n986, n987, n988, n989,
         n990, n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000,
         n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010,
         n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020,
         n1021, n1022, n1023, n1024;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  AND2_X1 U548 ( .A1(G2105), .A2(G2104), .ZN(n892) );
  AND2_X1 U549 ( .A1(n740), .A2(n739), .ZN(n741) );
  AND2_X1 U550 ( .A1(n605), .A2(n604), .ZN(n621) );
  NOR2_X2 U551 ( .A1(n563), .A2(n526), .ZN(n797) );
  OR2_X2 U552 ( .A1(n590), .A2(n769), .ZN(n686) );
  NAND2_X2 U553 ( .A1(n615), .A2(n614), .ZN(n970) );
  NOR2_X4 U554 ( .A1(G651), .A2(n563), .ZN(n592) );
  XOR2_X2 U555 ( .A(KEYINPUT0), .B(G543), .Z(n563) );
  INV_X1 U556 ( .A(KEYINPUT99), .ZN(n665) );
  OR2_X1 U557 ( .A1(n524), .A2(n523), .ZN(n582) );
  INV_X1 U558 ( .A(KEYINPUT95), .ZN(n627) );
  XNOR2_X1 U559 ( .A(n628), .B(n627), .ZN(n629) );
  XNOR2_X1 U560 ( .A(n668), .B(KEYINPUT32), .ZN(n676) );
  BUF_X2 U561 ( .A(n632), .Z(n622) );
  INV_X1 U562 ( .A(G1384), .ZN(n581) );
  INV_X1 U563 ( .A(KEYINPUT64), .ZN(n520) );
  AND2_X1 U564 ( .A1(n582), .A2(n581), .ZN(n687) );
  NAND2_X1 U565 ( .A1(G114), .A2(n892), .ZN(n513) );
  XNOR2_X1 U566 ( .A(n520), .B(KEYINPUT17), .ZN(n521) );
  AND2_X1 U567 ( .A1(n517), .A2(n516), .ZN(n518) );
  AND2_X2 U568 ( .A1(n515), .A2(G2104), .ZN(n895) );
  INV_X1 U569 ( .A(n582), .ZN(G164) );
  XOR2_X1 U570 ( .A(KEYINPUT87), .B(n513), .Z(n519) );
  INV_X1 U571 ( .A(G2105), .ZN(n515) );
  NOR2_X1 U572 ( .A1(G2104), .A2(n515), .ZN(n587) );
  NAND2_X1 U573 ( .A1(G126), .A2(n587), .ZN(n514) );
  XNOR2_X1 U574 ( .A(n514), .B(KEYINPUT86), .ZN(n517) );
  NAND2_X1 U575 ( .A1(n895), .A2(G102), .ZN(n516) );
  NAND2_X1 U576 ( .A1(n519), .A2(n518), .ZN(n524) );
  NOR2_X1 U577 ( .A1(G2105), .A2(G2104), .ZN(n522) );
  XNOR2_X2 U578 ( .A(n522), .B(n521), .ZN(n688) );
  AND2_X1 U579 ( .A1(G138), .A2(n688), .ZN(n523) );
  INV_X1 U580 ( .A(G651), .ZN(n526) );
  NOR2_X1 U581 ( .A1(G543), .A2(n526), .ZN(n525) );
  XOR2_X2 U582 ( .A(KEYINPUT1), .B(n525), .Z(n793) );
  NAND2_X1 U583 ( .A1(G65), .A2(n793), .ZN(n528) );
  NAND2_X1 U584 ( .A1(G78), .A2(n797), .ZN(n527) );
  NAND2_X1 U585 ( .A1(n528), .A2(n527), .ZN(n531) );
  NOR2_X2 U586 ( .A1(G651), .A2(G543), .ZN(n794) );
  NAND2_X1 U587 ( .A1(G91), .A2(n794), .ZN(n529) );
  XNOR2_X1 U588 ( .A(KEYINPUT65), .B(n529), .ZN(n530) );
  NOR2_X1 U589 ( .A1(n531), .A2(n530), .ZN(n533) );
  NAND2_X1 U590 ( .A1(n592), .A2(G53), .ZN(n532) );
  NAND2_X1 U591 ( .A1(n533), .A2(n532), .ZN(G299) );
  NAND2_X1 U592 ( .A1(G64), .A2(n793), .ZN(n535) );
  NAND2_X1 U593 ( .A1(G52), .A2(n592), .ZN(n534) );
  NAND2_X1 U594 ( .A1(n535), .A2(n534), .ZN(n540) );
  NAND2_X1 U595 ( .A1(G90), .A2(n794), .ZN(n537) );
  NAND2_X1 U596 ( .A1(G77), .A2(n797), .ZN(n536) );
  NAND2_X1 U597 ( .A1(n537), .A2(n536), .ZN(n538) );
  XOR2_X1 U598 ( .A(KEYINPUT9), .B(n538), .Z(n539) );
  NOR2_X1 U599 ( .A1(n540), .A2(n539), .ZN(G171) );
  INV_X1 U600 ( .A(G171), .ZN(G301) );
  NAND2_X1 U601 ( .A1(n794), .A2(G89), .ZN(n541) );
  XNOR2_X1 U602 ( .A(n541), .B(KEYINPUT4), .ZN(n543) );
  NAND2_X1 U603 ( .A1(G76), .A2(n797), .ZN(n542) );
  NAND2_X1 U604 ( .A1(n543), .A2(n542), .ZN(n544) );
  XNOR2_X1 U605 ( .A(n544), .B(KEYINPUT5), .ZN(n549) );
  NAND2_X1 U606 ( .A1(G63), .A2(n793), .ZN(n546) );
  NAND2_X1 U607 ( .A1(G51), .A2(n592), .ZN(n545) );
  NAND2_X1 U608 ( .A1(n546), .A2(n545), .ZN(n547) );
  XOR2_X1 U609 ( .A(KEYINPUT6), .B(n547), .Z(n548) );
  NAND2_X1 U610 ( .A1(n549), .A2(n548), .ZN(n550) );
  XNOR2_X1 U611 ( .A(n550), .B(KEYINPUT7), .ZN(G168) );
  XOR2_X1 U612 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U613 ( .A1(G62), .A2(n793), .ZN(n552) );
  NAND2_X1 U614 ( .A1(G50), .A2(n592), .ZN(n551) );
  NAND2_X1 U615 ( .A1(n552), .A2(n551), .ZN(n558) );
  NAND2_X1 U616 ( .A1(n794), .A2(G88), .ZN(n553) );
  XNOR2_X1 U617 ( .A(n553), .B(KEYINPUT78), .ZN(n555) );
  NAND2_X1 U618 ( .A1(G75), .A2(n797), .ZN(n554) );
  NAND2_X1 U619 ( .A1(n555), .A2(n554), .ZN(n556) );
  XOR2_X1 U620 ( .A(KEYINPUT79), .B(n556), .Z(n557) );
  NOR2_X1 U621 ( .A1(n558), .A2(n557), .ZN(G166) );
  INV_X1 U622 ( .A(G166), .ZN(G303) );
  NAND2_X1 U623 ( .A1(G49), .A2(n592), .ZN(n560) );
  NAND2_X1 U624 ( .A1(G74), .A2(G651), .ZN(n559) );
  NAND2_X1 U625 ( .A1(n560), .A2(n559), .ZN(n561) );
  XOR2_X1 U626 ( .A(KEYINPUT75), .B(n561), .Z(n562) );
  NOR2_X1 U627 ( .A1(n793), .A2(n562), .ZN(n565) );
  NAND2_X1 U628 ( .A1(n563), .A2(G87), .ZN(n564) );
  NAND2_X1 U629 ( .A1(n565), .A2(n564), .ZN(G288) );
  NAND2_X1 U630 ( .A1(G73), .A2(n797), .ZN(n566) );
  XNOR2_X1 U631 ( .A(n566), .B(KEYINPUT2), .ZN(n574) );
  NAND2_X1 U632 ( .A1(G61), .A2(n793), .ZN(n568) );
  NAND2_X1 U633 ( .A1(G86), .A2(n794), .ZN(n567) );
  NAND2_X1 U634 ( .A1(n568), .A2(n567), .ZN(n569) );
  XNOR2_X1 U635 ( .A(KEYINPUT76), .B(n569), .ZN(n572) );
  NAND2_X1 U636 ( .A1(G48), .A2(n592), .ZN(n570) );
  XNOR2_X1 U637 ( .A(KEYINPUT77), .B(n570), .ZN(n571) );
  NOR2_X1 U638 ( .A1(n572), .A2(n571), .ZN(n573) );
  NAND2_X1 U639 ( .A1(n574), .A2(n573), .ZN(G305) );
  NAND2_X1 U640 ( .A1(G85), .A2(n794), .ZN(n576) );
  NAND2_X1 U641 ( .A1(G72), .A2(n797), .ZN(n575) );
  NAND2_X1 U642 ( .A1(n576), .A2(n575), .ZN(n580) );
  NAND2_X1 U643 ( .A1(G60), .A2(n793), .ZN(n578) );
  NAND2_X1 U644 ( .A1(G47), .A2(n592), .ZN(n577) );
  NAND2_X1 U645 ( .A1(n578), .A2(n577), .ZN(n579) );
  OR2_X1 U646 ( .A1(n580), .A2(n579), .ZN(G290) );
  NAND2_X1 U647 ( .A1(n892), .A2(G113), .ZN(n585) );
  NAND2_X1 U648 ( .A1(G101), .A2(n895), .ZN(n583) );
  XOR2_X1 U649 ( .A(KEYINPUT23), .B(n583), .Z(n584) );
  NAND2_X1 U650 ( .A1(n585), .A2(n584), .ZN(n768) );
  INV_X1 U651 ( .A(n768), .ZN(n586) );
  NAND2_X1 U652 ( .A1(G40), .A2(n586), .ZN(n590) );
  BUF_X1 U653 ( .A(n587), .Z(n891) );
  NAND2_X1 U654 ( .A1(G125), .A2(n891), .ZN(n589) );
  NAND2_X1 U655 ( .A1(G137), .A2(n688), .ZN(n588) );
  NAND2_X1 U656 ( .A1(n589), .A2(n588), .ZN(n769) );
  INV_X1 U657 ( .A(n686), .ZN(n591) );
  NAND2_X2 U658 ( .A1(n687), .A2(n591), .ZN(n632) );
  NAND2_X2 U659 ( .A1(G8), .A2(n622), .ZN(n731) );
  NAND2_X1 U660 ( .A1(G79), .A2(n797), .ZN(n594) );
  NAND2_X1 U661 ( .A1(G54), .A2(n592), .ZN(n593) );
  NAND2_X1 U662 ( .A1(n594), .A2(n593), .ZN(n595) );
  XNOR2_X1 U663 ( .A(n595), .B(KEYINPUT69), .ZN(n600) );
  AND2_X1 U664 ( .A1(G66), .A2(n793), .ZN(n598) );
  NAND2_X1 U665 ( .A1(n794), .A2(G92), .ZN(n596) );
  XOR2_X1 U666 ( .A(KEYINPUT68), .B(n596), .Z(n597) );
  NOR2_X1 U667 ( .A1(n598), .A2(n597), .ZN(n599) );
  AND2_X1 U668 ( .A1(n600), .A2(n599), .ZN(n601) );
  XOR2_X1 U669 ( .A(KEYINPUT15), .B(n601), .Z(n618) );
  BUF_X1 U670 ( .A(n618), .Z(n965) );
  INV_X1 U671 ( .A(n632), .ZN(n602) );
  NAND2_X1 U672 ( .A1(n602), .A2(G1996), .ZN(n603) );
  XNOR2_X1 U673 ( .A(n603), .B(KEYINPUT26), .ZN(n605) );
  NAND2_X1 U674 ( .A1(n622), .A2(G1341), .ZN(n604) );
  NAND2_X1 U675 ( .A1(n793), .A2(G56), .ZN(n606) );
  XNOR2_X1 U676 ( .A(KEYINPUT14), .B(n606), .ZN(n612) );
  NAND2_X1 U677 ( .A1(n794), .A2(G81), .ZN(n607) );
  XNOR2_X1 U678 ( .A(n607), .B(KEYINPUT12), .ZN(n609) );
  NAND2_X1 U679 ( .A1(G68), .A2(n797), .ZN(n608) );
  NAND2_X1 U680 ( .A1(n609), .A2(n608), .ZN(n610) );
  XNOR2_X1 U681 ( .A(n610), .B(KEYINPUT13), .ZN(n611) );
  NAND2_X1 U682 ( .A1(n612), .A2(n611), .ZN(n613) );
  XNOR2_X1 U683 ( .A(n613), .B(KEYINPUT67), .ZN(n615) );
  NAND2_X1 U684 ( .A1(n592), .A2(G43), .ZN(n614) );
  INV_X1 U685 ( .A(n970), .ZN(n616) );
  AND2_X1 U686 ( .A1(n621), .A2(n616), .ZN(n617) );
  OR2_X1 U687 ( .A1(n965), .A2(n617), .ZN(n630) );
  INV_X1 U688 ( .A(n618), .ZN(n619) );
  NOR2_X1 U689 ( .A1(n970), .A2(n619), .ZN(n620) );
  NAND2_X1 U690 ( .A1(n621), .A2(n620), .ZN(n626) );
  NOR2_X1 U691 ( .A1(n643), .A2(G1348), .ZN(n624) );
  NOR2_X1 U692 ( .A1(G2067), .A2(n622), .ZN(n623) );
  NOR2_X1 U693 ( .A1(n624), .A2(n623), .ZN(n625) );
  NAND2_X1 U694 ( .A1(n626), .A2(n625), .ZN(n628) );
  NAND2_X1 U695 ( .A1(n630), .A2(n629), .ZN(n637) );
  INV_X1 U696 ( .A(G299), .ZN(n806) );
  INV_X1 U697 ( .A(n632), .ZN(n643) );
  NAND2_X1 U698 ( .A1(n643), .A2(G2072), .ZN(n631) );
  XNOR2_X1 U699 ( .A(KEYINPUT27), .B(n631), .ZN(n635) );
  NAND2_X1 U700 ( .A1(G1956), .A2(n632), .ZN(n633) );
  XOR2_X1 U701 ( .A(KEYINPUT94), .B(n633), .Z(n634) );
  NOR2_X1 U702 ( .A1(n635), .A2(n634), .ZN(n638) );
  NAND2_X1 U703 ( .A1(n806), .A2(n638), .ZN(n636) );
  NAND2_X1 U704 ( .A1(n637), .A2(n636), .ZN(n641) );
  NOR2_X1 U705 ( .A1(n806), .A2(n638), .ZN(n639) );
  XOR2_X1 U706 ( .A(n639), .B(KEYINPUT28), .Z(n640) );
  NAND2_X1 U707 ( .A1(n641), .A2(n640), .ZN(n642) );
  XNOR2_X1 U708 ( .A(n642), .B(KEYINPUT29), .ZN(n647) );
  NAND2_X1 U709 ( .A1(G1961), .A2(n622), .ZN(n645) );
  XOR2_X1 U710 ( .A(G2078), .B(KEYINPUT25), .Z(n945) );
  NAND2_X1 U711 ( .A1(n643), .A2(n945), .ZN(n644) );
  NAND2_X1 U712 ( .A1(n645), .A2(n644), .ZN(n648) );
  NOR2_X1 U713 ( .A1(G301), .A2(n648), .ZN(n646) );
  NOR2_X1 U714 ( .A1(n647), .A2(n646), .ZN(n657) );
  NAND2_X1 U715 ( .A1(G301), .A2(n648), .ZN(n649) );
  XOR2_X1 U716 ( .A(KEYINPUT96), .B(n649), .Z(n654) );
  NOR2_X1 U717 ( .A1(G1966), .A2(n731), .ZN(n672) );
  NOR2_X1 U718 ( .A1(G2084), .A2(n622), .ZN(n669) );
  NOR2_X1 U719 ( .A1(n672), .A2(n669), .ZN(n650) );
  NAND2_X1 U720 ( .A1(G8), .A2(n650), .ZN(n651) );
  XNOR2_X1 U721 ( .A(KEYINPUT30), .B(n651), .ZN(n652) );
  NOR2_X1 U722 ( .A1(G168), .A2(n652), .ZN(n653) );
  NOR2_X1 U723 ( .A1(n654), .A2(n653), .ZN(n655) );
  XNOR2_X1 U724 ( .A(n655), .B(KEYINPUT31), .ZN(n656) );
  NOR2_X1 U725 ( .A1(n657), .A2(n656), .ZN(n658) );
  XNOR2_X1 U726 ( .A(n658), .B(KEYINPUT97), .ZN(n670) );
  NAND2_X1 U727 ( .A1(n670), .A2(G286), .ZN(n664) );
  NOR2_X1 U728 ( .A1(G1971), .A2(n731), .ZN(n659) );
  XNOR2_X1 U729 ( .A(n659), .B(KEYINPUT98), .ZN(n661) );
  NOR2_X1 U730 ( .A1(n622), .A2(G2090), .ZN(n660) );
  NOR2_X1 U731 ( .A1(n661), .A2(n660), .ZN(n662) );
  NAND2_X1 U732 ( .A1(n662), .A2(G303), .ZN(n663) );
  NAND2_X1 U733 ( .A1(n664), .A2(n663), .ZN(n666) );
  XNOR2_X1 U734 ( .A(n666), .B(n665), .ZN(n667) );
  NAND2_X1 U735 ( .A1(n667), .A2(G8), .ZN(n668) );
  NAND2_X1 U736 ( .A1(G8), .A2(n669), .ZN(n674) );
  INV_X1 U737 ( .A(n670), .ZN(n671) );
  NOR2_X1 U738 ( .A1(n672), .A2(n671), .ZN(n673) );
  NAND2_X1 U739 ( .A1(n674), .A2(n673), .ZN(n675) );
  NAND2_X1 U740 ( .A1(n676), .A2(n675), .ZN(n724) );
  NOR2_X1 U741 ( .A1(G1971), .A2(G303), .ZN(n677) );
  NOR2_X1 U742 ( .A1(G1976), .A2(G288), .ZN(n973) );
  NOR2_X1 U743 ( .A1(n677), .A2(n973), .ZN(n678) );
  NAND2_X1 U744 ( .A1(n724), .A2(n678), .ZN(n679) );
  NAND2_X1 U745 ( .A1(G1976), .A2(G288), .ZN(n974) );
  NAND2_X1 U746 ( .A1(n679), .A2(n974), .ZN(n680) );
  XNOR2_X1 U747 ( .A(KEYINPUT100), .B(n680), .ZN(n681) );
  NOR2_X1 U748 ( .A1(n731), .A2(n681), .ZN(n682) );
  NOR2_X1 U749 ( .A1(KEYINPUT33), .A2(n682), .ZN(n685) );
  NAND2_X1 U750 ( .A1(n973), .A2(KEYINPUT33), .ZN(n683) );
  NOR2_X1 U751 ( .A1(n683), .A2(n731), .ZN(n684) );
  NOR2_X1 U752 ( .A1(n685), .A2(n684), .ZN(n723) );
  XOR2_X1 U753 ( .A(G1981), .B(G305), .Z(n987) );
  NOR2_X1 U754 ( .A1(n687), .A2(n686), .ZN(n753) );
  XNOR2_X1 U755 ( .A(G1986), .B(G290), .ZN(n967) );
  NAND2_X1 U756 ( .A1(n753), .A2(n967), .ZN(n734) );
  AND2_X1 U757 ( .A1(n987), .A2(n734), .ZN(n721) );
  NAND2_X1 U758 ( .A1(n895), .A2(G104), .ZN(n690) );
  NAND2_X1 U759 ( .A1(G140), .A2(n688), .ZN(n689) );
  NAND2_X1 U760 ( .A1(n690), .A2(n689), .ZN(n691) );
  XNOR2_X1 U761 ( .A(KEYINPUT34), .B(n691), .ZN(n696) );
  NAND2_X1 U762 ( .A1(G128), .A2(n891), .ZN(n693) );
  NAND2_X1 U763 ( .A1(G116), .A2(n892), .ZN(n692) );
  NAND2_X1 U764 ( .A1(n693), .A2(n692), .ZN(n694) );
  XOR2_X1 U765 ( .A(n694), .B(KEYINPUT35), .Z(n695) );
  NOR2_X1 U766 ( .A1(n696), .A2(n695), .ZN(n697) );
  XOR2_X1 U767 ( .A(KEYINPUT36), .B(n697), .Z(n698) );
  XOR2_X1 U768 ( .A(KEYINPUT88), .B(n698), .Z(n906) );
  XNOR2_X1 U769 ( .A(G2067), .B(KEYINPUT37), .ZN(n750) );
  NOR2_X1 U770 ( .A1(n906), .A2(n750), .ZN(n922) );
  NAND2_X1 U771 ( .A1(n753), .A2(n922), .ZN(n747) );
  INV_X1 U772 ( .A(n747), .ZN(n719) );
  NAND2_X1 U773 ( .A1(G105), .A2(n895), .ZN(n699) );
  XOR2_X1 U774 ( .A(KEYINPUT38), .B(n699), .Z(n704) );
  NAND2_X1 U775 ( .A1(G129), .A2(n891), .ZN(n701) );
  NAND2_X1 U776 ( .A1(G117), .A2(n892), .ZN(n700) );
  NAND2_X1 U777 ( .A1(n701), .A2(n700), .ZN(n702) );
  XOR2_X1 U778 ( .A(KEYINPUT91), .B(n702), .Z(n703) );
  NOR2_X1 U779 ( .A1(n704), .A2(n703), .ZN(n706) );
  NAND2_X1 U780 ( .A1(G141), .A2(n688), .ZN(n705) );
  NAND2_X1 U781 ( .A1(n706), .A2(n705), .ZN(n901) );
  NAND2_X1 U782 ( .A1(G1996), .A2(n901), .ZN(n707) );
  XNOR2_X1 U783 ( .A(n707), .B(KEYINPUT92), .ZN(n717) );
  NAND2_X1 U784 ( .A1(G95), .A2(n895), .ZN(n714) );
  NAND2_X1 U785 ( .A1(G119), .A2(n891), .ZN(n709) );
  NAND2_X1 U786 ( .A1(G107), .A2(n892), .ZN(n708) );
  NAND2_X1 U787 ( .A1(n709), .A2(n708), .ZN(n712) );
  NAND2_X1 U788 ( .A1(G131), .A2(n688), .ZN(n710) );
  XNOR2_X1 U789 ( .A(KEYINPUT89), .B(n710), .ZN(n711) );
  NOR2_X1 U790 ( .A1(n712), .A2(n711), .ZN(n713) );
  NAND2_X1 U791 ( .A1(n714), .A2(n713), .ZN(n715) );
  XNOR2_X1 U792 ( .A(n715), .B(KEYINPUT90), .ZN(n876) );
  NAND2_X1 U793 ( .A1(n876), .A2(G1991), .ZN(n716) );
  NAND2_X1 U794 ( .A1(n717), .A2(n716), .ZN(n928) );
  NAND2_X1 U795 ( .A1(n928), .A2(n753), .ZN(n718) );
  XNOR2_X1 U796 ( .A(n718), .B(KEYINPUT93), .ZN(n744) );
  OR2_X1 U797 ( .A1(n719), .A2(n744), .ZN(n736) );
  INV_X1 U798 ( .A(n736), .ZN(n720) );
  AND2_X1 U799 ( .A1(n721), .A2(n720), .ZN(n722) );
  NAND2_X1 U800 ( .A1(n723), .A2(n722), .ZN(n740) );
  NOR2_X1 U801 ( .A1(G2090), .A2(G303), .ZN(n725) );
  NAND2_X1 U802 ( .A1(G8), .A2(n725), .ZN(n726) );
  NAND2_X1 U803 ( .A1(n724), .A2(n726), .ZN(n727) );
  NAND2_X1 U804 ( .A1(n727), .A2(n731), .ZN(n728) );
  XNOR2_X1 U805 ( .A(n728), .B(KEYINPUT101), .ZN(n733) );
  NOR2_X1 U806 ( .A1(G1981), .A2(G305), .ZN(n729) );
  XOR2_X1 U807 ( .A(n729), .B(KEYINPUT24), .Z(n730) );
  NOR2_X1 U808 ( .A1(n731), .A2(n730), .ZN(n732) );
  OR2_X1 U809 ( .A1(n733), .A2(n732), .ZN(n738) );
  INV_X1 U810 ( .A(n734), .ZN(n735) );
  NOR2_X1 U811 ( .A1(n736), .A2(n735), .ZN(n737) );
  NAND2_X1 U812 ( .A1(n738), .A2(n737), .ZN(n739) );
  XNOR2_X1 U813 ( .A(n741), .B(KEYINPUT102), .ZN(n756) );
  NOR2_X1 U814 ( .A1(G1996), .A2(n901), .ZN(n932) );
  NOR2_X1 U815 ( .A1(G1991), .A2(n876), .ZN(n924) );
  NOR2_X1 U816 ( .A1(G1986), .A2(G290), .ZN(n742) );
  NOR2_X1 U817 ( .A1(n924), .A2(n742), .ZN(n743) );
  NOR2_X1 U818 ( .A1(n744), .A2(n743), .ZN(n745) );
  NOR2_X1 U819 ( .A1(n932), .A2(n745), .ZN(n746) );
  XNOR2_X1 U820 ( .A(n746), .B(KEYINPUT39), .ZN(n748) );
  NAND2_X1 U821 ( .A1(n748), .A2(n747), .ZN(n749) );
  XOR2_X1 U822 ( .A(KEYINPUT103), .B(n749), .Z(n752) );
  NAND2_X1 U823 ( .A1(n906), .A2(n750), .ZN(n751) );
  XNOR2_X1 U824 ( .A(n751), .B(KEYINPUT104), .ZN(n934) );
  NAND2_X1 U825 ( .A1(n752), .A2(n934), .ZN(n754) );
  NAND2_X1 U826 ( .A1(n754), .A2(n753), .ZN(n755) );
  NAND2_X1 U827 ( .A1(n756), .A2(n755), .ZN(n758) );
  XOR2_X1 U828 ( .A(KEYINPUT105), .B(KEYINPUT40), .Z(n757) );
  XNOR2_X1 U829 ( .A(n758), .B(n757), .ZN(G329) );
  XNOR2_X1 U830 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  XOR2_X1 U831 ( .A(G2443), .B(G2446), .Z(n760) );
  XNOR2_X1 U832 ( .A(G2427), .B(G2451), .ZN(n759) );
  XNOR2_X1 U833 ( .A(n760), .B(n759), .ZN(n766) );
  XOR2_X1 U834 ( .A(G2430), .B(G2454), .Z(n762) );
  XNOR2_X1 U835 ( .A(G1341), .B(G1348), .ZN(n761) );
  XNOR2_X1 U836 ( .A(n762), .B(n761), .ZN(n764) );
  XOR2_X1 U837 ( .A(G2435), .B(G2438), .Z(n763) );
  XNOR2_X1 U838 ( .A(n764), .B(n763), .ZN(n765) );
  XOR2_X1 U839 ( .A(n766), .B(n765), .Z(n767) );
  AND2_X1 U840 ( .A1(G14), .A2(n767), .ZN(G401) );
  AND2_X1 U841 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U842 ( .A(G132), .ZN(G219) );
  INV_X1 U843 ( .A(G82), .ZN(G220) );
  INV_X1 U844 ( .A(G120), .ZN(G236) );
  INV_X1 U845 ( .A(G69), .ZN(G235) );
  NOR2_X1 U846 ( .A1(n769), .A2(n768), .ZN(G160) );
  NAND2_X1 U847 ( .A1(G7), .A2(G661), .ZN(n770) );
  XNOR2_X1 U848 ( .A(n770), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U849 ( .A(G223), .ZN(n836) );
  NAND2_X1 U850 ( .A1(n836), .A2(G567), .ZN(n771) );
  XOR2_X1 U851 ( .A(KEYINPUT11), .B(n771), .Z(G234) );
  INV_X1 U852 ( .A(G860), .ZN(n803) );
  OR2_X1 U853 ( .A1(n970), .A2(n803), .ZN(G153) );
  NAND2_X1 U854 ( .A1(G868), .A2(G301), .ZN(n773) );
  INV_X1 U855 ( .A(G868), .ZN(n816) );
  NAND2_X1 U856 ( .A1(n619), .A2(n816), .ZN(n772) );
  NAND2_X1 U857 ( .A1(n773), .A2(n772), .ZN(G284) );
  NOR2_X1 U858 ( .A1(G868), .A2(G299), .ZN(n774) );
  XNOR2_X1 U859 ( .A(n774), .B(KEYINPUT70), .ZN(n776) );
  NOR2_X1 U860 ( .A1(n816), .A2(G286), .ZN(n775) );
  NOR2_X1 U861 ( .A1(n776), .A2(n775), .ZN(G297) );
  NAND2_X1 U862 ( .A1(n803), .A2(G559), .ZN(n777) );
  NAND2_X1 U863 ( .A1(n777), .A2(n965), .ZN(n778) );
  XNOR2_X1 U864 ( .A(n778), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U865 ( .A1(n619), .A2(n816), .ZN(n779) );
  XNOR2_X1 U866 ( .A(n779), .B(KEYINPUT71), .ZN(n780) );
  NOR2_X1 U867 ( .A1(G559), .A2(n780), .ZN(n782) );
  NOR2_X1 U868 ( .A1(G868), .A2(n970), .ZN(n781) );
  NOR2_X1 U869 ( .A1(n782), .A2(n781), .ZN(G282) );
  NAND2_X1 U870 ( .A1(G111), .A2(n892), .ZN(n784) );
  NAND2_X1 U871 ( .A1(G135), .A2(n688), .ZN(n783) );
  NAND2_X1 U872 ( .A1(n784), .A2(n783), .ZN(n787) );
  NAND2_X1 U873 ( .A1(n891), .A2(G123), .ZN(n785) );
  XOR2_X1 U874 ( .A(KEYINPUT18), .B(n785), .Z(n786) );
  NOR2_X1 U875 ( .A1(n787), .A2(n786), .ZN(n789) );
  NAND2_X1 U876 ( .A1(n895), .A2(G99), .ZN(n788) );
  NAND2_X1 U877 ( .A1(n789), .A2(n788), .ZN(n925) );
  XNOR2_X1 U878 ( .A(n925), .B(G2096), .ZN(n791) );
  XNOR2_X1 U879 ( .A(G2100), .B(KEYINPUT72), .ZN(n790) );
  NOR2_X1 U880 ( .A1(n791), .A2(n790), .ZN(n792) );
  XNOR2_X1 U881 ( .A(KEYINPUT73), .B(n792), .ZN(G156) );
  NAND2_X1 U882 ( .A1(G67), .A2(n793), .ZN(n796) );
  NAND2_X1 U883 ( .A1(G93), .A2(n794), .ZN(n795) );
  NAND2_X1 U884 ( .A1(n796), .A2(n795), .ZN(n801) );
  NAND2_X1 U885 ( .A1(G80), .A2(n797), .ZN(n799) );
  NAND2_X1 U886 ( .A1(G55), .A2(n592), .ZN(n798) );
  NAND2_X1 U887 ( .A1(n799), .A2(n798), .ZN(n800) );
  OR2_X1 U888 ( .A1(n801), .A2(n800), .ZN(n817) );
  XNOR2_X1 U889 ( .A(n817), .B(KEYINPUT74), .ZN(n805) );
  NAND2_X1 U890 ( .A1(G559), .A2(n965), .ZN(n802) );
  XOR2_X1 U891 ( .A(n970), .B(n802), .Z(n813) );
  NAND2_X1 U892 ( .A1(n813), .A2(n803), .ZN(n804) );
  XNOR2_X1 U893 ( .A(n805), .B(n804), .ZN(G145) );
  XNOR2_X1 U894 ( .A(KEYINPUT80), .B(KEYINPUT19), .ZN(n808) );
  XNOR2_X1 U895 ( .A(G290), .B(n806), .ZN(n807) );
  XNOR2_X1 U896 ( .A(n808), .B(n807), .ZN(n809) );
  XOR2_X1 U897 ( .A(n817), .B(n809), .Z(n811) );
  XNOR2_X1 U898 ( .A(G288), .B(G166), .ZN(n810) );
  XNOR2_X1 U899 ( .A(n811), .B(n810), .ZN(n812) );
  XNOR2_X1 U900 ( .A(n812), .B(G305), .ZN(n862) );
  XNOR2_X1 U901 ( .A(n813), .B(n862), .ZN(n814) );
  XNOR2_X1 U902 ( .A(KEYINPUT81), .B(n814), .ZN(n815) );
  NOR2_X1 U903 ( .A1(n816), .A2(n815), .ZN(n819) );
  NOR2_X1 U904 ( .A1(G868), .A2(n817), .ZN(n818) );
  NOR2_X1 U905 ( .A1(n819), .A2(n818), .ZN(G295) );
  NAND2_X1 U906 ( .A1(G2078), .A2(G2084), .ZN(n821) );
  XOR2_X1 U907 ( .A(KEYINPUT82), .B(KEYINPUT20), .Z(n820) );
  XNOR2_X1 U908 ( .A(n821), .B(n820), .ZN(n822) );
  NAND2_X1 U909 ( .A1(G2090), .A2(n822), .ZN(n823) );
  XNOR2_X1 U910 ( .A(KEYINPUT21), .B(n823), .ZN(n824) );
  NAND2_X1 U911 ( .A1(n824), .A2(G2072), .ZN(G158) );
  XOR2_X1 U912 ( .A(KEYINPUT66), .B(G57), .Z(G237) );
  NOR2_X1 U913 ( .A1(G235), .A2(G236), .ZN(n825) );
  XNOR2_X1 U914 ( .A(n825), .B(KEYINPUT83), .ZN(n826) );
  NOR2_X1 U915 ( .A1(G237), .A2(n826), .ZN(n827) );
  XNOR2_X1 U916 ( .A(KEYINPUT84), .B(n827), .ZN(n828) );
  NAND2_X1 U917 ( .A1(n828), .A2(G108), .ZN(n840) );
  NAND2_X1 U918 ( .A1(G567), .A2(n840), .ZN(n829) );
  XNOR2_X1 U919 ( .A(n829), .B(KEYINPUT85), .ZN(n834) );
  NOR2_X1 U920 ( .A1(G220), .A2(G219), .ZN(n830) );
  XNOR2_X1 U921 ( .A(KEYINPUT22), .B(n830), .ZN(n831) );
  NAND2_X1 U922 ( .A1(n831), .A2(G96), .ZN(n832) );
  OR2_X1 U923 ( .A1(G218), .A2(n832), .ZN(n841) );
  AND2_X1 U924 ( .A1(G2106), .A2(n841), .ZN(n833) );
  NOR2_X1 U925 ( .A1(n834), .A2(n833), .ZN(G319) );
  INV_X1 U926 ( .A(G319), .ZN(n912) );
  NAND2_X1 U927 ( .A1(G483), .A2(G661), .ZN(n835) );
  NOR2_X1 U928 ( .A1(n912), .A2(n835), .ZN(n839) );
  NAND2_X1 U929 ( .A1(n839), .A2(G36), .ZN(G176) );
  NAND2_X1 U930 ( .A1(G2106), .A2(n836), .ZN(G217) );
  AND2_X1 U931 ( .A1(G15), .A2(G2), .ZN(n837) );
  NAND2_X1 U932 ( .A1(G661), .A2(n837), .ZN(G259) );
  NAND2_X1 U933 ( .A1(G3), .A2(G1), .ZN(n838) );
  NAND2_X1 U934 ( .A1(n839), .A2(n838), .ZN(G188) );
  NOR2_X1 U936 ( .A1(n841), .A2(n840), .ZN(n842) );
  XNOR2_X1 U937 ( .A(KEYINPUT106), .B(n842), .ZN(G325) );
  XNOR2_X1 U938 ( .A(KEYINPUT107), .B(G325), .ZN(G261) );
  INV_X1 U939 ( .A(G108), .ZN(G238) );
  INV_X1 U940 ( .A(G96), .ZN(G221) );
  XOR2_X1 U941 ( .A(G2096), .B(KEYINPUT43), .Z(n844) );
  XNOR2_X1 U942 ( .A(G2090), .B(G2678), .ZN(n843) );
  XNOR2_X1 U943 ( .A(n844), .B(n843), .ZN(n845) );
  XOR2_X1 U944 ( .A(n845), .B(KEYINPUT42), .Z(n847) );
  XNOR2_X1 U945 ( .A(G2067), .B(G2072), .ZN(n846) );
  XNOR2_X1 U946 ( .A(n847), .B(n846), .ZN(n851) );
  XOR2_X1 U947 ( .A(KEYINPUT108), .B(G2100), .Z(n849) );
  XNOR2_X1 U948 ( .A(G2078), .B(G2084), .ZN(n848) );
  XNOR2_X1 U949 ( .A(n849), .B(n848), .ZN(n850) );
  XNOR2_X1 U950 ( .A(n851), .B(n850), .ZN(G227) );
  XOR2_X1 U951 ( .A(G1956), .B(G1966), .Z(n853) );
  XNOR2_X1 U952 ( .A(G1981), .B(G1976), .ZN(n852) );
  XNOR2_X1 U953 ( .A(n853), .B(n852), .ZN(n857) );
  XOR2_X1 U954 ( .A(G1971), .B(G1986), .Z(n855) );
  XNOR2_X1 U955 ( .A(G1996), .B(G1991), .ZN(n854) );
  XNOR2_X1 U956 ( .A(n855), .B(n854), .ZN(n856) );
  XOR2_X1 U957 ( .A(n857), .B(n856), .Z(n859) );
  XNOR2_X1 U958 ( .A(KEYINPUT109), .B(G2474), .ZN(n858) );
  XNOR2_X1 U959 ( .A(n859), .B(n858), .ZN(n861) );
  XOR2_X1 U960 ( .A(G1961), .B(KEYINPUT41), .Z(n860) );
  XNOR2_X1 U961 ( .A(n861), .B(n860), .ZN(G229) );
  XOR2_X1 U962 ( .A(n862), .B(G286), .Z(n864) );
  XNOR2_X1 U963 ( .A(G171), .B(n965), .ZN(n863) );
  XNOR2_X1 U964 ( .A(n864), .B(n863), .ZN(n865) );
  XNOR2_X1 U965 ( .A(n865), .B(n970), .ZN(n866) );
  NOR2_X1 U966 ( .A1(G37), .A2(n866), .ZN(G397) );
  NAND2_X1 U967 ( .A1(G112), .A2(n892), .ZN(n868) );
  NAND2_X1 U968 ( .A1(G100), .A2(n895), .ZN(n867) );
  NAND2_X1 U969 ( .A1(n868), .A2(n867), .ZN(n875) );
  NAND2_X1 U970 ( .A1(n891), .A2(G124), .ZN(n869) );
  XOR2_X1 U971 ( .A(KEYINPUT44), .B(n869), .Z(n872) );
  NAND2_X1 U972 ( .A1(G136), .A2(n688), .ZN(n870) );
  XOR2_X1 U973 ( .A(KEYINPUT110), .B(n870), .Z(n871) );
  NOR2_X1 U974 ( .A1(n872), .A2(n871), .ZN(n873) );
  XNOR2_X1 U975 ( .A(n873), .B(KEYINPUT111), .ZN(n874) );
  NOR2_X1 U976 ( .A1(n875), .A2(n874), .ZN(G162) );
  XNOR2_X1 U977 ( .A(G160), .B(n876), .ZN(n885) );
  NAND2_X1 U978 ( .A1(G127), .A2(n891), .ZN(n878) );
  NAND2_X1 U979 ( .A1(G115), .A2(n892), .ZN(n877) );
  NAND2_X1 U980 ( .A1(n878), .A2(n877), .ZN(n879) );
  XNOR2_X1 U981 ( .A(n879), .B(KEYINPUT47), .ZN(n881) );
  NAND2_X1 U982 ( .A1(G139), .A2(n688), .ZN(n880) );
  NAND2_X1 U983 ( .A1(n881), .A2(n880), .ZN(n884) );
  NAND2_X1 U984 ( .A1(n895), .A2(G103), .ZN(n882) );
  XOR2_X1 U985 ( .A(KEYINPUT112), .B(n882), .Z(n883) );
  NOR2_X1 U986 ( .A1(n884), .A2(n883), .ZN(n917) );
  XNOR2_X1 U987 ( .A(n885), .B(n917), .ZN(n890) );
  XOR2_X1 U988 ( .A(KEYINPUT113), .B(KEYINPUT114), .Z(n887) );
  XNOR2_X1 U989 ( .A(KEYINPUT46), .B(KEYINPUT48), .ZN(n886) );
  XNOR2_X1 U990 ( .A(n887), .B(n886), .ZN(n888) );
  XNOR2_X1 U991 ( .A(n888), .B(n925), .ZN(n889) );
  XOR2_X1 U992 ( .A(n890), .B(n889), .Z(n905) );
  NAND2_X1 U993 ( .A1(G130), .A2(n891), .ZN(n894) );
  NAND2_X1 U994 ( .A1(G118), .A2(n892), .ZN(n893) );
  NAND2_X1 U995 ( .A1(n894), .A2(n893), .ZN(n900) );
  NAND2_X1 U996 ( .A1(n895), .A2(G106), .ZN(n897) );
  NAND2_X1 U997 ( .A1(G142), .A2(n688), .ZN(n896) );
  NAND2_X1 U998 ( .A1(n897), .A2(n896), .ZN(n898) );
  XOR2_X1 U999 ( .A(n898), .B(KEYINPUT45), .Z(n899) );
  NOR2_X1 U1000 ( .A1(n900), .A2(n899), .ZN(n902) );
  XNOR2_X1 U1001 ( .A(n902), .B(n901), .ZN(n903) );
  XNOR2_X1 U1002 ( .A(G164), .B(n903), .ZN(n904) );
  XNOR2_X1 U1003 ( .A(n905), .B(n904), .ZN(n908) );
  XNOR2_X1 U1004 ( .A(G162), .B(n906), .ZN(n907) );
  XNOR2_X1 U1005 ( .A(n908), .B(n907), .ZN(n909) );
  NOR2_X1 U1006 ( .A1(G37), .A2(n909), .ZN(G395) );
  NOR2_X1 U1007 ( .A1(G227), .A2(G229), .ZN(n910) );
  XNOR2_X1 U1008 ( .A(KEYINPUT49), .B(n910), .ZN(n911) );
  NOR2_X1 U1009 ( .A1(G401), .A2(n911), .ZN(n914) );
  NOR2_X1 U1010 ( .A1(G397), .A2(n912), .ZN(n913) );
  NAND2_X1 U1011 ( .A1(n914), .A2(n913), .ZN(n915) );
  NOR2_X1 U1012 ( .A1(n915), .A2(G395), .ZN(n916) );
  XNOR2_X1 U1013 ( .A(n916), .B(KEYINPUT115), .ZN(G225) );
  INV_X1 U1014 ( .A(G225), .ZN(G308) );
  INV_X1 U1015 ( .A(KEYINPUT55), .ZN(n961) );
  XNOR2_X1 U1016 ( .A(KEYINPUT52), .B(KEYINPUT116), .ZN(n939) );
  XOR2_X1 U1017 ( .A(G2072), .B(n917), .Z(n919) );
  XOR2_X1 U1018 ( .A(G164), .B(G2078), .Z(n918) );
  NOR2_X1 U1019 ( .A1(n919), .A2(n918), .ZN(n920) );
  XOR2_X1 U1020 ( .A(KEYINPUT50), .B(n920), .Z(n921) );
  NOR2_X1 U1021 ( .A1(n922), .A2(n921), .ZN(n930) );
  XOR2_X1 U1022 ( .A(G160), .B(G2084), .Z(n923) );
  NOR2_X1 U1023 ( .A1(n924), .A2(n923), .ZN(n926) );
  NAND2_X1 U1024 ( .A1(n926), .A2(n925), .ZN(n927) );
  NOR2_X1 U1025 ( .A1(n928), .A2(n927), .ZN(n929) );
  NAND2_X1 U1026 ( .A1(n930), .A2(n929), .ZN(n937) );
  XOR2_X1 U1027 ( .A(G2090), .B(G162), .Z(n931) );
  NOR2_X1 U1028 ( .A1(n932), .A2(n931), .ZN(n933) );
  XOR2_X1 U1029 ( .A(KEYINPUT51), .B(n933), .Z(n935) );
  NAND2_X1 U1030 ( .A1(n935), .A2(n934), .ZN(n936) );
  NOR2_X1 U1031 ( .A1(n937), .A2(n936), .ZN(n938) );
  XNOR2_X1 U1032 ( .A(n939), .B(n938), .ZN(n940) );
  NAND2_X1 U1033 ( .A1(n961), .A2(n940), .ZN(n941) );
  NAND2_X1 U1034 ( .A1(n941), .A2(G29), .ZN(n997) );
  XNOR2_X1 U1035 ( .A(KEYINPUT117), .B(G2090), .ZN(n942) );
  XNOR2_X1 U1036 ( .A(n942), .B(G35), .ZN(n959) );
  XNOR2_X1 U1037 ( .A(G2084), .B(G34), .ZN(n943) );
  XNOR2_X1 U1038 ( .A(n943), .B(KEYINPUT54), .ZN(n957) );
  XOR2_X1 U1039 ( .A(G1991), .B(G25), .Z(n944) );
  NAND2_X1 U1040 ( .A1(n944), .A2(G28), .ZN(n954) );
  XNOR2_X1 U1041 ( .A(G1996), .B(G32), .ZN(n947) );
  XNOR2_X1 U1042 ( .A(n945), .B(G27), .ZN(n946) );
  NOR2_X1 U1043 ( .A1(n947), .A2(n946), .ZN(n948) );
  XNOR2_X1 U1044 ( .A(KEYINPUT118), .B(n948), .ZN(n952) );
  XNOR2_X1 U1045 ( .A(G2067), .B(G26), .ZN(n950) );
  XNOR2_X1 U1046 ( .A(G33), .B(G2072), .ZN(n949) );
  NOR2_X1 U1047 ( .A1(n950), .A2(n949), .ZN(n951) );
  NAND2_X1 U1048 ( .A1(n952), .A2(n951), .ZN(n953) );
  NOR2_X1 U1049 ( .A1(n954), .A2(n953), .ZN(n955) );
  XNOR2_X1 U1050 ( .A(n955), .B(KEYINPUT53), .ZN(n956) );
  NOR2_X1 U1051 ( .A1(n957), .A2(n956), .ZN(n958) );
  NAND2_X1 U1052 ( .A1(n959), .A2(n958), .ZN(n960) );
  XNOR2_X1 U1053 ( .A(n961), .B(n960), .ZN(n963) );
  INV_X1 U1054 ( .A(G29), .ZN(n962) );
  NAND2_X1 U1055 ( .A1(n963), .A2(n962), .ZN(n964) );
  NAND2_X1 U1056 ( .A1(G11), .A2(n964), .ZN(n995) );
  XNOR2_X1 U1057 ( .A(n965), .B(G1348), .ZN(n969) );
  XNOR2_X1 U1058 ( .A(G1961), .B(G301), .ZN(n966) );
  NOR2_X1 U1059 ( .A1(n967), .A2(n966), .ZN(n968) );
  NAND2_X1 U1060 ( .A1(n969), .A2(n968), .ZN(n983) );
  XOR2_X1 U1061 ( .A(n970), .B(G1341), .Z(n981) );
  XNOR2_X1 U1062 ( .A(G1956), .B(KEYINPUT120), .ZN(n971) );
  XNOR2_X1 U1063 ( .A(n971), .B(G299), .ZN(n972) );
  NOR2_X1 U1064 ( .A1(n973), .A2(n972), .ZN(n975) );
  NAND2_X1 U1065 ( .A1(n975), .A2(n974), .ZN(n978) );
  XNOR2_X1 U1066 ( .A(G166), .B(G1971), .ZN(n976) );
  XNOR2_X1 U1067 ( .A(KEYINPUT121), .B(n976), .ZN(n977) );
  NOR2_X1 U1068 ( .A1(n978), .A2(n977), .ZN(n979) );
  XNOR2_X1 U1069 ( .A(KEYINPUT122), .B(n979), .ZN(n980) );
  NAND2_X1 U1070 ( .A1(n981), .A2(n980), .ZN(n982) );
  NOR2_X1 U1071 ( .A1(n983), .A2(n982), .ZN(n984) );
  XNOR2_X1 U1072 ( .A(KEYINPUT123), .B(n984), .ZN(n990) );
  XOR2_X1 U1073 ( .A(G1966), .B(G168), .Z(n985) );
  XNOR2_X1 U1074 ( .A(KEYINPUT119), .B(n985), .ZN(n986) );
  NAND2_X1 U1075 ( .A1(n987), .A2(n986), .ZN(n988) );
  XOR2_X1 U1076 ( .A(KEYINPUT57), .B(n988), .Z(n989) );
  NOR2_X1 U1077 ( .A1(n990), .A2(n989), .ZN(n992) );
  XOR2_X1 U1078 ( .A(G16), .B(KEYINPUT56), .Z(n991) );
  NOR2_X1 U1079 ( .A1(n992), .A2(n991), .ZN(n993) );
  XNOR2_X1 U1080 ( .A(n993), .B(KEYINPUT124), .ZN(n994) );
  NOR2_X1 U1081 ( .A1(n995), .A2(n994), .ZN(n996) );
  NAND2_X1 U1082 ( .A1(n997), .A2(n996), .ZN(n1023) );
  XOR2_X1 U1083 ( .A(KEYINPUT125), .B(G16), .Z(n1021) );
  XOR2_X1 U1084 ( .A(G1976), .B(G23), .Z(n999) );
  XOR2_X1 U1085 ( .A(G1971), .B(G22), .Z(n998) );
  NAND2_X1 U1086 ( .A1(n999), .A2(n998), .ZN(n1001) );
  XNOR2_X1 U1087 ( .A(G24), .B(G1986), .ZN(n1000) );
  NOR2_X1 U1088 ( .A1(n1001), .A2(n1000), .ZN(n1002) );
  XOR2_X1 U1089 ( .A(KEYINPUT58), .B(n1002), .Z(n1018) );
  XOR2_X1 U1090 ( .A(G1961), .B(G5), .Z(n1013) );
  XOR2_X1 U1091 ( .A(G1956), .B(G20), .Z(n1007) );
  XNOR2_X1 U1092 ( .A(G1981), .B(G6), .ZN(n1004) );
  XNOR2_X1 U1093 ( .A(G19), .B(G1341), .ZN(n1003) );
  NOR2_X1 U1094 ( .A1(n1004), .A2(n1003), .ZN(n1005) );
  XNOR2_X1 U1095 ( .A(KEYINPUT126), .B(n1005), .ZN(n1006) );
  NAND2_X1 U1096 ( .A1(n1007), .A2(n1006), .ZN(n1010) );
  XOR2_X1 U1097 ( .A(KEYINPUT59), .B(G1348), .Z(n1008) );
  XNOR2_X1 U1098 ( .A(G4), .B(n1008), .ZN(n1009) );
  NOR2_X1 U1099 ( .A1(n1010), .A2(n1009), .ZN(n1011) );
  XNOR2_X1 U1100 ( .A(KEYINPUT60), .B(n1011), .ZN(n1012) );
  NAND2_X1 U1101 ( .A1(n1013), .A2(n1012), .ZN(n1015) );
  XNOR2_X1 U1102 ( .A(G21), .B(G1966), .ZN(n1014) );
  NOR2_X1 U1103 ( .A1(n1015), .A2(n1014), .ZN(n1016) );
  XNOR2_X1 U1104 ( .A(KEYINPUT127), .B(n1016), .ZN(n1017) );
  NOR2_X1 U1105 ( .A1(n1018), .A2(n1017), .ZN(n1019) );
  XOR2_X1 U1106 ( .A(KEYINPUT61), .B(n1019), .Z(n1020) );
  NOR2_X1 U1107 ( .A1(n1021), .A2(n1020), .ZN(n1022) );
  NOR2_X1 U1108 ( .A1(n1023), .A2(n1022), .ZN(n1024) );
  XNOR2_X1 U1109 ( .A(n1024), .B(KEYINPUT62), .ZN(G311) );
  INV_X1 U1110 ( .A(G311), .ZN(G150) );
endmodule

