//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 1 1 1 0 1 1 0 1 1 1 1 1 1 0 1 0 0 1 1 1 0 0 0 1 1 0 1 0 1 0 0 1 0 1 1 0 1 0 1 0 1 1 1 0 0 0 0 1 0 0 0 0 0 1 0 1 1 1 1 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:17:22 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n658, new_n659,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n696, new_n697, new_n698,
    new_n699, new_n701, new_n702, new_n703, new_n704, new_n705, new_n707,
    new_n708, new_n709, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n716, new_n718, new_n720, new_n721, new_n722, new_n723, new_n724,
    new_n725, new_n726, new_n727, new_n728, new_n729, new_n730, new_n731,
    new_n732, new_n733, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n755, new_n756, new_n757, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n809, new_n810, new_n812, new_n813, new_n814,
    new_n816, new_n817, new_n818, new_n819, new_n820, new_n821, new_n822,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n869, new_n870, new_n871, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n881, new_n882, new_n883, new_n884,
    new_n886, new_n887, new_n888, new_n889, new_n890, new_n891, new_n892,
    new_n893, new_n894, new_n895, new_n896, new_n897, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n920, new_n921, new_n922, new_n923,
    new_n925, new_n926, new_n927, new_n928, new_n929, new_n930, new_n932,
    new_n933, new_n934;
  INV_X1    g000(.A(KEYINPUT25), .ZN(new_n202));
  OAI21_X1  g001(.A(KEYINPUT64), .B1(G183gat), .B2(G190gat), .ZN(new_n203));
  INV_X1    g002(.A(KEYINPUT64), .ZN(new_n204));
  INV_X1    g003(.A(G183gat), .ZN(new_n205));
  INV_X1    g004(.A(G190gat), .ZN(new_n206));
  NAND3_X1  g005(.A1(new_n204), .A2(new_n205), .A3(new_n206), .ZN(new_n207));
  NAND2_X1  g006(.A1(G183gat), .A2(G190gat), .ZN(new_n208));
  INV_X1    g007(.A(KEYINPUT24), .ZN(new_n209));
  NAND2_X1  g008(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  NAND3_X1  g009(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n211));
  AND4_X1   g010(.A1(new_n203), .A2(new_n207), .A3(new_n210), .A4(new_n211), .ZN(new_n212));
  NOR2_X1   g011(.A1(G169gat), .A2(G176gat), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n213), .A2(KEYINPUT23), .ZN(new_n214));
  INV_X1    g013(.A(KEYINPUT23), .ZN(new_n215));
  AOI21_X1  g014(.A(new_n215), .B1(G169gat), .B2(G176gat), .ZN(new_n216));
  OAI21_X1  g015(.A(new_n214), .B1(new_n216), .B2(new_n213), .ZN(new_n217));
  OAI21_X1  g016(.A(new_n202), .B1(new_n212), .B2(new_n217), .ZN(new_n218));
  INV_X1    g017(.A(G169gat), .ZN(new_n219));
  INV_X1    g018(.A(G176gat), .ZN(new_n220));
  OAI21_X1  g019(.A(KEYINPUT23), .B1(new_n219), .B2(new_n220), .ZN(new_n221));
  INV_X1    g020(.A(new_n213), .ZN(new_n222));
  AOI21_X1  g021(.A(new_n202), .B1(new_n221), .B2(new_n222), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n213), .A2(KEYINPUT65), .ZN(new_n224));
  INV_X1    g023(.A(KEYINPUT65), .ZN(new_n225));
  OAI21_X1  g024(.A(new_n225), .B1(G169gat), .B2(G176gat), .ZN(new_n226));
  NAND3_X1  g025(.A1(new_n224), .A2(KEYINPUT23), .A3(new_n226), .ZN(new_n227));
  OAI21_X1  g026(.A(new_n208), .B1(KEYINPUT66), .B2(KEYINPUT24), .ZN(new_n228));
  AND2_X1   g027(.A1(KEYINPUT66), .A2(KEYINPUT24), .ZN(new_n229));
  NOR2_X1   g028(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  OAI21_X1  g029(.A(new_n211), .B1(G183gat), .B2(G190gat), .ZN(new_n231));
  OAI211_X1 g030(.A(new_n223), .B(new_n227), .C1(new_n230), .C2(new_n231), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n218), .A2(new_n232), .ZN(new_n233));
  INV_X1    g032(.A(KEYINPUT26), .ZN(new_n234));
  NAND3_X1  g033(.A1(new_n224), .A2(new_n234), .A3(new_n226), .ZN(new_n235));
  OAI21_X1  g034(.A(new_n234), .B1(new_n219), .B2(new_n220), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n236), .A2(new_n222), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n235), .A2(new_n237), .ZN(new_n238));
  INV_X1    g037(.A(KEYINPUT67), .ZN(new_n239));
  INV_X1    g038(.A(KEYINPUT27), .ZN(new_n240));
  OAI211_X1 g039(.A(new_n239), .B(new_n206), .C1(new_n240), .C2(G183gat), .ZN(new_n241));
  INV_X1    g040(.A(KEYINPUT28), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n241), .A2(new_n242), .ZN(new_n243));
  AOI21_X1  g042(.A(G190gat), .B1(new_n205), .B2(KEYINPUT27), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n240), .A2(G183gat), .ZN(new_n245));
  NAND2_X1  g044(.A1(new_n244), .A2(new_n245), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n243), .A2(new_n246), .ZN(new_n247));
  NAND4_X1  g046(.A1(new_n244), .A2(KEYINPUT67), .A3(new_n242), .A4(new_n245), .ZN(new_n248));
  NAND4_X1  g047(.A1(new_n238), .A2(new_n247), .A3(new_n208), .A4(new_n248), .ZN(new_n249));
  NOR2_X1   g048(.A1(new_n249), .A2(KEYINPUT68), .ZN(new_n250));
  INV_X1    g049(.A(KEYINPUT68), .ZN(new_n251));
  AND4_X1   g050(.A1(KEYINPUT67), .A2(new_n244), .A3(new_n242), .A4(new_n245), .ZN(new_n252));
  AOI22_X1  g051(.A1(new_n241), .A2(new_n242), .B1(new_n244), .B2(new_n245), .ZN(new_n253));
  NOR2_X1   g052(.A1(new_n252), .A2(new_n253), .ZN(new_n254));
  AOI22_X1  g053(.A1(new_n235), .A2(new_n237), .B1(G183gat), .B2(G190gat), .ZN(new_n255));
  AOI21_X1  g054(.A(new_n251), .B1(new_n254), .B2(new_n255), .ZN(new_n256));
  OAI21_X1  g055(.A(new_n233), .B1(new_n250), .B2(new_n256), .ZN(new_n257));
  INV_X1    g056(.A(KEYINPUT69), .ZN(new_n258));
  NAND2_X1  g057(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  XNOR2_X1  g058(.A(G113gat), .B(G120gat), .ZN(new_n260));
  NOR2_X1   g059(.A1(new_n260), .A2(KEYINPUT1), .ZN(new_n261));
  XNOR2_X1  g060(.A(G127gat), .B(G134gat), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  INV_X1    g062(.A(new_n262), .ZN(new_n264));
  OAI21_X1  g063(.A(new_n264), .B1(KEYINPUT1), .B2(new_n260), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n263), .A2(new_n265), .ZN(new_n266));
  OAI211_X1 g065(.A(KEYINPUT69), .B(new_n233), .C1(new_n250), .C2(new_n256), .ZN(new_n267));
  NAND3_X1  g066(.A1(new_n259), .A2(new_n266), .A3(new_n267), .ZN(new_n268));
  INV_X1    g067(.A(G227gat), .ZN(new_n269));
  INV_X1    g068(.A(G233gat), .ZN(new_n270));
  NOR2_X1   g069(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  NAND4_X1  g070(.A1(new_n257), .A2(new_n258), .A3(new_n263), .A4(new_n265), .ZN(new_n272));
  NAND3_X1  g071(.A1(new_n268), .A2(new_n271), .A3(new_n272), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n273), .A2(KEYINPUT70), .ZN(new_n274));
  INV_X1    g073(.A(KEYINPUT70), .ZN(new_n275));
  NAND4_X1  g074(.A1(new_n268), .A2(new_n275), .A3(new_n271), .A4(new_n272), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n274), .A2(new_n276), .ZN(new_n277));
  INV_X1    g076(.A(KEYINPUT33), .ZN(new_n278));
  XOR2_X1   g077(.A(G15gat), .B(G43gat), .Z(new_n279));
  XNOR2_X1  g078(.A(new_n279), .B(KEYINPUT72), .ZN(new_n280));
  XNOR2_X1  g079(.A(G71gat), .B(G99gat), .ZN(new_n281));
  XNOR2_X1  g080(.A(new_n280), .B(new_n281), .ZN(new_n282));
  OAI211_X1 g081(.A(new_n277), .B(KEYINPUT32), .C1(new_n278), .C2(new_n282), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n268), .A2(new_n272), .ZN(new_n284));
  INV_X1    g083(.A(new_n271), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  AND2_X1   g085(.A1(new_n286), .A2(KEYINPUT34), .ZN(new_n287));
  NOR2_X1   g086(.A1(new_n286), .A2(KEYINPUT34), .ZN(new_n288));
  NOR2_X1   g087(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  AOI21_X1  g088(.A(new_n282), .B1(new_n277), .B2(KEYINPUT32), .ZN(new_n290));
  NAND3_X1  g089(.A1(new_n277), .A2(KEYINPUT71), .A3(new_n278), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  AOI21_X1  g091(.A(KEYINPUT33), .B1(new_n274), .B2(new_n276), .ZN(new_n293));
  NOR2_X1   g092(.A1(new_n293), .A2(KEYINPUT71), .ZN(new_n294));
  OAI211_X1 g093(.A(new_n283), .B(new_n289), .C1(new_n292), .C2(new_n294), .ZN(new_n295));
  AND2_X1   g094(.A1(G226gat), .A2(G233gat), .ZN(new_n296));
  NOR2_X1   g095(.A1(new_n296), .A2(KEYINPUT29), .ZN(new_n297));
  INV_X1    g096(.A(new_n297), .ZN(new_n298));
  AOI21_X1  g097(.A(new_n298), .B1(new_n233), .B2(new_n249), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n249), .A2(KEYINPUT68), .ZN(new_n300));
  NAND3_X1  g099(.A1(new_n254), .A2(new_n251), .A3(new_n255), .ZN(new_n301));
  AOI22_X1  g100(.A1(new_n300), .A2(new_n301), .B1(new_n218), .B2(new_n232), .ZN(new_n302));
  AOI21_X1  g101(.A(new_n299), .B1(new_n302), .B2(new_n296), .ZN(new_n303));
  XNOR2_X1  g102(.A(G197gat), .B(G204gat), .ZN(new_n304));
  INV_X1    g103(.A(KEYINPUT22), .ZN(new_n305));
  INV_X1    g104(.A(G211gat), .ZN(new_n306));
  INV_X1    g105(.A(G218gat), .ZN(new_n307));
  OAI21_X1  g106(.A(new_n305), .B1(new_n306), .B2(new_n307), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n304), .A2(new_n308), .ZN(new_n309));
  XNOR2_X1  g108(.A(G211gat), .B(G218gat), .ZN(new_n310));
  INV_X1    g109(.A(new_n310), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n309), .A2(new_n311), .ZN(new_n312));
  NAND3_X1  g111(.A1(new_n310), .A2(new_n304), .A3(new_n308), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  INV_X1    g113(.A(new_n314), .ZN(new_n315));
  OAI21_X1  g114(.A(KEYINPUT75), .B1(new_n303), .B2(new_n315), .ZN(new_n316));
  OAI211_X1 g115(.A(new_n296), .B(new_n233), .C1(new_n250), .C2(new_n256), .ZN(new_n317));
  INV_X1    g116(.A(new_n299), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n317), .A2(new_n318), .ZN(new_n319));
  INV_X1    g118(.A(KEYINPUT75), .ZN(new_n320));
  NAND3_X1  g119(.A1(new_n319), .A2(new_n320), .A3(new_n314), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n316), .A2(new_n321), .ZN(new_n322));
  NAND3_X1  g121(.A1(new_n233), .A2(new_n296), .A3(new_n249), .ZN(new_n323));
  OAI211_X1 g122(.A(new_n315), .B(new_n323), .C1(new_n302), .C2(new_n298), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n324), .A2(KEYINPUT74), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n257), .A2(new_n297), .ZN(new_n326));
  INV_X1    g125(.A(KEYINPUT74), .ZN(new_n327));
  NAND4_X1  g126(.A1(new_n326), .A2(new_n327), .A3(new_n315), .A4(new_n323), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n325), .A2(new_n328), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n322), .A2(new_n329), .ZN(new_n330));
  XOR2_X1   g129(.A(G8gat), .B(G36gat), .Z(new_n331));
  XNOR2_X1  g130(.A(new_n331), .B(KEYINPUT76), .ZN(new_n332));
  XNOR2_X1  g131(.A(G64gat), .B(G92gat), .ZN(new_n333));
  XOR2_X1   g132(.A(new_n332), .B(new_n333), .Z(new_n334));
  NAND2_X1  g133(.A1(new_n330), .A2(new_n334), .ZN(new_n335));
  INV_X1    g134(.A(new_n334), .ZN(new_n336));
  NAND3_X1  g135(.A1(new_n322), .A2(new_n329), .A3(new_n336), .ZN(new_n337));
  INV_X1    g136(.A(KEYINPUT78), .ZN(new_n338));
  INV_X1    g137(.A(KEYINPUT30), .ZN(new_n339));
  AND3_X1   g138(.A1(new_n337), .A2(new_n338), .A3(new_n339), .ZN(new_n340));
  AOI21_X1  g139(.A(new_n338), .B1(new_n337), .B2(new_n339), .ZN(new_n341));
  OAI21_X1  g140(.A(new_n335), .B1(new_n340), .B2(new_n341), .ZN(new_n342));
  NAND4_X1  g141(.A1(new_n322), .A2(new_n329), .A3(KEYINPUT30), .A4(new_n336), .ZN(new_n343));
  INV_X1    g142(.A(KEYINPUT77), .ZN(new_n344));
  XNOR2_X1  g143(.A(new_n343), .B(new_n344), .ZN(new_n345));
  XOR2_X1   g144(.A(G141gat), .B(G148gat), .Z(new_n346));
  INV_X1    g145(.A(G155gat), .ZN(new_n347));
  INV_X1    g146(.A(G162gat), .ZN(new_n348));
  OAI21_X1  g147(.A(KEYINPUT2), .B1(new_n347), .B2(new_n348), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n346), .A2(new_n349), .ZN(new_n350));
  XNOR2_X1  g149(.A(G155gat), .B(G162gat), .ZN(new_n351));
  INV_X1    g150(.A(new_n351), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n350), .A2(new_n352), .ZN(new_n353));
  NAND3_X1  g152(.A1(new_n346), .A2(new_n351), .A3(new_n349), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n355), .A2(KEYINPUT3), .ZN(new_n356));
  INV_X1    g155(.A(KEYINPUT3), .ZN(new_n357));
  NAND3_X1  g156(.A1(new_n353), .A2(new_n357), .A3(new_n354), .ZN(new_n358));
  NAND3_X1  g157(.A1(new_n356), .A2(new_n266), .A3(new_n358), .ZN(new_n359));
  NAND4_X1  g158(.A1(new_n353), .A2(new_n263), .A3(new_n354), .A4(new_n265), .ZN(new_n360));
  INV_X1    g159(.A(new_n360), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n361), .A2(KEYINPUT4), .ZN(new_n362));
  NAND2_X1  g161(.A1(G225gat), .A2(G233gat), .ZN(new_n363));
  XNOR2_X1  g162(.A(new_n363), .B(KEYINPUT79), .ZN(new_n364));
  INV_X1    g163(.A(new_n364), .ZN(new_n365));
  INV_X1    g164(.A(KEYINPUT4), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n360), .A2(new_n366), .ZN(new_n367));
  NAND4_X1  g166(.A1(new_n359), .A2(new_n362), .A3(new_n365), .A4(new_n367), .ZN(new_n368));
  AOI22_X1  g167(.A1(new_n353), .A2(new_n354), .B1(new_n263), .B2(new_n265), .ZN(new_n369));
  OAI21_X1  g168(.A(new_n364), .B1(new_n361), .B2(new_n369), .ZN(new_n370));
  XOR2_X1   g169(.A(KEYINPUT80), .B(KEYINPUT5), .Z(new_n371));
  INV_X1    g170(.A(new_n371), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n370), .A2(new_n372), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n368), .A2(new_n373), .ZN(new_n374));
  XNOR2_X1  g173(.A(new_n360), .B(KEYINPUT4), .ZN(new_n375));
  NAND4_X1  g174(.A1(new_n375), .A2(new_n365), .A3(new_n359), .A4(new_n372), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n374), .A2(new_n376), .ZN(new_n377));
  XOR2_X1   g176(.A(G1gat), .B(G29gat), .Z(new_n378));
  XNOR2_X1  g177(.A(G57gat), .B(G85gat), .ZN(new_n379));
  XNOR2_X1  g178(.A(new_n378), .B(new_n379), .ZN(new_n380));
  XNOR2_X1  g179(.A(KEYINPUT81), .B(KEYINPUT0), .ZN(new_n381));
  XNOR2_X1  g180(.A(new_n380), .B(new_n381), .ZN(new_n382));
  INV_X1    g181(.A(new_n382), .ZN(new_n383));
  NOR2_X1   g182(.A1(new_n377), .A2(new_n383), .ZN(new_n384));
  AOI21_X1  g183(.A(new_n382), .B1(new_n374), .B2(new_n376), .ZN(new_n385));
  NOR3_X1   g184(.A1(new_n384), .A2(new_n385), .A3(KEYINPUT6), .ZN(new_n386));
  INV_X1    g185(.A(KEYINPUT6), .ZN(new_n387));
  NOR3_X1   g186(.A1(new_n377), .A2(new_n387), .A3(new_n383), .ZN(new_n388));
  NOR2_X1   g187(.A1(new_n386), .A2(new_n388), .ZN(new_n389));
  NOR4_X1   g188(.A1(new_n342), .A2(new_n345), .A3(KEYINPUT35), .A4(new_n389), .ZN(new_n390));
  OAI21_X1  g189(.A(new_n283), .B1(new_n292), .B2(new_n294), .ZN(new_n391));
  INV_X1    g190(.A(new_n289), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n391), .A2(new_n392), .ZN(new_n393));
  INV_X1    g192(.A(G228gat), .ZN(new_n394));
  NOR2_X1   g193(.A1(new_n394), .A2(new_n270), .ZN(new_n395));
  INV_X1    g194(.A(KEYINPUT29), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n358), .A2(new_n396), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n397), .A2(new_n315), .ZN(new_n398));
  INV_X1    g197(.A(KEYINPUT84), .ZN(new_n399));
  AOI21_X1  g198(.A(new_n395), .B1(new_n398), .B2(new_n399), .ZN(new_n400));
  AOI21_X1  g199(.A(KEYINPUT29), .B1(new_n312), .B2(new_n313), .ZN(new_n401));
  OAI21_X1  g200(.A(new_n355), .B1(new_n401), .B2(KEYINPUT3), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n398), .A2(new_n402), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n400), .A2(new_n403), .ZN(new_n404));
  INV_X1    g203(.A(G22gat), .ZN(new_n405));
  OAI211_X1 g204(.A(new_n398), .B(new_n402), .C1(new_n399), .C2(new_n395), .ZN(new_n406));
  NAND3_X1  g205(.A1(new_n404), .A2(new_n405), .A3(new_n406), .ZN(new_n407));
  INV_X1    g206(.A(KEYINPUT85), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n407), .A2(new_n408), .ZN(new_n409));
  NAND4_X1  g208(.A1(new_n404), .A2(KEYINPUT85), .A3(new_n405), .A4(new_n406), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n404), .A2(new_n406), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n411), .A2(G22gat), .ZN(new_n412));
  NAND3_X1  g211(.A1(new_n409), .A2(new_n410), .A3(new_n412), .ZN(new_n413));
  XNOR2_X1  g212(.A(G78gat), .B(G106gat), .ZN(new_n414));
  INV_X1    g213(.A(G50gat), .ZN(new_n415));
  XNOR2_X1  g214(.A(new_n414), .B(new_n415), .ZN(new_n416));
  XOR2_X1   g215(.A(KEYINPUT82), .B(KEYINPUT31), .Z(new_n417));
  XNOR2_X1  g216(.A(new_n416), .B(new_n417), .ZN(new_n418));
  XNOR2_X1  g217(.A(new_n418), .B(KEYINPUT83), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n413), .A2(new_n419), .ZN(new_n420));
  INV_X1    g219(.A(new_n418), .ZN(new_n421));
  NAND3_X1  g220(.A1(new_n412), .A2(new_n407), .A3(new_n421), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n420), .A2(new_n422), .ZN(new_n423));
  AND4_X1   g222(.A1(new_n295), .A2(new_n390), .A3(new_n393), .A4(new_n423), .ZN(new_n424));
  INV_X1    g223(.A(KEYINPUT73), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n391), .A2(new_n425), .ZN(new_n426));
  OR2_X1    g225(.A1(new_n293), .A2(KEYINPUT71), .ZN(new_n427));
  NAND3_X1  g226(.A1(new_n427), .A2(new_n291), .A3(new_n290), .ZN(new_n428));
  NAND3_X1  g227(.A1(new_n428), .A2(KEYINPUT73), .A3(new_n283), .ZN(new_n429));
  NAND3_X1  g228(.A1(new_n426), .A2(new_n429), .A3(new_n392), .ZN(new_n430));
  NOR2_X1   g229(.A1(new_n342), .A2(new_n345), .ZN(new_n431));
  INV_X1    g230(.A(new_n431), .ZN(new_n432));
  NOR2_X1   g231(.A1(new_n432), .A2(new_n389), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n295), .A2(new_n423), .ZN(new_n434));
  INV_X1    g233(.A(new_n434), .ZN(new_n435));
  NAND3_X1  g234(.A1(new_n430), .A2(new_n433), .A3(new_n435), .ZN(new_n436));
  AOI21_X1  g235(.A(new_n424), .B1(new_n436), .B2(KEYINPUT35), .ZN(new_n437));
  NOR4_X1   g236(.A1(new_n342), .A2(new_n345), .A3(new_n423), .A4(new_n389), .ZN(new_n438));
  INV_X1    g237(.A(KEYINPUT86), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n375), .A2(new_n359), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n440), .A2(new_n364), .ZN(new_n441));
  OAI21_X1  g240(.A(new_n383), .B1(new_n441), .B2(KEYINPUT39), .ZN(new_n442));
  OR2_X1    g241(.A1(new_n361), .A2(new_n369), .ZN(new_n443));
  OAI21_X1  g242(.A(KEYINPUT39), .B1(new_n443), .B2(new_n364), .ZN(new_n444));
  AOI21_X1  g243(.A(new_n444), .B1(new_n364), .B2(new_n440), .ZN(new_n445));
  OAI21_X1  g244(.A(new_n439), .B1(new_n442), .B2(new_n445), .ZN(new_n446));
  AOI21_X1  g245(.A(new_n384), .B1(new_n446), .B2(KEYINPUT40), .ZN(new_n447));
  INV_X1    g246(.A(KEYINPUT40), .ZN(new_n448));
  OAI211_X1 g247(.A(new_n439), .B(new_n448), .C1(new_n442), .C2(new_n445), .ZN(new_n449));
  AND2_X1   g248(.A1(new_n447), .A2(new_n449), .ZN(new_n450));
  OAI21_X1  g249(.A(new_n450), .B1(new_n342), .B2(new_n345), .ZN(new_n451));
  XNOR2_X1  g250(.A(KEYINPUT87), .B(KEYINPUT37), .ZN(new_n452));
  NAND3_X1  g251(.A1(new_n322), .A2(new_n329), .A3(new_n452), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n453), .A2(new_n334), .ZN(new_n454));
  INV_X1    g253(.A(KEYINPUT37), .ZN(new_n455));
  AOI21_X1  g254(.A(new_n455), .B1(new_n322), .B2(new_n329), .ZN(new_n456));
  OAI21_X1  g255(.A(KEYINPUT38), .B1(new_n454), .B2(new_n456), .ZN(new_n457));
  AOI21_X1  g256(.A(new_n455), .B1(new_n319), .B2(new_n315), .ZN(new_n458));
  NAND3_X1  g257(.A1(new_n326), .A2(new_n314), .A3(new_n323), .ZN(new_n459));
  AOI21_X1  g258(.A(KEYINPUT38), .B1(new_n458), .B2(new_n459), .ZN(new_n460));
  NAND3_X1  g259(.A1(new_n453), .A2(new_n334), .A3(new_n460), .ZN(new_n461));
  NAND4_X1  g260(.A1(new_n457), .A2(new_n389), .A3(new_n337), .A4(new_n461), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n451), .A2(new_n462), .ZN(new_n463));
  AOI21_X1  g262(.A(new_n438), .B1(new_n463), .B2(new_n423), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n295), .A2(KEYINPUT36), .ZN(new_n465));
  INV_X1    g264(.A(new_n465), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n430), .A2(new_n466), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n393), .A2(new_n295), .ZN(new_n468));
  INV_X1    g267(.A(KEYINPUT36), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  AOI21_X1  g269(.A(new_n464), .B1(new_n467), .B2(new_n470), .ZN(new_n471));
  NOR2_X1   g270(.A1(new_n437), .A2(new_n471), .ZN(new_n472));
  INV_X1    g271(.A(KEYINPUT14), .ZN(new_n473));
  INV_X1    g272(.A(G29gat), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  NAND2_X1  g274(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n476));
  AOI21_X1  g275(.A(G36gat), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  INV_X1    g276(.A(G36gat), .ZN(new_n478));
  NOR3_X1   g277(.A1(new_n473), .A2(new_n478), .A3(G29gat), .ZN(new_n479));
  OR3_X1    g278(.A1(new_n477), .A2(KEYINPUT15), .A3(new_n479), .ZN(new_n480));
  OAI21_X1  g279(.A(KEYINPUT15), .B1(new_n477), .B2(new_n479), .ZN(new_n481));
  XNOR2_X1  g280(.A(G43gat), .B(G50gat), .ZN(new_n482));
  NAND3_X1  g281(.A1(new_n480), .A2(new_n481), .A3(new_n482), .ZN(new_n483));
  OR2_X1    g282(.A1(new_n481), .A2(new_n482), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  INV_X1    g284(.A(KEYINPUT17), .ZN(new_n486));
  OAI21_X1  g285(.A(new_n485), .B1(KEYINPUT89), .B2(new_n486), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n486), .A2(KEYINPUT89), .ZN(new_n488));
  INV_X1    g287(.A(new_n488), .ZN(new_n489));
  XNOR2_X1  g288(.A(new_n487), .B(new_n489), .ZN(new_n490));
  XNOR2_X1  g289(.A(G15gat), .B(G22gat), .ZN(new_n491));
  INV_X1    g290(.A(KEYINPUT16), .ZN(new_n492));
  OAI21_X1  g291(.A(new_n491), .B1(new_n492), .B2(G1gat), .ZN(new_n493));
  OAI211_X1 g292(.A(new_n493), .B(KEYINPUT90), .C1(G1gat), .C2(new_n491), .ZN(new_n494));
  XOR2_X1   g293(.A(new_n494), .B(G8gat), .Z(new_n495));
  NAND2_X1  g294(.A1(new_n490), .A2(new_n495), .ZN(new_n496));
  NAND2_X1  g295(.A1(G229gat), .A2(G233gat), .ZN(new_n497));
  INV_X1    g296(.A(new_n495), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n498), .A2(new_n485), .ZN(new_n499));
  NAND3_X1  g298(.A1(new_n496), .A2(new_n497), .A3(new_n499), .ZN(new_n500));
  INV_X1    g299(.A(KEYINPUT18), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n502), .A2(KEYINPUT91), .ZN(new_n503));
  INV_X1    g302(.A(KEYINPUT91), .ZN(new_n504));
  NAND3_X1  g303(.A1(new_n500), .A2(new_n504), .A3(new_n501), .ZN(new_n505));
  AND2_X1   g304(.A1(new_n503), .A2(new_n505), .ZN(new_n506));
  XOR2_X1   g305(.A(new_n495), .B(new_n485), .Z(new_n507));
  XOR2_X1   g306(.A(new_n497), .B(KEYINPUT13), .Z(new_n508));
  NAND2_X1  g307(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  OAI21_X1  g308(.A(new_n509), .B1(new_n500), .B2(new_n501), .ZN(new_n510));
  XOR2_X1   g309(.A(G113gat), .B(G141gat), .Z(new_n511));
  XNOR2_X1  g310(.A(KEYINPUT88), .B(G197gat), .ZN(new_n512));
  XNOR2_X1  g311(.A(new_n511), .B(new_n512), .ZN(new_n513));
  XNOR2_X1  g312(.A(KEYINPUT11), .B(G169gat), .ZN(new_n514));
  XOR2_X1   g313(.A(new_n513), .B(new_n514), .Z(new_n515));
  XOR2_X1   g314(.A(new_n515), .B(KEYINPUT12), .Z(new_n516));
  NOR2_X1   g315(.A1(new_n510), .A2(new_n516), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n506), .A2(new_n517), .ZN(new_n518));
  INV_X1    g317(.A(new_n502), .ZN(new_n519));
  OAI21_X1  g318(.A(new_n516), .B1(new_n519), .B2(new_n510), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n518), .A2(new_n520), .ZN(new_n521));
  INV_X1    g320(.A(new_n521), .ZN(new_n522));
  NOR2_X1   g321(.A1(new_n472), .A2(new_n522), .ZN(new_n523));
  XNOR2_X1  g322(.A(KEYINPUT96), .B(KEYINPUT97), .ZN(new_n524));
  INV_X1    g323(.A(new_n524), .ZN(new_n525));
  NAND2_X1  g324(.A1(G85gat), .A2(G92gat), .ZN(new_n526));
  XNOR2_X1  g325(.A(new_n526), .B(KEYINPUT7), .ZN(new_n527));
  INV_X1    g326(.A(G99gat), .ZN(new_n528));
  INV_X1    g327(.A(G106gat), .ZN(new_n529));
  OAI21_X1  g328(.A(KEYINPUT8), .B1(new_n528), .B2(new_n529), .ZN(new_n530));
  XOR2_X1   g329(.A(KEYINPUT98), .B(G92gat), .Z(new_n531));
  OAI211_X1 g330(.A(new_n527), .B(new_n530), .C1(G85gat), .C2(new_n531), .ZN(new_n532));
  XOR2_X1   g331(.A(G99gat), .B(G106gat), .Z(new_n533));
  OR2_X1    g332(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n532), .A2(new_n533), .ZN(new_n535));
  NAND3_X1  g334(.A1(new_n534), .A2(KEYINPUT99), .A3(new_n535), .ZN(new_n536));
  INV_X1    g335(.A(KEYINPUT99), .ZN(new_n537));
  NAND3_X1  g336(.A1(new_n532), .A2(new_n537), .A3(new_n533), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n536), .A2(new_n538), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n539), .A2(new_n485), .ZN(new_n540));
  INV_X1    g339(.A(KEYINPUT41), .ZN(new_n541));
  INV_X1    g340(.A(G232gat), .ZN(new_n542));
  NOR3_X1   g341(.A1(new_n541), .A2(new_n542), .A3(new_n270), .ZN(new_n543));
  INV_X1    g342(.A(new_n543), .ZN(new_n544));
  NAND2_X1  g343(.A1(new_n540), .A2(new_n544), .ZN(new_n545));
  AND2_X1   g344(.A1(new_n545), .A2(KEYINPUT101), .ZN(new_n546));
  NOR2_X1   g345(.A1(new_n545), .A2(KEYINPUT101), .ZN(new_n547));
  OR2_X1    g346(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  NAND2_X1  g347(.A1(new_n539), .A2(KEYINPUT100), .ZN(new_n549));
  OR2_X1    g348(.A1(new_n539), .A2(KEYINPUT100), .ZN(new_n550));
  NAND3_X1  g349(.A1(new_n490), .A2(new_n549), .A3(new_n550), .ZN(new_n551));
  AOI21_X1  g350(.A(new_n525), .B1(new_n548), .B2(new_n551), .ZN(new_n552));
  INV_X1    g351(.A(new_n552), .ZN(new_n553));
  OAI211_X1 g352(.A(new_n551), .B(new_n525), .C1(new_n546), .C2(new_n547), .ZN(new_n554));
  XOR2_X1   g353(.A(G190gat), .B(G218gat), .Z(new_n555));
  XNOR2_X1  g354(.A(new_n555), .B(KEYINPUT102), .ZN(new_n556));
  XNOR2_X1  g355(.A(G134gat), .B(G162gat), .ZN(new_n557));
  OAI21_X1  g356(.A(new_n541), .B1(new_n542), .B2(new_n270), .ZN(new_n558));
  XNOR2_X1  g357(.A(new_n557), .B(new_n558), .ZN(new_n559));
  XOR2_X1   g358(.A(new_n556), .B(new_n559), .Z(new_n560));
  NAND3_X1  g359(.A1(new_n553), .A2(new_n554), .A3(new_n560), .ZN(new_n561));
  INV_X1    g360(.A(new_n560), .ZN(new_n562));
  INV_X1    g361(.A(new_n554), .ZN(new_n563));
  OAI21_X1  g362(.A(new_n562), .B1(new_n552), .B2(new_n563), .ZN(new_n564));
  NAND2_X1  g363(.A1(new_n561), .A2(new_n564), .ZN(new_n565));
  INV_X1    g364(.A(new_n565), .ZN(new_n566));
  INV_X1    g365(.A(KEYINPUT21), .ZN(new_n567));
  XOR2_X1   g366(.A(G57gat), .B(G64gat), .Z(new_n568));
  NAND2_X1  g367(.A1(G71gat), .A2(G78gat), .ZN(new_n569));
  INV_X1    g368(.A(new_n569), .ZN(new_n570));
  OAI21_X1  g369(.A(new_n568), .B1(KEYINPUT9), .B2(new_n570), .ZN(new_n571));
  NOR2_X1   g370(.A1(G71gat), .A2(G78gat), .ZN(new_n572));
  INV_X1    g371(.A(KEYINPUT92), .ZN(new_n573));
  AOI21_X1  g372(.A(new_n572), .B1(new_n573), .B2(new_n569), .ZN(new_n574));
  OAI211_X1 g373(.A(new_n571), .B(new_n574), .C1(new_n573), .C2(new_n569), .ZN(new_n575));
  INV_X1    g374(.A(G57gat), .ZN(new_n576));
  INV_X1    g375(.A(G64gat), .ZN(new_n577));
  OR3_X1    g376(.A1(new_n576), .A2(new_n577), .A3(KEYINPUT93), .ZN(new_n578));
  OAI21_X1  g377(.A(new_n577), .B1(new_n576), .B2(KEYINPUT93), .ZN(new_n579));
  AND2_X1   g378(.A1(new_n572), .A2(KEYINPUT9), .ZN(new_n580));
  OAI211_X1 g379(.A(new_n578), .B(new_n579), .C1(new_n580), .C2(new_n570), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n575), .A2(new_n581), .ZN(new_n582));
  OAI21_X1  g381(.A(new_n495), .B1(new_n567), .B2(new_n582), .ZN(new_n583));
  XNOR2_X1  g382(.A(new_n583), .B(KEYINPUT95), .ZN(new_n584));
  NAND2_X1  g383(.A1(G231gat), .A2(G233gat), .ZN(new_n585));
  XNOR2_X1  g384(.A(new_n585), .B(KEYINPUT94), .ZN(new_n586));
  XOR2_X1   g385(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n587));
  XOR2_X1   g386(.A(new_n586), .B(new_n587), .Z(new_n588));
  XNOR2_X1  g387(.A(new_n584), .B(new_n588), .ZN(new_n589));
  NAND2_X1  g388(.A1(new_n582), .A2(new_n567), .ZN(new_n590));
  XOR2_X1   g389(.A(G127gat), .B(G155gat), .Z(new_n591));
  XNOR2_X1  g390(.A(new_n590), .B(new_n591), .ZN(new_n592));
  XOR2_X1   g391(.A(G183gat), .B(G211gat), .Z(new_n593));
  XNOR2_X1  g392(.A(new_n592), .B(new_n593), .ZN(new_n594));
  INV_X1    g393(.A(new_n594), .ZN(new_n595));
  OR2_X1    g394(.A1(new_n589), .A2(new_n595), .ZN(new_n596));
  NAND2_X1  g395(.A1(new_n589), .A2(new_n595), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  INV_X1    g397(.A(new_n598), .ZN(new_n599));
  INV_X1    g398(.A(new_n539), .ZN(new_n600));
  NAND2_X1  g399(.A1(new_n600), .A2(new_n582), .ZN(new_n601));
  INV_X1    g400(.A(KEYINPUT10), .ZN(new_n602));
  INV_X1    g401(.A(new_n582), .ZN(new_n603));
  NAND3_X1  g402(.A1(new_n603), .A2(new_n535), .A3(new_n534), .ZN(new_n604));
  NAND3_X1  g403(.A1(new_n601), .A2(new_n602), .A3(new_n604), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n603), .A2(KEYINPUT10), .ZN(new_n606));
  OR3_X1    g405(.A1(new_n600), .A2(KEYINPUT103), .A3(new_n606), .ZN(new_n607));
  OAI21_X1  g406(.A(KEYINPUT103), .B1(new_n600), .B2(new_n606), .ZN(new_n608));
  NAND3_X1  g407(.A1(new_n605), .A2(new_n607), .A3(new_n608), .ZN(new_n609));
  NAND2_X1  g408(.A1(G230gat), .A2(G233gat), .ZN(new_n610));
  NAND2_X1  g409(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  NAND2_X1  g410(.A1(new_n601), .A2(new_n604), .ZN(new_n612));
  INV_X1    g411(.A(new_n610), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n611), .A2(new_n614), .ZN(new_n615));
  XNOR2_X1  g414(.A(G120gat), .B(G148gat), .ZN(new_n616));
  XNOR2_X1  g415(.A(G176gat), .B(G204gat), .ZN(new_n617));
  XOR2_X1   g416(.A(new_n616), .B(new_n617), .Z(new_n618));
  INV_X1    g417(.A(new_n618), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n615), .A2(new_n619), .ZN(new_n620));
  NAND3_X1  g419(.A1(new_n611), .A2(new_n614), .A3(new_n618), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  INV_X1    g421(.A(new_n622), .ZN(new_n623));
  NAND3_X1  g422(.A1(new_n566), .A2(new_n599), .A3(new_n623), .ZN(new_n624));
  INV_X1    g423(.A(new_n624), .ZN(new_n625));
  XNOR2_X1  g424(.A(new_n389), .B(KEYINPUT104), .ZN(new_n626));
  NAND3_X1  g425(.A1(new_n523), .A2(new_n625), .A3(new_n626), .ZN(new_n627));
  XNOR2_X1  g426(.A(new_n627), .B(G1gat), .ZN(G1324gat));
  XOR2_X1   g427(.A(KEYINPUT16), .B(G8gat), .Z(new_n629));
  NAND4_X1  g428(.A1(new_n523), .A2(new_n432), .A3(new_n625), .A4(new_n629), .ZN(new_n630));
  AOI21_X1  g429(.A(new_n289), .B1(new_n391), .B2(new_n425), .ZN(new_n631));
  AOI21_X1  g430(.A(new_n465), .B1(new_n631), .B2(new_n429), .ZN(new_n632));
  AOI21_X1  g431(.A(KEYINPUT36), .B1(new_n393), .B2(new_n295), .ZN(new_n633));
  INV_X1    g432(.A(new_n423), .ZN(new_n634));
  AOI21_X1  g433(.A(new_n634), .B1(new_n451), .B2(new_n462), .ZN(new_n635));
  OAI22_X1  g434(.A1(new_n632), .A2(new_n633), .B1(new_n635), .B2(new_n438), .ZN(new_n636));
  INV_X1    g435(.A(KEYINPUT35), .ZN(new_n637));
  AOI21_X1  g436(.A(new_n434), .B1(new_n631), .B2(new_n429), .ZN(new_n638));
  AOI21_X1  g437(.A(new_n637), .B1(new_n638), .B2(new_n433), .ZN(new_n639));
  OAI21_X1  g438(.A(new_n636), .B1(new_n639), .B2(new_n424), .ZN(new_n640));
  NAND3_X1  g439(.A1(new_n640), .A2(new_n432), .A3(new_n521), .ZN(new_n641));
  OAI21_X1  g440(.A(G8gat), .B1(new_n641), .B2(new_n624), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n630), .A2(new_n642), .ZN(new_n643));
  NAND2_X1  g442(.A1(new_n643), .A2(KEYINPUT42), .ZN(new_n644));
  INV_X1    g443(.A(KEYINPUT105), .ZN(new_n645));
  INV_X1    g444(.A(KEYINPUT42), .ZN(new_n646));
  NAND2_X1  g445(.A1(new_n630), .A2(new_n646), .ZN(new_n647));
  AND3_X1   g446(.A1(new_n644), .A2(new_n645), .A3(new_n647), .ZN(new_n648));
  AOI21_X1  g447(.A(new_n645), .B1(new_n644), .B2(new_n647), .ZN(new_n649));
  NOR2_X1   g448(.A1(new_n648), .A2(new_n649), .ZN(G1325gat));
  NAND2_X1  g449(.A1(new_n523), .A2(new_n625), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n467), .A2(new_n470), .ZN(new_n652));
  OAI21_X1  g451(.A(G15gat), .B1(new_n651), .B2(new_n652), .ZN(new_n653));
  INV_X1    g452(.A(new_n468), .ZN(new_n654));
  NOR2_X1   g453(.A1(new_n624), .A2(G15gat), .ZN(new_n655));
  NAND3_X1  g454(.A1(new_n523), .A2(new_n654), .A3(new_n655), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n653), .A2(new_n656), .ZN(G1326gat));
  NOR2_X1   g456(.A1(new_n651), .A2(new_n423), .ZN(new_n658));
  XOR2_X1   g457(.A(KEYINPUT43), .B(G22gat), .Z(new_n659));
  XNOR2_X1  g458(.A(new_n658), .B(new_n659), .ZN(G1327gat));
  NOR3_X1   g459(.A1(new_n522), .A2(new_n599), .A3(new_n622), .ZN(new_n661));
  NAND3_X1  g460(.A1(new_n640), .A2(new_n565), .A3(new_n661), .ZN(new_n662));
  INV_X1    g461(.A(new_n662), .ZN(new_n663));
  NAND3_X1  g462(.A1(new_n663), .A2(new_n474), .A3(new_n626), .ZN(new_n664));
  XNOR2_X1  g463(.A(new_n664), .B(KEYINPUT45), .ZN(new_n665));
  OAI21_X1  g464(.A(new_n565), .B1(new_n437), .B2(new_n471), .ZN(new_n666));
  INV_X1    g465(.A(KEYINPUT44), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  NAND3_X1  g467(.A1(new_n640), .A2(KEYINPUT44), .A3(new_n565), .ZN(new_n669));
  AND4_X1   g468(.A1(new_n626), .A2(new_n668), .A3(new_n661), .A4(new_n669), .ZN(new_n670));
  OAI21_X1  g469(.A(new_n665), .B1(new_n474), .B2(new_n670), .ZN(G1328gat));
  NOR3_X1   g470(.A1(new_n566), .A2(new_n599), .A3(new_n622), .ZN(new_n672));
  NAND4_X1  g471(.A1(new_n523), .A2(new_n478), .A3(new_n432), .A4(new_n672), .ZN(new_n673));
  OR2_X1    g472(.A1(new_n673), .A2(KEYINPUT46), .ZN(new_n674));
  NAND4_X1  g473(.A1(new_n668), .A2(new_n432), .A3(new_n669), .A4(new_n661), .ZN(new_n675));
  NAND2_X1  g474(.A1(new_n675), .A2(G36gat), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n673), .A2(KEYINPUT46), .ZN(new_n677));
  NAND3_X1  g476(.A1(new_n674), .A2(new_n676), .A3(new_n677), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n678), .A2(KEYINPUT106), .ZN(new_n679));
  INV_X1    g478(.A(KEYINPUT106), .ZN(new_n680));
  NAND4_X1  g479(.A1(new_n674), .A2(new_n680), .A3(new_n676), .A4(new_n677), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n679), .A2(new_n681), .ZN(G1329gat));
  INV_X1    g481(.A(G43gat), .ZN(new_n683));
  INV_X1    g482(.A(new_n652), .ZN(new_n684));
  NAND4_X1  g483(.A1(new_n668), .A2(new_n684), .A3(new_n669), .A4(new_n661), .ZN(new_n685));
  INV_X1    g484(.A(KEYINPUT108), .ZN(new_n686));
  AOI21_X1  g485(.A(new_n683), .B1(new_n685), .B2(new_n686), .ZN(new_n687));
  OAI21_X1  g486(.A(new_n687), .B1(new_n686), .B2(new_n685), .ZN(new_n688));
  NAND4_X1  g487(.A1(new_n523), .A2(new_n683), .A3(new_n654), .A4(new_n672), .ZN(new_n689));
  NAND3_X1  g488(.A1(new_n688), .A2(KEYINPUT47), .A3(new_n689), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n685), .A2(G43gat), .ZN(new_n691));
  NAND2_X1  g490(.A1(new_n691), .A2(new_n689), .ZN(new_n692));
  XOR2_X1   g491(.A(KEYINPUT107), .B(KEYINPUT47), .Z(new_n693));
  NAND2_X1  g492(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n690), .A2(new_n694), .ZN(G1330gat));
  NAND3_X1  g494(.A1(new_n663), .A2(new_n415), .A3(new_n634), .ZN(new_n696));
  AND4_X1   g495(.A1(new_n634), .A2(new_n668), .A3(new_n661), .A4(new_n669), .ZN(new_n697));
  OAI21_X1  g496(.A(new_n696), .B1(new_n697), .B2(new_n415), .ZN(new_n698));
  INV_X1    g497(.A(KEYINPUT48), .ZN(new_n699));
  XNOR2_X1  g498(.A(new_n698), .B(new_n699), .ZN(G1331gat));
  NAND2_X1  g499(.A1(new_n566), .A2(new_n599), .ZN(new_n701));
  NOR4_X1   g500(.A1(new_n472), .A2(new_n521), .A3(new_n701), .A4(new_n623), .ZN(new_n702));
  XNOR2_X1  g501(.A(new_n626), .B(KEYINPUT109), .ZN(new_n703));
  INV_X1    g502(.A(new_n703), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n702), .A2(new_n704), .ZN(new_n705));
  XNOR2_X1  g504(.A(new_n705), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g505(.A1(new_n702), .A2(new_n432), .ZN(new_n707));
  OAI21_X1  g506(.A(new_n707), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n708));
  XOR2_X1   g507(.A(KEYINPUT49), .B(G64gat), .Z(new_n709));
  OAI21_X1  g508(.A(new_n708), .B1(new_n707), .B2(new_n709), .ZN(G1333gat));
  INV_X1    g509(.A(G71gat), .ZN(new_n711));
  NAND3_X1  g510(.A1(new_n702), .A2(new_n711), .A3(new_n654), .ZN(new_n712));
  NAND2_X1  g511(.A1(new_n702), .A2(new_n684), .ZN(new_n713));
  INV_X1    g512(.A(new_n713), .ZN(new_n714));
  OAI21_X1  g513(.A(new_n712), .B1(new_n714), .B2(new_n711), .ZN(new_n715));
  XNOR2_X1  g514(.A(KEYINPUT110), .B(KEYINPUT50), .ZN(new_n716));
  XNOR2_X1  g515(.A(new_n715), .B(new_n716), .ZN(G1334gat));
  NAND2_X1  g516(.A1(new_n702), .A2(new_n634), .ZN(new_n718));
  XNOR2_X1  g517(.A(new_n718), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g518(.A1(new_n521), .A2(new_n599), .ZN(new_n720));
  OAI211_X1 g519(.A(new_n565), .B(new_n720), .C1(new_n437), .C2(new_n471), .ZN(new_n721));
  NAND2_X1  g520(.A1(new_n721), .A2(KEYINPUT51), .ZN(new_n722));
  INV_X1    g521(.A(KEYINPUT51), .ZN(new_n723));
  NAND4_X1  g522(.A1(new_n640), .A2(new_n723), .A3(new_n565), .A4(new_n720), .ZN(new_n724));
  AND2_X1   g523(.A1(new_n722), .A2(new_n724), .ZN(new_n725));
  NOR2_X1   g524(.A1(new_n623), .A2(G85gat), .ZN(new_n726));
  NAND3_X1  g525(.A1(new_n725), .A2(new_n626), .A3(new_n726), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n720), .A2(new_n622), .ZN(new_n728));
  XNOR2_X1  g527(.A(new_n728), .B(KEYINPUT111), .ZN(new_n729));
  NAND4_X1  g528(.A1(new_n668), .A2(new_n626), .A3(new_n669), .A4(new_n729), .ZN(new_n730));
  NAND2_X1  g529(.A1(new_n730), .A2(G85gat), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n727), .A2(new_n731), .ZN(new_n732));
  INV_X1    g531(.A(KEYINPUT112), .ZN(new_n733));
  XNOR2_X1  g532(.A(new_n732), .B(new_n733), .ZN(G1336gat));
  INV_X1    g533(.A(KEYINPUT114), .ZN(new_n735));
  NOR3_X1   g534(.A1(new_n431), .A2(new_n623), .A3(G92gat), .ZN(new_n736));
  NAND3_X1  g535(.A1(new_n722), .A2(new_n724), .A3(new_n736), .ZN(new_n737));
  INV_X1    g536(.A(KEYINPUT52), .ZN(new_n738));
  NAND2_X1  g537(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  NAND4_X1  g538(.A1(new_n668), .A2(new_n432), .A3(new_n669), .A4(new_n729), .ZN(new_n740));
  AOI21_X1  g539(.A(new_n739), .B1(new_n531), .B2(new_n740), .ZN(new_n741));
  NAND2_X1  g540(.A1(new_n740), .A2(new_n531), .ZN(new_n742));
  NAND2_X1  g541(.A1(new_n723), .A2(KEYINPUT113), .ZN(new_n743));
  INV_X1    g542(.A(new_n743), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n721), .A2(new_n744), .ZN(new_n745));
  NAND4_X1  g544(.A1(new_n640), .A2(new_n565), .A3(new_n720), .A4(new_n743), .ZN(new_n746));
  NAND2_X1  g545(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n747), .A2(new_n736), .ZN(new_n748));
  AOI21_X1  g547(.A(new_n738), .B1(new_n742), .B2(new_n748), .ZN(new_n749));
  OAI21_X1  g548(.A(new_n735), .B1(new_n741), .B2(new_n749), .ZN(new_n750));
  NAND3_X1  g549(.A1(new_n742), .A2(new_n738), .A3(new_n737), .ZN(new_n751));
  AOI22_X1  g550(.A1(new_n531), .A2(new_n740), .B1(new_n747), .B2(new_n736), .ZN(new_n752));
  OAI211_X1 g551(.A(new_n751), .B(KEYINPUT114), .C1(new_n738), .C2(new_n752), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n750), .A2(new_n753), .ZN(G1337gat));
  NAND4_X1  g553(.A1(new_n725), .A2(new_n528), .A3(new_n654), .A4(new_n622), .ZN(new_n755));
  NAND3_X1  g554(.A1(new_n668), .A2(new_n669), .A3(new_n729), .ZN(new_n756));
  OAI21_X1  g555(.A(G99gat), .B1(new_n756), .B2(new_n652), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n755), .A2(new_n757), .ZN(G1338gat));
  OAI21_X1  g557(.A(G106gat), .B1(new_n756), .B2(new_n423), .ZN(new_n759));
  INV_X1    g558(.A(new_n747), .ZN(new_n760));
  NOR3_X1   g559(.A1(new_n623), .A2(G106gat), .A3(new_n423), .ZN(new_n761));
  XNOR2_X1  g560(.A(new_n761), .B(KEYINPUT115), .ZN(new_n762));
  OAI21_X1  g561(.A(new_n759), .B1(new_n760), .B2(new_n762), .ZN(new_n763));
  NAND2_X1  g562(.A1(new_n763), .A2(KEYINPUT53), .ZN(new_n764));
  NAND3_X1  g563(.A1(new_n722), .A2(new_n724), .A3(new_n761), .ZN(new_n765));
  XNOR2_X1  g564(.A(new_n765), .B(KEYINPUT116), .ZN(new_n766));
  INV_X1    g565(.A(KEYINPUT53), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n759), .A2(new_n767), .ZN(new_n768));
  OAI21_X1  g567(.A(new_n764), .B1(new_n766), .B2(new_n768), .ZN(G1339gat));
  NOR2_X1   g568(.A1(new_n624), .A2(new_n521), .ZN(new_n770));
  INV_X1    g569(.A(KEYINPUT54), .ZN(new_n771));
  AOI21_X1  g570(.A(new_n771), .B1(new_n609), .B2(new_n610), .ZN(new_n772));
  OAI21_X1  g571(.A(new_n772), .B1(new_n610), .B2(new_n609), .ZN(new_n773));
  NAND3_X1  g572(.A1(new_n609), .A2(new_n771), .A3(new_n610), .ZN(new_n774));
  NAND4_X1  g573(.A1(new_n773), .A2(KEYINPUT55), .A3(new_n619), .A4(new_n774), .ZN(new_n775));
  AND2_X1   g574(.A1(new_n775), .A2(new_n621), .ZN(new_n776));
  NAND3_X1  g575(.A1(new_n773), .A2(new_n619), .A3(new_n774), .ZN(new_n777));
  INV_X1    g576(.A(KEYINPUT55), .ZN(new_n778));
  NAND2_X1  g577(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  NAND3_X1  g578(.A1(new_n776), .A2(new_n521), .A3(new_n779), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n496), .A2(new_n499), .ZN(new_n781));
  NAND3_X1  g580(.A1(new_n781), .A2(G229gat), .A3(G233gat), .ZN(new_n782));
  NOR2_X1   g581(.A1(new_n507), .A2(new_n508), .ZN(new_n783));
  INV_X1    g582(.A(new_n783), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n782), .A2(new_n784), .ZN(new_n785));
  AND2_X1   g584(.A1(new_n785), .A2(new_n515), .ZN(new_n786));
  AOI21_X1  g585(.A(new_n786), .B1(new_n506), .B2(new_n517), .ZN(new_n787));
  AOI21_X1  g586(.A(new_n565), .B1(new_n787), .B2(new_n622), .ZN(new_n788));
  AOI21_X1  g587(.A(new_n599), .B1(new_n780), .B2(new_n788), .ZN(new_n789));
  INV_X1    g588(.A(KEYINPUT117), .ZN(new_n790));
  OR2_X1    g589(.A1(new_n510), .A2(new_n516), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n503), .A2(new_n505), .ZN(new_n792));
  NOR2_X1   g591(.A1(new_n791), .A2(new_n792), .ZN(new_n793));
  OAI21_X1  g592(.A(new_n790), .B1(new_n793), .B2(new_n786), .ZN(new_n794));
  INV_X1    g593(.A(new_n786), .ZN(new_n795));
  NAND3_X1  g594(.A1(new_n518), .A2(KEYINPUT117), .A3(new_n795), .ZN(new_n796));
  NAND4_X1  g595(.A1(new_n794), .A2(new_n796), .A3(new_n776), .A4(new_n779), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n797), .A2(new_n565), .ZN(new_n798));
  AOI21_X1  g597(.A(new_n770), .B1(new_n789), .B2(new_n798), .ZN(new_n799));
  NOR2_X1   g598(.A1(new_n799), .A2(new_n703), .ZN(new_n800));
  AND2_X1   g599(.A1(new_n800), .A2(new_n638), .ZN(new_n801));
  AND2_X1   g600(.A1(new_n801), .A2(new_n431), .ZN(new_n802));
  AOI21_X1  g601(.A(G113gat), .B1(new_n802), .B2(new_n521), .ZN(new_n803));
  NAND2_X1  g602(.A1(new_n654), .A2(new_n423), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n626), .A2(new_n431), .ZN(new_n805));
  NOR3_X1   g604(.A1(new_n799), .A2(new_n804), .A3(new_n805), .ZN(new_n806));
  AND2_X1   g605(.A1(new_n521), .A2(G113gat), .ZN(new_n807));
  AOI21_X1  g606(.A(new_n803), .B1(new_n806), .B2(new_n807), .ZN(G1340gat));
  AOI21_X1  g607(.A(G120gat), .B1(new_n802), .B2(new_n622), .ZN(new_n809));
  AND2_X1   g608(.A1(new_n622), .A2(G120gat), .ZN(new_n810));
  AOI21_X1  g609(.A(new_n809), .B1(new_n806), .B2(new_n810), .ZN(G1341gat));
  NOR2_X1   g610(.A1(new_n598), .A2(G127gat), .ZN(new_n812));
  NAND2_X1  g611(.A1(new_n806), .A2(new_n599), .ZN(new_n813));
  AOI22_X1  g612(.A1(new_n802), .A2(new_n812), .B1(G127gat), .B2(new_n813), .ZN(new_n814));
  XNOR2_X1  g613(.A(new_n814), .B(KEYINPUT118), .ZN(G1342gat));
  NAND2_X1  g614(.A1(new_n565), .A2(new_n431), .ZN(new_n816));
  NOR2_X1   g615(.A1(new_n816), .A2(G134gat), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n801), .A2(new_n817), .ZN(new_n818));
  OR2_X1    g617(.A1(new_n818), .A2(KEYINPUT56), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n806), .A2(new_n565), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n820), .A2(G134gat), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n818), .A2(KEYINPUT56), .ZN(new_n822));
  NAND3_X1  g621(.A1(new_n819), .A2(new_n821), .A3(new_n822), .ZN(G1343gat));
  NAND2_X1  g622(.A1(new_n789), .A2(new_n798), .ZN(new_n824));
  INV_X1    g623(.A(new_n770), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n824), .A2(new_n825), .ZN(new_n826));
  NAND3_X1  g625(.A1(new_n826), .A2(KEYINPUT57), .A3(new_n634), .ZN(new_n827));
  INV_X1    g626(.A(KEYINPUT57), .ZN(new_n828));
  OAI21_X1  g627(.A(new_n828), .B1(new_n799), .B2(new_n423), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n827), .A2(new_n829), .ZN(new_n830));
  NOR2_X1   g629(.A1(new_n684), .A2(new_n805), .ZN(new_n831));
  NAND2_X1  g630(.A1(new_n830), .A2(new_n831), .ZN(new_n832));
  OAI21_X1  g631(.A(G141gat), .B1(new_n832), .B2(new_n522), .ZN(new_n833));
  NOR2_X1   g632(.A1(new_n684), .A2(new_n423), .ZN(new_n834));
  NAND2_X1  g633(.A1(new_n800), .A2(new_n834), .ZN(new_n835));
  INV_X1    g634(.A(new_n835), .ZN(new_n836));
  NAND2_X1  g635(.A1(new_n836), .A2(new_n431), .ZN(new_n837));
  OR2_X1    g636(.A1(new_n522), .A2(G141gat), .ZN(new_n838));
  OAI21_X1  g637(.A(new_n833), .B1(new_n837), .B2(new_n838), .ZN(new_n839));
  NAND2_X1  g638(.A1(new_n839), .A2(KEYINPUT58), .ZN(new_n840));
  INV_X1    g639(.A(KEYINPUT58), .ZN(new_n841));
  OAI211_X1 g640(.A(new_n833), .B(new_n841), .C1(new_n837), .C2(new_n838), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n840), .A2(new_n842), .ZN(G1344gat));
  NAND3_X1  g642(.A1(new_n830), .A2(new_n622), .A3(new_n831), .ZN(new_n844));
  INV_X1    g643(.A(KEYINPUT119), .ZN(new_n845));
  INV_X1    g644(.A(G148gat), .ZN(new_n846));
  NOR2_X1   g645(.A1(new_n846), .A2(KEYINPUT59), .ZN(new_n847));
  AND3_X1   g646(.A1(new_n844), .A2(new_n845), .A3(new_n847), .ZN(new_n848));
  AOI21_X1  g647(.A(new_n845), .B1(new_n844), .B2(new_n847), .ZN(new_n849));
  INV_X1    g648(.A(KEYINPUT121), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n827), .A2(new_n850), .ZN(new_n851));
  NOR3_X1   g650(.A1(new_n799), .A2(new_n828), .A3(new_n423), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n852), .A2(KEYINPUT121), .ZN(new_n853));
  NAND3_X1  g652(.A1(new_n851), .A2(new_n853), .A3(new_n829), .ZN(new_n854));
  NAND2_X1  g653(.A1(new_n831), .A2(new_n622), .ZN(new_n855));
  INV_X1    g654(.A(new_n855), .ZN(new_n856));
  AOI21_X1  g655(.A(new_n846), .B1(new_n854), .B2(new_n856), .ZN(new_n857));
  XNOR2_X1  g656(.A(KEYINPUT120), .B(KEYINPUT59), .ZN(new_n858));
  OAI22_X1  g657(.A1(new_n848), .A2(new_n849), .B1(new_n857), .B2(new_n858), .ZN(new_n859));
  NAND4_X1  g658(.A1(new_n836), .A2(new_n846), .A3(new_n431), .A4(new_n622), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n859), .A2(new_n860), .ZN(G1345gat));
  OAI21_X1  g660(.A(G155gat), .B1(new_n832), .B2(new_n598), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n599), .A2(new_n347), .ZN(new_n863));
  OAI21_X1  g662(.A(new_n862), .B1(new_n837), .B2(new_n863), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n864), .A2(KEYINPUT122), .ZN(new_n865));
  INV_X1    g664(.A(KEYINPUT122), .ZN(new_n866));
  OAI211_X1 g665(.A(new_n862), .B(new_n866), .C1(new_n837), .C2(new_n863), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n865), .A2(new_n867), .ZN(G1346gat));
  NOR3_X1   g667(.A1(new_n835), .A2(G162gat), .A3(new_n816), .ZN(new_n869));
  XOR2_X1   g668(.A(new_n869), .B(KEYINPUT123), .Z(new_n870));
  OAI21_X1  g669(.A(G162gat), .B1(new_n832), .B2(new_n566), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n870), .A2(new_n871), .ZN(G1347gat));
  NOR3_X1   g671(.A1(new_n799), .A2(new_n431), .A3(new_n626), .ZN(new_n873));
  NAND2_X1  g672(.A1(new_n873), .A2(new_n638), .ZN(new_n874));
  INV_X1    g673(.A(new_n874), .ZN(new_n875));
  AOI21_X1  g674(.A(G169gat), .B1(new_n875), .B2(new_n521), .ZN(new_n876));
  NAND2_X1  g675(.A1(new_n703), .A2(new_n432), .ZN(new_n877));
  NOR3_X1   g676(.A1(new_n799), .A2(new_n804), .A3(new_n877), .ZN(new_n878));
  NOR2_X1   g677(.A1(new_n522), .A2(new_n219), .ZN(new_n879));
  AOI21_X1  g678(.A(new_n876), .B1(new_n878), .B2(new_n879), .ZN(G1348gat));
  INV_X1    g679(.A(new_n877), .ZN(new_n881));
  NAND4_X1  g680(.A1(new_n826), .A2(new_n423), .A3(new_n654), .A4(new_n881), .ZN(new_n882));
  OAI21_X1  g681(.A(G176gat), .B1(new_n882), .B2(new_n623), .ZN(new_n883));
  NAND2_X1  g682(.A1(new_n622), .A2(new_n220), .ZN(new_n884));
  OAI21_X1  g683(.A(new_n883), .B1(new_n874), .B2(new_n884), .ZN(G1349gat));
  NAND2_X1  g684(.A1(new_n205), .A2(KEYINPUT27), .ZN(new_n886));
  NAND3_X1  g685(.A1(new_n599), .A2(new_n886), .A3(new_n245), .ZN(new_n887));
  INV_X1    g686(.A(new_n887), .ZN(new_n888));
  AND3_X1   g687(.A1(new_n873), .A2(new_n638), .A3(new_n888), .ZN(new_n889));
  AOI21_X1  g688(.A(new_n205), .B1(new_n878), .B2(new_n599), .ZN(new_n890));
  OAI21_X1  g689(.A(KEYINPUT125), .B1(new_n889), .B2(new_n890), .ZN(new_n891));
  OAI21_X1  g690(.A(G183gat), .B1(new_n882), .B2(new_n598), .ZN(new_n892));
  INV_X1    g691(.A(KEYINPUT125), .ZN(new_n893));
  NAND3_X1  g692(.A1(new_n873), .A2(new_n638), .A3(new_n888), .ZN(new_n894));
  NAND3_X1  g693(.A1(new_n892), .A2(new_n893), .A3(new_n894), .ZN(new_n895));
  NAND2_X1  g694(.A1(new_n891), .A2(new_n895), .ZN(new_n896));
  AND2_X1   g695(.A1(KEYINPUT124), .A2(KEYINPUT60), .ZN(new_n897));
  XNOR2_X1  g696(.A(new_n896), .B(new_n897), .ZN(G1350gat));
  NOR2_X1   g697(.A1(new_n566), .A2(G190gat), .ZN(new_n899));
  INV_X1    g698(.A(new_n899), .ZN(new_n900));
  OAI21_X1  g699(.A(KEYINPUT126), .B1(new_n874), .B2(new_n900), .ZN(new_n901));
  INV_X1    g700(.A(KEYINPUT126), .ZN(new_n902));
  NAND4_X1  g701(.A1(new_n873), .A2(new_n902), .A3(new_n638), .A4(new_n899), .ZN(new_n903));
  NAND2_X1  g702(.A1(new_n901), .A2(new_n903), .ZN(new_n904));
  AOI21_X1  g703(.A(new_n206), .B1(new_n878), .B2(new_n565), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n905), .A2(KEYINPUT61), .ZN(new_n906));
  OR2_X1    g705(.A1(new_n905), .A2(KEYINPUT61), .ZN(new_n907));
  NAND3_X1  g706(.A1(new_n904), .A2(new_n906), .A3(new_n907), .ZN(new_n908));
  INV_X1    g707(.A(KEYINPUT127), .ZN(new_n909));
  NAND2_X1  g708(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  NAND4_X1  g709(.A1(new_n904), .A2(new_n907), .A3(KEYINPUT127), .A4(new_n906), .ZN(new_n911));
  NAND2_X1  g710(.A1(new_n910), .A2(new_n911), .ZN(G1351gat));
  NAND2_X1  g711(.A1(new_n873), .A2(new_n834), .ZN(new_n913));
  INV_X1    g712(.A(new_n913), .ZN(new_n914));
  AOI21_X1  g713(.A(G197gat), .B1(new_n914), .B2(new_n521), .ZN(new_n915));
  NOR2_X1   g714(.A1(new_n684), .A2(new_n877), .ZN(new_n916));
  AND2_X1   g715(.A1(new_n854), .A2(new_n916), .ZN(new_n917));
  AND2_X1   g716(.A1(new_n521), .A2(G197gat), .ZN(new_n918));
  AOI21_X1  g717(.A(new_n915), .B1(new_n917), .B2(new_n918), .ZN(G1352gat));
  NOR3_X1   g718(.A1(new_n913), .A2(G204gat), .A3(new_n623), .ZN(new_n920));
  XNOR2_X1  g719(.A(new_n920), .B(KEYINPUT62), .ZN(new_n921));
  NAND3_X1  g720(.A1(new_n854), .A2(new_n622), .A3(new_n916), .ZN(new_n922));
  NAND2_X1  g721(.A1(new_n922), .A2(G204gat), .ZN(new_n923));
  NAND2_X1  g722(.A1(new_n921), .A2(new_n923), .ZN(G1353gat));
  NAND3_X1  g723(.A1(new_n914), .A2(new_n306), .A3(new_n599), .ZN(new_n925));
  OAI21_X1  g724(.A(new_n829), .B1(new_n852), .B2(KEYINPUT121), .ZN(new_n926));
  NOR2_X1   g725(.A1(new_n827), .A2(new_n850), .ZN(new_n927));
  OAI211_X1 g726(.A(new_n599), .B(new_n916), .C1(new_n926), .C2(new_n927), .ZN(new_n928));
  AND3_X1   g727(.A1(new_n928), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n929));
  AOI21_X1  g728(.A(KEYINPUT63), .B1(new_n928), .B2(G211gat), .ZN(new_n930));
  OAI21_X1  g729(.A(new_n925), .B1(new_n929), .B2(new_n930), .ZN(G1354gat));
  NAND3_X1  g730(.A1(new_n854), .A2(new_n565), .A3(new_n916), .ZN(new_n932));
  NAND2_X1  g731(.A1(new_n932), .A2(G218gat), .ZN(new_n933));
  NAND3_X1  g732(.A1(new_n914), .A2(new_n307), .A3(new_n565), .ZN(new_n934));
  NAND2_X1  g733(.A1(new_n933), .A2(new_n934), .ZN(G1355gat));
endmodule


