//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 1 0 1 0 1 1 1 1 0 0 0 1 1 0 0 1 0 1 1 0 1 0 1 1 0 0 1 1 0 1 1 0 0 1 1 1 1 1 0 0 0 0 1 1 0 1 1 0 1 0 1 0 0 1 1 1 0 0 0 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:16:52 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n683, new_n684, new_n685,
    new_n686, new_n687, new_n689, new_n690, new_n691, new_n693, new_n694,
    new_n695, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n719, new_n720, new_n721, new_n722, new_n723, new_n724,
    new_n725, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n753, new_n754, new_n755, new_n756,
    new_n757, new_n759, new_n760, new_n761, new_n762, new_n764, new_n765,
    new_n767, new_n768, new_n769, new_n770, new_n771, new_n772, new_n773,
    new_n774, new_n775, new_n776, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n787, new_n788, new_n789,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n862, new_n863,
    new_n864, new_n866, new_n867, new_n868, new_n869, new_n870, new_n871,
    new_n872, new_n873, new_n874, new_n875, new_n876, new_n877, new_n878,
    new_n879, new_n880, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n930,
    new_n931, new_n932, new_n933, new_n935, new_n936, new_n937, new_n938,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n951, new_n952, new_n953, new_n955,
    new_n956, new_n957, new_n958, new_n959, new_n960, new_n961, new_n963,
    new_n964, new_n965, new_n966, new_n967, new_n968, new_n969, new_n970,
    new_n971, new_n972, new_n973, new_n975, new_n976, new_n977, new_n978,
    new_n979, new_n980, new_n981, new_n982, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n990, new_n991, new_n992, new_n993, new_n994,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001;
  NAND2_X1  g000(.A1(G225gat), .A2(G233gat), .ZN(new_n202));
  INV_X1    g001(.A(KEYINPUT76), .ZN(new_n203));
  AND2_X1   g002(.A1(G155gat), .A2(G162gat), .ZN(new_n204));
  NOR2_X1   g003(.A1(G155gat), .A2(G162gat), .ZN(new_n205));
  OAI21_X1  g004(.A(new_n203), .B1(new_n204), .B2(new_n205), .ZN(new_n206));
  INV_X1    g005(.A(G141gat), .ZN(new_n207));
  INV_X1    g006(.A(G148gat), .ZN(new_n208));
  NAND2_X1  g007(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  INV_X1    g008(.A(KEYINPUT2), .ZN(new_n210));
  NAND2_X1  g009(.A1(G141gat), .A2(G148gat), .ZN(new_n211));
  NAND3_X1  g010(.A1(new_n209), .A2(new_n210), .A3(new_n211), .ZN(new_n212));
  OAI21_X1  g011(.A(KEYINPUT76), .B1(G155gat), .B2(G162gat), .ZN(new_n213));
  NAND3_X1  g012(.A1(new_n206), .A2(new_n212), .A3(new_n213), .ZN(new_n214));
  XNOR2_X1  g013(.A(KEYINPUT77), .B(G162gat), .ZN(new_n215));
  AOI21_X1  g014(.A(new_n210), .B1(new_n215), .B2(G155gat), .ZN(new_n216));
  XNOR2_X1  g015(.A(G155gat), .B(G162gat), .ZN(new_n217));
  NAND3_X1  g016(.A1(new_n217), .A2(new_n209), .A3(new_n211), .ZN(new_n218));
  OAI21_X1  g017(.A(new_n214), .B1(new_n216), .B2(new_n218), .ZN(new_n219));
  XOR2_X1   g018(.A(G127gat), .B(G134gat), .Z(new_n220));
  XNOR2_X1  g019(.A(G113gat), .B(G120gat), .ZN(new_n221));
  INV_X1    g020(.A(KEYINPUT1), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n222), .A2(KEYINPUT68), .ZN(new_n223));
  OAI21_X1  g022(.A(new_n220), .B1(new_n221), .B2(new_n223), .ZN(new_n224));
  INV_X1    g023(.A(G120gat), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n225), .A2(G113gat), .ZN(new_n226));
  INV_X1    g025(.A(G113gat), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n227), .A2(G120gat), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n226), .A2(new_n228), .ZN(new_n229));
  XNOR2_X1  g028(.A(G127gat), .B(G134gat), .ZN(new_n230));
  NAND4_X1  g029(.A1(new_n229), .A2(new_n230), .A3(KEYINPUT68), .A4(new_n222), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n224), .A2(new_n231), .ZN(new_n232));
  INV_X1    g031(.A(KEYINPUT4), .ZN(new_n233));
  NOR3_X1   g032(.A1(new_n219), .A2(new_n232), .A3(new_n233), .ZN(new_n234));
  INV_X1    g033(.A(KEYINPUT69), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n232), .A2(new_n235), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n215), .A2(G155gat), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n237), .A2(KEYINPUT2), .ZN(new_n238));
  AND3_X1   g037(.A1(new_n217), .A2(new_n209), .A3(new_n211), .ZN(new_n239));
  INV_X1    g038(.A(new_n213), .ZN(new_n240));
  AOI21_X1  g039(.A(new_n240), .B1(new_n217), .B2(new_n203), .ZN(new_n241));
  AOI22_X1  g040(.A1(new_n238), .A2(new_n239), .B1(new_n241), .B2(new_n212), .ZN(new_n242));
  NAND3_X1  g041(.A1(new_n224), .A2(new_n231), .A3(KEYINPUT69), .ZN(new_n243));
  NAND3_X1  g042(.A1(new_n236), .A2(new_n242), .A3(new_n243), .ZN(new_n244));
  AOI21_X1  g043(.A(new_n234), .B1(new_n244), .B2(new_n233), .ZN(new_n245));
  INV_X1    g044(.A(KEYINPUT78), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n219), .A2(new_n246), .ZN(new_n247));
  OAI211_X1 g046(.A(new_n214), .B(KEYINPUT78), .C1(new_n216), .C2(new_n218), .ZN(new_n248));
  NAND3_X1  g047(.A1(new_n247), .A2(KEYINPUT3), .A3(new_n248), .ZN(new_n249));
  INV_X1    g048(.A(KEYINPUT3), .ZN(new_n250));
  OAI211_X1 g049(.A(new_n214), .B(new_n250), .C1(new_n216), .C2(new_n218), .ZN(new_n251));
  AND2_X1   g050(.A1(new_n251), .A2(new_n232), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n249), .A2(new_n252), .ZN(new_n253));
  AOI21_X1  g052(.A(new_n202), .B1(new_n245), .B2(new_n253), .ZN(new_n254));
  NAND3_X1  g053(.A1(new_n247), .A2(new_n248), .A3(new_n232), .ZN(new_n255));
  NOR2_X1   g054(.A1(new_n219), .A2(new_n232), .ZN(new_n256));
  INV_X1    g055(.A(new_n256), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n255), .A2(new_n257), .ZN(new_n258));
  INV_X1    g057(.A(new_n202), .ZN(new_n259));
  OAI21_X1  g058(.A(KEYINPUT39), .B1(new_n258), .B2(new_n259), .ZN(new_n260));
  OR2_X1    g059(.A1(new_n254), .A2(new_n260), .ZN(new_n261));
  XOR2_X1   g060(.A(G1gat), .B(G29gat), .Z(new_n262));
  XNOR2_X1  g061(.A(G57gat), .B(G85gat), .ZN(new_n263));
  XNOR2_X1  g062(.A(new_n262), .B(new_n263), .ZN(new_n264));
  XNOR2_X1  g063(.A(KEYINPUT79), .B(KEYINPUT0), .ZN(new_n265));
  XNOR2_X1  g064(.A(new_n264), .B(new_n265), .ZN(new_n266));
  XNOR2_X1  g065(.A(KEYINPUT85), .B(KEYINPUT39), .ZN(new_n267));
  AOI21_X1  g066(.A(new_n266), .B1(new_n254), .B2(new_n267), .ZN(new_n268));
  INV_X1    g067(.A(KEYINPUT40), .ZN(new_n269));
  AND3_X1   g068(.A1(new_n261), .A2(new_n268), .A3(new_n269), .ZN(new_n270));
  AOI21_X1  g069(.A(new_n269), .B1(new_n261), .B2(new_n268), .ZN(new_n271));
  NOR2_X1   g070(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  INV_X1    g071(.A(KEYINPUT86), .ZN(new_n273));
  AOI21_X1  g072(.A(new_n259), .B1(new_n249), .B2(new_n252), .ZN(new_n274));
  INV_X1    g073(.A(KEYINPUT5), .ZN(new_n275));
  AND2_X1   g074(.A1(new_n245), .A2(new_n275), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n256), .A2(new_n233), .ZN(new_n277));
  AND3_X1   g076(.A1(new_n236), .A2(new_n242), .A3(new_n243), .ZN(new_n278));
  OAI21_X1  g077(.A(new_n277), .B1(new_n278), .B2(new_n233), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n279), .A2(new_n274), .ZN(new_n280));
  AOI21_X1  g079(.A(new_n275), .B1(new_n258), .B2(new_n259), .ZN(new_n281));
  AOI22_X1  g080(.A1(new_n274), .A2(new_n276), .B1(new_n280), .B2(new_n281), .ZN(new_n282));
  INV_X1    g081(.A(new_n266), .ZN(new_n283));
  OAI21_X1  g082(.A(new_n273), .B1(new_n282), .B2(new_n283), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n276), .A2(new_n274), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n280), .A2(new_n281), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  NAND3_X1  g086(.A1(new_n287), .A2(KEYINPUT86), .A3(new_n266), .ZN(new_n288));
  NAND2_X1  g087(.A1(new_n284), .A2(new_n288), .ZN(new_n289));
  NOR2_X1   g088(.A1(new_n272), .A2(new_n289), .ZN(new_n290));
  AND2_X1   g089(.A1(G211gat), .A2(G218gat), .ZN(new_n291));
  NOR2_X1   g090(.A1(G211gat), .A2(G218gat), .ZN(new_n292));
  NOR2_X1   g091(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  AND2_X1   g092(.A1(G197gat), .A2(G204gat), .ZN(new_n294));
  NOR2_X1   g093(.A1(G197gat), .A2(G204gat), .ZN(new_n295));
  NOR2_X1   g094(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  AOI21_X1  g095(.A(KEYINPUT22), .B1(G211gat), .B2(G218gat), .ZN(new_n297));
  OAI21_X1  g096(.A(new_n293), .B1(new_n296), .B2(new_n297), .ZN(new_n298));
  XNOR2_X1  g097(.A(G211gat), .B(G218gat), .ZN(new_n299));
  XNOR2_X1  g098(.A(G197gat), .B(G204gat), .ZN(new_n300));
  INV_X1    g099(.A(new_n297), .ZN(new_n301));
  NAND3_X1  g100(.A1(new_n299), .A2(new_n300), .A3(new_n301), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n298), .A2(new_n302), .ZN(new_n303));
  INV_X1    g102(.A(new_n303), .ZN(new_n304));
  NAND2_X1  g103(.A1(G226gat), .A2(G233gat), .ZN(new_n305));
  INV_X1    g104(.A(new_n305), .ZN(new_n306));
  INV_X1    g105(.A(G169gat), .ZN(new_n307));
  INV_X1    g106(.A(G176gat), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  INV_X1    g108(.A(KEYINPUT26), .ZN(new_n310));
  NOR2_X1   g109(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  AOI21_X1  g110(.A(new_n311), .B1(G183gat), .B2(G190gat), .ZN(new_n312));
  NAND2_X1  g111(.A1(G169gat), .A2(G176gat), .ZN(new_n313));
  NAND3_X1  g112(.A1(new_n309), .A2(new_n310), .A3(new_n313), .ZN(new_n314));
  AND2_X1   g113(.A1(KEYINPUT66), .A2(G190gat), .ZN(new_n315));
  NOR2_X1   g114(.A1(KEYINPUT66), .A2(G190gat), .ZN(new_n316));
  NOR2_X1   g115(.A1(new_n315), .A2(new_n316), .ZN(new_n317));
  XNOR2_X1  g116(.A(KEYINPUT27), .B(G183gat), .ZN(new_n318));
  AND3_X1   g117(.A1(new_n317), .A2(new_n318), .A3(KEYINPUT28), .ZN(new_n319));
  AOI21_X1  g118(.A(KEYINPUT28), .B1(new_n317), .B2(new_n318), .ZN(new_n320));
  OAI211_X1 g119(.A(new_n312), .B(new_n314), .C1(new_n319), .C2(new_n320), .ZN(new_n321));
  INV_X1    g120(.A(KEYINPUT65), .ZN(new_n322));
  INV_X1    g121(.A(KEYINPUT25), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n308), .A2(KEYINPUT64), .ZN(new_n324));
  INV_X1    g123(.A(KEYINPUT64), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n325), .A2(G176gat), .ZN(new_n326));
  NAND4_X1  g125(.A1(new_n324), .A2(new_n326), .A3(KEYINPUT23), .A4(new_n307), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n313), .A2(KEYINPUT23), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n328), .A2(new_n309), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n327), .A2(new_n329), .ZN(new_n330));
  NOR2_X1   g129(.A1(G183gat), .A2(G190gat), .ZN(new_n331));
  INV_X1    g130(.A(G183gat), .ZN(new_n332));
  INV_X1    g131(.A(G190gat), .ZN(new_n333));
  OAI21_X1  g132(.A(KEYINPUT24), .B1(new_n332), .B2(new_n333), .ZN(new_n334));
  INV_X1    g133(.A(KEYINPUT24), .ZN(new_n335));
  NAND3_X1  g134(.A1(new_n335), .A2(G183gat), .A3(G190gat), .ZN(new_n336));
  AOI21_X1  g135(.A(new_n331), .B1(new_n334), .B2(new_n336), .ZN(new_n337));
  OAI211_X1 g136(.A(new_n322), .B(new_n323), .C1(new_n330), .C2(new_n337), .ZN(new_n338));
  AOI22_X1  g137(.A1(new_n317), .A2(new_n332), .B1(new_n334), .B2(new_n336), .ZN(new_n339));
  NAND3_X1  g138(.A1(new_n307), .A2(new_n308), .A3(KEYINPUT23), .ZN(new_n340));
  NAND3_X1  g139(.A1(new_n329), .A2(KEYINPUT25), .A3(new_n340), .ZN(new_n341));
  OAI21_X1  g140(.A(KEYINPUT67), .B1(new_n339), .B2(new_n341), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n334), .A2(new_n336), .ZN(new_n343));
  INV_X1    g142(.A(new_n316), .ZN(new_n344));
  NAND2_X1  g143(.A1(KEYINPUT66), .A2(G190gat), .ZN(new_n345));
  NAND3_X1  g144(.A1(new_n344), .A2(new_n332), .A3(new_n345), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n343), .A2(new_n346), .ZN(new_n347));
  INV_X1    g146(.A(KEYINPUT67), .ZN(new_n348));
  AND2_X1   g147(.A1(new_n340), .A2(KEYINPUT25), .ZN(new_n349));
  NAND4_X1  g148(.A1(new_n347), .A2(new_n348), .A3(new_n329), .A4(new_n349), .ZN(new_n350));
  NAND3_X1  g149(.A1(new_n338), .A2(new_n342), .A3(new_n350), .ZN(new_n351));
  AND2_X1   g150(.A1(new_n334), .A2(new_n336), .ZN(new_n352));
  OAI211_X1 g151(.A(new_n327), .B(new_n329), .C1(new_n352), .C2(new_n331), .ZN(new_n353));
  AOI21_X1  g152(.A(new_n322), .B1(new_n353), .B2(new_n323), .ZN(new_n354));
  OAI21_X1  g153(.A(new_n321), .B1(new_n351), .B2(new_n354), .ZN(new_n355));
  INV_X1    g154(.A(KEYINPUT29), .ZN(new_n356));
  AOI21_X1  g155(.A(new_n306), .B1(new_n355), .B2(new_n356), .ZN(new_n357));
  OAI21_X1  g156(.A(new_n323), .B1(new_n330), .B2(new_n337), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n358), .A2(KEYINPUT65), .ZN(new_n359));
  NAND4_X1  g158(.A1(new_n359), .A2(new_n338), .A3(new_n342), .A4(new_n350), .ZN(new_n360));
  AOI21_X1  g159(.A(new_n305), .B1(new_n360), .B2(new_n321), .ZN(new_n361));
  OAI21_X1  g160(.A(new_n304), .B1(new_n357), .B2(new_n361), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n355), .A2(new_n306), .ZN(new_n363));
  AOI21_X1  g162(.A(KEYINPUT29), .B1(new_n360), .B2(new_n321), .ZN(new_n364));
  OAI211_X1 g163(.A(new_n363), .B(new_n303), .C1(new_n364), .C2(new_n306), .ZN(new_n365));
  AND2_X1   g164(.A1(new_n362), .A2(new_n365), .ZN(new_n366));
  INV_X1    g165(.A(KEYINPUT74), .ZN(new_n367));
  XOR2_X1   g166(.A(G8gat), .B(G36gat), .Z(new_n368));
  XOR2_X1   g167(.A(G64gat), .B(G92gat), .Z(new_n369));
  XOR2_X1   g168(.A(new_n368), .B(new_n369), .Z(new_n370));
  NAND4_X1  g169(.A1(new_n366), .A2(new_n367), .A3(KEYINPUT30), .A4(new_n370), .ZN(new_n371));
  NAND4_X1  g170(.A1(new_n362), .A2(KEYINPUT30), .A3(new_n365), .A4(new_n370), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n372), .A2(KEYINPUT74), .ZN(new_n373));
  INV_X1    g172(.A(KEYINPUT73), .ZN(new_n374));
  NAND2_X1  g173(.A1(new_n362), .A2(new_n365), .ZN(new_n375));
  XOR2_X1   g174(.A(new_n370), .B(KEYINPUT72), .Z(new_n376));
  AOI21_X1  g175(.A(new_n374), .B1(new_n375), .B2(new_n376), .ZN(new_n377));
  INV_X1    g176(.A(new_n376), .ZN(new_n378));
  AOI211_X1 g177(.A(KEYINPUT73), .B(new_n378), .C1(new_n362), .C2(new_n365), .ZN(new_n379));
  OAI211_X1 g178(.A(new_n371), .B(new_n373), .C1(new_n377), .C2(new_n379), .ZN(new_n380));
  INV_X1    g179(.A(new_n370), .ZN(new_n381));
  NOR2_X1   g180(.A1(new_n375), .A2(new_n381), .ZN(new_n382));
  NOR2_X1   g181(.A1(new_n382), .A2(KEYINPUT30), .ZN(new_n383));
  OAI21_X1  g182(.A(new_n290), .B1(new_n380), .B2(new_n383), .ZN(new_n384));
  XNOR2_X1  g183(.A(KEYINPUT81), .B(KEYINPUT31), .ZN(new_n385));
  INV_X1    g184(.A(new_n385), .ZN(new_n386));
  AOI21_X1  g185(.A(KEYINPUT29), .B1(new_n298), .B2(new_n302), .ZN(new_n387));
  OAI211_X1 g186(.A(new_n247), .B(new_n248), .C1(KEYINPUT3), .C2(new_n387), .ZN(new_n388));
  INV_X1    g187(.A(G228gat), .ZN(new_n389));
  INV_X1    g188(.A(G233gat), .ZN(new_n390));
  NOR2_X1   g189(.A1(new_n389), .A2(new_n390), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n251), .A2(new_n356), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n392), .A2(new_n304), .ZN(new_n393));
  NAND3_X1  g192(.A1(new_n388), .A2(new_n391), .A3(new_n393), .ZN(new_n394));
  INV_X1    g193(.A(KEYINPUT83), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n393), .A2(new_n395), .ZN(new_n396));
  NAND3_X1  g195(.A1(new_n392), .A2(KEYINPUT83), .A3(new_n304), .ZN(new_n397));
  INV_X1    g196(.A(KEYINPUT82), .ZN(new_n398));
  OAI21_X1  g197(.A(new_n250), .B1(new_n387), .B2(new_n398), .ZN(new_n399));
  AOI211_X1 g198(.A(KEYINPUT82), .B(KEYINPUT29), .C1(new_n298), .C2(new_n302), .ZN(new_n400));
  OAI21_X1  g199(.A(new_n219), .B1(new_n399), .B2(new_n400), .ZN(new_n401));
  NAND3_X1  g200(.A1(new_n396), .A2(new_n397), .A3(new_n401), .ZN(new_n402));
  INV_X1    g201(.A(KEYINPUT84), .ZN(new_n403));
  INV_X1    g202(.A(new_n391), .ZN(new_n404));
  AND3_X1   g203(.A1(new_n402), .A2(new_n403), .A3(new_n404), .ZN(new_n405));
  AOI21_X1  g204(.A(new_n403), .B1(new_n402), .B2(new_n404), .ZN(new_n406));
  OAI21_X1  g205(.A(new_n394), .B1(new_n405), .B2(new_n406), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n407), .A2(G22gat), .ZN(new_n408));
  XNOR2_X1  g207(.A(G78gat), .B(G106gat), .ZN(new_n409));
  INV_X1    g208(.A(G50gat), .ZN(new_n410));
  XNOR2_X1  g209(.A(new_n409), .B(new_n410), .ZN(new_n411));
  INV_X1    g210(.A(new_n411), .ZN(new_n412));
  INV_X1    g211(.A(G22gat), .ZN(new_n413));
  OAI211_X1 g212(.A(new_n413), .B(new_n394), .C1(new_n405), .C2(new_n406), .ZN(new_n414));
  AND3_X1   g213(.A1(new_n408), .A2(new_n412), .A3(new_n414), .ZN(new_n415));
  AOI21_X1  g214(.A(new_n412), .B1(new_n408), .B2(new_n414), .ZN(new_n416));
  OAI21_X1  g215(.A(new_n386), .B1(new_n415), .B2(new_n416), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n402), .A2(new_n404), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n418), .A2(KEYINPUT84), .ZN(new_n419));
  NAND3_X1  g218(.A1(new_n402), .A2(new_n403), .A3(new_n404), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  AOI21_X1  g220(.A(new_n413), .B1(new_n421), .B2(new_n394), .ZN(new_n422));
  INV_X1    g221(.A(new_n414), .ZN(new_n423));
  OAI21_X1  g222(.A(new_n411), .B1(new_n422), .B2(new_n423), .ZN(new_n424));
  NAND3_X1  g223(.A1(new_n408), .A2(new_n412), .A3(new_n414), .ZN(new_n425));
  NAND3_X1  g224(.A1(new_n424), .A2(new_n385), .A3(new_n425), .ZN(new_n426));
  INV_X1    g225(.A(KEYINPUT37), .ZN(new_n427));
  NAND3_X1  g226(.A1(new_n362), .A2(new_n427), .A3(new_n365), .ZN(new_n428));
  NOR2_X1   g227(.A1(new_n378), .A2(KEYINPUT38), .ZN(new_n429));
  AND2_X1   g228(.A1(new_n428), .A2(new_n429), .ZN(new_n430));
  AOI21_X1  g229(.A(new_n427), .B1(new_n362), .B2(new_n365), .ZN(new_n431));
  INV_X1    g230(.A(new_n431), .ZN(new_n432));
  AOI21_X1  g231(.A(new_n382), .B1(new_n430), .B2(new_n432), .ZN(new_n433));
  XNOR2_X1  g232(.A(KEYINPUT80), .B(KEYINPUT6), .ZN(new_n434));
  INV_X1    g233(.A(new_n434), .ZN(new_n435));
  NAND3_X1  g234(.A1(new_n287), .A2(new_n266), .A3(new_n435), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n428), .A2(new_n381), .ZN(new_n437));
  OAI21_X1  g236(.A(KEYINPUT38), .B1(new_n437), .B2(new_n431), .ZN(new_n438));
  AOI21_X1  g237(.A(new_n435), .B1(new_n282), .B2(new_n283), .ZN(new_n439));
  NAND3_X1  g238(.A1(new_n284), .A2(new_n439), .A3(new_n288), .ZN(new_n440));
  NAND4_X1  g239(.A1(new_n433), .A2(new_n436), .A3(new_n438), .A4(new_n440), .ZN(new_n441));
  NAND4_X1  g240(.A1(new_n384), .A2(new_n417), .A3(new_n426), .A4(new_n441), .ZN(new_n442));
  INV_X1    g241(.A(KEYINPUT36), .ZN(new_n443));
  INV_X1    g242(.A(G227gat), .ZN(new_n444));
  NOR2_X1   g243(.A1(new_n444), .A2(new_n390), .ZN(new_n445));
  INV_X1    g244(.A(new_n445), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n236), .A2(new_n243), .ZN(new_n447));
  OAI211_X1 g246(.A(new_n447), .B(new_n321), .C1(new_n351), .C2(new_n354), .ZN(new_n448));
  INV_X1    g247(.A(new_n448), .ZN(new_n449));
  AOI21_X1  g248(.A(new_n447), .B1(new_n360), .B2(new_n321), .ZN(new_n450));
  OAI21_X1  g249(.A(new_n446), .B1(new_n449), .B2(new_n450), .ZN(new_n451));
  INV_X1    g250(.A(KEYINPUT71), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n451), .A2(new_n452), .ZN(new_n453));
  INV_X1    g252(.A(new_n447), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n355), .A2(new_n454), .ZN(new_n455));
  AOI21_X1  g254(.A(new_n445), .B1(new_n455), .B2(new_n448), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n456), .A2(KEYINPUT71), .ZN(new_n457));
  INV_X1    g256(.A(KEYINPUT34), .ZN(new_n458));
  NAND3_X1  g257(.A1(new_n453), .A2(new_n457), .A3(new_n458), .ZN(new_n459));
  NAND3_X1  g258(.A1(new_n456), .A2(KEYINPUT71), .A3(KEYINPUT34), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  XNOR2_X1  g260(.A(G15gat), .B(G43gat), .ZN(new_n462));
  XNOR2_X1  g261(.A(G71gat), .B(G99gat), .ZN(new_n463));
  XNOR2_X1  g262(.A(new_n462), .B(new_n463), .ZN(new_n464));
  NAND3_X1  g263(.A1(new_n455), .A2(new_n445), .A3(new_n448), .ZN(new_n465));
  INV_X1    g264(.A(KEYINPUT33), .ZN(new_n466));
  AOI21_X1  g265(.A(new_n464), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  AOI22_X1  g266(.A1(new_n467), .A2(KEYINPUT70), .B1(KEYINPUT32), .B2(new_n465), .ZN(new_n468));
  NOR2_X1   g267(.A1(new_n464), .A2(new_n466), .ZN(new_n469));
  NAND3_X1  g268(.A1(new_n465), .A2(KEYINPUT32), .A3(new_n469), .ZN(new_n470));
  INV_X1    g269(.A(KEYINPUT70), .ZN(new_n471));
  AOI21_X1  g270(.A(new_n470), .B1(new_n467), .B2(new_n471), .ZN(new_n472));
  NOR3_X1   g271(.A1(new_n461), .A2(new_n468), .A3(new_n472), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n467), .A2(KEYINPUT70), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n465), .A2(KEYINPUT32), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n465), .A2(new_n466), .ZN(new_n477));
  INV_X1    g276(.A(new_n464), .ZN(new_n478));
  NAND3_X1  g277(.A1(new_n477), .A2(new_n471), .A3(new_n478), .ZN(new_n479));
  INV_X1    g278(.A(new_n470), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  AOI22_X1  g280(.A1(new_n476), .A2(new_n481), .B1(new_n460), .B2(new_n459), .ZN(new_n482));
  OAI21_X1  g281(.A(new_n443), .B1(new_n473), .B2(new_n482), .ZN(new_n483));
  OAI21_X1  g282(.A(new_n461), .B1(new_n468), .B2(new_n472), .ZN(new_n484));
  NAND4_X1  g283(.A1(new_n476), .A2(new_n481), .A3(new_n460), .A4(new_n459), .ZN(new_n485));
  NAND3_X1  g284(.A1(new_n484), .A2(new_n485), .A3(KEYINPUT36), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n483), .A2(new_n486), .ZN(new_n487));
  AND2_X1   g286(.A1(new_n442), .A2(new_n487), .ZN(new_n488));
  INV_X1    g287(.A(KEYINPUT75), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n371), .A2(new_n373), .ZN(new_n490));
  NOR2_X1   g289(.A1(new_n377), .A2(new_n379), .ZN(new_n491));
  OAI21_X1  g290(.A(new_n489), .B1(new_n490), .B2(new_n491), .ZN(new_n492));
  XNOR2_X1  g291(.A(new_n372), .B(new_n367), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n375), .A2(new_n376), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n494), .A2(KEYINPUT73), .ZN(new_n495));
  NAND3_X1  g294(.A1(new_n375), .A2(new_n374), .A3(new_n376), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  NAND3_X1  g296(.A1(new_n493), .A2(new_n497), .A3(KEYINPUT75), .ZN(new_n498));
  OAI21_X1  g297(.A(new_n439), .B1(new_n283), .B2(new_n282), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n499), .A2(new_n436), .ZN(new_n500));
  INV_X1    g299(.A(new_n383), .ZN(new_n501));
  NAND4_X1  g300(.A1(new_n492), .A2(new_n498), .A3(new_n500), .A4(new_n501), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n417), .A2(new_n426), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  NOR2_X1   g303(.A1(new_n473), .A2(new_n482), .ZN(new_n505));
  NAND3_X1  g304(.A1(new_n417), .A2(new_n426), .A3(new_n505), .ZN(new_n506));
  OAI21_X1  g305(.A(KEYINPUT35), .B1(new_n506), .B2(new_n502), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n440), .A2(new_n436), .ZN(new_n508));
  INV_X1    g307(.A(KEYINPUT35), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  NAND3_X1  g309(.A1(new_n501), .A2(new_n493), .A3(new_n497), .ZN(new_n511));
  NOR2_X1   g310(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  NAND4_X1  g311(.A1(new_n512), .A2(new_n426), .A3(new_n417), .A4(new_n505), .ZN(new_n513));
  AOI22_X1  g312(.A1(new_n488), .A2(new_n504), .B1(new_n507), .B2(new_n513), .ZN(new_n514));
  XNOR2_X1  g313(.A(G15gat), .B(G22gat), .ZN(new_n515));
  INV_X1    g314(.A(G1gat), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n516), .A2(KEYINPUT16), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n515), .A2(new_n517), .ZN(new_n518));
  OAI21_X1  g317(.A(new_n518), .B1(G1gat), .B2(new_n515), .ZN(new_n519));
  XNOR2_X1  g318(.A(new_n519), .B(G8gat), .ZN(new_n520));
  OAI21_X1  g319(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n521));
  INV_X1    g320(.A(new_n521), .ZN(new_n522));
  OR3_X1    g321(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n523));
  AOI21_X1  g322(.A(new_n522), .B1(new_n523), .B2(KEYINPUT87), .ZN(new_n524));
  OAI21_X1  g323(.A(new_n524), .B1(KEYINPUT87), .B2(new_n523), .ZN(new_n525));
  NAND2_X1  g324(.A1(G29gat), .A2(G36gat), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  INV_X1    g326(.A(G43gat), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n528), .A2(G50gat), .ZN(new_n529));
  NAND2_X1  g328(.A1(new_n410), .A2(G43gat), .ZN(new_n530));
  NAND3_X1  g329(.A1(new_n529), .A2(new_n530), .A3(KEYINPUT15), .ZN(new_n531));
  INV_X1    g330(.A(new_n531), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n527), .A2(new_n532), .ZN(new_n533));
  NOR2_X1   g332(.A1(new_n410), .A2(G43gat), .ZN(new_n534));
  INV_X1    g333(.A(KEYINPUT88), .ZN(new_n535));
  AOI21_X1  g334(.A(new_n534), .B1(new_n535), .B2(new_n530), .ZN(new_n536));
  NAND3_X1  g335(.A1(new_n410), .A2(KEYINPUT88), .A3(G43gat), .ZN(new_n537));
  AOI21_X1  g336(.A(KEYINPUT15), .B1(new_n536), .B2(new_n537), .ZN(new_n538));
  XNOR2_X1  g337(.A(new_n526), .B(KEYINPUT89), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n523), .A2(new_n521), .ZN(new_n540));
  NAND3_X1  g339(.A1(new_n539), .A2(new_n540), .A3(new_n531), .ZN(new_n541));
  NOR2_X1   g340(.A1(new_n538), .A2(new_n541), .ZN(new_n542));
  INV_X1    g341(.A(new_n542), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n533), .A2(new_n543), .ZN(new_n544));
  INV_X1    g343(.A(KEYINPUT17), .ZN(new_n545));
  AOI21_X1  g344(.A(new_n520), .B1(new_n544), .B2(new_n545), .ZN(new_n546));
  AND4_X1   g345(.A1(KEYINPUT90), .A2(new_n533), .A3(KEYINPUT17), .A4(new_n543), .ZN(new_n547));
  AOI21_X1  g346(.A(new_n542), .B1(new_n527), .B2(new_n532), .ZN(new_n548));
  AOI21_X1  g347(.A(KEYINPUT90), .B1(new_n548), .B2(KEYINPUT17), .ZN(new_n549));
  OAI21_X1  g348(.A(new_n546), .B1(new_n547), .B2(new_n549), .ZN(new_n550));
  NAND2_X1  g349(.A1(G229gat), .A2(G233gat), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n544), .A2(new_n520), .ZN(new_n552));
  NAND3_X1  g351(.A1(new_n550), .A2(new_n551), .A3(new_n552), .ZN(new_n553));
  INV_X1    g352(.A(KEYINPUT18), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  NAND4_X1  g354(.A1(new_n550), .A2(KEYINPUT18), .A3(new_n551), .A4(new_n552), .ZN(new_n556));
  INV_X1    g355(.A(new_n520), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n557), .A2(new_n548), .ZN(new_n558));
  OR2_X1    g357(.A1(new_n558), .A2(KEYINPUT91), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n558), .A2(KEYINPUT91), .ZN(new_n560));
  NAND3_X1  g359(.A1(new_n559), .A2(new_n552), .A3(new_n560), .ZN(new_n561));
  XOR2_X1   g360(.A(new_n551), .B(KEYINPUT13), .Z(new_n562));
  NAND2_X1  g361(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  NAND3_X1  g362(.A1(new_n555), .A2(new_n556), .A3(new_n563), .ZN(new_n564));
  XNOR2_X1  g363(.A(G113gat), .B(G141gat), .ZN(new_n565));
  XNOR2_X1  g364(.A(new_n565), .B(G197gat), .ZN(new_n566));
  XOR2_X1   g365(.A(KEYINPUT11), .B(G169gat), .Z(new_n567));
  XNOR2_X1  g366(.A(new_n566), .B(new_n567), .ZN(new_n568));
  XOR2_X1   g367(.A(new_n568), .B(KEYINPUT12), .Z(new_n569));
  NAND2_X1  g368(.A1(new_n564), .A2(new_n569), .ZN(new_n570));
  INV_X1    g369(.A(new_n569), .ZN(new_n571));
  NAND4_X1  g370(.A1(new_n555), .A2(new_n563), .A3(new_n571), .A4(new_n556), .ZN(new_n572));
  NAND3_X1  g371(.A1(new_n570), .A2(KEYINPUT92), .A3(new_n572), .ZN(new_n573));
  INV_X1    g372(.A(KEYINPUT92), .ZN(new_n574));
  NAND3_X1  g373(.A1(new_n564), .A2(new_n574), .A3(new_n569), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n573), .A2(new_n575), .ZN(new_n576));
  NOR2_X1   g375(.A1(new_n514), .A2(new_n576), .ZN(new_n577));
  NAND2_X1  g376(.A1(G232gat), .A2(G233gat), .ZN(new_n578));
  XNOR2_X1  g377(.A(new_n578), .B(KEYINPUT93), .ZN(new_n579));
  INV_X1    g378(.A(KEYINPUT41), .ZN(new_n580));
  NAND2_X1  g379(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  XOR2_X1   g380(.A(new_n581), .B(KEYINPUT94), .Z(new_n582));
  XNOR2_X1  g381(.A(G134gat), .B(G162gat), .ZN(new_n583));
  XOR2_X1   g382(.A(new_n582), .B(new_n583), .Z(new_n584));
  INV_X1    g383(.A(new_n584), .ZN(new_n585));
  XOR2_X1   g384(.A(G99gat), .B(G106gat), .Z(new_n586));
  XNOR2_X1  g385(.A(KEYINPUT95), .B(KEYINPUT7), .ZN(new_n587));
  INV_X1    g386(.A(G85gat), .ZN(new_n588));
  INV_X1    g387(.A(G92gat), .ZN(new_n589));
  NOR2_X1   g388(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  NAND2_X1  g389(.A1(new_n587), .A2(new_n590), .ZN(new_n591));
  NAND2_X1  g390(.A1(G99gat), .A2(G106gat), .ZN(new_n592));
  AOI22_X1  g391(.A1(KEYINPUT8), .A2(new_n592), .B1(new_n588), .B2(new_n589), .ZN(new_n593));
  NAND2_X1  g392(.A1(new_n591), .A2(new_n593), .ZN(new_n594));
  NOR2_X1   g393(.A1(new_n587), .A2(new_n590), .ZN(new_n595));
  OAI21_X1  g394(.A(new_n586), .B1(new_n594), .B2(new_n595), .ZN(new_n596));
  XOR2_X1   g395(.A(KEYINPUT95), .B(KEYINPUT7), .Z(new_n597));
  INV_X1    g396(.A(new_n590), .ZN(new_n598));
  NAND2_X1  g397(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  INV_X1    g398(.A(new_n586), .ZN(new_n600));
  NAND4_X1  g399(.A1(new_n599), .A2(new_n600), .A3(new_n591), .A4(new_n593), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n596), .A2(new_n601), .ZN(new_n602));
  INV_X1    g401(.A(new_n602), .ZN(new_n603));
  AOI21_X1  g402(.A(new_n603), .B1(new_n544), .B2(new_n545), .ZN(new_n604));
  OAI21_X1  g403(.A(new_n604), .B1(new_n547), .B2(new_n549), .ZN(new_n605));
  XNOR2_X1  g404(.A(G190gat), .B(G218gat), .ZN(new_n606));
  INV_X1    g405(.A(new_n606), .ZN(new_n607));
  NOR2_X1   g406(.A1(new_n579), .A2(new_n580), .ZN(new_n608));
  AOI21_X1  g407(.A(new_n608), .B1(new_n544), .B2(new_n603), .ZN(new_n609));
  NAND3_X1  g408(.A1(new_n605), .A2(new_n607), .A3(new_n609), .ZN(new_n610));
  INV_X1    g409(.A(new_n610), .ZN(new_n611));
  AOI21_X1  g410(.A(new_n607), .B1(new_n605), .B2(new_n609), .ZN(new_n612));
  XNOR2_X1  g411(.A(KEYINPUT96), .B(KEYINPUT97), .ZN(new_n613));
  INV_X1    g412(.A(new_n613), .ZN(new_n614));
  NOR3_X1   g413(.A1(new_n611), .A2(new_n612), .A3(new_n614), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n605), .A2(new_n609), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n616), .A2(new_n606), .ZN(new_n617));
  AOI21_X1  g416(.A(new_n613), .B1(new_n617), .B2(new_n610), .ZN(new_n618));
  OAI21_X1  g417(.A(new_n585), .B1(new_n615), .B2(new_n618), .ZN(new_n619));
  INV_X1    g418(.A(KEYINPUT98), .ZN(new_n620));
  NAND2_X1  g419(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  OAI211_X1 g420(.A(KEYINPUT98), .B(new_n585), .C1(new_n615), .C2(new_n618), .ZN(new_n622));
  OAI21_X1  g421(.A(new_n614), .B1(new_n611), .B2(new_n612), .ZN(new_n623));
  NAND3_X1  g422(.A1(new_n617), .A2(new_n610), .A3(new_n613), .ZN(new_n624));
  NAND3_X1  g423(.A1(new_n623), .A2(new_n624), .A3(new_n584), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n625), .A2(KEYINPUT99), .ZN(new_n626));
  INV_X1    g425(.A(KEYINPUT99), .ZN(new_n627));
  NAND4_X1  g426(.A1(new_n623), .A2(new_n624), .A3(new_n627), .A4(new_n584), .ZN(new_n628));
  AOI22_X1  g427(.A1(new_n621), .A2(new_n622), .B1(new_n626), .B2(new_n628), .ZN(new_n629));
  XNOR2_X1  g428(.A(G57gat), .B(G64gat), .ZN(new_n630));
  INV_X1    g429(.A(KEYINPUT9), .ZN(new_n631));
  NAND2_X1  g430(.A1(G71gat), .A2(G78gat), .ZN(new_n632));
  AOI21_X1  g431(.A(new_n630), .B1(new_n631), .B2(new_n632), .ZN(new_n633));
  OR2_X1    g432(.A1(G71gat), .A2(G78gat), .ZN(new_n634));
  NAND2_X1  g433(.A1(new_n634), .A2(new_n632), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n633), .A2(new_n635), .ZN(new_n636));
  OAI211_X1 g435(.A(new_n632), .B(new_n634), .C1(new_n630), .C2(new_n631), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  INV_X1    g437(.A(KEYINPUT21), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  NAND2_X1  g439(.A1(G231gat), .A2(G233gat), .ZN(new_n641));
  XNOR2_X1  g440(.A(new_n640), .B(new_n641), .ZN(new_n642));
  XNOR2_X1  g441(.A(new_n642), .B(G127gat), .ZN(new_n643));
  OAI21_X1  g442(.A(new_n557), .B1(new_n639), .B2(new_n638), .ZN(new_n644));
  XNOR2_X1  g443(.A(new_n643), .B(new_n644), .ZN(new_n645));
  XOR2_X1   g444(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n646));
  XNOR2_X1  g445(.A(new_n646), .B(G155gat), .ZN(new_n647));
  XOR2_X1   g446(.A(G183gat), .B(G211gat), .Z(new_n648));
  XNOR2_X1  g447(.A(new_n647), .B(new_n648), .ZN(new_n649));
  XNOR2_X1  g448(.A(new_n645), .B(new_n649), .ZN(new_n650));
  INV_X1    g449(.A(new_n650), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n629), .A2(new_n651), .ZN(new_n652));
  NAND2_X1  g451(.A1(G230gat), .A2(G233gat), .ZN(new_n653));
  INV_X1    g452(.A(new_n653), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n602), .A2(new_n638), .ZN(new_n655));
  INV_X1    g454(.A(KEYINPUT10), .ZN(new_n656));
  NAND4_X1  g455(.A1(new_n596), .A2(new_n637), .A3(new_n636), .A4(new_n601), .ZN(new_n657));
  NAND3_X1  g456(.A1(new_n655), .A2(new_n656), .A3(new_n657), .ZN(new_n658));
  OR2_X1    g457(.A1(new_n657), .A2(new_n656), .ZN(new_n659));
  AOI21_X1  g458(.A(new_n654), .B1(new_n658), .B2(new_n659), .ZN(new_n660));
  INV_X1    g459(.A(new_n660), .ZN(new_n661));
  NAND2_X1  g460(.A1(new_n655), .A2(new_n657), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n662), .A2(new_n654), .ZN(new_n663));
  XNOR2_X1  g462(.A(G120gat), .B(G148gat), .ZN(new_n664));
  XNOR2_X1  g463(.A(G176gat), .B(G204gat), .ZN(new_n665));
  XOR2_X1   g464(.A(new_n664), .B(new_n665), .Z(new_n666));
  NAND3_X1  g465(.A1(new_n661), .A2(new_n663), .A3(new_n666), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n667), .A2(KEYINPUT100), .ZN(new_n668));
  INV_X1    g467(.A(KEYINPUT100), .ZN(new_n669));
  NAND4_X1  g468(.A1(new_n661), .A2(new_n663), .A3(new_n669), .A4(new_n666), .ZN(new_n670));
  NAND2_X1  g469(.A1(new_n668), .A2(new_n670), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n661), .A2(new_n663), .ZN(new_n672));
  INV_X1    g471(.A(new_n666), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n671), .A2(new_n674), .ZN(new_n675));
  NOR2_X1   g474(.A1(new_n652), .A2(new_n675), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n577), .A2(new_n676), .ZN(new_n677));
  OR2_X1    g476(.A1(new_n500), .A2(KEYINPUT101), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n500), .A2(KEYINPUT101), .ZN(new_n679));
  NAND2_X1  g478(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  NOR2_X1   g479(.A1(new_n677), .A2(new_n680), .ZN(new_n681));
  XNOR2_X1  g480(.A(new_n681), .B(new_n516), .ZN(G1324gat));
  NAND3_X1  g481(.A1(new_n577), .A2(new_n511), .A3(new_n676), .ZN(new_n683));
  AND2_X1   g482(.A1(new_n683), .A2(G8gat), .ZN(new_n684));
  XNOR2_X1  g483(.A(KEYINPUT16), .B(G8gat), .ZN(new_n685));
  NOR2_X1   g484(.A1(new_n683), .A2(new_n685), .ZN(new_n686));
  OAI21_X1  g485(.A(KEYINPUT42), .B1(new_n684), .B2(new_n686), .ZN(new_n687));
  OAI21_X1  g486(.A(new_n687), .B1(KEYINPUT42), .B2(new_n686), .ZN(G1325gat));
  OAI21_X1  g487(.A(G15gat), .B1(new_n677), .B2(new_n487), .ZN(new_n689));
  INV_X1    g488(.A(new_n505), .ZN(new_n690));
  OR2_X1    g489(.A1(new_n690), .A2(G15gat), .ZN(new_n691));
  OAI21_X1  g490(.A(new_n689), .B1(new_n677), .B2(new_n691), .ZN(G1326gat));
  NAND3_X1  g491(.A1(new_n577), .A2(new_n503), .A3(new_n676), .ZN(new_n693));
  XNOR2_X1  g492(.A(new_n693), .B(KEYINPUT102), .ZN(new_n694));
  XNOR2_X1  g493(.A(KEYINPUT43), .B(G22gat), .ZN(new_n695));
  XNOR2_X1  g494(.A(new_n694), .B(new_n695), .ZN(G1327gat));
  NOR2_X1   g495(.A1(new_n651), .A2(new_n675), .ZN(new_n697));
  NAND2_X1  g496(.A1(new_n621), .A2(new_n622), .ZN(new_n698));
  NAND2_X1  g497(.A1(new_n626), .A2(new_n628), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n697), .A2(new_n700), .ZN(new_n701));
  NOR3_X1   g500(.A1(new_n701), .A2(G29gat), .A3(new_n680), .ZN(new_n702));
  NAND2_X1  g501(.A1(new_n577), .A2(new_n702), .ZN(new_n703));
  XNOR2_X1  g502(.A(new_n703), .B(KEYINPUT103), .ZN(new_n704));
  XNOR2_X1  g503(.A(new_n704), .B(KEYINPUT45), .ZN(new_n705));
  INV_X1    g504(.A(KEYINPUT44), .ZN(new_n706));
  OAI21_X1  g505(.A(new_n706), .B1(new_n514), .B2(new_n629), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n507), .A2(new_n513), .ZN(new_n708));
  NAND3_X1  g507(.A1(new_n504), .A2(new_n442), .A3(new_n487), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  NAND3_X1  g509(.A1(new_n710), .A2(KEYINPUT44), .A3(new_n700), .ZN(new_n711));
  AND2_X1   g510(.A1(new_n707), .A2(new_n711), .ZN(new_n712));
  NOR3_X1   g511(.A1(new_n651), .A2(new_n576), .A3(new_n675), .ZN(new_n713));
  NAND2_X1  g512(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  NOR3_X1   g513(.A1(new_n714), .A2(KEYINPUT104), .A3(new_n680), .ZN(new_n715));
  OAI21_X1  g514(.A(KEYINPUT104), .B1(new_n714), .B2(new_n680), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n716), .A2(G29gat), .ZN(new_n717));
  OAI21_X1  g516(.A(new_n705), .B1(new_n715), .B2(new_n717), .ZN(G1328gat));
  INV_X1    g517(.A(new_n511), .ZN(new_n719));
  NOR3_X1   g518(.A1(new_n701), .A2(G36gat), .A3(new_n719), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n577), .A2(new_n720), .ZN(new_n721));
  XOR2_X1   g520(.A(new_n721), .B(KEYINPUT46), .Z(new_n722));
  OAI21_X1  g521(.A(KEYINPUT105), .B1(new_n714), .B2(new_n719), .ZN(new_n723));
  NAND2_X1  g522(.A1(new_n723), .A2(G36gat), .ZN(new_n724));
  NOR3_X1   g523(.A1(new_n714), .A2(KEYINPUT105), .A3(new_n719), .ZN(new_n725));
  OAI21_X1  g524(.A(new_n722), .B1(new_n724), .B2(new_n725), .ZN(G1329gat));
  OAI21_X1  g525(.A(G43gat), .B1(new_n714), .B2(new_n487), .ZN(new_n727));
  INV_X1    g526(.A(new_n701), .ZN(new_n728));
  NAND4_X1  g527(.A1(new_n577), .A2(new_n528), .A3(new_n505), .A4(new_n728), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n727), .A2(new_n729), .ZN(new_n730));
  INV_X1    g529(.A(KEYINPUT47), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  NAND3_X1  g531(.A1(new_n727), .A2(KEYINPUT47), .A3(new_n729), .ZN(new_n733));
  NAND2_X1  g532(.A1(new_n732), .A2(new_n733), .ZN(G1330gat));
  INV_X1    g533(.A(KEYINPUT106), .ZN(new_n735));
  INV_X1    g534(.A(new_n503), .ZN(new_n736));
  OAI21_X1  g535(.A(new_n735), .B1(new_n736), .B2(G50gat), .ZN(new_n737));
  NAND3_X1  g536(.A1(new_n503), .A2(KEYINPUT106), .A3(new_n410), .ZN(new_n738));
  AND4_X1   g537(.A1(new_n577), .A2(new_n728), .A3(new_n737), .A4(new_n738), .ZN(new_n739));
  NAND3_X1  g538(.A1(new_n712), .A2(new_n503), .A3(new_n713), .ZN(new_n740));
  AOI21_X1  g539(.A(new_n739), .B1(new_n740), .B2(G50gat), .ZN(new_n741));
  XNOR2_X1  g540(.A(KEYINPUT107), .B(KEYINPUT48), .ZN(new_n742));
  XOR2_X1   g541(.A(new_n741), .B(new_n742), .Z(G1331gat));
  INV_X1    g542(.A(new_n576), .ZN(new_n744));
  INV_X1    g543(.A(new_n675), .ZN(new_n745));
  NOR4_X1   g544(.A1(new_n514), .A2(new_n744), .A3(new_n745), .A4(new_n652), .ZN(new_n746));
  INV_X1    g545(.A(KEYINPUT108), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n680), .A2(new_n747), .ZN(new_n748));
  NAND3_X1  g547(.A1(new_n678), .A2(KEYINPUT108), .A3(new_n679), .ZN(new_n749));
  NAND2_X1  g548(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  NAND2_X1  g549(.A1(new_n746), .A2(new_n750), .ZN(new_n751));
  XNOR2_X1  g550(.A(new_n751), .B(G57gat), .ZN(G1332gat));
  INV_X1    g551(.A(KEYINPUT49), .ZN(new_n753));
  INV_X1    g552(.A(G64gat), .ZN(new_n754));
  OAI211_X1 g553(.A(new_n746), .B(new_n511), .C1(new_n753), .C2(new_n754), .ZN(new_n755));
  XNOR2_X1  g554(.A(new_n755), .B(KEYINPUT109), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n753), .A2(new_n754), .ZN(new_n757));
  XNOR2_X1  g556(.A(new_n756), .B(new_n757), .ZN(G1333gat));
  INV_X1    g557(.A(new_n487), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n746), .A2(new_n759), .ZN(new_n760));
  NOR2_X1   g559(.A1(new_n690), .A2(G71gat), .ZN(new_n761));
  AOI22_X1  g560(.A1(new_n760), .A2(G71gat), .B1(new_n746), .B2(new_n761), .ZN(new_n762));
  XNOR2_X1  g561(.A(new_n762), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g562(.A1(new_n746), .A2(new_n503), .ZN(new_n764));
  XOR2_X1   g563(.A(KEYINPUT110), .B(G78gat), .Z(new_n765));
  XNOR2_X1  g564(.A(new_n764), .B(new_n765), .ZN(G1335gat));
  NOR3_X1   g565(.A1(new_n744), .A2(new_n651), .A3(new_n745), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n712), .A2(new_n767), .ZN(new_n768));
  OAI21_X1  g567(.A(G85gat), .B1(new_n768), .B2(new_n680), .ZN(new_n769));
  NOR2_X1   g568(.A1(new_n744), .A2(new_n651), .ZN(new_n770));
  AND4_X1   g569(.A1(KEYINPUT51), .A2(new_n710), .A3(new_n700), .A4(new_n770), .ZN(new_n771));
  AOI21_X1  g570(.A(new_n629), .B1(new_n708), .B2(new_n709), .ZN(new_n772));
  AOI21_X1  g571(.A(KEYINPUT51), .B1(new_n772), .B2(new_n770), .ZN(new_n773));
  OR2_X1    g572(.A1(new_n771), .A2(new_n773), .ZN(new_n774));
  INV_X1    g573(.A(new_n680), .ZN(new_n775));
  NAND4_X1  g574(.A1(new_n774), .A2(new_n588), .A3(new_n775), .A4(new_n675), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n769), .A2(new_n776), .ZN(G1336gat));
  INV_X1    g576(.A(KEYINPUT52), .ZN(new_n778));
  NAND4_X1  g577(.A1(new_n774), .A2(new_n589), .A3(new_n511), .A4(new_n675), .ZN(new_n779));
  INV_X1    g578(.A(KEYINPUT111), .ZN(new_n780));
  AOI21_X1  g579(.A(new_n778), .B1(new_n779), .B2(new_n780), .ZN(new_n781));
  OAI21_X1  g580(.A(G92gat), .B1(new_n768), .B2(new_n719), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n782), .A2(new_n779), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n781), .A2(new_n783), .ZN(new_n784));
  OAI211_X1 g583(.A(new_n782), .B(new_n779), .C1(new_n780), .C2(new_n778), .ZN(new_n785));
  NAND2_X1  g584(.A1(new_n784), .A2(new_n785), .ZN(G1337gat));
  OAI21_X1  g585(.A(G99gat), .B1(new_n768), .B2(new_n487), .ZN(new_n787));
  NOR3_X1   g586(.A1(new_n690), .A2(G99gat), .A3(new_n745), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n774), .A2(new_n788), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n787), .A2(new_n789), .ZN(G1338gat));
  NAND4_X1  g589(.A1(new_n707), .A2(new_n503), .A3(new_n711), .A4(new_n767), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n791), .A2(G106gat), .ZN(new_n792));
  INV_X1    g591(.A(KEYINPUT53), .ZN(new_n793));
  NOR3_X1   g592(.A1(new_n736), .A2(G106gat), .A3(new_n745), .ZN(new_n794));
  OAI21_X1  g593(.A(new_n794), .B1(new_n771), .B2(new_n773), .ZN(new_n795));
  NAND3_X1  g594(.A1(new_n792), .A2(new_n793), .A3(new_n795), .ZN(new_n796));
  INV_X1    g595(.A(KEYINPUT113), .ZN(new_n797));
  INV_X1    g596(.A(KEYINPUT112), .ZN(new_n798));
  AOI22_X1  g597(.A1(new_n795), .A2(new_n798), .B1(G106gat), .B2(new_n791), .ZN(new_n799));
  OAI211_X1 g598(.A(KEYINPUT112), .B(new_n794), .C1(new_n771), .C2(new_n773), .ZN(new_n800));
  AOI211_X1 g599(.A(new_n797), .B(new_n793), .C1(new_n799), .C2(new_n800), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n795), .A2(new_n798), .ZN(new_n802));
  NAND3_X1  g601(.A1(new_n802), .A2(new_n800), .A3(new_n792), .ZN(new_n803));
  AOI21_X1  g602(.A(KEYINPUT113), .B1(new_n803), .B2(KEYINPUT53), .ZN(new_n804));
  OAI21_X1  g603(.A(new_n796), .B1(new_n801), .B2(new_n804), .ZN(G1339gat));
  NAND4_X1  g604(.A1(new_n629), .A2(new_n576), .A3(new_n745), .A4(new_n651), .ZN(new_n806));
  XNOR2_X1  g605(.A(new_n806), .B(KEYINPUT114), .ZN(new_n807));
  NAND3_X1  g606(.A1(new_n658), .A2(new_n659), .A3(new_n654), .ZN(new_n808));
  NAND3_X1  g607(.A1(new_n661), .A2(KEYINPUT54), .A3(new_n808), .ZN(new_n809));
  INV_X1    g608(.A(KEYINPUT54), .ZN(new_n810));
  AOI211_X1 g609(.A(KEYINPUT115), .B(new_n666), .C1(new_n660), .C2(new_n810), .ZN(new_n811));
  INV_X1    g610(.A(KEYINPUT115), .ZN(new_n812));
  AND3_X1   g611(.A1(new_n655), .A2(new_n656), .A3(new_n657), .ZN(new_n813));
  NOR2_X1   g612(.A1(new_n657), .A2(new_n656), .ZN(new_n814));
  OAI211_X1 g613(.A(new_n810), .B(new_n653), .C1(new_n813), .C2(new_n814), .ZN(new_n815));
  AOI21_X1  g614(.A(new_n812), .B1(new_n815), .B2(new_n673), .ZN(new_n816));
  OAI211_X1 g615(.A(KEYINPUT55), .B(new_n809), .C1(new_n811), .C2(new_n816), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n817), .A2(new_n671), .ZN(new_n818));
  AOI211_X1 g617(.A(KEYINPUT54), .B(new_n654), .C1(new_n658), .C2(new_n659), .ZN(new_n819));
  OAI21_X1  g618(.A(KEYINPUT115), .B1(new_n819), .B2(new_n666), .ZN(new_n820));
  NAND3_X1  g619(.A1(new_n815), .A2(new_n812), .A3(new_n673), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  AOI21_X1  g621(.A(KEYINPUT55), .B1(new_n822), .B2(new_n809), .ZN(new_n823));
  OAI21_X1  g622(.A(KEYINPUT116), .B1(new_n818), .B2(new_n823), .ZN(new_n824));
  OAI21_X1  g623(.A(new_n809), .B1(new_n811), .B2(new_n816), .ZN(new_n825));
  INV_X1    g624(.A(KEYINPUT55), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n825), .A2(new_n826), .ZN(new_n827));
  INV_X1    g626(.A(KEYINPUT116), .ZN(new_n828));
  NAND4_X1  g627(.A1(new_n827), .A2(new_n828), .A3(new_n671), .A4(new_n817), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n824), .A2(new_n829), .ZN(new_n830));
  AOI21_X1  g629(.A(new_n551), .B1(new_n550), .B2(new_n552), .ZN(new_n831));
  INV_X1    g630(.A(KEYINPUT117), .ZN(new_n832));
  OAI22_X1  g631(.A1(new_n831), .A2(new_n832), .B1(new_n561), .B2(new_n562), .ZN(new_n833));
  AND2_X1   g632(.A1(new_n831), .A2(new_n832), .ZN(new_n834));
  OAI21_X1  g633(.A(new_n568), .B1(new_n833), .B2(new_n834), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n835), .A2(new_n572), .ZN(new_n836));
  NOR3_X1   g635(.A1(new_n629), .A2(new_n830), .A3(new_n836), .ZN(new_n837));
  NAND4_X1  g636(.A1(new_n824), .A2(new_n829), .A3(new_n575), .A4(new_n573), .ZN(new_n838));
  NAND3_X1  g637(.A1(new_n835), .A2(new_n675), .A3(new_n572), .ZN(new_n839));
  NAND2_X1  g638(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  AOI21_X1  g639(.A(new_n700), .B1(new_n840), .B2(KEYINPUT118), .ZN(new_n841));
  INV_X1    g640(.A(KEYINPUT118), .ZN(new_n842));
  NAND3_X1  g641(.A1(new_n838), .A2(new_n842), .A3(new_n839), .ZN(new_n843));
  AOI21_X1  g642(.A(new_n837), .B1(new_n841), .B2(new_n843), .ZN(new_n844));
  OAI21_X1  g643(.A(new_n807), .B1(new_n844), .B2(new_n651), .ZN(new_n845));
  INV_X1    g644(.A(new_n845), .ZN(new_n846));
  NOR2_X1   g645(.A1(new_n846), .A2(new_n503), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n775), .A2(new_n719), .ZN(new_n848));
  NOR2_X1   g647(.A1(new_n848), .A2(new_n690), .ZN(new_n849));
  NAND2_X1  g648(.A1(new_n847), .A2(new_n849), .ZN(new_n850));
  NOR3_X1   g649(.A1(new_n850), .A2(new_n227), .A3(new_n576), .ZN(new_n851));
  NAND2_X1  g650(.A1(new_n845), .A2(new_n750), .ZN(new_n852));
  NOR3_X1   g651(.A1(new_n852), .A2(new_n511), .A3(new_n506), .ZN(new_n853));
  AOI21_X1  g652(.A(G113gat), .B1(new_n853), .B2(new_n744), .ZN(new_n854));
  NOR2_X1   g653(.A1(new_n851), .A2(new_n854), .ZN(G1340gat));
  NAND3_X1  g654(.A1(new_n853), .A2(new_n225), .A3(new_n675), .ZN(new_n856));
  NAND3_X1  g655(.A1(new_n847), .A2(new_n675), .A3(new_n849), .ZN(new_n857));
  INV_X1    g656(.A(KEYINPUT119), .ZN(new_n858));
  AND3_X1   g657(.A1(new_n857), .A2(new_n858), .A3(G120gat), .ZN(new_n859));
  AOI21_X1  g658(.A(new_n858), .B1(new_n857), .B2(G120gat), .ZN(new_n860));
  OAI21_X1  g659(.A(new_n856), .B1(new_n859), .B2(new_n860), .ZN(G1341gat));
  OAI21_X1  g660(.A(G127gat), .B1(new_n850), .B2(new_n650), .ZN(new_n862));
  INV_X1    g661(.A(G127gat), .ZN(new_n863));
  NAND3_X1  g662(.A1(new_n853), .A2(new_n863), .A3(new_n651), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n862), .A2(new_n864), .ZN(G1342gat));
  NAND3_X1  g664(.A1(new_n847), .A2(new_n700), .A3(new_n849), .ZN(new_n866));
  INV_X1    g665(.A(new_n750), .ZN(new_n867));
  AND3_X1   g666(.A1(new_n838), .A2(new_n842), .A3(new_n839), .ZN(new_n868));
  AOI21_X1  g667(.A(new_n842), .B1(new_n838), .B2(new_n839), .ZN(new_n869));
  NOR3_X1   g668(.A1(new_n868), .A2(new_n869), .A3(new_n700), .ZN(new_n870));
  OAI21_X1  g669(.A(new_n650), .B1(new_n870), .B2(new_n837), .ZN(new_n871));
  AOI21_X1  g670(.A(new_n867), .B1(new_n871), .B2(new_n807), .ZN(new_n872));
  INV_X1    g671(.A(new_n506), .ZN(new_n873));
  NAND2_X1  g672(.A1(new_n700), .A2(new_n719), .ZN(new_n874));
  NOR2_X1   g673(.A1(new_n874), .A2(G134gat), .ZN(new_n875));
  NAND3_X1  g674(.A1(new_n872), .A2(new_n873), .A3(new_n875), .ZN(new_n876));
  AOI22_X1  g675(.A1(new_n866), .A2(G134gat), .B1(KEYINPUT56), .B2(new_n876), .ZN(new_n877));
  OR2_X1    g676(.A1(new_n876), .A2(KEYINPUT56), .ZN(new_n878));
  AND2_X1   g677(.A1(new_n878), .A2(KEYINPUT120), .ZN(new_n879));
  NOR2_X1   g678(.A1(new_n878), .A2(KEYINPUT120), .ZN(new_n880));
  OAI21_X1  g679(.A(new_n877), .B1(new_n879), .B2(new_n880), .ZN(G1343gat));
  NOR2_X1   g680(.A1(new_n848), .A2(new_n759), .ZN(new_n882));
  AOI21_X1  g681(.A(KEYINPUT57), .B1(new_n845), .B2(new_n503), .ZN(new_n883));
  NOR2_X1   g682(.A1(new_n818), .A2(new_n823), .ZN(new_n884));
  INV_X1    g683(.A(new_n884), .ZN(new_n885));
  OAI21_X1  g684(.A(new_n839), .B1(new_n885), .B2(new_n576), .ZN(new_n886));
  AND2_X1   g685(.A1(new_n886), .A2(new_n629), .ZN(new_n887));
  OAI21_X1  g686(.A(new_n650), .B1(new_n887), .B2(new_n837), .ZN(new_n888));
  NAND2_X1  g687(.A1(new_n807), .A2(new_n888), .ZN(new_n889));
  INV_X1    g688(.A(KEYINPUT57), .ZN(new_n890));
  NOR2_X1   g689(.A1(new_n736), .A2(new_n890), .ZN(new_n891));
  AND2_X1   g690(.A1(new_n889), .A2(new_n891), .ZN(new_n892));
  OAI211_X1 g691(.A(new_n744), .B(new_n882), .C1(new_n883), .C2(new_n892), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n893), .A2(G141gat), .ZN(new_n894));
  NOR2_X1   g693(.A1(new_n759), .A2(new_n736), .ZN(new_n895));
  INV_X1    g694(.A(new_n895), .ZN(new_n896));
  INV_X1    g695(.A(KEYINPUT121), .ZN(new_n897));
  AOI21_X1  g696(.A(new_n896), .B1(new_n872), .B2(new_n897), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n852), .A2(KEYINPUT121), .ZN(new_n899));
  NOR2_X1   g698(.A1(new_n576), .A2(G141gat), .ZN(new_n900));
  NAND4_X1  g699(.A1(new_n898), .A2(new_n719), .A3(new_n899), .A4(new_n900), .ZN(new_n901));
  NAND2_X1  g700(.A1(new_n894), .A2(new_n901), .ZN(new_n902));
  NAND2_X1  g701(.A1(new_n902), .A2(KEYINPUT58), .ZN(new_n903));
  INV_X1    g702(.A(KEYINPUT58), .ZN(new_n904));
  NAND3_X1  g703(.A1(new_n894), .A2(new_n904), .A3(new_n901), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n903), .A2(new_n905), .ZN(G1344gat));
  NOR2_X1   g705(.A1(new_n745), .A2(G148gat), .ZN(new_n907));
  NAND4_X1  g706(.A1(new_n898), .A2(new_n719), .A3(new_n899), .A4(new_n907), .ZN(new_n908));
  INV_X1    g707(.A(KEYINPUT59), .ZN(new_n909));
  NAND2_X1  g708(.A1(new_n882), .A2(new_n675), .ZN(new_n910));
  NAND2_X1  g709(.A1(new_n845), .A2(new_n891), .ZN(new_n911));
  NOR2_X1   g710(.A1(new_n629), .A2(new_n836), .ZN(new_n912));
  AOI22_X1  g711(.A1(new_n912), .A2(new_n884), .B1(new_n886), .B2(new_n629), .ZN(new_n913));
  OAI21_X1  g712(.A(new_n806), .B1(new_n913), .B2(new_n651), .ZN(new_n914));
  NAND2_X1  g713(.A1(new_n914), .A2(new_n503), .ZN(new_n915));
  NAND2_X1  g714(.A1(new_n915), .A2(new_n890), .ZN(new_n916));
  AOI21_X1  g715(.A(new_n910), .B1(new_n911), .B2(new_n916), .ZN(new_n917));
  INV_X1    g716(.A(KEYINPUT122), .ZN(new_n918));
  AOI21_X1  g717(.A(new_n208), .B1(new_n917), .B2(new_n918), .ZN(new_n919));
  AOI22_X1  g718(.A1(new_n845), .A2(new_n891), .B1(new_n915), .B2(new_n890), .ZN(new_n920));
  OAI21_X1  g719(.A(KEYINPUT122), .B1(new_n920), .B2(new_n910), .ZN(new_n921));
  AOI21_X1  g720(.A(new_n909), .B1(new_n919), .B2(new_n921), .ZN(new_n922));
  NAND2_X1  g721(.A1(new_n909), .A2(G148gat), .ZN(new_n923));
  INV_X1    g722(.A(new_n882), .ZN(new_n924));
  INV_X1    g723(.A(new_n883), .ZN(new_n925));
  INV_X1    g724(.A(new_n892), .ZN(new_n926));
  AOI21_X1  g725(.A(new_n924), .B1(new_n925), .B2(new_n926), .ZN(new_n927));
  AOI21_X1  g726(.A(new_n923), .B1(new_n927), .B2(new_n675), .ZN(new_n928));
  OAI21_X1  g727(.A(new_n908), .B1(new_n922), .B2(new_n928), .ZN(G1345gat));
  NAND2_X1  g728(.A1(new_n927), .A2(new_n651), .ZN(new_n930));
  NAND2_X1  g729(.A1(new_n930), .A2(G155gat), .ZN(new_n931));
  NOR2_X1   g730(.A1(new_n650), .A2(G155gat), .ZN(new_n932));
  NAND4_X1  g731(.A1(new_n898), .A2(new_n719), .A3(new_n899), .A4(new_n932), .ZN(new_n933));
  NAND2_X1  g732(.A1(new_n931), .A2(new_n933), .ZN(G1346gat));
  NAND2_X1  g733(.A1(new_n927), .A2(new_n700), .ZN(new_n935));
  NAND2_X1  g734(.A1(new_n935), .A2(new_n215), .ZN(new_n936));
  NAND2_X1  g735(.A1(new_n898), .A2(new_n899), .ZN(new_n937));
  OR2_X1    g736(.A1(new_n874), .A2(new_n215), .ZN(new_n938));
  OAI21_X1  g737(.A(new_n936), .B1(new_n937), .B2(new_n938), .ZN(G1347gat));
  NAND4_X1  g738(.A1(new_n748), .A2(new_n511), .A3(new_n505), .A4(new_n749), .ZN(new_n940));
  XNOR2_X1  g739(.A(new_n940), .B(KEYINPUT124), .ZN(new_n941));
  NAND2_X1  g740(.A1(new_n847), .A2(new_n941), .ZN(new_n942));
  NOR3_X1   g741(.A1(new_n942), .A2(new_n307), .A3(new_n576), .ZN(new_n943));
  NOR2_X1   g742(.A1(new_n846), .A2(new_n775), .ZN(new_n944));
  NAND2_X1  g743(.A1(new_n873), .A2(new_n511), .ZN(new_n945));
  XNOR2_X1  g744(.A(new_n945), .B(KEYINPUT123), .ZN(new_n946));
  NAND2_X1  g745(.A1(new_n944), .A2(new_n946), .ZN(new_n947));
  INV_X1    g746(.A(new_n947), .ZN(new_n948));
  NAND2_X1  g747(.A1(new_n948), .A2(new_n744), .ZN(new_n949));
  AOI21_X1  g748(.A(new_n943), .B1(new_n307), .B2(new_n949), .ZN(G1348gat));
  AOI21_X1  g749(.A(G176gat), .B1(new_n948), .B2(new_n675), .ZN(new_n951));
  INV_X1    g750(.A(new_n942), .ZN(new_n952));
  AOI21_X1  g751(.A(new_n745), .B1(new_n324), .B2(new_n326), .ZN(new_n953));
  AOI21_X1  g752(.A(new_n951), .B1(new_n952), .B2(new_n953), .ZN(G1349gat));
  NAND3_X1  g753(.A1(new_n847), .A2(new_n651), .A3(new_n941), .ZN(new_n955));
  NAND2_X1  g754(.A1(new_n955), .A2(G183gat), .ZN(new_n956));
  NAND4_X1  g755(.A1(new_n944), .A2(new_n318), .A3(new_n651), .A4(new_n946), .ZN(new_n957));
  NAND2_X1  g756(.A1(new_n956), .A2(new_n957), .ZN(new_n958));
  NAND2_X1  g757(.A1(new_n958), .A2(KEYINPUT60), .ZN(new_n959));
  INV_X1    g758(.A(KEYINPUT60), .ZN(new_n960));
  NAND3_X1  g759(.A1(new_n956), .A2(new_n960), .A3(new_n957), .ZN(new_n961));
  NAND2_X1  g760(.A1(new_n959), .A2(new_n961), .ZN(G1350gat));
  NAND4_X1  g761(.A1(new_n944), .A2(new_n317), .A3(new_n700), .A4(new_n946), .ZN(new_n963));
  INV_X1    g762(.A(KEYINPUT125), .ZN(new_n964));
  NAND4_X1  g763(.A1(new_n845), .A2(new_n941), .A3(new_n736), .A4(new_n700), .ZN(new_n965));
  INV_X1    g764(.A(KEYINPUT61), .ZN(new_n966));
  AND4_X1   g765(.A1(new_n964), .A2(new_n965), .A3(new_n966), .A4(G190gat), .ZN(new_n967));
  AOI21_X1  g766(.A(new_n333), .B1(KEYINPUT125), .B2(KEYINPUT61), .ZN(new_n968));
  AOI22_X1  g767(.A1(new_n965), .A2(new_n968), .B1(new_n964), .B2(new_n966), .ZN(new_n969));
  OAI21_X1  g768(.A(new_n963), .B1(new_n967), .B2(new_n969), .ZN(new_n970));
  NAND2_X1  g769(.A1(new_n970), .A2(KEYINPUT126), .ZN(new_n971));
  INV_X1    g770(.A(KEYINPUT126), .ZN(new_n972));
  OAI211_X1 g771(.A(new_n972), .B(new_n963), .C1(new_n967), .C2(new_n969), .ZN(new_n973));
  NAND2_X1  g772(.A1(new_n971), .A2(new_n973), .ZN(G1351gat));
  NOR2_X1   g773(.A1(new_n896), .A2(new_n719), .ZN(new_n975));
  NAND2_X1  g774(.A1(new_n944), .A2(new_n975), .ZN(new_n976));
  INV_X1    g775(.A(new_n976), .ZN(new_n977));
  AOI21_X1  g776(.A(G197gat), .B1(new_n977), .B2(new_n744), .ZN(new_n978));
  NOR3_X1   g777(.A1(new_n750), .A2(new_n719), .A3(new_n759), .ZN(new_n979));
  INV_X1    g778(.A(new_n979), .ZN(new_n980));
  NOR2_X1   g779(.A1(new_n920), .A2(new_n980), .ZN(new_n981));
  AND2_X1   g780(.A1(new_n744), .A2(G197gat), .ZN(new_n982));
  AOI21_X1  g781(.A(new_n978), .B1(new_n981), .B2(new_n982), .ZN(G1352gat));
  INV_X1    g782(.A(G204gat), .ZN(new_n984));
  NAND2_X1  g783(.A1(new_n675), .A2(new_n984), .ZN(new_n985));
  OR3_X1    g784(.A1(new_n976), .A2(KEYINPUT62), .A3(new_n985), .ZN(new_n986));
  OAI21_X1  g785(.A(KEYINPUT62), .B1(new_n976), .B2(new_n985), .ZN(new_n987));
  NOR3_X1   g786(.A1(new_n920), .A2(new_n745), .A3(new_n980), .ZN(new_n988));
  OAI211_X1 g787(.A(new_n986), .B(new_n987), .C1(new_n988), .C2(new_n984), .ZN(G1353gat));
  OR3_X1    g788(.A1(new_n976), .A2(G211gat), .A3(new_n650), .ZN(new_n990));
  NAND2_X1  g789(.A1(new_n911), .A2(new_n916), .ZN(new_n991));
  NAND3_X1  g790(.A1(new_n991), .A2(new_n651), .A3(new_n979), .ZN(new_n992));
  AND3_X1   g791(.A1(new_n992), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n993));
  AOI21_X1  g792(.A(KEYINPUT63), .B1(new_n992), .B2(G211gat), .ZN(new_n994));
  OAI21_X1  g793(.A(new_n990), .B1(new_n993), .B2(new_n994), .ZN(G1354gat));
  INV_X1    g794(.A(G218gat), .ZN(new_n996));
  NAND3_X1  g795(.A1(new_n977), .A2(new_n996), .A3(new_n700), .ZN(new_n997));
  INV_X1    g796(.A(KEYINPUT127), .ZN(new_n998));
  OAI21_X1  g797(.A(new_n998), .B1(new_n920), .B2(new_n980), .ZN(new_n999));
  NAND3_X1  g798(.A1(new_n991), .A2(KEYINPUT127), .A3(new_n979), .ZN(new_n1000));
  AND3_X1   g799(.A1(new_n999), .A2(new_n1000), .A3(new_n700), .ZN(new_n1001));
  OAI21_X1  g800(.A(new_n997), .B1(new_n1001), .B2(new_n996), .ZN(G1355gat));
endmodule


